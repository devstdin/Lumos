magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< nwell >>
rect -650 -650 650 650
<< psubdiff >>
rect -758 744 758 758
rect -758 712 -684 744
rect 684 712 758 744
rect -758 698 758 712
rect -758 684 -698 698
rect -758 -684 -744 684
rect -712 -684 -698 684
rect 698 684 758 698
rect -758 -698 -698 -684
rect 698 -684 712 684
rect 744 -684 758 684
rect 698 -698 758 -684
rect -758 -712 758 -698
rect -758 -744 -684 -712
rect 684 -744 758 -712
rect -758 -758 758 -744
<< nsubdiff >>
rect -602 588 602 602
rect -602 556 -528 588
rect 528 556 602 588
rect -602 542 602 556
rect -602 528 -542 542
rect -602 -528 -588 528
rect -556 -528 -542 528
rect 542 528 602 542
rect -602 -542 -542 -528
rect 542 -528 556 528
rect 588 -528 602 528
rect 542 -542 602 -528
rect -602 -556 602 -542
rect -602 -588 -528 -556
rect 528 -588 602 -556
rect -602 -602 602 -588
<< psubdiffcont >>
rect -684 712 684 744
rect -744 -684 -712 684
rect 712 -684 744 684
rect -684 -744 684 -712
<< nsubdiffcont >>
rect -528 556 528 588
rect -588 -528 -556 528
rect 556 -528 588 528
rect -528 -588 528 -556
<< pdiode >>
rect -500 461 500 500
rect -500 -462 -462 461
rect 461 -462 500 461
rect -500 -500 500 -462
<< pdiodecont >>
rect -462 -462 461 461
<< metal1 >>
rect -754 744 754 754
rect -754 712 -684 744
rect 684 712 754 744
rect -754 702 754 712
rect -754 684 -702 702
rect -754 -684 -744 684
rect -712 -684 -702 684
rect 702 684 754 702
rect -598 588 598 598
rect -598 556 -528 588
rect 528 556 598 588
rect -598 546 598 556
rect -598 528 -546 546
rect -598 -528 -588 528
rect -556 -528 -546 528
rect 546 528 598 546
rect -598 -546 -546 -528
rect 546 -528 556 528
rect 588 -528 598 528
rect 546 -546 598 -528
rect -598 -556 598 -546
rect -598 -588 -528 -556
rect 528 -588 598 -556
rect -598 -598 598 -588
rect -754 -702 -702 -684
rect 702 -684 712 684
rect 744 -684 754 684
rect 702 -702 754 -684
rect -754 -712 754 -702
rect -754 -744 -684 -712
rect 684 -744 754 -712
rect -754 -754 754 -744
<< properties >>
string gencell dpantenna
string library sg13g2_devstdin
string parameters w 5 l 5 nx 1 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class diode contcov 95 glc 1 grc 1 gtc 1 gbc 1
<< end >>
