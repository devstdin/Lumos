magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752516157
<< nwell >>
rect 312 312 2558 7098
<< pwell >>
rect 58 7198 2806 7346
rect 58 212 206 7198
rect 2658 212 2806 7198
rect 58 64 2806 212
<< pdiff >>
rect 846 6466 1098 6486
rect 846 6434 888 6466
rect 920 6434 960 6466
rect 992 6434 1032 6466
rect 1064 6434 1098 6466
rect 846 6394 1098 6434
rect 846 6362 888 6394
rect 920 6362 960 6394
rect 992 6362 1032 6394
rect 1064 6362 1098 6394
rect 846 6322 1098 6362
rect 846 6290 888 6322
rect 920 6290 960 6322
rect 992 6290 1032 6322
rect 1064 6290 1098 6322
rect 846 6250 1098 6290
rect 846 6218 888 6250
rect 920 6218 960 6250
rect 992 6218 1032 6250
rect 1064 6218 1098 6250
rect 846 6178 1098 6218
rect 846 6146 888 6178
rect 920 6146 960 6178
rect 992 6146 1032 6178
rect 1064 6146 1098 6178
rect 846 6106 1098 6146
rect 846 6074 888 6106
rect 920 6074 960 6106
rect 992 6074 1032 6106
rect 1064 6074 1098 6106
rect 846 6034 1098 6074
rect 846 6002 888 6034
rect 920 6002 960 6034
rect 992 6002 1032 6034
rect 1064 6002 1098 6034
rect 846 5962 1098 6002
rect 846 5930 888 5962
rect 920 5930 960 5962
rect 992 5930 1032 5962
rect 1064 5930 1098 5962
rect 846 5890 1098 5930
rect 846 5858 888 5890
rect 920 5858 960 5890
rect 992 5858 1032 5890
rect 1064 5858 1098 5890
rect 846 5818 1098 5858
rect 846 5786 888 5818
rect 920 5786 960 5818
rect 992 5786 1032 5818
rect 1064 5786 1098 5818
rect 846 5746 1098 5786
rect 846 5714 888 5746
rect 920 5714 960 5746
rect 992 5714 1032 5746
rect 1064 5714 1098 5746
rect 846 5674 1098 5714
rect 846 5642 888 5674
rect 920 5642 960 5674
rect 992 5642 1032 5674
rect 1064 5642 1098 5674
rect 846 5602 1098 5642
rect 846 5570 888 5602
rect 920 5570 960 5602
rect 992 5570 1032 5602
rect 1064 5570 1098 5602
rect 846 5530 1098 5570
rect 846 5498 888 5530
rect 920 5498 960 5530
rect 992 5498 1032 5530
rect 1064 5498 1098 5530
rect 846 5458 1098 5498
rect 846 5426 888 5458
rect 920 5426 960 5458
rect 992 5426 1032 5458
rect 1064 5426 1098 5458
rect 846 5386 1098 5426
rect 846 5354 888 5386
rect 920 5354 960 5386
rect 992 5354 1032 5386
rect 1064 5354 1098 5386
rect 846 5314 1098 5354
rect 846 5282 888 5314
rect 920 5282 960 5314
rect 992 5282 1032 5314
rect 1064 5282 1098 5314
rect 846 5242 1098 5282
rect 846 5210 888 5242
rect 920 5210 960 5242
rect 992 5210 1032 5242
rect 1064 5210 1098 5242
rect 846 5170 1098 5210
rect 846 5138 888 5170
rect 920 5138 960 5170
rect 992 5138 1032 5170
rect 1064 5138 1098 5170
rect 846 5098 1098 5138
rect 846 5066 888 5098
rect 920 5066 960 5098
rect 992 5066 1032 5098
rect 1064 5066 1098 5098
rect 846 5026 1098 5066
rect 846 4994 888 5026
rect 920 4994 960 5026
rect 992 4994 1032 5026
rect 1064 4994 1098 5026
rect 846 4954 1098 4994
rect 846 4922 888 4954
rect 920 4922 960 4954
rect 992 4922 1032 4954
rect 1064 4922 1098 4954
rect 846 4882 1098 4922
rect 846 4850 888 4882
rect 920 4850 960 4882
rect 992 4850 1032 4882
rect 1064 4850 1098 4882
rect 846 4810 1098 4850
rect 846 4778 888 4810
rect 920 4778 960 4810
rect 992 4778 1032 4810
rect 1064 4778 1098 4810
rect 846 4738 1098 4778
rect 846 4706 888 4738
rect 920 4706 960 4738
rect 992 4706 1032 4738
rect 1064 4706 1098 4738
rect 846 4666 1098 4706
rect 846 4634 888 4666
rect 920 4634 960 4666
rect 992 4634 1032 4666
rect 1064 4634 1098 4666
rect 846 4594 1098 4634
rect 846 4562 888 4594
rect 920 4562 960 4594
rect 992 4562 1032 4594
rect 1064 4562 1098 4594
rect 846 4522 1098 4562
rect 846 4490 888 4522
rect 920 4490 960 4522
rect 992 4490 1032 4522
rect 1064 4490 1098 4522
rect 846 4450 1098 4490
rect 846 4418 888 4450
rect 920 4418 960 4450
rect 992 4418 1032 4450
rect 1064 4418 1098 4450
rect 846 4378 1098 4418
rect 846 4346 888 4378
rect 920 4346 960 4378
rect 992 4346 1032 4378
rect 1064 4346 1098 4378
rect 846 4306 1098 4346
rect 846 4274 888 4306
rect 920 4274 960 4306
rect 992 4274 1032 4306
rect 1064 4274 1098 4306
rect 846 4234 1098 4274
rect 846 4202 888 4234
rect 920 4202 960 4234
rect 992 4202 1032 4234
rect 1064 4202 1098 4234
rect 846 4162 1098 4202
rect 846 4130 888 4162
rect 920 4130 960 4162
rect 992 4130 1032 4162
rect 1064 4130 1098 4162
rect 846 4090 1098 4130
rect 846 4058 888 4090
rect 920 4058 960 4090
rect 992 4058 1032 4090
rect 1064 4058 1098 4090
rect 846 4018 1098 4058
rect 846 3986 888 4018
rect 920 3986 960 4018
rect 992 3986 1032 4018
rect 1064 3986 1098 4018
rect 846 3946 1098 3986
rect 846 3914 888 3946
rect 920 3914 960 3946
rect 992 3914 1032 3946
rect 1064 3914 1098 3946
rect 846 3874 1098 3914
rect 846 3842 888 3874
rect 920 3842 960 3874
rect 992 3842 1032 3874
rect 1064 3842 1098 3874
rect 846 3802 1098 3842
rect 846 3770 888 3802
rect 920 3770 960 3802
rect 992 3770 1032 3802
rect 1064 3770 1098 3802
rect 846 3730 1098 3770
rect 846 3698 888 3730
rect 920 3698 960 3730
rect 992 3698 1032 3730
rect 1064 3698 1098 3730
rect 846 3658 1098 3698
rect 846 3626 888 3658
rect 920 3626 960 3658
rect 992 3626 1032 3658
rect 1064 3626 1098 3658
rect 846 3586 1098 3626
rect 846 3554 888 3586
rect 920 3554 960 3586
rect 992 3554 1032 3586
rect 1064 3554 1098 3586
rect 846 3514 1098 3554
rect 846 3482 888 3514
rect 920 3482 960 3514
rect 992 3482 1032 3514
rect 1064 3482 1098 3514
rect 846 3442 1098 3482
rect 846 3410 888 3442
rect 920 3410 960 3442
rect 992 3410 1032 3442
rect 1064 3410 1098 3442
rect 846 3370 1098 3410
rect 846 3338 888 3370
rect 920 3338 960 3370
rect 992 3338 1032 3370
rect 1064 3338 1098 3370
rect 846 3298 1098 3338
rect 846 3266 888 3298
rect 920 3266 960 3298
rect 992 3266 1032 3298
rect 1064 3266 1098 3298
rect 846 3226 1098 3266
rect 846 3194 888 3226
rect 920 3194 960 3226
rect 992 3194 1032 3226
rect 1064 3194 1098 3226
rect 846 3154 1098 3194
rect 846 3122 888 3154
rect 920 3122 960 3154
rect 992 3122 1032 3154
rect 1064 3122 1098 3154
rect 846 3082 1098 3122
rect 846 3050 888 3082
rect 920 3050 960 3082
rect 992 3050 1032 3082
rect 1064 3050 1098 3082
rect 846 3010 1098 3050
rect 846 2978 888 3010
rect 920 2978 960 3010
rect 992 2978 1032 3010
rect 1064 2978 1098 3010
rect 846 2938 1098 2978
rect 846 2906 888 2938
rect 920 2906 960 2938
rect 992 2906 1032 2938
rect 1064 2906 1098 2938
rect 846 2866 1098 2906
rect 846 2834 888 2866
rect 920 2834 960 2866
rect 992 2834 1032 2866
rect 1064 2834 1098 2866
rect 846 2794 1098 2834
rect 846 2762 888 2794
rect 920 2762 960 2794
rect 992 2762 1032 2794
rect 1064 2762 1098 2794
rect 846 2722 1098 2762
rect 846 2690 888 2722
rect 920 2690 960 2722
rect 992 2690 1032 2722
rect 1064 2690 1098 2722
rect 846 2650 1098 2690
rect 846 2618 888 2650
rect 920 2618 960 2650
rect 992 2618 1032 2650
rect 1064 2618 1098 2650
rect 846 2578 1098 2618
rect 846 2546 888 2578
rect 920 2546 960 2578
rect 992 2546 1032 2578
rect 1064 2546 1098 2578
rect 846 2506 1098 2546
rect 846 2474 888 2506
rect 920 2474 960 2506
rect 992 2474 1032 2506
rect 1064 2474 1098 2506
rect 846 2434 1098 2474
rect 846 2402 888 2434
rect 920 2402 960 2434
rect 992 2402 1032 2434
rect 1064 2402 1098 2434
rect 846 2362 1098 2402
rect 846 2330 888 2362
rect 920 2330 960 2362
rect 992 2330 1032 2362
rect 1064 2330 1098 2362
rect 846 2290 1098 2330
rect 846 2258 888 2290
rect 920 2258 960 2290
rect 992 2258 1032 2290
rect 1064 2258 1098 2290
rect 846 2218 1098 2258
rect 846 2186 888 2218
rect 920 2186 960 2218
rect 992 2186 1032 2218
rect 1064 2186 1098 2218
rect 846 2146 1098 2186
rect 846 2114 888 2146
rect 920 2114 960 2146
rect 992 2114 1032 2146
rect 1064 2114 1098 2146
rect 846 2074 1098 2114
rect 846 2042 888 2074
rect 920 2042 960 2074
rect 992 2042 1032 2074
rect 1064 2042 1098 2074
rect 846 2002 1098 2042
rect 846 1970 888 2002
rect 920 1970 960 2002
rect 992 1970 1032 2002
rect 1064 1970 1098 2002
rect 846 1930 1098 1970
rect 846 1898 888 1930
rect 920 1898 960 1930
rect 992 1898 1032 1930
rect 1064 1898 1098 1930
rect 846 1858 1098 1898
rect 846 1826 888 1858
rect 920 1826 960 1858
rect 992 1826 1032 1858
rect 1064 1826 1098 1858
rect 846 1786 1098 1826
rect 846 1754 888 1786
rect 920 1754 960 1786
rect 992 1754 1032 1786
rect 1064 1754 1098 1786
rect 846 1714 1098 1754
rect 846 1682 888 1714
rect 920 1682 960 1714
rect 992 1682 1032 1714
rect 1064 1682 1098 1714
rect 846 1642 1098 1682
rect 846 1610 888 1642
rect 920 1610 960 1642
rect 992 1610 1032 1642
rect 1064 1610 1098 1642
rect 846 1570 1098 1610
rect 846 1538 888 1570
rect 920 1538 960 1570
rect 992 1538 1032 1570
rect 1064 1538 1098 1570
rect 846 1498 1098 1538
rect 846 1466 888 1498
rect 920 1466 960 1498
rect 992 1466 1032 1498
rect 1064 1466 1098 1498
rect 846 1426 1098 1466
rect 846 1394 888 1426
rect 920 1394 960 1426
rect 992 1394 1032 1426
rect 1064 1394 1098 1426
rect 846 1354 1098 1394
rect 846 1322 888 1354
rect 920 1322 960 1354
rect 992 1322 1032 1354
rect 1064 1322 1098 1354
rect 846 1282 1098 1322
rect 846 1250 888 1282
rect 920 1250 960 1282
rect 992 1250 1032 1282
rect 1064 1250 1098 1282
rect 846 1210 1098 1250
rect 846 1178 888 1210
rect 920 1178 960 1210
rect 992 1178 1032 1210
rect 1064 1178 1098 1210
rect 846 1138 1098 1178
rect 846 1106 888 1138
rect 920 1106 960 1138
rect 992 1106 1032 1138
rect 1064 1106 1098 1138
rect 846 1066 1098 1106
rect 846 1034 888 1066
rect 920 1034 960 1066
rect 992 1034 1032 1066
rect 1064 1034 1098 1066
rect 846 994 1098 1034
rect 846 962 888 994
rect 920 962 960 994
rect 992 962 1032 994
rect 1064 962 1098 994
rect 846 930 1098 962
rect 1752 6466 2004 6486
rect 1752 6434 1794 6466
rect 1826 6434 1866 6466
rect 1898 6434 1938 6466
rect 1970 6434 2004 6466
rect 1752 6394 2004 6434
rect 1752 6362 1794 6394
rect 1826 6362 1866 6394
rect 1898 6362 1938 6394
rect 1970 6362 2004 6394
rect 1752 6322 2004 6362
rect 1752 6290 1794 6322
rect 1826 6290 1866 6322
rect 1898 6290 1938 6322
rect 1970 6290 2004 6322
rect 1752 6250 2004 6290
rect 1752 6218 1794 6250
rect 1826 6218 1866 6250
rect 1898 6218 1938 6250
rect 1970 6218 2004 6250
rect 1752 6178 2004 6218
rect 1752 6146 1794 6178
rect 1826 6146 1866 6178
rect 1898 6146 1938 6178
rect 1970 6146 2004 6178
rect 1752 6106 2004 6146
rect 1752 6074 1794 6106
rect 1826 6074 1866 6106
rect 1898 6074 1938 6106
rect 1970 6074 2004 6106
rect 1752 6034 2004 6074
rect 1752 6002 1794 6034
rect 1826 6002 1866 6034
rect 1898 6002 1938 6034
rect 1970 6002 2004 6034
rect 1752 5962 2004 6002
rect 1752 5930 1794 5962
rect 1826 5930 1866 5962
rect 1898 5930 1938 5962
rect 1970 5930 2004 5962
rect 1752 5890 2004 5930
rect 1752 5858 1794 5890
rect 1826 5858 1866 5890
rect 1898 5858 1938 5890
rect 1970 5858 2004 5890
rect 1752 5818 2004 5858
rect 1752 5786 1794 5818
rect 1826 5786 1866 5818
rect 1898 5786 1938 5818
rect 1970 5786 2004 5818
rect 1752 5746 2004 5786
rect 1752 5714 1794 5746
rect 1826 5714 1866 5746
rect 1898 5714 1938 5746
rect 1970 5714 2004 5746
rect 1752 5674 2004 5714
rect 1752 5642 1794 5674
rect 1826 5642 1866 5674
rect 1898 5642 1938 5674
rect 1970 5642 2004 5674
rect 1752 5602 2004 5642
rect 1752 5570 1794 5602
rect 1826 5570 1866 5602
rect 1898 5570 1938 5602
rect 1970 5570 2004 5602
rect 1752 5530 2004 5570
rect 1752 5498 1794 5530
rect 1826 5498 1866 5530
rect 1898 5498 1938 5530
rect 1970 5498 2004 5530
rect 1752 5458 2004 5498
rect 1752 5426 1794 5458
rect 1826 5426 1866 5458
rect 1898 5426 1938 5458
rect 1970 5426 2004 5458
rect 1752 5386 2004 5426
rect 1752 5354 1794 5386
rect 1826 5354 1866 5386
rect 1898 5354 1938 5386
rect 1970 5354 2004 5386
rect 1752 5314 2004 5354
rect 1752 5282 1794 5314
rect 1826 5282 1866 5314
rect 1898 5282 1938 5314
rect 1970 5282 2004 5314
rect 1752 5242 2004 5282
rect 1752 5210 1794 5242
rect 1826 5210 1866 5242
rect 1898 5210 1938 5242
rect 1970 5210 2004 5242
rect 1752 5170 2004 5210
rect 1752 5138 1794 5170
rect 1826 5138 1866 5170
rect 1898 5138 1938 5170
rect 1970 5138 2004 5170
rect 1752 5098 2004 5138
rect 1752 5066 1794 5098
rect 1826 5066 1866 5098
rect 1898 5066 1938 5098
rect 1970 5066 2004 5098
rect 1752 5026 2004 5066
rect 1752 4994 1794 5026
rect 1826 4994 1866 5026
rect 1898 4994 1938 5026
rect 1970 4994 2004 5026
rect 1752 4954 2004 4994
rect 1752 4922 1794 4954
rect 1826 4922 1866 4954
rect 1898 4922 1938 4954
rect 1970 4922 2004 4954
rect 1752 4882 2004 4922
rect 1752 4850 1794 4882
rect 1826 4850 1866 4882
rect 1898 4850 1938 4882
rect 1970 4850 2004 4882
rect 1752 4810 2004 4850
rect 1752 4778 1794 4810
rect 1826 4778 1866 4810
rect 1898 4778 1938 4810
rect 1970 4778 2004 4810
rect 1752 4738 2004 4778
rect 1752 4706 1794 4738
rect 1826 4706 1866 4738
rect 1898 4706 1938 4738
rect 1970 4706 2004 4738
rect 1752 4666 2004 4706
rect 1752 4634 1794 4666
rect 1826 4634 1866 4666
rect 1898 4634 1938 4666
rect 1970 4634 2004 4666
rect 1752 4594 2004 4634
rect 1752 4562 1794 4594
rect 1826 4562 1866 4594
rect 1898 4562 1938 4594
rect 1970 4562 2004 4594
rect 1752 4522 2004 4562
rect 1752 4490 1794 4522
rect 1826 4490 1866 4522
rect 1898 4490 1938 4522
rect 1970 4490 2004 4522
rect 1752 4450 2004 4490
rect 1752 4418 1794 4450
rect 1826 4418 1866 4450
rect 1898 4418 1938 4450
rect 1970 4418 2004 4450
rect 1752 4378 2004 4418
rect 1752 4346 1794 4378
rect 1826 4346 1866 4378
rect 1898 4346 1938 4378
rect 1970 4346 2004 4378
rect 1752 4306 2004 4346
rect 1752 4274 1794 4306
rect 1826 4274 1866 4306
rect 1898 4274 1938 4306
rect 1970 4274 2004 4306
rect 1752 4234 2004 4274
rect 1752 4202 1794 4234
rect 1826 4202 1866 4234
rect 1898 4202 1938 4234
rect 1970 4202 2004 4234
rect 1752 4162 2004 4202
rect 1752 4130 1794 4162
rect 1826 4130 1866 4162
rect 1898 4130 1938 4162
rect 1970 4130 2004 4162
rect 1752 4090 2004 4130
rect 1752 4058 1794 4090
rect 1826 4058 1866 4090
rect 1898 4058 1938 4090
rect 1970 4058 2004 4090
rect 1752 4018 2004 4058
rect 1752 3986 1794 4018
rect 1826 3986 1866 4018
rect 1898 3986 1938 4018
rect 1970 3986 2004 4018
rect 1752 3946 2004 3986
rect 1752 3914 1794 3946
rect 1826 3914 1866 3946
rect 1898 3914 1938 3946
rect 1970 3914 2004 3946
rect 1752 3874 2004 3914
rect 1752 3842 1794 3874
rect 1826 3842 1866 3874
rect 1898 3842 1938 3874
rect 1970 3842 2004 3874
rect 1752 3802 2004 3842
rect 1752 3770 1794 3802
rect 1826 3770 1866 3802
rect 1898 3770 1938 3802
rect 1970 3770 2004 3802
rect 1752 3730 2004 3770
rect 1752 3698 1794 3730
rect 1826 3698 1866 3730
rect 1898 3698 1938 3730
rect 1970 3698 2004 3730
rect 1752 3658 2004 3698
rect 1752 3626 1794 3658
rect 1826 3626 1866 3658
rect 1898 3626 1938 3658
rect 1970 3626 2004 3658
rect 1752 3586 2004 3626
rect 1752 3554 1794 3586
rect 1826 3554 1866 3586
rect 1898 3554 1938 3586
rect 1970 3554 2004 3586
rect 1752 3514 2004 3554
rect 1752 3482 1794 3514
rect 1826 3482 1866 3514
rect 1898 3482 1938 3514
rect 1970 3482 2004 3514
rect 1752 3442 2004 3482
rect 1752 3410 1794 3442
rect 1826 3410 1866 3442
rect 1898 3410 1938 3442
rect 1970 3410 2004 3442
rect 1752 3370 2004 3410
rect 1752 3338 1794 3370
rect 1826 3338 1866 3370
rect 1898 3338 1938 3370
rect 1970 3338 2004 3370
rect 1752 3298 2004 3338
rect 1752 3266 1794 3298
rect 1826 3266 1866 3298
rect 1898 3266 1938 3298
rect 1970 3266 2004 3298
rect 1752 3226 2004 3266
rect 1752 3194 1794 3226
rect 1826 3194 1866 3226
rect 1898 3194 1938 3226
rect 1970 3194 2004 3226
rect 1752 3154 2004 3194
rect 1752 3122 1794 3154
rect 1826 3122 1866 3154
rect 1898 3122 1938 3154
rect 1970 3122 2004 3154
rect 1752 3082 2004 3122
rect 1752 3050 1794 3082
rect 1826 3050 1866 3082
rect 1898 3050 1938 3082
rect 1970 3050 2004 3082
rect 1752 3010 2004 3050
rect 1752 2978 1794 3010
rect 1826 2978 1866 3010
rect 1898 2978 1938 3010
rect 1970 2978 2004 3010
rect 1752 2938 2004 2978
rect 1752 2906 1794 2938
rect 1826 2906 1866 2938
rect 1898 2906 1938 2938
rect 1970 2906 2004 2938
rect 1752 2866 2004 2906
rect 1752 2834 1794 2866
rect 1826 2834 1866 2866
rect 1898 2834 1938 2866
rect 1970 2834 2004 2866
rect 1752 2794 2004 2834
rect 1752 2762 1794 2794
rect 1826 2762 1866 2794
rect 1898 2762 1938 2794
rect 1970 2762 2004 2794
rect 1752 2722 2004 2762
rect 1752 2690 1794 2722
rect 1826 2690 1866 2722
rect 1898 2690 1938 2722
rect 1970 2690 2004 2722
rect 1752 2650 2004 2690
rect 1752 2618 1794 2650
rect 1826 2618 1866 2650
rect 1898 2618 1938 2650
rect 1970 2618 2004 2650
rect 1752 2578 2004 2618
rect 1752 2546 1794 2578
rect 1826 2546 1866 2578
rect 1898 2546 1938 2578
rect 1970 2546 2004 2578
rect 1752 2506 2004 2546
rect 1752 2474 1794 2506
rect 1826 2474 1866 2506
rect 1898 2474 1938 2506
rect 1970 2474 2004 2506
rect 1752 2434 2004 2474
rect 1752 2402 1794 2434
rect 1826 2402 1866 2434
rect 1898 2402 1938 2434
rect 1970 2402 2004 2434
rect 1752 2362 2004 2402
rect 1752 2330 1794 2362
rect 1826 2330 1866 2362
rect 1898 2330 1938 2362
rect 1970 2330 2004 2362
rect 1752 2290 2004 2330
rect 1752 2258 1794 2290
rect 1826 2258 1866 2290
rect 1898 2258 1938 2290
rect 1970 2258 2004 2290
rect 1752 2218 2004 2258
rect 1752 2186 1794 2218
rect 1826 2186 1866 2218
rect 1898 2186 1938 2218
rect 1970 2186 2004 2218
rect 1752 2146 2004 2186
rect 1752 2114 1794 2146
rect 1826 2114 1866 2146
rect 1898 2114 1938 2146
rect 1970 2114 2004 2146
rect 1752 2074 2004 2114
rect 1752 2042 1794 2074
rect 1826 2042 1866 2074
rect 1898 2042 1938 2074
rect 1970 2042 2004 2074
rect 1752 2002 2004 2042
rect 1752 1970 1794 2002
rect 1826 1970 1866 2002
rect 1898 1970 1938 2002
rect 1970 1970 2004 2002
rect 1752 1930 2004 1970
rect 1752 1898 1794 1930
rect 1826 1898 1866 1930
rect 1898 1898 1938 1930
rect 1970 1898 2004 1930
rect 1752 1858 2004 1898
rect 1752 1826 1794 1858
rect 1826 1826 1866 1858
rect 1898 1826 1938 1858
rect 1970 1826 2004 1858
rect 1752 1786 2004 1826
rect 1752 1754 1794 1786
rect 1826 1754 1866 1786
rect 1898 1754 1938 1786
rect 1970 1754 2004 1786
rect 1752 1714 2004 1754
rect 1752 1682 1794 1714
rect 1826 1682 1866 1714
rect 1898 1682 1938 1714
rect 1970 1682 2004 1714
rect 1752 1642 2004 1682
rect 1752 1610 1794 1642
rect 1826 1610 1866 1642
rect 1898 1610 1938 1642
rect 1970 1610 2004 1642
rect 1752 1570 2004 1610
rect 1752 1538 1794 1570
rect 1826 1538 1866 1570
rect 1898 1538 1938 1570
rect 1970 1538 2004 1570
rect 1752 1498 2004 1538
rect 1752 1466 1794 1498
rect 1826 1466 1866 1498
rect 1898 1466 1938 1498
rect 1970 1466 2004 1498
rect 1752 1426 2004 1466
rect 1752 1394 1794 1426
rect 1826 1394 1866 1426
rect 1898 1394 1938 1426
rect 1970 1394 2004 1426
rect 1752 1354 2004 1394
rect 1752 1322 1794 1354
rect 1826 1322 1866 1354
rect 1898 1322 1938 1354
rect 1970 1322 2004 1354
rect 1752 1282 2004 1322
rect 1752 1250 1794 1282
rect 1826 1250 1866 1282
rect 1898 1250 1938 1282
rect 1970 1250 2004 1282
rect 1752 1210 2004 1250
rect 1752 1178 1794 1210
rect 1826 1178 1866 1210
rect 1898 1178 1938 1210
rect 1970 1178 2004 1210
rect 1752 1138 2004 1178
rect 1752 1106 1794 1138
rect 1826 1106 1866 1138
rect 1898 1106 1938 1138
rect 1970 1106 2004 1138
rect 1752 1066 2004 1106
rect 1752 1034 1794 1066
rect 1826 1034 1866 1066
rect 1898 1034 1938 1066
rect 1970 1034 2004 1066
rect 1752 994 2004 1034
rect 1752 962 1794 994
rect 1826 962 1866 994
rect 1898 962 1938 994
rect 1970 962 2004 994
rect 1752 930 2004 962
<< pdiffc >>
rect 888 6434 920 6466
rect 960 6434 992 6466
rect 1032 6434 1064 6466
rect 888 6362 920 6394
rect 960 6362 992 6394
rect 1032 6362 1064 6394
rect 888 6290 920 6322
rect 960 6290 992 6322
rect 1032 6290 1064 6322
rect 888 6218 920 6250
rect 960 6218 992 6250
rect 1032 6218 1064 6250
rect 888 6146 920 6178
rect 960 6146 992 6178
rect 1032 6146 1064 6178
rect 888 6074 920 6106
rect 960 6074 992 6106
rect 1032 6074 1064 6106
rect 888 6002 920 6034
rect 960 6002 992 6034
rect 1032 6002 1064 6034
rect 888 5930 920 5962
rect 960 5930 992 5962
rect 1032 5930 1064 5962
rect 888 5858 920 5890
rect 960 5858 992 5890
rect 1032 5858 1064 5890
rect 888 5786 920 5818
rect 960 5786 992 5818
rect 1032 5786 1064 5818
rect 888 5714 920 5746
rect 960 5714 992 5746
rect 1032 5714 1064 5746
rect 888 5642 920 5674
rect 960 5642 992 5674
rect 1032 5642 1064 5674
rect 888 5570 920 5602
rect 960 5570 992 5602
rect 1032 5570 1064 5602
rect 888 5498 920 5530
rect 960 5498 992 5530
rect 1032 5498 1064 5530
rect 888 5426 920 5458
rect 960 5426 992 5458
rect 1032 5426 1064 5458
rect 888 5354 920 5386
rect 960 5354 992 5386
rect 1032 5354 1064 5386
rect 888 5282 920 5314
rect 960 5282 992 5314
rect 1032 5282 1064 5314
rect 888 5210 920 5242
rect 960 5210 992 5242
rect 1032 5210 1064 5242
rect 888 5138 920 5170
rect 960 5138 992 5170
rect 1032 5138 1064 5170
rect 888 5066 920 5098
rect 960 5066 992 5098
rect 1032 5066 1064 5098
rect 888 4994 920 5026
rect 960 4994 992 5026
rect 1032 4994 1064 5026
rect 888 4922 920 4954
rect 960 4922 992 4954
rect 1032 4922 1064 4954
rect 888 4850 920 4882
rect 960 4850 992 4882
rect 1032 4850 1064 4882
rect 888 4778 920 4810
rect 960 4778 992 4810
rect 1032 4778 1064 4810
rect 888 4706 920 4738
rect 960 4706 992 4738
rect 1032 4706 1064 4738
rect 888 4634 920 4666
rect 960 4634 992 4666
rect 1032 4634 1064 4666
rect 888 4562 920 4594
rect 960 4562 992 4594
rect 1032 4562 1064 4594
rect 888 4490 920 4522
rect 960 4490 992 4522
rect 1032 4490 1064 4522
rect 888 4418 920 4450
rect 960 4418 992 4450
rect 1032 4418 1064 4450
rect 888 4346 920 4378
rect 960 4346 992 4378
rect 1032 4346 1064 4378
rect 888 4274 920 4306
rect 960 4274 992 4306
rect 1032 4274 1064 4306
rect 888 4202 920 4234
rect 960 4202 992 4234
rect 1032 4202 1064 4234
rect 888 4130 920 4162
rect 960 4130 992 4162
rect 1032 4130 1064 4162
rect 888 4058 920 4090
rect 960 4058 992 4090
rect 1032 4058 1064 4090
rect 888 3986 920 4018
rect 960 3986 992 4018
rect 1032 3986 1064 4018
rect 888 3914 920 3946
rect 960 3914 992 3946
rect 1032 3914 1064 3946
rect 888 3842 920 3874
rect 960 3842 992 3874
rect 1032 3842 1064 3874
rect 888 3770 920 3802
rect 960 3770 992 3802
rect 1032 3770 1064 3802
rect 888 3698 920 3730
rect 960 3698 992 3730
rect 1032 3698 1064 3730
rect 888 3626 920 3658
rect 960 3626 992 3658
rect 1032 3626 1064 3658
rect 888 3554 920 3586
rect 960 3554 992 3586
rect 1032 3554 1064 3586
rect 888 3482 920 3514
rect 960 3482 992 3514
rect 1032 3482 1064 3514
rect 888 3410 920 3442
rect 960 3410 992 3442
rect 1032 3410 1064 3442
rect 888 3338 920 3370
rect 960 3338 992 3370
rect 1032 3338 1064 3370
rect 888 3266 920 3298
rect 960 3266 992 3298
rect 1032 3266 1064 3298
rect 888 3194 920 3226
rect 960 3194 992 3226
rect 1032 3194 1064 3226
rect 888 3122 920 3154
rect 960 3122 992 3154
rect 1032 3122 1064 3154
rect 888 3050 920 3082
rect 960 3050 992 3082
rect 1032 3050 1064 3082
rect 888 2978 920 3010
rect 960 2978 992 3010
rect 1032 2978 1064 3010
rect 888 2906 920 2938
rect 960 2906 992 2938
rect 1032 2906 1064 2938
rect 888 2834 920 2866
rect 960 2834 992 2866
rect 1032 2834 1064 2866
rect 888 2762 920 2794
rect 960 2762 992 2794
rect 1032 2762 1064 2794
rect 888 2690 920 2722
rect 960 2690 992 2722
rect 1032 2690 1064 2722
rect 888 2618 920 2650
rect 960 2618 992 2650
rect 1032 2618 1064 2650
rect 888 2546 920 2578
rect 960 2546 992 2578
rect 1032 2546 1064 2578
rect 888 2474 920 2506
rect 960 2474 992 2506
rect 1032 2474 1064 2506
rect 888 2402 920 2434
rect 960 2402 992 2434
rect 1032 2402 1064 2434
rect 888 2330 920 2362
rect 960 2330 992 2362
rect 1032 2330 1064 2362
rect 888 2258 920 2290
rect 960 2258 992 2290
rect 1032 2258 1064 2290
rect 888 2186 920 2218
rect 960 2186 992 2218
rect 1032 2186 1064 2218
rect 888 2114 920 2146
rect 960 2114 992 2146
rect 1032 2114 1064 2146
rect 888 2042 920 2074
rect 960 2042 992 2074
rect 1032 2042 1064 2074
rect 888 1970 920 2002
rect 960 1970 992 2002
rect 1032 1970 1064 2002
rect 888 1898 920 1930
rect 960 1898 992 1930
rect 1032 1898 1064 1930
rect 888 1826 920 1858
rect 960 1826 992 1858
rect 1032 1826 1064 1858
rect 888 1754 920 1786
rect 960 1754 992 1786
rect 1032 1754 1064 1786
rect 888 1682 920 1714
rect 960 1682 992 1714
rect 1032 1682 1064 1714
rect 888 1610 920 1642
rect 960 1610 992 1642
rect 1032 1610 1064 1642
rect 888 1538 920 1570
rect 960 1538 992 1570
rect 1032 1538 1064 1570
rect 888 1466 920 1498
rect 960 1466 992 1498
rect 1032 1466 1064 1498
rect 888 1394 920 1426
rect 960 1394 992 1426
rect 1032 1394 1064 1426
rect 888 1322 920 1354
rect 960 1322 992 1354
rect 1032 1322 1064 1354
rect 888 1250 920 1282
rect 960 1250 992 1282
rect 1032 1250 1064 1282
rect 888 1178 920 1210
rect 960 1178 992 1210
rect 1032 1178 1064 1210
rect 888 1106 920 1138
rect 960 1106 992 1138
rect 1032 1106 1064 1138
rect 888 1034 920 1066
rect 960 1034 992 1066
rect 1032 1034 1064 1066
rect 888 962 920 994
rect 960 962 992 994
rect 1032 962 1064 994
rect 1794 6434 1826 6466
rect 1866 6434 1898 6466
rect 1938 6434 1970 6466
rect 1794 6362 1826 6394
rect 1866 6362 1898 6394
rect 1938 6362 1970 6394
rect 1794 6290 1826 6322
rect 1866 6290 1898 6322
rect 1938 6290 1970 6322
rect 1794 6218 1826 6250
rect 1866 6218 1898 6250
rect 1938 6218 1970 6250
rect 1794 6146 1826 6178
rect 1866 6146 1898 6178
rect 1938 6146 1970 6178
rect 1794 6074 1826 6106
rect 1866 6074 1898 6106
rect 1938 6074 1970 6106
rect 1794 6002 1826 6034
rect 1866 6002 1898 6034
rect 1938 6002 1970 6034
rect 1794 5930 1826 5962
rect 1866 5930 1898 5962
rect 1938 5930 1970 5962
rect 1794 5858 1826 5890
rect 1866 5858 1898 5890
rect 1938 5858 1970 5890
rect 1794 5786 1826 5818
rect 1866 5786 1898 5818
rect 1938 5786 1970 5818
rect 1794 5714 1826 5746
rect 1866 5714 1898 5746
rect 1938 5714 1970 5746
rect 1794 5642 1826 5674
rect 1866 5642 1898 5674
rect 1938 5642 1970 5674
rect 1794 5570 1826 5602
rect 1866 5570 1898 5602
rect 1938 5570 1970 5602
rect 1794 5498 1826 5530
rect 1866 5498 1898 5530
rect 1938 5498 1970 5530
rect 1794 5426 1826 5458
rect 1866 5426 1898 5458
rect 1938 5426 1970 5458
rect 1794 5354 1826 5386
rect 1866 5354 1898 5386
rect 1938 5354 1970 5386
rect 1794 5282 1826 5314
rect 1866 5282 1898 5314
rect 1938 5282 1970 5314
rect 1794 5210 1826 5242
rect 1866 5210 1898 5242
rect 1938 5210 1970 5242
rect 1794 5138 1826 5170
rect 1866 5138 1898 5170
rect 1938 5138 1970 5170
rect 1794 5066 1826 5098
rect 1866 5066 1898 5098
rect 1938 5066 1970 5098
rect 1794 4994 1826 5026
rect 1866 4994 1898 5026
rect 1938 4994 1970 5026
rect 1794 4922 1826 4954
rect 1866 4922 1898 4954
rect 1938 4922 1970 4954
rect 1794 4850 1826 4882
rect 1866 4850 1898 4882
rect 1938 4850 1970 4882
rect 1794 4778 1826 4810
rect 1866 4778 1898 4810
rect 1938 4778 1970 4810
rect 1794 4706 1826 4738
rect 1866 4706 1898 4738
rect 1938 4706 1970 4738
rect 1794 4634 1826 4666
rect 1866 4634 1898 4666
rect 1938 4634 1970 4666
rect 1794 4562 1826 4594
rect 1866 4562 1898 4594
rect 1938 4562 1970 4594
rect 1794 4490 1826 4522
rect 1866 4490 1898 4522
rect 1938 4490 1970 4522
rect 1794 4418 1826 4450
rect 1866 4418 1898 4450
rect 1938 4418 1970 4450
rect 1794 4346 1826 4378
rect 1866 4346 1898 4378
rect 1938 4346 1970 4378
rect 1794 4274 1826 4306
rect 1866 4274 1898 4306
rect 1938 4274 1970 4306
rect 1794 4202 1826 4234
rect 1866 4202 1898 4234
rect 1938 4202 1970 4234
rect 1794 4130 1826 4162
rect 1866 4130 1898 4162
rect 1938 4130 1970 4162
rect 1794 4058 1826 4090
rect 1866 4058 1898 4090
rect 1938 4058 1970 4090
rect 1794 3986 1826 4018
rect 1866 3986 1898 4018
rect 1938 3986 1970 4018
rect 1794 3914 1826 3946
rect 1866 3914 1898 3946
rect 1938 3914 1970 3946
rect 1794 3842 1826 3874
rect 1866 3842 1898 3874
rect 1938 3842 1970 3874
rect 1794 3770 1826 3802
rect 1866 3770 1898 3802
rect 1938 3770 1970 3802
rect 1794 3698 1826 3730
rect 1866 3698 1898 3730
rect 1938 3698 1970 3730
rect 1794 3626 1826 3658
rect 1866 3626 1898 3658
rect 1938 3626 1970 3658
rect 1794 3554 1826 3586
rect 1866 3554 1898 3586
rect 1938 3554 1970 3586
rect 1794 3482 1826 3514
rect 1866 3482 1898 3514
rect 1938 3482 1970 3514
rect 1794 3410 1826 3442
rect 1866 3410 1898 3442
rect 1938 3410 1970 3442
rect 1794 3338 1826 3370
rect 1866 3338 1898 3370
rect 1938 3338 1970 3370
rect 1794 3266 1826 3298
rect 1866 3266 1898 3298
rect 1938 3266 1970 3298
rect 1794 3194 1826 3226
rect 1866 3194 1898 3226
rect 1938 3194 1970 3226
rect 1794 3122 1826 3154
rect 1866 3122 1898 3154
rect 1938 3122 1970 3154
rect 1794 3050 1826 3082
rect 1866 3050 1898 3082
rect 1938 3050 1970 3082
rect 1794 2978 1826 3010
rect 1866 2978 1898 3010
rect 1938 2978 1970 3010
rect 1794 2906 1826 2938
rect 1866 2906 1898 2938
rect 1938 2906 1970 2938
rect 1794 2834 1826 2866
rect 1866 2834 1898 2866
rect 1938 2834 1970 2866
rect 1794 2762 1826 2794
rect 1866 2762 1898 2794
rect 1938 2762 1970 2794
rect 1794 2690 1826 2722
rect 1866 2690 1898 2722
rect 1938 2690 1970 2722
rect 1794 2618 1826 2650
rect 1866 2618 1898 2650
rect 1938 2618 1970 2650
rect 1794 2546 1826 2578
rect 1866 2546 1898 2578
rect 1938 2546 1970 2578
rect 1794 2474 1826 2506
rect 1866 2474 1898 2506
rect 1938 2474 1970 2506
rect 1794 2402 1826 2434
rect 1866 2402 1898 2434
rect 1938 2402 1970 2434
rect 1794 2330 1826 2362
rect 1866 2330 1898 2362
rect 1938 2330 1970 2362
rect 1794 2258 1826 2290
rect 1866 2258 1898 2290
rect 1938 2258 1970 2290
rect 1794 2186 1826 2218
rect 1866 2186 1898 2218
rect 1938 2186 1970 2218
rect 1794 2114 1826 2146
rect 1866 2114 1898 2146
rect 1938 2114 1970 2146
rect 1794 2042 1826 2074
rect 1866 2042 1898 2074
rect 1938 2042 1970 2074
rect 1794 1970 1826 2002
rect 1866 1970 1898 2002
rect 1938 1970 1970 2002
rect 1794 1898 1826 1930
rect 1866 1898 1898 1930
rect 1938 1898 1970 1930
rect 1794 1826 1826 1858
rect 1866 1826 1898 1858
rect 1938 1826 1970 1858
rect 1794 1754 1826 1786
rect 1866 1754 1898 1786
rect 1938 1754 1970 1786
rect 1794 1682 1826 1714
rect 1866 1682 1898 1714
rect 1938 1682 1970 1714
rect 1794 1610 1826 1642
rect 1866 1610 1898 1642
rect 1938 1610 1970 1642
rect 1794 1538 1826 1570
rect 1866 1538 1898 1570
rect 1938 1538 1970 1570
rect 1794 1466 1826 1498
rect 1866 1466 1898 1498
rect 1938 1466 1970 1498
rect 1794 1394 1826 1426
rect 1866 1394 1898 1426
rect 1938 1394 1970 1426
rect 1794 1322 1826 1354
rect 1866 1322 1898 1354
rect 1938 1322 1970 1354
rect 1794 1250 1826 1282
rect 1866 1250 1898 1282
rect 1938 1250 1970 1282
rect 1794 1178 1826 1210
rect 1866 1178 1898 1210
rect 1938 1178 1970 1210
rect 1794 1106 1826 1138
rect 1866 1106 1898 1138
rect 1938 1106 1970 1138
rect 1794 1034 1826 1066
rect 1866 1034 1898 1066
rect 1938 1034 1970 1066
rect 1794 962 1826 994
rect 1866 962 1898 994
rect 1938 962 1970 994
<< psubdiff >>
rect 84 7288 2780 7320
rect 84 7256 124 7288
rect 156 7256 196 7288
rect 228 7256 268 7288
rect 300 7256 340 7288
rect 372 7256 412 7288
rect 444 7256 484 7288
rect 516 7256 556 7288
rect 588 7256 628 7288
rect 660 7256 700 7288
rect 732 7256 772 7288
rect 804 7256 844 7288
rect 876 7256 916 7288
rect 948 7256 988 7288
rect 1020 7256 1060 7288
rect 1092 7256 1132 7288
rect 1164 7256 1204 7288
rect 1236 7256 1276 7288
rect 1308 7256 1348 7288
rect 1380 7256 1420 7288
rect 1452 7256 1492 7288
rect 1524 7256 1564 7288
rect 1596 7256 1636 7288
rect 1668 7256 1708 7288
rect 1740 7256 1780 7288
rect 1812 7256 1852 7288
rect 1884 7256 1924 7288
rect 1956 7256 1996 7288
rect 2028 7256 2068 7288
rect 2100 7256 2140 7288
rect 2172 7256 2212 7288
rect 2244 7256 2284 7288
rect 2316 7256 2356 7288
rect 2388 7256 2428 7288
rect 2460 7256 2500 7288
rect 2532 7256 2572 7288
rect 2604 7256 2644 7288
rect 2676 7256 2716 7288
rect 2748 7256 2780 7288
rect 84 7224 2780 7256
rect 84 7165 180 7224
rect 84 7133 116 7165
rect 148 7133 180 7165
rect 84 7093 180 7133
rect 84 7061 116 7093
rect 148 7061 180 7093
rect 84 7021 180 7061
rect 84 6989 116 7021
rect 148 6989 180 7021
rect 2684 7165 2780 7224
rect 2684 7133 2708 7165
rect 2740 7133 2780 7165
rect 2684 7093 2780 7133
rect 2684 7061 2708 7093
rect 2740 7061 2780 7093
rect 2684 7021 2780 7061
rect 84 6949 180 6989
rect 84 6917 116 6949
rect 148 6917 180 6949
rect 84 6877 180 6917
rect 84 6845 116 6877
rect 148 6845 180 6877
rect 84 6805 180 6845
rect 84 6773 116 6805
rect 148 6773 180 6805
rect 84 6733 180 6773
rect 84 6701 116 6733
rect 148 6701 180 6733
rect 84 6661 180 6701
rect 84 6629 116 6661
rect 148 6629 180 6661
rect 84 6589 180 6629
rect 84 6557 116 6589
rect 148 6557 180 6589
rect 84 6517 180 6557
rect 84 6485 116 6517
rect 148 6485 180 6517
rect 84 6445 180 6485
rect 84 6413 116 6445
rect 148 6413 180 6445
rect 84 6373 180 6413
rect 84 6341 116 6373
rect 148 6341 180 6373
rect 84 6301 180 6341
rect 84 6269 116 6301
rect 148 6269 180 6301
rect 84 6229 180 6269
rect 84 6197 116 6229
rect 148 6197 180 6229
rect 84 6157 180 6197
rect 84 6125 116 6157
rect 148 6125 180 6157
rect 84 6085 180 6125
rect 84 6053 116 6085
rect 148 6053 180 6085
rect 84 6013 180 6053
rect 84 5981 116 6013
rect 148 5981 180 6013
rect 84 5941 180 5981
rect 84 5909 116 5941
rect 148 5909 180 5941
rect 84 5869 180 5909
rect 84 5837 116 5869
rect 148 5837 180 5869
rect 84 5797 180 5837
rect 84 5765 116 5797
rect 148 5765 180 5797
rect 84 5725 180 5765
rect 84 5693 116 5725
rect 148 5693 180 5725
rect 84 5653 180 5693
rect 84 5621 116 5653
rect 148 5621 180 5653
rect 84 5581 180 5621
rect 84 5549 116 5581
rect 148 5549 180 5581
rect 84 5509 180 5549
rect 84 5477 116 5509
rect 148 5477 180 5509
rect 84 5437 180 5477
rect 84 5405 116 5437
rect 148 5405 180 5437
rect 84 5365 180 5405
rect 84 5333 116 5365
rect 148 5333 180 5365
rect 84 5293 180 5333
rect 84 5261 116 5293
rect 148 5261 180 5293
rect 84 5221 180 5261
rect 84 5189 116 5221
rect 148 5189 180 5221
rect 84 5149 180 5189
rect 84 5117 116 5149
rect 148 5117 180 5149
rect 84 5077 180 5117
rect 84 5045 116 5077
rect 148 5045 180 5077
rect 84 5005 180 5045
rect 84 4973 116 5005
rect 148 4973 180 5005
rect 84 4933 180 4973
rect 84 4901 116 4933
rect 148 4901 180 4933
rect 84 4861 180 4901
rect 84 4829 116 4861
rect 148 4829 180 4861
rect 84 4789 180 4829
rect 84 4757 116 4789
rect 148 4757 180 4789
rect 84 4717 180 4757
rect 84 4685 116 4717
rect 148 4685 180 4717
rect 84 4645 180 4685
rect 84 4613 116 4645
rect 148 4613 180 4645
rect 84 4573 180 4613
rect 84 4541 116 4573
rect 148 4541 180 4573
rect 84 4501 180 4541
rect 84 4469 116 4501
rect 148 4469 180 4501
rect 84 4429 180 4469
rect 84 4397 116 4429
rect 148 4397 180 4429
rect 84 4357 180 4397
rect 84 4325 116 4357
rect 148 4325 180 4357
rect 84 4285 180 4325
rect 84 4253 116 4285
rect 148 4253 180 4285
rect 84 4213 180 4253
rect 84 4181 116 4213
rect 148 4181 180 4213
rect 84 4141 180 4181
rect 84 4109 116 4141
rect 148 4109 180 4141
rect 84 4069 180 4109
rect 84 4037 116 4069
rect 148 4037 180 4069
rect 84 3997 180 4037
rect 84 3965 116 3997
rect 148 3965 180 3997
rect 84 3925 180 3965
rect 84 3893 116 3925
rect 148 3893 180 3925
rect 84 3853 180 3893
rect 84 3821 116 3853
rect 148 3821 180 3853
rect 84 3781 180 3821
rect 84 3749 116 3781
rect 148 3749 180 3781
rect 84 3709 180 3749
rect 84 3677 116 3709
rect 148 3677 180 3709
rect 84 3637 180 3677
rect 84 3605 116 3637
rect 148 3605 180 3637
rect 84 3565 180 3605
rect 84 3533 116 3565
rect 148 3533 180 3565
rect 84 3493 180 3533
rect 84 3461 116 3493
rect 148 3461 180 3493
rect 84 3421 180 3461
rect 84 3389 116 3421
rect 148 3389 180 3421
rect 84 3349 180 3389
rect 84 3317 116 3349
rect 148 3317 180 3349
rect 84 3277 180 3317
rect 84 3245 116 3277
rect 148 3245 180 3277
rect 84 3205 180 3245
rect 84 3173 116 3205
rect 148 3173 180 3205
rect 84 3133 180 3173
rect 84 3101 116 3133
rect 148 3101 180 3133
rect 84 3061 180 3101
rect 84 3029 116 3061
rect 148 3029 180 3061
rect 84 2989 180 3029
rect 84 2957 116 2989
rect 148 2957 180 2989
rect 84 2917 180 2957
rect 84 2885 116 2917
rect 148 2885 180 2917
rect 84 2845 180 2885
rect 84 2813 116 2845
rect 148 2813 180 2845
rect 84 2773 180 2813
rect 84 2741 116 2773
rect 148 2741 180 2773
rect 84 2701 180 2741
rect 84 2669 116 2701
rect 148 2669 180 2701
rect 84 2629 180 2669
rect 84 2597 116 2629
rect 148 2597 180 2629
rect 84 2557 180 2597
rect 84 2525 116 2557
rect 148 2525 180 2557
rect 84 2485 180 2525
rect 84 2453 116 2485
rect 148 2453 180 2485
rect 84 2413 180 2453
rect 84 2381 116 2413
rect 148 2381 180 2413
rect 84 2341 180 2381
rect 84 2309 116 2341
rect 148 2309 180 2341
rect 84 2269 180 2309
rect 84 2237 116 2269
rect 148 2237 180 2269
rect 84 2197 180 2237
rect 84 2165 116 2197
rect 148 2165 180 2197
rect 84 2125 180 2165
rect 84 2093 116 2125
rect 148 2093 180 2125
rect 84 2053 180 2093
rect 84 2021 116 2053
rect 148 2021 180 2053
rect 84 1981 180 2021
rect 84 1949 116 1981
rect 148 1949 180 1981
rect 84 1909 180 1949
rect 84 1877 116 1909
rect 148 1877 180 1909
rect 84 1837 180 1877
rect 84 1805 116 1837
rect 148 1805 180 1837
rect 84 1765 180 1805
rect 84 1733 116 1765
rect 148 1733 180 1765
rect 84 1693 180 1733
rect 84 1661 116 1693
rect 148 1661 180 1693
rect 84 1621 180 1661
rect 84 1589 116 1621
rect 148 1589 180 1621
rect 84 1549 180 1589
rect 84 1517 116 1549
rect 148 1517 180 1549
rect 84 1477 180 1517
rect 84 1445 116 1477
rect 148 1445 180 1477
rect 84 1405 180 1445
rect 84 1373 116 1405
rect 148 1373 180 1405
rect 84 1333 180 1373
rect 84 1301 116 1333
rect 148 1301 180 1333
rect 84 1261 180 1301
rect 84 1229 116 1261
rect 148 1229 180 1261
rect 84 1189 180 1229
rect 84 1157 116 1189
rect 148 1157 180 1189
rect 84 1117 180 1157
rect 84 1085 116 1117
rect 148 1085 180 1117
rect 84 1045 180 1085
rect 84 1013 116 1045
rect 148 1013 180 1045
rect 84 973 180 1013
rect 84 941 116 973
rect 148 941 180 973
rect 84 901 180 941
rect 84 869 116 901
rect 148 869 180 901
rect 84 829 180 869
rect 84 797 116 829
rect 148 797 180 829
rect 84 757 180 797
rect 84 725 116 757
rect 148 725 180 757
rect 84 685 180 725
rect 84 653 116 685
rect 148 653 180 685
rect 84 613 180 653
rect 84 581 116 613
rect 148 581 180 613
rect 84 541 180 581
rect 84 509 116 541
rect 148 509 180 541
rect 84 469 180 509
rect 84 437 116 469
rect 148 437 180 469
rect 84 397 180 437
rect 84 365 116 397
rect 148 365 180 397
rect 2684 6989 2708 7021
rect 2740 6989 2780 7021
rect 2684 6949 2780 6989
rect 2684 6917 2708 6949
rect 2740 6917 2780 6949
rect 2684 6877 2780 6917
rect 2684 6845 2708 6877
rect 2740 6845 2780 6877
rect 2684 6805 2780 6845
rect 2684 6773 2708 6805
rect 2740 6773 2780 6805
rect 2684 6733 2780 6773
rect 2684 6701 2708 6733
rect 2740 6701 2780 6733
rect 2684 6661 2780 6701
rect 2684 6629 2708 6661
rect 2740 6629 2780 6661
rect 2684 6589 2780 6629
rect 2684 6557 2708 6589
rect 2740 6557 2780 6589
rect 2684 6517 2780 6557
rect 2684 6485 2708 6517
rect 2740 6485 2780 6517
rect 2684 6445 2780 6485
rect 2684 6413 2708 6445
rect 2740 6413 2780 6445
rect 2684 6373 2780 6413
rect 2684 6341 2708 6373
rect 2740 6341 2780 6373
rect 2684 6301 2780 6341
rect 2684 6269 2708 6301
rect 2740 6269 2780 6301
rect 2684 6229 2780 6269
rect 2684 6197 2708 6229
rect 2740 6197 2780 6229
rect 2684 6157 2780 6197
rect 2684 6125 2708 6157
rect 2740 6125 2780 6157
rect 2684 6085 2780 6125
rect 2684 6053 2708 6085
rect 2740 6053 2780 6085
rect 2684 6013 2780 6053
rect 2684 5981 2708 6013
rect 2740 5981 2780 6013
rect 2684 5941 2780 5981
rect 2684 5909 2708 5941
rect 2740 5909 2780 5941
rect 2684 5869 2780 5909
rect 2684 5837 2708 5869
rect 2740 5837 2780 5869
rect 2684 5797 2780 5837
rect 2684 5765 2708 5797
rect 2740 5765 2780 5797
rect 2684 5725 2780 5765
rect 2684 5693 2708 5725
rect 2740 5693 2780 5725
rect 2684 5653 2780 5693
rect 2684 5621 2708 5653
rect 2740 5621 2780 5653
rect 2684 5581 2780 5621
rect 2684 5549 2708 5581
rect 2740 5549 2780 5581
rect 2684 5509 2780 5549
rect 2684 5477 2708 5509
rect 2740 5477 2780 5509
rect 2684 5437 2780 5477
rect 2684 5405 2708 5437
rect 2740 5405 2780 5437
rect 2684 5365 2780 5405
rect 2684 5333 2708 5365
rect 2740 5333 2780 5365
rect 2684 5293 2780 5333
rect 2684 5261 2708 5293
rect 2740 5261 2780 5293
rect 2684 5221 2780 5261
rect 2684 5189 2708 5221
rect 2740 5189 2780 5221
rect 2684 5149 2780 5189
rect 2684 5117 2708 5149
rect 2740 5117 2780 5149
rect 2684 5077 2780 5117
rect 2684 5045 2708 5077
rect 2740 5045 2780 5077
rect 2684 5005 2780 5045
rect 2684 4973 2708 5005
rect 2740 4973 2780 5005
rect 2684 4933 2780 4973
rect 2684 4901 2708 4933
rect 2740 4901 2780 4933
rect 2684 4861 2780 4901
rect 2684 4829 2708 4861
rect 2740 4829 2780 4861
rect 2684 4789 2780 4829
rect 2684 4757 2708 4789
rect 2740 4757 2780 4789
rect 2684 4717 2780 4757
rect 2684 4685 2708 4717
rect 2740 4685 2780 4717
rect 2684 4645 2780 4685
rect 2684 4613 2708 4645
rect 2740 4613 2780 4645
rect 2684 4573 2780 4613
rect 2684 4541 2708 4573
rect 2740 4541 2780 4573
rect 2684 4501 2780 4541
rect 2684 4469 2708 4501
rect 2740 4469 2780 4501
rect 2684 4429 2780 4469
rect 2684 4397 2708 4429
rect 2740 4397 2780 4429
rect 2684 4357 2780 4397
rect 2684 4325 2708 4357
rect 2740 4325 2780 4357
rect 2684 4285 2780 4325
rect 2684 4253 2708 4285
rect 2740 4253 2780 4285
rect 2684 4213 2780 4253
rect 2684 4181 2708 4213
rect 2740 4181 2780 4213
rect 2684 4141 2780 4181
rect 2684 4109 2708 4141
rect 2740 4109 2780 4141
rect 2684 4069 2780 4109
rect 2684 4037 2708 4069
rect 2740 4037 2780 4069
rect 2684 3997 2780 4037
rect 2684 3965 2708 3997
rect 2740 3965 2780 3997
rect 2684 3925 2780 3965
rect 2684 3893 2708 3925
rect 2740 3893 2780 3925
rect 2684 3853 2780 3893
rect 2684 3821 2708 3853
rect 2740 3821 2780 3853
rect 2684 3781 2780 3821
rect 2684 3749 2708 3781
rect 2740 3749 2780 3781
rect 2684 3709 2780 3749
rect 2684 3677 2708 3709
rect 2740 3677 2780 3709
rect 2684 3637 2780 3677
rect 2684 3605 2708 3637
rect 2740 3605 2780 3637
rect 2684 3565 2780 3605
rect 2684 3533 2708 3565
rect 2740 3533 2780 3565
rect 2684 3493 2780 3533
rect 2684 3461 2708 3493
rect 2740 3461 2780 3493
rect 2684 3421 2780 3461
rect 2684 3389 2708 3421
rect 2740 3389 2780 3421
rect 2684 3349 2780 3389
rect 2684 3317 2708 3349
rect 2740 3317 2780 3349
rect 2684 3277 2780 3317
rect 2684 3245 2708 3277
rect 2740 3245 2780 3277
rect 2684 3205 2780 3245
rect 2684 3173 2708 3205
rect 2740 3173 2780 3205
rect 2684 3133 2780 3173
rect 2684 3101 2708 3133
rect 2740 3101 2780 3133
rect 2684 3061 2780 3101
rect 2684 3029 2708 3061
rect 2740 3029 2780 3061
rect 2684 2989 2780 3029
rect 2684 2957 2708 2989
rect 2740 2957 2780 2989
rect 2684 2917 2780 2957
rect 2684 2885 2708 2917
rect 2740 2885 2780 2917
rect 2684 2845 2780 2885
rect 2684 2813 2708 2845
rect 2740 2813 2780 2845
rect 2684 2773 2780 2813
rect 2684 2741 2708 2773
rect 2740 2741 2780 2773
rect 2684 2701 2780 2741
rect 2684 2669 2708 2701
rect 2740 2669 2780 2701
rect 2684 2629 2780 2669
rect 2684 2597 2708 2629
rect 2740 2597 2780 2629
rect 2684 2557 2780 2597
rect 2684 2525 2708 2557
rect 2740 2525 2780 2557
rect 2684 2485 2780 2525
rect 2684 2453 2708 2485
rect 2740 2453 2780 2485
rect 2684 2413 2780 2453
rect 2684 2381 2708 2413
rect 2740 2381 2780 2413
rect 2684 2341 2780 2381
rect 2684 2309 2708 2341
rect 2740 2309 2780 2341
rect 2684 2269 2780 2309
rect 2684 2237 2708 2269
rect 2740 2237 2780 2269
rect 2684 2197 2780 2237
rect 2684 2165 2708 2197
rect 2740 2165 2780 2197
rect 2684 2125 2780 2165
rect 2684 2093 2708 2125
rect 2740 2093 2780 2125
rect 2684 2053 2780 2093
rect 2684 2021 2708 2053
rect 2740 2021 2780 2053
rect 2684 1981 2780 2021
rect 2684 1949 2708 1981
rect 2740 1949 2780 1981
rect 2684 1909 2780 1949
rect 2684 1877 2708 1909
rect 2740 1877 2780 1909
rect 2684 1837 2780 1877
rect 2684 1805 2708 1837
rect 2740 1805 2780 1837
rect 2684 1765 2780 1805
rect 2684 1733 2708 1765
rect 2740 1733 2780 1765
rect 2684 1693 2780 1733
rect 2684 1661 2708 1693
rect 2740 1661 2780 1693
rect 2684 1621 2780 1661
rect 2684 1589 2708 1621
rect 2740 1589 2780 1621
rect 2684 1549 2780 1589
rect 2684 1517 2708 1549
rect 2740 1517 2780 1549
rect 2684 1477 2780 1517
rect 2684 1445 2708 1477
rect 2740 1445 2780 1477
rect 2684 1405 2780 1445
rect 2684 1373 2708 1405
rect 2740 1373 2780 1405
rect 2684 1333 2780 1373
rect 2684 1301 2708 1333
rect 2740 1301 2780 1333
rect 2684 1261 2780 1301
rect 2684 1229 2708 1261
rect 2740 1229 2780 1261
rect 2684 1189 2780 1229
rect 2684 1157 2708 1189
rect 2740 1157 2780 1189
rect 2684 1117 2780 1157
rect 2684 1085 2708 1117
rect 2740 1085 2780 1117
rect 2684 1045 2780 1085
rect 2684 1013 2708 1045
rect 2740 1013 2780 1045
rect 2684 973 2780 1013
rect 2684 941 2708 973
rect 2740 941 2780 973
rect 2684 901 2780 941
rect 2684 869 2708 901
rect 2740 869 2780 901
rect 2684 829 2780 869
rect 2684 797 2708 829
rect 2740 797 2780 829
rect 2684 757 2780 797
rect 2684 725 2708 757
rect 2740 725 2780 757
rect 2684 685 2780 725
rect 2684 653 2708 685
rect 2740 653 2780 685
rect 2684 613 2780 653
rect 2684 581 2708 613
rect 2740 581 2780 613
rect 2684 541 2780 581
rect 2684 509 2708 541
rect 2740 509 2780 541
rect 2684 469 2780 509
rect 2684 437 2708 469
rect 2740 437 2780 469
rect 2684 397 2780 437
rect 84 325 180 365
rect 84 293 116 325
rect 148 293 180 325
rect 84 253 180 293
rect 84 221 116 253
rect 148 221 180 253
rect 84 186 180 221
rect 2684 365 2708 397
rect 2740 365 2780 397
rect 2684 325 2780 365
rect 2684 293 2708 325
rect 2740 293 2780 325
rect 2684 253 2780 293
rect 2684 221 2708 253
rect 2740 221 2780 253
rect 2684 186 2780 221
rect 84 154 2780 186
rect 84 122 124 154
rect 156 122 196 154
rect 228 122 268 154
rect 300 122 340 154
rect 372 122 412 154
rect 444 122 484 154
rect 516 122 556 154
rect 588 122 628 154
rect 660 122 700 154
rect 732 122 772 154
rect 804 122 844 154
rect 876 122 916 154
rect 948 122 988 154
rect 1020 122 1060 154
rect 1092 122 1132 154
rect 1164 122 1204 154
rect 1236 122 1276 154
rect 1308 122 1348 154
rect 1380 122 1420 154
rect 1452 122 1492 154
rect 1524 122 1564 154
rect 1596 122 1636 154
rect 1668 122 1708 154
rect 1740 122 1780 154
rect 1812 122 1852 154
rect 1884 122 1924 154
rect 1956 122 1996 154
rect 2028 122 2068 154
rect 2100 122 2140 154
rect 2172 122 2212 154
rect 2244 122 2284 154
rect 2316 122 2356 154
rect 2388 122 2428 154
rect 2460 122 2500 154
rect 2532 122 2572 154
rect 2604 122 2644 154
rect 2676 122 2716 154
rect 2748 122 2780 154
rect 84 90 2780 122
<< nsubdiff >>
rect 396 6980 2462 7014
rect 396 6948 447 6980
rect 479 6948 519 6980
rect 551 6948 591 6980
rect 623 6948 663 6980
rect 695 6948 735 6980
rect 767 6948 807 6980
rect 839 6948 879 6980
rect 911 6948 951 6980
rect 983 6948 1023 6980
rect 1055 6948 1095 6980
rect 1127 6948 1167 6980
rect 1199 6948 1239 6980
rect 1271 6948 1311 6980
rect 1343 6948 1383 6980
rect 1415 6948 1455 6980
rect 1487 6948 1527 6980
rect 1559 6948 1599 6980
rect 1631 6948 1671 6980
rect 1703 6948 1743 6980
rect 1775 6948 1815 6980
rect 1847 6948 1887 6980
rect 1919 6948 1959 6980
rect 1991 6948 2031 6980
rect 2063 6948 2103 6980
rect 2135 6948 2175 6980
rect 2207 6948 2247 6980
rect 2279 6948 2319 6980
rect 2351 6948 2391 6980
rect 2423 6948 2462 6980
rect 396 6908 2462 6948
rect 396 6876 447 6908
rect 479 6876 519 6908
rect 551 6876 591 6908
rect 623 6876 663 6908
rect 695 6876 735 6908
rect 767 6876 807 6908
rect 839 6876 879 6908
rect 911 6876 951 6908
rect 983 6876 1023 6908
rect 1055 6876 1095 6908
rect 1127 6876 1167 6908
rect 1199 6876 1239 6908
rect 1271 6876 1311 6908
rect 1343 6876 1383 6908
rect 1415 6876 1455 6908
rect 1487 6876 1527 6908
rect 1559 6876 1599 6908
rect 1631 6876 1671 6908
rect 1703 6876 1743 6908
rect 1775 6876 1815 6908
rect 1847 6876 1887 6908
rect 1919 6876 1959 6908
rect 1991 6876 2031 6908
rect 2063 6876 2103 6908
rect 2135 6876 2175 6908
rect 2207 6876 2247 6908
rect 2279 6876 2319 6908
rect 2351 6876 2391 6908
rect 2423 6876 2462 6908
rect 396 6836 2462 6876
rect 396 6804 447 6836
rect 479 6804 519 6836
rect 551 6804 591 6836
rect 623 6804 663 6836
rect 695 6804 735 6836
rect 767 6804 807 6836
rect 839 6804 879 6836
rect 911 6804 951 6836
rect 983 6804 1023 6836
rect 1055 6804 1095 6836
rect 1127 6804 1167 6836
rect 1199 6804 1239 6836
rect 1271 6804 1311 6836
rect 1343 6804 1383 6836
rect 1415 6804 1455 6836
rect 1487 6804 1527 6836
rect 1559 6804 1599 6836
rect 1631 6804 1671 6836
rect 1703 6804 1743 6836
rect 1775 6804 1815 6836
rect 1847 6804 1887 6836
rect 1919 6804 1959 6836
rect 1991 6804 2031 6836
rect 2063 6804 2103 6836
rect 2135 6804 2175 6836
rect 2207 6804 2247 6836
rect 2279 6804 2319 6836
rect 2351 6804 2391 6836
rect 2423 6804 2462 6836
rect 396 6762 2462 6804
rect 396 6761 648 6762
rect 396 6729 433 6761
rect 465 6729 505 6761
rect 537 6729 577 6761
rect 609 6729 648 6761
rect 396 6689 648 6729
rect 396 6657 433 6689
rect 465 6657 505 6689
rect 537 6657 577 6689
rect 609 6657 648 6689
rect 396 6617 648 6657
rect 396 6585 433 6617
rect 465 6585 505 6617
rect 537 6585 577 6617
rect 609 6585 648 6617
rect 396 6545 648 6585
rect 396 6513 433 6545
rect 465 6513 505 6545
rect 537 6513 577 6545
rect 609 6513 648 6545
rect 396 6473 648 6513
rect 1302 6761 1554 6762
rect 1302 6729 1345 6761
rect 1377 6729 1417 6761
rect 1449 6729 1489 6761
rect 1521 6729 1554 6761
rect 1302 6689 1554 6729
rect 1302 6657 1345 6689
rect 1377 6657 1417 6689
rect 1449 6657 1489 6689
rect 1521 6657 1554 6689
rect 1302 6617 1554 6657
rect 1302 6585 1345 6617
rect 1377 6585 1417 6617
rect 1449 6585 1489 6617
rect 1521 6585 1554 6617
rect 1302 6545 1554 6585
rect 1302 6513 1345 6545
rect 1377 6513 1417 6545
rect 1449 6513 1489 6545
rect 1521 6513 1554 6545
rect 396 6441 433 6473
rect 465 6441 505 6473
rect 537 6441 577 6473
rect 609 6441 648 6473
rect 396 6401 648 6441
rect 396 6369 433 6401
rect 465 6369 505 6401
rect 537 6369 577 6401
rect 609 6369 648 6401
rect 396 6329 648 6369
rect 396 6297 433 6329
rect 465 6297 505 6329
rect 537 6297 577 6329
rect 609 6297 648 6329
rect 396 6257 648 6297
rect 396 6225 433 6257
rect 465 6225 505 6257
rect 537 6225 577 6257
rect 609 6225 648 6257
rect 396 6185 648 6225
rect 396 6153 433 6185
rect 465 6153 505 6185
rect 537 6153 577 6185
rect 609 6153 648 6185
rect 396 6113 648 6153
rect 396 6081 433 6113
rect 465 6081 505 6113
rect 537 6081 577 6113
rect 609 6081 648 6113
rect 396 6041 648 6081
rect 396 6009 433 6041
rect 465 6009 505 6041
rect 537 6009 577 6041
rect 609 6009 648 6041
rect 396 5969 648 6009
rect 396 5937 433 5969
rect 465 5937 505 5969
rect 537 5937 577 5969
rect 609 5937 648 5969
rect 396 5897 648 5937
rect 396 5865 433 5897
rect 465 5865 505 5897
rect 537 5865 577 5897
rect 609 5865 648 5897
rect 396 5825 648 5865
rect 396 5793 433 5825
rect 465 5793 505 5825
rect 537 5793 577 5825
rect 609 5793 648 5825
rect 396 5753 648 5793
rect 396 5721 433 5753
rect 465 5721 505 5753
rect 537 5721 577 5753
rect 609 5721 648 5753
rect 396 5681 648 5721
rect 396 5649 433 5681
rect 465 5649 505 5681
rect 537 5649 577 5681
rect 609 5649 648 5681
rect 396 5609 648 5649
rect 396 5577 433 5609
rect 465 5577 505 5609
rect 537 5577 577 5609
rect 609 5577 648 5609
rect 396 5537 648 5577
rect 396 5505 433 5537
rect 465 5505 505 5537
rect 537 5505 577 5537
rect 609 5505 648 5537
rect 396 5465 648 5505
rect 396 5433 433 5465
rect 465 5433 505 5465
rect 537 5433 577 5465
rect 609 5433 648 5465
rect 396 5393 648 5433
rect 396 5361 433 5393
rect 465 5361 505 5393
rect 537 5361 577 5393
rect 609 5361 648 5393
rect 396 5321 648 5361
rect 396 5289 433 5321
rect 465 5289 505 5321
rect 537 5289 577 5321
rect 609 5289 648 5321
rect 396 5249 648 5289
rect 396 5217 433 5249
rect 465 5217 505 5249
rect 537 5217 577 5249
rect 609 5217 648 5249
rect 396 5177 648 5217
rect 396 5145 433 5177
rect 465 5145 505 5177
rect 537 5145 577 5177
rect 609 5145 648 5177
rect 396 5105 648 5145
rect 396 5073 433 5105
rect 465 5073 505 5105
rect 537 5073 577 5105
rect 609 5073 648 5105
rect 396 5033 648 5073
rect 396 5001 433 5033
rect 465 5001 505 5033
rect 537 5001 577 5033
rect 609 5001 648 5033
rect 396 4961 648 5001
rect 396 4929 433 4961
rect 465 4929 505 4961
rect 537 4929 577 4961
rect 609 4929 648 4961
rect 396 4889 648 4929
rect 396 4857 433 4889
rect 465 4857 505 4889
rect 537 4857 577 4889
rect 609 4857 648 4889
rect 396 4817 648 4857
rect 396 4785 433 4817
rect 465 4785 505 4817
rect 537 4785 577 4817
rect 609 4785 648 4817
rect 396 4745 648 4785
rect 396 4713 433 4745
rect 465 4713 505 4745
rect 537 4713 577 4745
rect 609 4713 648 4745
rect 396 4673 648 4713
rect 396 4641 433 4673
rect 465 4641 505 4673
rect 537 4641 577 4673
rect 609 4641 648 4673
rect 396 4601 648 4641
rect 396 4569 433 4601
rect 465 4569 505 4601
rect 537 4569 577 4601
rect 609 4569 648 4601
rect 396 4529 648 4569
rect 396 4497 433 4529
rect 465 4497 505 4529
rect 537 4497 577 4529
rect 609 4497 648 4529
rect 396 4457 648 4497
rect 396 4425 433 4457
rect 465 4425 505 4457
rect 537 4425 577 4457
rect 609 4425 648 4457
rect 396 4385 648 4425
rect 396 4353 433 4385
rect 465 4353 505 4385
rect 537 4353 577 4385
rect 609 4353 648 4385
rect 396 4313 648 4353
rect 396 4281 433 4313
rect 465 4281 505 4313
rect 537 4281 577 4313
rect 609 4281 648 4313
rect 396 4241 648 4281
rect 396 4209 433 4241
rect 465 4209 505 4241
rect 537 4209 577 4241
rect 609 4209 648 4241
rect 396 4169 648 4209
rect 396 4137 433 4169
rect 465 4137 505 4169
rect 537 4137 577 4169
rect 609 4137 648 4169
rect 396 4097 648 4137
rect 396 4065 433 4097
rect 465 4065 505 4097
rect 537 4065 577 4097
rect 609 4065 648 4097
rect 396 4025 648 4065
rect 396 3993 433 4025
rect 465 3993 505 4025
rect 537 3993 577 4025
rect 609 3993 648 4025
rect 396 3953 648 3993
rect 396 3921 433 3953
rect 465 3921 505 3953
rect 537 3921 577 3953
rect 609 3921 648 3953
rect 396 3881 648 3921
rect 396 3849 433 3881
rect 465 3849 505 3881
rect 537 3849 577 3881
rect 609 3849 648 3881
rect 396 3809 648 3849
rect 396 3777 433 3809
rect 465 3777 505 3809
rect 537 3777 577 3809
rect 609 3777 648 3809
rect 396 3737 648 3777
rect 396 3705 433 3737
rect 465 3705 505 3737
rect 537 3705 577 3737
rect 609 3705 648 3737
rect 396 3665 648 3705
rect 396 3633 433 3665
rect 465 3633 505 3665
rect 537 3633 577 3665
rect 609 3633 648 3665
rect 396 3593 648 3633
rect 396 3561 433 3593
rect 465 3561 505 3593
rect 537 3561 577 3593
rect 609 3561 648 3593
rect 396 3521 648 3561
rect 396 3489 433 3521
rect 465 3489 505 3521
rect 537 3489 577 3521
rect 609 3489 648 3521
rect 396 3449 648 3489
rect 396 3417 433 3449
rect 465 3417 505 3449
rect 537 3417 577 3449
rect 609 3417 648 3449
rect 396 3377 648 3417
rect 396 3345 433 3377
rect 465 3345 505 3377
rect 537 3345 577 3377
rect 609 3345 648 3377
rect 396 3305 648 3345
rect 396 3273 433 3305
rect 465 3273 505 3305
rect 537 3273 577 3305
rect 609 3273 648 3305
rect 396 3233 648 3273
rect 396 3201 433 3233
rect 465 3201 505 3233
rect 537 3201 577 3233
rect 609 3201 648 3233
rect 396 3161 648 3201
rect 396 3129 433 3161
rect 465 3129 505 3161
rect 537 3129 577 3161
rect 609 3129 648 3161
rect 396 3089 648 3129
rect 396 3057 433 3089
rect 465 3057 505 3089
rect 537 3057 577 3089
rect 609 3057 648 3089
rect 396 3017 648 3057
rect 396 2985 433 3017
rect 465 2985 505 3017
rect 537 2985 577 3017
rect 609 2985 648 3017
rect 396 2945 648 2985
rect 396 2913 433 2945
rect 465 2913 505 2945
rect 537 2913 577 2945
rect 609 2913 648 2945
rect 396 2873 648 2913
rect 396 2841 433 2873
rect 465 2841 505 2873
rect 537 2841 577 2873
rect 609 2841 648 2873
rect 396 2801 648 2841
rect 396 2769 433 2801
rect 465 2769 505 2801
rect 537 2769 577 2801
rect 609 2769 648 2801
rect 396 2729 648 2769
rect 396 2697 433 2729
rect 465 2697 505 2729
rect 537 2697 577 2729
rect 609 2697 648 2729
rect 396 2657 648 2697
rect 396 2625 433 2657
rect 465 2625 505 2657
rect 537 2625 577 2657
rect 609 2625 648 2657
rect 396 2585 648 2625
rect 396 2553 433 2585
rect 465 2553 505 2585
rect 537 2553 577 2585
rect 609 2553 648 2585
rect 396 2513 648 2553
rect 396 2481 433 2513
rect 465 2481 505 2513
rect 537 2481 577 2513
rect 609 2481 648 2513
rect 396 2441 648 2481
rect 396 2409 433 2441
rect 465 2409 505 2441
rect 537 2409 577 2441
rect 609 2409 648 2441
rect 396 2369 648 2409
rect 396 2337 433 2369
rect 465 2337 505 2369
rect 537 2337 577 2369
rect 609 2337 648 2369
rect 396 2297 648 2337
rect 396 2265 433 2297
rect 465 2265 505 2297
rect 537 2265 577 2297
rect 609 2265 648 2297
rect 396 2225 648 2265
rect 396 2193 433 2225
rect 465 2193 505 2225
rect 537 2193 577 2225
rect 609 2193 648 2225
rect 396 2153 648 2193
rect 396 2121 433 2153
rect 465 2121 505 2153
rect 537 2121 577 2153
rect 609 2121 648 2153
rect 396 2081 648 2121
rect 396 2049 433 2081
rect 465 2049 505 2081
rect 537 2049 577 2081
rect 609 2049 648 2081
rect 396 2009 648 2049
rect 396 1977 433 2009
rect 465 1977 505 2009
rect 537 1977 577 2009
rect 609 1977 648 2009
rect 396 1937 648 1977
rect 396 1905 433 1937
rect 465 1905 505 1937
rect 537 1905 577 1937
rect 609 1905 648 1937
rect 396 1865 648 1905
rect 396 1833 433 1865
rect 465 1833 505 1865
rect 537 1833 577 1865
rect 609 1833 648 1865
rect 396 1793 648 1833
rect 396 1761 433 1793
rect 465 1761 505 1793
rect 537 1761 577 1793
rect 609 1761 648 1793
rect 396 1721 648 1761
rect 396 1689 433 1721
rect 465 1689 505 1721
rect 537 1689 577 1721
rect 609 1689 648 1721
rect 396 1649 648 1689
rect 396 1617 433 1649
rect 465 1617 505 1649
rect 537 1617 577 1649
rect 609 1617 648 1649
rect 396 1577 648 1617
rect 396 1545 433 1577
rect 465 1545 505 1577
rect 537 1545 577 1577
rect 609 1545 648 1577
rect 396 1505 648 1545
rect 396 1473 433 1505
rect 465 1473 505 1505
rect 537 1473 577 1505
rect 609 1473 648 1505
rect 396 1433 648 1473
rect 396 1401 433 1433
rect 465 1401 505 1433
rect 537 1401 577 1433
rect 609 1401 648 1433
rect 396 1361 648 1401
rect 396 1329 433 1361
rect 465 1329 505 1361
rect 537 1329 577 1361
rect 609 1329 648 1361
rect 396 1289 648 1329
rect 396 1257 433 1289
rect 465 1257 505 1289
rect 537 1257 577 1289
rect 609 1257 648 1289
rect 396 1217 648 1257
rect 396 1185 433 1217
rect 465 1185 505 1217
rect 537 1185 577 1217
rect 609 1185 648 1217
rect 396 1145 648 1185
rect 396 1113 433 1145
rect 465 1113 505 1145
rect 537 1113 577 1145
rect 609 1113 648 1145
rect 396 1073 648 1113
rect 396 1041 433 1073
rect 465 1041 505 1073
rect 537 1041 577 1073
rect 609 1041 648 1073
rect 396 1001 648 1041
rect 396 969 433 1001
rect 465 969 505 1001
rect 537 969 577 1001
rect 609 969 648 1001
rect 396 929 648 969
rect 1302 6473 1554 6513
rect 2210 6761 2462 6762
rect 2210 6729 2257 6761
rect 2289 6729 2329 6761
rect 2361 6729 2401 6761
rect 2433 6729 2462 6761
rect 2210 6689 2462 6729
rect 2210 6657 2257 6689
rect 2289 6657 2329 6689
rect 2361 6657 2401 6689
rect 2433 6657 2462 6689
rect 2210 6617 2462 6657
rect 2210 6585 2257 6617
rect 2289 6585 2329 6617
rect 2361 6585 2401 6617
rect 2433 6585 2462 6617
rect 2210 6545 2462 6585
rect 2210 6513 2257 6545
rect 2289 6513 2329 6545
rect 2361 6513 2401 6545
rect 2433 6513 2462 6545
rect 1302 6441 1345 6473
rect 1377 6441 1417 6473
rect 1449 6441 1489 6473
rect 1521 6441 1554 6473
rect 1302 6401 1554 6441
rect 1302 6369 1345 6401
rect 1377 6369 1417 6401
rect 1449 6369 1489 6401
rect 1521 6369 1554 6401
rect 1302 6329 1554 6369
rect 1302 6297 1345 6329
rect 1377 6297 1417 6329
rect 1449 6297 1489 6329
rect 1521 6297 1554 6329
rect 1302 6257 1554 6297
rect 1302 6225 1345 6257
rect 1377 6225 1417 6257
rect 1449 6225 1489 6257
rect 1521 6225 1554 6257
rect 1302 6185 1554 6225
rect 1302 6153 1345 6185
rect 1377 6153 1417 6185
rect 1449 6153 1489 6185
rect 1521 6153 1554 6185
rect 1302 6113 1554 6153
rect 1302 6081 1345 6113
rect 1377 6081 1417 6113
rect 1449 6081 1489 6113
rect 1521 6081 1554 6113
rect 1302 6041 1554 6081
rect 1302 6009 1345 6041
rect 1377 6009 1417 6041
rect 1449 6009 1489 6041
rect 1521 6009 1554 6041
rect 1302 5969 1554 6009
rect 1302 5937 1345 5969
rect 1377 5937 1417 5969
rect 1449 5937 1489 5969
rect 1521 5937 1554 5969
rect 1302 5897 1554 5937
rect 1302 5865 1345 5897
rect 1377 5865 1417 5897
rect 1449 5865 1489 5897
rect 1521 5865 1554 5897
rect 1302 5825 1554 5865
rect 1302 5793 1345 5825
rect 1377 5793 1417 5825
rect 1449 5793 1489 5825
rect 1521 5793 1554 5825
rect 1302 5753 1554 5793
rect 1302 5721 1345 5753
rect 1377 5721 1417 5753
rect 1449 5721 1489 5753
rect 1521 5721 1554 5753
rect 1302 5681 1554 5721
rect 1302 5649 1345 5681
rect 1377 5649 1417 5681
rect 1449 5649 1489 5681
rect 1521 5649 1554 5681
rect 1302 5609 1554 5649
rect 1302 5577 1345 5609
rect 1377 5577 1417 5609
rect 1449 5577 1489 5609
rect 1521 5577 1554 5609
rect 1302 5537 1554 5577
rect 1302 5505 1345 5537
rect 1377 5505 1417 5537
rect 1449 5505 1489 5537
rect 1521 5505 1554 5537
rect 1302 5465 1554 5505
rect 1302 5433 1345 5465
rect 1377 5433 1417 5465
rect 1449 5433 1489 5465
rect 1521 5433 1554 5465
rect 1302 5393 1554 5433
rect 1302 5361 1345 5393
rect 1377 5361 1417 5393
rect 1449 5361 1489 5393
rect 1521 5361 1554 5393
rect 1302 5321 1554 5361
rect 1302 5289 1345 5321
rect 1377 5289 1417 5321
rect 1449 5289 1489 5321
rect 1521 5289 1554 5321
rect 1302 5249 1554 5289
rect 1302 5217 1345 5249
rect 1377 5217 1417 5249
rect 1449 5217 1489 5249
rect 1521 5217 1554 5249
rect 1302 5177 1554 5217
rect 1302 5145 1345 5177
rect 1377 5145 1417 5177
rect 1449 5145 1489 5177
rect 1521 5145 1554 5177
rect 1302 5105 1554 5145
rect 1302 5073 1345 5105
rect 1377 5073 1417 5105
rect 1449 5073 1489 5105
rect 1521 5073 1554 5105
rect 1302 5033 1554 5073
rect 1302 5001 1345 5033
rect 1377 5001 1417 5033
rect 1449 5001 1489 5033
rect 1521 5001 1554 5033
rect 1302 4961 1554 5001
rect 1302 4929 1345 4961
rect 1377 4929 1417 4961
rect 1449 4929 1489 4961
rect 1521 4929 1554 4961
rect 1302 4889 1554 4929
rect 1302 4857 1345 4889
rect 1377 4857 1417 4889
rect 1449 4857 1489 4889
rect 1521 4857 1554 4889
rect 1302 4817 1554 4857
rect 1302 4785 1345 4817
rect 1377 4785 1417 4817
rect 1449 4785 1489 4817
rect 1521 4785 1554 4817
rect 1302 4745 1554 4785
rect 1302 4713 1345 4745
rect 1377 4713 1417 4745
rect 1449 4713 1489 4745
rect 1521 4713 1554 4745
rect 1302 4673 1554 4713
rect 1302 4641 1345 4673
rect 1377 4641 1417 4673
rect 1449 4641 1489 4673
rect 1521 4641 1554 4673
rect 1302 4601 1554 4641
rect 1302 4569 1345 4601
rect 1377 4569 1417 4601
rect 1449 4569 1489 4601
rect 1521 4569 1554 4601
rect 1302 4529 1554 4569
rect 1302 4497 1345 4529
rect 1377 4497 1417 4529
rect 1449 4497 1489 4529
rect 1521 4497 1554 4529
rect 1302 4457 1554 4497
rect 1302 4425 1345 4457
rect 1377 4425 1417 4457
rect 1449 4425 1489 4457
rect 1521 4425 1554 4457
rect 1302 4385 1554 4425
rect 1302 4353 1345 4385
rect 1377 4353 1417 4385
rect 1449 4353 1489 4385
rect 1521 4353 1554 4385
rect 1302 4313 1554 4353
rect 1302 4281 1345 4313
rect 1377 4281 1417 4313
rect 1449 4281 1489 4313
rect 1521 4281 1554 4313
rect 1302 4241 1554 4281
rect 1302 4209 1345 4241
rect 1377 4209 1417 4241
rect 1449 4209 1489 4241
rect 1521 4209 1554 4241
rect 1302 4169 1554 4209
rect 1302 4137 1345 4169
rect 1377 4137 1417 4169
rect 1449 4137 1489 4169
rect 1521 4137 1554 4169
rect 1302 4097 1554 4137
rect 1302 4065 1345 4097
rect 1377 4065 1417 4097
rect 1449 4065 1489 4097
rect 1521 4065 1554 4097
rect 1302 4025 1554 4065
rect 1302 3993 1345 4025
rect 1377 3993 1417 4025
rect 1449 3993 1489 4025
rect 1521 3993 1554 4025
rect 1302 3953 1554 3993
rect 1302 3921 1345 3953
rect 1377 3921 1417 3953
rect 1449 3921 1489 3953
rect 1521 3921 1554 3953
rect 1302 3881 1554 3921
rect 1302 3849 1345 3881
rect 1377 3849 1417 3881
rect 1449 3849 1489 3881
rect 1521 3849 1554 3881
rect 1302 3809 1554 3849
rect 1302 3777 1345 3809
rect 1377 3777 1417 3809
rect 1449 3777 1489 3809
rect 1521 3777 1554 3809
rect 1302 3737 1554 3777
rect 1302 3705 1345 3737
rect 1377 3705 1417 3737
rect 1449 3705 1489 3737
rect 1521 3705 1554 3737
rect 1302 3665 1554 3705
rect 1302 3633 1345 3665
rect 1377 3633 1417 3665
rect 1449 3633 1489 3665
rect 1521 3633 1554 3665
rect 1302 3593 1554 3633
rect 1302 3561 1345 3593
rect 1377 3561 1417 3593
rect 1449 3561 1489 3593
rect 1521 3561 1554 3593
rect 1302 3521 1554 3561
rect 1302 3489 1345 3521
rect 1377 3489 1417 3521
rect 1449 3489 1489 3521
rect 1521 3489 1554 3521
rect 1302 3449 1554 3489
rect 1302 3417 1345 3449
rect 1377 3417 1417 3449
rect 1449 3417 1489 3449
rect 1521 3417 1554 3449
rect 1302 3377 1554 3417
rect 1302 3345 1345 3377
rect 1377 3345 1417 3377
rect 1449 3345 1489 3377
rect 1521 3345 1554 3377
rect 1302 3305 1554 3345
rect 1302 3273 1345 3305
rect 1377 3273 1417 3305
rect 1449 3273 1489 3305
rect 1521 3273 1554 3305
rect 1302 3233 1554 3273
rect 1302 3201 1345 3233
rect 1377 3201 1417 3233
rect 1449 3201 1489 3233
rect 1521 3201 1554 3233
rect 1302 3161 1554 3201
rect 1302 3129 1345 3161
rect 1377 3129 1417 3161
rect 1449 3129 1489 3161
rect 1521 3129 1554 3161
rect 1302 3089 1554 3129
rect 1302 3057 1345 3089
rect 1377 3057 1417 3089
rect 1449 3057 1489 3089
rect 1521 3057 1554 3089
rect 1302 3017 1554 3057
rect 1302 2985 1345 3017
rect 1377 2985 1417 3017
rect 1449 2985 1489 3017
rect 1521 2985 1554 3017
rect 1302 2945 1554 2985
rect 1302 2913 1345 2945
rect 1377 2913 1417 2945
rect 1449 2913 1489 2945
rect 1521 2913 1554 2945
rect 1302 2873 1554 2913
rect 1302 2841 1345 2873
rect 1377 2841 1417 2873
rect 1449 2841 1489 2873
rect 1521 2841 1554 2873
rect 1302 2801 1554 2841
rect 1302 2769 1345 2801
rect 1377 2769 1417 2801
rect 1449 2769 1489 2801
rect 1521 2769 1554 2801
rect 1302 2729 1554 2769
rect 1302 2697 1345 2729
rect 1377 2697 1417 2729
rect 1449 2697 1489 2729
rect 1521 2697 1554 2729
rect 1302 2657 1554 2697
rect 1302 2625 1345 2657
rect 1377 2625 1417 2657
rect 1449 2625 1489 2657
rect 1521 2625 1554 2657
rect 1302 2585 1554 2625
rect 1302 2553 1345 2585
rect 1377 2553 1417 2585
rect 1449 2553 1489 2585
rect 1521 2553 1554 2585
rect 1302 2513 1554 2553
rect 1302 2481 1345 2513
rect 1377 2481 1417 2513
rect 1449 2481 1489 2513
rect 1521 2481 1554 2513
rect 1302 2441 1554 2481
rect 1302 2409 1345 2441
rect 1377 2409 1417 2441
rect 1449 2409 1489 2441
rect 1521 2409 1554 2441
rect 1302 2369 1554 2409
rect 1302 2337 1345 2369
rect 1377 2337 1417 2369
rect 1449 2337 1489 2369
rect 1521 2337 1554 2369
rect 1302 2297 1554 2337
rect 1302 2265 1345 2297
rect 1377 2265 1417 2297
rect 1449 2265 1489 2297
rect 1521 2265 1554 2297
rect 1302 2225 1554 2265
rect 1302 2193 1345 2225
rect 1377 2193 1417 2225
rect 1449 2193 1489 2225
rect 1521 2193 1554 2225
rect 1302 2153 1554 2193
rect 1302 2121 1345 2153
rect 1377 2121 1417 2153
rect 1449 2121 1489 2153
rect 1521 2121 1554 2153
rect 1302 2081 1554 2121
rect 1302 2049 1345 2081
rect 1377 2049 1417 2081
rect 1449 2049 1489 2081
rect 1521 2049 1554 2081
rect 1302 2009 1554 2049
rect 1302 1977 1345 2009
rect 1377 1977 1417 2009
rect 1449 1977 1489 2009
rect 1521 1977 1554 2009
rect 1302 1937 1554 1977
rect 1302 1905 1345 1937
rect 1377 1905 1417 1937
rect 1449 1905 1489 1937
rect 1521 1905 1554 1937
rect 1302 1865 1554 1905
rect 1302 1833 1345 1865
rect 1377 1833 1417 1865
rect 1449 1833 1489 1865
rect 1521 1833 1554 1865
rect 1302 1793 1554 1833
rect 1302 1761 1345 1793
rect 1377 1761 1417 1793
rect 1449 1761 1489 1793
rect 1521 1761 1554 1793
rect 1302 1721 1554 1761
rect 1302 1689 1345 1721
rect 1377 1689 1417 1721
rect 1449 1689 1489 1721
rect 1521 1689 1554 1721
rect 1302 1649 1554 1689
rect 1302 1617 1345 1649
rect 1377 1617 1417 1649
rect 1449 1617 1489 1649
rect 1521 1617 1554 1649
rect 1302 1577 1554 1617
rect 1302 1545 1345 1577
rect 1377 1545 1417 1577
rect 1449 1545 1489 1577
rect 1521 1545 1554 1577
rect 1302 1505 1554 1545
rect 1302 1473 1345 1505
rect 1377 1473 1417 1505
rect 1449 1473 1489 1505
rect 1521 1473 1554 1505
rect 1302 1433 1554 1473
rect 1302 1401 1345 1433
rect 1377 1401 1417 1433
rect 1449 1401 1489 1433
rect 1521 1401 1554 1433
rect 1302 1361 1554 1401
rect 1302 1329 1345 1361
rect 1377 1329 1417 1361
rect 1449 1329 1489 1361
rect 1521 1329 1554 1361
rect 1302 1289 1554 1329
rect 1302 1257 1345 1289
rect 1377 1257 1417 1289
rect 1449 1257 1489 1289
rect 1521 1257 1554 1289
rect 1302 1217 1554 1257
rect 1302 1185 1345 1217
rect 1377 1185 1417 1217
rect 1449 1185 1489 1217
rect 1521 1185 1554 1217
rect 1302 1145 1554 1185
rect 1302 1113 1345 1145
rect 1377 1113 1417 1145
rect 1449 1113 1489 1145
rect 1521 1113 1554 1145
rect 1302 1073 1554 1113
rect 1302 1041 1345 1073
rect 1377 1041 1417 1073
rect 1449 1041 1489 1073
rect 1521 1041 1554 1073
rect 1302 1001 1554 1041
rect 1302 969 1345 1001
rect 1377 969 1417 1001
rect 1449 969 1489 1001
rect 1521 969 1554 1001
rect 396 897 433 929
rect 465 897 505 929
rect 537 897 577 929
rect 609 897 648 929
rect 396 857 648 897
rect 396 825 433 857
rect 465 825 505 857
rect 537 825 577 857
rect 609 825 648 857
rect 396 785 648 825
rect 396 753 433 785
rect 465 753 505 785
rect 537 753 577 785
rect 609 753 648 785
rect 396 713 648 753
rect 396 681 433 713
rect 465 681 505 713
rect 537 681 577 713
rect 609 681 648 713
rect 396 648 648 681
rect 1302 929 1554 969
rect 2210 6473 2462 6513
rect 2210 6441 2257 6473
rect 2289 6441 2329 6473
rect 2361 6441 2401 6473
rect 2433 6441 2462 6473
rect 2210 6401 2462 6441
rect 2210 6369 2257 6401
rect 2289 6369 2329 6401
rect 2361 6369 2401 6401
rect 2433 6369 2462 6401
rect 2210 6329 2462 6369
rect 2210 6297 2257 6329
rect 2289 6297 2329 6329
rect 2361 6297 2401 6329
rect 2433 6297 2462 6329
rect 2210 6257 2462 6297
rect 2210 6225 2257 6257
rect 2289 6225 2329 6257
rect 2361 6225 2401 6257
rect 2433 6225 2462 6257
rect 2210 6185 2462 6225
rect 2210 6153 2257 6185
rect 2289 6153 2329 6185
rect 2361 6153 2401 6185
rect 2433 6153 2462 6185
rect 2210 6113 2462 6153
rect 2210 6081 2257 6113
rect 2289 6081 2329 6113
rect 2361 6081 2401 6113
rect 2433 6081 2462 6113
rect 2210 6041 2462 6081
rect 2210 6009 2257 6041
rect 2289 6009 2329 6041
rect 2361 6009 2401 6041
rect 2433 6009 2462 6041
rect 2210 5969 2462 6009
rect 2210 5937 2257 5969
rect 2289 5937 2329 5969
rect 2361 5937 2401 5969
rect 2433 5937 2462 5969
rect 2210 5897 2462 5937
rect 2210 5865 2257 5897
rect 2289 5865 2329 5897
rect 2361 5865 2401 5897
rect 2433 5865 2462 5897
rect 2210 5825 2462 5865
rect 2210 5793 2257 5825
rect 2289 5793 2329 5825
rect 2361 5793 2401 5825
rect 2433 5793 2462 5825
rect 2210 5753 2462 5793
rect 2210 5721 2257 5753
rect 2289 5721 2329 5753
rect 2361 5721 2401 5753
rect 2433 5721 2462 5753
rect 2210 5681 2462 5721
rect 2210 5649 2257 5681
rect 2289 5649 2329 5681
rect 2361 5649 2401 5681
rect 2433 5649 2462 5681
rect 2210 5609 2462 5649
rect 2210 5577 2257 5609
rect 2289 5577 2329 5609
rect 2361 5577 2401 5609
rect 2433 5577 2462 5609
rect 2210 5537 2462 5577
rect 2210 5505 2257 5537
rect 2289 5505 2329 5537
rect 2361 5505 2401 5537
rect 2433 5505 2462 5537
rect 2210 5465 2462 5505
rect 2210 5433 2257 5465
rect 2289 5433 2329 5465
rect 2361 5433 2401 5465
rect 2433 5433 2462 5465
rect 2210 5393 2462 5433
rect 2210 5361 2257 5393
rect 2289 5361 2329 5393
rect 2361 5361 2401 5393
rect 2433 5361 2462 5393
rect 2210 5321 2462 5361
rect 2210 5289 2257 5321
rect 2289 5289 2329 5321
rect 2361 5289 2401 5321
rect 2433 5289 2462 5321
rect 2210 5249 2462 5289
rect 2210 5217 2257 5249
rect 2289 5217 2329 5249
rect 2361 5217 2401 5249
rect 2433 5217 2462 5249
rect 2210 5177 2462 5217
rect 2210 5145 2257 5177
rect 2289 5145 2329 5177
rect 2361 5145 2401 5177
rect 2433 5145 2462 5177
rect 2210 5105 2462 5145
rect 2210 5073 2257 5105
rect 2289 5073 2329 5105
rect 2361 5073 2401 5105
rect 2433 5073 2462 5105
rect 2210 5033 2462 5073
rect 2210 5001 2257 5033
rect 2289 5001 2329 5033
rect 2361 5001 2401 5033
rect 2433 5001 2462 5033
rect 2210 4961 2462 5001
rect 2210 4929 2257 4961
rect 2289 4929 2329 4961
rect 2361 4929 2401 4961
rect 2433 4929 2462 4961
rect 2210 4889 2462 4929
rect 2210 4857 2257 4889
rect 2289 4857 2329 4889
rect 2361 4857 2401 4889
rect 2433 4857 2462 4889
rect 2210 4817 2462 4857
rect 2210 4785 2257 4817
rect 2289 4785 2329 4817
rect 2361 4785 2401 4817
rect 2433 4785 2462 4817
rect 2210 4745 2462 4785
rect 2210 4713 2257 4745
rect 2289 4713 2329 4745
rect 2361 4713 2401 4745
rect 2433 4713 2462 4745
rect 2210 4673 2462 4713
rect 2210 4641 2257 4673
rect 2289 4641 2329 4673
rect 2361 4641 2401 4673
rect 2433 4641 2462 4673
rect 2210 4601 2462 4641
rect 2210 4569 2257 4601
rect 2289 4569 2329 4601
rect 2361 4569 2401 4601
rect 2433 4569 2462 4601
rect 2210 4529 2462 4569
rect 2210 4497 2257 4529
rect 2289 4497 2329 4529
rect 2361 4497 2401 4529
rect 2433 4497 2462 4529
rect 2210 4457 2462 4497
rect 2210 4425 2257 4457
rect 2289 4425 2329 4457
rect 2361 4425 2401 4457
rect 2433 4425 2462 4457
rect 2210 4385 2462 4425
rect 2210 4353 2257 4385
rect 2289 4353 2329 4385
rect 2361 4353 2401 4385
rect 2433 4353 2462 4385
rect 2210 4313 2462 4353
rect 2210 4281 2257 4313
rect 2289 4281 2329 4313
rect 2361 4281 2401 4313
rect 2433 4281 2462 4313
rect 2210 4241 2462 4281
rect 2210 4209 2257 4241
rect 2289 4209 2329 4241
rect 2361 4209 2401 4241
rect 2433 4209 2462 4241
rect 2210 4169 2462 4209
rect 2210 4137 2257 4169
rect 2289 4137 2329 4169
rect 2361 4137 2401 4169
rect 2433 4137 2462 4169
rect 2210 4097 2462 4137
rect 2210 4065 2257 4097
rect 2289 4065 2329 4097
rect 2361 4065 2401 4097
rect 2433 4065 2462 4097
rect 2210 4025 2462 4065
rect 2210 3993 2257 4025
rect 2289 3993 2329 4025
rect 2361 3993 2401 4025
rect 2433 3993 2462 4025
rect 2210 3953 2462 3993
rect 2210 3921 2257 3953
rect 2289 3921 2329 3953
rect 2361 3921 2401 3953
rect 2433 3921 2462 3953
rect 2210 3881 2462 3921
rect 2210 3849 2257 3881
rect 2289 3849 2329 3881
rect 2361 3849 2401 3881
rect 2433 3849 2462 3881
rect 2210 3809 2462 3849
rect 2210 3777 2257 3809
rect 2289 3777 2329 3809
rect 2361 3777 2401 3809
rect 2433 3777 2462 3809
rect 2210 3737 2462 3777
rect 2210 3705 2257 3737
rect 2289 3705 2329 3737
rect 2361 3705 2401 3737
rect 2433 3705 2462 3737
rect 2210 3665 2462 3705
rect 2210 3633 2257 3665
rect 2289 3633 2329 3665
rect 2361 3633 2401 3665
rect 2433 3633 2462 3665
rect 2210 3593 2462 3633
rect 2210 3561 2257 3593
rect 2289 3561 2329 3593
rect 2361 3561 2401 3593
rect 2433 3561 2462 3593
rect 2210 3521 2462 3561
rect 2210 3489 2257 3521
rect 2289 3489 2329 3521
rect 2361 3489 2401 3521
rect 2433 3489 2462 3521
rect 2210 3449 2462 3489
rect 2210 3417 2257 3449
rect 2289 3417 2329 3449
rect 2361 3417 2401 3449
rect 2433 3417 2462 3449
rect 2210 3377 2462 3417
rect 2210 3345 2257 3377
rect 2289 3345 2329 3377
rect 2361 3345 2401 3377
rect 2433 3345 2462 3377
rect 2210 3305 2462 3345
rect 2210 3273 2257 3305
rect 2289 3273 2329 3305
rect 2361 3273 2401 3305
rect 2433 3273 2462 3305
rect 2210 3233 2462 3273
rect 2210 3201 2257 3233
rect 2289 3201 2329 3233
rect 2361 3201 2401 3233
rect 2433 3201 2462 3233
rect 2210 3161 2462 3201
rect 2210 3129 2257 3161
rect 2289 3129 2329 3161
rect 2361 3129 2401 3161
rect 2433 3129 2462 3161
rect 2210 3089 2462 3129
rect 2210 3057 2257 3089
rect 2289 3057 2329 3089
rect 2361 3057 2401 3089
rect 2433 3057 2462 3089
rect 2210 3017 2462 3057
rect 2210 2985 2257 3017
rect 2289 2985 2329 3017
rect 2361 2985 2401 3017
rect 2433 2985 2462 3017
rect 2210 2945 2462 2985
rect 2210 2913 2257 2945
rect 2289 2913 2329 2945
rect 2361 2913 2401 2945
rect 2433 2913 2462 2945
rect 2210 2873 2462 2913
rect 2210 2841 2257 2873
rect 2289 2841 2329 2873
rect 2361 2841 2401 2873
rect 2433 2841 2462 2873
rect 2210 2801 2462 2841
rect 2210 2769 2257 2801
rect 2289 2769 2329 2801
rect 2361 2769 2401 2801
rect 2433 2769 2462 2801
rect 2210 2729 2462 2769
rect 2210 2697 2257 2729
rect 2289 2697 2329 2729
rect 2361 2697 2401 2729
rect 2433 2697 2462 2729
rect 2210 2657 2462 2697
rect 2210 2625 2257 2657
rect 2289 2625 2329 2657
rect 2361 2625 2401 2657
rect 2433 2625 2462 2657
rect 2210 2585 2462 2625
rect 2210 2553 2257 2585
rect 2289 2553 2329 2585
rect 2361 2553 2401 2585
rect 2433 2553 2462 2585
rect 2210 2513 2462 2553
rect 2210 2481 2257 2513
rect 2289 2481 2329 2513
rect 2361 2481 2401 2513
rect 2433 2481 2462 2513
rect 2210 2441 2462 2481
rect 2210 2409 2257 2441
rect 2289 2409 2329 2441
rect 2361 2409 2401 2441
rect 2433 2409 2462 2441
rect 2210 2369 2462 2409
rect 2210 2337 2257 2369
rect 2289 2337 2329 2369
rect 2361 2337 2401 2369
rect 2433 2337 2462 2369
rect 2210 2297 2462 2337
rect 2210 2265 2257 2297
rect 2289 2265 2329 2297
rect 2361 2265 2401 2297
rect 2433 2265 2462 2297
rect 2210 2225 2462 2265
rect 2210 2193 2257 2225
rect 2289 2193 2329 2225
rect 2361 2193 2401 2225
rect 2433 2193 2462 2225
rect 2210 2153 2462 2193
rect 2210 2121 2257 2153
rect 2289 2121 2329 2153
rect 2361 2121 2401 2153
rect 2433 2121 2462 2153
rect 2210 2081 2462 2121
rect 2210 2049 2257 2081
rect 2289 2049 2329 2081
rect 2361 2049 2401 2081
rect 2433 2049 2462 2081
rect 2210 2009 2462 2049
rect 2210 1977 2257 2009
rect 2289 1977 2329 2009
rect 2361 1977 2401 2009
rect 2433 1977 2462 2009
rect 2210 1937 2462 1977
rect 2210 1905 2257 1937
rect 2289 1905 2329 1937
rect 2361 1905 2401 1937
rect 2433 1905 2462 1937
rect 2210 1865 2462 1905
rect 2210 1833 2257 1865
rect 2289 1833 2329 1865
rect 2361 1833 2401 1865
rect 2433 1833 2462 1865
rect 2210 1793 2462 1833
rect 2210 1761 2257 1793
rect 2289 1761 2329 1793
rect 2361 1761 2401 1793
rect 2433 1761 2462 1793
rect 2210 1721 2462 1761
rect 2210 1689 2257 1721
rect 2289 1689 2329 1721
rect 2361 1689 2401 1721
rect 2433 1689 2462 1721
rect 2210 1649 2462 1689
rect 2210 1617 2257 1649
rect 2289 1617 2329 1649
rect 2361 1617 2401 1649
rect 2433 1617 2462 1649
rect 2210 1577 2462 1617
rect 2210 1545 2257 1577
rect 2289 1545 2329 1577
rect 2361 1545 2401 1577
rect 2433 1545 2462 1577
rect 2210 1505 2462 1545
rect 2210 1473 2257 1505
rect 2289 1473 2329 1505
rect 2361 1473 2401 1505
rect 2433 1473 2462 1505
rect 2210 1433 2462 1473
rect 2210 1401 2257 1433
rect 2289 1401 2329 1433
rect 2361 1401 2401 1433
rect 2433 1401 2462 1433
rect 2210 1361 2462 1401
rect 2210 1329 2257 1361
rect 2289 1329 2329 1361
rect 2361 1329 2401 1361
rect 2433 1329 2462 1361
rect 2210 1289 2462 1329
rect 2210 1257 2257 1289
rect 2289 1257 2329 1289
rect 2361 1257 2401 1289
rect 2433 1257 2462 1289
rect 2210 1217 2462 1257
rect 2210 1185 2257 1217
rect 2289 1185 2329 1217
rect 2361 1185 2401 1217
rect 2433 1185 2462 1217
rect 2210 1145 2462 1185
rect 2210 1113 2257 1145
rect 2289 1113 2329 1145
rect 2361 1113 2401 1145
rect 2433 1113 2462 1145
rect 2210 1073 2462 1113
rect 2210 1041 2257 1073
rect 2289 1041 2329 1073
rect 2361 1041 2401 1073
rect 2433 1041 2462 1073
rect 2210 1001 2462 1041
rect 2210 969 2257 1001
rect 2289 969 2329 1001
rect 2361 969 2401 1001
rect 2433 969 2462 1001
rect 1302 897 1345 929
rect 1377 897 1417 929
rect 1449 897 1489 929
rect 1521 897 1554 929
rect 1302 857 1554 897
rect 1302 825 1345 857
rect 1377 825 1417 857
rect 1449 825 1489 857
rect 1521 825 1554 857
rect 1302 785 1554 825
rect 1302 753 1345 785
rect 1377 753 1417 785
rect 1449 753 1489 785
rect 1521 753 1554 785
rect 1302 713 1554 753
rect 1302 681 1345 713
rect 1377 681 1417 713
rect 1449 681 1489 713
rect 1521 681 1554 713
rect 1302 648 1554 681
rect 2210 929 2462 969
rect 2210 897 2257 929
rect 2289 897 2329 929
rect 2361 897 2401 929
rect 2433 897 2462 929
rect 2210 857 2462 897
rect 2210 825 2257 857
rect 2289 825 2329 857
rect 2361 825 2401 857
rect 2433 825 2462 857
rect 2210 785 2462 825
rect 2210 753 2257 785
rect 2289 753 2329 785
rect 2361 753 2401 785
rect 2433 753 2462 785
rect 2210 713 2462 753
rect 2210 681 2257 713
rect 2289 681 2329 713
rect 2361 681 2401 713
rect 2433 681 2462 713
rect 2210 648 2462 681
rect 396 614 2462 648
rect 396 582 447 614
rect 479 582 519 614
rect 551 582 591 614
rect 623 582 663 614
rect 695 582 735 614
rect 767 582 807 614
rect 839 582 879 614
rect 911 582 951 614
rect 983 582 1023 614
rect 1055 582 1095 614
rect 1127 582 1167 614
rect 1199 582 1239 614
rect 1271 582 1311 614
rect 1343 582 1383 614
rect 1415 582 1455 614
rect 1487 582 1527 614
rect 1559 582 1599 614
rect 1631 582 1671 614
rect 1703 582 1743 614
rect 1775 582 1815 614
rect 1847 582 1887 614
rect 1919 582 1959 614
rect 1991 582 2031 614
rect 2063 582 2103 614
rect 2135 582 2175 614
rect 2207 582 2247 614
rect 2279 582 2319 614
rect 2351 582 2391 614
rect 2423 582 2462 614
rect 396 542 2462 582
rect 396 510 447 542
rect 479 510 519 542
rect 551 510 591 542
rect 623 510 663 542
rect 695 510 735 542
rect 767 510 807 542
rect 839 510 879 542
rect 911 510 951 542
rect 983 510 1023 542
rect 1055 510 1095 542
rect 1127 510 1167 542
rect 1199 510 1239 542
rect 1271 510 1311 542
rect 1343 510 1383 542
rect 1415 510 1455 542
rect 1487 510 1527 542
rect 1559 510 1599 542
rect 1631 510 1671 542
rect 1703 510 1743 542
rect 1775 510 1815 542
rect 1847 510 1887 542
rect 1919 510 1959 542
rect 1991 510 2031 542
rect 2063 510 2103 542
rect 2135 510 2175 542
rect 2207 510 2247 542
rect 2279 510 2319 542
rect 2351 510 2391 542
rect 2423 510 2462 542
rect 396 470 2462 510
rect 396 438 447 470
rect 479 438 519 470
rect 551 438 591 470
rect 623 438 663 470
rect 695 438 735 470
rect 767 438 807 470
rect 839 438 879 470
rect 911 438 951 470
rect 983 438 1023 470
rect 1055 438 1095 470
rect 1127 438 1167 470
rect 1199 438 1239 470
rect 1271 438 1311 470
rect 1343 438 1383 470
rect 1415 438 1455 470
rect 1487 438 1527 470
rect 1559 438 1599 470
rect 1631 438 1671 470
rect 1703 438 1743 470
rect 1775 438 1815 470
rect 1847 438 1887 470
rect 1919 438 1959 470
rect 1991 438 2031 470
rect 2063 438 2103 470
rect 2135 438 2175 470
rect 2207 438 2247 470
rect 2279 438 2319 470
rect 2351 438 2391 470
rect 2423 438 2462 470
rect 396 396 2462 438
<< psubdiffcont >>
rect 124 7256 156 7288
rect 196 7256 228 7288
rect 268 7256 300 7288
rect 340 7256 372 7288
rect 412 7256 444 7288
rect 484 7256 516 7288
rect 556 7256 588 7288
rect 628 7256 660 7288
rect 700 7256 732 7288
rect 772 7256 804 7288
rect 844 7256 876 7288
rect 916 7256 948 7288
rect 988 7256 1020 7288
rect 1060 7256 1092 7288
rect 1132 7256 1164 7288
rect 1204 7256 1236 7288
rect 1276 7256 1308 7288
rect 1348 7256 1380 7288
rect 1420 7256 1452 7288
rect 1492 7256 1524 7288
rect 1564 7256 1596 7288
rect 1636 7256 1668 7288
rect 1708 7256 1740 7288
rect 1780 7256 1812 7288
rect 1852 7256 1884 7288
rect 1924 7256 1956 7288
rect 1996 7256 2028 7288
rect 2068 7256 2100 7288
rect 2140 7256 2172 7288
rect 2212 7256 2244 7288
rect 2284 7256 2316 7288
rect 2356 7256 2388 7288
rect 2428 7256 2460 7288
rect 2500 7256 2532 7288
rect 2572 7256 2604 7288
rect 2644 7256 2676 7288
rect 2716 7256 2748 7288
rect 116 7133 148 7165
rect 116 7061 148 7093
rect 116 6989 148 7021
rect 2708 7133 2740 7165
rect 2708 7061 2740 7093
rect 116 6917 148 6949
rect 116 6845 148 6877
rect 116 6773 148 6805
rect 116 6701 148 6733
rect 116 6629 148 6661
rect 116 6557 148 6589
rect 116 6485 148 6517
rect 116 6413 148 6445
rect 116 6341 148 6373
rect 116 6269 148 6301
rect 116 6197 148 6229
rect 116 6125 148 6157
rect 116 6053 148 6085
rect 116 5981 148 6013
rect 116 5909 148 5941
rect 116 5837 148 5869
rect 116 5765 148 5797
rect 116 5693 148 5725
rect 116 5621 148 5653
rect 116 5549 148 5581
rect 116 5477 148 5509
rect 116 5405 148 5437
rect 116 5333 148 5365
rect 116 5261 148 5293
rect 116 5189 148 5221
rect 116 5117 148 5149
rect 116 5045 148 5077
rect 116 4973 148 5005
rect 116 4901 148 4933
rect 116 4829 148 4861
rect 116 4757 148 4789
rect 116 4685 148 4717
rect 116 4613 148 4645
rect 116 4541 148 4573
rect 116 4469 148 4501
rect 116 4397 148 4429
rect 116 4325 148 4357
rect 116 4253 148 4285
rect 116 4181 148 4213
rect 116 4109 148 4141
rect 116 4037 148 4069
rect 116 3965 148 3997
rect 116 3893 148 3925
rect 116 3821 148 3853
rect 116 3749 148 3781
rect 116 3677 148 3709
rect 116 3605 148 3637
rect 116 3533 148 3565
rect 116 3461 148 3493
rect 116 3389 148 3421
rect 116 3317 148 3349
rect 116 3245 148 3277
rect 116 3173 148 3205
rect 116 3101 148 3133
rect 116 3029 148 3061
rect 116 2957 148 2989
rect 116 2885 148 2917
rect 116 2813 148 2845
rect 116 2741 148 2773
rect 116 2669 148 2701
rect 116 2597 148 2629
rect 116 2525 148 2557
rect 116 2453 148 2485
rect 116 2381 148 2413
rect 116 2309 148 2341
rect 116 2237 148 2269
rect 116 2165 148 2197
rect 116 2093 148 2125
rect 116 2021 148 2053
rect 116 1949 148 1981
rect 116 1877 148 1909
rect 116 1805 148 1837
rect 116 1733 148 1765
rect 116 1661 148 1693
rect 116 1589 148 1621
rect 116 1517 148 1549
rect 116 1445 148 1477
rect 116 1373 148 1405
rect 116 1301 148 1333
rect 116 1229 148 1261
rect 116 1157 148 1189
rect 116 1085 148 1117
rect 116 1013 148 1045
rect 116 941 148 973
rect 116 869 148 901
rect 116 797 148 829
rect 116 725 148 757
rect 116 653 148 685
rect 116 581 148 613
rect 116 509 148 541
rect 116 437 148 469
rect 116 365 148 397
rect 2708 6989 2740 7021
rect 2708 6917 2740 6949
rect 2708 6845 2740 6877
rect 2708 6773 2740 6805
rect 2708 6701 2740 6733
rect 2708 6629 2740 6661
rect 2708 6557 2740 6589
rect 2708 6485 2740 6517
rect 2708 6413 2740 6445
rect 2708 6341 2740 6373
rect 2708 6269 2740 6301
rect 2708 6197 2740 6229
rect 2708 6125 2740 6157
rect 2708 6053 2740 6085
rect 2708 5981 2740 6013
rect 2708 5909 2740 5941
rect 2708 5837 2740 5869
rect 2708 5765 2740 5797
rect 2708 5693 2740 5725
rect 2708 5621 2740 5653
rect 2708 5549 2740 5581
rect 2708 5477 2740 5509
rect 2708 5405 2740 5437
rect 2708 5333 2740 5365
rect 2708 5261 2740 5293
rect 2708 5189 2740 5221
rect 2708 5117 2740 5149
rect 2708 5045 2740 5077
rect 2708 4973 2740 5005
rect 2708 4901 2740 4933
rect 2708 4829 2740 4861
rect 2708 4757 2740 4789
rect 2708 4685 2740 4717
rect 2708 4613 2740 4645
rect 2708 4541 2740 4573
rect 2708 4469 2740 4501
rect 2708 4397 2740 4429
rect 2708 4325 2740 4357
rect 2708 4253 2740 4285
rect 2708 4181 2740 4213
rect 2708 4109 2740 4141
rect 2708 4037 2740 4069
rect 2708 3965 2740 3997
rect 2708 3893 2740 3925
rect 2708 3821 2740 3853
rect 2708 3749 2740 3781
rect 2708 3677 2740 3709
rect 2708 3605 2740 3637
rect 2708 3533 2740 3565
rect 2708 3461 2740 3493
rect 2708 3389 2740 3421
rect 2708 3317 2740 3349
rect 2708 3245 2740 3277
rect 2708 3173 2740 3205
rect 2708 3101 2740 3133
rect 2708 3029 2740 3061
rect 2708 2957 2740 2989
rect 2708 2885 2740 2917
rect 2708 2813 2740 2845
rect 2708 2741 2740 2773
rect 2708 2669 2740 2701
rect 2708 2597 2740 2629
rect 2708 2525 2740 2557
rect 2708 2453 2740 2485
rect 2708 2381 2740 2413
rect 2708 2309 2740 2341
rect 2708 2237 2740 2269
rect 2708 2165 2740 2197
rect 2708 2093 2740 2125
rect 2708 2021 2740 2053
rect 2708 1949 2740 1981
rect 2708 1877 2740 1909
rect 2708 1805 2740 1837
rect 2708 1733 2740 1765
rect 2708 1661 2740 1693
rect 2708 1589 2740 1621
rect 2708 1517 2740 1549
rect 2708 1445 2740 1477
rect 2708 1373 2740 1405
rect 2708 1301 2740 1333
rect 2708 1229 2740 1261
rect 2708 1157 2740 1189
rect 2708 1085 2740 1117
rect 2708 1013 2740 1045
rect 2708 941 2740 973
rect 2708 869 2740 901
rect 2708 797 2740 829
rect 2708 725 2740 757
rect 2708 653 2740 685
rect 2708 581 2740 613
rect 2708 509 2740 541
rect 2708 437 2740 469
rect 116 293 148 325
rect 116 221 148 253
rect 2708 365 2740 397
rect 2708 293 2740 325
rect 2708 221 2740 253
rect 124 122 156 154
rect 196 122 228 154
rect 268 122 300 154
rect 340 122 372 154
rect 412 122 444 154
rect 484 122 516 154
rect 556 122 588 154
rect 628 122 660 154
rect 700 122 732 154
rect 772 122 804 154
rect 844 122 876 154
rect 916 122 948 154
rect 988 122 1020 154
rect 1060 122 1092 154
rect 1132 122 1164 154
rect 1204 122 1236 154
rect 1276 122 1308 154
rect 1348 122 1380 154
rect 1420 122 1452 154
rect 1492 122 1524 154
rect 1564 122 1596 154
rect 1636 122 1668 154
rect 1708 122 1740 154
rect 1780 122 1812 154
rect 1852 122 1884 154
rect 1924 122 1956 154
rect 1996 122 2028 154
rect 2068 122 2100 154
rect 2140 122 2172 154
rect 2212 122 2244 154
rect 2284 122 2316 154
rect 2356 122 2388 154
rect 2428 122 2460 154
rect 2500 122 2532 154
rect 2572 122 2604 154
rect 2644 122 2676 154
rect 2716 122 2748 154
<< nsubdiffcont >>
rect 447 6948 479 6980
rect 519 6948 551 6980
rect 591 6948 623 6980
rect 663 6948 695 6980
rect 735 6948 767 6980
rect 807 6948 839 6980
rect 879 6948 911 6980
rect 951 6948 983 6980
rect 1023 6948 1055 6980
rect 1095 6948 1127 6980
rect 1167 6948 1199 6980
rect 1239 6948 1271 6980
rect 1311 6948 1343 6980
rect 1383 6948 1415 6980
rect 1455 6948 1487 6980
rect 1527 6948 1559 6980
rect 1599 6948 1631 6980
rect 1671 6948 1703 6980
rect 1743 6948 1775 6980
rect 1815 6948 1847 6980
rect 1887 6948 1919 6980
rect 1959 6948 1991 6980
rect 2031 6948 2063 6980
rect 2103 6948 2135 6980
rect 2175 6948 2207 6980
rect 2247 6948 2279 6980
rect 2319 6948 2351 6980
rect 2391 6948 2423 6980
rect 447 6876 479 6908
rect 519 6876 551 6908
rect 591 6876 623 6908
rect 663 6876 695 6908
rect 735 6876 767 6908
rect 807 6876 839 6908
rect 879 6876 911 6908
rect 951 6876 983 6908
rect 1023 6876 1055 6908
rect 1095 6876 1127 6908
rect 1167 6876 1199 6908
rect 1239 6876 1271 6908
rect 1311 6876 1343 6908
rect 1383 6876 1415 6908
rect 1455 6876 1487 6908
rect 1527 6876 1559 6908
rect 1599 6876 1631 6908
rect 1671 6876 1703 6908
rect 1743 6876 1775 6908
rect 1815 6876 1847 6908
rect 1887 6876 1919 6908
rect 1959 6876 1991 6908
rect 2031 6876 2063 6908
rect 2103 6876 2135 6908
rect 2175 6876 2207 6908
rect 2247 6876 2279 6908
rect 2319 6876 2351 6908
rect 2391 6876 2423 6908
rect 447 6804 479 6836
rect 519 6804 551 6836
rect 591 6804 623 6836
rect 663 6804 695 6836
rect 735 6804 767 6836
rect 807 6804 839 6836
rect 879 6804 911 6836
rect 951 6804 983 6836
rect 1023 6804 1055 6836
rect 1095 6804 1127 6836
rect 1167 6804 1199 6836
rect 1239 6804 1271 6836
rect 1311 6804 1343 6836
rect 1383 6804 1415 6836
rect 1455 6804 1487 6836
rect 1527 6804 1559 6836
rect 1599 6804 1631 6836
rect 1671 6804 1703 6836
rect 1743 6804 1775 6836
rect 1815 6804 1847 6836
rect 1887 6804 1919 6836
rect 1959 6804 1991 6836
rect 2031 6804 2063 6836
rect 2103 6804 2135 6836
rect 2175 6804 2207 6836
rect 2247 6804 2279 6836
rect 2319 6804 2351 6836
rect 2391 6804 2423 6836
rect 433 6729 465 6761
rect 505 6729 537 6761
rect 577 6729 609 6761
rect 433 6657 465 6689
rect 505 6657 537 6689
rect 577 6657 609 6689
rect 433 6585 465 6617
rect 505 6585 537 6617
rect 577 6585 609 6617
rect 433 6513 465 6545
rect 505 6513 537 6545
rect 577 6513 609 6545
rect 1345 6729 1377 6761
rect 1417 6729 1449 6761
rect 1489 6729 1521 6761
rect 1345 6657 1377 6689
rect 1417 6657 1449 6689
rect 1489 6657 1521 6689
rect 1345 6585 1377 6617
rect 1417 6585 1449 6617
rect 1489 6585 1521 6617
rect 1345 6513 1377 6545
rect 1417 6513 1449 6545
rect 1489 6513 1521 6545
rect 433 6441 465 6473
rect 505 6441 537 6473
rect 577 6441 609 6473
rect 433 6369 465 6401
rect 505 6369 537 6401
rect 577 6369 609 6401
rect 433 6297 465 6329
rect 505 6297 537 6329
rect 577 6297 609 6329
rect 433 6225 465 6257
rect 505 6225 537 6257
rect 577 6225 609 6257
rect 433 6153 465 6185
rect 505 6153 537 6185
rect 577 6153 609 6185
rect 433 6081 465 6113
rect 505 6081 537 6113
rect 577 6081 609 6113
rect 433 6009 465 6041
rect 505 6009 537 6041
rect 577 6009 609 6041
rect 433 5937 465 5969
rect 505 5937 537 5969
rect 577 5937 609 5969
rect 433 5865 465 5897
rect 505 5865 537 5897
rect 577 5865 609 5897
rect 433 5793 465 5825
rect 505 5793 537 5825
rect 577 5793 609 5825
rect 433 5721 465 5753
rect 505 5721 537 5753
rect 577 5721 609 5753
rect 433 5649 465 5681
rect 505 5649 537 5681
rect 577 5649 609 5681
rect 433 5577 465 5609
rect 505 5577 537 5609
rect 577 5577 609 5609
rect 433 5505 465 5537
rect 505 5505 537 5537
rect 577 5505 609 5537
rect 433 5433 465 5465
rect 505 5433 537 5465
rect 577 5433 609 5465
rect 433 5361 465 5393
rect 505 5361 537 5393
rect 577 5361 609 5393
rect 433 5289 465 5321
rect 505 5289 537 5321
rect 577 5289 609 5321
rect 433 5217 465 5249
rect 505 5217 537 5249
rect 577 5217 609 5249
rect 433 5145 465 5177
rect 505 5145 537 5177
rect 577 5145 609 5177
rect 433 5073 465 5105
rect 505 5073 537 5105
rect 577 5073 609 5105
rect 433 5001 465 5033
rect 505 5001 537 5033
rect 577 5001 609 5033
rect 433 4929 465 4961
rect 505 4929 537 4961
rect 577 4929 609 4961
rect 433 4857 465 4889
rect 505 4857 537 4889
rect 577 4857 609 4889
rect 433 4785 465 4817
rect 505 4785 537 4817
rect 577 4785 609 4817
rect 433 4713 465 4745
rect 505 4713 537 4745
rect 577 4713 609 4745
rect 433 4641 465 4673
rect 505 4641 537 4673
rect 577 4641 609 4673
rect 433 4569 465 4601
rect 505 4569 537 4601
rect 577 4569 609 4601
rect 433 4497 465 4529
rect 505 4497 537 4529
rect 577 4497 609 4529
rect 433 4425 465 4457
rect 505 4425 537 4457
rect 577 4425 609 4457
rect 433 4353 465 4385
rect 505 4353 537 4385
rect 577 4353 609 4385
rect 433 4281 465 4313
rect 505 4281 537 4313
rect 577 4281 609 4313
rect 433 4209 465 4241
rect 505 4209 537 4241
rect 577 4209 609 4241
rect 433 4137 465 4169
rect 505 4137 537 4169
rect 577 4137 609 4169
rect 433 4065 465 4097
rect 505 4065 537 4097
rect 577 4065 609 4097
rect 433 3993 465 4025
rect 505 3993 537 4025
rect 577 3993 609 4025
rect 433 3921 465 3953
rect 505 3921 537 3953
rect 577 3921 609 3953
rect 433 3849 465 3881
rect 505 3849 537 3881
rect 577 3849 609 3881
rect 433 3777 465 3809
rect 505 3777 537 3809
rect 577 3777 609 3809
rect 433 3705 465 3737
rect 505 3705 537 3737
rect 577 3705 609 3737
rect 433 3633 465 3665
rect 505 3633 537 3665
rect 577 3633 609 3665
rect 433 3561 465 3593
rect 505 3561 537 3593
rect 577 3561 609 3593
rect 433 3489 465 3521
rect 505 3489 537 3521
rect 577 3489 609 3521
rect 433 3417 465 3449
rect 505 3417 537 3449
rect 577 3417 609 3449
rect 433 3345 465 3377
rect 505 3345 537 3377
rect 577 3345 609 3377
rect 433 3273 465 3305
rect 505 3273 537 3305
rect 577 3273 609 3305
rect 433 3201 465 3233
rect 505 3201 537 3233
rect 577 3201 609 3233
rect 433 3129 465 3161
rect 505 3129 537 3161
rect 577 3129 609 3161
rect 433 3057 465 3089
rect 505 3057 537 3089
rect 577 3057 609 3089
rect 433 2985 465 3017
rect 505 2985 537 3017
rect 577 2985 609 3017
rect 433 2913 465 2945
rect 505 2913 537 2945
rect 577 2913 609 2945
rect 433 2841 465 2873
rect 505 2841 537 2873
rect 577 2841 609 2873
rect 433 2769 465 2801
rect 505 2769 537 2801
rect 577 2769 609 2801
rect 433 2697 465 2729
rect 505 2697 537 2729
rect 577 2697 609 2729
rect 433 2625 465 2657
rect 505 2625 537 2657
rect 577 2625 609 2657
rect 433 2553 465 2585
rect 505 2553 537 2585
rect 577 2553 609 2585
rect 433 2481 465 2513
rect 505 2481 537 2513
rect 577 2481 609 2513
rect 433 2409 465 2441
rect 505 2409 537 2441
rect 577 2409 609 2441
rect 433 2337 465 2369
rect 505 2337 537 2369
rect 577 2337 609 2369
rect 433 2265 465 2297
rect 505 2265 537 2297
rect 577 2265 609 2297
rect 433 2193 465 2225
rect 505 2193 537 2225
rect 577 2193 609 2225
rect 433 2121 465 2153
rect 505 2121 537 2153
rect 577 2121 609 2153
rect 433 2049 465 2081
rect 505 2049 537 2081
rect 577 2049 609 2081
rect 433 1977 465 2009
rect 505 1977 537 2009
rect 577 1977 609 2009
rect 433 1905 465 1937
rect 505 1905 537 1937
rect 577 1905 609 1937
rect 433 1833 465 1865
rect 505 1833 537 1865
rect 577 1833 609 1865
rect 433 1761 465 1793
rect 505 1761 537 1793
rect 577 1761 609 1793
rect 433 1689 465 1721
rect 505 1689 537 1721
rect 577 1689 609 1721
rect 433 1617 465 1649
rect 505 1617 537 1649
rect 577 1617 609 1649
rect 433 1545 465 1577
rect 505 1545 537 1577
rect 577 1545 609 1577
rect 433 1473 465 1505
rect 505 1473 537 1505
rect 577 1473 609 1505
rect 433 1401 465 1433
rect 505 1401 537 1433
rect 577 1401 609 1433
rect 433 1329 465 1361
rect 505 1329 537 1361
rect 577 1329 609 1361
rect 433 1257 465 1289
rect 505 1257 537 1289
rect 577 1257 609 1289
rect 433 1185 465 1217
rect 505 1185 537 1217
rect 577 1185 609 1217
rect 433 1113 465 1145
rect 505 1113 537 1145
rect 577 1113 609 1145
rect 433 1041 465 1073
rect 505 1041 537 1073
rect 577 1041 609 1073
rect 433 969 465 1001
rect 505 969 537 1001
rect 577 969 609 1001
rect 2257 6729 2289 6761
rect 2329 6729 2361 6761
rect 2401 6729 2433 6761
rect 2257 6657 2289 6689
rect 2329 6657 2361 6689
rect 2401 6657 2433 6689
rect 2257 6585 2289 6617
rect 2329 6585 2361 6617
rect 2401 6585 2433 6617
rect 2257 6513 2289 6545
rect 2329 6513 2361 6545
rect 2401 6513 2433 6545
rect 1345 6441 1377 6473
rect 1417 6441 1449 6473
rect 1489 6441 1521 6473
rect 1345 6369 1377 6401
rect 1417 6369 1449 6401
rect 1489 6369 1521 6401
rect 1345 6297 1377 6329
rect 1417 6297 1449 6329
rect 1489 6297 1521 6329
rect 1345 6225 1377 6257
rect 1417 6225 1449 6257
rect 1489 6225 1521 6257
rect 1345 6153 1377 6185
rect 1417 6153 1449 6185
rect 1489 6153 1521 6185
rect 1345 6081 1377 6113
rect 1417 6081 1449 6113
rect 1489 6081 1521 6113
rect 1345 6009 1377 6041
rect 1417 6009 1449 6041
rect 1489 6009 1521 6041
rect 1345 5937 1377 5969
rect 1417 5937 1449 5969
rect 1489 5937 1521 5969
rect 1345 5865 1377 5897
rect 1417 5865 1449 5897
rect 1489 5865 1521 5897
rect 1345 5793 1377 5825
rect 1417 5793 1449 5825
rect 1489 5793 1521 5825
rect 1345 5721 1377 5753
rect 1417 5721 1449 5753
rect 1489 5721 1521 5753
rect 1345 5649 1377 5681
rect 1417 5649 1449 5681
rect 1489 5649 1521 5681
rect 1345 5577 1377 5609
rect 1417 5577 1449 5609
rect 1489 5577 1521 5609
rect 1345 5505 1377 5537
rect 1417 5505 1449 5537
rect 1489 5505 1521 5537
rect 1345 5433 1377 5465
rect 1417 5433 1449 5465
rect 1489 5433 1521 5465
rect 1345 5361 1377 5393
rect 1417 5361 1449 5393
rect 1489 5361 1521 5393
rect 1345 5289 1377 5321
rect 1417 5289 1449 5321
rect 1489 5289 1521 5321
rect 1345 5217 1377 5249
rect 1417 5217 1449 5249
rect 1489 5217 1521 5249
rect 1345 5145 1377 5177
rect 1417 5145 1449 5177
rect 1489 5145 1521 5177
rect 1345 5073 1377 5105
rect 1417 5073 1449 5105
rect 1489 5073 1521 5105
rect 1345 5001 1377 5033
rect 1417 5001 1449 5033
rect 1489 5001 1521 5033
rect 1345 4929 1377 4961
rect 1417 4929 1449 4961
rect 1489 4929 1521 4961
rect 1345 4857 1377 4889
rect 1417 4857 1449 4889
rect 1489 4857 1521 4889
rect 1345 4785 1377 4817
rect 1417 4785 1449 4817
rect 1489 4785 1521 4817
rect 1345 4713 1377 4745
rect 1417 4713 1449 4745
rect 1489 4713 1521 4745
rect 1345 4641 1377 4673
rect 1417 4641 1449 4673
rect 1489 4641 1521 4673
rect 1345 4569 1377 4601
rect 1417 4569 1449 4601
rect 1489 4569 1521 4601
rect 1345 4497 1377 4529
rect 1417 4497 1449 4529
rect 1489 4497 1521 4529
rect 1345 4425 1377 4457
rect 1417 4425 1449 4457
rect 1489 4425 1521 4457
rect 1345 4353 1377 4385
rect 1417 4353 1449 4385
rect 1489 4353 1521 4385
rect 1345 4281 1377 4313
rect 1417 4281 1449 4313
rect 1489 4281 1521 4313
rect 1345 4209 1377 4241
rect 1417 4209 1449 4241
rect 1489 4209 1521 4241
rect 1345 4137 1377 4169
rect 1417 4137 1449 4169
rect 1489 4137 1521 4169
rect 1345 4065 1377 4097
rect 1417 4065 1449 4097
rect 1489 4065 1521 4097
rect 1345 3993 1377 4025
rect 1417 3993 1449 4025
rect 1489 3993 1521 4025
rect 1345 3921 1377 3953
rect 1417 3921 1449 3953
rect 1489 3921 1521 3953
rect 1345 3849 1377 3881
rect 1417 3849 1449 3881
rect 1489 3849 1521 3881
rect 1345 3777 1377 3809
rect 1417 3777 1449 3809
rect 1489 3777 1521 3809
rect 1345 3705 1377 3737
rect 1417 3705 1449 3737
rect 1489 3705 1521 3737
rect 1345 3633 1377 3665
rect 1417 3633 1449 3665
rect 1489 3633 1521 3665
rect 1345 3561 1377 3593
rect 1417 3561 1449 3593
rect 1489 3561 1521 3593
rect 1345 3489 1377 3521
rect 1417 3489 1449 3521
rect 1489 3489 1521 3521
rect 1345 3417 1377 3449
rect 1417 3417 1449 3449
rect 1489 3417 1521 3449
rect 1345 3345 1377 3377
rect 1417 3345 1449 3377
rect 1489 3345 1521 3377
rect 1345 3273 1377 3305
rect 1417 3273 1449 3305
rect 1489 3273 1521 3305
rect 1345 3201 1377 3233
rect 1417 3201 1449 3233
rect 1489 3201 1521 3233
rect 1345 3129 1377 3161
rect 1417 3129 1449 3161
rect 1489 3129 1521 3161
rect 1345 3057 1377 3089
rect 1417 3057 1449 3089
rect 1489 3057 1521 3089
rect 1345 2985 1377 3017
rect 1417 2985 1449 3017
rect 1489 2985 1521 3017
rect 1345 2913 1377 2945
rect 1417 2913 1449 2945
rect 1489 2913 1521 2945
rect 1345 2841 1377 2873
rect 1417 2841 1449 2873
rect 1489 2841 1521 2873
rect 1345 2769 1377 2801
rect 1417 2769 1449 2801
rect 1489 2769 1521 2801
rect 1345 2697 1377 2729
rect 1417 2697 1449 2729
rect 1489 2697 1521 2729
rect 1345 2625 1377 2657
rect 1417 2625 1449 2657
rect 1489 2625 1521 2657
rect 1345 2553 1377 2585
rect 1417 2553 1449 2585
rect 1489 2553 1521 2585
rect 1345 2481 1377 2513
rect 1417 2481 1449 2513
rect 1489 2481 1521 2513
rect 1345 2409 1377 2441
rect 1417 2409 1449 2441
rect 1489 2409 1521 2441
rect 1345 2337 1377 2369
rect 1417 2337 1449 2369
rect 1489 2337 1521 2369
rect 1345 2265 1377 2297
rect 1417 2265 1449 2297
rect 1489 2265 1521 2297
rect 1345 2193 1377 2225
rect 1417 2193 1449 2225
rect 1489 2193 1521 2225
rect 1345 2121 1377 2153
rect 1417 2121 1449 2153
rect 1489 2121 1521 2153
rect 1345 2049 1377 2081
rect 1417 2049 1449 2081
rect 1489 2049 1521 2081
rect 1345 1977 1377 2009
rect 1417 1977 1449 2009
rect 1489 1977 1521 2009
rect 1345 1905 1377 1937
rect 1417 1905 1449 1937
rect 1489 1905 1521 1937
rect 1345 1833 1377 1865
rect 1417 1833 1449 1865
rect 1489 1833 1521 1865
rect 1345 1761 1377 1793
rect 1417 1761 1449 1793
rect 1489 1761 1521 1793
rect 1345 1689 1377 1721
rect 1417 1689 1449 1721
rect 1489 1689 1521 1721
rect 1345 1617 1377 1649
rect 1417 1617 1449 1649
rect 1489 1617 1521 1649
rect 1345 1545 1377 1577
rect 1417 1545 1449 1577
rect 1489 1545 1521 1577
rect 1345 1473 1377 1505
rect 1417 1473 1449 1505
rect 1489 1473 1521 1505
rect 1345 1401 1377 1433
rect 1417 1401 1449 1433
rect 1489 1401 1521 1433
rect 1345 1329 1377 1361
rect 1417 1329 1449 1361
rect 1489 1329 1521 1361
rect 1345 1257 1377 1289
rect 1417 1257 1449 1289
rect 1489 1257 1521 1289
rect 1345 1185 1377 1217
rect 1417 1185 1449 1217
rect 1489 1185 1521 1217
rect 1345 1113 1377 1145
rect 1417 1113 1449 1145
rect 1489 1113 1521 1145
rect 1345 1041 1377 1073
rect 1417 1041 1449 1073
rect 1489 1041 1521 1073
rect 1345 969 1377 1001
rect 1417 969 1449 1001
rect 1489 969 1521 1001
rect 433 897 465 929
rect 505 897 537 929
rect 577 897 609 929
rect 433 825 465 857
rect 505 825 537 857
rect 577 825 609 857
rect 433 753 465 785
rect 505 753 537 785
rect 577 753 609 785
rect 433 681 465 713
rect 505 681 537 713
rect 577 681 609 713
rect 2257 6441 2289 6473
rect 2329 6441 2361 6473
rect 2401 6441 2433 6473
rect 2257 6369 2289 6401
rect 2329 6369 2361 6401
rect 2401 6369 2433 6401
rect 2257 6297 2289 6329
rect 2329 6297 2361 6329
rect 2401 6297 2433 6329
rect 2257 6225 2289 6257
rect 2329 6225 2361 6257
rect 2401 6225 2433 6257
rect 2257 6153 2289 6185
rect 2329 6153 2361 6185
rect 2401 6153 2433 6185
rect 2257 6081 2289 6113
rect 2329 6081 2361 6113
rect 2401 6081 2433 6113
rect 2257 6009 2289 6041
rect 2329 6009 2361 6041
rect 2401 6009 2433 6041
rect 2257 5937 2289 5969
rect 2329 5937 2361 5969
rect 2401 5937 2433 5969
rect 2257 5865 2289 5897
rect 2329 5865 2361 5897
rect 2401 5865 2433 5897
rect 2257 5793 2289 5825
rect 2329 5793 2361 5825
rect 2401 5793 2433 5825
rect 2257 5721 2289 5753
rect 2329 5721 2361 5753
rect 2401 5721 2433 5753
rect 2257 5649 2289 5681
rect 2329 5649 2361 5681
rect 2401 5649 2433 5681
rect 2257 5577 2289 5609
rect 2329 5577 2361 5609
rect 2401 5577 2433 5609
rect 2257 5505 2289 5537
rect 2329 5505 2361 5537
rect 2401 5505 2433 5537
rect 2257 5433 2289 5465
rect 2329 5433 2361 5465
rect 2401 5433 2433 5465
rect 2257 5361 2289 5393
rect 2329 5361 2361 5393
rect 2401 5361 2433 5393
rect 2257 5289 2289 5321
rect 2329 5289 2361 5321
rect 2401 5289 2433 5321
rect 2257 5217 2289 5249
rect 2329 5217 2361 5249
rect 2401 5217 2433 5249
rect 2257 5145 2289 5177
rect 2329 5145 2361 5177
rect 2401 5145 2433 5177
rect 2257 5073 2289 5105
rect 2329 5073 2361 5105
rect 2401 5073 2433 5105
rect 2257 5001 2289 5033
rect 2329 5001 2361 5033
rect 2401 5001 2433 5033
rect 2257 4929 2289 4961
rect 2329 4929 2361 4961
rect 2401 4929 2433 4961
rect 2257 4857 2289 4889
rect 2329 4857 2361 4889
rect 2401 4857 2433 4889
rect 2257 4785 2289 4817
rect 2329 4785 2361 4817
rect 2401 4785 2433 4817
rect 2257 4713 2289 4745
rect 2329 4713 2361 4745
rect 2401 4713 2433 4745
rect 2257 4641 2289 4673
rect 2329 4641 2361 4673
rect 2401 4641 2433 4673
rect 2257 4569 2289 4601
rect 2329 4569 2361 4601
rect 2401 4569 2433 4601
rect 2257 4497 2289 4529
rect 2329 4497 2361 4529
rect 2401 4497 2433 4529
rect 2257 4425 2289 4457
rect 2329 4425 2361 4457
rect 2401 4425 2433 4457
rect 2257 4353 2289 4385
rect 2329 4353 2361 4385
rect 2401 4353 2433 4385
rect 2257 4281 2289 4313
rect 2329 4281 2361 4313
rect 2401 4281 2433 4313
rect 2257 4209 2289 4241
rect 2329 4209 2361 4241
rect 2401 4209 2433 4241
rect 2257 4137 2289 4169
rect 2329 4137 2361 4169
rect 2401 4137 2433 4169
rect 2257 4065 2289 4097
rect 2329 4065 2361 4097
rect 2401 4065 2433 4097
rect 2257 3993 2289 4025
rect 2329 3993 2361 4025
rect 2401 3993 2433 4025
rect 2257 3921 2289 3953
rect 2329 3921 2361 3953
rect 2401 3921 2433 3953
rect 2257 3849 2289 3881
rect 2329 3849 2361 3881
rect 2401 3849 2433 3881
rect 2257 3777 2289 3809
rect 2329 3777 2361 3809
rect 2401 3777 2433 3809
rect 2257 3705 2289 3737
rect 2329 3705 2361 3737
rect 2401 3705 2433 3737
rect 2257 3633 2289 3665
rect 2329 3633 2361 3665
rect 2401 3633 2433 3665
rect 2257 3561 2289 3593
rect 2329 3561 2361 3593
rect 2401 3561 2433 3593
rect 2257 3489 2289 3521
rect 2329 3489 2361 3521
rect 2401 3489 2433 3521
rect 2257 3417 2289 3449
rect 2329 3417 2361 3449
rect 2401 3417 2433 3449
rect 2257 3345 2289 3377
rect 2329 3345 2361 3377
rect 2401 3345 2433 3377
rect 2257 3273 2289 3305
rect 2329 3273 2361 3305
rect 2401 3273 2433 3305
rect 2257 3201 2289 3233
rect 2329 3201 2361 3233
rect 2401 3201 2433 3233
rect 2257 3129 2289 3161
rect 2329 3129 2361 3161
rect 2401 3129 2433 3161
rect 2257 3057 2289 3089
rect 2329 3057 2361 3089
rect 2401 3057 2433 3089
rect 2257 2985 2289 3017
rect 2329 2985 2361 3017
rect 2401 2985 2433 3017
rect 2257 2913 2289 2945
rect 2329 2913 2361 2945
rect 2401 2913 2433 2945
rect 2257 2841 2289 2873
rect 2329 2841 2361 2873
rect 2401 2841 2433 2873
rect 2257 2769 2289 2801
rect 2329 2769 2361 2801
rect 2401 2769 2433 2801
rect 2257 2697 2289 2729
rect 2329 2697 2361 2729
rect 2401 2697 2433 2729
rect 2257 2625 2289 2657
rect 2329 2625 2361 2657
rect 2401 2625 2433 2657
rect 2257 2553 2289 2585
rect 2329 2553 2361 2585
rect 2401 2553 2433 2585
rect 2257 2481 2289 2513
rect 2329 2481 2361 2513
rect 2401 2481 2433 2513
rect 2257 2409 2289 2441
rect 2329 2409 2361 2441
rect 2401 2409 2433 2441
rect 2257 2337 2289 2369
rect 2329 2337 2361 2369
rect 2401 2337 2433 2369
rect 2257 2265 2289 2297
rect 2329 2265 2361 2297
rect 2401 2265 2433 2297
rect 2257 2193 2289 2225
rect 2329 2193 2361 2225
rect 2401 2193 2433 2225
rect 2257 2121 2289 2153
rect 2329 2121 2361 2153
rect 2401 2121 2433 2153
rect 2257 2049 2289 2081
rect 2329 2049 2361 2081
rect 2401 2049 2433 2081
rect 2257 1977 2289 2009
rect 2329 1977 2361 2009
rect 2401 1977 2433 2009
rect 2257 1905 2289 1937
rect 2329 1905 2361 1937
rect 2401 1905 2433 1937
rect 2257 1833 2289 1865
rect 2329 1833 2361 1865
rect 2401 1833 2433 1865
rect 2257 1761 2289 1793
rect 2329 1761 2361 1793
rect 2401 1761 2433 1793
rect 2257 1689 2289 1721
rect 2329 1689 2361 1721
rect 2401 1689 2433 1721
rect 2257 1617 2289 1649
rect 2329 1617 2361 1649
rect 2401 1617 2433 1649
rect 2257 1545 2289 1577
rect 2329 1545 2361 1577
rect 2401 1545 2433 1577
rect 2257 1473 2289 1505
rect 2329 1473 2361 1505
rect 2401 1473 2433 1505
rect 2257 1401 2289 1433
rect 2329 1401 2361 1433
rect 2401 1401 2433 1433
rect 2257 1329 2289 1361
rect 2329 1329 2361 1361
rect 2401 1329 2433 1361
rect 2257 1257 2289 1289
rect 2329 1257 2361 1289
rect 2401 1257 2433 1289
rect 2257 1185 2289 1217
rect 2329 1185 2361 1217
rect 2401 1185 2433 1217
rect 2257 1113 2289 1145
rect 2329 1113 2361 1145
rect 2401 1113 2433 1145
rect 2257 1041 2289 1073
rect 2329 1041 2361 1073
rect 2401 1041 2433 1073
rect 2257 969 2289 1001
rect 2329 969 2361 1001
rect 2401 969 2433 1001
rect 1345 897 1377 929
rect 1417 897 1449 929
rect 1489 897 1521 929
rect 1345 825 1377 857
rect 1417 825 1449 857
rect 1489 825 1521 857
rect 1345 753 1377 785
rect 1417 753 1449 785
rect 1489 753 1521 785
rect 1345 681 1377 713
rect 1417 681 1449 713
rect 1489 681 1521 713
rect 2257 897 2289 929
rect 2329 897 2361 929
rect 2401 897 2433 929
rect 2257 825 2289 857
rect 2329 825 2361 857
rect 2401 825 2433 857
rect 2257 753 2289 785
rect 2329 753 2361 785
rect 2401 753 2433 785
rect 2257 681 2289 713
rect 2329 681 2361 713
rect 2401 681 2433 713
rect 447 582 479 614
rect 519 582 551 614
rect 591 582 623 614
rect 663 582 695 614
rect 735 582 767 614
rect 807 582 839 614
rect 879 582 911 614
rect 951 582 983 614
rect 1023 582 1055 614
rect 1095 582 1127 614
rect 1167 582 1199 614
rect 1239 582 1271 614
rect 1311 582 1343 614
rect 1383 582 1415 614
rect 1455 582 1487 614
rect 1527 582 1559 614
rect 1599 582 1631 614
rect 1671 582 1703 614
rect 1743 582 1775 614
rect 1815 582 1847 614
rect 1887 582 1919 614
rect 1959 582 1991 614
rect 2031 582 2063 614
rect 2103 582 2135 614
rect 2175 582 2207 614
rect 2247 582 2279 614
rect 2319 582 2351 614
rect 2391 582 2423 614
rect 447 510 479 542
rect 519 510 551 542
rect 591 510 623 542
rect 663 510 695 542
rect 735 510 767 542
rect 807 510 839 542
rect 879 510 911 542
rect 951 510 983 542
rect 1023 510 1055 542
rect 1095 510 1127 542
rect 1167 510 1199 542
rect 1239 510 1271 542
rect 1311 510 1343 542
rect 1383 510 1415 542
rect 1455 510 1487 542
rect 1527 510 1559 542
rect 1599 510 1631 542
rect 1671 510 1703 542
rect 1743 510 1775 542
rect 1815 510 1847 542
rect 1887 510 1919 542
rect 1959 510 1991 542
rect 2031 510 2063 542
rect 2103 510 2135 542
rect 2175 510 2207 542
rect 2247 510 2279 542
rect 2319 510 2351 542
rect 2391 510 2423 542
rect 447 438 479 470
rect 519 438 551 470
rect 591 438 623 470
rect 663 438 695 470
rect 735 438 767 470
rect 807 438 839 470
rect 879 438 911 470
rect 951 438 983 470
rect 1023 438 1055 470
rect 1095 438 1127 470
rect 1167 438 1199 470
rect 1239 438 1271 470
rect 1311 438 1343 470
rect 1383 438 1415 470
rect 1455 438 1487 470
rect 1527 438 1559 470
rect 1599 438 1631 470
rect 1671 438 1703 470
rect 1743 438 1775 470
rect 1815 438 1847 470
rect 1887 438 1919 470
rect 1959 438 1991 470
rect 2031 438 2063 470
rect 2103 438 2135 470
rect 2175 438 2207 470
rect 2247 438 2279 470
rect 2319 438 2351 470
rect 2391 438 2423 470
<< metal1 >>
rect 0 7288 2864 7410
rect 0 7256 124 7288
rect 156 7256 196 7288
rect 228 7256 268 7288
rect 300 7256 340 7288
rect 372 7256 412 7288
rect 444 7256 484 7288
rect 516 7256 556 7288
rect 588 7256 628 7288
rect 660 7256 700 7288
rect 732 7256 772 7288
rect 804 7256 844 7288
rect 876 7256 916 7288
rect 948 7256 988 7288
rect 1020 7256 1060 7288
rect 1092 7256 1132 7288
rect 1164 7256 1204 7288
rect 1236 7256 1276 7288
rect 1308 7256 1348 7288
rect 1380 7256 1420 7288
rect 1452 7256 1492 7288
rect 1524 7256 1564 7288
rect 1596 7256 1636 7288
rect 1668 7256 1708 7288
rect 1740 7256 1780 7288
rect 1812 7256 1852 7288
rect 1884 7256 1924 7288
rect 1956 7256 1996 7288
rect 2028 7256 2068 7288
rect 2100 7256 2140 7288
rect 2172 7256 2212 7288
rect 2244 7256 2284 7288
rect 2316 7256 2356 7288
rect 2388 7256 2428 7288
rect 2460 7256 2500 7288
rect 2532 7256 2572 7288
rect 2604 7256 2644 7288
rect 2676 7256 2716 7288
rect 2748 7256 2864 7288
rect 0 7165 2864 7256
rect 0 7133 116 7165
rect 148 7140 2708 7165
rect 148 7133 270 7140
rect 0 7093 270 7133
rect 0 7061 116 7093
rect 148 7061 270 7093
rect 0 7021 270 7061
rect 2600 7133 2708 7140
rect 2740 7133 2864 7165
rect 2600 7093 2864 7133
rect 2600 7061 2708 7093
rect 2740 7061 2864 7093
rect 0 6989 116 7021
rect 148 6989 270 7021
rect 0 6949 270 6989
rect 0 6917 116 6949
rect 148 6917 270 6949
rect 0 6877 270 6917
rect 0 6845 116 6877
rect 148 6845 270 6877
rect 0 6805 270 6845
rect 0 6773 116 6805
rect 148 6773 270 6805
rect 0 6733 270 6773
rect 0 6701 116 6733
rect 148 6701 270 6733
rect 0 6661 270 6701
rect 0 6629 116 6661
rect 148 6629 270 6661
rect 0 6589 270 6629
rect 0 6557 116 6589
rect 148 6557 270 6589
rect 0 6517 270 6557
rect 0 6485 116 6517
rect 148 6485 270 6517
rect 0 6445 270 6485
rect 0 6413 116 6445
rect 148 6413 270 6445
rect 0 6373 270 6413
rect 0 6341 116 6373
rect 148 6341 270 6373
rect 0 6301 270 6341
rect 0 6269 116 6301
rect 148 6269 270 6301
rect 0 6229 270 6269
rect 0 6197 116 6229
rect 148 6197 270 6229
rect 0 6157 270 6197
rect 0 6125 116 6157
rect 148 6125 270 6157
rect 0 6085 270 6125
rect 0 6053 116 6085
rect 148 6053 270 6085
rect 0 6013 270 6053
rect 0 5981 116 6013
rect 148 5981 270 6013
rect 0 5941 270 5981
rect 0 5909 116 5941
rect 148 5909 270 5941
rect 0 5869 270 5909
rect 0 5837 116 5869
rect 148 5837 270 5869
rect 0 5797 270 5837
rect 0 5765 116 5797
rect 148 5765 270 5797
rect 0 5725 270 5765
rect 0 5693 116 5725
rect 148 5693 270 5725
rect 0 5653 270 5693
rect 0 5621 116 5653
rect 148 5621 270 5653
rect 0 5581 270 5621
rect 0 5549 116 5581
rect 148 5549 270 5581
rect 0 5509 270 5549
rect 0 5477 116 5509
rect 148 5477 270 5509
rect 0 5437 270 5477
rect 0 5405 116 5437
rect 148 5405 270 5437
rect 0 5365 270 5405
rect 0 5333 116 5365
rect 148 5333 270 5365
rect 0 5293 270 5333
rect 0 5261 116 5293
rect 148 5261 270 5293
rect 0 5221 270 5261
rect 0 5189 116 5221
rect 148 5189 270 5221
rect 0 5149 270 5189
rect 0 5117 116 5149
rect 148 5117 270 5149
rect 0 5077 270 5117
rect 0 5045 116 5077
rect 148 5045 270 5077
rect 0 5005 270 5045
rect 0 4973 116 5005
rect 148 4973 270 5005
rect 0 4933 270 4973
rect 0 4901 116 4933
rect 148 4901 270 4933
rect 0 4861 270 4901
rect 0 4829 116 4861
rect 148 4829 270 4861
rect 0 4789 270 4829
rect 0 4757 116 4789
rect 148 4757 270 4789
rect 0 4717 270 4757
rect 0 4685 116 4717
rect 148 4685 270 4717
rect 0 4645 270 4685
rect 0 4613 116 4645
rect 148 4613 270 4645
rect 0 4573 270 4613
rect 0 4541 116 4573
rect 148 4541 270 4573
rect 0 4501 270 4541
rect 0 4469 116 4501
rect 148 4469 270 4501
rect 0 4429 270 4469
rect 0 4397 116 4429
rect 148 4397 270 4429
rect 0 4357 270 4397
rect 0 4325 116 4357
rect 148 4325 270 4357
rect 0 4285 270 4325
rect 0 4253 116 4285
rect 148 4253 270 4285
rect 0 4213 270 4253
rect 0 4181 116 4213
rect 148 4181 270 4213
rect 0 4141 270 4181
rect 0 4109 116 4141
rect 148 4109 270 4141
rect 0 4069 270 4109
rect 0 4037 116 4069
rect 148 4037 270 4069
rect 0 3997 270 4037
rect 0 3965 116 3997
rect 148 3965 270 3997
rect 0 3925 270 3965
rect 0 3893 116 3925
rect 148 3893 270 3925
rect 0 3853 270 3893
rect 0 3821 116 3853
rect 148 3821 270 3853
rect 0 3781 270 3821
rect 0 3749 116 3781
rect 148 3749 270 3781
rect 0 3709 270 3749
rect 0 3677 116 3709
rect 148 3677 270 3709
rect 0 3637 270 3677
rect 0 3605 116 3637
rect 148 3605 270 3637
rect 0 3565 270 3605
rect 0 3533 116 3565
rect 148 3533 270 3565
rect 0 3493 270 3533
rect 0 3461 116 3493
rect 148 3461 270 3493
rect 0 3421 270 3461
rect 0 3389 116 3421
rect 148 3389 270 3421
rect 0 3349 270 3389
rect 0 3317 116 3349
rect 148 3317 270 3349
rect 0 3277 270 3317
rect 0 3245 116 3277
rect 148 3245 270 3277
rect 0 3205 270 3245
rect 0 3173 116 3205
rect 148 3173 270 3205
rect 0 3133 270 3173
rect 0 3101 116 3133
rect 148 3101 270 3133
rect 0 3061 270 3101
rect 0 3029 116 3061
rect 148 3029 270 3061
rect 0 2989 270 3029
rect 0 2957 116 2989
rect 148 2957 270 2989
rect 0 2917 270 2957
rect 0 2885 116 2917
rect 148 2885 270 2917
rect 0 2845 270 2885
rect 0 2813 116 2845
rect 148 2813 270 2845
rect 0 2773 270 2813
rect 0 2741 116 2773
rect 148 2741 270 2773
rect 0 2701 270 2741
rect 0 2669 116 2701
rect 148 2669 270 2701
rect 0 2629 270 2669
rect 0 2597 116 2629
rect 148 2597 270 2629
rect 0 2557 270 2597
rect 0 2525 116 2557
rect 148 2525 270 2557
rect 0 2485 270 2525
rect 0 2453 116 2485
rect 148 2453 270 2485
rect 0 2413 270 2453
rect 0 2381 116 2413
rect 148 2381 270 2413
rect 0 2341 270 2381
rect 0 2309 116 2341
rect 148 2309 270 2341
rect 0 2269 270 2309
rect 0 2237 116 2269
rect 148 2237 270 2269
rect 0 2197 270 2237
rect 0 2165 116 2197
rect 148 2165 270 2197
rect 0 2125 270 2165
rect 0 2093 116 2125
rect 148 2093 270 2125
rect 0 2053 270 2093
rect 0 2021 116 2053
rect 148 2021 270 2053
rect 0 1981 270 2021
rect 0 1949 116 1981
rect 148 1949 270 1981
rect 0 1909 270 1949
rect 0 1877 116 1909
rect 148 1877 270 1909
rect 0 1837 270 1877
rect 0 1805 116 1837
rect 148 1805 270 1837
rect 0 1765 270 1805
rect 0 1733 116 1765
rect 148 1733 270 1765
rect 0 1693 270 1733
rect 0 1661 116 1693
rect 148 1661 270 1693
rect 0 1621 270 1661
rect 0 1589 116 1621
rect 148 1589 270 1621
rect 0 1549 270 1589
rect 0 1517 116 1549
rect 148 1517 270 1549
rect 0 1477 270 1517
rect 0 1445 116 1477
rect 148 1445 270 1477
rect 0 1405 270 1445
rect 0 1373 116 1405
rect 148 1373 270 1405
rect 0 1333 270 1373
rect 0 1301 116 1333
rect 148 1301 270 1333
rect 0 1261 270 1301
rect 0 1229 116 1261
rect 148 1229 270 1261
rect 0 1189 270 1229
rect 0 1157 116 1189
rect 148 1157 270 1189
rect 0 1117 270 1157
rect 0 1085 116 1117
rect 148 1085 270 1117
rect 0 1045 270 1085
rect 0 1013 116 1045
rect 148 1013 270 1045
rect 0 973 270 1013
rect 0 941 116 973
rect 148 941 270 973
rect 0 901 270 941
rect 0 869 116 901
rect 148 869 270 901
rect 0 829 270 869
rect 0 797 116 829
rect 148 797 270 829
rect 0 757 270 797
rect 0 725 116 757
rect 148 725 270 757
rect 0 685 270 725
rect 0 653 116 685
rect 148 653 270 685
rect 0 613 270 653
rect 0 581 116 613
rect 148 581 270 613
rect 0 541 270 581
rect 0 509 116 541
rect 148 509 270 541
rect 0 469 270 509
rect 0 437 116 469
rect 148 437 270 469
rect 0 397 270 437
rect 0 365 116 397
rect 148 365 270 397
rect 366 6980 2492 7032
rect 366 6948 447 6980
rect 479 6948 519 6980
rect 551 6948 591 6980
rect 623 6948 663 6980
rect 695 6948 735 6980
rect 767 6948 807 6980
rect 839 6948 879 6980
rect 911 6948 951 6980
rect 983 6948 1023 6980
rect 1055 6948 1095 6980
rect 1127 6948 1167 6980
rect 1199 6948 1239 6980
rect 1271 6948 1311 6980
rect 1343 6948 1383 6980
rect 1415 6948 1455 6980
rect 1487 6948 1527 6980
rect 1559 6948 1599 6980
rect 1631 6948 1671 6980
rect 1703 6948 1743 6980
rect 1775 6948 1815 6980
rect 1847 6948 1887 6980
rect 1919 6948 1959 6980
rect 1991 6948 2031 6980
rect 2063 6948 2103 6980
rect 2135 6948 2175 6980
rect 2207 6948 2247 6980
rect 2279 6948 2319 6980
rect 2351 6948 2391 6980
rect 2423 6948 2492 6980
rect 366 6908 2492 6948
rect 366 6876 447 6908
rect 479 6876 519 6908
rect 551 6876 591 6908
rect 623 6876 663 6908
rect 695 6876 735 6908
rect 767 6876 807 6908
rect 839 6876 879 6908
rect 911 6876 951 6908
rect 983 6876 1023 6908
rect 1055 6876 1095 6908
rect 1127 6876 1167 6908
rect 1199 6876 1239 6908
rect 1271 6876 1311 6908
rect 1343 6876 1383 6908
rect 1415 6876 1455 6908
rect 1487 6876 1527 6908
rect 1559 6876 1599 6908
rect 1631 6876 1671 6908
rect 1703 6876 1743 6908
rect 1775 6876 1815 6908
rect 1847 6876 1887 6908
rect 1919 6876 1959 6908
rect 1991 6876 2031 6908
rect 2063 6876 2103 6908
rect 2135 6876 2175 6908
rect 2207 6876 2247 6908
rect 2279 6876 2319 6908
rect 2351 6876 2391 6908
rect 2423 6876 2492 6908
rect 366 6836 2492 6876
rect 366 6804 447 6836
rect 479 6804 519 6836
rect 551 6804 591 6836
rect 623 6804 663 6836
rect 695 6804 735 6836
rect 767 6804 807 6836
rect 839 6804 879 6836
rect 911 6804 951 6836
rect 983 6804 1023 6836
rect 1055 6804 1095 6836
rect 1127 6804 1167 6836
rect 1199 6804 1239 6836
rect 1271 6804 1311 6836
rect 1343 6804 1383 6836
rect 1415 6804 1455 6836
rect 1487 6804 1527 6836
rect 1559 6804 1599 6836
rect 1631 6804 1671 6836
rect 1703 6804 1743 6836
rect 1775 6804 1815 6836
rect 1847 6804 1887 6836
rect 1919 6804 1959 6836
rect 1991 6804 2031 6836
rect 2063 6804 2103 6836
rect 2135 6804 2175 6836
rect 2207 6804 2247 6836
rect 2279 6804 2319 6836
rect 2351 6804 2391 6836
rect 2423 6804 2492 6836
rect 366 6761 2492 6804
rect 366 6729 433 6761
rect 465 6729 505 6761
rect 537 6729 577 6761
rect 609 6750 1345 6761
rect 609 6729 672 6750
rect 366 6689 672 6729
rect 366 6663 433 6689
rect 465 6663 505 6689
rect 366 6623 400 6663
rect 465 6657 496 6663
rect 537 6657 577 6689
rect 609 6663 672 6689
rect 440 6623 496 6657
rect 536 6623 592 6657
rect 632 6623 672 6663
rect 366 6617 672 6623
rect 366 6585 433 6617
rect 465 6585 505 6617
rect 537 6585 577 6617
rect 609 6585 672 6617
rect 366 6567 672 6585
rect 366 6527 400 6567
rect 440 6545 496 6567
rect 536 6545 592 6567
rect 465 6527 496 6545
rect 366 6513 433 6527
rect 465 6513 505 6527
rect 537 6513 577 6545
rect 632 6527 672 6567
rect 1272 6729 1345 6750
rect 1377 6729 1417 6761
rect 1449 6729 1489 6761
rect 1521 6750 2257 6761
rect 1521 6729 1584 6750
rect 1272 6689 1584 6729
rect 1272 6663 1345 6689
rect 1377 6663 1417 6689
rect 1272 6623 1312 6663
rect 1377 6657 1408 6663
rect 1449 6657 1489 6689
rect 1521 6663 1584 6689
rect 1352 6623 1408 6657
rect 1448 6623 1504 6657
rect 1544 6623 1584 6663
rect 1272 6617 1584 6623
rect 1272 6585 1345 6617
rect 1377 6585 1417 6617
rect 1449 6585 1489 6617
rect 1521 6585 1584 6617
rect 1272 6567 1584 6585
rect 609 6513 672 6527
rect 366 6473 672 6513
rect 366 6471 433 6473
rect 465 6471 505 6473
rect 366 6431 400 6471
rect 465 6441 496 6471
rect 537 6441 577 6473
rect 609 6471 672 6473
rect 440 6431 496 6441
rect 536 6431 592 6441
rect 632 6431 672 6471
rect 366 6401 672 6431
rect 366 6375 433 6401
rect 465 6375 505 6401
rect 366 6335 400 6375
rect 465 6369 496 6375
rect 537 6369 577 6401
rect 609 6375 672 6401
rect 440 6335 496 6369
rect 536 6335 592 6369
rect 632 6335 672 6375
rect 366 6329 672 6335
rect 366 6297 433 6329
rect 465 6297 505 6329
rect 537 6297 577 6329
rect 609 6297 672 6329
rect 366 6279 672 6297
rect 366 6239 400 6279
rect 440 6257 496 6279
rect 536 6257 592 6279
rect 465 6239 496 6257
rect 366 6225 433 6239
rect 465 6225 505 6239
rect 537 6225 577 6257
rect 632 6239 672 6279
rect 609 6225 672 6239
rect 366 6185 672 6225
rect 366 6183 433 6185
rect 465 6183 505 6185
rect 366 6143 400 6183
rect 465 6153 496 6183
rect 537 6153 577 6185
rect 609 6183 672 6185
rect 440 6143 496 6153
rect 536 6143 592 6153
rect 632 6143 672 6183
rect 366 6113 672 6143
rect 366 6081 433 6113
rect 465 6081 505 6113
rect 537 6081 577 6113
rect 609 6081 672 6113
rect 366 6041 672 6081
rect 366 6009 433 6041
rect 465 6009 505 6041
rect 537 6009 577 6041
rect 609 6009 672 6041
rect 366 5969 672 6009
rect 366 5937 433 5969
rect 465 5937 505 5969
rect 537 5937 577 5969
rect 609 5937 672 5969
rect 366 5897 672 5937
rect 366 5865 433 5897
rect 465 5865 505 5897
rect 537 5865 577 5897
rect 609 5865 672 5897
rect 366 5825 672 5865
rect 366 5793 433 5825
rect 465 5793 505 5825
rect 537 5793 577 5825
rect 609 5793 672 5825
rect 366 5753 672 5793
rect 366 5721 433 5753
rect 465 5721 505 5753
rect 537 5721 577 5753
rect 609 5721 672 5753
rect 366 5681 672 5721
rect 366 5649 433 5681
rect 465 5649 505 5681
rect 537 5649 577 5681
rect 609 5649 672 5681
rect 366 5609 672 5649
rect 366 5577 433 5609
rect 465 5577 505 5609
rect 537 5577 577 5609
rect 609 5577 672 5609
rect 366 5537 672 5577
rect 366 5505 433 5537
rect 465 5505 505 5537
rect 537 5505 577 5537
rect 609 5505 672 5537
rect 366 5465 672 5505
rect 366 5433 433 5465
rect 465 5433 505 5465
rect 537 5433 577 5465
rect 609 5433 672 5465
rect 366 5393 672 5433
rect 366 5361 433 5393
rect 465 5361 505 5393
rect 537 5361 577 5393
rect 609 5361 672 5393
rect 366 5321 672 5361
rect 366 5289 433 5321
rect 465 5289 505 5321
rect 537 5289 577 5321
rect 609 5289 672 5321
rect 366 5249 672 5289
rect 366 5217 433 5249
rect 465 5217 505 5249
rect 537 5217 577 5249
rect 609 5217 672 5249
rect 366 5177 672 5217
rect 366 5145 433 5177
rect 465 5145 505 5177
rect 537 5145 577 5177
rect 609 5145 672 5177
rect 366 5105 672 5145
rect 366 5073 433 5105
rect 465 5073 505 5105
rect 537 5073 577 5105
rect 609 5073 672 5105
rect 366 5033 672 5073
rect 366 5001 433 5033
rect 465 5001 505 5033
rect 537 5001 577 5033
rect 609 5001 672 5033
rect 366 4961 672 5001
rect 366 4929 433 4961
rect 465 4929 505 4961
rect 537 4929 577 4961
rect 609 4929 672 4961
rect 366 4889 672 4929
rect 366 4863 433 4889
rect 465 4863 505 4889
rect 366 4823 400 4863
rect 465 4857 496 4863
rect 537 4857 577 4889
rect 609 4863 672 4889
rect 440 4823 496 4857
rect 536 4823 592 4857
rect 632 4823 672 4863
rect 366 4817 672 4823
rect 366 4785 433 4817
rect 465 4785 505 4817
rect 537 4785 577 4817
rect 609 4785 672 4817
rect 366 4767 672 4785
rect 366 4727 400 4767
rect 440 4745 496 4767
rect 536 4745 592 4767
rect 465 4727 496 4745
rect 366 4713 433 4727
rect 465 4713 505 4727
rect 537 4713 577 4745
rect 632 4727 672 4767
rect 609 4713 672 4727
rect 366 4673 672 4713
rect 366 4671 433 4673
rect 465 4671 505 4673
rect 366 4631 400 4671
rect 465 4641 496 4671
rect 537 4641 577 4673
rect 609 4671 672 4673
rect 440 4631 496 4641
rect 536 4631 592 4641
rect 632 4631 672 4671
rect 366 4601 672 4631
rect 366 4575 433 4601
rect 465 4575 505 4601
rect 366 4535 400 4575
rect 465 4569 496 4575
rect 537 4569 577 4601
rect 609 4575 672 4601
rect 440 4535 496 4569
rect 536 4535 592 4569
rect 632 4535 672 4575
rect 366 4529 672 4535
rect 366 4497 433 4529
rect 465 4497 505 4529
rect 537 4497 577 4529
rect 609 4497 672 4529
rect 366 4479 672 4497
rect 366 4439 400 4479
rect 440 4457 496 4479
rect 536 4457 592 4479
rect 465 4439 496 4457
rect 366 4425 433 4439
rect 465 4425 505 4439
rect 537 4425 577 4457
rect 632 4439 672 4479
rect 609 4425 672 4439
rect 366 4385 672 4425
rect 366 4383 433 4385
rect 465 4383 505 4385
rect 366 4343 400 4383
rect 465 4353 496 4383
rect 537 4353 577 4385
rect 609 4383 672 4385
rect 440 4343 496 4353
rect 536 4343 592 4353
rect 632 4343 672 4383
rect 366 4313 672 4343
rect 366 4281 433 4313
rect 465 4281 505 4313
rect 537 4281 577 4313
rect 609 4281 672 4313
rect 366 4241 672 4281
rect 366 4209 433 4241
rect 465 4209 505 4241
rect 537 4209 577 4241
rect 609 4209 672 4241
rect 366 4169 672 4209
rect 366 4137 433 4169
rect 465 4137 505 4169
rect 537 4137 577 4169
rect 609 4137 672 4169
rect 366 4097 672 4137
rect 366 4065 433 4097
rect 465 4065 505 4097
rect 537 4065 577 4097
rect 609 4065 672 4097
rect 366 4025 672 4065
rect 366 3993 433 4025
rect 465 3993 505 4025
rect 537 3993 577 4025
rect 609 3993 672 4025
rect 366 3953 672 3993
rect 366 3921 433 3953
rect 465 3921 505 3953
rect 537 3921 577 3953
rect 609 3921 672 3953
rect 366 3881 672 3921
rect 366 3849 433 3881
rect 465 3849 505 3881
rect 537 3849 577 3881
rect 609 3849 672 3881
rect 366 3809 672 3849
rect 366 3777 433 3809
rect 465 3777 505 3809
rect 537 3777 577 3809
rect 609 3777 672 3809
rect 366 3737 672 3777
rect 366 3705 433 3737
rect 465 3705 505 3737
rect 537 3705 577 3737
rect 609 3705 672 3737
rect 366 3665 672 3705
rect 366 3633 433 3665
rect 465 3633 505 3665
rect 537 3633 577 3665
rect 609 3633 672 3665
rect 366 3593 672 3633
rect 366 3561 433 3593
rect 465 3561 505 3593
rect 537 3561 577 3593
rect 609 3561 672 3593
rect 366 3521 672 3561
rect 366 3489 433 3521
rect 465 3489 505 3521
rect 537 3489 577 3521
rect 609 3489 672 3521
rect 366 3449 672 3489
rect 366 3417 433 3449
rect 465 3417 505 3449
rect 537 3417 577 3449
rect 609 3417 672 3449
rect 366 3377 672 3417
rect 366 3345 433 3377
rect 465 3345 505 3377
rect 537 3345 577 3377
rect 609 3345 672 3377
rect 366 3305 672 3345
rect 366 3273 433 3305
rect 465 3273 505 3305
rect 537 3273 577 3305
rect 609 3273 672 3305
rect 366 3233 672 3273
rect 366 3201 433 3233
rect 465 3201 505 3233
rect 537 3201 577 3233
rect 609 3201 672 3233
rect 366 3161 672 3201
rect 366 3129 433 3161
rect 465 3129 505 3161
rect 537 3129 577 3161
rect 609 3129 672 3161
rect 366 3089 672 3129
rect 366 3063 433 3089
rect 465 3063 505 3089
rect 366 3023 400 3063
rect 465 3057 496 3063
rect 537 3057 577 3089
rect 609 3063 672 3089
rect 440 3023 496 3057
rect 536 3023 592 3057
rect 632 3023 672 3063
rect 366 3017 672 3023
rect 366 2985 433 3017
rect 465 2985 505 3017
rect 537 2985 577 3017
rect 609 2985 672 3017
rect 366 2967 672 2985
rect 366 2927 400 2967
rect 440 2945 496 2967
rect 536 2945 592 2967
rect 465 2927 496 2945
rect 366 2913 433 2927
rect 465 2913 505 2927
rect 537 2913 577 2945
rect 632 2927 672 2967
rect 609 2913 672 2927
rect 366 2873 672 2913
rect 366 2871 433 2873
rect 465 2871 505 2873
rect 366 2831 400 2871
rect 465 2841 496 2871
rect 537 2841 577 2873
rect 609 2871 672 2873
rect 440 2831 496 2841
rect 536 2831 592 2841
rect 632 2831 672 2871
rect 366 2801 672 2831
rect 366 2775 433 2801
rect 465 2775 505 2801
rect 366 2735 400 2775
rect 465 2769 496 2775
rect 537 2769 577 2801
rect 609 2775 672 2801
rect 440 2735 496 2769
rect 536 2735 592 2769
rect 632 2735 672 2775
rect 366 2729 672 2735
rect 366 2697 433 2729
rect 465 2697 505 2729
rect 537 2697 577 2729
rect 609 2697 672 2729
rect 366 2679 672 2697
rect 366 2639 400 2679
rect 440 2657 496 2679
rect 536 2657 592 2679
rect 465 2639 496 2657
rect 366 2625 433 2639
rect 465 2625 505 2639
rect 537 2625 577 2657
rect 632 2639 672 2679
rect 609 2625 672 2639
rect 366 2585 672 2625
rect 366 2583 433 2585
rect 465 2583 505 2585
rect 366 2543 400 2583
rect 465 2553 496 2583
rect 537 2553 577 2585
rect 609 2583 672 2585
rect 440 2543 496 2553
rect 536 2543 592 2553
rect 632 2543 672 2583
rect 366 2513 672 2543
rect 366 2481 433 2513
rect 465 2481 505 2513
rect 537 2481 577 2513
rect 609 2481 672 2513
rect 366 2441 672 2481
rect 366 2409 433 2441
rect 465 2409 505 2441
rect 537 2409 577 2441
rect 609 2409 672 2441
rect 366 2369 672 2409
rect 366 2337 433 2369
rect 465 2337 505 2369
rect 537 2337 577 2369
rect 609 2337 672 2369
rect 366 2297 672 2337
rect 366 2265 433 2297
rect 465 2265 505 2297
rect 537 2265 577 2297
rect 609 2265 672 2297
rect 366 2225 672 2265
rect 366 2193 433 2225
rect 465 2193 505 2225
rect 537 2193 577 2225
rect 609 2193 672 2225
rect 366 2153 672 2193
rect 366 2121 433 2153
rect 465 2121 505 2153
rect 537 2121 577 2153
rect 609 2121 672 2153
rect 366 2081 672 2121
rect 366 2049 433 2081
rect 465 2049 505 2081
rect 537 2049 577 2081
rect 609 2049 672 2081
rect 366 2009 672 2049
rect 366 1977 433 2009
rect 465 1977 505 2009
rect 537 1977 577 2009
rect 609 1977 672 2009
rect 366 1937 672 1977
rect 366 1905 433 1937
rect 465 1905 505 1937
rect 537 1905 577 1937
rect 609 1905 672 1937
rect 366 1865 672 1905
rect 366 1833 433 1865
rect 465 1833 505 1865
rect 537 1833 577 1865
rect 609 1833 672 1865
rect 366 1793 672 1833
rect 366 1761 433 1793
rect 465 1761 505 1793
rect 537 1761 577 1793
rect 609 1761 672 1793
rect 366 1721 672 1761
rect 366 1689 433 1721
rect 465 1689 505 1721
rect 537 1689 577 1721
rect 609 1689 672 1721
rect 366 1649 672 1689
rect 366 1617 433 1649
rect 465 1617 505 1649
rect 537 1617 577 1649
rect 609 1617 672 1649
rect 366 1577 672 1617
rect 366 1545 433 1577
rect 465 1545 505 1577
rect 537 1545 577 1577
rect 609 1545 672 1577
rect 366 1505 672 1545
rect 366 1473 433 1505
rect 465 1473 505 1505
rect 537 1473 577 1505
rect 609 1473 672 1505
rect 366 1433 672 1473
rect 366 1401 433 1433
rect 465 1401 505 1433
rect 537 1401 577 1433
rect 609 1401 672 1433
rect 366 1361 672 1401
rect 366 1329 433 1361
rect 465 1329 505 1361
rect 537 1329 577 1361
rect 609 1329 672 1361
rect 366 1289 672 1329
rect 366 1263 433 1289
rect 465 1263 505 1289
rect 366 1223 400 1263
rect 465 1257 496 1263
rect 537 1257 577 1289
rect 609 1263 672 1289
rect 440 1223 496 1257
rect 536 1223 592 1257
rect 632 1223 672 1263
rect 366 1217 672 1223
rect 366 1185 433 1217
rect 465 1185 505 1217
rect 537 1185 577 1217
rect 609 1185 672 1217
rect 366 1167 672 1185
rect 366 1127 400 1167
rect 440 1145 496 1167
rect 536 1145 592 1167
rect 465 1127 496 1145
rect 366 1113 433 1127
rect 465 1113 505 1127
rect 537 1113 577 1145
rect 632 1127 672 1167
rect 609 1113 672 1127
rect 366 1073 672 1113
rect 366 1071 433 1073
rect 465 1071 505 1073
rect 366 1031 400 1071
rect 465 1041 496 1071
rect 537 1041 577 1073
rect 609 1071 672 1073
rect 440 1031 496 1041
rect 536 1031 592 1041
rect 632 1031 672 1071
rect 366 1001 672 1031
rect 366 975 433 1001
rect 465 975 505 1001
rect 366 935 400 975
rect 465 969 496 975
rect 537 969 577 1001
rect 609 975 672 1001
rect 440 935 496 969
rect 536 935 592 969
rect 632 935 672 975
rect 366 929 672 935
rect 366 897 433 929
rect 465 897 505 929
rect 537 897 577 929
rect 609 897 672 929
rect 366 879 672 897
rect 366 839 400 879
rect 440 857 496 879
rect 536 857 592 879
rect 465 839 496 857
rect 366 825 433 839
rect 465 825 505 839
rect 537 825 577 857
rect 632 839 672 879
rect 792 6466 1152 6540
rect 792 6434 888 6466
rect 920 6434 960 6466
rect 992 6434 1032 6466
rect 1064 6434 1152 6466
rect 792 6394 1152 6434
rect 792 6362 888 6394
rect 920 6362 960 6394
rect 992 6362 1032 6394
rect 1064 6362 1152 6394
rect 792 6322 1152 6362
rect 792 6290 888 6322
rect 920 6290 960 6322
rect 992 6290 1032 6322
rect 1064 6290 1152 6322
rect 792 6250 1152 6290
rect 792 6218 888 6250
rect 920 6218 960 6250
rect 992 6218 1032 6250
rect 1064 6218 1152 6250
rect 792 6178 1152 6218
rect 792 6146 888 6178
rect 920 6146 960 6178
rect 992 6146 1032 6178
rect 1064 6146 1152 6178
rect 792 6106 1152 6146
rect 792 6074 888 6106
rect 920 6074 960 6106
rect 992 6074 1032 6106
rect 1064 6074 1152 6106
rect 792 6034 1152 6074
rect 792 6002 888 6034
rect 920 6002 960 6034
rect 992 6002 1032 6034
rect 1064 6002 1152 6034
rect 792 5962 1152 6002
rect 792 5930 888 5962
rect 920 5930 960 5962
rect 992 5930 1032 5962
rect 1064 5930 1152 5962
rect 792 5890 1152 5930
rect 792 5858 888 5890
rect 920 5858 960 5890
rect 992 5858 1032 5890
rect 1064 5858 1152 5890
rect 792 5847 1152 5858
rect 792 5807 860 5847
rect 900 5818 956 5847
rect 996 5818 1052 5847
rect 920 5807 956 5818
rect 996 5807 1032 5818
rect 1092 5807 1152 5847
rect 792 5786 888 5807
rect 920 5786 960 5807
rect 992 5786 1032 5807
rect 1064 5786 1152 5807
rect 792 5751 1152 5786
rect 792 5711 860 5751
rect 900 5746 956 5751
rect 996 5746 1052 5751
rect 920 5714 956 5746
rect 996 5714 1032 5746
rect 900 5711 956 5714
rect 996 5711 1052 5714
rect 1092 5711 1152 5751
rect 792 5674 1152 5711
rect 792 5655 888 5674
rect 920 5655 960 5674
rect 992 5655 1032 5674
rect 1064 5655 1152 5674
rect 792 5615 860 5655
rect 920 5642 956 5655
rect 996 5642 1032 5655
rect 900 5615 956 5642
rect 996 5615 1052 5642
rect 1092 5615 1152 5655
rect 792 5602 1152 5615
rect 792 5570 888 5602
rect 920 5570 960 5602
rect 992 5570 1032 5602
rect 1064 5570 1152 5602
rect 792 5559 1152 5570
rect 792 5519 860 5559
rect 900 5530 956 5559
rect 996 5530 1052 5559
rect 920 5519 956 5530
rect 996 5519 1032 5530
rect 1092 5519 1152 5559
rect 792 5498 888 5519
rect 920 5498 960 5519
rect 992 5498 1032 5519
rect 1064 5498 1152 5519
rect 792 5463 1152 5498
rect 792 5423 860 5463
rect 900 5458 956 5463
rect 996 5458 1052 5463
rect 920 5426 956 5458
rect 996 5426 1032 5458
rect 900 5423 956 5426
rect 996 5423 1052 5426
rect 1092 5423 1152 5463
rect 792 5386 1152 5423
rect 792 5367 888 5386
rect 920 5367 960 5386
rect 992 5367 1032 5386
rect 1064 5367 1152 5386
rect 792 5327 860 5367
rect 920 5354 956 5367
rect 996 5354 1032 5367
rect 900 5327 956 5354
rect 996 5327 1052 5354
rect 1092 5327 1152 5367
rect 792 5314 1152 5327
rect 792 5282 888 5314
rect 920 5282 960 5314
rect 992 5282 1032 5314
rect 1064 5282 1152 5314
rect 792 5271 1152 5282
rect 792 5231 860 5271
rect 900 5242 956 5271
rect 996 5242 1052 5271
rect 920 5231 956 5242
rect 996 5231 1032 5242
rect 1092 5231 1152 5271
rect 792 5210 888 5231
rect 920 5210 960 5231
rect 992 5210 1032 5231
rect 1064 5210 1152 5231
rect 792 5175 1152 5210
rect 792 5135 860 5175
rect 900 5170 956 5175
rect 996 5170 1052 5175
rect 920 5138 956 5170
rect 996 5138 1032 5170
rect 900 5135 956 5138
rect 996 5135 1052 5138
rect 1092 5135 1152 5175
rect 792 5098 1152 5135
rect 792 5066 888 5098
rect 920 5066 960 5098
rect 992 5066 1032 5098
rect 1064 5066 1152 5098
rect 792 5026 1152 5066
rect 792 4994 888 5026
rect 920 4994 960 5026
rect 992 4994 1032 5026
rect 1064 4994 1152 5026
rect 792 4954 1152 4994
rect 792 4922 888 4954
rect 920 4922 960 4954
rect 992 4922 1032 4954
rect 1064 4922 1152 4954
rect 792 4882 1152 4922
rect 792 4850 888 4882
rect 920 4850 960 4882
rect 992 4850 1032 4882
rect 1064 4850 1152 4882
rect 792 4810 1152 4850
rect 792 4778 888 4810
rect 920 4778 960 4810
rect 992 4778 1032 4810
rect 1064 4778 1152 4810
rect 792 4738 1152 4778
rect 792 4706 888 4738
rect 920 4706 960 4738
rect 992 4706 1032 4738
rect 1064 4706 1152 4738
rect 792 4666 1152 4706
rect 792 4634 888 4666
rect 920 4634 960 4666
rect 992 4634 1032 4666
rect 1064 4634 1152 4666
rect 792 4594 1152 4634
rect 792 4562 888 4594
rect 920 4562 960 4594
rect 992 4562 1032 4594
rect 1064 4562 1152 4594
rect 792 4522 1152 4562
rect 792 4490 888 4522
rect 920 4490 960 4522
rect 992 4490 1032 4522
rect 1064 4490 1152 4522
rect 792 4450 1152 4490
rect 792 4418 888 4450
rect 920 4418 960 4450
rect 992 4418 1032 4450
rect 1064 4418 1152 4450
rect 792 4378 1152 4418
rect 792 4346 888 4378
rect 920 4346 960 4378
rect 992 4346 1032 4378
rect 1064 4346 1152 4378
rect 792 4306 1152 4346
rect 792 4274 888 4306
rect 920 4274 960 4306
rect 992 4274 1032 4306
rect 1064 4274 1152 4306
rect 792 4234 1152 4274
rect 792 4202 888 4234
rect 920 4202 960 4234
rect 992 4202 1032 4234
rect 1064 4202 1152 4234
rect 792 4162 1152 4202
rect 792 4130 888 4162
rect 920 4130 960 4162
rect 992 4130 1032 4162
rect 1064 4130 1152 4162
rect 792 4090 1152 4130
rect 792 4058 888 4090
rect 920 4058 960 4090
rect 992 4058 1032 4090
rect 1064 4058 1152 4090
rect 792 4047 1152 4058
rect 792 4007 860 4047
rect 900 4018 956 4047
rect 996 4018 1052 4047
rect 920 4007 956 4018
rect 996 4007 1032 4018
rect 1092 4007 1152 4047
rect 792 3986 888 4007
rect 920 3986 960 4007
rect 992 3986 1032 4007
rect 1064 3986 1152 4007
rect 792 3951 1152 3986
rect 792 3911 860 3951
rect 900 3946 956 3951
rect 996 3946 1052 3951
rect 920 3914 956 3946
rect 996 3914 1032 3946
rect 900 3911 956 3914
rect 996 3911 1052 3914
rect 1092 3911 1152 3951
rect 792 3874 1152 3911
rect 792 3855 888 3874
rect 920 3855 960 3874
rect 992 3855 1032 3874
rect 1064 3855 1152 3874
rect 792 3815 860 3855
rect 920 3842 956 3855
rect 996 3842 1032 3855
rect 900 3815 956 3842
rect 996 3815 1052 3842
rect 1092 3815 1152 3855
rect 792 3802 1152 3815
rect 792 3770 888 3802
rect 920 3770 960 3802
rect 992 3770 1032 3802
rect 1064 3770 1152 3802
rect 792 3759 1152 3770
rect 792 3719 860 3759
rect 900 3730 956 3759
rect 996 3730 1052 3759
rect 920 3719 956 3730
rect 996 3719 1032 3730
rect 1092 3719 1152 3759
rect 792 3698 888 3719
rect 920 3698 960 3719
rect 992 3698 1032 3719
rect 1064 3698 1152 3719
rect 792 3663 1152 3698
rect 792 3623 860 3663
rect 900 3658 956 3663
rect 996 3658 1052 3663
rect 920 3626 956 3658
rect 996 3626 1032 3658
rect 900 3623 956 3626
rect 996 3623 1052 3626
rect 1092 3623 1152 3663
rect 792 3586 1152 3623
rect 792 3567 888 3586
rect 920 3567 960 3586
rect 992 3567 1032 3586
rect 1064 3567 1152 3586
rect 792 3527 860 3567
rect 920 3554 956 3567
rect 996 3554 1032 3567
rect 900 3527 956 3554
rect 996 3527 1052 3554
rect 1092 3527 1152 3567
rect 792 3514 1152 3527
rect 792 3482 888 3514
rect 920 3482 960 3514
rect 992 3482 1032 3514
rect 1064 3482 1152 3514
rect 792 3471 1152 3482
rect 792 3431 860 3471
rect 900 3442 956 3471
rect 996 3442 1052 3471
rect 920 3431 956 3442
rect 996 3431 1032 3442
rect 1092 3431 1152 3471
rect 792 3410 888 3431
rect 920 3410 960 3431
rect 992 3410 1032 3431
rect 1064 3410 1152 3431
rect 792 3375 1152 3410
rect 792 3335 860 3375
rect 900 3370 956 3375
rect 996 3370 1052 3375
rect 920 3338 956 3370
rect 996 3338 1032 3370
rect 900 3335 956 3338
rect 996 3335 1052 3338
rect 1092 3335 1152 3375
rect 792 3298 1152 3335
rect 792 3266 888 3298
rect 920 3266 960 3298
rect 992 3266 1032 3298
rect 1064 3266 1152 3298
rect 792 3226 1152 3266
rect 792 3194 888 3226
rect 920 3194 960 3226
rect 992 3194 1032 3226
rect 1064 3194 1152 3226
rect 792 3154 1152 3194
rect 792 3122 888 3154
rect 920 3122 960 3154
rect 992 3122 1032 3154
rect 1064 3122 1152 3154
rect 792 3082 1152 3122
rect 792 3050 888 3082
rect 920 3050 960 3082
rect 992 3050 1032 3082
rect 1064 3050 1152 3082
rect 792 3010 1152 3050
rect 792 2978 888 3010
rect 920 2978 960 3010
rect 992 2978 1032 3010
rect 1064 2978 1152 3010
rect 792 2938 1152 2978
rect 792 2906 888 2938
rect 920 2906 960 2938
rect 992 2906 1032 2938
rect 1064 2906 1152 2938
rect 792 2866 1152 2906
rect 792 2834 888 2866
rect 920 2834 960 2866
rect 992 2834 1032 2866
rect 1064 2834 1152 2866
rect 792 2794 1152 2834
rect 792 2762 888 2794
rect 920 2762 960 2794
rect 992 2762 1032 2794
rect 1064 2762 1152 2794
rect 792 2722 1152 2762
rect 792 2690 888 2722
rect 920 2690 960 2722
rect 992 2690 1032 2722
rect 1064 2690 1152 2722
rect 792 2650 1152 2690
rect 792 2618 888 2650
rect 920 2618 960 2650
rect 992 2618 1032 2650
rect 1064 2618 1152 2650
rect 792 2578 1152 2618
rect 792 2546 888 2578
rect 920 2546 960 2578
rect 992 2546 1032 2578
rect 1064 2546 1152 2578
rect 792 2506 1152 2546
rect 792 2474 888 2506
rect 920 2474 960 2506
rect 992 2474 1032 2506
rect 1064 2474 1152 2506
rect 792 2434 1152 2474
rect 792 2402 888 2434
rect 920 2402 960 2434
rect 992 2402 1032 2434
rect 1064 2402 1152 2434
rect 792 2362 1152 2402
rect 792 2330 888 2362
rect 920 2330 960 2362
rect 992 2330 1032 2362
rect 1064 2330 1152 2362
rect 792 2290 1152 2330
rect 792 2258 888 2290
rect 920 2258 960 2290
rect 992 2258 1032 2290
rect 1064 2258 1152 2290
rect 792 2247 1152 2258
rect 792 2207 860 2247
rect 900 2218 956 2247
rect 996 2218 1052 2247
rect 920 2207 956 2218
rect 996 2207 1032 2218
rect 1092 2207 1152 2247
rect 792 2186 888 2207
rect 920 2186 960 2207
rect 992 2186 1032 2207
rect 1064 2186 1152 2207
rect 792 2151 1152 2186
rect 792 2111 860 2151
rect 900 2146 956 2151
rect 996 2146 1052 2151
rect 920 2114 956 2146
rect 996 2114 1032 2146
rect 900 2111 956 2114
rect 996 2111 1052 2114
rect 1092 2111 1152 2151
rect 792 2074 1152 2111
rect 792 2055 888 2074
rect 920 2055 960 2074
rect 992 2055 1032 2074
rect 1064 2055 1152 2074
rect 792 2015 860 2055
rect 920 2042 956 2055
rect 996 2042 1032 2055
rect 900 2015 956 2042
rect 996 2015 1052 2042
rect 1092 2015 1152 2055
rect 792 2002 1152 2015
rect 792 1970 888 2002
rect 920 1970 960 2002
rect 992 1970 1032 2002
rect 1064 1970 1152 2002
rect 792 1959 1152 1970
rect 792 1919 860 1959
rect 900 1930 956 1959
rect 996 1930 1052 1959
rect 920 1919 956 1930
rect 996 1919 1032 1930
rect 1092 1919 1152 1959
rect 792 1898 888 1919
rect 920 1898 960 1919
rect 992 1898 1032 1919
rect 1064 1898 1152 1919
rect 792 1863 1152 1898
rect 792 1823 860 1863
rect 900 1858 956 1863
rect 996 1858 1052 1863
rect 920 1826 956 1858
rect 996 1826 1032 1858
rect 900 1823 956 1826
rect 996 1823 1052 1826
rect 1092 1823 1152 1863
rect 792 1786 1152 1823
rect 792 1767 888 1786
rect 920 1767 960 1786
rect 992 1767 1032 1786
rect 1064 1767 1152 1786
rect 792 1727 860 1767
rect 920 1754 956 1767
rect 996 1754 1032 1767
rect 900 1727 956 1754
rect 996 1727 1052 1754
rect 1092 1727 1152 1767
rect 792 1714 1152 1727
rect 792 1682 888 1714
rect 920 1682 960 1714
rect 992 1682 1032 1714
rect 1064 1682 1152 1714
rect 792 1671 1152 1682
rect 792 1631 860 1671
rect 900 1642 956 1671
rect 996 1642 1052 1671
rect 920 1631 956 1642
rect 996 1631 1032 1642
rect 1092 1631 1152 1671
rect 792 1610 888 1631
rect 920 1610 960 1631
rect 992 1610 1032 1631
rect 1064 1610 1152 1631
rect 792 1575 1152 1610
rect 792 1535 860 1575
rect 900 1570 956 1575
rect 996 1570 1052 1575
rect 920 1538 956 1570
rect 996 1538 1032 1570
rect 900 1535 956 1538
rect 996 1535 1052 1538
rect 1092 1535 1152 1575
rect 792 1498 1152 1535
rect 792 1466 888 1498
rect 920 1466 960 1498
rect 992 1466 1032 1498
rect 1064 1466 1152 1498
rect 792 1426 1152 1466
rect 792 1394 888 1426
rect 920 1394 960 1426
rect 992 1394 1032 1426
rect 1064 1394 1152 1426
rect 792 1354 1152 1394
rect 792 1322 888 1354
rect 920 1322 960 1354
rect 992 1322 1032 1354
rect 1064 1322 1152 1354
rect 792 1282 1152 1322
rect 792 1250 888 1282
rect 920 1250 960 1282
rect 992 1250 1032 1282
rect 1064 1250 1152 1282
rect 792 1210 1152 1250
rect 792 1178 888 1210
rect 920 1178 960 1210
rect 992 1178 1032 1210
rect 1064 1178 1152 1210
rect 792 1138 1152 1178
rect 792 1106 888 1138
rect 920 1106 960 1138
rect 992 1106 1032 1138
rect 1064 1106 1152 1138
rect 792 1066 1152 1106
rect 792 1034 888 1066
rect 920 1034 960 1066
rect 992 1034 1032 1066
rect 1064 1034 1152 1066
rect 792 994 1152 1034
rect 792 962 888 994
rect 920 962 960 994
rect 992 962 1032 994
rect 1064 962 1152 994
rect 792 870 1152 962
rect 1272 6527 1312 6567
rect 1352 6545 1408 6567
rect 1448 6545 1504 6567
rect 1377 6527 1408 6545
rect 1272 6513 1345 6527
rect 1377 6513 1417 6527
rect 1449 6513 1489 6545
rect 1544 6527 1584 6567
rect 2180 6729 2257 6750
rect 2289 6729 2329 6761
rect 2361 6729 2401 6761
rect 2433 6729 2492 6761
rect 2180 6689 2492 6729
rect 2180 6663 2257 6689
rect 2289 6663 2329 6689
rect 2180 6623 2224 6663
rect 2289 6657 2320 6663
rect 2361 6657 2401 6689
rect 2433 6663 2492 6689
rect 2264 6623 2320 6657
rect 2360 6623 2416 6657
rect 2456 6623 2492 6663
rect 2180 6617 2492 6623
rect 2180 6585 2257 6617
rect 2289 6585 2329 6617
rect 2361 6585 2401 6617
rect 2433 6585 2492 6617
rect 2180 6567 2492 6585
rect 1521 6513 1584 6527
rect 1272 6473 1584 6513
rect 1272 6471 1345 6473
rect 1377 6471 1417 6473
rect 1272 6431 1312 6471
rect 1377 6441 1408 6471
rect 1449 6441 1489 6473
rect 1521 6471 1584 6473
rect 1352 6431 1408 6441
rect 1448 6431 1504 6441
rect 1544 6431 1584 6471
rect 1272 6401 1584 6431
rect 1272 6375 1345 6401
rect 1377 6375 1417 6401
rect 1272 6335 1312 6375
rect 1377 6369 1408 6375
rect 1449 6369 1489 6401
rect 1521 6375 1584 6401
rect 1352 6335 1408 6369
rect 1448 6335 1504 6369
rect 1544 6335 1584 6375
rect 1272 6329 1584 6335
rect 1272 6297 1345 6329
rect 1377 6297 1417 6329
rect 1449 6297 1489 6329
rect 1521 6297 1584 6329
rect 1272 6279 1584 6297
rect 1272 6239 1312 6279
rect 1352 6257 1408 6279
rect 1448 6257 1504 6279
rect 1377 6239 1408 6257
rect 1272 6225 1345 6239
rect 1377 6225 1417 6239
rect 1449 6225 1489 6257
rect 1544 6239 1584 6279
rect 1521 6225 1584 6239
rect 1272 6185 1584 6225
rect 1272 6183 1345 6185
rect 1377 6183 1417 6185
rect 1272 6143 1312 6183
rect 1377 6153 1408 6183
rect 1449 6153 1489 6185
rect 1521 6183 1584 6185
rect 1352 6143 1408 6153
rect 1448 6143 1504 6153
rect 1544 6143 1584 6183
rect 1272 6113 1584 6143
rect 1272 6081 1345 6113
rect 1377 6081 1417 6113
rect 1449 6081 1489 6113
rect 1521 6081 1584 6113
rect 1272 6041 1584 6081
rect 1272 6009 1345 6041
rect 1377 6009 1417 6041
rect 1449 6009 1489 6041
rect 1521 6009 1584 6041
rect 1272 5969 1584 6009
rect 1272 5937 1345 5969
rect 1377 5937 1417 5969
rect 1449 5937 1489 5969
rect 1521 5937 1584 5969
rect 1272 5897 1584 5937
rect 1272 5865 1345 5897
rect 1377 5865 1417 5897
rect 1449 5865 1489 5897
rect 1521 5865 1584 5897
rect 1272 5825 1584 5865
rect 1272 5793 1345 5825
rect 1377 5793 1417 5825
rect 1449 5793 1489 5825
rect 1521 5793 1584 5825
rect 1272 5753 1584 5793
rect 1272 5721 1345 5753
rect 1377 5721 1417 5753
rect 1449 5721 1489 5753
rect 1521 5721 1584 5753
rect 1272 5681 1584 5721
rect 1272 5649 1345 5681
rect 1377 5649 1417 5681
rect 1449 5649 1489 5681
rect 1521 5649 1584 5681
rect 1272 5609 1584 5649
rect 1272 5577 1345 5609
rect 1377 5577 1417 5609
rect 1449 5577 1489 5609
rect 1521 5577 1584 5609
rect 1272 5537 1584 5577
rect 1272 5505 1345 5537
rect 1377 5505 1417 5537
rect 1449 5505 1489 5537
rect 1521 5505 1584 5537
rect 1272 5465 1584 5505
rect 1272 5433 1345 5465
rect 1377 5433 1417 5465
rect 1449 5433 1489 5465
rect 1521 5433 1584 5465
rect 1272 5393 1584 5433
rect 1272 5361 1345 5393
rect 1377 5361 1417 5393
rect 1449 5361 1489 5393
rect 1521 5361 1584 5393
rect 1272 5321 1584 5361
rect 1272 5289 1345 5321
rect 1377 5289 1417 5321
rect 1449 5289 1489 5321
rect 1521 5289 1584 5321
rect 1272 5249 1584 5289
rect 1272 5217 1345 5249
rect 1377 5217 1417 5249
rect 1449 5217 1489 5249
rect 1521 5217 1584 5249
rect 1272 5177 1584 5217
rect 1272 5145 1345 5177
rect 1377 5145 1417 5177
rect 1449 5145 1489 5177
rect 1521 5145 1584 5177
rect 1272 5105 1584 5145
rect 1272 5073 1345 5105
rect 1377 5073 1417 5105
rect 1449 5073 1489 5105
rect 1521 5073 1584 5105
rect 1272 5033 1584 5073
rect 1272 5001 1345 5033
rect 1377 5001 1417 5033
rect 1449 5001 1489 5033
rect 1521 5001 1584 5033
rect 1272 4961 1584 5001
rect 1272 4929 1345 4961
rect 1377 4929 1417 4961
rect 1449 4929 1489 4961
rect 1521 4929 1584 4961
rect 1272 4889 1584 4929
rect 1272 4863 1345 4889
rect 1377 4863 1417 4889
rect 1272 4823 1312 4863
rect 1377 4857 1408 4863
rect 1449 4857 1489 4889
rect 1521 4863 1584 4889
rect 1352 4823 1408 4857
rect 1448 4823 1504 4857
rect 1544 4823 1584 4863
rect 1272 4817 1584 4823
rect 1272 4785 1345 4817
rect 1377 4785 1417 4817
rect 1449 4785 1489 4817
rect 1521 4785 1584 4817
rect 1272 4767 1584 4785
rect 1272 4727 1312 4767
rect 1352 4745 1408 4767
rect 1448 4745 1504 4767
rect 1377 4727 1408 4745
rect 1272 4713 1345 4727
rect 1377 4713 1417 4727
rect 1449 4713 1489 4745
rect 1544 4727 1584 4767
rect 1521 4713 1584 4727
rect 1272 4673 1584 4713
rect 1272 4671 1345 4673
rect 1377 4671 1417 4673
rect 1272 4631 1312 4671
rect 1377 4641 1408 4671
rect 1449 4641 1489 4673
rect 1521 4671 1584 4673
rect 1352 4631 1408 4641
rect 1448 4631 1504 4641
rect 1544 4631 1584 4671
rect 1272 4601 1584 4631
rect 1272 4575 1345 4601
rect 1377 4575 1417 4601
rect 1272 4535 1312 4575
rect 1377 4569 1408 4575
rect 1449 4569 1489 4601
rect 1521 4575 1584 4601
rect 1352 4535 1408 4569
rect 1448 4535 1504 4569
rect 1544 4535 1584 4575
rect 1272 4529 1584 4535
rect 1272 4497 1345 4529
rect 1377 4497 1417 4529
rect 1449 4497 1489 4529
rect 1521 4497 1584 4529
rect 1272 4479 1584 4497
rect 1272 4439 1312 4479
rect 1352 4457 1408 4479
rect 1448 4457 1504 4479
rect 1377 4439 1408 4457
rect 1272 4425 1345 4439
rect 1377 4425 1417 4439
rect 1449 4425 1489 4457
rect 1544 4439 1584 4479
rect 1521 4425 1584 4439
rect 1272 4385 1584 4425
rect 1272 4383 1345 4385
rect 1377 4383 1417 4385
rect 1272 4343 1312 4383
rect 1377 4353 1408 4383
rect 1449 4353 1489 4385
rect 1521 4383 1584 4385
rect 1352 4343 1408 4353
rect 1448 4343 1504 4353
rect 1544 4343 1584 4383
rect 1272 4313 1584 4343
rect 1272 4281 1345 4313
rect 1377 4281 1417 4313
rect 1449 4281 1489 4313
rect 1521 4281 1584 4313
rect 1272 4241 1584 4281
rect 1272 4209 1345 4241
rect 1377 4209 1417 4241
rect 1449 4209 1489 4241
rect 1521 4209 1584 4241
rect 1272 4169 1584 4209
rect 1272 4137 1345 4169
rect 1377 4137 1417 4169
rect 1449 4137 1489 4169
rect 1521 4137 1584 4169
rect 1272 4097 1584 4137
rect 1272 4065 1345 4097
rect 1377 4065 1417 4097
rect 1449 4065 1489 4097
rect 1521 4065 1584 4097
rect 1272 4025 1584 4065
rect 1272 3993 1345 4025
rect 1377 3993 1417 4025
rect 1449 3993 1489 4025
rect 1521 3993 1584 4025
rect 1272 3953 1584 3993
rect 1272 3921 1345 3953
rect 1377 3921 1417 3953
rect 1449 3921 1489 3953
rect 1521 3921 1584 3953
rect 1272 3881 1584 3921
rect 1272 3849 1345 3881
rect 1377 3849 1417 3881
rect 1449 3849 1489 3881
rect 1521 3849 1584 3881
rect 1272 3809 1584 3849
rect 1272 3777 1345 3809
rect 1377 3777 1417 3809
rect 1449 3777 1489 3809
rect 1521 3777 1584 3809
rect 1272 3737 1584 3777
rect 1272 3705 1345 3737
rect 1377 3705 1417 3737
rect 1449 3705 1489 3737
rect 1521 3705 1584 3737
rect 1272 3665 1584 3705
rect 1272 3633 1345 3665
rect 1377 3633 1417 3665
rect 1449 3633 1489 3665
rect 1521 3633 1584 3665
rect 1272 3593 1584 3633
rect 1272 3561 1345 3593
rect 1377 3561 1417 3593
rect 1449 3561 1489 3593
rect 1521 3561 1584 3593
rect 1272 3521 1584 3561
rect 1272 3489 1345 3521
rect 1377 3489 1417 3521
rect 1449 3489 1489 3521
rect 1521 3489 1584 3521
rect 1272 3449 1584 3489
rect 1272 3417 1345 3449
rect 1377 3417 1417 3449
rect 1449 3417 1489 3449
rect 1521 3417 1584 3449
rect 1272 3377 1584 3417
rect 1272 3345 1345 3377
rect 1377 3345 1417 3377
rect 1449 3345 1489 3377
rect 1521 3345 1584 3377
rect 1272 3305 1584 3345
rect 1272 3273 1345 3305
rect 1377 3273 1417 3305
rect 1449 3273 1489 3305
rect 1521 3273 1584 3305
rect 1272 3233 1584 3273
rect 1272 3201 1345 3233
rect 1377 3201 1417 3233
rect 1449 3201 1489 3233
rect 1521 3201 1584 3233
rect 1272 3161 1584 3201
rect 1272 3129 1345 3161
rect 1377 3129 1417 3161
rect 1449 3129 1489 3161
rect 1521 3129 1584 3161
rect 1272 3089 1584 3129
rect 1272 3063 1345 3089
rect 1377 3063 1417 3089
rect 1272 3023 1312 3063
rect 1377 3057 1408 3063
rect 1449 3057 1489 3089
rect 1521 3063 1584 3089
rect 1352 3023 1408 3057
rect 1448 3023 1504 3057
rect 1544 3023 1584 3063
rect 1272 3017 1584 3023
rect 1272 2985 1345 3017
rect 1377 2985 1417 3017
rect 1449 2985 1489 3017
rect 1521 2985 1584 3017
rect 1272 2967 1584 2985
rect 1272 2927 1312 2967
rect 1352 2945 1408 2967
rect 1448 2945 1504 2967
rect 1377 2927 1408 2945
rect 1272 2913 1345 2927
rect 1377 2913 1417 2927
rect 1449 2913 1489 2945
rect 1544 2927 1584 2967
rect 1521 2913 1584 2927
rect 1272 2873 1584 2913
rect 1272 2871 1345 2873
rect 1377 2871 1417 2873
rect 1272 2831 1312 2871
rect 1377 2841 1408 2871
rect 1449 2841 1489 2873
rect 1521 2871 1584 2873
rect 1352 2831 1408 2841
rect 1448 2831 1504 2841
rect 1544 2831 1584 2871
rect 1272 2801 1584 2831
rect 1272 2775 1345 2801
rect 1377 2775 1417 2801
rect 1272 2735 1312 2775
rect 1377 2769 1408 2775
rect 1449 2769 1489 2801
rect 1521 2775 1584 2801
rect 1352 2735 1408 2769
rect 1448 2735 1504 2769
rect 1544 2735 1584 2775
rect 1272 2729 1584 2735
rect 1272 2697 1345 2729
rect 1377 2697 1417 2729
rect 1449 2697 1489 2729
rect 1521 2697 1584 2729
rect 1272 2679 1584 2697
rect 1272 2639 1312 2679
rect 1352 2657 1408 2679
rect 1448 2657 1504 2679
rect 1377 2639 1408 2657
rect 1272 2625 1345 2639
rect 1377 2625 1417 2639
rect 1449 2625 1489 2657
rect 1544 2639 1584 2679
rect 1521 2625 1584 2639
rect 1272 2585 1584 2625
rect 1272 2583 1345 2585
rect 1377 2583 1417 2585
rect 1272 2543 1312 2583
rect 1377 2553 1408 2583
rect 1449 2553 1489 2585
rect 1521 2583 1584 2585
rect 1352 2543 1408 2553
rect 1448 2543 1504 2553
rect 1544 2543 1584 2583
rect 1272 2513 1584 2543
rect 1272 2481 1345 2513
rect 1377 2481 1417 2513
rect 1449 2481 1489 2513
rect 1521 2481 1584 2513
rect 1272 2441 1584 2481
rect 1272 2409 1345 2441
rect 1377 2409 1417 2441
rect 1449 2409 1489 2441
rect 1521 2409 1584 2441
rect 1272 2369 1584 2409
rect 1272 2337 1345 2369
rect 1377 2337 1417 2369
rect 1449 2337 1489 2369
rect 1521 2337 1584 2369
rect 1272 2297 1584 2337
rect 1272 2265 1345 2297
rect 1377 2265 1417 2297
rect 1449 2265 1489 2297
rect 1521 2265 1584 2297
rect 1272 2225 1584 2265
rect 1272 2193 1345 2225
rect 1377 2193 1417 2225
rect 1449 2193 1489 2225
rect 1521 2193 1584 2225
rect 1272 2153 1584 2193
rect 1272 2121 1345 2153
rect 1377 2121 1417 2153
rect 1449 2121 1489 2153
rect 1521 2121 1584 2153
rect 1272 2081 1584 2121
rect 1272 2049 1345 2081
rect 1377 2049 1417 2081
rect 1449 2049 1489 2081
rect 1521 2049 1584 2081
rect 1272 2009 1584 2049
rect 1272 1977 1345 2009
rect 1377 1977 1417 2009
rect 1449 1977 1489 2009
rect 1521 1977 1584 2009
rect 1272 1937 1584 1977
rect 1272 1905 1345 1937
rect 1377 1905 1417 1937
rect 1449 1905 1489 1937
rect 1521 1905 1584 1937
rect 1272 1865 1584 1905
rect 1272 1833 1345 1865
rect 1377 1833 1417 1865
rect 1449 1833 1489 1865
rect 1521 1833 1584 1865
rect 1272 1793 1584 1833
rect 1272 1761 1345 1793
rect 1377 1761 1417 1793
rect 1449 1761 1489 1793
rect 1521 1761 1584 1793
rect 1272 1721 1584 1761
rect 1272 1689 1345 1721
rect 1377 1689 1417 1721
rect 1449 1689 1489 1721
rect 1521 1689 1584 1721
rect 1272 1649 1584 1689
rect 1272 1617 1345 1649
rect 1377 1617 1417 1649
rect 1449 1617 1489 1649
rect 1521 1617 1584 1649
rect 1272 1577 1584 1617
rect 1272 1545 1345 1577
rect 1377 1545 1417 1577
rect 1449 1545 1489 1577
rect 1521 1545 1584 1577
rect 1272 1505 1584 1545
rect 1272 1473 1345 1505
rect 1377 1473 1417 1505
rect 1449 1473 1489 1505
rect 1521 1473 1584 1505
rect 1272 1433 1584 1473
rect 1272 1401 1345 1433
rect 1377 1401 1417 1433
rect 1449 1401 1489 1433
rect 1521 1401 1584 1433
rect 1272 1361 1584 1401
rect 1272 1329 1345 1361
rect 1377 1329 1417 1361
rect 1449 1329 1489 1361
rect 1521 1329 1584 1361
rect 1272 1289 1584 1329
rect 1272 1263 1345 1289
rect 1377 1263 1417 1289
rect 1272 1223 1312 1263
rect 1377 1257 1408 1263
rect 1449 1257 1489 1289
rect 1521 1263 1584 1289
rect 1352 1223 1408 1257
rect 1448 1223 1504 1257
rect 1544 1223 1584 1263
rect 1272 1217 1584 1223
rect 1272 1185 1345 1217
rect 1377 1185 1417 1217
rect 1449 1185 1489 1217
rect 1521 1185 1584 1217
rect 1272 1167 1584 1185
rect 1272 1127 1312 1167
rect 1352 1145 1408 1167
rect 1448 1145 1504 1167
rect 1377 1127 1408 1145
rect 1272 1113 1345 1127
rect 1377 1113 1417 1127
rect 1449 1113 1489 1145
rect 1544 1127 1584 1167
rect 1521 1113 1584 1127
rect 1272 1073 1584 1113
rect 1272 1071 1345 1073
rect 1377 1071 1417 1073
rect 1272 1031 1312 1071
rect 1377 1041 1408 1071
rect 1449 1041 1489 1073
rect 1521 1071 1584 1073
rect 1352 1031 1408 1041
rect 1448 1031 1504 1041
rect 1544 1031 1584 1071
rect 1272 1001 1584 1031
rect 1272 975 1345 1001
rect 1377 975 1417 1001
rect 1272 935 1312 975
rect 1377 969 1408 975
rect 1449 969 1489 1001
rect 1521 975 1584 1001
rect 1352 935 1408 969
rect 1448 935 1504 969
rect 1544 935 1584 975
rect 1272 929 1584 935
rect 1272 897 1345 929
rect 1377 897 1417 929
rect 1449 897 1489 929
rect 1521 897 1584 929
rect 1272 879 1584 897
rect 609 825 672 839
rect 366 785 672 825
rect 366 783 433 785
rect 465 783 505 785
rect 366 743 400 783
rect 465 753 496 783
rect 537 753 577 785
rect 609 783 672 785
rect 440 743 496 753
rect 536 743 592 753
rect 632 743 672 783
rect 366 713 672 743
rect 366 681 433 713
rect 465 681 505 713
rect 537 681 577 713
rect 609 681 672 713
rect 366 660 672 681
rect 1272 839 1312 879
rect 1352 857 1408 879
rect 1448 857 1504 879
rect 1377 839 1408 857
rect 1272 825 1345 839
rect 1377 825 1417 839
rect 1449 825 1489 857
rect 1544 839 1584 879
rect 1698 6466 2058 6540
rect 1698 6434 1794 6466
rect 1826 6434 1866 6466
rect 1898 6434 1938 6466
rect 1970 6434 2058 6466
rect 1698 6394 2058 6434
rect 1698 6362 1794 6394
rect 1826 6362 1866 6394
rect 1898 6362 1938 6394
rect 1970 6362 2058 6394
rect 1698 6322 2058 6362
rect 1698 6290 1794 6322
rect 1826 6290 1866 6322
rect 1898 6290 1938 6322
rect 1970 6290 2058 6322
rect 1698 6250 2058 6290
rect 1698 6218 1794 6250
rect 1826 6218 1866 6250
rect 1898 6218 1938 6250
rect 1970 6218 2058 6250
rect 1698 6178 2058 6218
rect 1698 6146 1794 6178
rect 1826 6146 1866 6178
rect 1898 6146 1938 6178
rect 1970 6146 2058 6178
rect 1698 6106 2058 6146
rect 1698 6074 1794 6106
rect 1826 6074 1866 6106
rect 1898 6074 1938 6106
rect 1970 6074 2058 6106
rect 1698 6034 2058 6074
rect 1698 6002 1794 6034
rect 1826 6002 1866 6034
rect 1898 6002 1938 6034
rect 1970 6002 2058 6034
rect 1698 5962 2058 6002
rect 1698 5930 1794 5962
rect 1826 5930 1866 5962
rect 1898 5930 1938 5962
rect 1970 5930 2058 5962
rect 1698 5890 2058 5930
rect 1698 5858 1794 5890
rect 1826 5858 1866 5890
rect 1898 5858 1938 5890
rect 1970 5858 2058 5890
rect 1698 5847 2058 5858
rect 1698 5807 1766 5847
rect 1806 5818 1862 5847
rect 1902 5818 1958 5847
rect 1826 5807 1862 5818
rect 1902 5807 1938 5818
rect 1998 5807 2058 5847
rect 1698 5786 1794 5807
rect 1826 5786 1866 5807
rect 1898 5786 1938 5807
rect 1970 5786 2058 5807
rect 1698 5751 2058 5786
rect 1698 5711 1766 5751
rect 1806 5746 1862 5751
rect 1902 5746 1958 5751
rect 1826 5714 1862 5746
rect 1902 5714 1938 5746
rect 1806 5711 1862 5714
rect 1902 5711 1958 5714
rect 1998 5711 2058 5751
rect 1698 5674 2058 5711
rect 1698 5655 1794 5674
rect 1826 5655 1866 5674
rect 1898 5655 1938 5674
rect 1970 5655 2058 5674
rect 1698 5615 1766 5655
rect 1826 5642 1862 5655
rect 1902 5642 1938 5655
rect 1806 5615 1862 5642
rect 1902 5615 1958 5642
rect 1998 5615 2058 5655
rect 1698 5602 2058 5615
rect 1698 5570 1794 5602
rect 1826 5570 1866 5602
rect 1898 5570 1938 5602
rect 1970 5570 2058 5602
rect 1698 5559 2058 5570
rect 1698 5519 1766 5559
rect 1806 5530 1862 5559
rect 1902 5530 1958 5559
rect 1826 5519 1862 5530
rect 1902 5519 1938 5530
rect 1998 5519 2058 5559
rect 1698 5498 1794 5519
rect 1826 5498 1866 5519
rect 1898 5498 1938 5519
rect 1970 5498 2058 5519
rect 1698 5463 2058 5498
rect 1698 5423 1766 5463
rect 1806 5458 1862 5463
rect 1902 5458 1958 5463
rect 1826 5426 1862 5458
rect 1902 5426 1938 5458
rect 1806 5423 1862 5426
rect 1902 5423 1958 5426
rect 1998 5423 2058 5463
rect 1698 5386 2058 5423
rect 1698 5367 1794 5386
rect 1826 5367 1866 5386
rect 1898 5367 1938 5386
rect 1970 5367 2058 5386
rect 1698 5327 1766 5367
rect 1826 5354 1862 5367
rect 1902 5354 1938 5367
rect 1806 5327 1862 5354
rect 1902 5327 1958 5354
rect 1998 5327 2058 5367
rect 1698 5314 2058 5327
rect 1698 5282 1794 5314
rect 1826 5282 1866 5314
rect 1898 5282 1938 5314
rect 1970 5282 2058 5314
rect 1698 5271 2058 5282
rect 1698 5231 1766 5271
rect 1806 5242 1862 5271
rect 1902 5242 1958 5271
rect 1826 5231 1862 5242
rect 1902 5231 1938 5242
rect 1998 5231 2058 5271
rect 1698 5210 1794 5231
rect 1826 5210 1866 5231
rect 1898 5210 1938 5231
rect 1970 5210 2058 5231
rect 1698 5175 2058 5210
rect 1698 5135 1766 5175
rect 1806 5170 1862 5175
rect 1902 5170 1958 5175
rect 1826 5138 1862 5170
rect 1902 5138 1938 5170
rect 1806 5135 1862 5138
rect 1902 5135 1958 5138
rect 1998 5135 2058 5175
rect 1698 5098 2058 5135
rect 1698 5066 1794 5098
rect 1826 5066 1866 5098
rect 1898 5066 1938 5098
rect 1970 5066 2058 5098
rect 1698 5026 2058 5066
rect 1698 4994 1794 5026
rect 1826 4994 1866 5026
rect 1898 4994 1938 5026
rect 1970 4994 2058 5026
rect 1698 4954 2058 4994
rect 1698 4922 1794 4954
rect 1826 4922 1866 4954
rect 1898 4922 1938 4954
rect 1970 4922 2058 4954
rect 1698 4882 2058 4922
rect 1698 4850 1794 4882
rect 1826 4850 1866 4882
rect 1898 4850 1938 4882
rect 1970 4850 2058 4882
rect 1698 4810 2058 4850
rect 1698 4778 1794 4810
rect 1826 4778 1866 4810
rect 1898 4778 1938 4810
rect 1970 4778 2058 4810
rect 1698 4738 2058 4778
rect 1698 4706 1794 4738
rect 1826 4706 1866 4738
rect 1898 4706 1938 4738
rect 1970 4706 2058 4738
rect 1698 4666 2058 4706
rect 1698 4634 1794 4666
rect 1826 4634 1866 4666
rect 1898 4634 1938 4666
rect 1970 4634 2058 4666
rect 1698 4594 2058 4634
rect 1698 4562 1794 4594
rect 1826 4562 1866 4594
rect 1898 4562 1938 4594
rect 1970 4562 2058 4594
rect 1698 4522 2058 4562
rect 1698 4490 1794 4522
rect 1826 4490 1866 4522
rect 1898 4490 1938 4522
rect 1970 4490 2058 4522
rect 1698 4450 2058 4490
rect 1698 4418 1794 4450
rect 1826 4418 1866 4450
rect 1898 4418 1938 4450
rect 1970 4418 2058 4450
rect 1698 4378 2058 4418
rect 1698 4346 1794 4378
rect 1826 4346 1866 4378
rect 1898 4346 1938 4378
rect 1970 4346 2058 4378
rect 1698 4306 2058 4346
rect 1698 4274 1794 4306
rect 1826 4274 1866 4306
rect 1898 4274 1938 4306
rect 1970 4274 2058 4306
rect 1698 4234 2058 4274
rect 1698 4202 1794 4234
rect 1826 4202 1866 4234
rect 1898 4202 1938 4234
rect 1970 4202 2058 4234
rect 1698 4162 2058 4202
rect 1698 4130 1794 4162
rect 1826 4130 1866 4162
rect 1898 4130 1938 4162
rect 1970 4130 2058 4162
rect 1698 4090 2058 4130
rect 1698 4058 1794 4090
rect 1826 4058 1866 4090
rect 1898 4058 1938 4090
rect 1970 4058 2058 4090
rect 1698 4047 2058 4058
rect 1698 4007 1766 4047
rect 1806 4018 1862 4047
rect 1902 4018 1958 4047
rect 1826 4007 1862 4018
rect 1902 4007 1938 4018
rect 1998 4007 2058 4047
rect 1698 3986 1794 4007
rect 1826 3986 1866 4007
rect 1898 3986 1938 4007
rect 1970 3986 2058 4007
rect 1698 3951 2058 3986
rect 1698 3911 1766 3951
rect 1806 3946 1862 3951
rect 1902 3946 1958 3951
rect 1826 3914 1862 3946
rect 1902 3914 1938 3946
rect 1806 3911 1862 3914
rect 1902 3911 1958 3914
rect 1998 3911 2058 3951
rect 1698 3874 2058 3911
rect 1698 3855 1794 3874
rect 1826 3855 1866 3874
rect 1898 3855 1938 3874
rect 1970 3855 2058 3874
rect 1698 3815 1766 3855
rect 1826 3842 1862 3855
rect 1902 3842 1938 3855
rect 1806 3815 1862 3842
rect 1902 3815 1958 3842
rect 1998 3815 2058 3855
rect 1698 3802 2058 3815
rect 1698 3770 1794 3802
rect 1826 3770 1866 3802
rect 1898 3770 1938 3802
rect 1970 3770 2058 3802
rect 1698 3759 2058 3770
rect 1698 3719 1766 3759
rect 1806 3730 1862 3759
rect 1902 3730 1958 3759
rect 1826 3719 1862 3730
rect 1902 3719 1938 3730
rect 1998 3719 2058 3759
rect 1698 3698 1794 3719
rect 1826 3698 1866 3719
rect 1898 3698 1938 3719
rect 1970 3698 2058 3719
rect 1698 3663 2058 3698
rect 1698 3623 1766 3663
rect 1806 3658 1862 3663
rect 1902 3658 1958 3663
rect 1826 3626 1862 3658
rect 1902 3626 1938 3658
rect 1806 3623 1862 3626
rect 1902 3623 1958 3626
rect 1998 3623 2058 3663
rect 1698 3586 2058 3623
rect 1698 3567 1794 3586
rect 1826 3567 1866 3586
rect 1898 3567 1938 3586
rect 1970 3567 2058 3586
rect 1698 3527 1766 3567
rect 1826 3554 1862 3567
rect 1902 3554 1938 3567
rect 1806 3527 1862 3554
rect 1902 3527 1958 3554
rect 1998 3527 2058 3567
rect 1698 3514 2058 3527
rect 1698 3482 1794 3514
rect 1826 3482 1866 3514
rect 1898 3482 1938 3514
rect 1970 3482 2058 3514
rect 1698 3471 2058 3482
rect 1698 3431 1766 3471
rect 1806 3442 1862 3471
rect 1902 3442 1958 3471
rect 1826 3431 1862 3442
rect 1902 3431 1938 3442
rect 1998 3431 2058 3471
rect 1698 3410 1794 3431
rect 1826 3410 1866 3431
rect 1898 3410 1938 3431
rect 1970 3410 2058 3431
rect 1698 3375 2058 3410
rect 1698 3335 1766 3375
rect 1806 3370 1862 3375
rect 1902 3370 1958 3375
rect 1826 3338 1862 3370
rect 1902 3338 1938 3370
rect 1806 3335 1862 3338
rect 1902 3335 1958 3338
rect 1998 3335 2058 3375
rect 1698 3298 2058 3335
rect 1698 3266 1794 3298
rect 1826 3266 1866 3298
rect 1898 3266 1938 3298
rect 1970 3266 2058 3298
rect 1698 3226 2058 3266
rect 1698 3194 1794 3226
rect 1826 3194 1866 3226
rect 1898 3194 1938 3226
rect 1970 3194 2058 3226
rect 1698 3154 2058 3194
rect 1698 3122 1794 3154
rect 1826 3122 1866 3154
rect 1898 3122 1938 3154
rect 1970 3122 2058 3154
rect 1698 3082 2058 3122
rect 1698 3050 1794 3082
rect 1826 3050 1866 3082
rect 1898 3050 1938 3082
rect 1970 3050 2058 3082
rect 1698 3010 2058 3050
rect 1698 2978 1794 3010
rect 1826 2978 1866 3010
rect 1898 2978 1938 3010
rect 1970 2978 2058 3010
rect 1698 2938 2058 2978
rect 1698 2906 1794 2938
rect 1826 2906 1866 2938
rect 1898 2906 1938 2938
rect 1970 2906 2058 2938
rect 1698 2866 2058 2906
rect 1698 2834 1794 2866
rect 1826 2834 1866 2866
rect 1898 2834 1938 2866
rect 1970 2834 2058 2866
rect 1698 2794 2058 2834
rect 1698 2762 1794 2794
rect 1826 2762 1866 2794
rect 1898 2762 1938 2794
rect 1970 2762 2058 2794
rect 1698 2722 2058 2762
rect 1698 2690 1794 2722
rect 1826 2690 1866 2722
rect 1898 2690 1938 2722
rect 1970 2690 2058 2722
rect 1698 2650 2058 2690
rect 1698 2618 1794 2650
rect 1826 2618 1866 2650
rect 1898 2618 1938 2650
rect 1970 2618 2058 2650
rect 1698 2578 2058 2618
rect 1698 2546 1794 2578
rect 1826 2546 1866 2578
rect 1898 2546 1938 2578
rect 1970 2546 2058 2578
rect 1698 2506 2058 2546
rect 1698 2474 1794 2506
rect 1826 2474 1866 2506
rect 1898 2474 1938 2506
rect 1970 2474 2058 2506
rect 1698 2434 2058 2474
rect 1698 2402 1794 2434
rect 1826 2402 1866 2434
rect 1898 2402 1938 2434
rect 1970 2402 2058 2434
rect 1698 2362 2058 2402
rect 1698 2330 1794 2362
rect 1826 2330 1866 2362
rect 1898 2330 1938 2362
rect 1970 2330 2058 2362
rect 1698 2290 2058 2330
rect 1698 2258 1794 2290
rect 1826 2258 1866 2290
rect 1898 2258 1938 2290
rect 1970 2258 2058 2290
rect 1698 2247 2058 2258
rect 1698 2207 1766 2247
rect 1806 2218 1862 2247
rect 1902 2218 1958 2247
rect 1826 2207 1862 2218
rect 1902 2207 1938 2218
rect 1998 2207 2058 2247
rect 1698 2186 1794 2207
rect 1826 2186 1866 2207
rect 1898 2186 1938 2207
rect 1970 2186 2058 2207
rect 1698 2151 2058 2186
rect 1698 2111 1766 2151
rect 1806 2146 1862 2151
rect 1902 2146 1958 2151
rect 1826 2114 1862 2146
rect 1902 2114 1938 2146
rect 1806 2111 1862 2114
rect 1902 2111 1958 2114
rect 1998 2111 2058 2151
rect 1698 2074 2058 2111
rect 1698 2055 1794 2074
rect 1826 2055 1866 2074
rect 1898 2055 1938 2074
rect 1970 2055 2058 2074
rect 1698 2015 1766 2055
rect 1826 2042 1862 2055
rect 1902 2042 1938 2055
rect 1806 2015 1862 2042
rect 1902 2015 1958 2042
rect 1998 2015 2058 2055
rect 1698 2002 2058 2015
rect 1698 1970 1794 2002
rect 1826 1970 1866 2002
rect 1898 1970 1938 2002
rect 1970 1970 2058 2002
rect 1698 1959 2058 1970
rect 1698 1919 1766 1959
rect 1806 1930 1862 1959
rect 1902 1930 1958 1959
rect 1826 1919 1862 1930
rect 1902 1919 1938 1930
rect 1998 1919 2058 1959
rect 1698 1898 1794 1919
rect 1826 1898 1866 1919
rect 1898 1898 1938 1919
rect 1970 1898 2058 1919
rect 1698 1863 2058 1898
rect 1698 1823 1766 1863
rect 1806 1858 1862 1863
rect 1902 1858 1958 1863
rect 1826 1826 1862 1858
rect 1902 1826 1938 1858
rect 1806 1823 1862 1826
rect 1902 1823 1958 1826
rect 1998 1823 2058 1863
rect 1698 1786 2058 1823
rect 1698 1767 1794 1786
rect 1826 1767 1866 1786
rect 1898 1767 1938 1786
rect 1970 1767 2058 1786
rect 1698 1727 1766 1767
rect 1826 1754 1862 1767
rect 1902 1754 1938 1767
rect 1806 1727 1862 1754
rect 1902 1727 1958 1754
rect 1998 1727 2058 1767
rect 1698 1714 2058 1727
rect 1698 1682 1794 1714
rect 1826 1682 1866 1714
rect 1898 1682 1938 1714
rect 1970 1682 2058 1714
rect 1698 1671 2058 1682
rect 1698 1631 1766 1671
rect 1806 1642 1862 1671
rect 1902 1642 1958 1671
rect 1826 1631 1862 1642
rect 1902 1631 1938 1642
rect 1998 1631 2058 1671
rect 1698 1610 1794 1631
rect 1826 1610 1866 1631
rect 1898 1610 1938 1631
rect 1970 1610 2058 1631
rect 1698 1575 2058 1610
rect 1698 1535 1766 1575
rect 1806 1570 1862 1575
rect 1902 1570 1958 1575
rect 1826 1538 1862 1570
rect 1902 1538 1938 1570
rect 1806 1535 1862 1538
rect 1902 1535 1958 1538
rect 1998 1535 2058 1575
rect 1698 1498 2058 1535
rect 1698 1466 1794 1498
rect 1826 1466 1866 1498
rect 1898 1466 1938 1498
rect 1970 1466 2058 1498
rect 1698 1426 2058 1466
rect 1698 1394 1794 1426
rect 1826 1394 1866 1426
rect 1898 1394 1938 1426
rect 1970 1394 2058 1426
rect 1698 1354 2058 1394
rect 1698 1322 1794 1354
rect 1826 1322 1866 1354
rect 1898 1322 1938 1354
rect 1970 1322 2058 1354
rect 1698 1282 2058 1322
rect 1698 1250 1794 1282
rect 1826 1250 1866 1282
rect 1898 1250 1938 1282
rect 1970 1250 2058 1282
rect 1698 1210 2058 1250
rect 1698 1178 1794 1210
rect 1826 1178 1866 1210
rect 1898 1178 1938 1210
rect 1970 1178 2058 1210
rect 1698 1138 2058 1178
rect 1698 1106 1794 1138
rect 1826 1106 1866 1138
rect 1898 1106 1938 1138
rect 1970 1106 2058 1138
rect 1698 1066 2058 1106
rect 1698 1034 1794 1066
rect 1826 1034 1866 1066
rect 1898 1034 1938 1066
rect 1970 1034 2058 1066
rect 1698 994 2058 1034
rect 1698 962 1794 994
rect 1826 962 1866 994
rect 1898 962 1938 994
rect 1970 962 2058 994
rect 1698 870 2058 962
rect 2180 6527 2224 6567
rect 2264 6545 2320 6567
rect 2360 6545 2416 6567
rect 2289 6527 2320 6545
rect 2180 6513 2257 6527
rect 2289 6513 2329 6527
rect 2361 6513 2401 6545
rect 2456 6527 2492 6567
rect 2433 6513 2492 6527
rect 2180 6473 2492 6513
rect 2180 6471 2257 6473
rect 2289 6471 2329 6473
rect 2180 6431 2224 6471
rect 2289 6441 2320 6471
rect 2361 6441 2401 6473
rect 2433 6471 2492 6473
rect 2264 6431 2320 6441
rect 2360 6431 2416 6441
rect 2456 6431 2492 6471
rect 2180 6401 2492 6431
rect 2180 6375 2257 6401
rect 2289 6375 2329 6401
rect 2180 6335 2224 6375
rect 2289 6369 2320 6375
rect 2361 6369 2401 6401
rect 2433 6375 2492 6401
rect 2264 6335 2320 6369
rect 2360 6335 2416 6369
rect 2456 6335 2492 6375
rect 2180 6329 2492 6335
rect 2180 6297 2257 6329
rect 2289 6297 2329 6329
rect 2361 6297 2401 6329
rect 2433 6297 2492 6329
rect 2180 6279 2492 6297
rect 2180 6239 2224 6279
rect 2264 6257 2320 6279
rect 2360 6257 2416 6279
rect 2289 6239 2320 6257
rect 2180 6225 2257 6239
rect 2289 6225 2329 6239
rect 2361 6225 2401 6257
rect 2456 6239 2492 6279
rect 2433 6225 2492 6239
rect 2180 6185 2492 6225
rect 2180 6183 2257 6185
rect 2289 6183 2329 6185
rect 2180 6143 2224 6183
rect 2289 6153 2320 6183
rect 2361 6153 2401 6185
rect 2433 6183 2492 6185
rect 2264 6143 2320 6153
rect 2360 6143 2416 6153
rect 2456 6143 2492 6183
rect 2180 6113 2492 6143
rect 2180 6081 2257 6113
rect 2289 6081 2329 6113
rect 2361 6081 2401 6113
rect 2433 6081 2492 6113
rect 2180 6041 2492 6081
rect 2180 6009 2257 6041
rect 2289 6009 2329 6041
rect 2361 6009 2401 6041
rect 2433 6009 2492 6041
rect 2180 5969 2492 6009
rect 2180 5937 2257 5969
rect 2289 5937 2329 5969
rect 2361 5937 2401 5969
rect 2433 5937 2492 5969
rect 2180 5897 2492 5937
rect 2180 5865 2257 5897
rect 2289 5865 2329 5897
rect 2361 5865 2401 5897
rect 2433 5865 2492 5897
rect 2180 5825 2492 5865
rect 2180 5793 2257 5825
rect 2289 5793 2329 5825
rect 2361 5793 2401 5825
rect 2433 5793 2492 5825
rect 2180 5753 2492 5793
rect 2180 5721 2257 5753
rect 2289 5721 2329 5753
rect 2361 5721 2401 5753
rect 2433 5721 2492 5753
rect 2180 5681 2492 5721
rect 2180 5649 2257 5681
rect 2289 5649 2329 5681
rect 2361 5649 2401 5681
rect 2433 5649 2492 5681
rect 2180 5609 2492 5649
rect 2180 5577 2257 5609
rect 2289 5577 2329 5609
rect 2361 5577 2401 5609
rect 2433 5577 2492 5609
rect 2180 5537 2492 5577
rect 2180 5505 2257 5537
rect 2289 5505 2329 5537
rect 2361 5505 2401 5537
rect 2433 5505 2492 5537
rect 2180 5465 2492 5505
rect 2180 5433 2257 5465
rect 2289 5433 2329 5465
rect 2361 5433 2401 5465
rect 2433 5433 2492 5465
rect 2180 5393 2492 5433
rect 2180 5361 2257 5393
rect 2289 5361 2329 5393
rect 2361 5361 2401 5393
rect 2433 5361 2492 5393
rect 2180 5321 2492 5361
rect 2180 5289 2257 5321
rect 2289 5289 2329 5321
rect 2361 5289 2401 5321
rect 2433 5289 2492 5321
rect 2180 5249 2492 5289
rect 2180 5217 2257 5249
rect 2289 5217 2329 5249
rect 2361 5217 2401 5249
rect 2433 5217 2492 5249
rect 2180 5177 2492 5217
rect 2180 5145 2257 5177
rect 2289 5145 2329 5177
rect 2361 5145 2401 5177
rect 2433 5145 2492 5177
rect 2180 5105 2492 5145
rect 2180 5073 2257 5105
rect 2289 5073 2329 5105
rect 2361 5073 2401 5105
rect 2433 5073 2492 5105
rect 2180 5033 2492 5073
rect 2180 5001 2257 5033
rect 2289 5001 2329 5033
rect 2361 5001 2401 5033
rect 2433 5001 2492 5033
rect 2180 4961 2492 5001
rect 2180 4929 2257 4961
rect 2289 4929 2329 4961
rect 2361 4929 2401 4961
rect 2433 4929 2492 4961
rect 2180 4889 2492 4929
rect 2180 4863 2257 4889
rect 2289 4863 2329 4889
rect 2180 4823 2224 4863
rect 2289 4857 2320 4863
rect 2361 4857 2401 4889
rect 2433 4863 2492 4889
rect 2264 4823 2320 4857
rect 2360 4823 2416 4857
rect 2456 4823 2492 4863
rect 2180 4817 2492 4823
rect 2180 4785 2257 4817
rect 2289 4785 2329 4817
rect 2361 4785 2401 4817
rect 2433 4785 2492 4817
rect 2180 4767 2492 4785
rect 2180 4727 2224 4767
rect 2264 4745 2320 4767
rect 2360 4745 2416 4767
rect 2289 4727 2320 4745
rect 2180 4713 2257 4727
rect 2289 4713 2329 4727
rect 2361 4713 2401 4745
rect 2456 4727 2492 4767
rect 2433 4713 2492 4727
rect 2180 4673 2492 4713
rect 2180 4671 2257 4673
rect 2289 4671 2329 4673
rect 2180 4631 2224 4671
rect 2289 4641 2320 4671
rect 2361 4641 2401 4673
rect 2433 4671 2492 4673
rect 2264 4631 2320 4641
rect 2360 4631 2416 4641
rect 2456 4631 2492 4671
rect 2180 4601 2492 4631
rect 2180 4575 2257 4601
rect 2289 4575 2329 4601
rect 2180 4535 2224 4575
rect 2289 4569 2320 4575
rect 2361 4569 2401 4601
rect 2433 4575 2492 4601
rect 2264 4535 2320 4569
rect 2360 4535 2416 4569
rect 2456 4535 2492 4575
rect 2180 4529 2492 4535
rect 2180 4497 2257 4529
rect 2289 4497 2329 4529
rect 2361 4497 2401 4529
rect 2433 4497 2492 4529
rect 2180 4479 2492 4497
rect 2180 4439 2224 4479
rect 2264 4457 2320 4479
rect 2360 4457 2416 4479
rect 2289 4439 2320 4457
rect 2180 4425 2257 4439
rect 2289 4425 2329 4439
rect 2361 4425 2401 4457
rect 2456 4439 2492 4479
rect 2433 4425 2492 4439
rect 2180 4385 2492 4425
rect 2180 4383 2257 4385
rect 2289 4383 2329 4385
rect 2180 4343 2224 4383
rect 2289 4353 2320 4383
rect 2361 4353 2401 4385
rect 2433 4383 2492 4385
rect 2264 4343 2320 4353
rect 2360 4343 2416 4353
rect 2456 4343 2492 4383
rect 2180 4313 2492 4343
rect 2180 4281 2257 4313
rect 2289 4281 2329 4313
rect 2361 4281 2401 4313
rect 2433 4281 2492 4313
rect 2180 4241 2492 4281
rect 2180 4209 2257 4241
rect 2289 4209 2329 4241
rect 2361 4209 2401 4241
rect 2433 4209 2492 4241
rect 2180 4169 2492 4209
rect 2180 4137 2257 4169
rect 2289 4137 2329 4169
rect 2361 4137 2401 4169
rect 2433 4137 2492 4169
rect 2180 4097 2492 4137
rect 2180 4065 2257 4097
rect 2289 4065 2329 4097
rect 2361 4065 2401 4097
rect 2433 4065 2492 4097
rect 2180 4025 2492 4065
rect 2180 3993 2257 4025
rect 2289 3993 2329 4025
rect 2361 3993 2401 4025
rect 2433 3993 2492 4025
rect 2180 3953 2492 3993
rect 2180 3921 2257 3953
rect 2289 3921 2329 3953
rect 2361 3921 2401 3953
rect 2433 3921 2492 3953
rect 2180 3881 2492 3921
rect 2180 3849 2257 3881
rect 2289 3849 2329 3881
rect 2361 3849 2401 3881
rect 2433 3849 2492 3881
rect 2180 3809 2492 3849
rect 2180 3777 2257 3809
rect 2289 3777 2329 3809
rect 2361 3777 2401 3809
rect 2433 3777 2492 3809
rect 2180 3737 2492 3777
rect 2180 3705 2257 3737
rect 2289 3705 2329 3737
rect 2361 3705 2401 3737
rect 2433 3705 2492 3737
rect 2180 3665 2492 3705
rect 2180 3633 2257 3665
rect 2289 3633 2329 3665
rect 2361 3633 2401 3665
rect 2433 3633 2492 3665
rect 2180 3593 2492 3633
rect 2180 3561 2257 3593
rect 2289 3561 2329 3593
rect 2361 3561 2401 3593
rect 2433 3561 2492 3593
rect 2180 3521 2492 3561
rect 2180 3489 2257 3521
rect 2289 3489 2329 3521
rect 2361 3489 2401 3521
rect 2433 3489 2492 3521
rect 2180 3449 2492 3489
rect 2180 3417 2257 3449
rect 2289 3417 2329 3449
rect 2361 3417 2401 3449
rect 2433 3417 2492 3449
rect 2180 3377 2492 3417
rect 2180 3345 2257 3377
rect 2289 3345 2329 3377
rect 2361 3345 2401 3377
rect 2433 3345 2492 3377
rect 2180 3305 2492 3345
rect 2180 3273 2257 3305
rect 2289 3273 2329 3305
rect 2361 3273 2401 3305
rect 2433 3273 2492 3305
rect 2180 3233 2492 3273
rect 2180 3201 2257 3233
rect 2289 3201 2329 3233
rect 2361 3201 2401 3233
rect 2433 3201 2492 3233
rect 2180 3161 2492 3201
rect 2180 3129 2257 3161
rect 2289 3129 2329 3161
rect 2361 3129 2401 3161
rect 2433 3129 2492 3161
rect 2180 3089 2492 3129
rect 2180 3063 2257 3089
rect 2289 3063 2329 3089
rect 2180 3023 2224 3063
rect 2289 3057 2320 3063
rect 2361 3057 2401 3089
rect 2433 3063 2492 3089
rect 2264 3023 2320 3057
rect 2360 3023 2416 3057
rect 2456 3023 2492 3063
rect 2180 3017 2492 3023
rect 2180 2985 2257 3017
rect 2289 2985 2329 3017
rect 2361 2985 2401 3017
rect 2433 2985 2492 3017
rect 2180 2967 2492 2985
rect 2180 2927 2224 2967
rect 2264 2945 2320 2967
rect 2360 2945 2416 2967
rect 2289 2927 2320 2945
rect 2180 2913 2257 2927
rect 2289 2913 2329 2927
rect 2361 2913 2401 2945
rect 2456 2927 2492 2967
rect 2433 2913 2492 2927
rect 2180 2873 2492 2913
rect 2180 2871 2257 2873
rect 2289 2871 2329 2873
rect 2180 2831 2224 2871
rect 2289 2841 2320 2871
rect 2361 2841 2401 2873
rect 2433 2871 2492 2873
rect 2264 2831 2320 2841
rect 2360 2831 2416 2841
rect 2456 2831 2492 2871
rect 2180 2801 2492 2831
rect 2180 2775 2257 2801
rect 2289 2775 2329 2801
rect 2180 2735 2224 2775
rect 2289 2769 2320 2775
rect 2361 2769 2401 2801
rect 2433 2775 2492 2801
rect 2264 2735 2320 2769
rect 2360 2735 2416 2769
rect 2456 2735 2492 2775
rect 2180 2729 2492 2735
rect 2180 2697 2257 2729
rect 2289 2697 2329 2729
rect 2361 2697 2401 2729
rect 2433 2697 2492 2729
rect 2180 2679 2492 2697
rect 2180 2639 2224 2679
rect 2264 2657 2320 2679
rect 2360 2657 2416 2679
rect 2289 2639 2320 2657
rect 2180 2625 2257 2639
rect 2289 2625 2329 2639
rect 2361 2625 2401 2657
rect 2456 2639 2492 2679
rect 2433 2625 2492 2639
rect 2180 2585 2492 2625
rect 2180 2583 2257 2585
rect 2289 2583 2329 2585
rect 2180 2543 2224 2583
rect 2289 2553 2320 2583
rect 2361 2553 2401 2585
rect 2433 2583 2492 2585
rect 2264 2543 2320 2553
rect 2360 2543 2416 2553
rect 2456 2543 2492 2583
rect 2180 2513 2492 2543
rect 2180 2481 2257 2513
rect 2289 2481 2329 2513
rect 2361 2481 2401 2513
rect 2433 2481 2492 2513
rect 2180 2441 2492 2481
rect 2180 2409 2257 2441
rect 2289 2409 2329 2441
rect 2361 2409 2401 2441
rect 2433 2409 2492 2441
rect 2180 2369 2492 2409
rect 2180 2337 2257 2369
rect 2289 2337 2329 2369
rect 2361 2337 2401 2369
rect 2433 2337 2492 2369
rect 2180 2297 2492 2337
rect 2180 2265 2257 2297
rect 2289 2265 2329 2297
rect 2361 2265 2401 2297
rect 2433 2265 2492 2297
rect 2180 2225 2492 2265
rect 2180 2193 2257 2225
rect 2289 2193 2329 2225
rect 2361 2193 2401 2225
rect 2433 2193 2492 2225
rect 2180 2153 2492 2193
rect 2180 2121 2257 2153
rect 2289 2121 2329 2153
rect 2361 2121 2401 2153
rect 2433 2121 2492 2153
rect 2180 2081 2492 2121
rect 2180 2049 2257 2081
rect 2289 2049 2329 2081
rect 2361 2049 2401 2081
rect 2433 2049 2492 2081
rect 2180 2009 2492 2049
rect 2180 1977 2257 2009
rect 2289 1977 2329 2009
rect 2361 1977 2401 2009
rect 2433 1977 2492 2009
rect 2180 1937 2492 1977
rect 2180 1905 2257 1937
rect 2289 1905 2329 1937
rect 2361 1905 2401 1937
rect 2433 1905 2492 1937
rect 2180 1865 2492 1905
rect 2180 1833 2257 1865
rect 2289 1833 2329 1865
rect 2361 1833 2401 1865
rect 2433 1833 2492 1865
rect 2180 1793 2492 1833
rect 2180 1761 2257 1793
rect 2289 1761 2329 1793
rect 2361 1761 2401 1793
rect 2433 1761 2492 1793
rect 2180 1721 2492 1761
rect 2180 1689 2257 1721
rect 2289 1689 2329 1721
rect 2361 1689 2401 1721
rect 2433 1689 2492 1721
rect 2180 1649 2492 1689
rect 2180 1617 2257 1649
rect 2289 1617 2329 1649
rect 2361 1617 2401 1649
rect 2433 1617 2492 1649
rect 2180 1577 2492 1617
rect 2180 1545 2257 1577
rect 2289 1545 2329 1577
rect 2361 1545 2401 1577
rect 2433 1545 2492 1577
rect 2180 1505 2492 1545
rect 2180 1473 2257 1505
rect 2289 1473 2329 1505
rect 2361 1473 2401 1505
rect 2433 1473 2492 1505
rect 2180 1433 2492 1473
rect 2180 1401 2257 1433
rect 2289 1401 2329 1433
rect 2361 1401 2401 1433
rect 2433 1401 2492 1433
rect 2180 1361 2492 1401
rect 2180 1329 2257 1361
rect 2289 1329 2329 1361
rect 2361 1329 2401 1361
rect 2433 1329 2492 1361
rect 2180 1289 2492 1329
rect 2180 1263 2257 1289
rect 2289 1263 2329 1289
rect 2180 1223 2224 1263
rect 2289 1257 2320 1263
rect 2361 1257 2401 1289
rect 2433 1263 2492 1289
rect 2264 1223 2320 1257
rect 2360 1223 2416 1257
rect 2456 1223 2492 1263
rect 2180 1217 2492 1223
rect 2180 1185 2257 1217
rect 2289 1185 2329 1217
rect 2361 1185 2401 1217
rect 2433 1185 2492 1217
rect 2180 1167 2492 1185
rect 2180 1127 2224 1167
rect 2264 1145 2320 1167
rect 2360 1145 2416 1167
rect 2289 1127 2320 1145
rect 2180 1113 2257 1127
rect 2289 1113 2329 1127
rect 2361 1113 2401 1145
rect 2456 1127 2492 1167
rect 2433 1113 2492 1127
rect 2180 1073 2492 1113
rect 2180 1071 2257 1073
rect 2289 1071 2329 1073
rect 2180 1031 2224 1071
rect 2289 1041 2320 1071
rect 2361 1041 2401 1073
rect 2433 1071 2492 1073
rect 2264 1031 2320 1041
rect 2360 1031 2416 1041
rect 2456 1031 2492 1071
rect 2180 1001 2492 1031
rect 2180 975 2257 1001
rect 2289 975 2329 1001
rect 2180 935 2224 975
rect 2289 969 2320 975
rect 2361 969 2401 1001
rect 2433 975 2492 1001
rect 2264 935 2320 969
rect 2360 935 2416 969
rect 2456 935 2492 975
rect 2180 929 2492 935
rect 2180 897 2257 929
rect 2289 897 2329 929
rect 2361 897 2401 929
rect 2433 897 2492 929
rect 2180 879 2492 897
rect 1521 825 1584 839
rect 1272 785 1584 825
rect 1272 783 1345 785
rect 1377 783 1417 785
rect 1272 743 1312 783
rect 1377 753 1408 783
rect 1449 753 1489 785
rect 1521 783 1584 785
rect 1352 743 1408 753
rect 1448 743 1504 753
rect 1544 743 1584 783
rect 1272 713 1584 743
rect 1272 681 1345 713
rect 1377 681 1417 713
rect 1449 681 1489 713
rect 1521 681 1584 713
rect 1272 660 1584 681
rect 2180 839 2224 879
rect 2264 857 2320 879
rect 2360 857 2416 879
rect 2289 839 2320 857
rect 2180 825 2257 839
rect 2289 825 2329 839
rect 2361 825 2401 857
rect 2456 839 2492 879
rect 2433 825 2492 839
rect 2180 785 2492 825
rect 2180 783 2257 785
rect 2289 783 2329 785
rect 2180 743 2224 783
rect 2289 753 2320 783
rect 2361 753 2401 785
rect 2433 783 2492 785
rect 2264 743 2320 753
rect 2360 743 2416 753
rect 2456 743 2492 783
rect 2180 713 2492 743
rect 2180 681 2257 713
rect 2289 681 2329 713
rect 2361 681 2401 713
rect 2433 681 2492 713
rect 2180 660 2492 681
rect 366 614 2492 660
rect 366 582 447 614
rect 479 582 519 614
rect 551 582 591 614
rect 623 582 663 614
rect 695 582 735 614
rect 767 582 807 614
rect 839 582 879 614
rect 911 582 951 614
rect 983 582 1023 614
rect 1055 582 1095 614
rect 1127 582 1167 614
rect 1199 582 1239 614
rect 1271 582 1311 614
rect 1343 582 1383 614
rect 1415 582 1455 614
rect 1487 582 1527 614
rect 1559 582 1599 614
rect 1631 582 1671 614
rect 1703 582 1743 614
rect 1775 582 1815 614
rect 1847 582 1887 614
rect 1919 582 1959 614
rect 1991 582 2031 614
rect 2063 582 2103 614
rect 2135 582 2175 614
rect 2207 582 2247 614
rect 2279 582 2319 614
rect 2351 582 2391 614
rect 2423 582 2492 614
rect 366 542 2492 582
rect 366 510 447 542
rect 479 510 519 542
rect 551 510 591 542
rect 623 510 663 542
rect 695 510 735 542
rect 767 510 807 542
rect 839 510 879 542
rect 911 510 951 542
rect 983 510 1023 542
rect 1055 510 1095 542
rect 1127 510 1167 542
rect 1199 510 1239 542
rect 1271 510 1311 542
rect 1343 510 1383 542
rect 1415 510 1455 542
rect 1487 510 1527 542
rect 1559 510 1599 542
rect 1631 510 1671 542
rect 1703 510 1743 542
rect 1775 510 1815 542
rect 1847 510 1887 542
rect 1919 510 1959 542
rect 1991 510 2031 542
rect 2063 510 2103 542
rect 2135 510 2175 542
rect 2207 510 2247 542
rect 2279 510 2319 542
rect 2351 510 2391 542
rect 2423 510 2492 542
rect 366 470 2492 510
rect 366 438 447 470
rect 479 438 519 470
rect 551 438 591 470
rect 623 438 663 470
rect 695 438 735 470
rect 767 438 807 470
rect 839 438 879 470
rect 911 438 951 470
rect 983 438 1023 470
rect 1055 438 1095 470
rect 1127 438 1167 470
rect 1199 438 1239 470
rect 1271 438 1311 470
rect 1343 438 1383 470
rect 1415 438 1455 470
rect 1487 438 1527 470
rect 1559 438 1599 470
rect 1631 438 1671 470
rect 1703 438 1743 470
rect 1775 438 1815 470
rect 1847 438 1887 470
rect 1919 438 1959 470
rect 1991 438 2031 470
rect 2063 438 2103 470
rect 2135 438 2175 470
rect 2207 438 2247 470
rect 2279 438 2319 470
rect 2351 438 2391 470
rect 2423 438 2492 470
rect 366 378 2492 438
rect 2600 7021 2864 7061
rect 2600 6989 2708 7021
rect 2740 6989 2864 7021
rect 2600 6949 2864 6989
rect 2600 6917 2708 6949
rect 2740 6917 2864 6949
rect 2600 6877 2864 6917
rect 2600 6845 2708 6877
rect 2740 6845 2864 6877
rect 2600 6805 2864 6845
rect 2600 6773 2708 6805
rect 2740 6773 2864 6805
rect 2600 6733 2864 6773
rect 2600 6701 2708 6733
rect 2740 6701 2864 6733
rect 2600 6661 2864 6701
rect 2600 6629 2708 6661
rect 2740 6629 2864 6661
rect 2600 6589 2864 6629
rect 2600 6557 2708 6589
rect 2740 6557 2864 6589
rect 2600 6517 2864 6557
rect 2600 6485 2708 6517
rect 2740 6485 2864 6517
rect 2600 6445 2864 6485
rect 2600 6413 2708 6445
rect 2740 6413 2864 6445
rect 2600 6373 2864 6413
rect 2600 6341 2708 6373
rect 2740 6341 2864 6373
rect 2600 6301 2864 6341
rect 2600 6269 2708 6301
rect 2740 6269 2864 6301
rect 2600 6229 2864 6269
rect 2600 6197 2708 6229
rect 2740 6197 2864 6229
rect 2600 6157 2864 6197
rect 2600 6125 2708 6157
rect 2740 6125 2864 6157
rect 2600 6085 2864 6125
rect 2600 6053 2708 6085
rect 2740 6053 2864 6085
rect 2600 6013 2864 6053
rect 2600 5981 2708 6013
rect 2740 5981 2864 6013
rect 2600 5941 2864 5981
rect 2600 5909 2708 5941
rect 2740 5909 2864 5941
rect 2600 5869 2864 5909
rect 2600 5837 2708 5869
rect 2740 5837 2864 5869
rect 2600 5797 2864 5837
rect 2600 5765 2708 5797
rect 2740 5765 2864 5797
rect 2600 5725 2864 5765
rect 2600 5693 2708 5725
rect 2740 5693 2864 5725
rect 2600 5653 2864 5693
rect 2600 5621 2708 5653
rect 2740 5621 2864 5653
rect 2600 5581 2864 5621
rect 2600 5549 2708 5581
rect 2740 5549 2864 5581
rect 2600 5509 2864 5549
rect 2600 5477 2708 5509
rect 2740 5477 2864 5509
rect 2600 5437 2864 5477
rect 2600 5405 2708 5437
rect 2740 5405 2864 5437
rect 2600 5365 2864 5405
rect 2600 5333 2708 5365
rect 2740 5333 2864 5365
rect 2600 5293 2864 5333
rect 2600 5261 2708 5293
rect 2740 5261 2864 5293
rect 2600 5221 2864 5261
rect 2600 5189 2708 5221
rect 2740 5189 2864 5221
rect 2600 5149 2864 5189
rect 2600 5117 2708 5149
rect 2740 5117 2864 5149
rect 2600 5077 2864 5117
rect 2600 5045 2708 5077
rect 2740 5045 2864 5077
rect 2600 5005 2864 5045
rect 2600 4973 2708 5005
rect 2740 4973 2864 5005
rect 2600 4933 2864 4973
rect 2600 4901 2708 4933
rect 2740 4901 2864 4933
rect 2600 4861 2864 4901
rect 2600 4829 2708 4861
rect 2740 4829 2864 4861
rect 2600 4789 2864 4829
rect 2600 4757 2708 4789
rect 2740 4757 2864 4789
rect 2600 4717 2864 4757
rect 2600 4685 2708 4717
rect 2740 4685 2864 4717
rect 2600 4645 2864 4685
rect 2600 4613 2708 4645
rect 2740 4613 2864 4645
rect 2600 4573 2864 4613
rect 2600 4541 2708 4573
rect 2740 4541 2864 4573
rect 2600 4501 2864 4541
rect 2600 4469 2708 4501
rect 2740 4469 2864 4501
rect 2600 4429 2864 4469
rect 2600 4397 2708 4429
rect 2740 4397 2864 4429
rect 2600 4357 2864 4397
rect 2600 4325 2708 4357
rect 2740 4325 2864 4357
rect 2600 4285 2864 4325
rect 2600 4253 2708 4285
rect 2740 4253 2864 4285
rect 2600 4213 2864 4253
rect 2600 4181 2708 4213
rect 2740 4181 2864 4213
rect 2600 4141 2864 4181
rect 2600 4109 2708 4141
rect 2740 4109 2864 4141
rect 2600 4069 2864 4109
rect 2600 4037 2708 4069
rect 2740 4037 2864 4069
rect 2600 3997 2864 4037
rect 2600 3965 2708 3997
rect 2740 3965 2864 3997
rect 2600 3925 2864 3965
rect 2600 3893 2708 3925
rect 2740 3893 2864 3925
rect 2600 3853 2864 3893
rect 2600 3821 2708 3853
rect 2740 3821 2864 3853
rect 2600 3781 2864 3821
rect 2600 3749 2708 3781
rect 2740 3749 2864 3781
rect 2600 3709 2864 3749
rect 2600 3677 2708 3709
rect 2740 3677 2864 3709
rect 2600 3637 2864 3677
rect 2600 3605 2708 3637
rect 2740 3605 2864 3637
rect 2600 3565 2864 3605
rect 2600 3533 2708 3565
rect 2740 3533 2864 3565
rect 2600 3493 2864 3533
rect 2600 3461 2708 3493
rect 2740 3461 2864 3493
rect 2600 3421 2864 3461
rect 2600 3389 2708 3421
rect 2740 3389 2864 3421
rect 2600 3349 2864 3389
rect 2600 3317 2708 3349
rect 2740 3317 2864 3349
rect 2600 3277 2864 3317
rect 2600 3245 2708 3277
rect 2740 3245 2864 3277
rect 2600 3205 2864 3245
rect 2600 3173 2708 3205
rect 2740 3173 2864 3205
rect 2600 3133 2864 3173
rect 2600 3101 2708 3133
rect 2740 3101 2864 3133
rect 2600 3061 2864 3101
rect 2600 3029 2708 3061
rect 2740 3029 2864 3061
rect 2600 2989 2864 3029
rect 2600 2957 2708 2989
rect 2740 2957 2864 2989
rect 2600 2917 2864 2957
rect 2600 2885 2708 2917
rect 2740 2885 2864 2917
rect 2600 2845 2864 2885
rect 2600 2813 2708 2845
rect 2740 2813 2864 2845
rect 2600 2773 2864 2813
rect 2600 2741 2708 2773
rect 2740 2741 2864 2773
rect 2600 2701 2864 2741
rect 2600 2669 2708 2701
rect 2740 2669 2864 2701
rect 2600 2629 2864 2669
rect 2600 2597 2708 2629
rect 2740 2597 2864 2629
rect 2600 2557 2864 2597
rect 2600 2525 2708 2557
rect 2740 2525 2864 2557
rect 2600 2485 2864 2525
rect 2600 2453 2708 2485
rect 2740 2453 2864 2485
rect 2600 2413 2864 2453
rect 2600 2381 2708 2413
rect 2740 2381 2864 2413
rect 2600 2341 2864 2381
rect 2600 2309 2708 2341
rect 2740 2309 2864 2341
rect 2600 2269 2864 2309
rect 2600 2237 2708 2269
rect 2740 2237 2864 2269
rect 2600 2197 2864 2237
rect 2600 2165 2708 2197
rect 2740 2165 2864 2197
rect 2600 2125 2864 2165
rect 2600 2093 2708 2125
rect 2740 2093 2864 2125
rect 2600 2053 2864 2093
rect 2600 2021 2708 2053
rect 2740 2021 2864 2053
rect 2600 1981 2864 2021
rect 2600 1949 2708 1981
rect 2740 1949 2864 1981
rect 2600 1909 2864 1949
rect 2600 1877 2708 1909
rect 2740 1877 2864 1909
rect 2600 1837 2864 1877
rect 2600 1805 2708 1837
rect 2740 1805 2864 1837
rect 2600 1765 2864 1805
rect 2600 1733 2708 1765
rect 2740 1733 2864 1765
rect 2600 1693 2864 1733
rect 2600 1661 2708 1693
rect 2740 1661 2864 1693
rect 2600 1621 2864 1661
rect 2600 1589 2708 1621
rect 2740 1589 2864 1621
rect 2600 1549 2864 1589
rect 2600 1517 2708 1549
rect 2740 1517 2864 1549
rect 2600 1477 2864 1517
rect 2600 1445 2708 1477
rect 2740 1445 2864 1477
rect 2600 1405 2864 1445
rect 2600 1373 2708 1405
rect 2740 1373 2864 1405
rect 2600 1333 2864 1373
rect 2600 1301 2708 1333
rect 2740 1301 2864 1333
rect 2600 1261 2864 1301
rect 2600 1229 2708 1261
rect 2740 1229 2864 1261
rect 2600 1189 2864 1229
rect 2600 1157 2708 1189
rect 2740 1157 2864 1189
rect 2600 1117 2864 1157
rect 2600 1085 2708 1117
rect 2740 1085 2864 1117
rect 2600 1045 2864 1085
rect 2600 1013 2708 1045
rect 2740 1013 2864 1045
rect 2600 973 2864 1013
rect 2600 941 2708 973
rect 2740 941 2864 973
rect 2600 901 2864 941
rect 2600 869 2708 901
rect 2740 869 2864 901
rect 2600 829 2864 869
rect 2600 797 2708 829
rect 2740 797 2864 829
rect 2600 757 2864 797
rect 2600 725 2708 757
rect 2740 725 2864 757
rect 2600 685 2864 725
rect 2600 653 2708 685
rect 2740 653 2864 685
rect 2600 613 2864 653
rect 2600 581 2708 613
rect 2740 581 2864 613
rect 2600 541 2864 581
rect 2600 509 2708 541
rect 2740 509 2864 541
rect 2600 469 2864 509
rect 2600 437 2708 469
rect 2740 437 2864 469
rect 2600 397 2864 437
rect 0 325 270 365
rect 0 293 116 325
rect 148 293 270 325
rect 0 270 270 293
rect 2600 365 2708 397
rect 2740 365 2864 397
rect 2600 325 2864 365
rect 2600 293 2708 325
rect 2740 293 2864 325
rect 2600 270 2864 293
rect 0 253 2864 270
rect 0 221 116 253
rect 148 221 2708 253
rect 2740 221 2864 253
rect 0 154 2864 221
rect 0 122 124 154
rect 156 122 196 154
rect 228 122 268 154
rect 300 122 340 154
rect 372 122 412 154
rect 444 122 484 154
rect 516 122 556 154
rect 588 122 628 154
rect 660 122 700 154
rect 732 122 772 154
rect 804 122 844 154
rect 876 122 916 154
rect 948 122 988 154
rect 1020 122 1060 154
rect 1092 122 1132 154
rect 1164 122 1204 154
rect 1236 122 1276 154
rect 1308 122 1348 154
rect 1380 122 1420 154
rect 1452 122 1492 154
rect 1524 122 1564 154
rect 1596 122 1636 154
rect 1668 122 1708 154
rect 1740 122 1780 154
rect 1812 122 1852 154
rect 1884 122 1924 154
rect 1956 122 1996 154
rect 2028 122 2068 154
rect 2100 122 2140 154
rect 2172 122 2212 154
rect 2244 122 2284 154
rect 2316 122 2356 154
rect 2388 122 2428 154
rect 2460 122 2500 154
rect 2532 122 2572 154
rect 2604 122 2644 154
rect 2676 122 2716 154
rect 2748 122 2864 154
rect 0 0 2864 122
<< via1 >>
rect 400 6657 433 6663
rect 433 6657 440 6663
rect 496 6657 505 6663
rect 505 6657 536 6663
rect 592 6657 609 6663
rect 609 6657 632 6663
rect 400 6623 440 6657
rect 496 6623 536 6657
rect 592 6623 632 6657
rect 400 6545 440 6567
rect 496 6545 536 6567
rect 592 6545 632 6567
rect 400 6527 433 6545
rect 433 6527 440 6545
rect 496 6527 505 6545
rect 505 6527 536 6545
rect 592 6527 609 6545
rect 609 6527 632 6545
rect 1312 6657 1345 6663
rect 1345 6657 1352 6663
rect 1408 6657 1417 6663
rect 1417 6657 1448 6663
rect 1504 6657 1521 6663
rect 1521 6657 1544 6663
rect 1312 6623 1352 6657
rect 1408 6623 1448 6657
rect 1504 6623 1544 6657
rect 400 6441 433 6471
rect 433 6441 440 6471
rect 496 6441 505 6471
rect 505 6441 536 6471
rect 592 6441 609 6471
rect 609 6441 632 6471
rect 400 6431 440 6441
rect 496 6431 536 6441
rect 592 6431 632 6441
rect 400 6369 433 6375
rect 433 6369 440 6375
rect 496 6369 505 6375
rect 505 6369 536 6375
rect 592 6369 609 6375
rect 609 6369 632 6375
rect 400 6335 440 6369
rect 496 6335 536 6369
rect 592 6335 632 6369
rect 400 6257 440 6279
rect 496 6257 536 6279
rect 592 6257 632 6279
rect 400 6239 433 6257
rect 433 6239 440 6257
rect 496 6239 505 6257
rect 505 6239 536 6257
rect 592 6239 609 6257
rect 609 6239 632 6257
rect 400 6153 433 6183
rect 433 6153 440 6183
rect 496 6153 505 6183
rect 505 6153 536 6183
rect 592 6153 609 6183
rect 609 6153 632 6183
rect 400 6143 440 6153
rect 496 6143 536 6153
rect 592 6143 632 6153
rect 400 4857 433 4863
rect 433 4857 440 4863
rect 496 4857 505 4863
rect 505 4857 536 4863
rect 592 4857 609 4863
rect 609 4857 632 4863
rect 400 4823 440 4857
rect 496 4823 536 4857
rect 592 4823 632 4857
rect 400 4745 440 4767
rect 496 4745 536 4767
rect 592 4745 632 4767
rect 400 4727 433 4745
rect 433 4727 440 4745
rect 496 4727 505 4745
rect 505 4727 536 4745
rect 592 4727 609 4745
rect 609 4727 632 4745
rect 400 4641 433 4671
rect 433 4641 440 4671
rect 496 4641 505 4671
rect 505 4641 536 4671
rect 592 4641 609 4671
rect 609 4641 632 4671
rect 400 4631 440 4641
rect 496 4631 536 4641
rect 592 4631 632 4641
rect 400 4569 433 4575
rect 433 4569 440 4575
rect 496 4569 505 4575
rect 505 4569 536 4575
rect 592 4569 609 4575
rect 609 4569 632 4575
rect 400 4535 440 4569
rect 496 4535 536 4569
rect 592 4535 632 4569
rect 400 4457 440 4479
rect 496 4457 536 4479
rect 592 4457 632 4479
rect 400 4439 433 4457
rect 433 4439 440 4457
rect 496 4439 505 4457
rect 505 4439 536 4457
rect 592 4439 609 4457
rect 609 4439 632 4457
rect 400 4353 433 4383
rect 433 4353 440 4383
rect 496 4353 505 4383
rect 505 4353 536 4383
rect 592 4353 609 4383
rect 609 4353 632 4383
rect 400 4343 440 4353
rect 496 4343 536 4353
rect 592 4343 632 4353
rect 400 3057 433 3063
rect 433 3057 440 3063
rect 496 3057 505 3063
rect 505 3057 536 3063
rect 592 3057 609 3063
rect 609 3057 632 3063
rect 400 3023 440 3057
rect 496 3023 536 3057
rect 592 3023 632 3057
rect 400 2945 440 2967
rect 496 2945 536 2967
rect 592 2945 632 2967
rect 400 2927 433 2945
rect 433 2927 440 2945
rect 496 2927 505 2945
rect 505 2927 536 2945
rect 592 2927 609 2945
rect 609 2927 632 2945
rect 400 2841 433 2871
rect 433 2841 440 2871
rect 496 2841 505 2871
rect 505 2841 536 2871
rect 592 2841 609 2871
rect 609 2841 632 2871
rect 400 2831 440 2841
rect 496 2831 536 2841
rect 592 2831 632 2841
rect 400 2769 433 2775
rect 433 2769 440 2775
rect 496 2769 505 2775
rect 505 2769 536 2775
rect 592 2769 609 2775
rect 609 2769 632 2775
rect 400 2735 440 2769
rect 496 2735 536 2769
rect 592 2735 632 2769
rect 400 2657 440 2679
rect 496 2657 536 2679
rect 592 2657 632 2679
rect 400 2639 433 2657
rect 433 2639 440 2657
rect 496 2639 505 2657
rect 505 2639 536 2657
rect 592 2639 609 2657
rect 609 2639 632 2657
rect 400 2553 433 2583
rect 433 2553 440 2583
rect 496 2553 505 2583
rect 505 2553 536 2583
rect 592 2553 609 2583
rect 609 2553 632 2583
rect 400 2543 440 2553
rect 496 2543 536 2553
rect 592 2543 632 2553
rect 400 1257 433 1263
rect 433 1257 440 1263
rect 496 1257 505 1263
rect 505 1257 536 1263
rect 592 1257 609 1263
rect 609 1257 632 1263
rect 400 1223 440 1257
rect 496 1223 536 1257
rect 592 1223 632 1257
rect 400 1145 440 1167
rect 496 1145 536 1167
rect 592 1145 632 1167
rect 400 1127 433 1145
rect 433 1127 440 1145
rect 496 1127 505 1145
rect 505 1127 536 1145
rect 592 1127 609 1145
rect 609 1127 632 1145
rect 400 1041 433 1071
rect 433 1041 440 1071
rect 496 1041 505 1071
rect 505 1041 536 1071
rect 592 1041 609 1071
rect 609 1041 632 1071
rect 400 1031 440 1041
rect 496 1031 536 1041
rect 592 1031 632 1041
rect 400 969 433 975
rect 433 969 440 975
rect 496 969 505 975
rect 505 969 536 975
rect 592 969 609 975
rect 609 969 632 975
rect 400 935 440 969
rect 496 935 536 969
rect 592 935 632 969
rect 400 857 440 879
rect 496 857 536 879
rect 592 857 632 879
rect 400 839 433 857
rect 433 839 440 857
rect 496 839 505 857
rect 505 839 536 857
rect 592 839 609 857
rect 609 839 632 857
rect 860 5818 900 5847
rect 956 5818 996 5847
rect 1052 5818 1092 5847
rect 860 5807 888 5818
rect 888 5807 900 5818
rect 956 5807 960 5818
rect 960 5807 992 5818
rect 992 5807 996 5818
rect 1052 5807 1064 5818
rect 1064 5807 1092 5818
rect 860 5746 900 5751
rect 956 5746 996 5751
rect 1052 5746 1092 5751
rect 860 5714 888 5746
rect 888 5714 900 5746
rect 956 5714 960 5746
rect 960 5714 992 5746
rect 992 5714 996 5746
rect 1052 5714 1064 5746
rect 1064 5714 1092 5746
rect 860 5711 900 5714
rect 956 5711 996 5714
rect 1052 5711 1092 5714
rect 860 5642 888 5655
rect 888 5642 900 5655
rect 956 5642 960 5655
rect 960 5642 992 5655
rect 992 5642 996 5655
rect 1052 5642 1064 5655
rect 1064 5642 1092 5655
rect 860 5615 900 5642
rect 956 5615 996 5642
rect 1052 5615 1092 5642
rect 860 5530 900 5559
rect 956 5530 996 5559
rect 1052 5530 1092 5559
rect 860 5519 888 5530
rect 888 5519 900 5530
rect 956 5519 960 5530
rect 960 5519 992 5530
rect 992 5519 996 5530
rect 1052 5519 1064 5530
rect 1064 5519 1092 5530
rect 860 5458 900 5463
rect 956 5458 996 5463
rect 1052 5458 1092 5463
rect 860 5426 888 5458
rect 888 5426 900 5458
rect 956 5426 960 5458
rect 960 5426 992 5458
rect 992 5426 996 5458
rect 1052 5426 1064 5458
rect 1064 5426 1092 5458
rect 860 5423 900 5426
rect 956 5423 996 5426
rect 1052 5423 1092 5426
rect 860 5354 888 5367
rect 888 5354 900 5367
rect 956 5354 960 5367
rect 960 5354 992 5367
rect 992 5354 996 5367
rect 1052 5354 1064 5367
rect 1064 5354 1092 5367
rect 860 5327 900 5354
rect 956 5327 996 5354
rect 1052 5327 1092 5354
rect 860 5242 900 5271
rect 956 5242 996 5271
rect 1052 5242 1092 5271
rect 860 5231 888 5242
rect 888 5231 900 5242
rect 956 5231 960 5242
rect 960 5231 992 5242
rect 992 5231 996 5242
rect 1052 5231 1064 5242
rect 1064 5231 1092 5242
rect 860 5170 900 5175
rect 956 5170 996 5175
rect 1052 5170 1092 5175
rect 860 5138 888 5170
rect 888 5138 900 5170
rect 956 5138 960 5170
rect 960 5138 992 5170
rect 992 5138 996 5170
rect 1052 5138 1064 5170
rect 1064 5138 1092 5170
rect 860 5135 900 5138
rect 956 5135 996 5138
rect 1052 5135 1092 5138
rect 860 4018 900 4047
rect 956 4018 996 4047
rect 1052 4018 1092 4047
rect 860 4007 888 4018
rect 888 4007 900 4018
rect 956 4007 960 4018
rect 960 4007 992 4018
rect 992 4007 996 4018
rect 1052 4007 1064 4018
rect 1064 4007 1092 4018
rect 860 3946 900 3951
rect 956 3946 996 3951
rect 1052 3946 1092 3951
rect 860 3914 888 3946
rect 888 3914 900 3946
rect 956 3914 960 3946
rect 960 3914 992 3946
rect 992 3914 996 3946
rect 1052 3914 1064 3946
rect 1064 3914 1092 3946
rect 860 3911 900 3914
rect 956 3911 996 3914
rect 1052 3911 1092 3914
rect 860 3842 888 3855
rect 888 3842 900 3855
rect 956 3842 960 3855
rect 960 3842 992 3855
rect 992 3842 996 3855
rect 1052 3842 1064 3855
rect 1064 3842 1092 3855
rect 860 3815 900 3842
rect 956 3815 996 3842
rect 1052 3815 1092 3842
rect 860 3730 900 3759
rect 956 3730 996 3759
rect 1052 3730 1092 3759
rect 860 3719 888 3730
rect 888 3719 900 3730
rect 956 3719 960 3730
rect 960 3719 992 3730
rect 992 3719 996 3730
rect 1052 3719 1064 3730
rect 1064 3719 1092 3730
rect 860 3658 900 3663
rect 956 3658 996 3663
rect 1052 3658 1092 3663
rect 860 3626 888 3658
rect 888 3626 900 3658
rect 956 3626 960 3658
rect 960 3626 992 3658
rect 992 3626 996 3658
rect 1052 3626 1064 3658
rect 1064 3626 1092 3658
rect 860 3623 900 3626
rect 956 3623 996 3626
rect 1052 3623 1092 3626
rect 860 3554 888 3567
rect 888 3554 900 3567
rect 956 3554 960 3567
rect 960 3554 992 3567
rect 992 3554 996 3567
rect 1052 3554 1064 3567
rect 1064 3554 1092 3567
rect 860 3527 900 3554
rect 956 3527 996 3554
rect 1052 3527 1092 3554
rect 860 3442 900 3471
rect 956 3442 996 3471
rect 1052 3442 1092 3471
rect 860 3431 888 3442
rect 888 3431 900 3442
rect 956 3431 960 3442
rect 960 3431 992 3442
rect 992 3431 996 3442
rect 1052 3431 1064 3442
rect 1064 3431 1092 3442
rect 860 3370 900 3375
rect 956 3370 996 3375
rect 1052 3370 1092 3375
rect 860 3338 888 3370
rect 888 3338 900 3370
rect 956 3338 960 3370
rect 960 3338 992 3370
rect 992 3338 996 3370
rect 1052 3338 1064 3370
rect 1064 3338 1092 3370
rect 860 3335 900 3338
rect 956 3335 996 3338
rect 1052 3335 1092 3338
rect 860 2218 900 2247
rect 956 2218 996 2247
rect 1052 2218 1092 2247
rect 860 2207 888 2218
rect 888 2207 900 2218
rect 956 2207 960 2218
rect 960 2207 992 2218
rect 992 2207 996 2218
rect 1052 2207 1064 2218
rect 1064 2207 1092 2218
rect 860 2146 900 2151
rect 956 2146 996 2151
rect 1052 2146 1092 2151
rect 860 2114 888 2146
rect 888 2114 900 2146
rect 956 2114 960 2146
rect 960 2114 992 2146
rect 992 2114 996 2146
rect 1052 2114 1064 2146
rect 1064 2114 1092 2146
rect 860 2111 900 2114
rect 956 2111 996 2114
rect 1052 2111 1092 2114
rect 860 2042 888 2055
rect 888 2042 900 2055
rect 956 2042 960 2055
rect 960 2042 992 2055
rect 992 2042 996 2055
rect 1052 2042 1064 2055
rect 1064 2042 1092 2055
rect 860 2015 900 2042
rect 956 2015 996 2042
rect 1052 2015 1092 2042
rect 860 1930 900 1959
rect 956 1930 996 1959
rect 1052 1930 1092 1959
rect 860 1919 888 1930
rect 888 1919 900 1930
rect 956 1919 960 1930
rect 960 1919 992 1930
rect 992 1919 996 1930
rect 1052 1919 1064 1930
rect 1064 1919 1092 1930
rect 860 1858 900 1863
rect 956 1858 996 1863
rect 1052 1858 1092 1863
rect 860 1826 888 1858
rect 888 1826 900 1858
rect 956 1826 960 1858
rect 960 1826 992 1858
rect 992 1826 996 1858
rect 1052 1826 1064 1858
rect 1064 1826 1092 1858
rect 860 1823 900 1826
rect 956 1823 996 1826
rect 1052 1823 1092 1826
rect 860 1754 888 1767
rect 888 1754 900 1767
rect 956 1754 960 1767
rect 960 1754 992 1767
rect 992 1754 996 1767
rect 1052 1754 1064 1767
rect 1064 1754 1092 1767
rect 860 1727 900 1754
rect 956 1727 996 1754
rect 1052 1727 1092 1754
rect 860 1642 900 1671
rect 956 1642 996 1671
rect 1052 1642 1092 1671
rect 860 1631 888 1642
rect 888 1631 900 1642
rect 956 1631 960 1642
rect 960 1631 992 1642
rect 992 1631 996 1642
rect 1052 1631 1064 1642
rect 1064 1631 1092 1642
rect 860 1570 900 1575
rect 956 1570 996 1575
rect 1052 1570 1092 1575
rect 860 1538 888 1570
rect 888 1538 900 1570
rect 956 1538 960 1570
rect 960 1538 992 1570
rect 992 1538 996 1570
rect 1052 1538 1064 1570
rect 1064 1538 1092 1570
rect 860 1535 900 1538
rect 956 1535 996 1538
rect 1052 1535 1092 1538
rect 1312 6545 1352 6567
rect 1408 6545 1448 6567
rect 1504 6545 1544 6567
rect 1312 6527 1345 6545
rect 1345 6527 1352 6545
rect 1408 6527 1417 6545
rect 1417 6527 1448 6545
rect 1504 6527 1521 6545
rect 1521 6527 1544 6545
rect 2224 6657 2257 6663
rect 2257 6657 2264 6663
rect 2320 6657 2329 6663
rect 2329 6657 2360 6663
rect 2416 6657 2433 6663
rect 2433 6657 2456 6663
rect 2224 6623 2264 6657
rect 2320 6623 2360 6657
rect 2416 6623 2456 6657
rect 1312 6441 1345 6471
rect 1345 6441 1352 6471
rect 1408 6441 1417 6471
rect 1417 6441 1448 6471
rect 1504 6441 1521 6471
rect 1521 6441 1544 6471
rect 1312 6431 1352 6441
rect 1408 6431 1448 6441
rect 1504 6431 1544 6441
rect 1312 6369 1345 6375
rect 1345 6369 1352 6375
rect 1408 6369 1417 6375
rect 1417 6369 1448 6375
rect 1504 6369 1521 6375
rect 1521 6369 1544 6375
rect 1312 6335 1352 6369
rect 1408 6335 1448 6369
rect 1504 6335 1544 6369
rect 1312 6257 1352 6279
rect 1408 6257 1448 6279
rect 1504 6257 1544 6279
rect 1312 6239 1345 6257
rect 1345 6239 1352 6257
rect 1408 6239 1417 6257
rect 1417 6239 1448 6257
rect 1504 6239 1521 6257
rect 1521 6239 1544 6257
rect 1312 6153 1345 6183
rect 1345 6153 1352 6183
rect 1408 6153 1417 6183
rect 1417 6153 1448 6183
rect 1504 6153 1521 6183
rect 1521 6153 1544 6183
rect 1312 6143 1352 6153
rect 1408 6143 1448 6153
rect 1504 6143 1544 6153
rect 1312 4857 1345 4863
rect 1345 4857 1352 4863
rect 1408 4857 1417 4863
rect 1417 4857 1448 4863
rect 1504 4857 1521 4863
rect 1521 4857 1544 4863
rect 1312 4823 1352 4857
rect 1408 4823 1448 4857
rect 1504 4823 1544 4857
rect 1312 4745 1352 4767
rect 1408 4745 1448 4767
rect 1504 4745 1544 4767
rect 1312 4727 1345 4745
rect 1345 4727 1352 4745
rect 1408 4727 1417 4745
rect 1417 4727 1448 4745
rect 1504 4727 1521 4745
rect 1521 4727 1544 4745
rect 1312 4641 1345 4671
rect 1345 4641 1352 4671
rect 1408 4641 1417 4671
rect 1417 4641 1448 4671
rect 1504 4641 1521 4671
rect 1521 4641 1544 4671
rect 1312 4631 1352 4641
rect 1408 4631 1448 4641
rect 1504 4631 1544 4641
rect 1312 4569 1345 4575
rect 1345 4569 1352 4575
rect 1408 4569 1417 4575
rect 1417 4569 1448 4575
rect 1504 4569 1521 4575
rect 1521 4569 1544 4575
rect 1312 4535 1352 4569
rect 1408 4535 1448 4569
rect 1504 4535 1544 4569
rect 1312 4457 1352 4479
rect 1408 4457 1448 4479
rect 1504 4457 1544 4479
rect 1312 4439 1345 4457
rect 1345 4439 1352 4457
rect 1408 4439 1417 4457
rect 1417 4439 1448 4457
rect 1504 4439 1521 4457
rect 1521 4439 1544 4457
rect 1312 4353 1345 4383
rect 1345 4353 1352 4383
rect 1408 4353 1417 4383
rect 1417 4353 1448 4383
rect 1504 4353 1521 4383
rect 1521 4353 1544 4383
rect 1312 4343 1352 4353
rect 1408 4343 1448 4353
rect 1504 4343 1544 4353
rect 1312 3057 1345 3063
rect 1345 3057 1352 3063
rect 1408 3057 1417 3063
rect 1417 3057 1448 3063
rect 1504 3057 1521 3063
rect 1521 3057 1544 3063
rect 1312 3023 1352 3057
rect 1408 3023 1448 3057
rect 1504 3023 1544 3057
rect 1312 2945 1352 2967
rect 1408 2945 1448 2967
rect 1504 2945 1544 2967
rect 1312 2927 1345 2945
rect 1345 2927 1352 2945
rect 1408 2927 1417 2945
rect 1417 2927 1448 2945
rect 1504 2927 1521 2945
rect 1521 2927 1544 2945
rect 1312 2841 1345 2871
rect 1345 2841 1352 2871
rect 1408 2841 1417 2871
rect 1417 2841 1448 2871
rect 1504 2841 1521 2871
rect 1521 2841 1544 2871
rect 1312 2831 1352 2841
rect 1408 2831 1448 2841
rect 1504 2831 1544 2841
rect 1312 2769 1345 2775
rect 1345 2769 1352 2775
rect 1408 2769 1417 2775
rect 1417 2769 1448 2775
rect 1504 2769 1521 2775
rect 1521 2769 1544 2775
rect 1312 2735 1352 2769
rect 1408 2735 1448 2769
rect 1504 2735 1544 2769
rect 1312 2657 1352 2679
rect 1408 2657 1448 2679
rect 1504 2657 1544 2679
rect 1312 2639 1345 2657
rect 1345 2639 1352 2657
rect 1408 2639 1417 2657
rect 1417 2639 1448 2657
rect 1504 2639 1521 2657
rect 1521 2639 1544 2657
rect 1312 2553 1345 2583
rect 1345 2553 1352 2583
rect 1408 2553 1417 2583
rect 1417 2553 1448 2583
rect 1504 2553 1521 2583
rect 1521 2553 1544 2583
rect 1312 2543 1352 2553
rect 1408 2543 1448 2553
rect 1504 2543 1544 2553
rect 1312 1257 1345 1263
rect 1345 1257 1352 1263
rect 1408 1257 1417 1263
rect 1417 1257 1448 1263
rect 1504 1257 1521 1263
rect 1521 1257 1544 1263
rect 1312 1223 1352 1257
rect 1408 1223 1448 1257
rect 1504 1223 1544 1257
rect 1312 1145 1352 1167
rect 1408 1145 1448 1167
rect 1504 1145 1544 1167
rect 1312 1127 1345 1145
rect 1345 1127 1352 1145
rect 1408 1127 1417 1145
rect 1417 1127 1448 1145
rect 1504 1127 1521 1145
rect 1521 1127 1544 1145
rect 1312 1041 1345 1071
rect 1345 1041 1352 1071
rect 1408 1041 1417 1071
rect 1417 1041 1448 1071
rect 1504 1041 1521 1071
rect 1521 1041 1544 1071
rect 1312 1031 1352 1041
rect 1408 1031 1448 1041
rect 1504 1031 1544 1041
rect 1312 969 1345 975
rect 1345 969 1352 975
rect 1408 969 1417 975
rect 1417 969 1448 975
rect 1504 969 1521 975
rect 1521 969 1544 975
rect 1312 935 1352 969
rect 1408 935 1448 969
rect 1504 935 1544 969
rect 400 753 433 783
rect 433 753 440 783
rect 496 753 505 783
rect 505 753 536 783
rect 592 753 609 783
rect 609 753 632 783
rect 400 743 440 753
rect 496 743 536 753
rect 592 743 632 753
rect 1312 857 1352 879
rect 1408 857 1448 879
rect 1504 857 1544 879
rect 1312 839 1345 857
rect 1345 839 1352 857
rect 1408 839 1417 857
rect 1417 839 1448 857
rect 1504 839 1521 857
rect 1521 839 1544 857
rect 1766 5818 1806 5847
rect 1862 5818 1902 5847
rect 1958 5818 1998 5847
rect 1766 5807 1794 5818
rect 1794 5807 1806 5818
rect 1862 5807 1866 5818
rect 1866 5807 1898 5818
rect 1898 5807 1902 5818
rect 1958 5807 1970 5818
rect 1970 5807 1998 5818
rect 1766 5746 1806 5751
rect 1862 5746 1902 5751
rect 1958 5746 1998 5751
rect 1766 5714 1794 5746
rect 1794 5714 1806 5746
rect 1862 5714 1866 5746
rect 1866 5714 1898 5746
rect 1898 5714 1902 5746
rect 1958 5714 1970 5746
rect 1970 5714 1998 5746
rect 1766 5711 1806 5714
rect 1862 5711 1902 5714
rect 1958 5711 1998 5714
rect 1766 5642 1794 5655
rect 1794 5642 1806 5655
rect 1862 5642 1866 5655
rect 1866 5642 1898 5655
rect 1898 5642 1902 5655
rect 1958 5642 1970 5655
rect 1970 5642 1998 5655
rect 1766 5615 1806 5642
rect 1862 5615 1902 5642
rect 1958 5615 1998 5642
rect 1766 5530 1806 5559
rect 1862 5530 1902 5559
rect 1958 5530 1998 5559
rect 1766 5519 1794 5530
rect 1794 5519 1806 5530
rect 1862 5519 1866 5530
rect 1866 5519 1898 5530
rect 1898 5519 1902 5530
rect 1958 5519 1970 5530
rect 1970 5519 1998 5530
rect 1766 5458 1806 5463
rect 1862 5458 1902 5463
rect 1958 5458 1998 5463
rect 1766 5426 1794 5458
rect 1794 5426 1806 5458
rect 1862 5426 1866 5458
rect 1866 5426 1898 5458
rect 1898 5426 1902 5458
rect 1958 5426 1970 5458
rect 1970 5426 1998 5458
rect 1766 5423 1806 5426
rect 1862 5423 1902 5426
rect 1958 5423 1998 5426
rect 1766 5354 1794 5367
rect 1794 5354 1806 5367
rect 1862 5354 1866 5367
rect 1866 5354 1898 5367
rect 1898 5354 1902 5367
rect 1958 5354 1970 5367
rect 1970 5354 1998 5367
rect 1766 5327 1806 5354
rect 1862 5327 1902 5354
rect 1958 5327 1998 5354
rect 1766 5242 1806 5271
rect 1862 5242 1902 5271
rect 1958 5242 1998 5271
rect 1766 5231 1794 5242
rect 1794 5231 1806 5242
rect 1862 5231 1866 5242
rect 1866 5231 1898 5242
rect 1898 5231 1902 5242
rect 1958 5231 1970 5242
rect 1970 5231 1998 5242
rect 1766 5170 1806 5175
rect 1862 5170 1902 5175
rect 1958 5170 1998 5175
rect 1766 5138 1794 5170
rect 1794 5138 1806 5170
rect 1862 5138 1866 5170
rect 1866 5138 1898 5170
rect 1898 5138 1902 5170
rect 1958 5138 1970 5170
rect 1970 5138 1998 5170
rect 1766 5135 1806 5138
rect 1862 5135 1902 5138
rect 1958 5135 1998 5138
rect 1766 4018 1806 4047
rect 1862 4018 1902 4047
rect 1958 4018 1998 4047
rect 1766 4007 1794 4018
rect 1794 4007 1806 4018
rect 1862 4007 1866 4018
rect 1866 4007 1898 4018
rect 1898 4007 1902 4018
rect 1958 4007 1970 4018
rect 1970 4007 1998 4018
rect 1766 3946 1806 3951
rect 1862 3946 1902 3951
rect 1958 3946 1998 3951
rect 1766 3914 1794 3946
rect 1794 3914 1806 3946
rect 1862 3914 1866 3946
rect 1866 3914 1898 3946
rect 1898 3914 1902 3946
rect 1958 3914 1970 3946
rect 1970 3914 1998 3946
rect 1766 3911 1806 3914
rect 1862 3911 1902 3914
rect 1958 3911 1998 3914
rect 1766 3842 1794 3855
rect 1794 3842 1806 3855
rect 1862 3842 1866 3855
rect 1866 3842 1898 3855
rect 1898 3842 1902 3855
rect 1958 3842 1970 3855
rect 1970 3842 1998 3855
rect 1766 3815 1806 3842
rect 1862 3815 1902 3842
rect 1958 3815 1998 3842
rect 1766 3730 1806 3759
rect 1862 3730 1902 3759
rect 1958 3730 1998 3759
rect 1766 3719 1794 3730
rect 1794 3719 1806 3730
rect 1862 3719 1866 3730
rect 1866 3719 1898 3730
rect 1898 3719 1902 3730
rect 1958 3719 1970 3730
rect 1970 3719 1998 3730
rect 1766 3658 1806 3663
rect 1862 3658 1902 3663
rect 1958 3658 1998 3663
rect 1766 3626 1794 3658
rect 1794 3626 1806 3658
rect 1862 3626 1866 3658
rect 1866 3626 1898 3658
rect 1898 3626 1902 3658
rect 1958 3626 1970 3658
rect 1970 3626 1998 3658
rect 1766 3623 1806 3626
rect 1862 3623 1902 3626
rect 1958 3623 1998 3626
rect 1766 3554 1794 3567
rect 1794 3554 1806 3567
rect 1862 3554 1866 3567
rect 1866 3554 1898 3567
rect 1898 3554 1902 3567
rect 1958 3554 1970 3567
rect 1970 3554 1998 3567
rect 1766 3527 1806 3554
rect 1862 3527 1902 3554
rect 1958 3527 1998 3554
rect 1766 3442 1806 3471
rect 1862 3442 1902 3471
rect 1958 3442 1998 3471
rect 1766 3431 1794 3442
rect 1794 3431 1806 3442
rect 1862 3431 1866 3442
rect 1866 3431 1898 3442
rect 1898 3431 1902 3442
rect 1958 3431 1970 3442
rect 1970 3431 1998 3442
rect 1766 3370 1806 3375
rect 1862 3370 1902 3375
rect 1958 3370 1998 3375
rect 1766 3338 1794 3370
rect 1794 3338 1806 3370
rect 1862 3338 1866 3370
rect 1866 3338 1898 3370
rect 1898 3338 1902 3370
rect 1958 3338 1970 3370
rect 1970 3338 1998 3370
rect 1766 3335 1806 3338
rect 1862 3335 1902 3338
rect 1958 3335 1998 3338
rect 1766 2218 1806 2247
rect 1862 2218 1902 2247
rect 1958 2218 1998 2247
rect 1766 2207 1794 2218
rect 1794 2207 1806 2218
rect 1862 2207 1866 2218
rect 1866 2207 1898 2218
rect 1898 2207 1902 2218
rect 1958 2207 1970 2218
rect 1970 2207 1998 2218
rect 1766 2146 1806 2151
rect 1862 2146 1902 2151
rect 1958 2146 1998 2151
rect 1766 2114 1794 2146
rect 1794 2114 1806 2146
rect 1862 2114 1866 2146
rect 1866 2114 1898 2146
rect 1898 2114 1902 2146
rect 1958 2114 1970 2146
rect 1970 2114 1998 2146
rect 1766 2111 1806 2114
rect 1862 2111 1902 2114
rect 1958 2111 1998 2114
rect 1766 2042 1794 2055
rect 1794 2042 1806 2055
rect 1862 2042 1866 2055
rect 1866 2042 1898 2055
rect 1898 2042 1902 2055
rect 1958 2042 1970 2055
rect 1970 2042 1998 2055
rect 1766 2015 1806 2042
rect 1862 2015 1902 2042
rect 1958 2015 1998 2042
rect 1766 1930 1806 1959
rect 1862 1930 1902 1959
rect 1958 1930 1998 1959
rect 1766 1919 1794 1930
rect 1794 1919 1806 1930
rect 1862 1919 1866 1930
rect 1866 1919 1898 1930
rect 1898 1919 1902 1930
rect 1958 1919 1970 1930
rect 1970 1919 1998 1930
rect 1766 1858 1806 1863
rect 1862 1858 1902 1863
rect 1958 1858 1998 1863
rect 1766 1826 1794 1858
rect 1794 1826 1806 1858
rect 1862 1826 1866 1858
rect 1866 1826 1898 1858
rect 1898 1826 1902 1858
rect 1958 1826 1970 1858
rect 1970 1826 1998 1858
rect 1766 1823 1806 1826
rect 1862 1823 1902 1826
rect 1958 1823 1998 1826
rect 1766 1754 1794 1767
rect 1794 1754 1806 1767
rect 1862 1754 1866 1767
rect 1866 1754 1898 1767
rect 1898 1754 1902 1767
rect 1958 1754 1970 1767
rect 1970 1754 1998 1767
rect 1766 1727 1806 1754
rect 1862 1727 1902 1754
rect 1958 1727 1998 1754
rect 1766 1642 1806 1671
rect 1862 1642 1902 1671
rect 1958 1642 1998 1671
rect 1766 1631 1794 1642
rect 1794 1631 1806 1642
rect 1862 1631 1866 1642
rect 1866 1631 1898 1642
rect 1898 1631 1902 1642
rect 1958 1631 1970 1642
rect 1970 1631 1998 1642
rect 1766 1570 1806 1575
rect 1862 1570 1902 1575
rect 1958 1570 1998 1575
rect 1766 1538 1794 1570
rect 1794 1538 1806 1570
rect 1862 1538 1866 1570
rect 1866 1538 1898 1570
rect 1898 1538 1902 1570
rect 1958 1538 1970 1570
rect 1970 1538 1998 1570
rect 1766 1535 1806 1538
rect 1862 1535 1902 1538
rect 1958 1535 1998 1538
rect 2224 6545 2264 6567
rect 2320 6545 2360 6567
rect 2416 6545 2456 6567
rect 2224 6527 2257 6545
rect 2257 6527 2264 6545
rect 2320 6527 2329 6545
rect 2329 6527 2360 6545
rect 2416 6527 2433 6545
rect 2433 6527 2456 6545
rect 2224 6441 2257 6471
rect 2257 6441 2264 6471
rect 2320 6441 2329 6471
rect 2329 6441 2360 6471
rect 2416 6441 2433 6471
rect 2433 6441 2456 6471
rect 2224 6431 2264 6441
rect 2320 6431 2360 6441
rect 2416 6431 2456 6441
rect 2224 6369 2257 6375
rect 2257 6369 2264 6375
rect 2320 6369 2329 6375
rect 2329 6369 2360 6375
rect 2416 6369 2433 6375
rect 2433 6369 2456 6375
rect 2224 6335 2264 6369
rect 2320 6335 2360 6369
rect 2416 6335 2456 6369
rect 2224 6257 2264 6279
rect 2320 6257 2360 6279
rect 2416 6257 2456 6279
rect 2224 6239 2257 6257
rect 2257 6239 2264 6257
rect 2320 6239 2329 6257
rect 2329 6239 2360 6257
rect 2416 6239 2433 6257
rect 2433 6239 2456 6257
rect 2224 6153 2257 6183
rect 2257 6153 2264 6183
rect 2320 6153 2329 6183
rect 2329 6153 2360 6183
rect 2416 6153 2433 6183
rect 2433 6153 2456 6183
rect 2224 6143 2264 6153
rect 2320 6143 2360 6153
rect 2416 6143 2456 6153
rect 2224 4857 2257 4863
rect 2257 4857 2264 4863
rect 2320 4857 2329 4863
rect 2329 4857 2360 4863
rect 2416 4857 2433 4863
rect 2433 4857 2456 4863
rect 2224 4823 2264 4857
rect 2320 4823 2360 4857
rect 2416 4823 2456 4857
rect 2224 4745 2264 4767
rect 2320 4745 2360 4767
rect 2416 4745 2456 4767
rect 2224 4727 2257 4745
rect 2257 4727 2264 4745
rect 2320 4727 2329 4745
rect 2329 4727 2360 4745
rect 2416 4727 2433 4745
rect 2433 4727 2456 4745
rect 2224 4641 2257 4671
rect 2257 4641 2264 4671
rect 2320 4641 2329 4671
rect 2329 4641 2360 4671
rect 2416 4641 2433 4671
rect 2433 4641 2456 4671
rect 2224 4631 2264 4641
rect 2320 4631 2360 4641
rect 2416 4631 2456 4641
rect 2224 4569 2257 4575
rect 2257 4569 2264 4575
rect 2320 4569 2329 4575
rect 2329 4569 2360 4575
rect 2416 4569 2433 4575
rect 2433 4569 2456 4575
rect 2224 4535 2264 4569
rect 2320 4535 2360 4569
rect 2416 4535 2456 4569
rect 2224 4457 2264 4479
rect 2320 4457 2360 4479
rect 2416 4457 2456 4479
rect 2224 4439 2257 4457
rect 2257 4439 2264 4457
rect 2320 4439 2329 4457
rect 2329 4439 2360 4457
rect 2416 4439 2433 4457
rect 2433 4439 2456 4457
rect 2224 4353 2257 4383
rect 2257 4353 2264 4383
rect 2320 4353 2329 4383
rect 2329 4353 2360 4383
rect 2416 4353 2433 4383
rect 2433 4353 2456 4383
rect 2224 4343 2264 4353
rect 2320 4343 2360 4353
rect 2416 4343 2456 4353
rect 2224 3057 2257 3063
rect 2257 3057 2264 3063
rect 2320 3057 2329 3063
rect 2329 3057 2360 3063
rect 2416 3057 2433 3063
rect 2433 3057 2456 3063
rect 2224 3023 2264 3057
rect 2320 3023 2360 3057
rect 2416 3023 2456 3057
rect 2224 2945 2264 2967
rect 2320 2945 2360 2967
rect 2416 2945 2456 2967
rect 2224 2927 2257 2945
rect 2257 2927 2264 2945
rect 2320 2927 2329 2945
rect 2329 2927 2360 2945
rect 2416 2927 2433 2945
rect 2433 2927 2456 2945
rect 2224 2841 2257 2871
rect 2257 2841 2264 2871
rect 2320 2841 2329 2871
rect 2329 2841 2360 2871
rect 2416 2841 2433 2871
rect 2433 2841 2456 2871
rect 2224 2831 2264 2841
rect 2320 2831 2360 2841
rect 2416 2831 2456 2841
rect 2224 2769 2257 2775
rect 2257 2769 2264 2775
rect 2320 2769 2329 2775
rect 2329 2769 2360 2775
rect 2416 2769 2433 2775
rect 2433 2769 2456 2775
rect 2224 2735 2264 2769
rect 2320 2735 2360 2769
rect 2416 2735 2456 2769
rect 2224 2657 2264 2679
rect 2320 2657 2360 2679
rect 2416 2657 2456 2679
rect 2224 2639 2257 2657
rect 2257 2639 2264 2657
rect 2320 2639 2329 2657
rect 2329 2639 2360 2657
rect 2416 2639 2433 2657
rect 2433 2639 2456 2657
rect 2224 2553 2257 2583
rect 2257 2553 2264 2583
rect 2320 2553 2329 2583
rect 2329 2553 2360 2583
rect 2416 2553 2433 2583
rect 2433 2553 2456 2583
rect 2224 2543 2264 2553
rect 2320 2543 2360 2553
rect 2416 2543 2456 2553
rect 2224 1257 2257 1263
rect 2257 1257 2264 1263
rect 2320 1257 2329 1263
rect 2329 1257 2360 1263
rect 2416 1257 2433 1263
rect 2433 1257 2456 1263
rect 2224 1223 2264 1257
rect 2320 1223 2360 1257
rect 2416 1223 2456 1257
rect 2224 1145 2264 1167
rect 2320 1145 2360 1167
rect 2416 1145 2456 1167
rect 2224 1127 2257 1145
rect 2257 1127 2264 1145
rect 2320 1127 2329 1145
rect 2329 1127 2360 1145
rect 2416 1127 2433 1145
rect 2433 1127 2456 1145
rect 2224 1041 2257 1071
rect 2257 1041 2264 1071
rect 2320 1041 2329 1071
rect 2329 1041 2360 1071
rect 2416 1041 2433 1071
rect 2433 1041 2456 1071
rect 2224 1031 2264 1041
rect 2320 1031 2360 1041
rect 2416 1031 2456 1041
rect 2224 969 2257 975
rect 2257 969 2264 975
rect 2320 969 2329 975
rect 2329 969 2360 975
rect 2416 969 2433 975
rect 2433 969 2456 975
rect 2224 935 2264 969
rect 2320 935 2360 969
rect 2416 935 2456 969
rect 1312 753 1345 783
rect 1345 753 1352 783
rect 1408 753 1417 783
rect 1417 753 1448 783
rect 1504 753 1521 783
rect 1521 753 1544 783
rect 1312 743 1352 753
rect 1408 743 1448 753
rect 1504 743 1544 753
rect 2224 857 2264 879
rect 2320 857 2360 879
rect 2416 857 2456 879
rect 2224 839 2257 857
rect 2257 839 2264 857
rect 2320 839 2329 857
rect 2329 839 2360 857
rect 2416 839 2433 857
rect 2433 839 2456 857
rect 2224 753 2257 783
rect 2257 753 2264 783
rect 2320 753 2329 783
rect 2329 753 2360 783
rect 2416 753 2433 783
rect 2433 753 2456 783
rect 2224 743 2264 753
rect 2320 743 2360 753
rect 2416 743 2456 753
<< metal2 >>
rect 391 6623 400 6663
rect 440 6623 496 6663
rect 536 6623 592 6663
rect 632 6623 1312 6663
rect 1352 6623 1408 6663
rect 1448 6623 1504 6663
rect 1544 6623 2224 6663
rect 2264 6623 2320 6663
rect 2360 6623 2416 6663
rect 2456 6623 3101 6663
rect 391 6567 3101 6623
rect 391 6527 400 6567
rect 440 6527 496 6567
rect 536 6527 592 6567
rect 632 6527 1312 6567
rect 1352 6527 1408 6567
rect 1448 6527 1504 6567
rect 1544 6527 2224 6567
rect 2264 6527 2320 6567
rect 2360 6527 2416 6567
rect 2456 6527 3101 6567
rect 391 6471 3101 6527
rect 391 6431 400 6471
rect 440 6431 496 6471
rect 536 6431 592 6471
rect 632 6431 1312 6471
rect 1352 6431 1408 6471
rect 1448 6431 1504 6471
rect 1544 6431 2224 6471
rect 2264 6431 2320 6471
rect 2360 6431 2416 6471
rect 2456 6431 3101 6471
rect 391 6375 3101 6431
rect 391 6335 400 6375
rect 440 6335 496 6375
rect 536 6335 592 6375
rect 632 6335 1312 6375
rect 1352 6335 1408 6375
rect 1448 6335 1504 6375
rect 1544 6335 2224 6375
rect 2264 6335 2320 6375
rect 2360 6335 2416 6375
rect 2456 6335 3101 6375
rect 391 6279 3101 6335
rect 391 6239 400 6279
rect 440 6239 496 6279
rect 536 6239 592 6279
rect 632 6239 1312 6279
rect 1352 6239 1408 6279
rect 1448 6239 1504 6279
rect 1544 6239 2224 6279
rect 2264 6239 2320 6279
rect 2360 6239 2416 6279
rect 2456 6239 3101 6279
rect 391 6183 3101 6239
rect 391 6143 400 6183
rect 440 6143 496 6183
rect 536 6143 592 6183
rect 632 6143 1312 6183
rect 1352 6143 1408 6183
rect 1448 6143 1504 6183
rect 1544 6143 2224 6183
rect 2264 6143 2320 6183
rect 2360 6143 2416 6183
rect 2456 6143 3101 6183
rect -460 5847 1908 5859
rect -460 5807 860 5847
rect 900 5807 956 5847
rect 996 5807 1052 5847
rect 1092 5807 1766 5847
rect 1806 5807 1862 5847
rect 1902 5807 1958 5847
rect 1998 5807 2007 5847
rect -460 5751 2007 5807
rect -460 5711 860 5751
rect 900 5711 956 5751
rect 996 5711 1052 5751
rect 1092 5711 1766 5751
rect 1806 5711 1862 5751
rect 1902 5711 1958 5751
rect 1998 5711 2007 5751
rect -460 5655 2007 5711
rect -460 5615 860 5655
rect 900 5615 956 5655
rect 996 5615 1052 5655
rect 1092 5615 1766 5655
rect 1806 5615 1862 5655
rect 1902 5615 1958 5655
rect 1998 5615 2007 5655
rect -460 5559 2007 5615
rect -460 5519 860 5559
rect 900 5519 956 5559
rect 996 5519 1052 5559
rect 1092 5519 1766 5559
rect 1806 5519 1862 5559
rect 1902 5519 1958 5559
rect 1998 5519 2007 5559
rect -460 5463 2007 5519
rect -460 5423 860 5463
rect 900 5423 956 5463
rect 996 5423 1052 5463
rect 1092 5423 1766 5463
rect 1806 5423 1862 5463
rect 1902 5423 1958 5463
rect 1998 5423 2007 5463
rect -460 5367 2007 5423
rect -460 5327 860 5367
rect 900 5327 956 5367
rect 996 5327 1052 5367
rect 1092 5327 1766 5367
rect 1806 5327 1862 5367
rect 1902 5327 1958 5367
rect 1998 5327 2007 5367
rect -460 5271 2007 5327
rect -460 5231 860 5271
rect 900 5231 956 5271
rect 996 5231 1052 5271
rect 1092 5231 1766 5271
rect 1806 5231 1862 5271
rect 1902 5231 1958 5271
rect 1998 5231 2007 5271
rect -460 5175 2007 5231
rect -460 5147 860 5175
rect -460 4059 261 5147
rect 851 5135 860 5147
rect 900 5135 956 5175
rect 996 5135 1052 5175
rect 1092 5147 1766 5175
rect 1092 5135 1101 5147
rect 1757 5135 1766 5147
rect 1806 5135 1862 5175
rect 1902 5135 1958 5175
rect 1998 5135 2007 5175
rect 2372 4863 3101 6143
rect 391 4823 400 4863
rect 440 4823 496 4863
rect 536 4823 592 4863
rect 632 4823 1312 4863
rect 1352 4823 1408 4863
rect 1448 4823 1504 4863
rect 1544 4823 2224 4863
rect 2264 4823 2320 4863
rect 2360 4823 2416 4863
rect 2456 4823 3101 4863
rect 391 4767 3101 4823
rect 391 4727 400 4767
rect 440 4727 496 4767
rect 536 4727 592 4767
rect 632 4727 1312 4767
rect 1352 4727 1408 4767
rect 1448 4727 1504 4767
rect 1544 4727 2224 4767
rect 2264 4727 2320 4767
rect 2360 4727 2416 4767
rect 2456 4727 3101 4767
rect 391 4671 3101 4727
rect 391 4631 400 4671
rect 440 4631 496 4671
rect 536 4631 592 4671
rect 632 4631 1312 4671
rect 1352 4631 1408 4671
rect 1448 4631 1504 4671
rect 1544 4631 2224 4671
rect 2264 4631 2320 4671
rect 2360 4631 2416 4671
rect 2456 4631 3101 4671
rect 391 4575 3101 4631
rect 391 4535 400 4575
rect 440 4535 496 4575
rect 536 4535 592 4575
rect 632 4535 1312 4575
rect 1352 4535 1408 4575
rect 1448 4535 1504 4575
rect 1544 4535 2224 4575
rect 2264 4535 2320 4575
rect 2360 4535 2416 4575
rect 2456 4535 3101 4575
rect 391 4479 3101 4535
rect 391 4439 400 4479
rect 440 4439 496 4479
rect 536 4439 592 4479
rect 632 4439 1312 4479
rect 1352 4439 1408 4479
rect 1448 4439 1504 4479
rect 1544 4439 2224 4479
rect 2264 4439 2320 4479
rect 2360 4439 2416 4479
rect 2456 4439 3101 4479
rect 391 4383 3101 4439
rect 391 4343 400 4383
rect 440 4343 496 4383
rect 536 4343 592 4383
rect 632 4343 1312 4383
rect 1352 4343 1408 4383
rect 1448 4343 1504 4383
rect 1544 4343 2224 4383
rect 2264 4343 2320 4383
rect 2360 4343 2416 4383
rect 2456 4343 3101 4383
rect -460 4047 1908 4059
rect -460 4007 860 4047
rect 900 4007 956 4047
rect 996 4007 1052 4047
rect 1092 4007 1766 4047
rect 1806 4007 1862 4047
rect 1902 4007 1958 4047
rect 1998 4007 2007 4047
rect -460 3951 2007 4007
rect -460 3911 860 3951
rect 900 3911 956 3951
rect 996 3911 1052 3951
rect 1092 3911 1766 3951
rect 1806 3911 1862 3951
rect 1902 3911 1958 3951
rect 1998 3911 2007 3951
rect -460 3855 2007 3911
rect -460 3815 860 3855
rect 900 3815 956 3855
rect 996 3815 1052 3855
rect 1092 3815 1766 3855
rect 1806 3815 1862 3855
rect 1902 3815 1958 3855
rect 1998 3815 2007 3855
rect -460 3759 2007 3815
rect -460 3719 860 3759
rect 900 3719 956 3759
rect 996 3719 1052 3759
rect 1092 3719 1766 3759
rect 1806 3719 1862 3759
rect 1902 3719 1958 3759
rect 1998 3719 2007 3759
rect -460 3663 2007 3719
rect -460 3623 860 3663
rect 900 3623 956 3663
rect 996 3623 1052 3663
rect 1092 3623 1766 3663
rect 1806 3623 1862 3663
rect 1902 3623 1958 3663
rect 1998 3623 2007 3663
rect -460 3567 2007 3623
rect -460 3527 860 3567
rect 900 3527 956 3567
rect 996 3527 1052 3567
rect 1092 3527 1766 3567
rect 1806 3527 1862 3567
rect 1902 3527 1958 3567
rect 1998 3527 2007 3567
rect -460 3471 2007 3527
rect -460 3431 860 3471
rect 900 3431 956 3471
rect 996 3431 1052 3471
rect 1092 3431 1766 3471
rect 1806 3431 1862 3471
rect 1902 3431 1958 3471
rect 1998 3431 2007 3471
rect -460 3375 2007 3431
rect -460 3347 860 3375
rect -460 2259 261 3347
rect 851 3335 860 3347
rect 900 3335 956 3375
rect 996 3335 1052 3375
rect 1092 3347 1766 3375
rect 1092 3335 1101 3347
rect 1757 3335 1766 3347
rect 1806 3335 1862 3375
rect 1902 3335 1958 3375
rect 1998 3335 2007 3375
rect 2372 3063 3101 4343
rect 391 3023 400 3063
rect 440 3023 496 3063
rect 536 3023 592 3063
rect 632 3023 1312 3063
rect 1352 3023 1408 3063
rect 1448 3023 1504 3063
rect 1544 3023 2224 3063
rect 2264 3023 2320 3063
rect 2360 3023 2416 3063
rect 2456 3023 3101 3063
rect 391 2967 3101 3023
rect 391 2927 400 2967
rect 440 2927 496 2967
rect 536 2927 592 2967
rect 632 2927 1312 2967
rect 1352 2927 1408 2967
rect 1448 2927 1504 2967
rect 1544 2927 2224 2967
rect 2264 2927 2320 2967
rect 2360 2927 2416 2967
rect 2456 2927 3101 2967
rect 391 2871 3101 2927
rect 391 2831 400 2871
rect 440 2831 496 2871
rect 536 2831 592 2871
rect 632 2831 1312 2871
rect 1352 2831 1408 2871
rect 1448 2831 1504 2871
rect 1544 2831 2224 2871
rect 2264 2831 2320 2871
rect 2360 2831 2416 2871
rect 2456 2831 3101 2871
rect 391 2775 3101 2831
rect 391 2735 400 2775
rect 440 2735 496 2775
rect 536 2735 592 2775
rect 632 2735 1312 2775
rect 1352 2735 1408 2775
rect 1448 2735 1504 2775
rect 1544 2735 2224 2775
rect 2264 2735 2320 2775
rect 2360 2735 2416 2775
rect 2456 2735 3101 2775
rect 391 2679 3101 2735
rect 391 2639 400 2679
rect 440 2639 496 2679
rect 536 2639 592 2679
rect 632 2639 1312 2679
rect 1352 2639 1408 2679
rect 1448 2639 1504 2679
rect 1544 2639 2224 2679
rect 2264 2639 2320 2679
rect 2360 2639 2416 2679
rect 2456 2639 3101 2679
rect 391 2583 3101 2639
rect 391 2543 400 2583
rect 440 2543 496 2583
rect 536 2543 592 2583
rect 632 2543 1312 2583
rect 1352 2543 1408 2583
rect 1448 2543 1504 2583
rect 1544 2543 2224 2583
rect 2264 2543 2320 2583
rect 2360 2543 2416 2583
rect 2456 2543 3101 2583
rect -460 2247 1908 2259
rect -460 2207 860 2247
rect 900 2207 956 2247
rect 996 2207 1052 2247
rect 1092 2207 1766 2247
rect 1806 2207 1862 2247
rect 1902 2207 1958 2247
rect 1998 2207 2007 2247
rect -460 2151 2007 2207
rect -460 2111 860 2151
rect 900 2111 956 2151
rect 996 2111 1052 2151
rect 1092 2111 1766 2151
rect 1806 2111 1862 2151
rect 1902 2111 1958 2151
rect 1998 2111 2007 2151
rect -460 2055 2007 2111
rect -460 2015 860 2055
rect 900 2015 956 2055
rect 996 2015 1052 2055
rect 1092 2015 1766 2055
rect 1806 2015 1862 2055
rect 1902 2015 1958 2055
rect 1998 2015 2007 2055
rect -460 1959 2007 2015
rect -460 1919 860 1959
rect 900 1919 956 1959
rect 996 1919 1052 1959
rect 1092 1919 1766 1959
rect 1806 1919 1862 1959
rect 1902 1919 1958 1959
rect 1998 1919 2007 1959
rect -460 1863 2007 1919
rect -460 1823 860 1863
rect 900 1823 956 1863
rect 996 1823 1052 1863
rect 1092 1823 1766 1863
rect 1806 1823 1862 1863
rect 1902 1823 1958 1863
rect 1998 1823 2007 1863
rect -460 1767 2007 1823
rect -460 1727 860 1767
rect 900 1727 956 1767
rect 996 1727 1052 1767
rect 1092 1727 1766 1767
rect 1806 1727 1862 1767
rect 1902 1727 1958 1767
rect 1998 1727 2007 1767
rect -460 1671 2007 1727
rect -460 1631 860 1671
rect 900 1631 956 1671
rect 996 1631 1052 1671
rect 1092 1631 1766 1671
rect 1806 1631 1862 1671
rect 1902 1631 1958 1671
rect 1998 1631 2007 1671
rect -460 1575 2007 1631
rect -460 1547 860 1575
rect 851 1535 860 1547
rect 900 1535 956 1575
rect 996 1535 1052 1575
rect 1092 1547 1766 1575
rect 1092 1535 1101 1547
rect 1757 1535 1766 1547
rect 1806 1535 1862 1575
rect 1902 1535 1958 1575
rect 1998 1535 2007 1575
rect 2372 1263 3101 2543
rect 391 1223 400 1263
rect 440 1223 496 1263
rect 536 1223 592 1263
rect 632 1223 1312 1263
rect 1352 1223 1408 1263
rect 1448 1223 1504 1263
rect 1544 1223 2224 1263
rect 2264 1223 2320 1263
rect 2360 1223 2416 1263
rect 2456 1223 3101 1263
rect 391 1167 3101 1223
rect 391 1127 400 1167
rect 440 1127 496 1167
rect 536 1127 592 1167
rect 632 1127 1312 1167
rect 1352 1127 1408 1167
rect 1448 1127 1504 1167
rect 1544 1127 2224 1167
rect 2264 1127 2320 1167
rect 2360 1127 2416 1167
rect 2456 1127 3101 1167
rect 391 1071 3101 1127
rect 391 1031 400 1071
rect 440 1031 496 1071
rect 536 1031 592 1071
rect 632 1031 1312 1071
rect 1352 1031 1408 1071
rect 1448 1031 1504 1071
rect 1544 1031 2224 1071
rect 2264 1031 2320 1071
rect 2360 1031 2416 1071
rect 2456 1031 3101 1071
rect 391 975 3101 1031
rect 391 935 400 975
rect 440 935 496 975
rect 536 935 592 975
rect 632 935 1312 975
rect 1352 935 1408 975
rect 1448 935 1504 975
rect 1544 935 2224 975
rect 2264 935 2320 975
rect 2360 935 2416 975
rect 2456 935 3101 975
rect 391 879 3101 935
rect 391 839 400 879
rect 440 839 496 879
rect 536 839 592 879
rect 632 839 1312 879
rect 1352 839 1408 879
rect 1448 839 1504 879
rect 1544 839 2224 879
rect 2264 839 2320 879
rect 2360 839 2416 879
rect 2456 839 3101 879
rect 391 783 3101 839
rect 391 743 400 783
rect 440 743 496 783
rect 536 743 592 783
rect 632 743 1312 783
rect 1352 743 1408 783
rect 1448 743 1504 783
rect 1544 743 2224 783
rect 2264 743 2320 783
rect 2360 743 2416 783
rect 2456 743 3101 783
<< labels >>
flabel comment s -102 3688 -102 3688 0 FreeSans 400 0 0 0 PAD
flabel comment s 2728 3705 2728 3705 0 FreeSans 400 0 0 0 VDD
flabel comment s 1432 7275 1432 7275 0 FreeSans 400 0 0 0 VSS
flabel comment s 689 99 689 99 0 FreeSans 400 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 131812
string GDS_FILE diodevdd_4kv.gds
string GDS_START 272
<< end >>
