magic
tech ihp-sg13g2
timestamp 1749416725
<< error_p >>
rect -93 530 -88 535
rect 88 530 93 535
rect 225 530 230 535
rect 406 530 411 535
rect -98 525 -93 530
rect 93 525 98 530
rect 220 525 225 530
rect 411 525 416 530
rect -98 514 -93 519
rect 93 514 98 519
rect 220 514 225 519
rect 411 514 416 519
rect -93 509 -88 514
rect 88 509 93 514
rect 225 509 230 514
rect 406 509 411 514
rect -127 493 -122 498
rect -116 493 -111 498
rect 111 493 116 498
rect 122 493 127 498
rect 191 493 196 498
rect 202 493 207 498
rect 429 493 434 498
rect 440 493 445 498
rect -132 488 -127 493
rect -111 488 -106 493
rect 106 488 111 493
rect 127 488 132 493
rect 186 488 191 493
rect 207 488 212 493
rect 424 488 429 493
rect 445 488 450 493
rect -132 -493 -127 -488
rect -111 -493 -106 -488
rect 106 -493 111 -488
rect 127 -493 132 -488
rect 186 -493 191 -488
rect 207 -493 212 -488
rect 424 -493 429 -488
rect 445 -493 450 -488
rect -127 -498 -122 -493
rect -116 -498 -111 -493
rect 111 -498 116 -493
rect 122 -498 127 -493
rect 191 -498 196 -493
rect 202 -498 207 -493
rect 429 -498 434 -493
rect 440 -498 445 -493
rect -93 -514 -88 -509
rect 88 -514 93 -509
rect 225 -514 230 -509
rect 406 -514 411 -509
rect -98 -519 -93 -514
rect 93 -519 98 -514
rect 220 -519 225 -514
rect 411 -519 416 -514
rect -98 -530 -93 -525
rect 93 -530 98 -525
rect 220 -530 225 -525
rect 411 -530 416 -525
rect -93 -535 -88 -530
rect 88 -535 93 -530
rect 225 -535 230 -530
rect 406 -535 411 -530
<< nwell >>
rect -280 -651 598 651
<< hvpmos >>
rect -100 -500 100 500
rect 218 -500 418 500
<< hvpdiff >>
rect -134 493 -100 500
rect -134 -493 -127 493
rect -111 -493 -100 493
rect -134 -500 -100 -493
rect 100 493 134 500
rect 100 -493 111 493
rect 127 -493 134 493
rect 100 -500 134 -493
rect 184 493 218 500
rect 184 -493 191 493
rect 207 -493 218 493
rect 184 -500 218 -493
rect 418 493 452 500
rect 418 -493 429 493
rect 445 -493 452 493
rect 418 -500 452 -493
<< hvpdiffc >>
rect -127 -493 -111 493
rect 111 -493 127 493
rect 191 -493 207 493
rect 429 -493 445 493
<< nsubdiff >>
rect -218 582 536 589
rect -218 566 -181 582
rect 499 566 536 582
rect -218 559 536 566
rect -218 552 -188 559
rect -218 -552 -211 552
rect -195 -552 -188 552
rect 506 552 536 559
rect -218 -559 -188 -552
rect 506 -552 513 552
rect 529 -552 536 552
rect 506 -559 536 -552
rect -218 -566 536 -559
rect -218 -582 -181 -566
rect 499 -582 536 -566
rect -218 -589 536 -582
<< nsubdiffcont >>
rect -181 566 499 582
rect -211 -552 -195 552
rect 513 -552 529 552
rect -181 -582 499 -566
<< poly >>
rect -100 530 100 537
rect -100 514 -93 530
rect 93 514 100 530
rect -100 500 100 514
rect 218 530 418 537
rect 218 514 225 530
rect 411 514 418 530
rect 218 500 418 514
rect -100 -514 100 -500
rect -100 -530 -93 -514
rect 93 -530 100 -514
rect -100 -537 100 -530
rect 218 -514 418 -500
rect 218 -530 225 -514
rect 411 -530 418 -514
rect 218 -537 418 -530
<< polycont >>
rect -93 514 93 530
rect 225 514 411 530
rect -93 -530 93 -514
rect 225 -530 411 -514
<< metal1 >>
rect -216 582 534 587
rect -216 566 -181 582
rect 499 566 534 582
rect -216 561 534 566
rect -216 552 -190 561
rect -216 -552 -211 552
rect -195 -552 -190 552
rect 508 552 534 561
rect -216 -561 -190 -552
rect 508 -552 513 552
rect 529 -552 534 552
rect 508 -561 534 -552
rect -216 -566 534 -561
rect -216 -582 -181 -566
rect 499 -582 534 -566
rect -216 -587 534 -582
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 10 l 2 nf 1 nx 2 dx 0.5 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
