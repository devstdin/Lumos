magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 14 56 348 288
rect -26 -56 410 56
<< nmos >>
rect 108 152 134 262
rect 218 114 244 262
<< pmos >>
rect 108 468 134 636
rect 218 412 244 636
<< ndiff >>
rect 40 247 108 262
rect 40 215 54 247
rect 86 215 108 247
rect 40 152 108 215
rect 134 202 218 262
rect 134 170 164 202
rect 196 170 218 202
rect 134 152 218 170
rect 148 114 218 152
rect 244 245 322 262
rect 244 213 276 245
rect 308 213 322 245
rect 244 162 322 213
rect 244 130 276 162
rect 308 130 322 162
rect 244 114 322 130
<< pdiff >>
rect 40 622 108 636
rect 40 590 54 622
rect 86 590 108 622
rect 40 554 108 590
rect 40 522 54 554
rect 86 522 108 554
rect 40 468 108 522
rect 134 622 218 636
rect 134 590 164 622
rect 196 590 218 622
rect 134 468 218 590
rect 168 412 218 468
rect 244 622 319 636
rect 244 590 273 622
rect 305 590 319 622
rect 244 554 319 590
rect 244 522 273 554
rect 305 522 319 554
rect 244 486 319 522
rect 244 454 273 486
rect 305 454 319 486
rect 244 412 319 454
<< ndiffc >>
rect 54 215 86 247
rect 164 170 196 202
rect 276 213 308 245
rect 276 130 308 162
<< pdiffc >>
rect 54 590 86 622
rect 54 522 86 554
rect 164 590 196 622
rect 273 590 305 622
rect 273 522 305 554
rect 273 454 305 486
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 108 636 134 672
rect 218 636 244 672
rect 108 446 134 468
rect 73 432 134 446
rect 73 400 87 432
rect 119 400 134 432
rect 73 386 134 400
rect 108 262 134 386
rect 218 366 244 412
rect 184 349 244 366
rect 184 317 198 349
rect 230 317 244 349
rect 184 300 244 317
rect 218 262 244 300
rect 108 116 134 152
rect 218 78 244 114
<< polycont >>
rect 87 400 119 432
rect 198 317 230 349
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 48 622 102 636
rect 48 590 54 622
rect 86 590 102 622
rect 48 554 102 590
rect 154 622 206 712
rect 154 590 164 622
rect 196 590 206 622
rect 154 578 206 590
rect 260 622 320 636
rect 260 590 273 622
rect 305 590 320 622
rect 48 522 54 554
rect 86 524 102 554
rect 260 554 320 590
rect 86 522 214 524
rect 48 488 214 522
rect 57 432 136 452
rect 57 400 87 432
rect 119 400 136 432
rect 57 386 136 400
rect 180 366 214 488
rect 260 522 273 554
rect 305 522 320 554
rect 260 486 320 522
rect 260 454 273 486
rect 305 454 320 486
rect 260 404 320 454
rect 180 349 245 366
rect 180 317 198 349
rect 230 317 245 349
rect 180 300 245 317
rect 180 293 214 300
rect 43 258 214 293
rect 282 258 320 404
rect 43 247 103 258
rect 43 215 54 247
rect 86 215 103 247
rect 43 200 103 215
rect 262 245 320 258
rect 153 202 203 214
rect 153 170 164 202
rect 196 170 203 202
rect 153 44 203 170
rect 262 213 276 245
rect 308 213 320 245
rect 262 162 320 213
rect 262 130 276 162
rect 308 130 320 162
rect 262 110 320 130
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 263 414 316 589 0 FreeSans 340 0 0 0 X
port 2 nsew
flabel metal1 s 57 386 136 452 0 FreeSans 340 0 0 0 A
port 3 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 111510
string GDS_FILE 6_final.gds
string GDS_START 108382
<< end >>
