magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 443 2736 834
rect -48 370 454 443
rect -48 350 187 370
rect 1044 367 2736 443
rect 1044 348 1463 367
rect 2019 350 2736 367
rect 2019 330 2514 350
<< pwell >>
rect 755 382 855 384
rect 669 358 998 382
rect 223 237 426 333
rect 647 309 998 358
rect 647 301 1435 309
rect 647 246 1790 301
rect 2356 268 2673 288
rect 647 237 715 246
rect 223 224 715 237
rect 12 56 715 224
rect 1001 224 1790 246
rect 2150 224 2673 268
rect 1001 56 2673 224
rect -26 -56 2714 56
<< nmos >>
rect 106 114 132 198
rect 190 114 216 198
rect 306 159 332 307
rect 741 272 767 356
rect 843 272 869 356
rect 524 127 550 211
rect 587 127 613 211
rect 1095 135 1121 283
rect 1315 135 1341 283
rect 1557 191 1583 275
rect 1664 127 1690 275
rect 1874 114 1900 198
rect 1976 114 2002 198
rect 2038 114 2064 198
rect 2244 114 2270 242
rect 2450 114 2476 262
rect 2553 114 2579 262
<< pmos >>
rect 106 432 132 516
rect 208 432 234 516
rect 298 432 324 632
rect 508 505 534 589
rect 655 505 681 589
rect 733 505 759 589
rect 835 505 861 589
rect 1175 410 1201 634
rect 1320 410 1346 634
rect 1607 429 1633 629
rect 1746 429 1772 513
rect 1822 429 1848 513
rect 1944 429 1970 513
rect 2046 429 2072 513
rect 2160 429 2186 629
rect 2450 412 2476 636
rect 2553 412 2579 636
<< ndiff >>
rect 249 198 306 307
rect 38 167 106 198
rect 38 135 52 167
rect 84 135 106 167
rect 38 114 106 135
rect 132 114 190 198
rect 216 167 306 198
rect 216 135 238 167
rect 270 159 306 167
rect 332 208 400 307
rect 781 356 829 358
rect 695 332 741 356
rect 673 318 741 332
rect 673 286 687 318
rect 719 286 741 318
rect 673 272 741 286
rect 767 344 843 356
rect 767 312 789 344
rect 821 312 843 344
rect 767 272 843 312
rect 869 330 972 356
rect 869 298 926 330
rect 958 298 972 330
rect 869 272 972 298
rect 332 176 354 208
rect 386 176 400 208
rect 332 159 400 176
rect 443 173 524 211
rect 270 135 289 159
rect 216 114 289 135
rect 443 141 457 173
rect 489 141 524 173
rect 443 127 524 141
rect 550 127 587 211
rect 613 191 689 211
rect 613 159 643 191
rect 675 159 689 191
rect 613 127 689 159
rect 1027 269 1095 283
rect 1027 237 1041 269
rect 1073 237 1095 269
rect 1027 135 1095 237
rect 1121 135 1315 283
rect 1341 204 1409 283
rect 1341 172 1363 204
rect 1395 172 1409 204
rect 1489 247 1557 275
rect 1489 215 1503 247
rect 1535 215 1557 247
rect 1489 191 1557 215
rect 1583 261 1664 275
rect 1583 229 1605 261
rect 1637 229 1664 261
rect 1583 191 1664 229
rect 1341 135 1409 172
rect 1136 36 1196 135
rect 1612 127 1664 191
rect 1690 127 1764 275
rect 2176 228 2244 242
rect 1704 124 1764 127
rect 1704 92 1718 124
rect 1750 92 1764 124
rect 1806 167 1874 198
rect 1806 135 1820 167
rect 1852 135 1874 167
rect 1806 114 1874 135
rect 1900 167 1976 198
rect 1900 135 1922 167
rect 1954 135 1976 167
rect 1900 114 1976 135
rect 2002 114 2038 198
rect 2064 167 2132 198
rect 2064 135 2086 167
rect 2118 135 2132 167
rect 2064 114 2132 135
rect 2176 196 2190 228
rect 2222 196 2244 228
rect 2176 160 2244 196
rect 2176 128 2190 160
rect 2222 128 2244 160
rect 2176 114 2244 128
rect 2270 228 2338 242
rect 2270 196 2292 228
rect 2324 196 2338 228
rect 2270 160 2338 196
rect 2270 128 2292 160
rect 2324 128 2338 160
rect 2270 114 2338 128
rect 2382 228 2450 262
rect 2382 196 2396 228
rect 2428 196 2450 228
rect 2382 160 2450 196
rect 2382 128 2396 160
rect 2428 128 2450 160
rect 2382 114 2450 128
rect 2476 228 2553 262
rect 2476 196 2498 228
rect 2530 196 2553 228
rect 2476 160 2553 196
rect 2476 128 2498 160
rect 2530 128 2553 160
rect 2476 114 2553 128
rect 2579 228 2647 262
rect 2579 196 2601 228
rect 2633 196 2647 228
rect 2579 160 2647 196
rect 2579 128 2601 160
rect 2633 128 2647 160
rect 2579 114 2647 128
rect 1704 78 1764 92
<< pdiff >>
rect 38 665 283 679
rect 38 633 53 665
rect 85 633 283 665
rect 38 632 283 633
rect 38 602 298 632
rect 248 516 298 602
rect 38 490 106 516
rect 38 458 52 490
rect 84 458 106 490
rect 38 432 106 458
rect 132 491 208 516
rect 132 459 154 491
rect 186 459 208 491
rect 132 432 208 459
rect 234 432 298 516
rect 324 570 392 632
rect 576 614 636 628
rect 576 589 590 614
rect 324 538 346 570
rect 378 538 392 570
rect 324 432 392 538
rect 438 570 508 589
rect 438 538 452 570
rect 484 538 508 570
rect 438 505 508 538
rect 534 582 590 589
rect 622 589 636 614
rect 1215 634 1306 720
rect 622 582 655 589
rect 534 505 655 582
rect 681 505 733 589
rect 759 551 835 589
rect 759 519 781 551
rect 813 519 835 551
rect 759 505 835 519
rect 861 573 929 589
rect 861 541 883 573
rect 915 541 929 573
rect 861 505 929 541
rect 1106 540 1175 634
rect 1106 508 1120 540
rect 1152 508 1175 540
rect 1106 459 1175 508
rect 1106 427 1120 459
rect 1152 427 1175 459
rect 1106 410 1175 427
rect 1201 410 1320 634
rect 1346 467 1414 634
rect 1539 475 1607 629
rect 1346 435 1368 467
rect 1400 435 1414 467
rect 1346 410 1414 435
rect 1539 443 1553 475
rect 1585 443 1607 475
rect 1539 429 1607 443
rect 1633 513 1683 629
rect 1862 513 1922 720
rect 2086 670 2146 720
rect 2086 638 2100 670
rect 2132 638 2146 670
rect 2086 629 2146 638
rect 2086 602 2160 629
rect 2086 570 2100 602
rect 2132 570 2160 602
rect 2086 534 2160 570
rect 2086 513 2100 534
rect 1633 487 1746 513
rect 1633 455 1692 487
rect 1724 455 1746 487
rect 1633 429 1746 455
rect 1772 429 1822 513
rect 1848 429 1944 513
rect 1970 489 2046 513
rect 1970 457 1992 489
rect 2024 457 2046 489
rect 1970 429 2046 457
rect 2072 502 2100 513
rect 2132 502 2160 534
rect 2072 429 2160 502
rect 2186 611 2254 629
rect 2186 579 2208 611
rect 2240 579 2254 611
rect 2186 543 2254 579
rect 2186 511 2208 543
rect 2240 511 2254 543
rect 2186 475 2254 511
rect 2186 443 2208 475
rect 2240 443 2254 475
rect 2186 429 2254 443
rect 2382 622 2450 636
rect 2382 590 2396 622
rect 2428 590 2450 622
rect 2382 554 2450 590
rect 2382 522 2396 554
rect 2428 522 2450 554
rect 2382 486 2450 522
rect 2382 454 2396 486
rect 2428 454 2450 486
rect 2382 412 2450 454
rect 2476 622 2553 636
rect 2476 590 2498 622
rect 2530 590 2553 622
rect 2476 554 2553 590
rect 2476 522 2498 554
rect 2530 522 2553 554
rect 2476 486 2553 522
rect 2476 454 2498 486
rect 2530 454 2553 486
rect 2476 412 2553 454
rect 2579 622 2647 636
rect 2579 590 2601 622
rect 2633 590 2647 622
rect 2579 554 2647 590
rect 2579 522 2601 554
rect 2633 522 2647 554
rect 2579 486 2647 522
rect 2579 454 2601 486
rect 2633 454 2647 486
rect 2579 412 2647 454
<< ndiffc >>
rect 52 135 84 167
rect 238 135 270 167
rect 687 286 719 318
rect 789 312 821 344
rect 926 298 958 330
rect 354 176 386 208
rect 457 141 489 173
rect 643 159 675 191
rect 1041 237 1073 269
rect 1363 172 1395 204
rect 1503 215 1535 247
rect 1605 229 1637 261
rect 1718 92 1750 124
rect 1820 135 1852 167
rect 1922 135 1954 167
rect 2086 135 2118 167
rect 2190 196 2222 228
rect 2190 128 2222 160
rect 2292 196 2324 228
rect 2292 128 2324 160
rect 2396 196 2428 228
rect 2396 128 2428 160
rect 2498 196 2530 228
rect 2498 128 2530 160
rect 2601 196 2633 228
rect 2601 128 2633 160
<< pdiffc >>
rect 53 633 85 665
rect 52 458 84 490
rect 154 459 186 491
rect 346 538 378 570
rect 452 538 484 570
rect 590 582 622 614
rect 781 519 813 551
rect 883 541 915 573
rect 1120 508 1152 540
rect 1120 427 1152 459
rect 1368 435 1400 467
rect 1553 443 1585 475
rect 2100 638 2132 670
rect 2100 570 2132 602
rect 1692 455 1724 487
rect 1992 457 2024 489
rect 2100 502 2132 534
rect 2208 579 2240 611
rect 2208 511 2240 543
rect 2208 443 2240 475
rect 2396 590 2428 622
rect 2396 522 2428 554
rect 2396 454 2428 486
rect 2498 590 2530 622
rect 2498 522 2530 554
rect 2498 454 2530 486
rect 2601 590 2633 622
rect 2601 522 2633 554
rect 2601 454 2633 486
<< psubdiff >>
rect 1136 30 1196 36
rect 0 16 2688 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2528 16
rect 2560 -16 2624 16
rect 2656 -16 2688 16
rect 0 -30 2688 -16
<< nsubdiff >>
rect 0 772 2688 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2528 772
rect 2560 740 2624 772
rect 2656 740 2688 772
rect 0 726 2688 740
rect 1215 720 1306 726
rect 1862 720 1922 726
rect 2086 720 2146 726
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
rect 1280 -16 1312 16
rect 1376 -16 1408 16
rect 1472 -16 1504 16
rect 1568 -16 1600 16
rect 1664 -16 1696 16
rect 1760 -16 1792 16
rect 1856 -16 1888 16
rect 1952 -16 1984 16
rect 2048 -16 2080 16
rect 2144 -16 2176 16
rect 2240 -16 2272 16
rect 2336 -16 2368 16
rect 2432 -16 2464 16
rect 2528 -16 2560 16
rect 2624 -16 2656 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
rect 1280 740 1312 772
rect 1376 740 1408 772
rect 1472 740 1504 772
rect 1568 740 1600 772
rect 1664 740 1696 772
rect 1760 740 1792 772
rect 1856 740 1888 772
rect 1952 740 1984 772
rect 2048 740 2080 772
rect 2144 740 2176 772
rect 2240 740 2272 772
rect 2336 740 2368 772
rect 2432 740 2464 772
rect 2528 740 2560 772
rect 2624 740 2656 772
<< poly >>
rect 298 632 324 668
rect 508 661 1027 687
rect 106 516 132 552
rect 208 516 234 552
rect 508 589 534 661
rect 967 647 1027 661
rect 655 589 681 625
rect 733 589 759 625
rect 835 589 861 625
rect 967 615 981 647
rect 1013 615 1027 647
rect 1175 634 1201 670
rect 1320 634 1346 670
rect 967 601 1027 615
rect 106 354 132 432
rect 208 396 234 432
rect 47 340 132 354
rect 47 308 61 340
rect 93 308 132 340
rect 47 294 132 308
rect 106 198 132 294
rect 190 330 234 396
rect 298 397 324 432
rect 508 397 534 505
rect 655 397 681 505
rect 298 383 373 397
rect 298 351 327 383
rect 359 351 373 383
rect 298 337 373 351
rect 490 383 550 397
rect 490 351 504 383
rect 536 351 550 383
rect 490 337 550 351
rect 190 198 216 330
rect 306 307 332 337
rect 524 211 550 337
rect 587 383 681 397
rect 587 351 601 383
rect 633 371 681 383
rect 733 401 759 505
rect 835 488 861 505
rect 835 472 1060 488
rect 835 458 1014 472
rect 733 371 767 401
rect 633 351 647 371
rect 741 356 767 371
rect 843 356 869 458
rect 1000 440 1014 458
rect 1046 440 1060 472
rect 1000 425 1060 440
rect 1607 629 1633 665
rect 1449 457 1509 471
rect 1449 425 1463 457
rect 1495 425 1509 457
rect 1746 513 1772 549
rect 1822 513 1848 549
rect 1979 647 2039 661
rect 1979 628 1993 647
rect 1944 615 1993 628
rect 2025 615 2039 647
rect 1944 601 2039 615
rect 2160 629 2186 665
rect 2450 636 2476 672
rect 2553 636 2579 672
rect 1944 513 1970 601
rect 2046 513 2072 549
rect 1449 414 1509 425
rect 1607 414 1633 429
rect 1449 411 1633 414
rect 1175 374 1201 410
rect 1320 374 1346 410
rect 1480 384 1633 411
rect 1095 357 1210 374
rect 587 337 647 351
rect 587 211 613 337
rect 1095 325 1147 357
rect 1179 325 1210 357
rect 1320 357 1404 374
rect 1320 338 1355 357
rect 1095 308 1210 325
rect 1315 325 1355 338
rect 1387 325 1404 357
rect 1315 308 1404 325
rect 1095 283 1121 308
rect 1315 283 1341 308
rect 306 123 332 159
rect 106 78 132 114
rect 190 86 216 114
rect 524 86 550 127
rect 190 59 550 86
rect 587 85 613 127
rect 741 121 767 272
rect 843 236 869 272
rect 1557 275 1583 384
rect 1746 361 1772 429
rect 1822 397 1848 429
rect 1664 344 1772 361
rect 1664 312 1678 344
rect 1710 335 1772 344
rect 1811 380 1877 397
rect 1811 348 1828 380
rect 1860 348 1877 380
rect 1710 312 1724 335
rect 1811 331 1877 348
rect 1944 363 1970 429
rect 1664 295 1724 312
rect 1664 275 1690 295
rect 1557 153 1583 191
rect 1095 121 1121 135
rect 741 93 1121 121
rect 1315 99 1341 135
rect 1841 243 1871 331
rect 1944 330 1983 363
rect 2046 337 2072 429
rect 2160 337 2186 429
rect 2328 349 2388 363
rect 1841 213 1900 243
rect 1874 198 1900 213
rect 1957 239 1983 330
rect 2030 323 2270 337
rect 2030 291 2044 323
rect 2076 311 2270 323
rect 2076 291 2090 311
rect 2030 277 2090 291
rect 1957 212 2002 239
rect 1976 198 2002 212
rect 2038 198 2064 277
rect 2244 242 2270 311
rect 2328 317 2342 349
rect 2374 330 2388 349
rect 2450 330 2476 412
rect 2553 330 2579 412
rect 2374 317 2579 330
rect 2328 303 2579 317
rect 2450 262 2476 303
rect 2553 262 2579 303
rect 1664 89 1690 127
rect 1874 78 1900 114
rect 1976 78 2002 114
rect 2038 78 2064 114
rect 2244 78 2270 114
rect 2450 78 2476 114
rect 2553 78 2579 114
<< polycont >>
rect 981 615 1013 647
rect 61 308 93 340
rect 327 351 359 383
rect 504 351 536 383
rect 601 351 633 383
rect 1014 440 1046 472
rect 1463 425 1495 457
rect 1993 615 2025 647
rect 1147 325 1179 357
rect 1355 325 1387 357
rect 1678 312 1710 344
rect 1828 348 1860 380
rect 2044 291 2076 323
rect 2342 317 2374 349
<< metal1 >>
rect 0 772 2688 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2528 772
rect 2560 740 2624 772
rect 2656 740 2688 772
rect 0 712 2688 740
rect 43 665 94 712
rect 43 633 53 665
rect 85 633 94 665
rect 43 490 94 633
rect 158 616 553 648
rect 158 504 196 616
rect 43 458 52 490
rect 84 458 94 490
rect 43 443 94 458
rect 144 491 196 504
rect 144 459 154 491
rect 186 459 196 491
rect 144 448 196 459
rect 240 570 388 580
rect 240 538 346 570
rect 378 538 388 570
rect 240 528 388 538
rect 449 570 485 580
rect 449 538 452 570
rect 484 538 485 570
rect 51 340 122 371
rect 51 308 61 340
rect 93 308 122 340
rect 51 275 122 308
rect 158 168 190 448
rect 240 266 272 528
rect 449 463 485 538
rect 521 536 553 616
rect 589 614 623 712
rect 2090 670 2142 712
rect 971 647 1023 657
rect 1982 647 2036 657
rect 589 582 590 614
rect 622 582 623 614
rect 589 572 623 582
rect 691 597 925 629
rect 971 615 981 647
rect 1013 615 1993 647
rect 2025 615 2036 647
rect 971 605 1023 615
rect 1982 605 2036 615
rect 2090 638 2100 670
rect 2132 638 2142 670
rect 691 536 723 597
rect 858 573 925 597
rect 521 504 723 536
rect 778 551 815 561
rect 778 519 781 551
rect 813 519 815 551
rect 778 463 815 519
rect 449 461 815 463
rect 317 429 815 461
rect 317 383 369 429
rect 317 351 327 383
rect 359 351 369 383
rect 317 341 369 351
rect 440 383 550 393
rect 440 351 504 383
rect 536 351 550 383
rect 440 302 550 351
rect 587 383 643 393
rect 587 351 601 383
rect 633 351 643 383
rect 778 362 815 429
rect 858 541 883 573
rect 915 541 925 573
rect 2090 602 2142 638
rect 2386 622 2438 712
rect 2090 570 2100 602
rect 2132 570 2142 602
rect 858 537 925 541
rect 1085 540 1655 558
rect 587 266 619 351
rect 778 344 822 362
rect 240 234 619 266
rect 677 318 729 328
rect 677 286 687 318
rect 719 286 729 318
rect 778 312 789 344
rect 821 312 822 344
rect 778 302 822 312
rect 677 266 729 286
rect 858 266 890 537
rect 1085 508 1120 540
rect 1152 526 1655 540
rect 1152 508 1157 526
rect 1085 482 1157 508
rect 1004 472 1157 482
rect 1549 475 1587 490
rect 1004 440 1014 472
rect 1046 459 1157 472
rect 1046 440 1120 459
rect 1004 430 1120 440
rect 1031 427 1120 430
rect 1152 427 1157 459
rect 1031 412 1157 427
rect 1193 467 1505 474
rect 1193 435 1368 467
rect 1400 457 1505 467
rect 1400 435 1463 457
rect 1193 429 1463 435
rect 926 330 979 340
rect 958 298 979 330
rect 926 288 979 298
rect 677 245 890 266
rect 693 234 890 245
rect 937 260 979 288
rect 1031 269 1083 412
rect 1193 374 1225 429
rect 1453 425 1463 429
rect 1495 425 1505 457
rect 1453 415 1505 425
rect 1549 443 1553 475
rect 1585 443 1587 475
rect 1130 357 1225 374
rect 1130 325 1147 357
rect 1179 325 1225 357
rect 1130 308 1225 325
rect 344 208 396 234
rect 42 167 190 168
rect 42 135 52 167
rect 84 135 190 167
rect 42 129 190 135
rect 228 167 280 177
rect 228 135 238 167
rect 270 135 280 167
rect 344 176 354 208
rect 386 176 396 208
rect 344 163 396 176
rect 447 173 499 183
rect 228 44 280 135
rect 447 141 457 173
rect 489 141 499 173
rect 447 44 499 141
rect 541 121 575 234
rect 937 192 973 260
rect 1031 237 1041 269
rect 1073 237 1083 269
rect 1031 227 1083 237
rect 633 191 973 192
rect 633 159 643 191
rect 675 159 973 191
rect 1193 205 1225 308
rect 1273 357 1398 387
rect 1273 325 1355 357
rect 1387 325 1398 357
rect 1549 345 1587 443
rect 1273 267 1398 325
rect 1434 311 1587 345
rect 1623 354 1655 526
rect 2090 534 2142 570
rect 2090 502 2100 534
rect 2132 502 2142 534
rect 1691 487 1732 500
rect 1691 455 1692 487
rect 1724 459 1732 487
rect 1982 489 2034 499
rect 2090 492 2142 502
rect 2198 611 2250 621
rect 2198 579 2208 611
rect 2240 579 2250 611
rect 2198 543 2250 579
rect 2198 511 2208 543
rect 2240 511 2250 543
rect 1724 455 1790 459
rect 1691 425 1790 455
rect 1982 457 1992 489
rect 2024 457 2034 489
rect 1982 452 2034 457
rect 2198 475 2250 511
rect 1623 344 1720 354
rect 1623 312 1678 344
rect 1710 312 1720 344
rect 1351 205 1398 214
rect 1193 204 1398 205
rect 1193 172 1363 204
rect 1395 172 1398 204
rect 1193 171 1398 172
rect 1351 162 1398 171
rect 633 157 973 159
rect 1434 121 1466 311
rect 1623 302 1720 312
rect 1758 293 1790 425
rect 1826 420 2146 452
rect 1826 380 1877 420
rect 1826 348 1828 380
rect 1860 348 1877 380
rect 1826 331 1877 348
rect 2033 323 2078 333
rect 2033 293 2044 323
rect 1758 291 2044 293
rect 2076 291 2078 323
rect 1758 263 2078 291
rect 1502 247 1536 262
rect 1502 215 1503 247
rect 1535 215 1536 247
rect 1592 261 2078 263
rect 1592 229 1605 261
rect 1637 255 2078 261
rect 1637 229 1794 255
rect 1502 193 1536 215
rect 1502 167 1862 193
rect 2114 177 2146 420
rect 2198 443 2208 475
rect 2240 443 2250 475
rect 2198 359 2250 443
rect 2386 590 2396 622
rect 2428 590 2438 622
rect 2386 554 2438 590
rect 2386 522 2396 554
rect 2428 522 2438 554
rect 2386 486 2438 522
rect 2386 454 2396 486
rect 2428 454 2438 486
rect 2386 438 2438 454
rect 2488 622 2540 632
rect 2488 590 2498 622
rect 2530 590 2540 622
rect 2488 554 2540 590
rect 2488 522 2498 554
rect 2530 522 2540 554
rect 2488 486 2540 522
rect 2488 454 2498 486
rect 2530 454 2540 486
rect 2488 369 2540 454
rect 2591 622 2643 712
rect 2591 590 2601 622
rect 2633 590 2643 622
rect 2591 554 2643 590
rect 2591 522 2601 554
rect 2633 522 2643 554
rect 2591 486 2643 522
rect 2591 454 2601 486
rect 2633 454 2643 486
rect 2591 444 2643 454
rect 2198 349 2384 359
rect 2198 317 2342 349
rect 2374 317 2384 349
rect 2198 311 2384 317
rect 2282 308 2384 311
rect 1502 161 1820 167
rect 1810 135 1820 161
rect 1852 135 1862 167
rect 1810 125 1862 135
rect 1912 167 1964 177
rect 1912 135 1922 167
rect 1954 135 1964 167
rect 1708 124 1760 125
rect 1708 121 1718 124
rect 541 92 1718 121
rect 1750 92 1760 124
rect 541 88 1760 92
rect 1912 44 1964 135
rect 2076 167 2146 177
rect 2076 135 2086 167
rect 2118 135 2146 167
rect 2076 125 2146 135
rect 2185 228 2232 238
rect 2185 196 2190 228
rect 2222 196 2232 228
rect 2185 160 2232 196
rect 2185 128 2190 160
rect 2222 128 2232 160
rect 2185 44 2232 128
rect 2282 228 2334 308
rect 2488 301 2630 369
rect 2282 196 2292 228
rect 2324 196 2334 228
rect 2282 160 2334 196
rect 2282 128 2292 160
rect 2324 128 2334 160
rect 2282 118 2334 128
rect 2387 228 2440 240
rect 2387 196 2396 228
rect 2428 196 2440 228
rect 2387 160 2440 196
rect 2387 128 2396 160
rect 2428 128 2440 160
rect 2387 44 2440 128
rect 2488 228 2540 301
rect 2488 196 2498 228
rect 2530 196 2540 228
rect 2488 160 2540 196
rect 2488 128 2498 160
rect 2530 128 2540 160
rect 2488 119 2540 128
rect 2592 228 2643 240
rect 2592 196 2601 228
rect 2633 196 2643 228
rect 2592 160 2643 196
rect 2592 128 2601 160
rect 2633 128 2643 160
rect 2592 44 2643 128
rect 0 16 2688 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2528 16
rect 2560 -16 2624 16
rect 2656 -16 2688 16
rect 0 -44 2688 -16
<< labels >>
flabel metal1 s 1273 267 1398 387 0 FreeSans 400 0 0 0 CLK
port 2 nsew
flabel metal1 s 0 -44 2688 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 51 275 122 371 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel metal1 s 2488 301 2630 369 0 FreeSans 340 0 0 0 Q
port 5 nsew
flabel metal1 s 0 712 2688 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s 440 302 550 393 0 FreeSans 400 0 0 0 RESET_B
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 756
string GDS_END 94406
string GDS_FILE 6_final.gds
string GDS_START 79402
<< end >>
