magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< error_p >>
rect -2110 15430 -2101 15439
rect 2101 15430 2110 15439
rect 2330 15430 2339 15439
rect 6541 15430 6550 15439
rect -2119 15421 -2110 15430
rect 2110 15421 2119 15430
rect -2119 11210 -2110 11219
rect 2110 11210 2119 11219
rect 2321 11210 2330 11219
rect 6550 11210 6559 11219
rect -2110 11201 -2101 11210
rect 2101 11201 2110 11210
rect 2330 11201 2339 11210
rect 6541 11201 6550 11210
rect -2110 10990 -2101 10999
rect 2101 10990 2110 10999
rect 2330 10990 2339 10999
rect 6541 10990 6550 10999
rect -2119 10981 -2110 10990
rect 2110 10981 2119 10990
rect -2119 6770 -2110 6779
rect 2110 6770 2119 6779
rect 2321 6770 2330 6779
rect 6550 6770 6559 6779
rect -2110 6761 -2101 6770
rect 2101 6761 2110 6770
rect 2330 6761 2339 6770
rect 6541 6761 6550 6770
rect -2110 6550 -2101 6559
rect 2101 6550 2110 6559
rect 2330 6550 2339 6559
rect 6541 6550 6550 6559
rect -2119 6541 -2110 6550
rect 2110 6541 2119 6550
rect -2119 2330 -2110 2339
rect 2110 2330 2119 2339
rect 2321 2330 2330 2339
rect 6550 2330 6559 2339
rect -2110 2321 -2101 2330
rect 2101 2321 2110 2330
rect 2330 2321 2339 2330
rect 6541 2321 6550 2330
rect -2110 2110 -2101 2119
rect 2101 2110 2110 2119
rect 2330 2110 2339 2119
rect 6541 2110 6550 2119
rect -2119 2101 -2110 2110
rect 2110 2101 2119 2110
rect -2119 -2110 -2110 -2101
rect 2110 -2110 2119 -2101
rect 2321 -2110 2330 -2101
rect 6550 -2110 6559 -2101
rect -2110 -2119 -2101 -2110
rect 2101 -2119 2110 -2110
rect 2330 -2119 2339 -2110
rect 6541 -2119 6550 -2110
<< via4 >>
rect -2110 11210 2110 15430
rect 2330 11210 6550 15430
rect -2110 6770 2110 10990
rect 2330 6770 6550 10990
rect -2110 2330 2110 6550
rect 2330 2330 6550 6550
rect -2110 -2110 2110 2110
rect 2330 -2110 6550 2110
<< metal5 >>
rect -2120 15430 2120 15440
rect -2120 11210 -2110 15430
rect 2110 11210 2120 15430
rect -2120 11200 2120 11210
rect 2320 15430 6560 15440
rect 2320 11210 2330 15430
rect 6550 11210 6560 15430
rect 2320 11200 6560 11210
rect -2120 10990 2120 11000
rect -2120 6770 -2110 10990
rect 2110 6770 2120 10990
rect -2120 6760 2120 6770
rect 2320 10990 6560 11000
rect 2320 6770 2330 10990
rect 6550 6770 6560 10990
rect 2320 6760 6560 6770
rect -2120 6550 2120 6560
rect -2120 2330 -2110 6550
rect 2110 2330 2120 6550
rect -2120 2320 2120 2330
rect 2320 6550 6560 6560
rect 2320 2330 2330 6550
rect 6550 2330 6560 6550
rect 2320 2320 6560 2330
rect -2120 2110 2120 2120
rect -2120 -2110 -2110 2110
rect 2110 -2110 2120 2110
rect -2120 -2120 2120 -2110
rect 2320 2110 6560 2120
rect 2320 -2110 2330 2110
rect 6550 -2110 6560 2110
rect 2320 -2120 6560 -2110
<< mimcap >>
rect -2000 15248 2000 15320
rect -2000 11392 -1928 15248
rect 1928 11392 2000 15248
rect -2000 11320 2000 11392
rect 2440 15248 6440 15320
rect 2440 11392 2512 15248
rect 6368 11392 6440 15248
rect 2440 11320 6440 11392
rect -2000 10808 2000 10880
rect -2000 6952 -1928 10808
rect 1928 6952 2000 10808
rect -2000 6880 2000 6952
rect 2440 10808 6440 10880
rect 2440 6952 2512 10808
rect 6368 6952 6440 10808
rect 2440 6880 6440 6952
rect -2000 6368 2000 6440
rect -2000 2512 -1928 6368
rect 1928 2512 2000 6368
rect -2000 2440 2000 2512
rect 2440 6368 6440 6440
rect 2440 2512 2512 6368
rect 6368 2512 6440 6368
rect 2440 2440 6440 2512
rect -2000 1928 2000 2000
rect -2000 -1928 -1928 1928
rect 1928 -1928 2000 1928
rect -2000 -2000 2000 -1928
rect 2440 1928 6440 2000
rect 2440 -1928 2512 1928
rect 6368 -1928 6440 1928
rect 2440 -2000 6440 -1928
<< mimcapcontact >>
rect -1928 11392 1928 15248
rect 2512 11392 6368 15248
rect -1928 6952 1928 10808
rect 2512 6952 6368 10808
rect -1928 2512 1928 6368
rect 2512 2512 6368 6368
rect -1928 -1928 1928 1928
rect 2512 -1928 6368 1928
<< properties >>
string gencell cmim
string library sg13g2_devstdin
string parameters w 20 l 20 nx 2 dx 1 ny 4 dy 1 wmin 1.14 lmin 1.14 class capacitor topcc 100 botcc 100
<< end >>
