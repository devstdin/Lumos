magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect -3 56 342 281
rect -26 -56 410 56
<< nmos >>
rect 97 195 123 255
rect 221 96 247 255
<< pmos >>
rect 97 429 123 561
rect 222 429 248 660
<< ndiff >>
rect 23 241 97 255
rect 23 209 37 241
rect 69 209 97 241
rect 23 195 97 209
rect 123 195 221 255
rect 148 142 221 195
rect 148 110 162 142
rect 194 110 221 142
rect 148 96 221 110
rect 247 239 316 255
rect 247 207 270 239
rect 302 207 316 239
rect 247 96 316 207
rect 148 36 202 96
<< pdiff >>
rect 23 661 204 720
rect 23 629 37 661
rect 69 660 204 661
rect 69 629 222 660
rect 23 615 222 629
rect 141 561 222 615
rect 23 480 97 561
rect 23 448 37 480
rect 69 448 97 480
rect 23 429 97 448
rect 123 429 222 561
rect 248 563 316 660
rect 248 531 270 563
rect 302 531 316 563
rect 248 475 316 531
rect 248 443 270 475
rect 302 443 316 475
rect 248 429 316 443
<< ndiffc >>
rect 37 209 69 241
rect 162 110 194 142
rect 270 207 302 239
<< pdiffc >>
rect 37 629 69 661
rect 37 448 69 480
rect 270 531 302 563
rect 270 443 302 475
<< psubdiff >>
rect 148 30 202 36
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
rect 23 720 204 726
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 222 660 248 698
rect 97 561 123 599
rect 97 331 123 429
rect 222 395 248 429
rect 222 381 326 395
rect 222 366 280 381
rect 266 349 280 366
rect 312 349 326 381
rect 266 335 326 349
rect 23 317 123 331
rect 23 285 37 317
rect 69 285 123 317
rect 23 271 123 285
rect 97 255 123 271
rect 169 315 229 329
rect 169 283 183 315
rect 215 298 229 315
rect 215 283 247 298
rect 169 269 247 283
rect 221 255 247 269
rect 97 157 123 195
rect 221 60 247 96
<< polycont >>
rect 280 349 312 381
rect 37 285 69 317
rect 183 283 215 315
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 27 661 79 712
rect 27 629 37 661
rect 69 629 79 661
rect 27 619 79 629
rect 260 563 317 582
rect 260 531 270 563
rect 302 531 317 563
rect 27 480 79 490
rect 27 448 37 480
rect 69 448 79 480
rect 27 438 79 448
rect 39 406 79 438
rect 260 475 317 531
rect 260 443 270 475
rect 302 443 317 475
rect 260 433 317 443
rect 39 363 224 406
rect 27 317 79 327
rect 27 285 37 317
rect 69 285 79 317
rect 27 241 79 285
rect 174 315 224 363
rect 174 283 183 315
rect 215 283 224 315
rect 174 271 224 283
rect 260 381 315 391
rect 260 349 280 381
rect 312 349 315 381
rect 27 209 37 241
rect 69 209 79 241
rect 27 199 79 209
rect 260 239 315 349
rect 260 207 270 239
rect 302 207 315 239
rect 260 197 315 207
rect 152 142 204 152
rect 152 110 162 142
rect 194 110 204 142
rect 152 44 204 110
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 260 433 317 582 0 FreeSans 400 0 0 0 L_HI
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 75094
string GDS_FILE 6_final.gds
string GDS_START 71706
<< end >>
