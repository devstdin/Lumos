magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2026 3448 3820
<< nwell >>
rect -124 1116 1448 1820
<< pwell >>
rect -26 854 602 974
rect -26 94 94 854
rect 482 94 602 854
rect -26 -26 602 94
rect 842 -26 1350 974
<< psubdiff >>
rect 0 930 576 948
rect 0 898 34 930
rect 66 898 102 930
rect 134 898 170 930
rect 202 898 238 930
rect 270 898 306 930
rect 338 898 374 930
rect 406 898 442 930
rect 474 898 510 930
rect 542 898 576 930
rect 0 880 576 898
rect 0 830 68 880
rect 0 798 18 830
rect 50 798 68 830
rect 0 762 68 798
rect 0 730 18 762
rect 50 730 68 762
rect 508 830 576 880
rect 508 798 526 830
rect 558 798 576 830
rect 508 762 576 798
rect 0 694 68 730
rect 0 662 18 694
rect 50 662 68 694
rect 0 626 68 662
rect 0 594 18 626
rect 50 594 68 626
rect 0 558 68 594
rect 0 526 18 558
rect 50 526 68 558
rect 0 490 68 526
rect 0 458 18 490
rect 50 458 68 490
rect 0 422 68 458
rect 0 390 18 422
rect 50 390 68 422
rect 0 354 68 390
rect 0 322 18 354
rect 50 322 68 354
rect 0 286 68 322
rect 0 254 18 286
rect 50 254 68 286
rect 0 218 68 254
rect 0 186 18 218
rect 50 186 68 218
rect 508 730 526 762
rect 558 730 576 762
rect 508 694 576 730
rect 508 662 526 694
rect 558 662 576 694
rect 508 626 576 662
rect 508 594 526 626
rect 558 594 576 626
rect 508 558 576 594
rect 508 526 526 558
rect 558 526 576 558
rect 508 490 576 526
rect 508 458 526 490
rect 558 458 576 490
rect 508 422 576 458
rect 508 390 526 422
rect 558 390 576 422
rect 508 354 576 390
rect 508 322 526 354
rect 558 322 576 354
rect 508 286 576 322
rect 508 254 526 286
rect 558 254 576 286
rect 508 218 576 254
rect 0 150 68 186
rect 0 118 18 150
rect 50 118 68 150
rect 0 68 68 118
rect 508 186 526 218
rect 558 186 576 218
rect 508 150 576 186
rect 508 118 526 150
rect 558 118 576 150
rect 508 68 576 118
rect 0 50 576 68
rect 0 18 34 50
rect 66 18 102 50
rect 134 18 170 50
rect 202 18 238 50
rect 270 18 306 50
rect 338 18 374 50
rect 406 18 442 50
rect 474 18 510 50
rect 542 18 576 50
rect 0 0 576 18
rect 868 930 1324 948
rect 868 898 910 930
rect 942 898 978 930
rect 1010 898 1046 930
rect 1078 898 1114 930
rect 1146 898 1182 930
rect 1214 898 1250 930
rect 1282 898 1324 930
rect 868 880 1324 898
rect 868 830 936 880
rect 868 798 886 830
rect 918 798 936 830
rect 868 762 936 798
rect 1256 830 1324 880
rect 1256 798 1274 830
rect 1306 798 1324 830
rect 868 730 886 762
rect 918 730 936 762
rect 868 694 936 730
rect 868 662 886 694
rect 918 662 936 694
rect 868 626 936 662
rect 868 594 886 626
rect 918 594 936 626
rect 868 558 936 594
rect 868 526 886 558
rect 918 526 936 558
rect 868 490 936 526
rect 868 458 886 490
rect 918 458 936 490
rect 868 422 936 458
rect 868 390 886 422
rect 918 390 936 422
rect 868 354 936 390
rect 868 322 886 354
rect 918 322 936 354
rect 868 286 936 322
rect 868 254 886 286
rect 918 254 936 286
rect 868 218 936 254
rect 868 186 886 218
rect 918 186 936 218
rect 868 150 936 186
rect 1256 762 1324 798
rect 1256 730 1274 762
rect 1306 730 1324 762
rect 1256 694 1324 730
rect 1256 662 1274 694
rect 1306 662 1324 694
rect 1256 626 1324 662
rect 1256 594 1274 626
rect 1306 594 1324 626
rect 1256 558 1324 594
rect 1256 526 1274 558
rect 1306 526 1324 558
rect 1256 490 1324 526
rect 1256 458 1274 490
rect 1306 458 1324 490
rect 1256 422 1324 458
rect 1256 390 1274 422
rect 1306 390 1324 422
rect 1256 354 1324 390
rect 1256 322 1274 354
rect 1306 322 1324 354
rect 1256 286 1324 322
rect 1256 254 1274 286
rect 1306 254 1324 286
rect 1256 218 1324 254
rect 1256 186 1274 218
rect 1306 186 1324 218
rect 868 118 886 150
rect 918 118 936 150
rect 868 68 936 118
rect 1256 150 1324 186
rect 1256 118 1274 150
rect 1306 118 1324 150
rect 1256 68 1324 118
rect 868 50 1324 68
rect 868 18 910 50
rect 942 18 978 50
rect 1010 18 1046 50
rect 1078 18 1114 50
rect 1146 18 1182 50
rect 1214 18 1250 50
rect 1282 18 1324 50
rect 868 0 1324 18
<< nsubdiff >>
rect 0 1678 1324 1696
rect 0 1646 34 1678
rect 66 1646 102 1678
rect 134 1646 170 1678
rect 202 1646 238 1678
rect 270 1646 306 1678
rect 338 1646 374 1678
rect 406 1646 442 1678
rect 474 1646 510 1678
rect 542 1646 578 1678
rect 610 1646 646 1678
rect 678 1646 714 1678
rect 746 1646 782 1678
rect 814 1646 850 1678
rect 882 1646 918 1678
rect 950 1646 986 1678
rect 1018 1646 1054 1678
rect 1086 1646 1122 1678
rect 1154 1646 1190 1678
rect 1222 1646 1258 1678
rect 1290 1646 1324 1678
rect 0 1628 1324 1646
rect 0 1586 68 1628
rect 0 1554 18 1586
rect 50 1554 68 1586
rect 0 1518 68 1554
rect 1256 1586 1324 1628
rect 1256 1554 1274 1586
rect 1306 1554 1324 1586
rect 0 1486 18 1518
rect 50 1486 68 1518
rect 0 1450 68 1486
rect 0 1418 18 1450
rect 50 1418 68 1450
rect 0 1382 68 1418
rect 1256 1518 1324 1554
rect 1256 1486 1274 1518
rect 1306 1486 1324 1518
rect 1256 1450 1324 1486
rect 1256 1418 1274 1450
rect 1306 1418 1324 1450
rect 0 1350 18 1382
rect 50 1350 68 1382
rect 0 1308 68 1350
rect 1256 1382 1324 1418
rect 1256 1350 1274 1382
rect 1306 1350 1324 1382
rect 1256 1308 1324 1350
rect 0 1290 1324 1308
rect 0 1258 34 1290
rect 66 1258 102 1290
rect 134 1258 170 1290
rect 202 1258 238 1290
rect 270 1258 306 1290
rect 338 1258 374 1290
rect 406 1258 442 1290
rect 474 1258 510 1290
rect 542 1258 578 1290
rect 610 1258 646 1290
rect 678 1258 714 1290
rect 746 1258 782 1290
rect 814 1258 850 1290
rect 882 1258 918 1290
rect 950 1258 986 1290
rect 1018 1258 1054 1290
rect 1086 1258 1122 1290
rect 1154 1258 1190 1290
rect 1222 1258 1258 1290
rect 1290 1258 1324 1290
rect 0 1240 1324 1258
<< psubdiffcont >>
rect 34 898 66 930
rect 102 898 134 930
rect 170 898 202 930
rect 238 898 270 930
rect 306 898 338 930
rect 374 898 406 930
rect 442 898 474 930
rect 510 898 542 930
rect 18 798 50 830
rect 18 730 50 762
rect 526 798 558 830
rect 18 662 50 694
rect 18 594 50 626
rect 18 526 50 558
rect 18 458 50 490
rect 18 390 50 422
rect 18 322 50 354
rect 18 254 50 286
rect 18 186 50 218
rect 526 730 558 762
rect 526 662 558 694
rect 526 594 558 626
rect 526 526 558 558
rect 526 458 558 490
rect 526 390 558 422
rect 526 322 558 354
rect 526 254 558 286
rect 18 118 50 150
rect 526 186 558 218
rect 526 118 558 150
rect 34 18 66 50
rect 102 18 134 50
rect 170 18 202 50
rect 238 18 270 50
rect 306 18 338 50
rect 374 18 406 50
rect 442 18 474 50
rect 510 18 542 50
rect 910 898 942 930
rect 978 898 1010 930
rect 1046 898 1078 930
rect 1114 898 1146 930
rect 1182 898 1214 930
rect 1250 898 1282 930
rect 886 798 918 830
rect 1274 798 1306 830
rect 886 730 918 762
rect 886 662 918 694
rect 886 594 918 626
rect 886 526 918 558
rect 886 458 918 490
rect 886 390 918 422
rect 886 322 918 354
rect 886 254 918 286
rect 886 186 918 218
rect 1274 730 1306 762
rect 1274 662 1306 694
rect 1274 594 1306 626
rect 1274 526 1306 558
rect 1274 458 1306 490
rect 1274 390 1306 422
rect 1274 322 1306 354
rect 1274 254 1306 286
rect 1274 186 1306 218
rect 886 118 918 150
rect 1274 118 1306 150
rect 910 18 942 50
rect 978 18 1010 50
rect 1046 18 1078 50
rect 1114 18 1146 50
rect 1182 18 1214 50
rect 1250 18 1282 50
<< nsubdiffcont >>
rect 34 1646 66 1678
rect 102 1646 134 1678
rect 170 1646 202 1678
rect 238 1646 270 1678
rect 306 1646 338 1678
rect 374 1646 406 1678
rect 442 1646 474 1678
rect 510 1646 542 1678
rect 578 1646 610 1678
rect 646 1646 678 1678
rect 714 1646 746 1678
rect 782 1646 814 1678
rect 850 1646 882 1678
rect 918 1646 950 1678
rect 986 1646 1018 1678
rect 1054 1646 1086 1678
rect 1122 1646 1154 1678
rect 1190 1646 1222 1678
rect 1258 1646 1290 1678
rect 18 1554 50 1586
rect 1274 1554 1306 1586
rect 18 1486 50 1518
rect 18 1418 50 1450
rect 1274 1486 1306 1518
rect 1274 1418 1306 1450
rect 18 1350 50 1382
rect 1274 1350 1306 1382
rect 34 1258 66 1290
rect 102 1258 134 1290
rect 170 1258 202 1290
rect 238 1258 270 1290
rect 306 1258 338 1290
rect 374 1258 406 1290
rect 442 1258 474 1290
rect 510 1258 542 1290
rect 578 1258 610 1290
rect 646 1258 678 1290
rect 714 1258 746 1290
rect 782 1258 814 1290
rect 850 1258 882 1290
rect 918 1258 950 1290
rect 986 1258 1018 1290
rect 1054 1258 1086 1290
rect 1122 1258 1154 1290
rect 1190 1258 1222 1290
rect 1258 1258 1290 1290
<< poly >>
rect 188 746 388 760
rect 188 714 204 746
rect 236 714 272 746
rect 304 714 340 746
rect 372 714 388 746
rect 188 674 388 714
rect 188 234 388 274
rect 188 202 204 234
rect 236 202 272 234
rect 304 202 340 234
rect 372 202 388 234
rect 188 188 388 202
<< polycont >>
rect 204 714 236 746
rect 272 714 304 746
rect 340 714 372 746
rect 204 202 236 234
rect 272 202 304 234
rect 340 202 372 234
<< ppolyres >>
rect 188 274 388 674
<< pdiode >>
rect 164 1518 1160 1532
rect 164 1486 204 1518
rect 236 1486 272 1518
rect 304 1486 340 1518
rect 372 1486 408 1518
rect 440 1486 476 1518
rect 508 1486 544 1518
rect 576 1486 612 1518
rect 644 1486 680 1518
rect 712 1486 748 1518
rect 780 1486 816 1518
rect 848 1486 884 1518
rect 916 1486 952 1518
rect 984 1486 1020 1518
rect 1052 1486 1088 1518
rect 1120 1486 1160 1518
rect 164 1450 1160 1486
rect 164 1418 204 1450
rect 236 1418 272 1450
rect 304 1418 340 1450
rect 372 1418 408 1450
rect 440 1418 476 1450
rect 508 1418 544 1450
rect 576 1418 612 1450
rect 644 1418 680 1450
rect 712 1418 748 1450
rect 780 1418 816 1450
rect 848 1418 884 1450
rect 916 1418 952 1450
rect 984 1418 1020 1450
rect 1052 1418 1088 1450
rect 1120 1418 1160 1450
rect 164 1404 1160 1418
<< ndiode >>
rect 1032 762 1160 784
rect 1032 730 1046 762
rect 1078 730 1114 762
rect 1146 730 1160 762
rect 1032 694 1160 730
rect 1032 662 1046 694
rect 1078 662 1114 694
rect 1146 662 1160 694
rect 1032 626 1160 662
rect 1032 594 1046 626
rect 1078 594 1114 626
rect 1146 594 1160 626
rect 1032 558 1160 594
rect 1032 526 1046 558
rect 1078 526 1114 558
rect 1146 526 1160 558
rect 1032 490 1160 526
rect 1032 458 1046 490
rect 1078 458 1114 490
rect 1146 458 1160 490
rect 1032 422 1160 458
rect 1032 390 1046 422
rect 1078 390 1114 422
rect 1146 390 1160 422
rect 1032 354 1160 390
rect 1032 322 1046 354
rect 1078 322 1114 354
rect 1146 322 1160 354
rect 1032 286 1160 322
rect 1032 254 1046 286
rect 1078 254 1114 286
rect 1146 254 1160 286
rect 1032 218 1160 254
rect 1032 186 1046 218
rect 1078 186 1114 218
rect 1146 186 1160 218
rect 1032 164 1160 186
<< pdiodecont >>
rect 204 1486 236 1518
rect 272 1486 304 1518
rect 340 1486 372 1518
rect 408 1486 440 1518
rect 476 1486 508 1518
rect 544 1486 576 1518
rect 612 1486 644 1518
rect 680 1486 712 1518
rect 748 1486 780 1518
rect 816 1486 848 1518
rect 884 1486 916 1518
rect 952 1486 984 1518
rect 1020 1486 1052 1518
rect 1088 1486 1120 1518
rect 204 1418 236 1450
rect 272 1418 304 1450
rect 340 1418 372 1450
rect 408 1418 440 1450
rect 476 1418 508 1450
rect 544 1418 576 1450
rect 612 1418 644 1450
rect 680 1418 712 1450
rect 748 1418 780 1450
rect 816 1418 848 1450
rect 884 1418 916 1450
rect 952 1418 984 1450
rect 1020 1418 1052 1450
rect 1088 1418 1120 1450
<< ndiodecont >>
rect 1046 730 1078 762
rect 1114 730 1146 762
rect 1046 662 1078 694
rect 1114 662 1146 694
rect 1046 594 1078 626
rect 1114 594 1146 626
rect 1046 526 1078 558
rect 1114 526 1146 558
rect 1046 458 1078 490
rect 1114 458 1146 490
rect 1046 390 1078 422
rect 1114 390 1146 422
rect 1046 322 1078 354
rect 1114 322 1146 354
rect 1046 254 1078 286
rect 1114 254 1146 286
rect 1046 186 1078 218
rect 1114 186 1146 218
<< metal1 >>
rect 0 1678 1324 1696
rect 0 1646 34 1678
rect 66 1646 102 1678
rect 134 1646 170 1678
rect 202 1646 238 1678
rect 270 1646 306 1678
rect 338 1646 374 1678
rect 406 1646 442 1678
rect 474 1646 510 1678
rect 542 1646 578 1678
rect 610 1646 646 1678
rect 678 1646 714 1678
rect 746 1646 782 1678
rect 814 1646 850 1678
rect 882 1646 918 1678
rect 950 1646 986 1678
rect 1018 1646 1054 1678
rect 1086 1646 1122 1678
rect 1154 1646 1190 1678
rect 1222 1646 1258 1678
rect 1290 1646 1324 1678
rect 0 1628 1324 1646
rect 0 1586 68 1628
rect 0 1554 18 1586
rect 50 1554 68 1586
rect 0 1518 68 1554
rect 1256 1586 1324 1628
rect 1256 1554 1274 1586
rect 1306 1554 1324 1586
rect 0 1486 18 1518
rect 50 1486 68 1518
rect 0 1450 68 1486
rect 0 1418 18 1450
rect 50 1418 68 1450
rect 0 1382 68 1418
rect 204 1488 1120 1534
rect 204 1448 232 1488
rect 1092 1448 1120 1488
rect 204 1402 1120 1448
rect 1256 1518 1324 1554
rect 1256 1486 1274 1518
rect 1306 1486 1324 1518
rect 1256 1450 1324 1486
rect 1256 1418 1274 1450
rect 1306 1418 1324 1450
rect 0 1350 18 1382
rect 50 1350 68 1382
rect 0 1308 68 1350
rect 1256 1382 1324 1418
rect 1256 1350 1274 1382
rect 1306 1350 1324 1382
rect 1256 1308 1324 1350
rect 0 1290 1324 1308
rect 0 1258 34 1290
rect 66 1258 102 1290
rect 134 1258 170 1290
rect 202 1258 238 1290
rect 270 1258 306 1290
rect 338 1258 374 1290
rect 406 1258 442 1290
rect 474 1258 510 1290
rect 542 1258 578 1290
rect 610 1258 646 1290
rect 678 1258 714 1290
rect 746 1258 782 1290
rect 814 1258 850 1290
rect 882 1258 918 1290
rect 950 1258 986 1290
rect 1018 1258 1054 1290
rect 1086 1258 1122 1290
rect 1154 1258 1190 1290
rect 1222 1258 1258 1290
rect 1290 1258 1324 1290
rect 0 1240 1324 1258
rect 0 930 576 948
rect 0 898 34 930
rect 66 898 102 930
rect 134 898 170 930
rect 202 898 238 930
rect 270 898 306 930
rect 338 898 374 930
rect 406 898 442 930
rect 474 898 510 930
rect 542 898 576 930
rect 0 880 576 898
rect 0 830 68 880
rect 0 798 18 830
rect 50 798 68 830
rect 0 762 68 798
rect 508 830 576 880
rect 508 798 526 830
rect 558 798 576 830
rect 508 762 576 798
rect 0 730 18 762
rect 50 730 68 762
rect 0 694 68 730
rect 204 747 372 762
rect 204 746 227 747
rect 349 746 372 747
rect 204 707 227 714
rect 349 707 372 714
rect 204 698 372 707
rect 508 730 526 762
rect 558 730 576 762
rect 0 662 18 694
rect 50 662 68 694
rect 0 626 68 662
rect 0 594 18 626
rect 50 594 68 626
rect 0 558 68 594
rect 0 526 18 558
rect 50 526 68 558
rect 0 490 68 526
rect 0 458 18 490
rect 50 458 68 490
rect 0 422 68 458
rect 0 390 18 422
rect 50 390 68 422
rect 0 354 68 390
rect 0 322 18 354
rect 50 322 68 354
rect 0 286 68 322
rect 0 254 18 286
rect 50 254 68 286
rect 0 218 68 254
rect 508 694 576 730
rect 508 662 526 694
rect 558 662 576 694
rect 508 626 576 662
rect 508 594 526 626
rect 558 594 576 626
rect 508 558 576 594
rect 508 526 526 558
rect 558 526 576 558
rect 508 490 576 526
rect 508 458 526 490
rect 558 458 576 490
rect 508 422 576 458
rect 508 390 526 422
rect 558 390 576 422
rect 508 354 576 390
rect 508 322 526 354
rect 558 322 576 354
rect 508 297 576 322
rect 508 286 535 297
rect 508 254 526 286
rect 0 186 18 218
rect 50 186 68 218
rect 204 241 372 250
rect 204 234 227 241
rect 349 234 372 241
rect 204 201 227 202
rect 349 201 372 202
rect 204 186 372 201
rect 508 218 535 254
rect 508 186 526 218
rect 0 150 68 186
rect 0 118 18 150
rect 50 118 68 150
rect 0 68 68 118
rect 508 150 535 186
rect 508 118 526 150
rect 508 93 535 118
rect 575 93 576 297
rect 508 68 576 93
rect 0 50 576 68
rect 0 18 34 50
rect 66 18 102 50
rect 134 18 170 50
rect 202 18 238 50
rect 270 18 306 50
rect 338 18 374 50
rect 406 18 442 50
rect 474 18 510 50
rect 542 18 576 50
rect 0 0 576 18
rect 868 930 1324 948
rect 868 898 910 930
rect 942 898 978 930
rect 1010 898 1046 930
rect 1078 898 1114 930
rect 1146 898 1182 930
rect 1214 898 1250 930
rect 1282 898 1324 930
rect 868 880 1324 898
rect 868 830 936 880
rect 868 798 886 830
rect 918 798 936 830
rect 868 762 936 798
rect 1256 830 1324 880
rect 1256 798 1274 830
rect 1306 798 1324 830
rect 868 730 886 762
rect 918 730 936 762
rect 868 694 936 730
rect 868 662 886 694
rect 918 662 936 694
rect 868 626 936 662
rect 868 594 886 626
rect 918 594 936 626
rect 868 558 936 594
rect 868 526 886 558
rect 918 526 936 558
rect 868 490 936 526
rect 868 458 886 490
rect 918 458 936 490
rect 868 422 936 458
rect 868 390 886 422
rect 918 390 936 422
rect 868 354 936 390
rect 868 322 886 354
rect 918 322 936 354
rect 868 297 936 322
rect 868 93 869 297
rect 909 286 936 297
rect 918 254 936 286
rect 909 218 936 254
rect 918 186 936 218
rect 909 150 936 186
rect 1046 740 1146 778
rect 1046 208 1076 740
rect 1116 208 1146 740
rect 1046 170 1146 208
rect 1256 762 1324 798
rect 1256 730 1274 762
rect 1306 730 1324 762
rect 1256 694 1324 730
rect 1256 662 1274 694
rect 1306 662 1324 694
rect 1256 626 1324 662
rect 1256 594 1274 626
rect 1306 594 1324 626
rect 1256 558 1324 594
rect 1256 526 1274 558
rect 1306 526 1324 558
rect 1256 490 1324 526
rect 1256 458 1274 490
rect 1306 458 1324 490
rect 1256 422 1324 458
rect 1256 390 1274 422
rect 1306 390 1324 422
rect 1256 354 1324 390
rect 1256 322 1274 354
rect 1306 322 1324 354
rect 1256 286 1324 322
rect 1256 254 1274 286
rect 1306 254 1324 286
rect 1256 218 1324 254
rect 1256 186 1274 218
rect 1306 186 1324 218
rect 918 118 936 150
rect 909 93 936 118
rect 868 68 936 93
rect 1256 150 1324 186
rect 1256 118 1274 150
rect 1306 118 1324 150
rect 1256 68 1324 118
rect 868 50 1324 68
rect 868 18 910 50
rect 942 18 978 50
rect 1010 18 1046 50
rect 1078 18 1114 50
rect 1146 18 1182 50
rect 1214 18 1250 50
rect 1282 18 1324 50
rect 868 0 1324 18
<< via1 >>
rect 232 1448 1092 1488
rect 227 746 349 747
rect 227 714 236 746
rect 236 714 272 746
rect 272 714 304 746
rect 304 714 340 746
rect 340 714 349 746
rect 227 707 349 714
rect 535 286 575 297
rect 535 254 558 286
rect 558 254 575 286
rect 227 234 349 241
rect 227 202 236 234
rect 236 202 272 234
rect 272 202 304 234
rect 304 202 340 234
rect 340 202 349 234
rect 227 201 349 202
rect 535 218 575 254
rect 535 186 558 218
rect 558 186 575 218
rect 535 150 575 186
rect 535 118 558 150
rect 558 118 575 150
rect 535 93 575 118
rect 869 286 909 297
rect 869 254 886 286
rect 886 254 909 286
rect 869 218 909 254
rect 869 186 886 218
rect 886 186 909 218
rect 869 150 909 186
rect 1076 208 1116 740
rect 869 118 886 150
rect 886 118 909 150
rect 869 93 909 118
<< metal2 >>
rect 204 1488 1120 1696
rect 204 1448 232 1488
rect 1092 1448 1120 1488
rect 204 1402 1120 1448
rect 204 778 372 1402
rect 204 747 1146 778
rect 204 707 227 747
rect 349 740 1146 747
rect 349 707 1076 740
rect 204 698 1076 707
rect 535 297 909 306
rect 204 241 372 250
rect 204 201 227 241
rect 349 201 372 241
rect 204 0 372 201
rect 575 93 869 297
rect 1046 208 1076 698
rect 1116 208 1146 740
rect 1046 170 1146 208
rect 535 84 909 93
<< labels >>
rlabel comment s 902 34 902 34 4 sub!
rlabel comment s 34 34 34 34 4 sub!
rlabel comment s 662 1468 662 1468 4 dpant
rlabel comment s 288 474 288 474 4 rppd r=793.834
rlabel comment s 1096 474 1096 474 4 dant
flabel metal1 s 0 1628 1324 1696 0 FreeSans 800 0 0 0 iovdd
port 1 nsew
flabel metal2 s 535 84 909 306 0 FreeSans 800 0 0 0 iovss
port 2 nsew
rlabel metal2 s 204 1402 1120 1696 4 core
port 4 nsew
rlabel metal2 s 204 0 372 250 4 pad
port 3 nsew
<< properties >>
string device primitive
string GDS_END 17350994
string GDS_FILE sg13g2_io.gds
string GDS_START 17335126
<< end >>
