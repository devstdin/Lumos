magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< nwell >>
rect -23 149 17525 199
<< poly >>
rect -1600 -243 -1550 -201
<< metal1 >>
rect -1948 13357 17939 14105
rect -1948 13355 855 13357
rect -1948 1715 -813 13214
rect -678 12981 -386 13033
rect -678 1855 -586 1921
rect -678 1798 -668 1855
rect -596 1798 -586 1855
rect -678 1788 -586 1798
rect -478 1855 -386 1921
rect -478 1798 -468 1855
rect -396 1798 -386 1855
rect -478 1788 -386 1798
rect -230 1715 -25 13213
rect 105 13179 291 13355
rect 369 13211 3341 13263
rect 105 11207 343 13179
rect 105 10995 291 11207
rect 1755 11175 1955 13211
rect 3553 13179 3739 13357
rect 3817 13211 6789 13263
rect 3367 11207 3499 13179
rect 369 11027 3341 11175
rect 105 9023 343 10995
rect 105 8811 291 9023
rect 1755 8991 1955 11027
rect 3419 10995 3499 11207
rect 3367 9023 3499 10995
rect 369 8843 3341 8991
rect 105 6839 343 8811
rect 105 6627 291 6839
rect 1755 6807 1955 8843
rect 3419 8811 3499 9023
rect 3367 6839 3499 8811
rect 369 6659 3341 6807
rect 105 4655 343 6627
rect 105 4443 291 4655
rect 1755 4623 1955 6659
rect 3419 6627 3499 6839
rect 3367 4655 3499 6627
rect 369 4475 3341 4623
rect 105 2471 343 4443
rect 105 2259 291 2471
rect 1755 2439 1955 4475
rect 3419 4443 3499 4655
rect 3367 2471 3499 4443
rect 369 2291 3341 2439
rect 105 1865 343 2259
rect 18 1855 343 1865
rect 18 1798 28 1855
rect 91 1798 343 1855
rect 18 1788 343 1798
rect -1948 1574 -25 1715
rect -1948 162 -1684 1574
rect -1625 365 -1505 375
rect -1625 281 -1615 365
rect -1515 281 -1505 365
rect -1625 271 -1505 281
rect -230 162 -25 1574
rect 105 287 343 1788
rect 1755 255 1955 2291
rect 3419 2259 3499 2471
rect 3367 287 3499 2259
rect 3553 11207 3791 13179
rect 3553 10995 3739 11207
rect 5203 11175 5403 13211
rect 7001 13179 7187 13357
rect 7265 13211 10237 13263
rect 6815 11207 6947 13179
rect 3817 11027 6789 11175
rect 3553 9023 3791 10995
rect 3553 8811 3739 9023
rect 5203 8991 5403 11027
rect 6867 10995 6947 11207
rect 6815 9023 6947 10995
rect 3817 8843 6789 8991
rect 3553 6839 3791 8811
rect 3553 6627 3739 6839
rect 5203 6807 5403 8843
rect 6867 8811 6947 9023
rect 6815 6839 6947 8811
rect 3817 6659 6789 6807
rect 3553 4655 3791 6627
rect 3553 4443 3739 4655
rect 5203 4623 5403 6659
rect 6867 6627 6947 6839
rect 6815 4655 6947 6627
rect 3817 4475 6789 4623
rect 3553 2471 3791 4443
rect 3553 2259 3739 2471
rect 5203 2439 5403 4475
rect 6867 4443 6947 4655
rect 6815 2471 6947 4443
rect 3817 2291 6789 2439
rect 3553 287 3791 2259
rect 369 203 3341 255
rect -1948 119 -25 162
rect 1755 138 1955 203
rect -1948 14 673 119
rect -1948 -456 -1669 14
rect -1526 -110 446 -108
rect -1526 -150 -668 -110
rect -596 -150 446 -110
rect -1526 -160 446 -150
rect -1610 -196 -1558 -186
rect -1610 -201 -1540 -196
rect -1610 -243 -1600 -201
rect -1550 -206 -1540 -201
rect 488 -206 530 -176
rect -1550 -238 530 -206
rect -1550 -243 -1540 -238
rect -1610 -248 -1540 -243
rect -1610 -258 -1558 -248
rect 488 -268 530 -238
rect -1526 -456 446 -284
rect -1948 -457 446 -456
rect 586 -369 673 14
rect 1755 -16 1765 138
rect 1945 -16 1955 138
rect 1755 -26 1955 -16
rect 3419 -111 3499 287
rect 5203 255 5403 2291
rect 6867 2259 6947 2471
rect 6815 287 6947 2259
rect 7001 11207 7239 13179
rect 7001 10995 7187 11207
rect 8651 11175 8851 13211
rect 10449 13179 10635 13357
rect 10713 13211 13685 13263
rect 10263 11207 10395 13179
rect 7265 11027 10237 11175
rect 7001 9023 7239 10995
rect 7001 8811 7187 9023
rect 8651 8991 8851 11027
rect 10315 10995 10395 11207
rect 10263 9023 10395 10995
rect 7265 8843 10237 8991
rect 7001 6839 7239 8811
rect 7001 6627 7187 6839
rect 8651 6807 8851 8843
rect 10315 8811 10395 9023
rect 10263 6839 10395 8811
rect 7265 6659 10237 6807
rect 7001 4655 7239 6627
rect 7001 4443 7187 4655
rect 8651 4623 8851 6659
rect 10315 6627 10395 6839
rect 10263 4655 10395 6627
rect 7265 4475 10237 4623
rect 7001 2471 7239 4443
rect 7001 2259 7187 2471
rect 8651 2439 8851 4475
rect 10315 4443 10395 4655
rect 10263 2471 10395 4443
rect 7265 2291 10237 2439
rect 7001 287 7239 2259
rect 3817 203 6789 255
rect 5203 138 5403 203
rect 5203 -16 5213 138
rect 5393 -16 5403 138
rect 5203 -26 5403 -16
rect 6867 148 6947 287
rect 8651 255 8851 2291
rect 10315 2259 10395 2471
rect 10263 287 10395 2259
rect 10449 11207 10687 13179
rect 10449 10995 10635 11207
rect 12099 11175 12299 13211
rect 13897 13179 14083 13357
rect 14161 13211 17133 13263
rect 13711 11207 13843 13179
rect 10713 11027 13685 11175
rect 10449 9023 10687 10995
rect 10449 8811 10635 9023
rect 12099 8991 12299 11027
rect 13763 10995 13843 11207
rect 13711 9023 13843 10995
rect 10713 8843 13685 8991
rect 10449 6839 10687 8811
rect 10449 6627 10635 6839
rect 12099 6807 12299 8843
rect 13763 8811 13843 9023
rect 13711 6839 13843 8811
rect 10713 6659 13685 6807
rect 10449 4655 10687 6627
rect 10449 4443 10635 4655
rect 12099 4623 12299 6659
rect 13763 6627 13843 6839
rect 13711 4655 13843 6627
rect 10713 4475 13685 4623
rect 10449 2471 10687 4443
rect 10449 2259 10635 2471
rect 12099 2439 12299 4475
rect 13763 4443 13843 4655
rect 13711 2471 13843 4443
rect 10713 2291 13685 2439
rect 10449 287 10687 2259
rect 7265 203 10237 255
rect 6867 138 7054 148
rect 6867 -16 6877 138
rect 7044 -16 7054 138
rect 6867 -26 7054 -16
rect 8651 138 8851 203
rect 8651 -16 8661 138
rect 8841 -16 8851 138
rect 10315 111 10395 287
rect 12099 255 12299 2291
rect 13763 2259 13843 2471
rect 13711 287 13843 2259
rect 13897 11207 14135 13179
rect 13897 10995 14083 11207
rect 15547 11175 15747 13211
rect 17159 11207 17291 13179
rect 14161 11027 17133 11175
rect 13897 9023 14135 10995
rect 13897 8811 14083 9023
rect 15547 8991 15747 11027
rect 17211 10995 17291 11207
rect 17159 9023 17291 10995
rect 14161 8843 17133 8991
rect 13897 6839 14135 8811
rect 13897 6627 14083 6839
rect 15547 6807 15747 8843
rect 17211 8811 17291 9023
rect 17159 6839 17291 8811
rect 14161 6659 17133 6807
rect 13897 4655 14135 6627
rect 13897 4443 14083 4655
rect 15547 4623 15747 6659
rect 17211 6627 17291 6839
rect 17159 4655 17291 6627
rect 14161 4475 17133 4623
rect 13897 2471 14135 4443
rect 13897 2259 14083 2471
rect 15547 2439 15747 4475
rect 17211 4443 17291 4655
rect 17159 2471 17291 4443
rect 14161 2291 17133 2439
rect 13897 287 14135 2259
rect 10713 203 13685 255
rect 8651 -26 8851 -16
rect 10069 101 10395 111
rect 10069 -73 10079 101
rect 10259 -73 10395 101
rect 12099 138 12299 203
rect 12099 -16 12109 138
rect 12289 -16 12299 138
rect 12099 -26 12299 -16
rect 13763 148 13843 287
rect 15547 255 15747 2291
rect 17211 2259 17291 2471
rect 17159 287 17291 2259
rect 17366 327 17939 13357
rect 14161 203 17133 255
rect 13763 138 13950 148
rect 13763 -16 13773 138
rect 13940 -16 13950 138
rect 13763 -26 13950 -16
rect 15547 138 15747 203
rect 15547 -16 15557 138
rect 15737 -16 15747 138
rect 15547 -26 15747 -16
rect 17211 149 17291 287
rect 10069 -83 10395 -73
rect 1845 -121 4351 -111
rect 17211 -120 17398 149
rect 1845 -238 1855 -121
rect 1959 -238 4161 -121
rect 4341 -238 4351 -121
rect 1845 -248 4351 -238
rect 586 -439 6489 -369
rect 586 -457 2359 -439
rect -1948 -773 2359 -457
rect 4151 -491 4351 -481
rect 4151 -541 4161 -491
rect 2665 -583 4161 -541
rect 4341 -541 4351 -491
rect 5915 -492 6034 -481
rect 4341 -583 5837 -541
rect 2665 -593 5837 -583
rect 5915 -589 5925 -492
rect 6024 -589 6034 -492
rect -1948 -994 -1483 -773
rect 1845 -852 1969 -842
rect -1405 -962 1767 -910
rect 1845 -950 1855 -852
rect 1959 -950 1969 -852
rect -1948 -1966 -1431 -994
rect -1948 -2178 -1483 -1966
rect 81 -1998 281 -962
rect 1845 -994 1969 -950
rect 1793 -1966 1969 -994
rect -1405 -2050 1767 -1998
rect 81 -2094 281 -2050
rect -1405 -2146 1767 -2094
rect -1948 -3150 -1431 -2178
rect -1948 -3362 -1483 -3150
rect 81 -3182 281 -2146
rect 1845 -2178 1969 -1966
rect 1793 -3150 1969 -2178
rect -1405 -3234 1767 -3182
rect 81 -3278 281 -3234
rect -1405 -3330 1767 -3278
rect -1948 -4334 -1431 -3362
rect -1948 -4546 -1483 -4334
rect 81 -4366 281 -3330
rect 1845 -3362 1969 -3150
rect 1793 -4334 1969 -3362
rect -1405 -4418 1767 -4366
rect 81 -4462 281 -4418
rect -1405 -4514 1767 -4462
rect -1948 -5518 -1431 -4546
rect -1948 -5730 -1483 -5518
rect 81 -5550 281 -4514
rect 1845 -4546 1969 -4334
rect 1793 -5518 1969 -4546
rect -1405 -5602 1767 -5550
rect 81 -5646 281 -5602
rect -1405 -5698 1767 -5646
rect -1948 -6702 -1431 -5730
rect -1948 -6914 -1483 -6702
rect 81 -6734 281 -5698
rect 1845 -5730 1969 -5518
rect 1793 -6702 1969 -5730
rect -1405 -6786 1767 -6734
rect 81 -6830 281 -6786
rect -1405 -6882 1767 -6830
rect -1948 -7886 -1431 -6914
rect -1948 -8098 -1483 -7886
rect 81 -7918 281 -6882
rect 1845 -6914 1969 -6702
rect 1793 -7886 1969 -6914
rect -1405 -7970 1767 -7918
rect 81 -8014 281 -7970
rect -1405 -8066 1767 -8014
rect -1948 -9070 -1431 -8098
rect -1948 -9282 -1483 -9070
rect 81 -9102 281 -8066
rect 1845 -8098 1969 -7886
rect 1793 -9070 1969 -8098
rect -1405 -9154 1767 -9102
rect 81 -9198 281 -9154
rect -1405 -9250 1767 -9198
rect -1948 -10254 -1431 -9282
rect -1948 -10466 -1483 -10254
rect 81 -10286 281 -9250
rect 1845 -9282 1969 -9070
rect 1793 -10254 1969 -9282
rect -1405 -10338 1767 -10286
rect 81 -10382 281 -10338
rect -1405 -10434 1767 -10382
rect -1948 -11438 -1431 -10466
rect -1948 -11650 -1483 -11438
rect 81 -11470 281 -10434
rect 1845 -10466 1969 -10254
rect 1793 -11438 1969 -10466
rect -1405 -11522 1767 -11470
rect 81 -11566 281 -11522
rect -1405 -11618 1767 -11566
rect -1948 -12622 -1431 -11650
rect -1948 -12834 -1483 -12622
rect 81 -12654 281 -11618
rect 1845 -11650 1969 -11438
rect 1793 -12622 1969 -11650
rect -1405 -12706 1767 -12654
rect 81 -12750 281 -12706
rect -1405 -12802 1767 -12750
rect -1948 -13806 -1431 -12834
rect -1948 -14018 -1483 -13806
rect 81 -13838 281 -12802
rect 1845 -12834 1969 -12622
rect 1793 -13806 1969 -12834
rect -1405 -13890 1767 -13838
rect 81 -13934 281 -13890
rect -1405 -13986 1767 -13934
rect -1948 -14990 -1431 -14018
rect -1948 -15202 -1483 -14990
rect 81 -15022 281 -13986
rect 1845 -14018 1969 -13806
rect 1793 -14990 1969 -14018
rect -1405 -15074 1767 -15022
rect 81 -15118 281 -15074
rect -1405 -15170 1767 -15118
rect -1948 -16174 -1431 -15202
rect -1948 -16388 -1684 -16174
rect 81 -16204 281 -15170
rect 1845 -15202 1969 -14990
rect 1793 -16174 1969 -15202
rect 81 -16206 91 -16204
rect -1405 -16258 91 -16206
rect 81 -16326 91 -16258
rect 271 -16206 281 -16204
rect 271 -16258 1767 -16206
rect 271 -16326 281 -16258
rect 81 -16336 281 -16326
rect 2050 -16388 2359 -773
rect 2477 -1597 2639 -625
rect 2477 -1809 2587 -1597
rect 4151 -1629 4351 -593
rect 5915 -625 6034 -589
rect 5863 -1597 6034 -625
rect 2665 -1777 5837 -1629
rect 2477 -2781 2639 -1809
rect 2477 -2993 2587 -2781
rect 4151 -2813 4351 -1777
rect 5915 -1809 6034 -1597
rect 5863 -2781 6034 -1809
rect 2665 -2961 5837 -2813
rect 2477 -3965 2639 -2993
rect 2477 -4177 2587 -3965
rect 4151 -3997 4351 -2961
rect 5915 -2993 6034 -2781
rect 5863 -3965 6034 -2993
rect 2665 -4145 5837 -3997
rect 2477 -5149 2639 -4177
rect 2477 -5361 2587 -5149
rect 4151 -5181 4351 -4145
rect 5915 -4177 6034 -3965
rect 5863 -5149 6034 -4177
rect 2665 -5329 5837 -5181
rect 2477 -6333 2639 -5361
rect 2477 -6545 2587 -6333
rect 4151 -6365 4351 -5329
rect 5915 -5361 6034 -5149
rect 5863 -6333 6034 -5361
rect 2665 -6513 5837 -6365
rect 2477 -7517 2639 -6545
rect 2477 -7729 2587 -7517
rect 4151 -7549 4351 -6513
rect 5915 -6545 6034 -6333
rect 5863 -7517 6034 -6545
rect 2665 -7697 5837 -7549
rect 2477 -8701 2639 -7729
rect 2477 -8913 2587 -8701
rect 4151 -8733 4351 -7697
rect 5915 -7729 6034 -7517
rect 5863 -8701 6034 -7729
rect 2665 -8881 5837 -8733
rect 2477 -9885 2639 -8913
rect 2477 -10097 2587 -9885
rect 4151 -9917 4351 -8881
rect 5915 -8913 6034 -8701
rect 5863 -9885 6034 -8913
rect 2665 -10065 5837 -9917
rect 2477 -11069 2639 -10097
rect 2477 -11281 2587 -11069
rect 4151 -11101 4351 -10065
rect 5915 -10097 6034 -9885
rect 5863 -11069 6034 -10097
rect 2665 -11249 5837 -11101
rect 2477 -12253 2639 -11281
rect 2477 -12465 2587 -12253
rect 4151 -12285 4351 -11249
rect 5915 -11281 6034 -11069
rect 5863 -12253 6034 -11281
rect 2665 -12433 5837 -12285
rect 2477 -13437 2639 -12465
rect 2477 -13649 2587 -13437
rect 4151 -13469 4351 -12433
rect 5915 -12465 6034 -12253
rect 5863 -13437 6034 -12465
rect 2665 -13617 5837 -13469
rect 2477 -14621 2639 -13649
rect 2477 -14833 2587 -14621
rect 4151 -14653 4351 -13617
rect 5915 -13649 6034 -13437
rect 5863 -14621 6034 -13649
rect 2665 -14801 5837 -14653
rect 2477 -15805 2639 -14833
rect 2477 -15829 2589 -15805
rect 2477 -15940 2487 -15829
rect 2579 -15940 2589 -15829
rect 4151 -15837 4351 -14801
rect 5915 -14833 6034 -14621
rect 5863 -15805 6034 -14833
rect 2665 -15889 5837 -15837
rect 2477 -15948 2589 -15940
rect 2477 -16158 3023 -16148
rect 2477 -16305 2487 -16158
rect 2579 -16305 3023 -16158
rect 2477 -16315 3023 -16305
rect 5483 -16317 5712 -16150
rect 5592 -16388 5712 -16317
rect 6132 -16388 6489 -439
rect 6711 -469 16789 -201
rect 6711 -2811 7036 -469
rect 7355 -621 7727 -569
rect 8051 -621 8423 -569
rect 8747 -621 9119 -569
rect 9443 -621 9815 -569
rect 10803 -621 11175 -569
rect 11499 -621 11871 -569
rect 12195 -621 12567 -569
rect 12891 -621 13263 -569
rect 14251 -621 14623 -569
rect 14947 -621 15319 -569
rect 15643 -621 16015 -569
rect 16339 -621 16711 -569
rect 7225 -1006 7329 -653
rect 7225 -1186 7235 -1006
rect 7319 -1186 7329 -1006
rect 7225 -2625 7329 -1186
rect 7491 -1549 7591 -621
rect 7491 -1729 7501 -1549
rect 7582 -1729 7591 -1549
rect 7491 -2657 7591 -1729
rect 7753 -2092 7857 -653
rect 7753 -2272 7763 -2092
rect 7847 -2272 7857 -2092
rect 7753 -2625 7857 -2272
rect 7921 -1006 8025 -653
rect 7921 -1186 7931 -1006
rect 8015 -1186 8025 -1006
rect 7921 -2625 8025 -1186
rect 8187 -1549 8287 -621
rect 8187 -1729 8197 -1549
rect 8277 -1729 8287 -1549
rect 8187 -2657 8287 -1729
rect 8449 -2092 8553 -653
rect 8449 -2272 8459 -2092
rect 8543 -2272 8553 -2092
rect 8449 -2625 8553 -2272
rect 8617 -1006 8721 -653
rect 8617 -1186 8627 -1006
rect 8711 -1186 8721 -1006
rect 8617 -2625 8721 -1186
rect 8883 -1549 8983 -621
rect 8883 -1729 8893 -1549
rect 8973 -1729 8983 -1549
rect 8883 -2657 8983 -1729
rect 9145 -2092 9249 -653
rect 9145 -2272 9155 -2092
rect 9239 -2272 9249 -2092
rect 9145 -2625 9249 -2272
rect 9313 -1006 9417 -653
rect 9313 -1186 9323 -1006
rect 9407 -1186 9417 -1006
rect 9313 -2625 9417 -1186
rect 9579 -1549 9679 -621
rect 9579 -1729 9589 -1549
rect 9669 -1729 9679 -1549
rect 9579 -2657 9679 -1729
rect 9841 -2092 9945 -653
rect 9841 -2272 9851 -2092
rect 9935 -2272 9945 -2092
rect 9841 -2625 9945 -2272
rect 10673 -1006 10777 -653
rect 10673 -1186 10683 -1006
rect 10767 -1186 10777 -1006
rect 10673 -2625 10777 -1186
rect 10939 -1549 11039 -621
rect 10939 -1729 10949 -1549
rect 11030 -1729 11039 -1549
rect 10939 -2657 11039 -1729
rect 11201 -2092 11305 -653
rect 11201 -2272 11211 -2092
rect 11295 -2272 11305 -2092
rect 11201 -2625 11305 -2272
rect 11369 -1006 11473 -653
rect 11369 -1186 11379 -1006
rect 11463 -1186 11473 -1006
rect 11369 -2625 11473 -1186
rect 11635 -1549 11735 -621
rect 11635 -1729 11645 -1549
rect 11726 -1729 11735 -1549
rect 11635 -2657 11735 -1729
rect 11897 -2092 12001 -653
rect 11897 -2272 11907 -2092
rect 11991 -2272 12001 -2092
rect 11897 -2625 12001 -2272
rect 12065 -1006 12169 -653
rect 12065 -1186 12075 -1006
rect 12159 -1186 12169 -1006
rect 12065 -2625 12169 -1186
rect 12331 -1549 12431 -621
rect 12331 -1729 12341 -1549
rect 12422 -1729 12431 -1549
rect 12331 -2657 12431 -1729
rect 12593 -2092 12697 -653
rect 12593 -2272 12603 -2092
rect 12687 -2272 12697 -2092
rect 12593 -2625 12697 -2272
rect 12761 -1006 12865 -653
rect 12761 -1186 12771 -1006
rect 12855 -1186 12865 -1006
rect 12761 -2625 12865 -1186
rect 13027 -1549 13127 -621
rect 13027 -1729 13037 -1549
rect 13118 -1729 13127 -1549
rect 13027 -2657 13127 -1729
rect 13289 -2092 13393 -653
rect 13289 -2272 13299 -2092
rect 13383 -2272 13393 -2092
rect 13289 -2625 13393 -2272
rect 14121 -1006 14225 -653
rect 14121 -1186 14131 -1006
rect 14215 -1186 14225 -1006
rect 14121 -2625 14225 -1186
rect 14387 -1549 14487 -621
rect 14387 -1729 14397 -1549
rect 14478 -1729 14487 -1549
rect 14387 -2657 14487 -1729
rect 14649 -2092 14753 -653
rect 14649 -2272 14659 -2092
rect 14743 -2272 14753 -2092
rect 14649 -2625 14753 -2272
rect 14817 -1006 14921 -653
rect 14817 -1186 14827 -1006
rect 14911 -1186 14921 -1006
rect 14817 -2625 14921 -1186
rect 15083 -1549 15183 -621
rect 15083 -1729 15093 -1549
rect 15174 -1729 15183 -1549
rect 15083 -2657 15183 -1729
rect 15345 -2092 15449 -653
rect 15345 -2272 15355 -2092
rect 15439 -2272 15449 -2092
rect 15345 -2625 15449 -2272
rect 15513 -1006 15617 -653
rect 15513 -1186 15523 -1006
rect 15607 -1186 15617 -1006
rect 15513 -2625 15617 -1186
rect 15779 -1549 15879 -621
rect 15779 -1729 15789 -1549
rect 15870 -1729 15879 -1549
rect 15779 -2657 15879 -1729
rect 16041 -2092 16145 -653
rect 16041 -2272 16051 -2092
rect 16135 -2272 16145 -2092
rect 16041 -2625 16145 -2272
rect 16209 -1006 16313 -653
rect 16209 -1186 16219 -1006
rect 16303 -1186 16313 -1006
rect 16209 -2625 16313 -1186
rect 16475 -1549 16575 -621
rect 17049 -637 17939 -120
rect 16475 -1729 16485 -1549
rect 16566 -1729 16575 -1549
rect 16475 -2657 16575 -1729
rect 16737 -2092 16841 -653
rect 16737 -2272 16747 -2092
rect 16831 -2272 16841 -2092
rect 16737 -2625 16841 -2272
rect 7355 -2709 7727 -2657
rect 8051 -2709 8423 -2657
rect 8747 -2709 9119 -2657
rect 9443 -2709 9815 -2657
rect 10803 -2709 11175 -2657
rect 11499 -2709 11871 -2657
rect 12195 -2709 12567 -2657
rect 12891 -2709 13263 -2657
rect 14251 -2709 14623 -2657
rect 14947 -2709 15319 -2657
rect 15643 -2709 16015 -2657
rect 16339 -2709 16711 -2657
rect 6711 -3152 9893 -2811
rect 10069 -2998 10398 -2988
rect 10069 -3142 10079 -2998
rect 10259 -3142 10398 -2998
rect 10069 -3152 10398 -3142
rect 6711 -3308 7187 -3152
rect 7265 -3276 10237 -3224
rect 6711 -5280 7239 -3308
rect 8651 -4204 8851 -3276
rect 10315 -3308 10398 -3152
rect 8651 -4384 8661 -4204
rect 8841 -4384 8851 -4204
rect 6711 -5492 7187 -5280
rect 8651 -5312 8851 -4384
rect 10263 -4204 10398 -3308
rect 10263 -4384 10283 -4204
rect 10388 -4384 10398 -4204
rect 10263 -5280 10398 -4384
rect 7265 -5460 10237 -5312
rect 6711 -7464 7239 -5492
rect 6711 -7676 7187 -7464
rect 8651 -7496 8851 -5460
rect 10315 -5492 10398 -5280
rect 10263 -7464 10398 -5492
rect 7265 -7644 10237 -7496
rect 6711 -9648 7239 -7676
rect 6711 -9860 7187 -9648
rect 8651 -9680 8851 -7644
rect 10315 -7676 10398 -7464
rect 10263 -9648 10398 -7676
rect 7265 -9828 10237 -9680
rect 6711 -11832 7239 -9860
rect 6711 -12044 7187 -11832
rect 8651 -11864 8851 -9828
rect 10315 -9860 10398 -9648
rect 10263 -11832 10398 -9860
rect 7265 -12012 10237 -11864
rect 6711 -14016 7239 -12044
rect 6711 -14228 7187 -14016
rect 8651 -14048 8851 -12012
rect 10315 -12044 10398 -11832
rect 10263 -14016 10398 -12044
rect 7265 -14196 10237 -14048
rect 6711 -16200 7239 -14228
rect 6711 -16388 7183 -16200
rect 8651 -16232 8851 -14196
rect 10315 -14228 10398 -14016
rect 10263 -16200 10398 -14228
rect 10449 -3152 13341 -2810
rect 13517 -2998 13846 -2988
rect 13517 -3142 13527 -2998
rect 13707 -3142 13846 -2998
rect 13517 -3152 13846 -3142
rect 10449 -3308 10635 -3152
rect 10713 -3276 13685 -3224
rect 10449 -5280 10687 -3308
rect 12099 -4204 12299 -3276
rect 13763 -3308 13846 -3152
rect 12099 -4384 12109 -4204
rect 12289 -4384 12299 -4204
rect 10449 -5492 10635 -5280
rect 12099 -5312 12299 -4384
rect 13711 -5280 13846 -3308
rect 10713 -5460 13685 -5312
rect 10449 -7464 10687 -5492
rect 10449 -7676 10635 -7464
rect 12099 -7496 12299 -5460
rect 13763 -5492 13846 -5280
rect 13711 -7464 13846 -5492
rect 10713 -7644 13685 -7496
rect 10449 -9648 10687 -7676
rect 10449 -9860 10635 -9648
rect 12099 -9680 12299 -7644
rect 13763 -7676 13846 -7464
rect 13711 -9648 13846 -7676
rect 10713 -9828 13685 -9680
rect 10449 -11832 10687 -9860
rect 10449 -12044 10635 -11832
rect 12099 -11864 12299 -9828
rect 13763 -9860 13846 -9648
rect 13711 -11832 13846 -9860
rect 10713 -12012 13685 -11864
rect 10449 -14016 10687 -12044
rect 10449 -14228 10635 -14016
rect 12099 -14048 12299 -12012
rect 13763 -12044 13846 -11832
rect 13711 -14016 13846 -12044
rect 10713 -14196 13685 -14048
rect 10449 -16200 10687 -14228
rect 7265 -16284 10237 -16232
rect 10449 -16388 10631 -16200
rect 12099 -16232 12299 -14196
rect 13763 -14228 13846 -14016
rect 13711 -16200 13846 -14228
rect 13897 -3152 16789 -2812
rect 16965 -2998 17294 -2988
rect 16965 -3142 16975 -2998
rect 17155 -3142 17294 -2998
rect 16965 -3152 17294 -3142
rect 13897 -3308 14083 -3152
rect 14161 -3276 17133 -3224
rect 13897 -5280 14135 -3308
rect 15547 -4204 15747 -3276
rect 17211 -3308 17294 -3152
rect 15547 -4384 15557 -4204
rect 15737 -4384 15747 -4204
rect 13897 -5492 14083 -5280
rect 15547 -5312 15747 -4384
rect 17159 -5280 17294 -3308
rect 14161 -5460 17133 -5312
rect 13897 -7464 14135 -5492
rect 13897 -7676 14083 -7464
rect 15547 -7496 15747 -5460
rect 17211 -5492 17294 -5280
rect 17159 -7464 17294 -5492
rect 14161 -7644 17133 -7496
rect 13897 -9648 14135 -7676
rect 13897 -9860 14083 -9648
rect 15547 -9680 15747 -7644
rect 17211 -7676 17294 -7464
rect 17159 -9648 17294 -7676
rect 14161 -9828 17133 -9680
rect 13897 -11832 14135 -9860
rect 13897 -12044 14083 -11832
rect 15547 -11864 15747 -9828
rect 17211 -9860 17294 -9648
rect 17159 -11832 17294 -9860
rect 14161 -12012 17133 -11864
rect 13897 -14016 14135 -12044
rect 13897 -14228 14083 -14016
rect 15547 -14048 15747 -12012
rect 17211 -12044 17294 -11832
rect 17159 -14016 17294 -12044
rect 14161 -14196 17133 -14048
rect 13897 -16200 14135 -14228
rect 10713 -16284 13685 -16232
rect 13897 -16388 14079 -16200
rect 15547 -16232 15747 -14196
rect 17211 -14228 17294 -14016
rect 17159 -16200 17294 -14228
rect 14161 -16284 17133 -16232
rect 17380 -16388 17938 -2852
rect -1948 -17053 17938 -16388
<< via1 >>
rect -668 1798 -596 1855
rect -468 1798 -396 1855
rect 28 1798 91 1855
rect -668 422 -596 1314
rect -1615 281 -1515 365
rect -668 -150 -596 -110
rect -1600 -243 -1550 -201
rect 1765 -16 1945 138
rect 5213 -16 5393 138
rect 6877 -16 7044 138
rect 8661 -16 8841 138
rect 10079 -73 10259 101
rect 12109 -16 12289 138
rect 13773 -16 13940 138
rect 15557 -16 15737 138
rect 1855 -238 1959 -121
rect 4161 -238 4341 -121
rect 4161 -583 4341 -491
rect 5925 -589 6024 -492
rect 1855 -950 1959 -852
rect 91 -16326 271 -16204
rect 2487 -15940 2579 -15829
rect 2487 -16305 2579 -16158
rect 7235 -1186 7319 -1006
rect 7501 -1729 7582 -1549
rect 7763 -2272 7847 -2092
rect 7931 -1186 8015 -1006
rect 8197 -1729 8277 -1549
rect 8459 -2272 8543 -2092
rect 8627 -1186 8711 -1006
rect 8893 -1729 8973 -1549
rect 9155 -2272 9239 -2092
rect 9323 -1186 9407 -1006
rect 9589 -1729 9669 -1549
rect 9851 -2272 9935 -2092
rect 10683 -1186 10767 -1006
rect 10949 -1729 11030 -1549
rect 11211 -2272 11295 -2092
rect 11379 -1186 11463 -1006
rect 11645 -1729 11726 -1549
rect 11907 -2272 11991 -2092
rect 12075 -1186 12159 -1006
rect 12341 -1729 12422 -1549
rect 12603 -2272 12687 -2092
rect 12771 -1186 12855 -1006
rect 13037 -1729 13118 -1549
rect 13299 -2272 13383 -2092
rect 14131 -1186 14215 -1006
rect 14397 -1729 14478 -1549
rect 14659 -2272 14743 -2092
rect 14827 -1186 14911 -1006
rect 15093 -1729 15174 -1549
rect 15355 -2272 15439 -2092
rect 15523 -1186 15607 -1006
rect 15789 -1729 15870 -1549
rect 16051 -2272 16135 -2092
rect 16219 -1186 16303 -1006
rect 16485 -1729 16566 -1549
rect 16747 -2272 16831 -2092
rect 10079 -3142 10259 -2998
rect 8661 -4384 8841 -4204
rect 10283 -4384 10388 -4204
rect 13527 -3142 13707 -2998
rect 12109 -4384 12289 -4204
rect 16975 -3142 17155 -2998
rect 15557 -4384 15737 -4204
<< metal2 >>
rect -678 1855 -586 1865
rect -678 1798 -668 1855
rect -596 1798 -586 1855
rect -678 1314 -586 1798
rect -478 1855 101 1865
rect -478 1798 -468 1855
rect -396 1798 28 1855
rect 91 1798 101 1855
rect -478 1788 101 1798
rect -678 422 -668 1314
rect -596 422 -586 1314
rect -1625 365 -1505 375
rect -1625 281 -1615 365
rect -1515 281 -1505 365
rect -1625 -201 -1505 281
rect -678 -110 -586 422
rect 1755 138 8851 148
rect 1755 -16 1765 138
rect 1945 -16 5213 138
rect 5393 -16 6877 138
rect 7044 -16 8661 138
rect 8841 -16 8851 138
rect 12099 138 17938 148
rect 1755 -26 8851 -16
rect 10069 101 10269 111
rect -678 -150 -668 -110
rect -596 -150 -586 -110
rect -678 -160 -586 -150
rect 1845 -121 1969 -111
rect -1625 -243 -1600 -201
rect -1550 -243 -1505 -201
rect -1625 -495 -1505 -243
rect 1845 -238 1855 -121
rect 1959 -238 1969 -121
rect 1845 -495 1969 -238
rect -1625 -613 1969 -495
rect 4151 -121 4351 -111
rect 4151 -238 4161 -121
rect 4341 -238 4351 -121
rect 4151 -491 4351 -238
rect 4151 -583 4161 -491
rect 4341 -583 4351 -491
rect 4151 -593 4351 -583
rect 5915 -492 6034 -26
rect 5915 -589 5925 -492
rect 6024 -589 6034 -492
rect 5915 -599 6034 -589
rect 10069 -73 10079 101
rect 10259 -73 10269 101
rect 12099 -16 12109 138
rect 12289 -16 13773 138
rect 13940 -16 15557 138
rect 15737 -16 17938 138
rect 12099 -26 17938 -16
rect 1845 -852 1969 -613
rect 1845 -950 1855 -852
rect 1959 -950 1969 -852
rect 1845 -960 1969 -950
rect 10069 -996 10269 -73
rect 13517 -996 13717 -26
rect 17053 -995 17940 -810
rect 16965 -996 17940 -995
rect 7225 -1006 10269 -996
rect 7225 -1186 7235 -1006
rect 7319 -1186 7931 -1006
rect 8015 -1186 8627 -1006
rect 8711 -1186 9323 -1006
rect 9407 -1186 10269 -1006
rect 7225 -1196 10269 -1186
rect 10673 -1006 13717 -996
rect 10673 -1186 10683 -1006
rect 10767 -1186 11379 -1006
rect 11463 -1186 12075 -1006
rect 12159 -1186 12771 -1006
rect 12855 -1186 13717 -1006
rect 10673 -1196 13717 -1186
rect 14121 -1006 17940 -996
rect 14121 -1186 14131 -1006
rect 14215 -1186 14827 -1006
rect 14911 -1186 15523 -1006
rect 15607 -1186 16219 -1006
rect 16303 -1186 17940 -1006
rect 14121 -1196 17940 -1186
rect 10069 -1539 10269 -1196
rect 17053 -1384 17940 -1196
rect 7225 -1549 17938 -1539
rect 7225 -1729 7501 -1549
rect 7582 -1729 8197 -1549
rect 8277 -1729 8893 -1549
rect 8973 -1729 9589 -1549
rect 9669 -1729 10949 -1549
rect 11030 -1729 11645 -1549
rect 11726 -1729 12341 -1549
rect 12422 -1729 13037 -1549
rect 13118 -1729 14397 -1549
rect 14478 -1729 15093 -1549
rect 15174 -1729 15789 -1549
rect 15870 -1729 16485 -1549
rect 16566 -1729 17938 -1549
rect 7225 -1739 17938 -1729
rect 7225 -2092 10269 -2082
rect 7225 -2272 7763 -2092
rect 7847 -2272 8459 -2092
rect 8543 -2272 9155 -2092
rect 9239 -2272 9851 -2092
rect 9935 -2272 10269 -2092
rect 7225 -2282 10269 -2272
rect 10673 -2092 13717 -2082
rect 10673 -2272 11211 -2092
rect 11295 -2272 11907 -2092
rect 11991 -2272 12603 -2092
rect 12687 -2272 13299 -2092
rect 13383 -2272 13717 -2092
rect 10673 -2282 13717 -2272
rect 14121 -2092 17165 -2082
rect 14121 -2272 14659 -2092
rect 14743 -2272 15355 -2092
rect 15439 -2272 16051 -2092
rect 16135 -2272 16747 -2092
rect 16831 -2272 17165 -2092
rect 14121 -2282 17165 -2272
rect 10069 -2998 10269 -2282
rect 10069 -3142 10079 -2998
rect 10259 -3142 10269 -2998
rect 10069 -3152 10269 -3142
rect 13517 -2998 13717 -2282
rect 13517 -3142 13527 -2998
rect 13707 -3142 13717 -2998
rect 13517 -3152 13717 -3142
rect 16965 -2998 17165 -2282
rect 16965 -3142 16975 -2998
rect 17155 -3142 17165 -2998
rect 16965 -3152 17165 -3142
rect 7197 -4204 17938 -4194
rect 7197 -4384 8661 -4204
rect 8841 -4384 10283 -4204
rect 10388 -4384 12109 -4204
rect 12289 -4384 15557 -4204
rect 15737 -4384 17938 -4204
rect 7197 -4394 17938 -4384
rect 2477 -15829 2589 -15819
rect 2477 -15940 2487 -15829
rect 2579 -15940 2589 -15829
rect 2477 -16158 2589 -15940
rect 81 -16204 281 -16194
rect 81 -16326 91 -16204
rect 271 -16235 281 -16204
rect 2477 -16235 2487 -16158
rect 271 -16305 2487 -16235
rect 2579 -16305 2589 -16158
rect 271 -16326 2589 -16305
rect 81 -16336 2589 -16326
use dpantenna_C8WG83  dpantenna_C8WG83_0
timestamp 1757240632
transform 1 0 -959 0 1 869
box -758 -758 758 758
use hvnmos_4SLWUS  hvnmos_4SLWUS_0
timestamp 1757240632
transform 0 1 -540 -1 0 -222
box -286 -1178 286 1178
use hvnmos_QQE73P  hvnmos_QQE73P_0
timestamp 1757240632
transform 1 0 7541 0 1 -1639
box -544 -1222 2356 1222
use hvnmos_QQE73P  hvnmos_QQE73P_1
timestamp 1757240632
transform 1 0 10989 0 1 -1639
box -544 -1222 2356 1222
use hvnmos_QQE73P  hvnmos_QQE73P_2
timestamp 1757240632
transform 1 0 14437 0 1 -1639
box -544 -1222 2356 1222
use hvnmos_RVVQDP  hvnmos_RVVQDP_0
timestamp 1757240632
transform 1 0 4251 0 1 -15319
box -1944 -722 1944 14930
use hvpmos_NE86AY  hvpmos_NE86AY_0
timestamp 1757240632
transform 1 0 1855 0 1 1273
box -1878 -1124 1878 12229
use hvpmos_NE86AY  hvpmos_NE86AY_1
timestamp 1757240632
transform 1 0 5303 0 1 1273
box -1878 -1124 1878 12229
use hvpmos_NE86AY  hvpmos_NE86AY_2
timestamp 1757240632
transform 1 0 8751 0 1 1273
box -1878 -1124 1878 12229
use hvpmos_NE86AY  hvpmos_NE86AY_3
timestamp 1757240632
transform 1 0 12199 0 1 1273
box -1878 -1124 1878 12229
use hvpmos_NE86AY  hvpmos_NE86AY_4
timestamp 1757240632
transform 1 0 15647 0 1 1273
box -1878 -1124 1878 12229
use lvnmos_533TXK  lvnmos_533TXK_0
timestamp 1757240632
transform 1 0 8751 0 1 -15214
box -1754 -1218 1754 11994
use lvnmos_533TXK  lvnmos_533TXK_1
timestamp 1757240632
transform 1 0 12199 0 1 -15214
box -1754 -1218 1754 11994
use lvnmos_533TXK  lvnmos_533TXK_2
timestamp 1757240632
transform 1 0 15647 0 1 -15214
box -1754 -1218 1754 11994
use lvnmos_RVV4EF  lvnmos_RVV4EF_0
timestamp 1757240632
transform 1 0 181 0 1 -15688
box -1896 -746 1896 14954
use rhigh_65D4BW  rhigh_65D4BW_0
timestamp 1757240632
transform 0 1 4253 -1 0 -16235
box -50 -1286 230 1286
use rhigh_RJR7YG  rhigh_RJR7YG_0
timestamp 1757240632
transform 1 0 -632 0 1 7451
box -230 -5766 430 5766
<< labels >>
flabel metal1 -1948 13355 -1198 14105 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 -1948 12464 -1198 13214 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal2 17545 -26 17938 148 0 FreeSans 800 0 0 0 VSOURCE
port 4 nsew
flabel metal1 17422 -637 17939 -120 0 FreeSans 800 0 0 0 ISOURCE
port 5 nsew
flabel metal2 17366 -1384 17940 -810 0 FreeSans 800 0 0 0 ISINK
port 6 nsew
flabel metal2 17549 -1739 17938 -1539 0 FreeSans 800 0 0 0 VSINKT
port 7 nsew
flabel metal2 17567 -4394 17938 -4194 0 FreeSans 800 0 0 0 VSINKB
port 9 nsew
flabel metal2 -635 1763 -635 1763 0 FreeSans 480 0 0 0 vs
flabel metal2 1910 -313 1910 -313 0 FreeSans 480 0 0 0 vp
flabel metal2 1891 -16291 1891 -16291 0 FreeSans 480 0 0 0 vth
flabel metal2 5973 -195 5973 -195 0 FreeSans 480 0 0 0 vm
<< end >>
