magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -924 6124 37600
<< isosubstrate >>
rect 50 23124 3950 28034
rect 50 18112 3950 22924
rect 50 13000 3950 17912
<< nwell >>
rect -124 33246 4124 33554
rect -124 29546 4124 29854
rect -124 1076 4124 12324
<< pwell >>
rect 24 31344 3976 31456
rect 24 12974 3976 28060
<< psubdiff >>
rect 184 31384 216 31416
rect 256 31384 288 31416
rect 328 31384 360 31416
rect 400 31384 432 31416
rect 472 31384 504 31416
rect 544 31384 576 31416
rect 616 31384 648 31416
rect 688 31384 720 31416
rect 760 31384 792 31416
rect 832 31384 864 31416
rect 904 31384 936 31416
rect 976 31384 1008 31416
rect 1048 31384 1080 31416
rect 1120 31384 1152 31416
rect 1192 31384 1224 31416
rect 1264 31384 1296 31416
rect 1336 31384 1368 31416
rect 1408 31384 1440 31416
rect 1480 31384 1512 31416
rect 1552 31384 1584 31416
rect 1624 31384 1656 31416
rect 1696 31384 1728 31416
rect 1768 31384 1800 31416
rect 1840 31384 1872 31416
rect 1912 31384 1944 31416
rect 1984 31384 2016 31416
rect 2056 31384 2088 31416
rect 2128 31384 2160 31416
rect 2200 31384 2232 31416
rect 2272 31384 2304 31416
rect 2344 31384 2376 31416
rect 2416 31384 2448 31416
rect 2488 31384 2520 31416
rect 2560 31384 2592 31416
rect 2632 31384 2664 31416
rect 2704 31384 2736 31416
rect 2776 31384 2808 31416
rect 2848 31384 2880 31416
rect 2920 31384 2952 31416
rect 2992 31384 3024 31416
rect 3064 31384 3096 31416
rect 3136 31384 3168 31416
rect 3208 31384 3240 31416
rect 3280 31384 3312 31416
rect 3352 31384 3384 31416
rect 3424 31384 3456 31416
rect 3496 31384 3528 31416
rect 3568 31384 3600 31416
rect 3640 31384 3672 31416
rect 3712 31384 3744 31416
rect 3784 31384 3816 31416
rect 3856 31384 3888 31416
rect 184 27939 216 27971
rect 256 27939 288 27971
rect 328 27939 360 27971
rect 400 27939 432 27971
rect 472 27939 504 27971
rect 544 27939 576 27971
rect 616 27939 648 27971
rect 688 27939 720 27971
rect 760 27939 792 27971
rect 832 27939 864 27971
rect 904 27939 936 27971
rect 976 27939 1008 27971
rect 1048 27939 1080 27971
rect 1120 27939 1152 27971
rect 1192 27939 1224 27971
rect 1264 27939 1296 27971
rect 1336 27939 1368 27971
rect 1408 27939 1440 27971
rect 1480 27939 1512 27971
rect 1552 27939 1584 27971
rect 1624 27939 1656 27971
rect 1696 27939 1728 27971
rect 1768 27939 1800 27971
rect 1840 27939 1872 27971
rect 1912 27939 1944 27971
rect 1984 27939 2016 27971
rect 2056 27939 2088 27971
rect 2128 27939 2160 27971
rect 2200 27939 2232 27971
rect 2272 27939 2304 27971
rect 2344 27939 2376 27971
rect 2416 27939 2448 27971
rect 2488 27939 2520 27971
rect 2560 27939 2592 27971
rect 2632 27939 2664 27971
rect 2704 27939 2736 27971
rect 2776 27939 2808 27971
rect 2848 27939 2880 27971
rect 2920 27939 2952 27971
rect 2992 27939 3024 27971
rect 3064 27939 3096 27971
rect 3136 27939 3168 27971
rect 3208 27939 3240 27971
rect 3280 27939 3312 27971
rect 3352 27939 3384 27971
rect 3424 27939 3456 27971
rect 3496 27939 3528 27971
rect 3568 27939 3600 27971
rect 3640 27939 3672 27971
rect 3712 27939 3744 27971
rect 3784 27939 3816 27971
rect 3856 27939 3888 27971
rect 112 27867 144 27899
rect 184 27867 216 27899
rect 256 27867 288 27899
rect 328 27867 360 27899
rect 400 27867 432 27899
rect 472 27867 504 27899
rect 544 27867 576 27899
rect 616 27867 648 27899
rect 688 27867 720 27899
rect 760 27867 792 27899
rect 832 27867 864 27899
rect 904 27867 936 27899
rect 976 27867 1008 27899
rect 1048 27867 1080 27899
rect 1120 27867 1152 27899
rect 1192 27867 1224 27899
rect 1264 27867 1296 27899
rect 1336 27867 1368 27899
rect 1408 27867 1440 27899
rect 1480 27867 1512 27899
rect 1552 27867 1584 27899
rect 1624 27867 1656 27899
rect 1696 27867 1728 27899
rect 1768 27867 1800 27899
rect 1840 27867 1872 27899
rect 1912 27867 1944 27899
rect 1984 27867 2016 27899
rect 2056 27867 2088 27899
rect 2128 27867 2160 27899
rect 2200 27867 2232 27899
rect 2272 27867 2304 27899
rect 2344 27867 2376 27899
rect 2416 27867 2448 27899
rect 2488 27867 2520 27899
rect 2560 27867 2592 27899
rect 2632 27867 2664 27899
rect 2704 27867 2736 27899
rect 2776 27867 2808 27899
rect 2848 27867 2880 27899
rect 2920 27867 2952 27899
rect 2992 27867 3024 27899
rect 3064 27867 3096 27899
rect 3136 27867 3168 27899
rect 3208 27867 3240 27899
rect 3280 27867 3312 27899
rect 3352 27867 3384 27899
rect 3424 27867 3456 27899
rect 3496 27867 3528 27899
rect 3568 27867 3600 27899
rect 3640 27867 3672 27899
rect 3712 27867 3744 27899
rect 3784 27867 3816 27899
rect 3856 27867 3888 27899
rect 112 27795 144 27827
rect 184 27795 216 27827
rect 256 27795 288 27827
rect 328 27795 360 27827
rect 400 27795 432 27827
rect 472 27795 504 27827
rect 544 27795 576 27827
rect 616 27795 648 27827
rect 688 27795 720 27827
rect 760 27795 792 27827
rect 832 27795 864 27827
rect 904 27795 936 27827
rect 976 27795 1008 27827
rect 1048 27795 1080 27827
rect 1120 27795 1152 27827
rect 1192 27795 1224 27827
rect 1264 27795 1296 27827
rect 1336 27795 1368 27827
rect 1408 27795 1440 27827
rect 1480 27795 1512 27827
rect 1552 27795 1584 27827
rect 1624 27795 1656 27827
rect 1696 27795 1728 27827
rect 1768 27795 1800 27827
rect 1840 27795 1872 27827
rect 1912 27795 1944 27827
rect 1984 27795 2016 27827
rect 2056 27795 2088 27827
rect 2128 27795 2160 27827
rect 2200 27795 2232 27827
rect 2272 27795 2304 27827
rect 2344 27795 2376 27827
rect 2416 27795 2448 27827
rect 2488 27795 2520 27827
rect 2560 27795 2592 27827
rect 2632 27795 2664 27827
rect 2704 27795 2736 27827
rect 2776 27795 2808 27827
rect 2848 27795 2880 27827
rect 2920 27795 2952 27827
rect 2992 27795 3024 27827
rect 3064 27795 3096 27827
rect 3136 27795 3168 27827
rect 3208 27795 3240 27827
rect 3280 27795 3312 27827
rect 3352 27795 3384 27827
rect 3424 27795 3456 27827
rect 3496 27795 3528 27827
rect 3568 27795 3600 27827
rect 3640 27795 3672 27827
rect 3712 27795 3744 27827
rect 3784 27795 3816 27827
rect 3856 27795 3888 27827
rect 112 27723 144 27755
rect 184 27723 216 27755
rect 256 27723 288 27755
rect 328 27723 360 27755
rect 400 27723 432 27755
rect 472 27723 504 27755
rect 544 27723 576 27755
rect 616 27723 648 27755
rect 688 27723 720 27755
rect 760 27723 792 27755
rect 832 27723 864 27755
rect 904 27723 936 27755
rect 976 27723 1008 27755
rect 1048 27723 1080 27755
rect 1120 27723 1152 27755
rect 1192 27723 1224 27755
rect 1264 27723 1296 27755
rect 1336 27723 1368 27755
rect 1408 27723 1440 27755
rect 1480 27723 1512 27755
rect 1552 27723 1584 27755
rect 1624 27723 1656 27755
rect 1696 27723 1728 27755
rect 1768 27723 1800 27755
rect 1840 27723 1872 27755
rect 1912 27723 1944 27755
rect 1984 27723 2016 27755
rect 2056 27723 2088 27755
rect 2128 27723 2160 27755
rect 2200 27723 2232 27755
rect 2272 27723 2304 27755
rect 2344 27723 2376 27755
rect 2416 27723 2448 27755
rect 2488 27723 2520 27755
rect 2560 27723 2592 27755
rect 2632 27723 2664 27755
rect 2704 27723 2736 27755
rect 2776 27723 2808 27755
rect 2848 27723 2880 27755
rect 2920 27723 2952 27755
rect 2992 27723 3024 27755
rect 3064 27723 3096 27755
rect 3136 27723 3168 27755
rect 3208 27723 3240 27755
rect 3280 27723 3312 27755
rect 3352 27723 3384 27755
rect 3424 27723 3456 27755
rect 3496 27723 3528 27755
rect 3568 27723 3600 27755
rect 3640 27723 3672 27755
rect 3712 27723 3744 27755
rect 3784 27723 3816 27755
rect 3856 27723 3888 27755
rect 112 27651 144 27683
rect 184 27651 216 27683
rect 256 27651 288 27683
rect 328 27651 360 27683
rect 400 27651 432 27683
rect 472 27651 504 27683
rect 544 27651 576 27683
rect 616 27651 648 27683
rect 688 27651 720 27683
rect 760 27651 792 27683
rect 832 27651 864 27683
rect 904 27651 936 27683
rect 976 27651 1008 27683
rect 1048 27651 1080 27683
rect 1120 27651 1152 27683
rect 1192 27651 1224 27683
rect 1264 27651 1296 27683
rect 1336 27651 1368 27683
rect 1408 27651 1440 27683
rect 1480 27651 1512 27683
rect 1552 27651 1584 27683
rect 1624 27651 1656 27683
rect 1696 27651 1728 27683
rect 1768 27651 1800 27683
rect 1840 27651 1872 27683
rect 1912 27651 1944 27683
rect 1984 27651 2016 27683
rect 2056 27651 2088 27683
rect 2128 27651 2160 27683
rect 2200 27651 2232 27683
rect 2272 27651 2304 27683
rect 2344 27651 2376 27683
rect 2416 27651 2448 27683
rect 2488 27651 2520 27683
rect 2560 27651 2592 27683
rect 2632 27651 2664 27683
rect 2704 27651 2736 27683
rect 2776 27651 2808 27683
rect 2848 27651 2880 27683
rect 2920 27651 2952 27683
rect 2992 27651 3024 27683
rect 3064 27651 3096 27683
rect 3136 27651 3168 27683
rect 3208 27651 3240 27683
rect 3280 27651 3312 27683
rect 3352 27651 3384 27683
rect 3424 27651 3456 27683
rect 3496 27651 3528 27683
rect 3568 27651 3600 27683
rect 3640 27651 3672 27683
rect 3712 27651 3744 27683
rect 3784 27651 3816 27683
rect 3856 27651 3888 27683
rect 112 27579 144 27611
rect 184 27579 216 27611
rect 256 27579 288 27611
rect 328 27579 360 27611
rect 400 27579 432 27611
rect 472 27579 504 27611
rect 544 27579 576 27611
rect 616 27579 648 27611
rect 688 27579 720 27611
rect 760 27579 792 27611
rect 832 27579 864 27611
rect 904 27579 936 27611
rect 976 27579 1008 27611
rect 1048 27579 1080 27611
rect 1120 27579 1152 27611
rect 1192 27579 1224 27611
rect 1264 27579 1296 27611
rect 1336 27579 1368 27611
rect 1408 27579 1440 27611
rect 1480 27579 1512 27611
rect 1552 27579 1584 27611
rect 1624 27579 1656 27611
rect 1696 27579 1728 27611
rect 1768 27579 1800 27611
rect 1840 27579 1872 27611
rect 1912 27579 1944 27611
rect 1984 27579 2016 27611
rect 2056 27579 2088 27611
rect 2128 27579 2160 27611
rect 2200 27579 2232 27611
rect 2272 27579 2304 27611
rect 2344 27579 2376 27611
rect 2416 27579 2448 27611
rect 2488 27579 2520 27611
rect 2560 27579 2592 27611
rect 2632 27579 2664 27611
rect 2704 27579 2736 27611
rect 2776 27579 2808 27611
rect 2848 27579 2880 27611
rect 2920 27579 2952 27611
rect 2992 27579 3024 27611
rect 3064 27579 3096 27611
rect 3136 27579 3168 27611
rect 3208 27579 3240 27611
rect 3280 27579 3312 27611
rect 3352 27579 3384 27611
rect 3424 27579 3456 27611
rect 3496 27579 3528 27611
rect 3568 27579 3600 27611
rect 3640 27579 3672 27611
rect 3712 27579 3744 27611
rect 3784 27579 3816 27611
rect 3856 27579 3888 27611
rect 112 27507 144 27539
rect 184 27507 216 27539
rect 256 27507 288 27539
rect 328 27507 360 27539
rect 400 27507 432 27539
rect 472 27507 504 27539
rect 544 27507 576 27539
rect 616 27507 648 27539
rect 688 27507 720 27539
rect 760 27507 792 27539
rect 832 27507 864 27539
rect 904 27507 936 27539
rect 976 27507 1008 27539
rect 1048 27507 1080 27539
rect 1120 27507 1152 27539
rect 1192 27507 1224 27539
rect 1264 27507 1296 27539
rect 1336 27507 1368 27539
rect 1408 27507 1440 27539
rect 1480 27507 1512 27539
rect 1552 27507 1584 27539
rect 1624 27507 1656 27539
rect 1696 27507 1728 27539
rect 1768 27507 1800 27539
rect 1840 27507 1872 27539
rect 1912 27507 1944 27539
rect 1984 27507 2016 27539
rect 2056 27507 2088 27539
rect 2128 27507 2160 27539
rect 2200 27507 2232 27539
rect 2272 27507 2304 27539
rect 2344 27507 2376 27539
rect 2416 27507 2448 27539
rect 2488 27507 2520 27539
rect 2560 27507 2592 27539
rect 2632 27507 2664 27539
rect 2704 27507 2736 27539
rect 2776 27507 2808 27539
rect 2848 27507 2880 27539
rect 2920 27507 2952 27539
rect 2992 27507 3024 27539
rect 3064 27507 3096 27539
rect 3136 27507 3168 27539
rect 3208 27507 3240 27539
rect 3280 27507 3312 27539
rect 3352 27507 3384 27539
rect 3424 27507 3456 27539
rect 3496 27507 3528 27539
rect 3568 27507 3600 27539
rect 3640 27507 3672 27539
rect 3712 27507 3744 27539
rect 3784 27507 3816 27539
rect 3856 27507 3888 27539
rect 112 27435 144 27467
rect 184 27435 216 27467
rect 256 27435 288 27467
rect 328 27435 360 27467
rect 400 27435 432 27467
rect 472 27435 504 27467
rect 544 27435 576 27467
rect 616 27435 648 27467
rect 688 27435 720 27467
rect 760 27435 792 27467
rect 832 27435 864 27467
rect 904 27435 936 27467
rect 976 27435 1008 27467
rect 1048 27435 1080 27467
rect 1120 27435 1152 27467
rect 1192 27435 1224 27467
rect 1264 27435 1296 27467
rect 1336 27435 1368 27467
rect 1408 27435 1440 27467
rect 1480 27435 1512 27467
rect 1552 27435 1584 27467
rect 1624 27435 1656 27467
rect 1696 27435 1728 27467
rect 1768 27435 1800 27467
rect 1840 27435 1872 27467
rect 1912 27435 1944 27467
rect 1984 27435 2016 27467
rect 2056 27435 2088 27467
rect 2128 27435 2160 27467
rect 2200 27435 2232 27467
rect 2272 27435 2304 27467
rect 2344 27435 2376 27467
rect 2416 27435 2448 27467
rect 2488 27435 2520 27467
rect 2560 27435 2592 27467
rect 2632 27435 2664 27467
rect 2704 27435 2736 27467
rect 2776 27435 2808 27467
rect 2848 27435 2880 27467
rect 2920 27435 2952 27467
rect 2992 27435 3024 27467
rect 3064 27435 3096 27467
rect 3136 27435 3168 27467
rect 3208 27435 3240 27467
rect 3280 27435 3312 27467
rect 3352 27435 3384 27467
rect 3424 27435 3456 27467
rect 3496 27435 3528 27467
rect 3568 27435 3600 27467
rect 3640 27435 3672 27467
rect 3712 27435 3744 27467
rect 3784 27435 3816 27467
rect 3856 27435 3888 27467
rect 112 27363 144 27395
rect 184 27363 216 27395
rect 256 27363 288 27395
rect 328 27363 360 27395
rect 400 27363 432 27395
rect 472 27363 504 27395
rect 544 27363 576 27395
rect 616 27363 648 27395
rect 688 27363 720 27395
rect 760 27363 792 27395
rect 832 27363 864 27395
rect 904 27363 936 27395
rect 976 27363 1008 27395
rect 1048 27363 1080 27395
rect 1120 27363 1152 27395
rect 1192 27363 1224 27395
rect 1264 27363 1296 27395
rect 1336 27363 1368 27395
rect 1408 27363 1440 27395
rect 1480 27363 1512 27395
rect 1552 27363 1584 27395
rect 1624 27363 1656 27395
rect 1696 27363 1728 27395
rect 1768 27363 1800 27395
rect 1840 27363 1872 27395
rect 1912 27363 1944 27395
rect 1984 27363 2016 27395
rect 2056 27363 2088 27395
rect 2128 27363 2160 27395
rect 2200 27363 2232 27395
rect 2272 27363 2304 27395
rect 2344 27363 2376 27395
rect 2416 27363 2448 27395
rect 2488 27363 2520 27395
rect 2560 27363 2592 27395
rect 2632 27363 2664 27395
rect 2704 27363 2736 27395
rect 2776 27363 2808 27395
rect 2848 27363 2880 27395
rect 2920 27363 2952 27395
rect 2992 27363 3024 27395
rect 3064 27363 3096 27395
rect 3136 27363 3168 27395
rect 3208 27363 3240 27395
rect 3280 27363 3312 27395
rect 3352 27363 3384 27395
rect 3424 27363 3456 27395
rect 3496 27363 3528 27395
rect 3568 27363 3600 27395
rect 3640 27363 3672 27395
rect 3712 27363 3744 27395
rect 3784 27363 3816 27395
rect 3856 27363 3888 27395
rect 112 27291 144 27323
rect 184 27291 216 27323
rect 256 27291 288 27323
rect 328 27291 360 27323
rect 400 27291 432 27323
rect 472 27291 504 27323
rect 544 27291 576 27323
rect 616 27291 648 27323
rect 688 27291 720 27323
rect 760 27291 792 27323
rect 832 27291 864 27323
rect 904 27291 936 27323
rect 976 27291 1008 27323
rect 1048 27291 1080 27323
rect 1120 27291 1152 27323
rect 1192 27291 1224 27323
rect 1264 27291 1296 27323
rect 1336 27291 1368 27323
rect 1408 27291 1440 27323
rect 1480 27291 1512 27323
rect 1552 27291 1584 27323
rect 1624 27291 1656 27323
rect 1696 27291 1728 27323
rect 1768 27291 1800 27323
rect 1840 27291 1872 27323
rect 1912 27291 1944 27323
rect 1984 27291 2016 27323
rect 2056 27291 2088 27323
rect 2128 27291 2160 27323
rect 2200 27291 2232 27323
rect 2272 27291 2304 27323
rect 2344 27291 2376 27323
rect 2416 27291 2448 27323
rect 2488 27291 2520 27323
rect 2560 27291 2592 27323
rect 2632 27291 2664 27323
rect 2704 27291 2736 27323
rect 2776 27291 2808 27323
rect 2848 27291 2880 27323
rect 2920 27291 2952 27323
rect 2992 27291 3024 27323
rect 3064 27291 3096 27323
rect 3136 27291 3168 27323
rect 3208 27291 3240 27323
rect 3280 27291 3312 27323
rect 3352 27291 3384 27323
rect 3424 27291 3456 27323
rect 3496 27291 3528 27323
rect 3568 27291 3600 27323
rect 3640 27291 3672 27323
rect 3712 27291 3744 27323
rect 3784 27291 3816 27323
rect 3856 27291 3888 27323
rect 112 27219 144 27251
rect 184 27219 216 27251
rect 256 27219 288 27251
rect 328 27219 360 27251
rect 400 27219 432 27251
rect 472 27219 504 27251
rect 544 27219 576 27251
rect 616 27219 648 27251
rect 688 27219 720 27251
rect 760 27219 792 27251
rect 832 27219 864 27251
rect 904 27219 936 27251
rect 976 27219 1008 27251
rect 1048 27219 1080 27251
rect 1120 27219 1152 27251
rect 1192 27219 1224 27251
rect 1264 27219 1296 27251
rect 1336 27219 1368 27251
rect 1408 27219 1440 27251
rect 1480 27219 1512 27251
rect 1552 27219 1584 27251
rect 1624 27219 1656 27251
rect 1696 27219 1728 27251
rect 1768 27219 1800 27251
rect 1840 27219 1872 27251
rect 1912 27219 1944 27251
rect 1984 27219 2016 27251
rect 2056 27219 2088 27251
rect 2128 27219 2160 27251
rect 2200 27219 2232 27251
rect 2272 27219 2304 27251
rect 2344 27219 2376 27251
rect 2416 27219 2448 27251
rect 2488 27219 2520 27251
rect 2560 27219 2592 27251
rect 2632 27219 2664 27251
rect 2704 27219 2736 27251
rect 2776 27219 2808 27251
rect 2848 27219 2880 27251
rect 2920 27219 2952 27251
rect 2992 27219 3024 27251
rect 3064 27219 3096 27251
rect 3136 27219 3168 27251
rect 3208 27219 3240 27251
rect 3280 27219 3312 27251
rect 3352 27219 3384 27251
rect 3424 27219 3456 27251
rect 3496 27219 3528 27251
rect 3568 27219 3600 27251
rect 3640 27219 3672 27251
rect 3712 27219 3744 27251
rect 3784 27219 3816 27251
rect 3856 27219 3888 27251
rect 112 27147 144 27179
rect 184 27147 216 27179
rect 256 27147 288 27179
rect 328 27147 360 27179
rect 400 27147 432 27179
rect 472 27147 504 27179
rect 544 27147 576 27179
rect 616 27147 648 27179
rect 688 27147 720 27179
rect 760 27147 792 27179
rect 832 27147 864 27179
rect 904 27147 936 27179
rect 976 27147 1008 27179
rect 1048 27147 1080 27179
rect 1120 27147 1152 27179
rect 1192 27147 1224 27179
rect 1264 27147 1296 27179
rect 1336 27147 1368 27179
rect 1408 27147 1440 27179
rect 1480 27147 1512 27179
rect 1552 27147 1584 27179
rect 1624 27147 1656 27179
rect 1696 27147 1728 27179
rect 1768 27147 1800 27179
rect 1840 27147 1872 27179
rect 1912 27147 1944 27179
rect 1984 27147 2016 27179
rect 2056 27147 2088 27179
rect 2128 27147 2160 27179
rect 2200 27147 2232 27179
rect 2272 27147 2304 27179
rect 2344 27147 2376 27179
rect 2416 27147 2448 27179
rect 2488 27147 2520 27179
rect 2560 27147 2592 27179
rect 2632 27147 2664 27179
rect 2704 27147 2736 27179
rect 2776 27147 2808 27179
rect 2848 27147 2880 27179
rect 2920 27147 2952 27179
rect 2992 27147 3024 27179
rect 3064 27147 3096 27179
rect 3136 27147 3168 27179
rect 3208 27147 3240 27179
rect 3280 27147 3312 27179
rect 3352 27147 3384 27179
rect 3424 27147 3456 27179
rect 3496 27147 3528 27179
rect 3568 27147 3600 27179
rect 3640 27147 3672 27179
rect 3712 27147 3744 27179
rect 3784 27147 3816 27179
rect 3856 27147 3888 27179
rect 112 27075 144 27107
rect 184 27075 216 27107
rect 256 27075 288 27107
rect 328 27075 360 27107
rect 400 27075 432 27107
rect 472 27075 504 27107
rect 544 27075 576 27107
rect 616 27075 648 27107
rect 688 27075 720 27107
rect 760 27075 792 27107
rect 832 27075 864 27107
rect 904 27075 936 27107
rect 976 27075 1008 27107
rect 1048 27075 1080 27107
rect 1120 27075 1152 27107
rect 1192 27075 1224 27107
rect 1264 27075 1296 27107
rect 1336 27075 1368 27107
rect 1408 27075 1440 27107
rect 1480 27075 1512 27107
rect 1552 27075 1584 27107
rect 1624 27075 1656 27107
rect 1696 27075 1728 27107
rect 1768 27075 1800 27107
rect 1840 27075 1872 27107
rect 1912 27075 1944 27107
rect 1984 27075 2016 27107
rect 2056 27075 2088 27107
rect 2128 27075 2160 27107
rect 2200 27075 2232 27107
rect 2272 27075 2304 27107
rect 2344 27075 2376 27107
rect 2416 27075 2448 27107
rect 2488 27075 2520 27107
rect 2560 27075 2592 27107
rect 2632 27075 2664 27107
rect 2704 27075 2736 27107
rect 2776 27075 2808 27107
rect 2848 27075 2880 27107
rect 2920 27075 2952 27107
rect 2992 27075 3024 27107
rect 3064 27075 3096 27107
rect 3136 27075 3168 27107
rect 3208 27075 3240 27107
rect 3280 27075 3312 27107
rect 3352 27075 3384 27107
rect 3424 27075 3456 27107
rect 3496 27075 3528 27107
rect 3568 27075 3600 27107
rect 3640 27075 3672 27107
rect 3712 27075 3744 27107
rect 3784 27075 3816 27107
rect 3856 27075 3888 27107
rect 112 27003 144 27035
rect 184 27003 216 27035
rect 256 27003 288 27035
rect 328 27003 360 27035
rect 400 27003 432 27035
rect 472 27003 504 27035
rect 544 27003 576 27035
rect 616 27003 648 27035
rect 688 27003 720 27035
rect 760 27003 792 27035
rect 832 27003 864 27035
rect 904 27003 936 27035
rect 976 27003 1008 27035
rect 1048 27003 1080 27035
rect 1120 27003 1152 27035
rect 1192 27003 1224 27035
rect 1264 27003 1296 27035
rect 1336 27003 1368 27035
rect 1408 27003 1440 27035
rect 1480 27003 1512 27035
rect 1552 27003 1584 27035
rect 1624 27003 1656 27035
rect 1696 27003 1728 27035
rect 1768 27003 1800 27035
rect 1840 27003 1872 27035
rect 1912 27003 1944 27035
rect 1984 27003 2016 27035
rect 2056 27003 2088 27035
rect 2128 27003 2160 27035
rect 2200 27003 2232 27035
rect 2272 27003 2304 27035
rect 2344 27003 2376 27035
rect 2416 27003 2448 27035
rect 2488 27003 2520 27035
rect 2560 27003 2592 27035
rect 2632 27003 2664 27035
rect 2704 27003 2736 27035
rect 2776 27003 2808 27035
rect 2848 27003 2880 27035
rect 2920 27003 2952 27035
rect 2992 27003 3024 27035
rect 3064 27003 3096 27035
rect 3136 27003 3168 27035
rect 3208 27003 3240 27035
rect 3280 27003 3312 27035
rect 3352 27003 3384 27035
rect 3424 27003 3456 27035
rect 3496 27003 3528 27035
rect 3568 27003 3600 27035
rect 3640 27003 3672 27035
rect 3712 27003 3744 27035
rect 3784 27003 3816 27035
rect 3856 27003 3888 27035
rect 112 26931 144 26963
rect 184 26931 216 26963
rect 256 26931 288 26963
rect 328 26931 360 26963
rect 400 26931 432 26963
rect 472 26931 504 26963
rect 544 26931 576 26963
rect 616 26931 648 26963
rect 688 26931 720 26963
rect 760 26931 792 26963
rect 832 26931 864 26963
rect 904 26931 936 26963
rect 976 26931 1008 26963
rect 1048 26931 1080 26963
rect 1120 26931 1152 26963
rect 1192 26931 1224 26963
rect 1264 26931 1296 26963
rect 1336 26931 1368 26963
rect 1408 26931 1440 26963
rect 1480 26931 1512 26963
rect 1552 26931 1584 26963
rect 1624 26931 1656 26963
rect 1696 26931 1728 26963
rect 1768 26931 1800 26963
rect 1840 26931 1872 26963
rect 1912 26931 1944 26963
rect 1984 26931 2016 26963
rect 2056 26931 2088 26963
rect 2128 26931 2160 26963
rect 2200 26931 2232 26963
rect 2272 26931 2304 26963
rect 2344 26931 2376 26963
rect 2416 26931 2448 26963
rect 2488 26931 2520 26963
rect 2560 26931 2592 26963
rect 2632 26931 2664 26963
rect 2704 26931 2736 26963
rect 2776 26931 2808 26963
rect 2848 26931 2880 26963
rect 2920 26931 2952 26963
rect 2992 26931 3024 26963
rect 3064 26931 3096 26963
rect 3136 26931 3168 26963
rect 3208 26931 3240 26963
rect 3280 26931 3312 26963
rect 3352 26931 3384 26963
rect 3424 26931 3456 26963
rect 3496 26931 3528 26963
rect 3568 26931 3600 26963
rect 3640 26931 3672 26963
rect 3712 26931 3744 26963
rect 3784 26931 3816 26963
rect 3856 26931 3888 26963
rect 112 26859 144 26891
rect 184 26859 216 26891
rect 256 26859 288 26891
rect 328 26859 360 26891
rect 400 26859 432 26891
rect 472 26859 504 26891
rect 544 26859 576 26891
rect 616 26859 648 26891
rect 688 26859 720 26891
rect 760 26859 792 26891
rect 832 26859 864 26891
rect 904 26859 936 26891
rect 976 26859 1008 26891
rect 1048 26859 1080 26891
rect 1120 26859 1152 26891
rect 1192 26859 1224 26891
rect 1264 26859 1296 26891
rect 1336 26859 1368 26891
rect 1408 26859 1440 26891
rect 1480 26859 1512 26891
rect 1552 26859 1584 26891
rect 1624 26859 1656 26891
rect 1696 26859 1728 26891
rect 1768 26859 1800 26891
rect 1840 26859 1872 26891
rect 1912 26859 1944 26891
rect 1984 26859 2016 26891
rect 2056 26859 2088 26891
rect 2128 26859 2160 26891
rect 2200 26859 2232 26891
rect 2272 26859 2304 26891
rect 2344 26859 2376 26891
rect 2416 26859 2448 26891
rect 2488 26859 2520 26891
rect 2560 26859 2592 26891
rect 2632 26859 2664 26891
rect 2704 26859 2736 26891
rect 2776 26859 2808 26891
rect 2848 26859 2880 26891
rect 2920 26859 2952 26891
rect 2992 26859 3024 26891
rect 3064 26859 3096 26891
rect 3136 26859 3168 26891
rect 3208 26859 3240 26891
rect 3280 26859 3312 26891
rect 3352 26859 3384 26891
rect 3424 26859 3456 26891
rect 3496 26859 3528 26891
rect 3568 26859 3600 26891
rect 3640 26859 3672 26891
rect 3712 26859 3744 26891
rect 3784 26859 3816 26891
rect 3856 26859 3888 26891
rect 112 26787 144 26819
rect 184 26787 216 26819
rect 256 26787 288 26819
rect 328 26787 360 26819
rect 400 26787 432 26819
rect 472 26787 504 26819
rect 544 26787 576 26819
rect 616 26787 648 26819
rect 688 26787 720 26819
rect 760 26787 792 26819
rect 832 26787 864 26819
rect 904 26787 936 26819
rect 976 26787 1008 26819
rect 1048 26787 1080 26819
rect 1120 26787 1152 26819
rect 1192 26787 1224 26819
rect 1264 26787 1296 26819
rect 1336 26787 1368 26819
rect 1408 26787 1440 26819
rect 1480 26787 1512 26819
rect 1552 26787 1584 26819
rect 1624 26787 1656 26819
rect 1696 26787 1728 26819
rect 1768 26787 1800 26819
rect 1840 26787 1872 26819
rect 1912 26787 1944 26819
rect 1984 26787 2016 26819
rect 2056 26787 2088 26819
rect 2128 26787 2160 26819
rect 2200 26787 2232 26819
rect 2272 26787 2304 26819
rect 2344 26787 2376 26819
rect 2416 26787 2448 26819
rect 2488 26787 2520 26819
rect 2560 26787 2592 26819
rect 2632 26787 2664 26819
rect 2704 26787 2736 26819
rect 2776 26787 2808 26819
rect 2848 26787 2880 26819
rect 2920 26787 2952 26819
rect 2992 26787 3024 26819
rect 3064 26787 3096 26819
rect 3136 26787 3168 26819
rect 3208 26787 3240 26819
rect 3280 26787 3312 26819
rect 3352 26787 3384 26819
rect 3424 26787 3456 26819
rect 3496 26787 3528 26819
rect 3568 26787 3600 26819
rect 3640 26787 3672 26819
rect 3712 26787 3744 26819
rect 3784 26787 3816 26819
rect 3856 26787 3888 26819
rect 112 26715 144 26747
rect 184 26715 216 26747
rect 256 26715 288 26747
rect 328 26715 360 26747
rect 400 26715 432 26747
rect 472 26715 504 26747
rect 544 26715 576 26747
rect 616 26715 648 26747
rect 688 26715 720 26747
rect 760 26715 792 26747
rect 832 26715 864 26747
rect 904 26715 936 26747
rect 976 26715 1008 26747
rect 1048 26715 1080 26747
rect 1120 26715 1152 26747
rect 1192 26715 1224 26747
rect 1264 26715 1296 26747
rect 1336 26715 1368 26747
rect 1408 26715 1440 26747
rect 1480 26715 1512 26747
rect 1552 26715 1584 26747
rect 1624 26715 1656 26747
rect 1696 26715 1728 26747
rect 1768 26715 1800 26747
rect 1840 26715 1872 26747
rect 1912 26715 1944 26747
rect 1984 26715 2016 26747
rect 2056 26715 2088 26747
rect 2128 26715 2160 26747
rect 2200 26715 2232 26747
rect 2272 26715 2304 26747
rect 2344 26715 2376 26747
rect 2416 26715 2448 26747
rect 2488 26715 2520 26747
rect 2560 26715 2592 26747
rect 2632 26715 2664 26747
rect 2704 26715 2736 26747
rect 2776 26715 2808 26747
rect 2848 26715 2880 26747
rect 2920 26715 2952 26747
rect 2992 26715 3024 26747
rect 3064 26715 3096 26747
rect 3136 26715 3168 26747
rect 3208 26715 3240 26747
rect 3280 26715 3312 26747
rect 3352 26715 3384 26747
rect 3424 26715 3456 26747
rect 3496 26715 3528 26747
rect 3568 26715 3600 26747
rect 3640 26715 3672 26747
rect 3712 26715 3744 26747
rect 3784 26715 3816 26747
rect 3856 26715 3888 26747
rect 112 26643 144 26675
rect 184 26643 216 26675
rect 256 26643 288 26675
rect 328 26643 360 26675
rect 400 26643 432 26675
rect 472 26643 504 26675
rect 544 26643 576 26675
rect 616 26643 648 26675
rect 688 26643 720 26675
rect 760 26643 792 26675
rect 832 26643 864 26675
rect 904 26643 936 26675
rect 976 26643 1008 26675
rect 1048 26643 1080 26675
rect 1120 26643 1152 26675
rect 1192 26643 1224 26675
rect 1264 26643 1296 26675
rect 1336 26643 1368 26675
rect 1408 26643 1440 26675
rect 1480 26643 1512 26675
rect 1552 26643 1584 26675
rect 1624 26643 1656 26675
rect 1696 26643 1728 26675
rect 1768 26643 1800 26675
rect 1840 26643 1872 26675
rect 1912 26643 1944 26675
rect 1984 26643 2016 26675
rect 2056 26643 2088 26675
rect 2128 26643 2160 26675
rect 2200 26643 2232 26675
rect 2272 26643 2304 26675
rect 2344 26643 2376 26675
rect 2416 26643 2448 26675
rect 2488 26643 2520 26675
rect 2560 26643 2592 26675
rect 2632 26643 2664 26675
rect 2704 26643 2736 26675
rect 2776 26643 2808 26675
rect 2848 26643 2880 26675
rect 2920 26643 2952 26675
rect 2992 26643 3024 26675
rect 3064 26643 3096 26675
rect 3136 26643 3168 26675
rect 3208 26643 3240 26675
rect 3280 26643 3312 26675
rect 3352 26643 3384 26675
rect 3424 26643 3456 26675
rect 3496 26643 3528 26675
rect 3568 26643 3600 26675
rect 3640 26643 3672 26675
rect 3712 26643 3744 26675
rect 3784 26643 3816 26675
rect 3856 26643 3888 26675
rect 112 26571 144 26603
rect 184 26571 216 26603
rect 256 26571 288 26603
rect 328 26571 360 26603
rect 400 26571 432 26603
rect 472 26571 504 26603
rect 544 26571 576 26603
rect 616 26571 648 26603
rect 688 26571 720 26603
rect 760 26571 792 26603
rect 832 26571 864 26603
rect 904 26571 936 26603
rect 976 26571 1008 26603
rect 1048 26571 1080 26603
rect 1120 26571 1152 26603
rect 1192 26571 1224 26603
rect 1264 26571 1296 26603
rect 1336 26571 1368 26603
rect 1408 26571 1440 26603
rect 1480 26571 1512 26603
rect 1552 26571 1584 26603
rect 1624 26571 1656 26603
rect 1696 26571 1728 26603
rect 1768 26571 1800 26603
rect 1840 26571 1872 26603
rect 1912 26571 1944 26603
rect 1984 26571 2016 26603
rect 2056 26571 2088 26603
rect 2128 26571 2160 26603
rect 2200 26571 2232 26603
rect 2272 26571 2304 26603
rect 2344 26571 2376 26603
rect 2416 26571 2448 26603
rect 2488 26571 2520 26603
rect 2560 26571 2592 26603
rect 2632 26571 2664 26603
rect 2704 26571 2736 26603
rect 2776 26571 2808 26603
rect 2848 26571 2880 26603
rect 2920 26571 2952 26603
rect 2992 26571 3024 26603
rect 3064 26571 3096 26603
rect 3136 26571 3168 26603
rect 3208 26571 3240 26603
rect 3280 26571 3312 26603
rect 3352 26571 3384 26603
rect 3424 26571 3456 26603
rect 3496 26571 3528 26603
rect 3568 26571 3600 26603
rect 3640 26571 3672 26603
rect 3712 26571 3744 26603
rect 3784 26571 3816 26603
rect 3856 26571 3888 26603
rect 112 26499 144 26531
rect 184 26499 216 26531
rect 256 26499 288 26531
rect 328 26499 360 26531
rect 400 26499 432 26531
rect 472 26499 504 26531
rect 544 26499 576 26531
rect 616 26499 648 26531
rect 688 26499 720 26531
rect 760 26499 792 26531
rect 832 26499 864 26531
rect 904 26499 936 26531
rect 976 26499 1008 26531
rect 1048 26499 1080 26531
rect 1120 26499 1152 26531
rect 1192 26499 1224 26531
rect 1264 26499 1296 26531
rect 1336 26499 1368 26531
rect 1408 26499 1440 26531
rect 1480 26499 1512 26531
rect 1552 26499 1584 26531
rect 1624 26499 1656 26531
rect 1696 26499 1728 26531
rect 1768 26499 1800 26531
rect 1840 26499 1872 26531
rect 1912 26499 1944 26531
rect 1984 26499 2016 26531
rect 2056 26499 2088 26531
rect 2128 26499 2160 26531
rect 2200 26499 2232 26531
rect 2272 26499 2304 26531
rect 2344 26499 2376 26531
rect 2416 26499 2448 26531
rect 2488 26499 2520 26531
rect 2560 26499 2592 26531
rect 2632 26499 2664 26531
rect 2704 26499 2736 26531
rect 2776 26499 2808 26531
rect 2848 26499 2880 26531
rect 2920 26499 2952 26531
rect 2992 26499 3024 26531
rect 3064 26499 3096 26531
rect 3136 26499 3168 26531
rect 3208 26499 3240 26531
rect 3280 26499 3312 26531
rect 3352 26499 3384 26531
rect 3424 26499 3456 26531
rect 3496 26499 3528 26531
rect 3568 26499 3600 26531
rect 3640 26499 3672 26531
rect 3712 26499 3744 26531
rect 3784 26499 3816 26531
rect 3856 26499 3888 26531
rect 112 26427 144 26459
rect 184 26427 216 26459
rect 256 26427 288 26459
rect 328 26427 360 26459
rect 400 26427 432 26459
rect 472 26427 504 26459
rect 544 26427 576 26459
rect 616 26427 648 26459
rect 688 26427 720 26459
rect 760 26427 792 26459
rect 832 26427 864 26459
rect 904 26427 936 26459
rect 976 26427 1008 26459
rect 1048 26427 1080 26459
rect 1120 26427 1152 26459
rect 1192 26427 1224 26459
rect 1264 26427 1296 26459
rect 1336 26427 1368 26459
rect 1408 26427 1440 26459
rect 1480 26427 1512 26459
rect 1552 26427 1584 26459
rect 1624 26427 1656 26459
rect 1696 26427 1728 26459
rect 1768 26427 1800 26459
rect 1840 26427 1872 26459
rect 1912 26427 1944 26459
rect 1984 26427 2016 26459
rect 2056 26427 2088 26459
rect 2128 26427 2160 26459
rect 2200 26427 2232 26459
rect 2272 26427 2304 26459
rect 2344 26427 2376 26459
rect 2416 26427 2448 26459
rect 2488 26427 2520 26459
rect 2560 26427 2592 26459
rect 2632 26427 2664 26459
rect 2704 26427 2736 26459
rect 2776 26427 2808 26459
rect 2848 26427 2880 26459
rect 2920 26427 2952 26459
rect 2992 26427 3024 26459
rect 3064 26427 3096 26459
rect 3136 26427 3168 26459
rect 3208 26427 3240 26459
rect 3280 26427 3312 26459
rect 3352 26427 3384 26459
rect 3424 26427 3456 26459
rect 3496 26427 3528 26459
rect 3568 26427 3600 26459
rect 3640 26427 3672 26459
rect 3712 26427 3744 26459
rect 3784 26427 3816 26459
rect 3856 26427 3888 26459
rect 112 26355 144 26387
rect 184 26355 216 26387
rect 256 26355 288 26387
rect 328 26355 360 26387
rect 400 26355 432 26387
rect 472 26355 504 26387
rect 544 26355 576 26387
rect 616 26355 648 26387
rect 688 26355 720 26387
rect 760 26355 792 26387
rect 832 26355 864 26387
rect 904 26355 936 26387
rect 976 26355 1008 26387
rect 1048 26355 1080 26387
rect 1120 26355 1152 26387
rect 1192 26355 1224 26387
rect 1264 26355 1296 26387
rect 1336 26355 1368 26387
rect 1408 26355 1440 26387
rect 1480 26355 1512 26387
rect 1552 26355 1584 26387
rect 1624 26355 1656 26387
rect 1696 26355 1728 26387
rect 1768 26355 1800 26387
rect 1840 26355 1872 26387
rect 1912 26355 1944 26387
rect 1984 26355 2016 26387
rect 2056 26355 2088 26387
rect 2128 26355 2160 26387
rect 2200 26355 2232 26387
rect 2272 26355 2304 26387
rect 2344 26355 2376 26387
rect 2416 26355 2448 26387
rect 2488 26355 2520 26387
rect 2560 26355 2592 26387
rect 2632 26355 2664 26387
rect 2704 26355 2736 26387
rect 2776 26355 2808 26387
rect 2848 26355 2880 26387
rect 2920 26355 2952 26387
rect 2992 26355 3024 26387
rect 3064 26355 3096 26387
rect 3136 26355 3168 26387
rect 3208 26355 3240 26387
rect 3280 26355 3312 26387
rect 3352 26355 3384 26387
rect 3424 26355 3456 26387
rect 3496 26355 3528 26387
rect 3568 26355 3600 26387
rect 3640 26355 3672 26387
rect 3712 26355 3744 26387
rect 3784 26355 3816 26387
rect 3856 26355 3888 26387
rect 112 26283 144 26315
rect 184 26283 216 26315
rect 256 26283 288 26315
rect 328 26283 360 26315
rect 400 26283 432 26315
rect 472 26283 504 26315
rect 544 26283 576 26315
rect 616 26283 648 26315
rect 688 26283 720 26315
rect 760 26283 792 26315
rect 832 26283 864 26315
rect 904 26283 936 26315
rect 976 26283 1008 26315
rect 1048 26283 1080 26315
rect 1120 26283 1152 26315
rect 1192 26283 1224 26315
rect 1264 26283 1296 26315
rect 1336 26283 1368 26315
rect 1408 26283 1440 26315
rect 1480 26283 1512 26315
rect 1552 26283 1584 26315
rect 1624 26283 1656 26315
rect 1696 26283 1728 26315
rect 1768 26283 1800 26315
rect 1840 26283 1872 26315
rect 1912 26283 1944 26315
rect 1984 26283 2016 26315
rect 2056 26283 2088 26315
rect 2128 26283 2160 26315
rect 2200 26283 2232 26315
rect 2272 26283 2304 26315
rect 2344 26283 2376 26315
rect 2416 26283 2448 26315
rect 2488 26283 2520 26315
rect 2560 26283 2592 26315
rect 2632 26283 2664 26315
rect 2704 26283 2736 26315
rect 2776 26283 2808 26315
rect 2848 26283 2880 26315
rect 2920 26283 2952 26315
rect 2992 26283 3024 26315
rect 3064 26283 3096 26315
rect 3136 26283 3168 26315
rect 3208 26283 3240 26315
rect 3280 26283 3312 26315
rect 3352 26283 3384 26315
rect 3424 26283 3456 26315
rect 3496 26283 3528 26315
rect 3568 26283 3600 26315
rect 3640 26283 3672 26315
rect 3712 26283 3744 26315
rect 3784 26283 3816 26315
rect 3856 26283 3888 26315
rect 112 26211 144 26243
rect 184 26211 216 26243
rect 256 26211 288 26243
rect 328 26211 360 26243
rect 400 26211 432 26243
rect 472 26211 504 26243
rect 544 26211 576 26243
rect 616 26211 648 26243
rect 688 26211 720 26243
rect 760 26211 792 26243
rect 832 26211 864 26243
rect 904 26211 936 26243
rect 976 26211 1008 26243
rect 1048 26211 1080 26243
rect 1120 26211 1152 26243
rect 1192 26211 1224 26243
rect 1264 26211 1296 26243
rect 1336 26211 1368 26243
rect 1408 26211 1440 26243
rect 1480 26211 1512 26243
rect 1552 26211 1584 26243
rect 1624 26211 1656 26243
rect 1696 26211 1728 26243
rect 1768 26211 1800 26243
rect 1840 26211 1872 26243
rect 1912 26211 1944 26243
rect 1984 26211 2016 26243
rect 2056 26211 2088 26243
rect 2128 26211 2160 26243
rect 2200 26211 2232 26243
rect 2272 26211 2304 26243
rect 2344 26211 2376 26243
rect 2416 26211 2448 26243
rect 2488 26211 2520 26243
rect 2560 26211 2592 26243
rect 2632 26211 2664 26243
rect 2704 26211 2736 26243
rect 2776 26211 2808 26243
rect 2848 26211 2880 26243
rect 2920 26211 2952 26243
rect 2992 26211 3024 26243
rect 3064 26211 3096 26243
rect 3136 26211 3168 26243
rect 3208 26211 3240 26243
rect 3280 26211 3312 26243
rect 3352 26211 3384 26243
rect 3424 26211 3456 26243
rect 3496 26211 3528 26243
rect 3568 26211 3600 26243
rect 3640 26211 3672 26243
rect 3712 26211 3744 26243
rect 3784 26211 3816 26243
rect 3856 26211 3888 26243
rect 112 26139 144 26171
rect 184 26139 216 26171
rect 256 26139 288 26171
rect 328 26139 360 26171
rect 400 26139 432 26171
rect 472 26139 504 26171
rect 544 26139 576 26171
rect 616 26139 648 26171
rect 688 26139 720 26171
rect 760 26139 792 26171
rect 832 26139 864 26171
rect 904 26139 936 26171
rect 976 26139 1008 26171
rect 1048 26139 1080 26171
rect 1120 26139 1152 26171
rect 1192 26139 1224 26171
rect 1264 26139 1296 26171
rect 1336 26139 1368 26171
rect 1408 26139 1440 26171
rect 1480 26139 1512 26171
rect 1552 26139 1584 26171
rect 1624 26139 1656 26171
rect 1696 26139 1728 26171
rect 1768 26139 1800 26171
rect 1840 26139 1872 26171
rect 1912 26139 1944 26171
rect 1984 26139 2016 26171
rect 2056 26139 2088 26171
rect 2128 26139 2160 26171
rect 2200 26139 2232 26171
rect 2272 26139 2304 26171
rect 2344 26139 2376 26171
rect 2416 26139 2448 26171
rect 2488 26139 2520 26171
rect 2560 26139 2592 26171
rect 2632 26139 2664 26171
rect 2704 26139 2736 26171
rect 2776 26139 2808 26171
rect 2848 26139 2880 26171
rect 2920 26139 2952 26171
rect 2992 26139 3024 26171
rect 3064 26139 3096 26171
rect 3136 26139 3168 26171
rect 3208 26139 3240 26171
rect 3280 26139 3312 26171
rect 3352 26139 3384 26171
rect 3424 26139 3456 26171
rect 3496 26139 3528 26171
rect 3568 26139 3600 26171
rect 3640 26139 3672 26171
rect 3712 26139 3744 26171
rect 3784 26139 3816 26171
rect 3856 26139 3888 26171
rect 112 26067 144 26099
rect 184 26067 216 26099
rect 256 26067 288 26099
rect 328 26067 360 26099
rect 400 26067 432 26099
rect 472 26067 504 26099
rect 544 26067 576 26099
rect 616 26067 648 26099
rect 688 26067 720 26099
rect 760 26067 792 26099
rect 832 26067 864 26099
rect 904 26067 936 26099
rect 976 26067 1008 26099
rect 1048 26067 1080 26099
rect 1120 26067 1152 26099
rect 1192 26067 1224 26099
rect 1264 26067 1296 26099
rect 1336 26067 1368 26099
rect 1408 26067 1440 26099
rect 1480 26067 1512 26099
rect 1552 26067 1584 26099
rect 1624 26067 1656 26099
rect 1696 26067 1728 26099
rect 1768 26067 1800 26099
rect 1840 26067 1872 26099
rect 1912 26067 1944 26099
rect 1984 26067 2016 26099
rect 2056 26067 2088 26099
rect 2128 26067 2160 26099
rect 2200 26067 2232 26099
rect 2272 26067 2304 26099
rect 2344 26067 2376 26099
rect 2416 26067 2448 26099
rect 2488 26067 2520 26099
rect 2560 26067 2592 26099
rect 2632 26067 2664 26099
rect 2704 26067 2736 26099
rect 2776 26067 2808 26099
rect 2848 26067 2880 26099
rect 2920 26067 2952 26099
rect 2992 26067 3024 26099
rect 3064 26067 3096 26099
rect 3136 26067 3168 26099
rect 3208 26067 3240 26099
rect 3280 26067 3312 26099
rect 3352 26067 3384 26099
rect 3424 26067 3456 26099
rect 3496 26067 3528 26099
rect 3568 26067 3600 26099
rect 3640 26067 3672 26099
rect 3712 26067 3744 26099
rect 3784 26067 3816 26099
rect 3856 26067 3888 26099
rect 112 25995 144 26027
rect 184 25995 216 26027
rect 256 25995 288 26027
rect 328 25995 360 26027
rect 400 25995 432 26027
rect 472 25995 504 26027
rect 544 25995 576 26027
rect 616 25995 648 26027
rect 688 25995 720 26027
rect 760 25995 792 26027
rect 832 25995 864 26027
rect 904 25995 936 26027
rect 976 25995 1008 26027
rect 1048 25995 1080 26027
rect 1120 25995 1152 26027
rect 1192 25995 1224 26027
rect 1264 25995 1296 26027
rect 1336 25995 1368 26027
rect 1408 25995 1440 26027
rect 1480 25995 1512 26027
rect 1552 25995 1584 26027
rect 1624 25995 1656 26027
rect 1696 25995 1728 26027
rect 1768 25995 1800 26027
rect 1840 25995 1872 26027
rect 1912 25995 1944 26027
rect 1984 25995 2016 26027
rect 2056 25995 2088 26027
rect 2128 25995 2160 26027
rect 2200 25995 2232 26027
rect 2272 25995 2304 26027
rect 2344 25995 2376 26027
rect 2416 25995 2448 26027
rect 2488 25995 2520 26027
rect 2560 25995 2592 26027
rect 2632 25995 2664 26027
rect 2704 25995 2736 26027
rect 2776 25995 2808 26027
rect 2848 25995 2880 26027
rect 2920 25995 2952 26027
rect 2992 25995 3024 26027
rect 3064 25995 3096 26027
rect 3136 25995 3168 26027
rect 3208 25995 3240 26027
rect 3280 25995 3312 26027
rect 3352 25995 3384 26027
rect 3424 25995 3456 26027
rect 3496 25995 3528 26027
rect 3568 25995 3600 26027
rect 3640 25995 3672 26027
rect 3712 25995 3744 26027
rect 3784 25995 3816 26027
rect 3856 25995 3888 26027
rect 112 25923 144 25955
rect 184 25923 216 25955
rect 256 25923 288 25955
rect 328 25923 360 25955
rect 400 25923 432 25955
rect 472 25923 504 25955
rect 544 25923 576 25955
rect 616 25923 648 25955
rect 688 25923 720 25955
rect 760 25923 792 25955
rect 832 25923 864 25955
rect 904 25923 936 25955
rect 976 25923 1008 25955
rect 1048 25923 1080 25955
rect 1120 25923 1152 25955
rect 1192 25923 1224 25955
rect 1264 25923 1296 25955
rect 1336 25923 1368 25955
rect 1408 25923 1440 25955
rect 1480 25923 1512 25955
rect 1552 25923 1584 25955
rect 1624 25923 1656 25955
rect 1696 25923 1728 25955
rect 1768 25923 1800 25955
rect 1840 25923 1872 25955
rect 1912 25923 1944 25955
rect 1984 25923 2016 25955
rect 2056 25923 2088 25955
rect 2128 25923 2160 25955
rect 2200 25923 2232 25955
rect 2272 25923 2304 25955
rect 2344 25923 2376 25955
rect 2416 25923 2448 25955
rect 2488 25923 2520 25955
rect 2560 25923 2592 25955
rect 2632 25923 2664 25955
rect 2704 25923 2736 25955
rect 2776 25923 2808 25955
rect 2848 25923 2880 25955
rect 2920 25923 2952 25955
rect 2992 25923 3024 25955
rect 3064 25923 3096 25955
rect 3136 25923 3168 25955
rect 3208 25923 3240 25955
rect 3280 25923 3312 25955
rect 3352 25923 3384 25955
rect 3424 25923 3456 25955
rect 3496 25923 3528 25955
rect 3568 25923 3600 25955
rect 3640 25923 3672 25955
rect 3712 25923 3744 25955
rect 3784 25923 3816 25955
rect 3856 25923 3888 25955
rect 112 25851 144 25883
rect 184 25851 216 25883
rect 256 25851 288 25883
rect 328 25851 360 25883
rect 400 25851 432 25883
rect 472 25851 504 25883
rect 544 25851 576 25883
rect 616 25851 648 25883
rect 688 25851 720 25883
rect 760 25851 792 25883
rect 832 25851 864 25883
rect 904 25851 936 25883
rect 976 25851 1008 25883
rect 1048 25851 1080 25883
rect 1120 25851 1152 25883
rect 1192 25851 1224 25883
rect 1264 25851 1296 25883
rect 1336 25851 1368 25883
rect 1408 25851 1440 25883
rect 1480 25851 1512 25883
rect 1552 25851 1584 25883
rect 1624 25851 1656 25883
rect 1696 25851 1728 25883
rect 1768 25851 1800 25883
rect 1840 25851 1872 25883
rect 1912 25851 1944 25883
rect 1984 25851 2016 25883
rect 2056 25851 2088 25883
rect 2128 25851 2160 25883
rect 2200 25851 2232 25883
rect 2272 25851 2304 25883
rect 2344 25851 2376 25883
rect 2416 25851 2448 25883
rect 2488 25851 2520 25883
rect 2560 25851 2592 25883
rect 2632 25851 2664 25883
rect 2704 25851 2736 25883
rect 2776 25851 2808 25883
rect 2848 25851 2880 25883
rect 2920 25851 2952 25883
rect 2992 25851 3024 25883
rect 3064 25851 3096 25883
rect 3136 25851 3168 25883
rect 3208 25851 3240 25883
rect 3280 25851 3312 25883
rect 3352 25851 3384 25883
rect 3424 25851 3456 25883
rect 3496 25851 3528 25883
rect 3568 25851 3600 25883
rect 3640 25851 3672 25883
rect 3712 25851 3744 25883
rect 3784 25851 3816 25883
rect 3856 25851 3888 25883
rect 112 25779 144 25811
rect 184 25779 216 25811
rect 256 25779 288 25811
rect 328 25779 360 25811
rect 400 25779 432 25811
rect 472 25779 504 25811
rect 544 25779 576 25811
rect 616 25779 648 25811
rect 688 25779 720 25811
rect 760 25779 792 25811
rect 832 25779 864 25811
rect 904 25779 936 25811
rect 976 25779 1008 25811
rect 1048 25779 1080 25811
rect 1120 25779 1152 25811
rect 1192 25779 1224 25811
rect 1264 25779 1296 25811
rect 1336 25779 1368 25811
rect 1408 25779 1440 25811
rect 1480 25779 1512 25811
rect 1552 25779 1584 25811
rect 1624 25779 1656 25811
rect 1696 25779 1728 25811
rect 1768 25779 1800 25811
rect 1840 25779 1872 25811
rect 1912 25779 1944 25811
rect 1984 25779 2016 25811
rect 2056 25779 2088 25811
rect 2128 25779 2160 25811
rect 2200 25779 2232 25811
rect 2272 25779 2304 25811
rect 2344 25779 2376 25811
rect 2416 25779 2448 25811
rect 2488 25779 2520 25811
rect 2560 25779 2592 25811
rect 2632 25779 2664 25811
rect 2704 25779 2736 25811
rect 2776 25779 2808 25811
rect 2848 25779 2880 25811
rect 2920 25779 2952 25811
rect 2992 25779 3024 25811
rect 3064 25779 3096 25811
rect 3136 25779 3168 25811
rect 3208 25779 3240 25811
rect 3280 25779 3312 25811
rect 3352 25779 3384 25811
rect 3424 25779 3456 25811
rect 3496 25779 3528 25811
rect 3568 25779 3600 25811
rect 3640 25779 3672 25811
rect 3712 25779 3744 25811
rect 3784 25779 3816 25811
rect 3856 25779 3888 25811
rect 112 25707 144 25739
rect 184 25707 216 25739
rect 256 25707 288 25739
rect 328 25707 360 25739
rect 400 25707 432 25739
rect 472 25707 504 25739
rect 544 25707 576 25739
rect 616 25707 648 25739
rect 688 25707 720 25739
rect 760 25707 792 25739
rect 832 25707 864 25739
rect 904 25707 936 25739
rect 976 25707 1008 25739
rect 1048 25707 1080 25739
rect 1120 25707 1152 25739
rect 1192 25707 1224 25739
rect 1264 25707 1296 25739
rect 1336 25707 1368 25739
rect 1408 25707 1440 25739
rect 1480 25707 1512 25739
rect 1552 25707 1584 25739
rect 1624 25707 1656 25739
rect 1696 25707 1728 25739
rect 1768 25707 1800 25739
rect 1840 25707 1872 25739
rect 1912 25707 1944 25739
rect 1984 25707 2016 25739
rect 2056 25707 2088 25739
rect 2128 25707 2160 25739
rect 2200 25707 2232 25739
rect 2272 25707 2304 25739
rect 2344 25707 2376 25739
rect 2416 25707 2448 25739
rect 2488 25707 2520 25739
rect 2560 25707 2592 25739
rect 2632 25707 2664 25739
rect 2704 25707 2736 25739
rect 2776 25707 2808 25739
rect 2848 25707 2880 25739
rect 2920 25707 2952 25739
rect 2992 25707 3024 25739
rect 3064 25707 3096 25739
rect 3136 25707 3168 25739
rect 3208 25707 3240 25739
rect 3280 25707 3312 25739
rect 3352 25707 3384 25739
rect 3424 25707 3456 25739
rect 3496 25707 3528 25739
rect 3568 25707 3600 25739
rect 3640 25707 3672 25739
rect 3712 25707 3744 25739
rect 3784 25707 3816 25739
rect 3856 25707 3888 25739
rect 112 25635 144 25667
rect 184 25635 216 25667
rect 256 25635 288 25667
rect 328 25635 360 25667
rect 400 25635 432 25667
rect 472 25635 504 25667
rect 544 25635 576 25667
rect 616 25635 648 25667
rect 688 25635 720 25667
rect 760 25635 792 25667
rect 832 25635 864 25667
rect 904 25635 936 25667
rect 976 25635 1008 25667
rect 1048 25635 1080 25667
rect 1120 25635 1152 25667
rect 1192 25635 1224 25667
rect 1264 25635 1296 25667
rect 1336 25635 1368 25667
rect 1408 25635 1440 25667
rect 1480 25635 1512 25667
rect 1552 25635 1584 25667
rect 1624 25635 1656 25667
rect 1696 25635 1728 25667
rect 1768 25635 1800 25667
rect 1840 25635 1872 25667
rect 1912 25635 1944 25667
rect 1984 25635 2016 25667
rect 2056 25635 2088 25667
rect 2128 25635 2160 25667
rect 2200 25635 2232 25667
rect 2272 25635 2304 25667
rect 2344 25635 2376 25667
rect 2416 25635 2448 25667
rect 2488 25635 2520 25667
rect 2560 25635 2592 25667
rect 2632 25635 2664 25667
rect 2704 25635 2736 25667
rect 2776 25635 2808 25667
rect 2848 25635 2880 25667
rect 2920 25635 2952 25667
rect 2992 25635 3024 25667
rect 3064 25635 3096 25667
rect 3136 25635 3168 25667
rect 3208 25635 3240 25667
rect 3280 25635 3312 25667
rect 3352 25635 3384 25667
rect 3424 25635 3456 25667
rect 3496 25635 3528 25667
rect 3568 25635 3600 25667
rect 3640 25635 3672 25667
rect 3712 25635 3744 25667
rect 3784 25635 3816 25667
rect 3856 25635 3888 25667
rect 112 25563 144 25595
rect 184 25563 216 25595
rect 256 25563 288 25595
rect 328 25563 360 25595
rect 400 25563 432 25595
rect 472 25563 504 25595
rect 544 25563 576 25595
rect 616 25563 648 25595
rect 688 25563 720 25595
rect 760 25563 792 25595
rect 832 25563 864 25595
rect 904 25563 936 25595
rect 976 25563 1008 25595
rect 1048 25563 1080 25595
rect 1120 25563 1152 25595
rect 1192 25563 1224 25595
rect 1264 25563 1296 25595
rect 1336 25563 1368 25595
rect 1408 25563 1440 25595
rect 1480 25563 1512 25595
rect 1552 25563 1584 25595
rect 1624 25563 1656 25595
rect 1696 25563 1728 25595
rect 1768 25563 1800 25595
rect 1840 25563 1872 25595
rect 1912 25563 1944 25595
rect 1984 25563 2016 25595
rect 2056 25563 2088 25595
rect 2128 25563 2160 25595
rect 2200 25563 2232 25595
rect 2272 25563 2304 25595
rect 2344 25563 2376 25595
rect 2416 25563 2448 25595
rect 2488 25563 2520 25595
rect 2560 25563 2592 25595
rect 2632 25563 2664 25595
rect 2704 25563 2736 25595
rect 2776 25563 2808 25595
rect 2848 25563 2880 25595
rect 2920 25563 2952 25595
rect 2992 25563 3024 25595
rect 3064 25563 3096 25595
rect 3136 25563 3168 25595
rect 3208 25563 3240 25595
rect 3280 25563 3312 25595
rect 3352 25563 3384 25595
rect 3424 25563 3456 25595
rect 3496 25563 3528 25595
rect 3568 25563 3600 25595
rect 3640 25563 3672 25595
rect 3712 25563 3744 25595
rect 3784 25563 3816 25595
rect 3856 25563 3888 25595
rect 112 25491 144 25523
rect 184 25491 216 25523
rect 256 25491 288 25523
rect 328 25491 360 25523
rect 400 25491 432 25523
rect 472 25491 504 25523
rect 544 25491 576 25523
rect 616 25491 648 25523
rect 688 25491 720 25523
rect 760 25491 792 25523
rect 832 25491 864 25523
rect 904 25491 936 25523
rect 976 25491 1008 25523
rect 1048 25491 1080 25523
rect 1120 25491 1152 25523
rect 1192 25491 1224 25523
rect 1264 25491 1296 25523
rect 1336 25491 1368 25523
rect 1408 25491 1440 25523
rect 1480 25491 1512 25523
rect 1552 25491 1584 25523
rect 1624 25491 1656 25523
rect 1696 25491 1728 25523
rect 1768 25491 1800 25523
rect 1840 25491 1872 25523
rect 1912 25491 1944 25523
rect 1984 25491 2016 25523
rect 2056 25491 2088 25523
rect 2128 25491 2160 25523
rect 2200 25491 2232 25523
rect 2272 25491 2304 25523
rect 2344 25491 2376 25523
rect 2416 25491 2448 25523
rect 2488 25491 2520 25523
rect 2560 25491 2592 25523
rect 2632 25491 2664 25523
rect 2704 25491 2736 25523
rect 2776 25491 2808 25523
rect 2848 25491 2880 25523
rect 2920 25491 2952 25523
rect 2992 25491 3024 25523
rect 3064 25491 3096 25523
rect 3136 25491 3168 25523
rect 3208 25491 3240 25523
rect 3280 25491 3312 25523
rect 3352 25491 3384 25523
rect 3424 25491 3456 25523
rect 3496 25491 3528 25523
rect 3568 25491 3600 25523
rect 3640 25491 3672 25523
rect 3712 25491 3744 25523
rect 3784 25491 3816 25523
rect 3856 25491 3888 25523
rect 112 25419 144 25451
rect 184 25419 216 25451
rect 256 25419 288 25451
rect 328 25419 360 25451
rect 400 25419 432 25451
rect 472 25419 504 25451
rect 544 25419 576 25451
rect 616 25419 648 25451
rect 688 25419 720 25451
rect 760 25419 792 25451
rect 832 25419 864 25451
rect 904 25419 936 25451
rect 976 25419 1008 25451
rect 1048 25419 1080 25451
rect 1120 25419 1152 25451
rect 1192 25419 1224 25451
rect 1264 25419 1296 25451
rect 1336 25419 1368 25451
rect 1408 25419 1440 25451
rect 1480 25419 1512 25451
rect 1552 25419 1584 25451
rect 1624 25419 1656 25451
rect 1696 25419 1728 25451
rect 1768 25419 1800 25451
rect 1840 25419 1872 25451
rect 1912 25419 1944 25451
rect 1984 25419 2016 25451
rect 2056 25419 2088 25451
rect 2128 25419 2160 25451
rect 2200 25419 2232 25451
rect 2272 25419 2304 25451
rect 2344 25419 2376 25451
rect 2416 25419 2448 25451
rect 2488 25419 2520 25451
rect 2560 25419 2592 25451
rect 2632 25419 2664 25451
rect 2704 25419 2736 25451
rect 2776 25419 2808 25451
rect 2848 25419 2880 25451
rect 2920 25419 2952 25451
rect 2992 25419 3024 25451
rect 3064 25419 3096 25451
rect 3136 25419 3168 25451
rect 3208 25419 3240 25451
rect 3280 25419 3312 25451
rect 3352 25419 3384 25451
rect 3424 25419 3456 25451
rect 3496 25419 3528 25451
rect 3568 25419 3600 25451
rect 3640 25419 3672 25451
rect 3712 25419 3744 25451
rect 3784 25419 3816 25451
rect 3856 25419 3888 25451
rect 112 25347 144 25379
rect 184 25347 216 25379
rect 256 25347 288 25379
rect 328 25347 360 25379
rect 400 25347 432 25379
rect 472 25347 504 25379
rect 544 25347 576 25379
rect 616 25347 648 25379
rect 688 25347 720 25379
rect 760 25347 792 25379
rect 832 25347 864 25379
rect 904 25347 936 25379
rect 976 25347 1008 25379
rect 1048 25347 1080 25379
rect 1120 25347 1152 25379
rect 1192 25347 1224 25379
rect 1264 25347 1296 25379
rect 1336 25347 1368 25379
rect 1408 25347 1440 25379
rect 1480 25347 1512 25379
rect 1552 25347 1584 25379
rect 1624 25347 1656 25379
rect 1696 25347 1728 25379
rect 1768 25347 1800 25379
rect 1840 25347 1872 25379
rect 1912 25347 1944 25379
rect 1984 25347 2016 25379
rect 2056 25347 2088 25379
rect 2128 25347 2160 25379
rect 2200 25347 2232 25379
rect 2272 25347 2304 25379
rect 2344 25347 2376 25379
rect 2416 25347 2448 25379
rect 2488 25347 2520 25379
rect 2560 25347 2592 25379
rect 2632 25347 2664 25379
rect 2704 25347 2736 25379
rect 2776 25347 2808 25379
rect 2848 25347 2880 25379
rect 2920 25347 2952 25379
rect 2992 25347 3024 25379
rect 3064 25347 3096 25379
rect 3136 25347 3168 25379
rect 3208 25347 3240 25379
rect 3280 25347 3312 25379
rect 3352 25347 3384 25379
rect 3424 25347 3456 25379
rect 3496 25347 3528 25379
rect 3568 25347 3600 25379
rect 3640 25347 3672 25379
rect 3712 25347 3744 25379
rect 3784 25347 3816 25379
rect 3856 25347 3888 25379
rect 112 25275 144 25307
rect 184 25275 216 25307
rect 256 25275 288 25307
rect 328 25275 360 25307
rect 400 25275 432 25307
rect 472 25275 504 25307
rect 544 25275 576 25307
rect 616 25275 648 25307
rect 688 25275 720 25307
rect 760 25275 792 25307
rect 832 25275 864 25307
rect 904 25275 936 25307
rect 976 25275 1008 25307
rect 1048 25275 1080 25307
rect 1120 25275 1152 25307
rect 1192 25275 1224 25307
rect 1264 25275 1296 25307
rect 1336 25275 1368 25307
rect 1408 25275 1440 25307
rect 1480 25275 1512 25307
rect 1552 25275 1584 25307
rect 1624 25275 1656 25307
rect 1696 25275 1728 25307
rect 1768 25275 1800 25307
rect 1840 25275 1872 25307
rect 1912 25275 1944 25307
rect 1984 25275 2016 25307
rect 2056 25275 2088 25307
rect 2128 25275 2160 25307
rect 2200 25275 2232 25307
rect 2272 25275 2304 25307
rect 2344 25275 2376 25307
rect 2416 25275 2448 25307
rect 2488 25275 2520 25307
rect 2560 25275 2592 25307
rect 2632 25275 2664 25307
rect 2704 25275 2736 25307
rect 2776 25275 2808 25307
rect 2848 25275 2880 25307
rect 2920 25275 2952 25307
rect 2992 25275 3024 25307
rect 3064 25275 3096 25307
rect 3136 25275 3168 25307
rect 3208 25275 3240 25307
rect 3280 25275 3312 25307
rect 3352 25275 3384 25307
rect 3424 25275 3456 25307
rect 3496 25275 3528 25307
rect 3568 25275 3600 25307
rect 3640 25275 3672 25307
rect 3712 25275 3744 25307
rect 3784 25275 3816 25307
rect 3856 25275 3888 25307
rect 112 25203 144 25235
rect 184 25203 216 25235
rect 256 25203 288 25235
rect 328 25203 360 25235
rect 400 25203 432 25235
rect 472 25203 504 25235
rect 544 25203 576 25235
rect 616 25203 648 25235
rect 688 25203 720 25235
rect 760 25203 792 25235
rect 832 25203 864 25235
rect 904 25203 936 25235
rect 976 25203 1008 25235
rect 1048 25203 1080 25235
rect 1120 25203 1152 25235
rect 1192 25203 1224 25235
rect 1264 25203 1296 25235
rect 1336 25203 1368 25235
rect 1408 25203 1440 25235
rect 1480 25203 1512 25235
rect 1552 25203 1584 25235
rect 1624 25203 1656 25235
rect 1696 25203 1728 25235
rect 1768 25203 1800 25235
rect 1840 25203 1872 25235
rect 1912 25203 1944 25235
rect 1984 25203 2016 25235
rect 2056 25203 2088 25235
rect 2128 25203 2160 25235
rect 2200 25203 2232 25235
rect 2272 25203 2304 25235
rect 2344 25203 2376 25235
rect 2416 25203 2448 25235
rect 2488 25203 2520 25235
rect 2560 25203 2592 25235
rect 2632 25203 2664 25235
rect 2704 25203 2736 25235
rect 2776 25203 2808 25235
rect 2848 25203 2880 25235
rect 2920 25203 2952 25235
rect 2992 25203 3024 25235
rect 3064 25203 3096 25235
rect 3136 25203 3168 25235
rect 3208 25203 3240 25235
rect 3280 25203 3312 25235
rect 3352 25203 3384 25235
rect 3424 25203 3456 25235
rect 3496 25203 3528 25235
rect 3568 25203 3600 25235
rect 3640 25203 3672 25235
rect 3712 25203 3744 25235
rect 3784 25203 3816 25235
rect 3856 25203 3888 25235
rect 112 25131 144 25163
rect 184 25131 216 25163
rect 256 25131 288 25163
rect 328 25131 360 25163
rect 400 25131 432 25163
rect 472 25131 504 25163
rect 544 25131 576 25163
rect 616 25131 648 25163
rect 688 25131 720 25163
rect 760 25131 792 25163
rect 832 25131 864 25163
rect 904 25131 936 25163
rect 976 25131 1008 25163
rect 1048 25131 1080 25163
rect 1120 25131 1152 25163
rect 1192 25131 1224 25163
rect 1264 25131 1296 25163
rect 1336 25131 1368 25163
rect 1408 25131 1440 25163
rect 1480 25131 1512 25163
rect 1552 25131 1584 25163
rect 1624 25131 1656 25163
rect 1696 25131 1728 25163
rect 1768 25131 1800 25163
rect 1840 25131 1872 25163
rect 1912 25131 1944 25163
rect 1984 25131 2016 25163
rect 2056 25131 2088 25163
rect 2128 25131 2160 25163
rect 2200 25131 2232 25163
rect 2272 25131 2304 25163
rect 2344 25131 2376 25163
rect 2416 25131 2448 25163
rect 2488 25131 2520 25163
rect 2560 25131 2592 25163
rect 2632 25131 2664 25163
rect 2704 25131 2736 25163
rect 2776 25131 2808 25163
rect 2848 25131 2880 25163
rect 2920 25131 2952 25163
rect 2992 25131 3024 25163
rect 3064 25131 3096 25163
rect 3136 25131 3168 25163
rect 3208 25131 3240 25163
rect 3280 25131 3312 25163
rect 3352 25131 3384 25163
rect 3424 25131 3456 25163
rect 3496 25131 3528 25163
rect 3568 25131 3600 25163
rect 3640 25131 3672 25163
rect 3712 25131 3744 25163
rect 3784 25131 3816 25163
rect 3856 25131 3888 25163
rect 112 25059 144 25091
rect 184 25059 216 25091
rect 256 25059 288 25091
rect 328 25059 360 25091
rect 400 25059 432 25091
rect 472 25059 504 25091
rect 544 25059 576 25091
rect 616 25059 648 25091
rect 688 25059 720 25091
rect 760 25059 792 25091
rect 832 25059 864 25091
rect 904 25059 936 25091
rect 976 25059 1008 25091
rect 1048 25059 1080 25091
rect 1120 25059 1152 25091
rect 1192 25059 1224 25091
rect 1264 25059 1296 25091
rect 1336 25059 1368 25091
rect 1408 25059 1440 25091
rect 1480 25059 1512 25091
rect 1552 25059 1584 25091
rect 1624 25059 1656 25091
rect 1696 25059 1728 25091
rect 1768 25059 1800 25091
rect 1840 25059 1872 25091
rect 1912 25059 1944 25091
rect 1984 25059 2016 25091
rect 2056 25059 2088 25091
rect 2128 25059 2160 25091
rect 2200 25059 2232 25091
rect 2272 25059 2304 25091
rect 2344 25059 2376 25091
rect 2416 25059 2448 25091
rect 2488 25059 2520 25091
rect 2560 25059 2592 25091
rect 2632 25059 2664 25091
rect 2704 25059 2736 25091
rect 2776 25059 2808 25091
rect 2848 25059 2880 25091
rect 2920 25059 2952 25091
rect 2992 25059 3024 25091
rect 3064 25059 3096 25091
rect 3136 25059 3168 25091
rect 3208 25059 3240 25091
rect 3280 25059 3312 25091
rect 3352 25059 3384 25091
rect 3424 25059 3456 25091
rect 3496 25059 3528 25091
rect 3568 25059 3600 25091
rect 3640 25059 3672 25091
rect 3712 25059 3744 25091
rect 3784 25059 3816 25091
rect 3856 25059 3888 25091
rect 112 24987 144 25019
rect 184 24987 216 25019
rect 256 24987 288 25019
rect 328 24987 360 25019
rect 400 24987 432 25019
rect 472 24987 504 25019
rect 544 24987 576 25019
rect 616 24987 648 25019
rect 688 24987 720 25019
rect 760 24987 792 25019
rect 832 24987 864 25019
rect 904 24987 936 25019
rect 976 24987 1008 25019
rect 1048 24987 1080 25019
rect 1120 24987 1152 25019
rect 1192 24987 1224 25019
rect 1264 24987 1296 25019
rect 1336 24987 1368 25019
rect 1408 24987 1440 25019
rect 1480 24987 1512 25019
rect 1552 24987 1584 25019
rect 1624 24987 1656 25019
rect 1696 24987 1728 25019
rect 1768 24987 1800 25019
rect 1840 24987 1872 25019
rect 1912 24987 1944 25019
rect 1984 24987 2016 25019
rect 2056 24987 2088 25019
rect 2128 24987 2160 25019
rect 2200 24987 2232 25019
rect 2272 24987 2304 25019
rect 2344 24987 2376 25019
rect 2416 24987 2448 25019
rect 2488 24987 2520 25019
rect 2560 24987 2592 25019
rect 2632 24987 2664 25019
rect 2704 24987 2736 25019
rect 2776 24987 2808 25019
rect 2848 24987 2880 25019
rect 2920 24987 2952 25019
rect 2992 24987 3024 25019
rect 3064 24987 3096 25019
rect 3136 24987 3168 25019
rect 3208 24987 3240 25019
rect 3280 24987 3312 25019
rect 3352 24987 3384 25019
rect 3424 24987 3456 25019
rect 3496 24987 3528 25019
rect 3568 24987 3600 25019
rect 3640 24987 3672 25019
rect 3712 24987 3744 25019
rect 3784 24987 3816 25019
rect 3856 24987 3888 25019
rect 112 24915 144 24947
rect 184 24915 216 24947
rect 256 24915 288 24947
rect 328 24915 360 24947
rect 400 24915 432 24947
rect 472 24915 504 24947
rect 544 24915 576 24947
rect 616 24915 648 24947
rect 688 24915 720 24947
rect 760 24915 792 24947
rect 832 24915 864 24947
rect 904 24915 936 24947
rect 976 24915 1008 24947
rect 1048 24915 1080 24947
rect 1120 24915 1152 24947
rect 1192 24915 1224 24947
rect 1264 24915 1296 24947
rect 1336 24915 1368 24947
rect 1408 24915 1440 24947
rect 1480 24915 1512 24947
rect 1552 24915 1584 24947
rect 1624 24915 1656 24947
rect 1696 24915 1728 24947
rect 1768 24915 1800 24947
rect 1840 24915 1872 24947
rect 1912 24915 1944 24947
rect 1984 24915 2016 24947
rect 2056 24915 2088 24947
rect 2128 24915 2160 24947
rect 2200 24915 2232 24947
rect 2272 24915 2304 24947
rect 2344 24915 2376 24947
rect 2416 24915 2448 24947
rect 2488 24915 2520 24947
rect 2560 24915 2592 24947
rect 2632 24915 2664 24947
rect 2704 24915 2736 24947
rect 2776 24915 2808 24947
rect 2848 24915 2880 24947
rect 2920 24915 2952 24947
rect 2992 24915 3024 24947
rect 3064 24915 3096 24947
rect 3136 24915 3168 24947
rect 3208 24915 3240 24947
rect 3280 24915 3312 24947
rect 3352 24915 3384 24947
rect 3424 24915 3456 24947
rect 3496 24915 3528 24947
rect 3568 24915 3600 24947
rect 3640 24915 3672 24947
rect 3712 24915 3744 24947
rect 3784 24915 3816 24947
rect 3856 24915 3888 24947
rect 112 24843 144 24875
rect 184 24843 216 24875
rect 256 24843 288 24875
rect 328 24843 360 24875
rect 400 24843 432 24875
rect 472 24843 504 24875
rect 544 24843 576 24875
rect 616 24843 648 24875
rect 688 24843 720 24875
rect 760 24843 792 24875
rect 832 24843 864 24875
rect 904 24843 936 24875
rect 976 24843 1008 24875
rect 1048 24843 1080 24875
rect 1120 24843 1152 24875
rect 1192 24843 1224 24875
rect 1264 24843 1296 24875
rect 1336 24843 1368 24875
rect 1408 24843 1440 24875
rect 1480 24843 1512 24875
rect 1552 24843 1584 24875
rect 1624 24843 1656 24875
rect 1696 24843 1728 24875
rect 1768 24843 1800 24875
rect 1840 24843 1872 24875
rect 1912 24843 1944 24875
rect 1984 24843 2016 24875
rect 2056 24843 2088 24875
rect 2128 24843 2160 24875
rect 2200 24843 2232 24875
rect 2272 24843 2304 24875
rect 2344 24843 2376 24875
rect 2416 24843 2448 24875
rect 2488 24843 2520 24875
rect 2560 24843 2592 24875
rect 2632 24843 2664 24875
rect 2704 24843 2736 24875
rect 2776 24843 2808 24875
rect 2848 24843 2880 24875
rect 2920 24843 2952 24875
rect 2992 24843 3024 24875
rect 3064 24843 3096 24875
rect 3136 24843 3168 24875
rect 3208 24843 3240 24875
rect 3280 24843 3312 24875
rect 3352 24843 3384 24875
rect 3424 24843 3456 24875
rect 3496 24843 3528 24875
rect 3568 24843 3600 24875
rect 3640 24843 3672 24875
rect 3712 24843 3744 24875
rect 3784 24843 3816 24875
rect 3856 24843 3888 24875
rect 112 24771 144 24803
rect 184 24771 216 24803
rect 256 24771 288 24803
rect 328 24771 360 24803
rect 400 24771 432 24803
rect 472 24771 504 24803
rect 544 24771 576 24803
rect 616 24771 648 24803
rect 688 24771 720 24803
rect 760 24771 792 24803
rect 832 24771 864 24803
rect 904 24771 936 24803
rect 976 24771 1008 24803
rect 1048 24771 1080 24803
rect 1120 24771 1152 24803
rect 1192 24771 1224 24803
rect 1264 24771 1296 24803
rect 1336 24771 1368 24803
rect 1408 24771 1440 24803
rect 1480 24771 1512 24803
rect 1552 24771 1584 24803
rect 1624 24771 1656 24803
rect 1696 24771 1728 24803
rect 1768 24771 1800 24803
rect 1840 24771 1872 24803
rect 1912 24771 1944 24803
rect 1984 24771 2016 24803
rect 2056 24771 2088 24803
rect 2128 24771 2160 24803
rect 2200 24771 2232 24803
rect 2272 24771 2304 24803
rect 2344 24771 2376 24803
rect 2416 24771 2448 24803
rect 2488 24771 2520 24803
rect 2560 24771 2592 24803
rect 2632 24771 2664 24803
rect 2704 24771 2736 24803
rect 2776 24771 2808 24803
rect 2848 24771 2880 24803
rect 2920 24771 2952 24803
rect 2992 24771 3024 24803
rect 3064 24771 3096 24803
rect 3136 24771 3168 24803
rect 3208 24771 3240 24803
rect 3280 24771 3312 24803
rect 3352 24771 3384 24803
rect 3424 24771 3456 24803
rect 3496 24771 3528 24803
rect 3568 24771 3600 24803
rect 3640 24771 3672 24803
rect 3712 24771 3744 24803
rect 3784 24771 3816 24803
rect 3856 24771 3888 24803
rect 112 24699 144 24731
rect 184 24699 216 24731
rect 256 24699 288 24731
rect 328 24699 360 24731
rect 400 24699 432 24731
rect 472 24699 504 24731
rect 544 24699 576 24731
rect 616 24699 648 24731
rect 688 24699 720 24731
rect 760 24699 792 24731
rect 832 24699 864 24731
rect 904 24699 936 24731
rect 976 24699 1008 24731
rect 1048 24699 1080 24731
rect 1120 24699 1152 24731
rect 1192 24699 1224 24731
rect 1264 24699 1296 24731
rect 1336 24699 1368 24731
rect 1408 24699 1440 24731
rect 1480 24699 1512 24731
rect 1552 24699 1584 24731
rect 1624 24699 1656 24731
rect 1696 24699 1728 24731
rect 1768 24699 1800 24731
rect 1840 24699 1872 24731
rect 1912 24699 1944 24731
rect 1984 24699 2016 24731
rect 2056 24699 2088 24731
rect 2128 24699 2160 24731
rect 2200 24699 2232 24731
rect 2272 24699 2304 24731
rect 2344 24699 2376 24731
rect 2416 24699 2448 24731
rect 2488 24699 2520 24731
rect 2560 24699 2592 24731
rect 2632 24699 2664 24731
rect 2704 24699 2736 24731
rect 2776 24699 2808 24731
rect 2848 24699 2880 24731
rect 2920 24699 2952 24731
rect 2992 24699 3024 24731
rect 3064 24699 3096 24731
rect 3136 24699 3168 24731
rect 3208 24699 3240 24731
rect 3280 24699 3312 24731
rect 3352 24699 3384 24731
rect 3424 24699 3456 24731
rect 3496 24699 3528 24731
rect 3568 24699 3600 24731
rect 3640 24699 3672 24731
rect 3712 24699 3744 24731
rect 3784 24699 3816 24731
rect 3856 24699 3888 24731
rect 112 24627 144 24659
rect 184 24627 216 24659
rect 256 24627 288 24659
rect 328 24627 360 24659
rect 400 24627 432 24659
rect 472 24627 504 24659
rect 544 24627 576 24659
rect 616 24627 648 24659
rect 688 24627 720 24659
rect 760 24627 792 24659
rect 832 24627 864 24659
rect 904 24627 936 24659
rect 976 24627 1008 24659
rect 1048 24627 1080 24659
rect 1120 24627 1152 24659
rect 1192 24627 1224 24659
rect 1264 24627 1296 24659
rect 1336 24627 1368 24659
rect 1408 24627 1440 24659
rect 1480 24627 1512 24659
rect 1552 24627 1584 24659
rect 1624 24627 1656 24659
rect 1696 24627 1728 24659
rect 1768 24627 1800 24659
rect 1840 24627 1872 24659
rect 1912 24627 1944 24659
rect 1984 24627 2016 24659
rect 2056 24627 2088 24659
rect 2128 24627 2160 24659
rect 2200 24627 2232 24659
rect 2272 24627 2304 24659
rect 2344 24627 2376 24659
rect 2416 24627 2448 24659
rect 2488 24627 2520 24659
rect 2560 24627 2592 24659
rect 2632 24627 2664 24659
rect 2704 24627 2736 24659
rect 2776 24627 2808 24659
rect 2848 24627 2880 24659
rect 2920 24627 2952 24659
rect 2992 24627 3024 24659
rect 3064 24627 3096 24659
rect 3136 24627 3168 24659
rect 3208 24627 3240 24659
rect 3280 24627 3312 24659
rect 3352 24627 3384 24659
rect 3424 24627 3456 24659
rect 3496 24627 3528 24659
rect 3568 24627 3600 24659
rect 3640 24627 3672 24659
rect 3712 24627 3744 24659
rect 3784 24627 3816 24659
rect 3856 24627 3888 24659
rect 112 24555 144 24587
rect 184 24555 216 24587
rect 256 24555 288 24587
rect 328 24555 360 24587
rect 400 24555 432 24587
rect 472 24555 504 24587
rect 544 24555 576 24587
rect 616 24555 648 24587
rect 688 24555 720 24587
rect 760 24555 792 24587
rect 832 24555 864 24587
rect 904 24555 936 24587
rect 976 24555 1008 24587
rect 1048 24555 1080 24587
rect 1120 24555 1152 24587
rect 1192 24555 1224 24587
rect 1264 24555 1296 24587
rect 1336 24555 1368 24587
rect 1408 24555 1440 24587
rect 1480 24555 1512 24587
rect 1552 24555 1584 24587
rect 1624 24555 1656 24587
rect 1696 24555 1728 24587
rect 1768 24555 1800 24587
rect 1840 24555 1872 24587
rect 1912 24555 1944 24587
rect 1984 24555 2016 24587
rect 2056 24555 2088 24587
rect 2128 24555 2160 24587
rect 2200 24555 2232 24587
rect 2272 24555 2304 24587
rect 2344 24555 2376 24587
rect 2416 24555 2448 24587
rect 2488 24555 2520 24587
rect 2560 24555 2592 24587
rect 2632 24555 2664 24587
rect 2704 24555 2736 24587
rect 2776 24555 2808 24587
rect 2848 24555 2880 24587
rect 2920 24555 2952 24587
rect 2992 24555 3024 24587
rect 3064 24555 3096 24587
rect 3136 24555 3168 24587
rect 3208 24555 3240 24587
rect 3280 24555 3312 24587
rect 3352 24555 3384 24587
rect 3424 24555 3456 24587
rect 3496 24555 3528 24587
rect 3568 24555 3600 24587
rect 3640 24555 3672 24587
rect 3712 24555 3744 24587
rect 3784 24555 3816 24587
rect 3856 24555 3888 24587
rect 112 24483 144 24515
rect 184 24483 216 24515
rect 256 24483 288 24515
rect 328 24483 360 24515
rect 400 24483 432 24515
rect 472 24483 504 24515
rect 544 24483 576 24515
rect 616 24483 648 24515
rect 688 24483 720 24515
rect 760 24483 792 24515
rect 832 24483 864 24515
rect 904 24483 936 24515
rect 976 24483 1008 24515
rect 1048 24483 1080 24515
rect 1120 24483 1152 24515
rect 1192 24483 1224 24515
rect 1264 24483 1296 24515
rect 1336 24483 1368 24515
rect 1408 24483 1440 24515
rect 1480 24483 1512 24515
rect 1552 24483 1584 24515
rect 1624 24483 1656 24515
rect 1696 24483 1728 24515
rect 1768 24483 1800 24515
rect 1840 24483 1872 24515
rect 1912 24483 1944 24515
rect 1984 24483 2016 24515
rect 2056 24483 2088 24515
rect 2128 24483 2160 24515
rect 2200 24483 2232 24515
rect 2272 24483 2304 24515
rect 2344 24483 2376 24515
rect 2416 24483 2448 24515
rect 2488 24483 2520 24515
rect 2560 24483 2592 24515
rect 2632 24483 2664 24515
rect 2704 24483 2736 24515
rect 2776 24483 2808 24515
rect 2848 24483 2880 24515
rect 2920 24483 2952 24515
rect 2992 24483 3024 24515
rect 3064 24483 3096 24515
rect 3136 24483 3168 24515
rect 3208 24483 3240 24515
rect 3280 24483 3312 24515
rect 3352 24483 3384 24515
rect 3424 24483 3456 24515
rect 3496 24483 3528 24515
rect 3568 24483 3600 24515
rect 3640 24483 3672 24515
rect 3712 24483 3744 24515
rect 3784 24483 3816 24515
rect 3856 24483 3888 24515
rect 112 24411 144 24443
rect 184 24411 216 24443
rect 256 24411 288 24443
rect 328 24411 360 24443
rect 400 24411 432 24443
rect 472 24411 504 24443
rect 544 24411 576 24443
rect 616 24411 648 24443
rect 688 24411 720 24443
rect 760 24411 792 24443
rect 832 24411 864 24443
rect 904 24411 936 24443
rect 976 24411 1008 24443
rect 1048 24411 1080 24443
rect 1120 24411 1152 24443
rect 1192 24411 1224 24443
rect 1264 24411 1296 24443
rect 1336 24411 1368 24443
rect 1408 24411 1440 24443
rect 1480 24411 1512 24443
rect 1552 24411 1584 24443
rect 1624 24411 1656 24443
rect 1696 24411 1728 24443
rect 1768 24411 1800 24443
rect 1840 24411 1872 24443
rect 1912 24411 1944 24443
rect 1984 24411 2016 24443
rect 2056 24411 2088 24443
rect 2128 24411 2160 24443
rect 2200 24411 2232 24443
rect 2272 24411 2304 24443
rect 2344 24411 2376 24443
rect 2416 24411 2448 24443
rect 2488 24411 2520 24443
rect 2560 24411 2592 24443
rect 2632 24411 2664 24443
rect 2704 24411 2736 24443
rect 2776 24411 2808 24443
rect 2848 24411 2880 24443
rect 2920 24411 2952 24443
rect 2992 24411 3024 24443
rect 3064 24411 3096 24443
rect 3136 24411 3168 24443
rect 3208 24411 3240 24443
rect 3280 24411 3312 24443
rect 3352 24411 3384 24443
rect 3424 24411 3456 24443
rect 3496 24411 3528 24443
rect 3568 24411 3600 24443
rect 3640 24411 3672 24443
rect 3712 24411 3744 24443
rect 3784 24411 3816 24443
rect 3856 24411 3888 24443
rect 112 24339 144 24371
rect 184 24339 216 24371
rect 256 24339 288 24371
rect 328 24339 360 24371
rect 400 24339 432 24371
rect 472 24339 504 24371
rect 544 24339 576 24371
rect 616 24339 648 24371
rect 688 24339 720 24371
rect 760 24339 792 24371
rect 832 24339 864 24371
rect 904 24339 936 24371
rect 976 24339 1008 24371
rect 1048 24339 1080 24371
rect 1120 24339 1152 24371
rect 1192 24339 1224 24371
rect 1264 24339 1296 24371
rect 1336 24339 1368 24371
rect 1408 24339 1440 24371
rect 1480 24339 1512 24371
rect 1552 24339 1584 24371
rect 1624 24339 1656 24371
rect 1696 24339 1728 24371
rect 1768 24339 1800 24371
rect 1840 24339 1872 24371
rect 1912 24339 1944 24371
rect 1984 24339 2016 24371
rect 2056 24339 2088 24371
rect 2128 24339 2160 24371
rect 2200 24339 2232 24371
rect 2272 24339 2304 24371
rect 2344 24339 2376 24371
rect 2416 24339 2448 24371
rect 2488 24339 2520 24371
rect 2560 24339 2592 24371
rect 2632 24339 2664 24371
rect 2704 24339 2736 24371
rect 2776 24339 2808 24371
rect 2848 24339 2880 24371
rect 2920 24339 2952 24371
rect 2992 24339 3024 24371
rect 3064 24339 3096 24371
rect 3136 24339 3168 24371
rect 3208 24339 3240 24371
rect 3280 24339 3312 24371
rect 3352 24339 3384 24371
rect 3424 24339 3456 24371
rect 3496 24339 3528 24371
rect 3568 24339 3600 24371
rect 3640 24339 3672 24371
rect 3712 24339 3744 24371
rect 3784 24339 3816 24371
rect 3856 24339 3888 24371
rect 112 24267 144 24299
rect 184 24267 216 24299
rect 256 24267 288 24299
rect 328 24267 360 24299
rect 400 24267 432 24299
rect 472 24267 504 24299
rect 544 24267 576 24299
rect 616 24267 648 24299
rect 688 24267 720 24299
rect 760 24267 792 24299
rect 832 24267 864 24299
rect 904 24267 936 24299
rect 976 24267 1008 24299
rect 1048 24267 1080 24299
rect 1120 24267 1152 24299
rect 1192 24267 1224 24299
rect 1264 24267 1296 24299
rect 1336 24267 1368 24299
rect 1408 24267 1440 24299
rect 1480 24267 1512 24299
rect 1552 24267 1584 24299
rect 1624 24267 1656 24299
rect 1696 24267 1728 24299
rect 1768 24267 1800 24299
rect 1840 24267 1872 24299
rect 1912 24267 1944 24299
rect 1984 24267 2016 24299
rect 2056 24267 2088 24299
rect 2128 24267 2160 24299
rect 2200 24267 2232 24299
rect 2272 24267 2304 24299
rect 2344 24267 2376 24299
rect 2416 24267 2448 24299
rect 2488 24267 2520 24299
rect 2560 24267 2592 24299
rect 2632 24267 2664 24299
rect 2704 24267 2736 24299
rect 2776 24267 2808 24299
rect 2848 24267 2880 24299
rect 2920 24267 2952 24299
rect 2992 24267 3024 24299
rect 3064 24267 3096 24299
rect 3136 24267 3168 24299
rect 3208 24267 3240 24299
rect 3280 24267 3312 24299
rect 3352 24267 3384 24299
rect 3424 24267 3456 24299
rect 3496 24267 3528 24299
rect 3568 24267 3600 24299
rect 3640 24267 3672 24299
rect 3712 24267 3744 24299
rect 3784 24267 3816 24299
rect 3856 24267 3888 24299
rect 112 24195 144 24227
rect 184 24195 216 24227
rect 256 24195 288 24227
rect 328 24195 360 24227
rect 400 24195 432 24227
rect 472 24195 504 24227
rect 544 24195 576 24227
rect 616 24195 648 24227
rect 688 24195 720 24227
rect 760 24195 792 24227
rect 832 24195 864 24227
rect 904 24195 936 24227
rect 976 24195 1008 24227
rect 1048 24195 1080 24227
rect 1120 24195 1152 24227
rect 1192 24195 1224 24227
rect 1264 24195 1296 24227
rect 1336 24195 1368 24227
rect 1408 24195 1440 24227
rect 1480 24195 1512 24227
rect 1552 24195 1584 24227
rect 1624 24195 1656 24227
rect 1696 24195 1728 24227
rect 1768 24195 1800 24227
rect 1840 24195 1872 24227
rect 1912 24195 1944 24227
rect 1984 24195 2016 24227
rect 2056 24195 2088 24227
rect 2128 24195 2160 24227
rect 2200 24195 2232 24227
rect 2272 24195 2304 24227
rect 2344 24195 2376 24227
rect 2416 24195 2448 24227
rect 2488 24195 2520 24227
rect 2560 24195 2592 24227
rect 2632 24195 2664 24227
rect 2704 24195 2736 24227
rect 2776 24195 2808 24227
rect 2848 24195 2880 24227
rect 2920 24195 2952 24227
rect 2992 24195 3024 24227
rect 3064 24195 3096 24227
rect 3136 24195 3168 24227
rect 3208 24195 3240 24227
rect 3280 24195 3312 24227
rect 3352 24195 3384 24227
rect 3424 24195 3456 24227
rect 3496 24195 3528 24227
rect 3568 24195 3600 24227
rect 3640 24195 3672 24227
rect 3712 24195 3744 24227
rect 3784 24195 3816 24227
rect 3856 24195 3888 24227
rect 112 24123 144 24155
rect 184 24123 216 24155
rect 256 24123 288 24155
rect 328 24123 360 24155
rect 400 24123 432 24155
rect 472 24123 504 24155
rect 544 24123 576 24155
rect 616 24123 648 24155
rect 688 24123 720 24155
rect 760 24123 792 24155
rect 832 24123 864 24155
rect 904 24123 936 24155
rect 976 24123 1008 24155
rect 1048 24123 1080 24155
rect 1120 24123 1152 24155
rect 1192 24123 1224 24155
rect 1264 24123 1296 24155
rect 1336 24123 1368 24155
rect 1408 24123 1440 24155
rect 1480 24123 1512 24155
rect 1552 24123 1584 24155
rect 1624 24123 1656 24155
rect 1696 24123 1728 24155
rect 1768 24123 1800 24155
rect 1840 24123 1872 24155
rect 1912 24123 1944 24155
rect 1984 24123 2016 24155
rect 2056 24123 2088 24155
rect 2128 24123 2160 24155
rect 2200 24123 2232 24155
rect 2272 24123 2304 24155
rect 2344 24123 2376 24155
rect 2416 24123 2448 24155
rect 2488 24123 2520 24155
rect 2560 24123 2592 24155
rect 2632 24123 2664 24155
rect 2704 24123 2736 24155
rect 2776 24123 2808 24155
rect 2848 24123 2880 24155
rect 2920 24123 2952 24155
rect 2992 24123 3024 24155
rect 3064 24123 3096 24155
rect 3136 24123 3168 24155
rect 3208 24123 3240 24155
rect 3280 24123 3312 24155
rect 3352 24123 3384 24155
rect 3424 24123 3456 24155
rect 3496 24123 3528 24155
rect 3568 24123 3600 24155
rect 3640 24123 3672 24155
rect 3712 24123 3744 24155
rect 3784 24123 3816 24155
rect 3856 24123 3888 24155
rect 112 24051 144 24083
rect 184 24051 216 24083
rect 256 24051 288 24083
rect 328 24051 360 24083
rect 400 24051 432 24083
rect 472 24051 504 24083
rect 544 24051 576 24083
rect 616 24051 648 24083
rect 688 24051 720 24083
rect 760 24051 792 24083
rect 832 24051 864 24083
rect 904 24051 936 24083
rect 976 24051 1008 24083
rect 1048 24051 1080 24083
rect 1120 24051 1152 24083
rect 1192 24051 1224 24083
rect 1264 24051 1296 24083
rect 1336 24051 1368 24083
rect 1408 24051 1440 24083
rect 1480 24051 1512 24083
rect 1552 24051 1584 24083
rect 1624 24051 1656 24083
rect 1696 24051 1728 24083
rect 1768 24051 1800 24083
rect 1840 24051 1872 24083
rect 1912 24051 1944 24083
rect 1984 24051 2016 24083
rect 2056 24051 2088 24083
rect 2128 24051 2160 24083
rect 2200 24051 2232 24083
rect 2272 24051 2304 24083
rect 2344 24051 2376 24083
rect 2416 24051 2448 24083
rect 2488 24051 2520 24083
rect 2560 24051 2592 24083
rect 2632 24051 2664 24083
rect 2704 24051 2736 24083
rect 2776 24051 2808 24083
rect 2848 24051 2880 24083
rect 2920 24051 2952 24083
rect 2992 24051 3024 24083
rect 3064 24051 3096 24083
rect 3136 24051 3168 24083
rect 3208 24051 3240 24083
rect 3280 24051 3312 24083
rect 3352 24051 3384 24083
rect 3424 24051 3456 24083
rect 3496 24051 3528 24083
rect 3568 24051 3600 24083
rect 3640 24051 3672 24083
rect 3712 24051 3744 24083
rect 3784 24051 3816 24083
rect 3856 24051 3888 24083
rect 112 23979 144 24011
rect 184 23979 216 24011
rect 256 23979 288 24011
rect 328 23979 360 24011
rect 400 23979 432 24011
rect 472 23979 504 24011
rect 544 23979 576 24011
rect 616 23979 648 24011
rect 688 23979 720 24011
rect 760 23979 792 24011
rect 832 23979 864 24011
rect 904 23979 936 24011
rect 976 23979 1008 24011
rect 1048 23979 1080 24011
rect 1120 23979 1152 24011
rect 1192 23979 1224 24011
rect 1264 23979 1296 24011
rect 1336 23979 1368 24011
rect 1408 23979 1440 24011
rect 1480 23979 1512 24011
rect 1552 23979 1584 24011
rect 1624 23979 1656 24011
rect 1696 23979 1728 24011
rect 1768 23979 1800 24011
rect 1840 23979 1872 24011
rect 1912 23979 1944 24011
rect 1984 23979 2016 24011
rect 2056 23979 2088 24011
rect 2128 23979 2160 24011
rect 2200 23979 2232 24011
rect 2272 23979 2304 24011
rect 2344 23979 2376 24011
rect 2416 23979 2448 24011
rect 2488 23979 2520 24011
rect 2560 23979 2592 24011
rect 2632 23979 2664 24011
rect 2704 23979 2736 24011
rect 2776 23979 2808 24011
rect 2848 23979 2880 24011
rect 2920 23979 2952 24011
rect 2992 23979 3024 24011
rect 3064 23979 3096 24011
rect 3136 23979 3168 24011
rect 3208 23979 3240 24011
rect 3280 23979 3312 24011
rect 3352 23979 3384 24011
rect 3424 23979 3456 24011
rect 3496 23979 3528 24011
rect 3568 23979 3600 24011
rect 3640 23979 3672 24011
rect 3712 23979 3744 24011
rect 3784 23979 3816 24011
rect 3856 23979 3888 24011
rect 112 23907 144 23939
rect 184 23907 216 23939
rect 256 23907 288 23939
rect 328 23907 360 23939
rect 400 23907 432 23939
rect 472 23907 504 23939
rect 544 23907 576 23939
rect 616 23907 648 23939
rect 688 23907 720 23939
rect 760 23907 792 23939
rect 832 23907 864 23939
rect 904 23907 936 23939
rect 976 23907 1008 23939
rect 1048 23907 1080 23939
rect 1120 23907 1152 23939
rect 1192 23907 1224 23939
rect 1264 23907 1296 23939
rect 1336 23907 1368 23939
rect 1408 23907 1440 23939
rect 1480 23907 1512 23939
rect 1552 23907 1584 23939
rect 1624 23907 1656 23939
rect 1696 23907 1728 23939
rect 1768 23907 1800 23939
rect 1840 23907 1872 23939
rect 1912 23907 1944 23939
rect 1984 23907 2016 23939
rect 2056 23907 2088 23939
rect 2128 23907 2160 23939
rect 2200 23907 2232 23939
rect 2272 23907 2304 23939
rect 2344 23907 2376 23939
rect 2416 23907 2448 23939
rect 2488 23907 2520 23939
rect 2560 23907 2592 23939
rect 2632 23907 2664 23939
rect 2704 23907 2736 23939
rect 2776 23907 2808 23939
rect 2848 23907 2880 23939
rect 2920 23907 2952 23939
rect 2992 23907 3024 23939
rect 3064 23907 3096 23939
rect 3136 23907 3168 23939
rect 3208 23907 3240 23939
rect 3280 23907 3312 23939
rect 3352 23907 3384 23939
rect 3424 23907 3456 23939
rect 3496 23907 3528 23939
rect 3568 23907 3600 23939
rect 3640 23907 3672 23939
rect 3712 23907 3744 23939
rect 3784 23907 3816 23939
rect 3856 23907 3888 23939
rect 112 23835 144 23867
rect 184 23835 216 23867
rect 256 23835 288 23867
rect 328 23835 360 23867
rect 400 23835 432 23867
rect 472 23835 504 23867
rect 544 23835 576 23867
rect 616 23835 648 23867
rect 688 23835 720 23867
rect 760 23835 792 23867
rect 832 23835 864 23867
rect 904 23835 936 23867
rect 976 23835 1008 23867
rect 1048 23835 1080 23867
rect 1120 23835 1152 23867
rect 1192 23835 1224 23867
rect 1264 23835 1296 23867
rect 1336 23835 1368 23867
rect 1408 23835 1440 23867
rect 1480 23835 1512 23867
rect 1552 23835 1584 23867
rect 1624 23835 1656 23867
rect 1696 23835 1728 23867
rect 1768 23835 1800 23867
rect 1840 23835 1872 23867
rect 1912 23835 1944 23867
rect 1984 23835 2016 23867
rect 2056 23835 2088 23867
rect 2128 23835 2160 23867
rect 2200 23835 2232 23867
rect 2272 23835 2304 23867
rect 2344 23835 2376 23867
rect 2416 23835 2448 23867
rect 2488 23835 2520 23867
rect 2560 23835 2592 23867
rect 2632 23835 2664 23867
rect 2704 23835 2736 23867
rect 2776 23835 2808 23867
rect 2848 23835 2880 23867
rect 2920 23835 2952 23867
rect 2992 23835 3024 23867
rect 3064 23835 3096 23867
rect 3136 23835 3168 23867
rect 3208 23835 3240 23867
rect 3280 23835 3312 23867
rect 3352 23835 3384 23867
rect 3424 23835 3456 23867
rect 3496 23835 3528 23867
rect 3568 23835 3600 23867
rect 3640 23835 3672 23867
rect 3712 23835 3744 23867
rect 3784 23835 3816 23867
rect 3856 23835 3888 23867
rect 112 23763 144 23795
rect 184 23763 216 23795
rect 256 23763 288 23795
rect 328 23763 360 23795
rect 400 23763 432 23795
rect 472 23763 504 23795
rect 544 23763 576 23795
rect 616 23763 648 23795
rect 688 23763 720 23795
rect 760 23763 792 23795
rect 832 23763 864 23795
rect 904 23763 936 23795
rect 976 23763 1008 23795
rect 1048 23763 1080 23795
rect 1120 23763 1152 23795
rect 1192 23763 1224 23795
rect 1264 23763 1296 23795
rect 1336 23763 1368 23795
rect 1408 23763 1440 23795
rect 1480 23763 1512 23795
rect 1552 23763 1584 23795
rect 1624 23763 1656 23795
rect 1696 23763 1728 23795
rect 1768 23763 1800 23795
rect 1840 23763 1872 23795
rect 1912 23763 1944 23795
rect 1984 23763 2016 23795
rect 2056 23763 2088 23795
rect 2128 23763 2160 23795
rect 2200 23763 2232 23795
rect 2272 23763 2304 23795
rect 2344 23763 2376 23795
rect 2416 23763 2448 23795
rect 2488 23763 2520 23795
rect 2560 23763 2592 23795
rect 2632 23763 2664 23795
rect 2704 23763 2736 23795
rect 2776 23763 2808 23795
rect 2848 23763 2880 23795
rect 2920 23763 2952 23795
rect 2992 23763 3024 23795
rect 3064 23763 3096 23795
rect 3136 23763 3168 23795
rect 3208 23763 3240 23795
rect 3280 23763 3312 23795
rect 3352 23763 3384 23795
rect 3424 23763 3456 23795
rect 3496 23763 3528 23795
rect 3568 23763 3600 23795
rect 3640 23763 3672 23795
rect 3712 23763 3744 23795
rect 3784 23763 3816 23795
rect 3856 23763 3888 23795
rect 112 23691 144 23723
rect 184 23691 216 23723
rect 256 23691 288 23723
rect 328 23691 360 23723
rect 400 23691 432 23723
rect 472 23691 504 23723
rect 544 23691 576 23723
rect 616 23691 648 23723
rect 688 23691 720 23723
rect 760 23691 792 23723
rect 832 23691 864 23723
rect 904 23691 936 23723
rect 976 23691 1008 23723
rect 1048 23691 1080 23723
rect 1120 23691 1152 23723
rect 1192 23691 1224 23723
rect 1264 23691 1296 23723
rect 1336 23691 1368 23723
rect 1408 23691 1440 23723
rect 1480 23691 1512 23723
rect 1552 23691 1584 23723
rect 1624 23691 1656 23723
rect 1696 23691 1728 23723
rect 1768 23691 1800 23723
rect 1840 23691 1872 23723
rect 1912 23691 1944 23723
rect 1984 23691 2016 23723
rect 2056 23691 2088 23723
rect 2128 23691 2160 23723
rect 2200 23691 2232 23723
rect 2272 23691 2304 23723
rect 2344 23691 2376 23723
rect 2416 23691 2448 23723
rect 2488 23691 2520 23723
rect 2560 23691 2592 23723
rect 2632 23691 2664 23723
rect 2704 23691 2736 23723
rect 2776 23691 2808 23723
rect 2848 23691 2880 23723
rect 2920 23691 2952 23723
rect 2992 23691 3024 23723
rect 3064 23691 3096 23723
rect 3136 23691 3168 23723
rect 3208 23691 3240 23723
rect 3280 23691 3312 23723
rect 3352 23691 3384 23723
rect 3424 23691 3456 23723
rect 3496 23691 3528 23723
rect 3568 23691 3600 23723
rect 3640 23691 3672 23723
rect 3712 23691 3744 23723
rect 3784 23691 3816 23723
rect 3856 23691 3888 23723
rect 112 23619 144 23651
rect 184 23619 216 23651
rect 256 23619 288 23651
rect 328 23619 360 23651
rect 400 23619 432 23651
rect 472 23619 504 23651
rect 544 23619 576 23651
rect 616 23619 648 23651
rect 688 23619 720 23651
rect 760 23619 792 23651
rect 832 23619 864 23651
rect 904 23619 936 23651
rect 976 23619 1008 23651
rect 1048 23619 1080 23651
rect 1120 23619 1152 23651
rect 1192 23619 1224 23651
rect 1264 23619 1296 23651
rect 1336 23619 1368 23651
rect 1408 23619 1440 23651
rect 1480 23619 1512 23651
rect 1552 23619 1584 23651
rect 1624 23619 1656 23651
rect 1696 23619 1728 23651
rect 1768 23619 1800 23651
rect 1840 23619 1872 23651
rect 1912 23619 1944 23651
rect 1984 23619 2016 23651
rect 2056 23619 2088 23651
rect 2128 23619 2160 23651
rect 2200 23619 2232 23651
rect 2272 23619 2304 23651
rect 2344 23619 2376 23651
rect 2416 23619 2448 23651
rect 2488 23619 2520 23651
rect 2560 23619 2592 23651
rect 2632 23619 2664 23651
rect 2704 23619 2736 23651
rect 2776 23619 2808 23651
rect 2848 23619 2880 23651
rect 2920 23619 2952 23651
rect 2992 23619 3024 23651
rect 3064 23619 3096 23651
rect 3136 23619 3168 23651
rect 3208 23619 3240 23651
rect 3280 23619 3312 23651
rect 3352 23619 3384 23651
rect 3424 23619 3456 23651
rect 3496 23619 3528 23651
rect 3568 23619 3600 23651
rect 3640 23619 3672 23651
rect 3712 23619 3744 23651
rect 3784 23619 3816 23651
rect 3856 23619 3888 23651
rect 112 23547 144 23579
rect 184 23547 216 23579
rect 256 23547 288 23579
rect 328 23547 360 23579
rect 400 23547 432 23579
rect 472 23547 504 23579
rect 544 23547 576 23579
rect 616 23547 648 23579
rect 688 23547 720 23579
rect 760 23547 792 23579
rect 832 23547 864 23579
rect 904 23547 936 23579
rect 976 23547 1008 23579
rect 1048 23547 1080 23579
rect 1120 23547 1152 23579
rect 1192 23547 1224 23579
rect 1264 23547 1296 23579
rect 1336 23547 1368 23579
rect 1408 23547 1440 23579
rect 1480 23547 1512 23579
rect 1552 23547 1584 23579
rect 1624 23547 1656 23579
rect 1696 23547 1728 23579
rect 1768 23547 1800 23579
rect 1840 23547 1872 23579
rect 1912 23547 1944 23579
rect 1984 23547 2016 23579
rect 2056 23547 2088 23579
rect 2128 23547 2160 23579
rect 2200 23547 2232 23579
rect 2272 23547 2304 23579
rect 2344 23547 2376 23579
rect 2416 23547 2448 23579
rect 2488 23547 2520 23579
rect 2560 23547 2592 23579
rect 2632 23547 2664 23579
rect 2704 23547 2736 23579
rect 2776 23547 2808 23579
rect 2848 23547 2880 23579
rect 2920 23547 2952 23579
rect 2992 23547 3024 23579
rect 3064 23547 3096 23579
rect 3136 23547 3168 23579
rect 3208 23547 3240 23579
rect 3280 23547 3312 23579
rect 3352 23547 3384 23579
rect 3424 23547 3456 23579
rect 3496 23547 3528 23579
rect 3568 23547 3600 23579
rect 3640 23547 3672 23579
rect 3712 23547 3744 23579
rect 3784 23547 3816 23579
rect 3856 23547 3888 23579
rect 112 23475 144 23507
rect 184 23475 216 23507
rect 256 23475 288 23507
rect 328 23475 360 23507
rect 400 23475 432 23507
rect 472 23475 504 23507
rect 544 23475 576 23507
rect 616 23475 648 23507
rect 688 23475 720 23507
rect 760 23475 792 23507
rect 832 23475 864 23507
rect 904 23475 936 23507
rect 976 23475 1008 23507
rect 1048 23475 1080 23507
rect 1120 23475 1152 23507
rect 1192 23475 1224 23507
rect 1264 23475 1296 23507
rect 1336 23475 1368 23507
rect 1408 23475 1440 23507
rect 1480 23475 1512 23507
rect 1552 23475 1584 23507
rect 1624 23475 1656 23507
rect 1696 23475 1728 23507
rect 1768 23475 1800 23507
rect 1840 23475 1872 23507
rect 1912 23475 1944 23507
rect 1984 23475 2016 23507
rect 2056 23475 2088 23507
rect 2128 23475 2160 23507
rect 2200 23475 2232 23507
rect 2272 23475 2304 23507
rect 2344 23475 2376 23507
rect 2416 23475 2448 23507
rect 2488 23475 2520 23507
rect 2560 23475 2592 23507
rect 2632 23475 2664 23507
rect 2704 23475 2736 23507
rect 2776 23475 2808 23507
rect 2848 23475 2880 23507
rect 2920 23475 2952 23507
rect 2992 23475 3024 23507
rect 3064 23475 3096 23507
rect 3136 23475 3168 23507
rect 3208 23475 3240 23507
rect 3280 23475 3312 23507
rect 3352 23475 3384 23507
rect 3424 23475 3456 23507
rect 3496 23475 3528 23507
rect 3568 23475 3600 23507
rect 3640 23475 3672 23507
rect 3712 23475 3744 23507
rect 3784 23475 3816 23507
rect 3856 23475 3888 23507
rect 112 23403 144 23435
rect 184 23403 216 23435
rect 256 23403 288 23435
rect 328 23403 360 23435
rect 400 23403 432 23435
rect 472 23403 504 23435
rect 544 23403 576 23435
rect 616 23403 648 23435
rect 688 23403 720 23435
rect 760 23403 792 23435
rect 832 23403 864 23435
rect 904 23403 936 23435
rect 976 23403 1008 23435
rect 1048 23403 1080 23435
rect 1120 23403 1152 23435
rect 1192 23403 1224 23435
rect 1264 23403 1296 23435
rect 1336 23403 1368 23435
rect 1408 23403 1440 23435
rect 1480 23403 1512 23435
rect 1552 23403 1584 23435
rect 1624 23403 1656 23435
rect 1696 23403 1728 23435
rect 1768 23403 1800 23435
rect 1840 23403 1872 23435
rect 1912 23403 1944 23435
rect 1984 23403 2016 23435
rect 2056 23403 2088 23435
rect 2128 23403 2160 23435
rect 2200 23403 2232 23435
rect 2272 23403 2304 23435
rect 2344 23403 2376 23435
rect 2416 23403 2448 23435
rect 2488 23403 2520 23435
rect 2560 23403 2592 23435
rect 2632 23403 2664 23435
rect 2704 23403 2736 23435
rect 2776 23403 2808 23435
rect 2848 23403 2880 23435
rect 2920 23403 2952 23435
rect 2992 23403 3024 23435
rect 3064 23403 3096 23435
rect 3136 23403 3168 23435
rect 3208 23403 3240 23435
rect 3280 23403 3312 23435
rect 3352 23403 3384 23435
rect 3424 23403 3456 23435
rect 3496 23403 3528 23435
rect 3568 23403 3600 23435
rect 3640 23403 3672 23435
rect 3712 23403 3744 23435
rect 3784 23403 3816 23435
rect 3856 23403 3888 23435
rect 112 23331 144 23363
rect 184 23331 216 23363
rect 256 23331 288 23363
rect 328 23331 360 23363
rect 400 23331 432 23363
rect 472 23331 504 23363
rect 544 23331 576 23363
rect 616 23331 648 23363
rect 688 23331 720 23363
rect 760 23331 792 23363
rect 832 23331 864 23363
rect 904 23331 936 23363
rect 976 23331 1008 23363
rect 1048 23331 1080 23363
rect 1120 23331 1152 23363
rect 1192 23331 1224 23363
rect 1264 23331 1296 23363
rect 1336 23331 1368 23363
rect 1408 23331 1440 23363
rect 1480 23331 1512 23363
rect 1552 23331 1584 23363
rect 1624 23331 1656 23363
rect 1696 23331 1728 23363
rect 1768 23331 1800 23363
rect 1840 23331 1872 23363
rect 1912 23331 1944 23363
rect 1984 23331 2016 23363
rect 2056 23331 2088 23363
rect 2128 23331 2160 23363
rect 2200 23331 2232 23363
rect 2272 23331 2304 23363
rect 2344 23331 2376 23363
rect 2416 23331 2448 23363
rect 2488 23331 2520 23363
rect 2560 23331 2592 23363
rect 2632 23331 2664 23363
rect 2704 23331 2736 23363
rect 2776 23331 2808 23363
rect 2848 23331 2880 23363
rect 2920 23331 2952 23363
rect 2992 23331 3024 23363
rect 3064 23331 3096 23363
rect 3136 23331 3168 23363
rect 3208 23331 3240 23363
rect 3280 23331 3312 23363
rect 3352 23331 3384 23363
rect 3424 23331 3456 23363
rect 3496 23331 3528 23363
rect 3568 23331 3600 23363
rect 3640 23331 3672 23363
rect 3712 23331 3744 23363
rect 3784 23331 3816 23363
rect 3856 23331 3888 23363
rect 112 23259 144 23291
rect 184 23259 216 23291
rect 256 23259 288 23291
rect 328 23259 360 23291
rect 400 23259 432 23291
rect 472 23259 504 23291
rect 544 23259 576 23291
rect 616 23259 648 23291
rect 688 23259 720 23291
rect 760 23259 792 23291
rect 832 23259 864 23291
rect 904 23259 936 23291
rect 976 23259 1008 23291
rect 1048 23259 1080 23291
rect 1120 23259 1152 23291
rect 1192 23259 1224 23291
rect 1264 23259 1296 23291
rect 1336 23259 1368 23291
rect 1408 23259 1440 23291
rect 1480 23259 1512 23291
rect 1552 23259 1584 23291
rect 1624 23259 1656 23291
rect 1696 23259 1728 23291
rect 1768 23259 1800 23291
rect 1840 23259 1872 23291
rect 1912 23259 1944 23291
rect 1984 23259 2016 23291
rect 2056 23259 2088 23291
rect 2128 23259 2160 23291
rect 2200 23259 2232 23291
rect 2272 23259 2304 23291
rect 2344 23259 2376 23291
rect 2416 23259 2448 23291
rect 2488 23259 2520 23291
rect 2560 23259 2592 23291
rect 2632 23259 2664 23291
rect 2704 23259 2736 23291
rect 2776 23259 2808 23291
rect 2848 23259 2880 23291
rect 2920 23259 2952 23291
rect 2992 23259 3024 23291
rect 3064 23259 3096 23291
rect 3136 23259 3168 23291
rect 3208 23259 3240 23291
rect 3280 23259 3312 23291
rect 3352 23259 3384 23291
rect 3424 23259 3456 23291
rect 3496 23259 3528 23291
rect 3568 23259 3600 23291
rect 3640 23259 3672 23291
rect 3712 23259 3744 23291
rect 3784 23259 3816 23291
rect 3856 23259 3888 23291
rect 112 23187 144 23219
rect 184 23187 216 23219
rect 256 23187 288 23219
rect 328 23187 360 23219
rect 400 23187 432 23219
rect 472 23187 504 23219
rect 544 23187 576 23219
rect 616 23187 648 23219
rect 688 23187 720 23219
rect 760 23187 792 23219
rect 832 23187 864 23219
rect 904 23187 936 23219
rect 976 23187 1008 23219
rect 1048 23187 1080 23219
rect 1120 23187 1152 23219
rect 1192 23187 1224 23219
rect 1264 23187 1296 23219
rect 1336 23187 1368 23219
rect 1408 23187 1440 23219
rect 1480 23187 1512 23219
rect 1552 23187 1584 23219
rect 1624 23187 1656 23219
rect 1696 23187 1728 23219
rect 1768 23187 1800 23219
rect 1840 23187 1872 23219
rect 1912 23187 1944 23219
rect 1984 23187 2016 23219
rect 2056 23187 2088 23219
rect 2128 23187 2160 23219
rect 2200 23187 2232 23219
rect 2272 23187 2304 23219
rect 2344 23187 2376 23219
rect 2416 23187 2448 23219
rect 2488 23187 2520 23219
rect 2560 23187 2592 23219
rect 2632 23187 2664 23219
rect 2704 23187 2736 23219
rect 2776 23187 2808 23219
rect 2848 23187 2880 23219
rect 2920 23187 2952 23219
rect 2992 23187 3024 23219
rect 3064 23187 3096 23219
rect 3136 23187 3168 23219
rect 3208 23187 3240 23219
rect 3280 23187 3312 23219
rect 3352 23187 3384 23219
rect 3424 23187 3456 23219
rect 3496 23187 3528 23219
rect 3568 23187 3600 23219
rect 3640 23187 3672 23219
rect 3712 23187 3744 23219
rect 3784 23187 3816 23219
rect 3856 23187 3888 23219
rect 184 22842 216 22874
rect 256 22842 288 22874
rect 328 22842 360 22874
rect 400 22842 432 22874
rect 472 22842 504 22874
rect 544 22842 576 22874
rect 616 22842 648 22874
rect 688 22842 720 22874
rect 760 22842 792 22874
rect 832 22842 864 22874
rect 904 22842 936 22874
rect 976 22842 1008 22874
rect 1048 22842 1080 22874
rect 1120 22842 1152 22874
rect 1192 22842 1224 22874
rect 1264 22842 1296 22874
rect 1336 22842 1368 22874
rect 1408 22842 1440 22874
rect 1480 22842 1512 22874
rect 1552 22842 1584 22874
rect 1624 22842 1656 22874
rect 1696 22842 1728 22874
rect 1768 22842 1800 22874
rect 1840 22842 1872 22874
rect 1912 22842 1944 22874
rect 1984 22842 2016 22874
rect 2056 22842 2088 22874
rect 2128 22842 2160 22874
rect 2200 22842 2232 22874
rect 2272 22842 2304 22874
rect 2344 22842 2376 22874
rect 2416 22842 2448 22874
rect 2488 22842 2520 22874
rect 2560 22842 2592 22874
rect 2632 22842 2664 22874
rect 2704 22842 2736 22874
rect 2776 22842 2808 22874
rect 2848 22842 2880 22874
rect 2920 22842 2952 22874
rect 2992 22842 3024 22874
rect 3064 22842 3096 22874
rect 3136 22842 3168 22874
rect 3208 22842 3240 22874
rect 3280 22842 3312 22874
rect 3352 22842 3384 22874
rect 3424 22842 3456 22874
rect 3496 22842 3528 22874
rect 3568 22842 3600 22874
rect 3640 22842 3672 22874
rect 3712 22842 3744 22874
rect 3784 22842 3816 22874
rect 3856 22842 3888 22874
rect 112 22770 144 22802
rect 184 22770 216 22802
rect 256 22770 288 22802
rect 328 22770 360 22802
rect 400 22770 432 22802
rect 472 22770 504 22802
rect 544 22770 576 22802
rect 616 22770 648 22802
rect 688 22770 720 22802
rect 760 22770 792 22802
rect 832 22770 864 22802
rect 904 22770 936 22802
rect 976 22770 1008 22802
rect 1048 22770 1080 22802
rect 1120 22770 1152 22802
rect 1192 22770 1224 22802
rect 1264 22770 1296 22802
rect 1336 22770 1368 22802
rect 1408 22770 1440 22802
rect 1480 22770 1512 22802
rect 1552 22770 1584 22802
rect 1624 22770 1656 22802
rect 1696 22770 1728 22802
rect 1768 22770 1800 22802
rect 1840 22770 1872 22802
rect 1912 22770 1944 22802
rect 1984 22770 2016 22802
rect 2056 22770 2088 22802
rect 2128 22770 2160 22802
rect 2200 22770 2232 22802
rect 2272 22770 2304 22802
rect 2344 22770 2376 22802
rect 2416 22770 2448 22802
rect 2488 22770 2520 22802
rect 2560 22770 2592 22802
rect 2632 22770 2664 22802
rect 2704 22770 2736 22802
rect 2776 22770 2808 22802
rect 2848 22770 2880 22802
rect 2920 22770 2952 22802
rect 2992 22770 3024 22802
rect 3064 22770 3096 22802
rect 3136 22770 3168 22802
rect 3208 22770 3240 22802
rect 3280 22770 3312 22802
rect 3352 22770 3384 22802
rect 3424 22770 3456 22802
rect 3496 22770 3528 22802
rect 3568 22770 3600 22802
rect 3640 22770 3672 22802
rect 3712 22770 3744 22802
rect 3784 22770 3816 22802
rect 3856 22770 3888 22802
rect 112 22698 144 22730
rect 184 22698 216 22730
rect 256 22698 288 22730
rect 328 22698 360 22730
rect 400 22698 432 22730
rect 472 22698 504 22730
rect 544 22698 576 22730
rect 616 22698 648 22730
rect 688 22698 720 22730
rect 760 22698 792 22730
rect 832 22698 864 22730
rect 904 22698 936 22730
rect 976 22698 1008 22730
rect 1048 22698 1080 22730
rect 1120 22698 1152 22730
rect 1192 22698 1224 22730
rect 1264 22698 1296 22730
rect 1336 22698 1368 22730
rect 1408 22698 1440 22730
rect 1480 22698 1512 22730
rect 1552 22698 1584 22730
rect 1624 22698 1656 22730
rect 1696 22698 1728 22730
rect 1768 22698 1800 22730
rect 1840 22698 1872 22730
rect 1912 22698 1944 22730
rect 1984 22698 2016 22730
rect 2056 22698 2088 22730
rect 2128 22698 2160 22730
rect 2200 22698 2232 22730
rect 2272 22698 2304 22730
rect 2344 22698 2376 22730
rect 2416 22698 2448 22730
rect 2488 22698 2520 22730
rect 2560 22698 2592 22730
rect 2632 22698 2664 22730
rect 2704 22698 2736 22730
rect 2776 22698 2808 22730
rect 2848 22698 2880 22730
rect 2920 22698 2952 22730
rect 2992 22698 3024 22730
rect 3064 22698 3096 22730
rect 3136 22698 3168 22730
rect 3208 22698 3240 22730
rect 3280 22698 3312 22730
rect 3352 22698 3384 22730
rect 3424 22698 3456 22730
rect 3496 22698 3528 22730
rect 3568 22698 3600 22730
rect 3640 22698 3672 22730
rect 3712 22698 3744 22730
rect 3784 22698 3816 22730
rect 3856 22698 3888 22730
rect 112 22626 144 22658
rect 184 22626 216 22658
rect 256 22626 288 22658
rect 328 22626 360 22658
rect 400 22626 432 22658
rect 472 22626 504 22658
rect 544 22626 576 22658
rect 616 22626 648 22658
rect 688 22626 720 22658
rect 760 22626 792 22658
rect 832 22626 864 22658
rect 904 22626 936 22658
rect 976 22626 1008 22658
rect 1048 22626 1080 22658
rect 1120 22626 1152 22658
rect 1192 22626 1224 22658
rect 1264 22626 1296 22658
rect 1336 22626 1368 22658
rect 1408 22626 1440 22658
rect 1480 22626 1512 22658
rect 1552 22626 1584 22658
rect 1624 22626 1656 22658
rect 1696 22626 1728 22658
rect 1768 22626 1800 22658
rect 1840 22626 1872 22658
rect 1912 22626 1944 22658
rect 1984 22626 2016 22658
rect 2056 22626 2088 22658
rect 2128 22626 2160 22658
rect 2200 22626 2232 22658
rect 2272 22626 2304 22658
rect 2344 22626 2376 22658
rect 2416 22626 2448 22658
rect 2488 22626 2520 22658
rect 2560 22626 2592 22658
rect 2632 22626 2664 22658
rect 2704 22626 2736 22658
rect 2776 22626 2808 22658
rect 2848 22626 2880 22658
rect 2920 22626 2952 22658
rect 2992 22626 3024 22658
rect 3064 22626 3096 22658
rect 3136 22626 3168 22658
rect 3208 22626 3240 22658
rect 3280 22626 3312 22658
rect 3352 22626 3384 22658
rect 3424 22626 3456 22658
rect 3496 22626 3528 22658
rect 3568 22626 3600 22658
rect 3640 22626 3672 22658
rect 3712 22626 3744 22658
rect 3784 22626 3816 22658
rect 3856 22626 3888 22658
rect 112 22554 144 22586
rect 184 22554 216 22586
rect 256 22554 288 22586
rect 328 22554 360 22586
rect 400 22554 432 22586
rect 472 22554 504 22586
rect 544 22554 576 22586
rect 616 22554 648 22586
rect 688 22554 720 22586
rect 760 22554 792 22586
rect 832 22554 864 22586
rect 904 22554 936 22586
rect 976 22554 1008 22586
rect 1048 22554 1080 22586
rect 1120 22554 1152 22586
rect 1192 22554 1224 22586
rect 1264 22554 1296 22586
rect 1336 22554 1368 22586
rect 1408 22554 1440 22586
rect 1480 22554 1512 22586
rect 1552 22554 1584 22586
rect 1624 22554 1656 22586
rect 1696 22554 1728 22586
rect 1768 22554 1800 22586
rect 1840 22554 1872 22586
rect 1912 22554 1944 22586
rect 1984 22554 2016 22586
rect 2056 22554 2088 22586
rect 2128 22554 2160 22586
rect 2200 22554 2232 22586
rect 2272 22554 2304 22586
rect 2344 22554 2376 22586
rect 2416 22554 2448 22586
rect 2488 22554 2520 22586
rect 2560 22554 2592 22586
rect 2632 22554 2664 22586
rect 2704 22554 2736 22586
rect 2776 22554 2808 22586
rect 2848 22554 2880 22586
rect 2920 22554 2952 22586
rect 2992 22554 3024 22586
rect 3064 22554 3096 22586
rect 3136 22554 3168 22586
rect 3208 22554 3240 22586
rect 3280 22554 3312 22586
rect 3352 22554 3384 22586
rect 3424 22554 3456 22586
rect 3496 22554 3528 22586
rect 3568 22554 3600 22586
rect 3640 22554 3672 22586
rect 3712 22554 3744 22586
rect 3784 22554 3816 22586
rect 3856 22554 3888 22586
rect 112 22482 144 22514
rect 184 22482 216 22514
rect 256 22482 288 22514
rect 328 22482 360 22514
rect 400 22482 432 22514
rect 472 22482 504 22514
rect 544 22482 576 22514
rect 616 22482 648 22514
rect 688 22482 720 22514
rect 760 22482 792 22514
rect 832 22482 864 22514
rect 904 22482 936 22514
rect 976 22482 1008 22514
rect 1048 22482 1080 22514
rect 1120 22482 1152 22514
rect 1192 22482 1224 22514
rect 1264 22482 1296 22514
rect 1336 22482 1368 22514
rect 1408 22482 1440 22514
rect 1480 22482 1512 22514
rect 1552 22482 1584 22514
rect 1624 22482 1656 22514
rect 1696 22482 1728 22514
rect 1768 22482 1800 22514
rect 1840 22482 1872 22514
rect 1912 22482 1944 22514
rect 1984 22482 2016 22514
rect 2056 22482 2088 22514
rect 2128 22482 2160 22514
rect 2200 22482 2232 22514
rect 2272 22482 2304 22514
rect 2344 22482 2376 22514
rect 2416 22482 2448 22514
rect 2488 22482 2520 22514
rect 2560 22482 2592 22514
rect 2632 22482 2664 22514
rect 2704 22482 2736 22514
rect 2776 22482 2808 22514
rect 2848 22482 2880 22514
rect 2920 22482 2952 22514
rect 2992 22482 3024 22514
rect 3064 22482 3096 22514
rect 3136 22482 3168 22514
rect 3208 22482 3240 22514
rect 3280 22482 3312 22514
rect 3352 22482 3384 22514
rect 3424 22482 3456 22514
rect 3496 22482 3528 22514
rect 3568 22482 3600 22514
rect 3640 22482 3672 22514
rect 3712 22482 3744 22514
rect 3784 22482 3816 22514
rect 3856 22482 3888 22514
rect 112 22410 144 22442
rect 184 22410 216 22442
rect 256 22410 288 22442
rect 328 22410 360 22442
rect 400 22410 432 22442
rect 472 22410 504 22442
rect 544 22410 576 22442
rect 616 22410 648 22442
rect 688 22410 720 22442
rect 760 22410 792 22442
rect 832 22410 864 22442
rect 904 22410 936 22442
rect 976 22410 1008 22442
rect 1048 22410 1080 22442
rect 1120 22410 1152 22442
rect 1192 22410 1224 22442
rect 1264 22410 1296 22442
rect 1336 22410 1368 22442
rect 1408 22410 1440 22442
rect 1480 22410 1512 22442
rect 1552 22410 1584 22442
rect 1624 22410 1656 22442
rect 1696 22410 1728 22442
rect 1768 22410 1800 22442
rect 1840 22410 1872 22442
rect 1912 22410 1944 22442
rect 1984 22410 2016 22442
rect 2056 22410 2088 22442
rect 2128 22410 2160 22442
rect 2200 22410 2232 22442
rect 2272 22410 2304 22442
rect 2344 22410 2376 22442
rect 2416 22410 2448 22442
rect 2488 22410 2520 22442
rect 2560 22410 2592 22442
rect 2632 22410 2664 22442
rect 2704 22410 2736 22442
rect 2776 22410 2808 22442
rect 2848 22410 2880 22442
rect 2920 22410 2952 22442
rect 2992 22410 3024 22442
rect 3064 22410 3096 22442
rect 3136 22410 3168 22442
rect 3208 22410 3240 22442
rect 3280 22410 3312 22442
rect 3352 22410 3384 22442
rect 3424 22410 3456 22442
rect 3496 22410 3528 22442
rect 3568 22410 3600 22442
rect 3640 22410 3672 22442
rect 3712 22410 3744 22442
rect 3784 22410 3816 22442
rect 3856 22410 3888 22442
rect 112 22338 144 22370
rect 184 22338 216 22370
rect 256 22338 288 22370
rect 328 22338 360 22370
rect 400 22338 432 22370
rect 472 22338 504 22370
rect 544 22338 576 22370
rect 616 22338 648 22370
rect 688 22338 720 22370
rect 760 22338 792 22370
rect 832 22338 864 22370
rect 904 22338 936 22370
rect 976 22338 1008 22370
rect 1048 22338 1080 22370
rect 1120 22338 1152 22370
rect 1192 22338 1224 22370
rect 1264 22338 1296 22370
rect 1336 22338 1368 22370
rect 1408 22338 1440 22370
rect 1480 22338 1512 22370
rect 1552 22338 1584 22370
rect 1624 22338 1656 22370
rect 1696 22338 1728 22370
rect 1768 22338 1800 22370
rect 1840 22338 1872 22370
rect 1912 22338 1944 22370
rect 1984 22338 2016 22370
rect 2056 22338 2088 22370
rect 2128 22338 2160 22370
rect 2200 22338 2232 22370
rect 2272 22338 2304 22370
rect 2344 22338 2376 22370
rect 2416 22338 2448 22370
rect 2488 22338 2520 22370
rect 2560 22338 2592 22370
rect 2632 22338 2664 22370
rect 2704 22338 2736 22370
rect 2776 22338 2808 22370
rect 2848 22338 2880 22370
rect 2920 22338 2952 22370
rect 2992 22338 3024 22370
rect 3064 22338 3096 22370
rect 3136 22338 3168 22370
rect 3208 22338 3240 22370
rect 3280 22338 3312 22370
rect 3352 22338 3384 22370
rect 3424 22338 3456 22370
rect 3496 22338 3528 22370
rect 3568 22338 3600 22370
rect 3640 22338 3672 22370
rect 3712 22338 3744 22370
rect 3784 22338 3816 22370
rect 3856 22338 3888 22370
rect 112 22266 144 22298
rect 184 22266 216 22298
rect 256 22266 288 22298
rect 328 22266 360 22298
rect 400 22266 432 22298
rect 472 22266 504 22298
rect 544 22266 576 22298
rect 616 22266 648 22298
rect 688 22266 720 22298
rect 760 22266 792 22298
rect 832 22266 864 22298
rect 904 22266 936 22298
rect 976 22266 1008 22298
rect 1048 22266 1080 22298
rect 1120 22266 1152 22298
rect 1192 22266 1224 22298
rect 1264 22266 1296 22298
rect 1336 22266 1368 22298
rect 1408 22266 1440 22298
rect 1480 22266 1512 22298
rect 1552 22266 1584 22298
rect 1624 22266 1656 22298
rect 1696 22266 1728 22298
rect 1768 22266 1800 22298
rect 1840 22266 1872 22298
rect 1912 22266 1944 22298
rect 1984 22266 2016 22298
rect 2056 22266 2088 22298
rect 2128 22266 2160 22298
rect 2200 22266 2232 22298
rect 2272 22266 2304 22298
rect 2344 22266 2376 22298
rect 2416 22266 2448 22298
rect 2488 22266 2520 22298
rect 2560 22266 2592 22298
rect 2632 22266 2664 22298
rect 2704 22266 2736 22298
rect 2776 22266 2808 22298
rect 2848 22266 2880 22298
rect 2920 22266 2952 22298
rect 2992 22266 3024 22298
rect 3064 22266 3096 22298
rect 3136 22266 3168 22298
rect 3208 22266 3240 22298
rect 3280 22266 3312 22298
rect 3352 22266 3384 22298
rect 3424 22266 3456 22298
rect 3496 22266 3528 22298
rect 3568 22266 3600 22298
rect 3640 22266 3672 22298
rect 3712 22266 3744 22298
rect 3784 22266 3816 22298
rect 3856 22266 3888 22298
rect 112 22194 144 22226
rect 184 22194 216 22226
rect 256 22194 288 22226
rect 328 22194 360 22226
rect 400 22194 432 22226
rect 472 22194 504 22226
rect 544 22194 576 22226
rect 616 22194 648 22226
rect 688 22194 720 22226
rect 760 22194 792 22226
rect 832 22194 864 22226
rect 904 22194 936 22226
rect 976 22194 1008 22226
rect 1048 22194 1080 22226
rect 1120 22194 1152 22226
rect 1192 22194 1224 22226
rect 1264 22194 1296 22226
rect 1336 22194 1368 22226
rect 1408 22194 1440 22226
rect 1480 22194 1512 22226
rect 1552 22194 1584 22226
rect 1624 22194 1656 22226
rect 1696 22194 1728 22226
rect 1768 22194 1800 22226
rect 1840 22194 1872 22226
rect 1912 22194 1944 22226
rect 1984 22194 2016 22226
rect 2056 22194 2088 22226
rect 2128 22194 2160 22226
rect 2200 22194 2232 22226
rect 2272 22194 2304 22226
rect 2344 22194 2376 22226
rect 2416 22194 2448 22226
rect 2488 22194 2520 22226
rect 2560 22194 2592 22226
rect 2632 22194 2664 22226
rect 2704 22194 2736 22226
rect 2776 22194 2808 22226
rect 2848 22194 2880 22226
rect 2920 22194 2952 22226
rect 2992 22194 3024 22226
rect 3064 22194 3096 22226
rect 3136 22194 3168 22226
rect 3208 22194 3240 22226
rect 3280 22194 3312 22226
rect 3352 22194 3384 22226
rect 3424 22194 3456 22226
rect 3496 22194 3528 22226
rect 3568 22194 3600 22226
rect 3640 22194 3672 22226
rect 3712 22194 3744 22226
rect 3784 22194 3816 22226
rect 3856 22194 3888 22226
rect 112 22122 144 22154
rect 184 22122 216 22154
rect 256 22122 288 22154
rect 328 22122 360 22154
rect 400 22122 432 22154
rect 472 22122 504 22154
rect 544 22122 576 22154
rect 616 22122 648 22154
rect 688 22122 720 22154
rect 760 22122 792 22154
rect 832 22122 864 22154
rect 904 22122 936 22154
rect 976 22122 1008 22154
rect 1048 22122 1080 22154
rect 1120 22122 1152 22154
rect 1192 22122 1224 22154
rect 1264 22122 1296 22154
rect 1336 22122 1368 22154
rect 1408 22122 1440 22154
rect 1480 22122 1512 22154
rect 1552 22122 1584 22154
rect 1624 22122 1656 22154
rect 1696 22122 1728 22154
rect 1768 22122 1800 22154
rect 1840 22122 1872 22154
rect 1912 22122 1944 22154
rect 1984 22122 2016 22154
rect 2056 22122 2088 22154
rect 2128 22122 2160 22154
rect 2200 22122 2232 22154
rect 2272 22122 2304 22154
rect 2344 22122 2376 22154
rect 2416 22122 2448 22154
rect 2488 22122 2520 22154
rect 2560 22122 2592 22154
rect 2632 22122 2664 22154
rect 2704 22122 2736 22154
rect 2776 22122 2808 22154
rect 2848 22122 2880 22154
rect 2920 22122 2952 22154
rect 2992 22122 3024 22154
rect 3064 22122 3096 22154
rect 3136 22122 3168 22154
rect 3208 22122 3240 22154
rect 3280 22122 3312 22154
rect 3352 22122 3384 22154
rect 3424 22122 3456 22154
rect 3496 22122 3528 22154
rect 3568 22122 3600 22154
rect 3640 22122 3672 22154
rect 3712 22122 3744 22154
rect 3784 22122 3816 22154
rect 3856 22122 3888 22154
rect 112 22050 144 22082
rect 184 22050 216 22082
rect 256 22050 288 22082
rect 328 22050 360 22082
rect 400 22050 432 22082
rect 472 22050 504 22082
rect 544 22050 576 22082
rect 616 22050 648 22082
rect 688 22050 720 22082
rect 760 22050 792 22082
rect 832 22050 864 22082
rect 904 22050 936 22082
rect 976 22050 1008 22082
rect 1048 22050 1080 22082
rect 1120 22050 1152 22082
rect 1192 22050 1224 22082
rect 1264 22050 1296 22082
rect 1336 22050 1368 22082
rect 1408 22050 1440 22082
rect 1480 22050 1512 22082
rect 1552 22050 1584 22082
rect 1624 22050 1656 22082
rect 1696 22050 1728 22082
rect 1768 22050 1800 22082
rect 1840 22050 1872 22082
rect 1912 22050 1944 22082
rect 1984 22050 2016 22082
rect 2056 22050 2088 22082
rect 2128 22050 2160 22082
rect 2200 22050 2232 22082
rect 2272 22050 2304 22082
rect 2344 22050 2376 22082
rect 2416 22050 2448 22082
rect 2488 22050 2520 22082
rect 2560 22050 2592 22082
rect 2632 22050 2664 22082
rect 2704 22050 2736 22082
rect 2776 22050 2808 22082
rect 2848 22050 2880 22082
rect 2920 22050 2952 22082
rect 2992 22050 3024 22082
rect 3064 22050 3096 22082
rect 3136 22050 3168 22082
rect 3208 22050 3240 22082
rect 3280 22050 3312 22082
rect 3352 22050 3384 22082
rect 3424 22050 3456 22082
rect 3496 22050 3528 22082
rect 3568 22050 3600 22082
rect 3640 22050 3672 22082
rect 3712 22050 3744 22082
rect 3784 22050 3816 22082
rect 3856 22050 3888 22082
rect 112 21978 144 22010
rect 184 21978 216 22010
rect 256 21978 288 22010
rect 328 21978 360 22010
rect 400 21978 432 22010
rect 472 21978 504 22010
rect 544 21978 576 22010
rect 616 21978 648 22010
rect 688 21978 720 22010
rect 760 21978 792 22010
rect 832 21978 864 22010
rect 904 21978 936 22010
rect 976 21978 1008 22010
rect 1048 21978 1080 22010
rect 1120 21978 1152 22010
rect 1192 21978 1224 22010
rect 1264 21978 1296 22010
rect 1336 21978 1368 22010
rect 1408 21978 1440 22010
rect 1480 21978 1512 22010
rect 1552 21978 1584 22010
rect 1624 21978 1656 22010
rect 1696 21978 1728 22010
rect 1768 21978 1800 22010
rect 1840 21978 1872 22010
rect 1912 21978 1944 22010
rect 1984 21978 2016 22010
rect 2056 21978 2088 22010
rect 2128 21978 2160 22010
rect 2200 21978 2232 22010
rect 2272 21978 2304 22010
rect 2344 21978 2376 22010
rect 2416 21978 2448 22010
rect 2488 21978 2520 22010
rect 2560 21978 2592 22010
rect 2632 21978 2664 22010
rect 2704 21978 2736 22010
rect 2776 21978 2808 22010
rect 2848 21978 2880 22010
rect 2920 21978 2952 22010
rect 2992 21978 3024 22010
rect 3064 21978 3096 22010
rect 3136 21978 3168 22010
rect 3208 21978 3240 22010
rect 3280 21978 3312 22010
rect 3352 21978 3384 22010
rect 3424 21978 3456 22010
rect 3496 21978 3528 22010
rect 3568 21978 3600 22010
rect 3640 21978 3672 22010
rect 3712 21978 3744 22010
rect 3784 21978 3816 22010
rect 3856 21978 3888 22010
rect 112 21906 144 21938
rect 184 21906 216 21938
rect 256 21906 288 21938
rect 328 21906 360 21938
rect 400 21906 432 21938
rect 472 21906 504 21938
rect 544 21906 576 21938
rect 616 21906 648 21938
rect 688 21906 720 21938
rect 760 21906 792 21938
rect 832 21906 864 21938
rect 904 21906 936 21938
rect 976 21906 1008 21938
rect 1048 21906 1080 21938
rect 1120 21906 1152 21938
rect 1192 21906 1224 21938
rect 1264 21906 1296 21938
rect 1336 21906 1368 21938
rect 1408 21906 1440 21938
rect 1480 21906 1512 21938
rect 1552 21906 1584 21938
rect 1624 21906 1656 21938
rect 1696 21906 1728 21938
rect 1768 21906 1800 21938
rect 1840 21906 1872 21938
rect 1912 21906 1944 21938
rect 1984 21906 2016 21938
rect 2056 21906 2088 21938
rect 2128 21906 2160 21938
rect 2200 21906 2232 21938
rect 2272 21906 2304 21938
rect 2344 21906 2376 21938
rect 2416 21906 2448 21938
rect 2488 21906 2520 21938
rect 2560 21906 2592 21938
rect 2632 21906 2664 21938
rect 2704 21906 2736 21938
rect 2776 21906 2808 21938
rect 2848 21906 2880 21938
rect 2920 21906 2952 21938
rect 2992 21906 3024 21938
rect 3064 21906 3096 21938
rect 3136 21906 3168 21938
rect 3208 21906 3240 21938
rect 3280 21906 3312 21938
rect 3352 21906 3384 21938
rect 3424 21906 3456 21938
rect 3496 21906 3528 21938
rect 3568 21906 3600 21938
rect 3640 21906 3672 21938
rect 3712 21906 3744 21938
rect 3784 21906 3816 21938
rect 3856 21906 3888 21938
rect 112 21834 144 21866
rect 184 21834 216 21866
rect 256 21834 288 21866
rect 328 21834 360 21866
rect 400 21834 432 21866
rect 472 21834 504 21866
rect 544 21834 576 21866
rect 616 21834 648 21866
rect 688 21834 720 21866
rect 760 21834 792 21866
rect 832 21834 864 21866
rect 904 21834 936 21866
rect 976 21834 1008 21866
rect 1048 21834 1080 21866
rect 1120 21834 1152 21866
rect 1192 21834 1224 21866
rect 1264 21834 1296 21866
rect 1336 21834 1368 21866
rect 1408 21834 1440 21866
rect 1480 21834 1512 21866
rect 1552 21834 1584 21866
rect 1624 21834 1656 21866
rect 1696 21834 1728 21866
rect 1768 21834 1800 21866
rect 1840 21834 1872 21866
rect 1912 21834 1944 21866
rect 1984 21834 2016 21866
rect 2056 21834 2088 21866
rect 2128 21834 2160 21866
rect 2200 21834 2232 21866
rect 2272 21834 2304 21866
rect 2344 21834 2376 21866
rect 2416 21834 2448 21866
rect 2488 21834 2520 21866
rect 2560 21834 2592 21866
rect 2632 21834 2664 21866
rect 2704 21834 2736 21866
rect 2776 21834 2808 21866
rect 2848 21834 2880 21866
rect 2920 21834 2952 21866
rect 2992 21834 3024 21866
rect 3064 21834 3096 21866
rect 3136 21834 3168 21866
rect 3208 21834 3240 21866
rect 3280 21834 3312 21866
rect 3352 21834 3384 21866
rect 3424 21834 3456 21866
rect 3496 21834 3528 21866
rect 3568 21834 3600 21866
rect 3640 21834 3672 21866
rect 3712 21834 3744 21866
rect 3784 21834 3816 21866
rect 3856 21834 3888 21866
rect 112 21762 144 21794
rect 184 21762 216 21794
rect 256 21762 288 21794
rect 328 21762 360 21794
rect 400 21762 432 21794
rect 472 21762 504 21794
rect 544 21762 576 21794
rect 616 21762 648 21794
rect 688 21762 720 21794
rect 760 21762 792 21794
rect 832 21762 864 21794
rect 904 21762 936 21794
rect 976 21762 1008 21794
rect 1048 21762 1080 21794
rect 1120 21762 1152 21794
rect 1192 21762 1224 21794
rect 1264 21762 1296 21794
rect 1336 21762 1368 21794
rect 1408 21762 1440 21794
rect 1480 21762 1512 21794
rect 1552 21762 1584 21794
rect 1624 21762 1656 21794
rect 1696 21762 1728 21794
rect 1768 21762 1800 21794
rect 1840 21762 1872 21794
rect 1912 21762 1944 21794
rect 1984 21762 2016 21794
rect 2056 21762 2088 21794
rect 2128 21762 2160 21794
rect 2200 21762 2232 21794
rect 2272 21762 2304 21794
rect 2344 21762 2376 21794
rect 2416 21762 2448 21794
rect 2488 21762 2520 21794
rect 2560 21762 2592 21794
rect 2632 21762 2664 21794
rect 2704 21762 2736 21794
rect 2776 21762 2808 21794
rect 2848 21762 2880 21794
rect 2920 21762 2952 21794
rect 2992 21762 3024 21794
rect 3064 21762 3096 21794
rect 3136 21762 3168 21794
rect 3208 21762 3240 21794
rect 3280 21762 3312 21794
rect 3352 21762 3384 21794
rect 3424 21762 3456 21794
rect 3496 21762 3528 21794
rect 3568 21762 3600 21794
rect 3640 21762 3672 21794
rect 3712 21762 3744 21794
rect 3784 21762 3816 21794
rect 3856 21762 3888 21794
rect 112 21690 144 21722
rect 184 21690 216 21722
rect 256 21690 288 21722
rect 328 21690 360 21722
rect 400 21690 432 21722
rect 472 21690 504 21722
rect 544 21690 576 21722
rect 616 21690 648 21722
rect 688 21690 720 21722
rect 760 21690 792 21722
rect 832 21690 864 21722
rect 904 21690 936 21722
rect 976 21690 1008 21722
rect 1048 21690 1080 21722
rect 1120 21690 1152 21722
rect 1192 21690 1224 21722
rect 1264 21690 1296 21722
rect 1336 21690 1368 21722
rect 1408 21690 1440 21722
rect 1480 21690 1512 21722
rect 1552 21690 1584 21722
rect 1624 21690 1656 21722
rect 1696 21690 1728 21722
rect 1768 21690 1800 21722
rect 1840 21690 1872 21722
rect 1912 21690 1944 21722
rect 1984 21690 2016 21722
rect 2056 21690 2088 21722
rect 2128 21690 2160 21722
rect 2200 21690 2232 21722
rect 2272 21690 2304 21722
rect 2344 21690 2376 21722
rect 2416 21690 2448 21722
rect 2488 21690 2520 21722
rect 2560 21690 2592 21722
rect 2632 21690 2664 21722
rect 2704 21690 2736 21722
rect 2776 21690 2808 21722
rect 2848 21690 2880 21722
rect 2920 21690 2952 21722
rect 2992 21690 3024 21722
rect 3064 21690 3096 21722
rect 3136 21690 3168 21722
rect 3208 21690 3240 21722
rect 3280 21690 3312 21722
rect 3352 21690 3384 21722
rect 3424 21690 3456 21722
rect 3496 21690 3528 21722
rect 3568 21690 3600 21722
rect 3640 21690 3672 21722
rect 3712 21690 3744 21722
rect 3784 21690 3816 21722
rect 3856 21690 3888 21722
rect 112 21618 144 21650
rect 184 21618 216 21650
rect 256 21618 288 21650
rect 328 21618 360 21650
rect 400 21618 432 21650
rect 472 21618 504 21650
rect 544 21618 576 21650
rect 616 21618 648 21650
rect 688 21618 720 21650
rect 760 21618 792 21650
rect 832 21618 864 21650
rect 904 21618 936 21650
rect 976 21618 1008 21650
rect 1048 21618 1080 21650
rect 1120 21618 1152 21650
rect 1192 21618 1224 21650
rect 1264 21618 1296 21650
rect 1336 21618 1368 21650
rect 1408 21618 1440 21650
rect 1480 21618 1512 21650
rect 1552 21618 1584 21650
rect 1624 21618 1656 21650
rect 1696 21618 1728 21650
rect 1768 21618 1800 21650
rect 1840 21618 1872 21650
rect 1912 21618 1944 21650
rect 1984 21618 2016 21650
rect 2056 21618 2088 21650
rect 2128 21618 2160 21650
rect 2200 21618 2232 21650
rect 2272 21618 2304 21650
rect 2344 21618 2376 21650
rect 2416 21618 2448 21650
rect 2488 21618 2520 21650
rect 2560 21618 2592 21650
rect 2632 21618 2664 21650
rect 2704 21618 2736 21650
rect 2776 21618 2808 21650
rect 2848 21618 2880 21650
rect 2920 21618 2952 21650
rect 2992 21618 3024 21650
rect 3064 21618 3096 21650
rect 3136 21618 3168 21650
rect 3208 21618 3240 21650
rect 3280 21618 3312 21650
rect 3352 21618 3384 21650
rect 3424 21618 3456 21650
rect 3496 21618 3528 21650
rect 3568 21618 3600 21650
rect 3640 21618 3672 21650
rect 3712 21618 3744 21650
rect 3784 21618 3816 21650
rect 3856 21618 3888 21650
rect 112 21546 144 21578
rect 184 21546 216 21578
rect 256 21546 288 21578
rect 328 21546 360 21578
rect 400 21546 432 21578
rect 472 21546 504 21578
rect 544 21546 576 21578
rect 616 21546 648 21578
rect 688 21546 720 21578
rect 760 21546 792 21578
rect 832 21546 864 21578
rect 904 21546 936 21578
rect 976 21546 1008 21578
rect 1048 21546 1080 21578
rect 1120 21546 1152 21578
rect 1192 21546 1224 21578
rect 1264 21546 1296 21578
rect 1336 21546 1368 21578
rect 1408 21546 1440 21578
rect 1480 21546 1512 21578
rect 1552 21546 1584 21578
rect 1624 21546 1656 21578
rect 1696 21546 1728 21578
rect 1768 21546 1800 21578
rect 1840 21546 1872 21578
rect 1912 21546 1944 21578
rect 1984 21546 2016 21578
rect 2056 21546 2088 21578
rect 2128 21546 2160 21578
rect 2200 21546 2232 21578
rect 2272 21546 2304 21578
rect 2344 21546 2376 21578
rect 2416 21546 2448 21578
rect 2488 21546 2520 21578
rect 2560 21546 2592 21578
rect 2632 21546 2664 21578
rect 2704 21546 2736 21578
rect 2776 21546 2808 21578
rect 2848 21546 2880 21578
rect 2920 21546 2952 21578
rect 2992 21546 3024 21578
rect 3064 21546 3096 21578
rect 3136 21546 3168 21578
rect 3208 21546 3240 21578
rect 3280 21546 3312 21578
rect 3352 21546 3384 21578
rect 3424 21546 3456 21578
rect 3496 21546 3528 21578
rect 3568 21546 3600 21578
rect 3640 21546 3672 21578
rect 3712 21546 3744 21578
rect 3784 21546 3816 21578
rect 3856 21546 3888 21578
rect 112 21474 144 21506
rect 184 21474 216 21506
rect 256 21474 288 21506
rect 328 21474 360 21506
rect 400 21474 432 21506
rect 472 21474 504 21506
rect 544 21474 576 21506
rect 616 21474 648 21506
rect 688 21474 720 21506
rect 760 21474 792 21506
rect 832 21474 864 21506
rect 904 21474 936 21506
rect 976 21474 1008 21506
rect 1048 21474 1080 21506
rect 1120 21474 1152 21506
rect 1192 21474 1224 21506
rect 1264 21474 1296 21506
rect 1336 21474 1368 21506
rect 1408 21474 1440 21506
rect 1480 21474 1512 21506
rect 1552 21474 1584 21506
rect 1624 21474 1656 21506
rect 1696 21474 1728 21506
rect 1768 21474 1800 21506
rect 1840 21474 1872 21506
rect 1912 21474 1944 21506
rect 1984 21474 2016 21506
rect 2056 21474 2088 21506
rect 2128 21474 2160 21506
rect 2200 21474 2232 21506
rect 2272 21474 2304 21506
rect 2344 21474 2376 21506
rect 2416 21474 2448 21506
rect 2488 21474 2520 21506
rect 2560 21474 2592 21506
rect 2632 21474 2664 21506
rect 2704 21474 2736 21506
rect 2776 21474 2808 21506
rect 2848 21474 2880 21506
rect 2920 21474 2952 21506
rect 2992 21474 3024 21506
rect 3064 21474 3096 21506
rect 3136 21474 3168 21506
rect 3208 21474 3240 21506
rect 3280 21474 3312 21506
rect 3352 21474 3384 21506
rect 3424 21474 3456 21506
rect 3496 21474 3528 21506
rect 3568 21474 3600 21506
rect 3640 21474 3672 21506
rect 3712 21474 3744 21506
rect 3784 21474 3816 21506
rect 3856 21474 3888 21506
rect 112 21402 144 21434
rect 184 21402 216 21434
rect 256 21402 288 21434
rect 328 21402 360 21434
rect 400 21402 432 21434
rect 472 21402 504 21434
rect 544 21402 576 21434
rect 616 21402 648 21434
rect 688 21402 720 21434
rect 760 21402 792 21434
rect 832 21402 864 21434
rect 904 21402 936 21434
rect 976 21402 1008 21434
rect 1048 21402 1080 21434
rect 1120 21402 1152 21434
rect 1192 21402 1224 21434
rect 1264 21402 1296 21434
rect 1336 21402 1368 21434
rect 1408 21402 1440 21434
rect 1480 21402 1512 21434
rect 1552 21402 1584 21434
rect 1624 21402 1656 21434
rect 1696 21402 1728 21434
rect 1768 21402 1800 21434
rect 1840 21402 1872 21434
rect 1912 21402 1944 21434
rect 1984 21402 2016 21434
rect 2056 21402 2088 21434
rect 2128 21402 2160 21434
rect 2200 21402 2232 21434
rect 2272 21402 2304 21434
rect 2344 21402 2376 21434
rect 2416 21402 2448 21434
rect 2488 21402 2520 21434
rect 2560 21402 2592 21434
rect 2632 21402 2664 21434
rect 2704 21402 2736 21434
rect 2776 21402 2808 21434
rect 2848 21402 2880 21434
rect 2920 21402 2952 21434
rect 2992 21402 3024 21434
rect 3064 21402 3096 21434
rect 3136 21402 3168 21434
rect 3208 21402 3240 21434
rect 3280 21402 3312 21434
rect 3352 21402 3384 21434
rect 3424 21402 3456 21434
rect 3496 21402 3528 21434
rect 3568 21402 3600 21434
rect 3640 21402 3672 21434
rect 3712 21402 3744 21434
rect 3784 21402 3816 21434
rect 3856 21402 3888 21434
rect 112 21330 144 21362
rect 184 21330 216 21362
rect 256 21330 288 21362
rect 328 21330 360 21362
rect 400 21330 432 21362
rect 472 21330 504 21362
rect 544 21330 576 21362
rect 616 21330 648 21362
rect 688 21330 720 21362
rect 760 21330 792 21362
rect 832 21330 864 21362
rect 904 21330 936 21362
rect 976 21330 1008 21362
rect 1048 21330 1080 21362
rect 1120 21330 1152 21362
rect 1192 21330 1224 21362
rect 1264 21330 1296 21362
rect 1336 21330 1368 21362
rect 1408 21330 1440 21362
rect 1480 21330 1512 21362
rect 1552 21330 1584 21362
rect 1624 21330 1656 21362
rect 1696 21330 1728 21362
rect 1768 21330 1800 21362
rect 1840 21330 1872 21362
rect 1912 21330 1944 21362
rect 1984 21330 2016 21362
rect 2056 21330 2088 21362
rect 2128 21330 2160 21362
rect 2200 21330 2232 21362
rect 2272 21330 2304 21362
rect 2344 21330 2376 21362
rect 2416 21330 2448 21362
rect 2488 21330 2520 21362
rect 2560 21330 2592 21362
rect 2632 21330 2664 21362
rect 2704 21330 2736 21362
rect 2776 21330 2808 21362
rect 2848 21330 2880 21362
rect 2920 21330 2952 21362
rect 2992 21330 3024 21362
rect 3064 21330 3096 21362
rect 3136 21330 3168 21362
rect 3208 21330 3240 21362
rect 3280 21330 3312 21362
rect 3352 21330 3384 21362
rect 3424 21330 3456 21362
rect 3496 21330 3528 21362
rect 3568 21330 3600 21362
rect 3640 21330 3672 21362
rect 3712 21330 3744 21362
rect 3784 21330 3816 21362
rect 3856 21330 3888 21362
rect 112 21258 144 21290
rect 184 21258 216 21290
rect 256 21258 288 21290
rect 328 21258 360 21290
rect 400 21258 432 21290
rect 472 21258 504 21290
rect 544 21258 576 21290
rect 616 21258 648 21290
rect 688 21258 720 21290
rect 760 21258 792 21290
rect 832 21258 864 21290
rect 904 21258 936 21290
rect 976 21258 1008 21290
rect 1048 21258 1080 21290
rect 1120 21258 1152 21290
rect 1192 21258 1224 21290
rect 1264 21258 1296 21290
rect 1336 21258 1368 21290
rect 1408 21258 1440 21290
rect 1480 21258 1512 21290
rect 1552 21258 1584 21290
rect 1624 21258 1656 21290
rect 1696 21258 1728 21290
rect 1768 21258 1800 21290
rect 1840 21258 1872 21290
rect 1912 21258 1944 21290
rect 1984 21258 2016 21290
rect 2056 21258 2088 21290
rect 2128 21258 2160 21290
rect 2200 21258 2232 21290
rect 2272 21258 2304 21290
rect 2344 21258 2376 21290
rect 2416 21258 2448 21290
rect 2488 21258 2520 21290
rect 2560 21258 2592 21290
rect 2632 21258 2664 21290
rect 2704 21258 2736 21290
rect 2776 21258 2808 21290
rect 2848 21258 2880 21290
rect 2920 21258 2952 21290
rect 2992 21258 3024 21290
rect 3064 21258 3096 21290
rect 3136 21258 3168 21290
rect 3208 21258 3240 21290
rect 3280 21258 3312 21290
rect 3352 21258 3384 21290
rect 3424 21258 3456 21290
rect 3496 21258 3528 21290
rect 3568 21258 3600 21290
rect 3640 21258 3672 21290
rect 3712 21258 3744 21290
rect 3784 21258 3816 21290
rect 3856 21258 3888 21290
rect 112 21186 144 21218
rect 184 21186 216 21218
rect 256 21186 288 21218
rect 328 21186 360 21218
rect 400 21186 432 21218
rect 472 21186 504 21218
rect 544 21186 576 21218
rect 616 21186 648 21218
rect 688 21186 720 21218
rect 760 21186 792 21218
rect 832 21186 864 21218
rect 904 21186 936 21218
rect 976 21186 1008 21218
rect 1048 21186 1080 21218
rect 1120 21186 1152 21218
rect 1192 21186 1224 21218
rect 1264 21186 1296 21218
rect 1336 21186 1368 21218
rect 1408 21186 1440 21218
rect 1480 21186 1512 21218
rect 1552 21186 1584 21218
rect 1624 21186 1656 21218
rect 1696 21186 1728 21218
rect 1768 21186 1800 21218
rect 1840 21186 1872 21218
rect 1912 21186 1944 21218
rect 1984 21186 2016 21218
rect 2056 21186 2088 21218
rect 2128 21186 2160 21218
rect 2200 21186 2232 21218
rect 2272 21186 2304 21218
rect 2344 21186 2376 21218
rect 2416 21186 2448 21218
rect 2488 21186 2520 21218
rect 2560 21186 2592 21218
rect 2632 21186 2664 21218
rect 2704 21186 2736 21218
rect 2776 21186 2808 21218
rect 2848 21186 2880 21218
rect 2920 21186 2952 21218
rect 2992 21186 3024 21218
rect 3064 21186 3096 21218
rect 3136 21186 3168 21218
rect 3208 21186 3240 21218
rect 3280 21186 3312 21218
rect 3352 21186 3384 21218
rect 3424 21186 3456 21218
rect 3496 21186 3528 21218
rect 3568 21186 3600 21218
rect 3640 21186 3672 21218
rect 3712 21186 3744 21218
rect 3784 21186 3816 21218
rect 3856 21186 3888 21218
rect 112 21114 144 21146
rect 184 21114 216 21146
rect 256 21114 288 21146
rect 328 21114 360 21146
rect 400 21114 432 21146
rect 472 21114 504 21146
rect 544 21114 576 21146
rect 616 21114 648 21146
rect 688 21114 720 21146
rect 760 21114 792 21146
rect 832 21114 864 21146
rect 904 21114 936 21146
rect 976 21114 1008 21146
rect 1048 21114 1080 21146
rect 1120 21114 1152 21146
rect 1192 21114 1224 21146
rect 1264 21114 1296 21146
rect 1336 21114 1368 21146
rect 1408 21114 1440 21146
rect 1480 21114 1512 21146
rect 1552 21114 1584 21146
rect 1624 21114 1656 21146
rect 1696 21114 1728 21146
rect 1768 21114 1800 21146
rect 1840 21114 1872 21146
rect 1912 21114 1944 21146
rect 1984 21114 2016 21146
rect 2056 21114 2088 21146
rect 2128 21114 2160 21146
rect 2200 21114 2232 21146
rect 2272 21114 2304 21146
rect 2344 21114 2376 21146
rect 2416 21114 2448 21146
rect 2488 21114 2520 21146
rect 2560 21114 2592 21146
rect 2632 21114 2664 21146
rect 2704 21114 2736 21146
rect 2776 21114 2808 21146
rect 2848 21114 2880 21146
rect 2920 21114 2952 21146
rect 2992 21114 3024 21146
rect 3064 21114 3096 21146
rect 3136 21114 3168 21146
rect 3208 21114 3240 21146
rect 3280 21114 3312 21146
rect 3352 21114 3384 21146
rect 3424 21114 3456 21146
rect 3496 21114 3528 21146
rect 3568 21114 3600 21146
rect 3640 21114 3672 21146
rect 3712 21114 3744 21146
rect 3784 21114 3816 21146
rect 3856 21114 3888 21146
rect 112 21042 144 21074
rect 184 21042 216 21074
rect 256 21042 288 21074
rect 328 21042 360 21074
rect 400 21042 432 21074
rect 472 21042 504 21074
rect 544 21042 576 21074
rect 616 21042 648 21074
rect 688 21042 720 21074
rect 760 21042 792 21074
rect 832 21042 864 21074
rect 904 21042 936 21074
rect 976 21042 1008 21074
rect 1048 21042 1080 21074
rect 1120 21042 1152 21074
rect 1192 21042 1224 21074
rect 1264 21042 1296 21074
rect 1336 21042 1368 21074
rect 1408 21042 1440 21074
rect 1480 21042 1512 21074
rect 1552 21042 1584 21074
rect 1624 21042 1656 21074
rect 1696 21042 1728 21074
rect 1768 21042 1800 21074
rect 1840 21042 1872 21074
rect 1912 21042 1944 21074
rect 1984 21042 2016 21074
rect 2056 21042 2088 21074
rect 2128 21042 2160 21074
rect 2200 21042 2232 21074
rect 2272 21042 2304 21074
rect 2344 21042 2376 21074
rect 2416 21042 2448 21074
rect 2488 21042 2520 21074
rect 2560 21042 2592 21074
rect 2632 21042 2664 21074
rect 2704 21042 2736 21074
rect 2776 21042 2808 21074
rect 2848 21042 2880 21074
rect 2920 21042 2952 21074
rect 2992 21042 3024 21074
rect 3064 21042 3096 21074
rect 3136 21042 3168 21074
rect 3208 21042 3240 21074
rect 3280 21042 3312 21074
rect 3352 21042 3384 21074
rect 3424 21042 3456 21074
rect 3496 21042 3528 21074
rect 3568 21042 3600 21074
rect 3640 21042 3672 21074
rect 3712 21042 3744 21074
rect 3784 21042 3816 21074
rect 3856 21042 3888 21074
rect 112 20970 144 21002
rect 184 20970 216 21002
rect 256 20970 288 21002
rect 328 20970 360 21002
rect 400 20970 432 21002
rect 472 20970 504 21002
rect 544 20970 576 21002
rect 616 20970 648 21002
rect 688 20970 720 21002
rect 760 20970 792 21002
rect 832 20970 864 21002
rect 904 20970 936 21002
rect 976 20970 1008 21002
rect 1048 20970 1080 21002
rect 1120 20970 1152 21002
rect 1192 20970 1224 21002
rect 1264 20970 1296 21002
rect 1336 20970 1368 21002
rect 1408 20970 1440 21002
rect 1480 20970 1512 21002
rect 1552 20970 1584 21002
rect 1624 20970 1656 21002
rect 1696 20970 1728 21002
rect 1768 20970 1800 21002
rect 1840 20970 1872 21002
rect 1912 20970 1944 21002
rect 1984 20970 2016 21002
rect 2056 20970 2088 21002
rect 2128 20970 2160 21002
rect 2200 20970 2232 21002
rect 2272 20970 2304 21002
rect 2344 20970 2376 21002
rect 2416 20970 2448 21002
rect 2488 20970 2520 21002
rect 2560 20970 2592 21002
rect 2632 20970 2664 21002
rect 2704 20970 2736 21002
rect 2776 20970 2808 21002
rect 2848 20970 2880 21002
rect 2920 20970 2952 21002
rect 2992 20970 3024 21002
rect 3064 20970 3096 21002
rect 3136 20970 3168 21002
rect 3208 20970 3240 21002
rect 3280 20970 3312 21002
rect 3352 20970 3384 21002
rect 3424 20970 3456 21002
rect 3496 20970 3528 21002
rect 3568 20970 3600 21002
rect 3640 20970 3672 21002
rect 3712 20970 3744 21002
rect 3784 20970 3816 21002
rect 3856 20970 3888 21002
rect 112 20898 144 20930
rect 184 20898 216 20930
rect 256 20898 288 20930
rect 328 20898 360 20930
rect 400 20898 432 20930
rect 472 20898 504 20930
rect 544 20898 576 20930
rect 616 20898 648 20930
rect 688 20898 720 20930
rect 760 20898 792 20930
rect 832 20898 864 20930
rect 904 20898 936 20930
rect 976 20898 1008 20930
rect 1048 20898 1080 20930
rect 1120 20898 1152 20930
rect 1192 20898 1224 20930
rect 1264 20898 1296 20930
rect 1336 20898 1368 20930
rect 1408 20898 1440 20930
rect 1480 20898 1512 20930
rect 1552 20898 1584 20930
rect 1624 20898 1656 20930
rect 1696 20898 1728 20930
rect 1768 20898 1800 20930
rect 1840 20898 1872 20930
rect 1912 20898 1944 20930
rect 1984 20898 2016 20930
rect 2056 20898 2088 20930
rect 2128 20898 2160 20930
rect 2200 20898 2232 20930
rect 2272 20898 2304 20930
rect 2344 20898 2376 20930
rect 2416 20898 2448 20930
rect 2488 20898 2520 20930
rect 2560 20898 2592 20930
rect 2632 20898 2664 20930
rect 2704 20898 2736 20930
rect 2776 20898 2808 20930
rect 2848 20898 2880 20930
rect 2920 20898 2952 20930
rect 2992 20898 3024 20930
rect 3064 20898 3096 20930
rect 3136 20898 3168 20930
rect 3208 20898 3240 20930
rect 3280 20898 3312 20930
rect 3352 20898 3384 20930
rect 3424 20898 3456 20930
rect 3496 20898 3528 20930
rect 3568 20898 3600 20930
rect 3640 20898 3672 20930
rect 3712 20898 3744 20930
rect 3784 20898 3816 20930
rect 3856 20898 3888 20930
rect 112 20826 144 20858
rect 184 20826 216 20858
rect 256 20826 288 20858
rect 328 20826 360 20858
rect 400 20826 432 20858
rect 472 20826 504 20858
rect 544 20826 576 20858
rect 616 20826 648 20858
rect 688 20826 720 20858
rect 760 20826 792 20858
rect 832 20826 864 20858
rect 904 20826 936 20858
rect 976 20826 1008 20858
rect 1048 20826 1080 20858
rect 1120 20826 1152 20858
rect 1192 20826 1224 20858
rect 1264 20826 1296 20858
rect 1336 20826 1368 20858
rect 1408 20826 1440 20858
rect 1480 20826 1512 20858
rect 1552 20826 1584 20858
rect 1624 20826 1656 20858
rect 1696 20826 1728 20858
rect 1768 20826 1800 20858
rect 1840 20826 1872 20858
rect 1912 20826 1944 20858
rect 1984 20826 2016 20858
rect 2056 20826 2088 20858
rect 2128 20826 2160 20858
rect 2200 20826 2232 20858
rect 2272 20826 2304 20858
rect 2344 20826 2376 20858
rect 2416 20826 2448 20858
rect 2488 20826 2520 20858
rect 2560 20826 2592 20858
rect 2632 20826 2664 20858
rect 2704 20826 2736 20858
rect 2776 20826 2808 20858
rect 2848 20826 2880 20858
rect 2920 20826 2952 20858
rect 2992 20826 3024 20858
rect 3064 20826 3096 20858
rect 3136 20826 3168 20858
rect 3208 20826 3240 20858
rect 3280 20826 3312 20858
rect 3352 20826 3384 20858
rect 3424 20826 3456 20858
rect 3496 20826 3528 20858
rect 3568 20826 3600 20858
rect 3640 20826 3672 20858
rect 3712 20826 3744 20858
rect 3784 20826 3816 20858
rect 3856 20826 3888 20858
rect 112 20754 144 20786
rect 184 20754 216 20786
rect 256 20754 288 20786
rect 328 20754 360 20786
rect 400 20754 432 20786
rect 472 20754 504 20786
rect 544 20754 576 20786
rect 616 20754 648 20786
rect 688 20754 720 20786
rect 760 20754 792 20786
rect 832 20754 864 20786
rect 904 20754 936 20786
rect 976 20754 1008 20786
rect 1048 20754 1080 20786
rect 1120 20754 1152 20786
rect 1192 20754 1224 20786
rect 1264 20754 1296 20786
rect 1336 20754 1368 20786
rect 1408 20754 1440 20786
rect 1480 20754 1512 20786
rect 1552 20754 1584 20786
rect 1624 20754 1656 20786
rect 1696 20754 1728 20786
rect 1768 20754 1800 20786
rect 1840 20754 1872 20786
rect 1912 20754 1944 20786
rect 1984 20754 2016 20786
rect 2056 20754 2088 20786
rect 2128 20754 2160 20786
rect 2200 20754 2232 20786
rect 2272 20754 2304 20786
rect 2344 20754 2376 20786
rect 2416 20754 2448 20786
rect 2488 20754 2520 20786
rect 2560 20754 2592 20786
rect 2632 20754 2664 20786
rect 2704 20754 2736 20786
rect 2776 20754 2808 20786
rect 2848 20754 2880 20786
rect 2920 20754 2952 20786
rect 2992 20754 3024 20786
rect 3064 20754 3096 20786
rect 3136 20754 3168 20786
rect 3208 20754 3240 20786
rect 3280 20754 3312 20786
rect 3352 20754 3384 20786
rect 3424 20754 3456 20786
rect 3496 20754 3528 20786
rect 3568 20754 3600 20786
rect 3640 20754 3672 20786
rect 3712 20754 3744 20786
rect 3784 20754 3816 20786
rect 3856 20754 3888 20786
rect 112 20682 144 20714
rect 184 20682 216 20714
rect 256 20682 288 20714
rect 328 20682 360 20714
rect 400 20682 432 20714
rect 472 20682 504 20714
rect 544 20682 576 20714
rect 616 20682 648 20714
rect 688 20682 720 20714
rect 760 20682 792 20714
rect 832 20682 864 20714
rect 904 20682 936 20714
rect 976 20682 1008 20714
rect 1048 20682 1080 20714
rect 1120 20682 1152 20714
rect 1192 20682 1224 20714
rect 1264 20682 1296 20714
rect 1336 20682 1368 20714
rect 1408 20682 1440 20714
rect 1480 20682 1512 20714
rect 1552 20682 1584 20714
rect 1624 20682 1656 20714
rect 1696 20682 1728 20714
rect 1768 20682 1800 20714
rect 1840 20682 1872 20714
rect 1912 20682 1944 20714
rect 1984 20682 2016 20714
rect 2056 20682 2088 20714
rect 2128 20682 2160 20714
rect 2200 20682 2232 20714
rect 2272 20682 2304 20714
rect 2344 20682 2376 20714
rect 2416 20682 2448 20714
rect 2488 20682 2520 20714
rect 2560 20682 2592 20714
rect 2632 20682 2664 20714
rect 2704 20682 2736 20714
rect 2776 20682 2808 20714
rect 2848 20682 2880 20714
rect 2920 20682 2952 20714
rect 2992 20682 3024 20714
rect 3064 20682 3096 20714
rect 3136 20682 3168 20714
rect 3208 20682 3240 20714
rect 3280 20682 3312 20714
rect 3352 20682 3384 20714
rect 3424 20682 3456 20714
rect 3496 20682 3528 20714
rect 3568 20682 3600 20714
rect 3640 20682 3672 20714
rect 3712 20682 3744 20714
rect 3784 20682 3816 20714
rect 3856 20682 3888 20714
rect 112 20610 144 20642
rect 184 20610 216 20642
rect 256 20610 288 20642
rect 328 20610 360 20642
rect 400 20610 432 20642
rect 472 20610 504 20642
rect 544 20610 576 20642
rect 616 20610 648 20642
rect 688 20610 720 20642
rect 760 20610 792 20642
rect 832 20610 864 20642
rect 904 20610 936 20642
rect 976 20610 1008 20642
rect 1048 20610 1080 20642
rect 1120 20610 1152 20642
rect 1192 20610 1224 20642
rect 1264 20610 1296 20642
rect 1336 20610 1368 20642
rect 1408 20610 1440 20642
rect 1480 20610 1512 20642
rect 1552 20610 1584 20642
rect 1624 20610 1656 20642
rect 1696 20610 1728 20642
rect 1768 20610 1800 20642
rect 1840 20610 1872 20642
rect 1912 20610 1944 20642
rect 1984 20610 2016 20642
rect 2056 20610 2088 20642
rect 2128 20610 2160 20642
rect 2200 20610 2232 20642
rect 2272 20610 2304 20642
rect 2344 20610 2376 20642
rect 2416 20610 2448 20642
rect 2488 20610 2520 20642
rect 2560 20610 2592 20642
rect 2632 20610 2664 20642
rect 2704 20610 2736 20642
rect 2776 20610 2808 20642
rect 2848 20610 2880 20642
rect 2920 20610 2952 20642
rect 2992 20610 3024 20642
rect 3064 20610 3096 20642
rect 3136 20610 3168 20642
rect 3208 20610 3240 20642
rect 3280 20610 3312 20642
rect 3352 20610 3384 20642
rect 3424 20610 3456 20642
rect 3496 20610 3528 20642
rect 3568 20610 3600 20642
rect 3640 20610 3672 20642
rect 3712 20610 3744 20642
rect 3784 20610 3816 20642
rect 3856 20610 3888 20642
rect 112 20538 144 20570
rect 184 20538 216 20570
rect 256 20538 288 20570
rect 328 20538 360 20570
rect 400 20538 432 20570
rect 472 20538 504 20570
rect 544 20538 576 20570
rect 616 20538 648 20570
rect 688 20538 720 20570
rect 760 20538 792 20570
rect 832 20538 864 20570
rect 904 20538 936 20570
rect 976 20538 1008 20570
rect 1048 20538 1080 20570
rect 1120 20538 1152 20570
rect 1192 20538 1224 20570
rect 1264 20538 1296 20570
rect 1336 20538 1368 20570
rect 1408 20538 1440 20570
rect 1480 20538 1512 20570
rect 1552 20538 1584 20570
rect 1624 20538 1656 20570
rect 1696 20538 1728 20570
rect 1768 20538 1800 20570
rect 1840 20538 1872 20570
rect 1912 20538 1944 20570
rect 1984 20538 2016 20570
rect 2056 20538 2088 20570
rect 2128 20538 2160 20570
rect 2200 20538 2232 20570
rect 2272 20538 2304 20570
rect 2344 20538 2376 20570
rect 2416 20538 2448 20570
rect 2488 20538 2520 20570
rect 2560 20538 2592 20570
rect 2632 20538 2664 20570
rect 2704 20538 2736 20570
rect 2776 20538 2808 20570
rect 2848 20538 2880 20570
rect 2920 20538 2952 20570
rect 2992 20538 3024 20570
rect 3064 20538 3096 20570
rect 3136 20538 3168 20570
rect 3208 20538 3240 20570
rect 3280 20538 3312 20570
rect 3352 20538 3384 20570
rect 3424 20538 3456 20570
rect 3496 20538 3528 20570
rect 3568 20538 3600 20570
rect 3640 20538 3672 20570
rect 3712 20538 3744 20570
rect 3784 20538 3816 20570
rect 3856 20538 3888 20570
rect 112 20466 144 20498
rect 184 20466 216 20498
rect 256 20466 288 20498
rect 328 20466 360 20498
rect 400 20466 432 20498
rect 472 20466 504 20498
rect 544 20466 576 20498
rect 616 20466 648 20498
rect 688 20466 720 20498
rect 760 20466 792 20498
rect 832 20466 864 20498
rect 904 20466 936 20498
rect 976 20466 1008 20498
rect 1048 20466 1080 20498
rect 1120 20466 1152 20498
rect 1192 20466 1224 20498
rect 1264 20466 1296 20498
rect 1336 20466 1368 20498
rect 1408 20466 1440 20498
rect 1480 20466 1512 20498
rect 1552 20466 1584 20498
rect 1624 20466 1656 20498
rect 1696 20466 1728 20498
rect 1768 20466 1800 20498
rect 1840 20466 1872 20498
rect 1912 20466 1944 20498
rect 1984 20466 2016 20498
rect 2056 20466 2088 20498
rect 2128 20466 2160 20498
rect 2200 20466 2232 20498
rect 2272 20466 2304 20498
rect 2344 20466 2376 20498
rect 2416 20466 2448 20498
rect 2488 20466 2520 20498
rect 2560 20466 2592 20498
rect 2632 20466 2664 20498
rect 2704 20466 2736 20498
rect 2776 20466 2808 20498
rect 2848 20466 2880 20498
rect 2920 20466 2952 20498
rect 2992 20466 3024 20498
rect 3064 20466 3096 20498
rect 3136 20466 3168 20498
rect 3208 20466 3240 20498
rect 3280 20466 3312 20498
rect 3352 20466 3384 20498
rect 3424 20466 3456 20498
rect 3496 20466 3528 20498
rect 3568 20466 3600 20498
rect 3640 20466 3672 20498
rect 3712 20466 3744 20498
rect 3784 20466 3816 20498
rect 3856 20466 3888 20498
rect 112 20394 144 20426
rect 184 20394 216 20426
rect 256 20394 288 20426
rect 328 20394 360 20426
rect 400 20394 432 20426
rect 472 20394 504 20426
rect 544 20394 576 20426
rect 616 20394 648 20426
rect 688 20394 720 20426
rect 760 20394 792 20426
rect 832 20394 864 20426
rect 904 20394 936 20426
rect 976 20394 1008 20426
rect 1048 20394 1080 20426
rect 1120 20394 1152 20426
rect 1192 20394 1224 20426
rect 1264 20394 1296 20426
rect 1336 20394 1368 20426
rect 1408 20394 1440 20426
rect 1480 20394 1512 20426
rect 1552 20394 1584 20426
rect 1624 20394 1656 20426
rect 1696 20394 1728 20426
rect 1768 20394 1800 20426
rect 1840 20394 1872 20426
rect 1912 20394 1944 20426
rect 1984 20394 2016 20426
rect 2056 20394 2088 20426
rect 2128 20394 2160 20426
rect 2200 20394 2232 20426
rect 2272 20394 2304 20426
rect 2344 20394 2376 20426
rect 2416 20394 2448 20426
rect 2488 20394 2520 20426
rect 2560 20394 2592 20426
rect 2632 20394 2664 20426
rect 2704 20394 2736 20426
rect 2776 20394 2808 20426
rect 2848 20394 2880 20426
rect 2920 20394 2952 20426
rect 2992 20394 3024 20426
rect 3064 20394 3096 20426
rect 3136 20394 3168 20426
rect 3208 20394 3240 20426
rect 3280 20394 3312 20426
rect 3352 20394 3384 20426
rect 3424 20394 3456 20426
rect 3496 20394 3528 20426
rect 3568 20394 3600 20426
rect 3640 20394 3672 20426
rect 3712 20394 3744 20426
rect 3784 20394 3816 20426
rect 3856 20394 3888 20426
rect 112 20322 144 20354
rect 184 20322 216 20354
rect 256 20322 288 20354
rect 328 20322 360 20354
rect 400 20322 432 20354
rect 472 20322 504 20354
rect 544 20322 576 20354
rect 616 20322 648 20354
rect 688 20322 720 20354
rect 760 20322 792 20354
rect 832 20322 864 20354
rect 904 20322 936 20354
rect 976 20322 1008 20354
rect 1048 20322 1080 20354
rect 1120 20322 1152 20354
rect 1192 20322 1224 20354
rect 1264 20322 1296 20354
rect 1336 20322 1368 20354
rect 1408 20322 1440 20354
rect 1480 20322 1512 20354
rect 1552 20322 1584 20354
rect 1624 20322 1656 20354
rect 1696 20322 1728 20354
rect 1768 20322 1800 20354
rect 1840 20322 1872 20354
rect 1912 20322 1944 20354
rect 1984 20322 2016 20354
rect 2056 20322 2088 20354
rect 2128 20322 2160 20354
rect 2200 20322 2232 20354
rect 2272 20322 2304 20354
rect 2344 20322 2376 20354
rect 2416 20322 2448 20354
rect 2488 20322 2520 20354
rect 2560 20322 2592 20354
rect 2632 20322 2664 20354
rect 2704 20322 2736 20354
rect 2776 20322 2808 20354
rect 2848 20322 2880 20354
rect 2920 20322 2952 20354
rect 2992 20322 3024 20354
rect 3064 20322 3096 20354
rect 3136 20322 3168 20354
rect 3208 20322 3240 20354
rect 3280 20322 3312 20354
rect 3352 20322 3384 20354
rect 3424 20322 3456 20354
rect 3496 20322 3528 20354
rect 3568 20322 3600 20354
rect 3640 20322 3672 20354
rect 3712 20322 3744 20354
rect 3784 20322 3816 20354
rect 3856 20322 3888 20354
rect 112 20250 144 20282
rect 184 20250 216 20282
rect 256 20250 288 20282
rect 328 20250 360 20282
rect 400 20250 432 20282
rect 472 20250 504 20282
rect 544 20250 576 20282
rect 616 20250 648 20282
rect 688 20250 720 20282
rect 760 20250 792 20282
rect 832 20250 864 20282
rect 904 20250 936 20282
rect 976 20250 1008 20282
rect 1048 20250 1080 20282
rect 1120 20250 1152 20282
rect 1192 20250 1224 20282
rect 1264 20250 1296 20282
rect 1336 20250 1368 20282
rect 1408 20250 1440 20282
rect 1480 20250 1512 20282
rect 1552 20250 1584 20282
rect 1624 20250 1656 20282
rect 1696 20250 1728 20282
rect 1768 20250 1800 20282
rect 1840 20250 1872 20282
rect 1912 20250 1944 20282
rect 1984 20250 2016 20282
rect 2056 20250 2088 20282
rect 2128 20250 2160 20282
rect 2200 20250 2232 20282
rect 2272 20250 2304 20282
rect 2344 20250 2376 20282
rect 2416 20250 2448 20282
rect 2488 20250 2520 20282
rect 2560 20250 2592 20282
rect 2632 20250 2664 20282
rect 2704 20250 2736 20282
rect 2776 20250 2808 20282
rect 2848 20250 2880 20282
rect 2920 20250 2952 20282
rect 2992 20250 3024 20282
rect 3064 20250 3096 20282
rect 3136 20250 3168 20282
rect 3208 20250 3240 20282
rect 3280 20250 3312 20282
rect 3352 20250 3384 20282
rect 3424 20250 3456 20282
rect 3496 20250 3528 20282
rect 3568 20250 3600 20282
rect 3640 20250 3672 20282
rect 3712 20250 3744 20282
rect 3784 20250 3816 20282
rect 3856 20250 3888 20282
rect 112 20178 144 20210
rect 184 20178 216 20210
rect 256 20178 288 20210
rect 328 20178 360 20210
rect 400 20178 432 20210
rect 472 20178 504 20210
rect 544 20178 576 20210
rect 616 20178 648 20210
rect 688 20178 720 20210
rect 760 20178 792 20210
rect 832 20178 864 20210
rect 904 20178 936 20210
rect 976 20178 1008 20210
rect 1048 20178 1080 20210
rect 1120 20178 1152 20210
rect 1192 20178 1224 20210
rect 1264 20178 1296 20210
rect 1336 20178 1368 20210
rect 1408 20178 1440 20210
rect 1480 20178 1512 20210
rect 1552 20178 1584 20210
rect 1624 20178 1656 20210
rect 1696 20178 1728 20210
rect 1768 20178 1800 20210
rect 1840 20178 1872 20210
rect 1912 20178 1944 20210
rect 1984 20178 2016 20210
rect 2056 20178 2088 20210
rect 2128 20178 2160 20210
rect 2200 20178 2232 20210
rect 2272 20178 2304 20210
rect 2344 20178 2376 20210
rect 2416 20178 2448 20210
rect 2488 20178 2520 20210
rect 2560 20178 2592 20210
rect 2632 20178 2664 20210
rect 2704 20178 2736 20210
rect 2776 20178 2808 20210
rect 2848 20178 2880 20210
rect 2920 20178 2952 20210
rect 2992 20178 3024 20210
rect 3064 20178 3096 20210
rect 3136 20178 3168 20210
rect 3208 20178 3240 20210
rect 3280 20178 3312 20210
rect 3352 20178 3384 20210
rect 3424 20178 3456 20210
rect 3496 20178 3528 20210
rect 3568 20178 3600 20210
rect 3640 20178 3672 20210
rect 3712 20178 3744 20210
rect 3784 20178 3816 20210
rect 3856 20178 3888 20210
rect 112 20106 144 20138
rect 184 20106 216 20138
rect 256 20106 288 20138
rect 328 20106 360 20138
rect 400 20106 432 20138
rect 472 20106 504 20138
rect 544 20106 576 20138
rect 616 20106 648 20138
rect 688 20106 720 20138
rect 760 20106 792 20138
rect 832 20106 864 20138
rect 904 20106 936 20138
rect 976 20106 1008 20138
rect 1048 20106 1080 20138
rect 1120 20106 1152 20138
rect 1192 20106 1224 20138
rect 1264 20106 1296 20138
rect 1336 20106 1368 20138
rect 1408 20106 1440 20138
rect 1480 20106 1512 20138
rect 1552 20106 1584 20138
rect 1624 20106 1656 20138
rect 1696 20106 1728 20138
rect 1768 20106 1800 20138
rect 1840 20106 1872 20138
rect 1912 20106 1944 20138
rect 1984 20106 2016 20138
rect 2056 20106 2088 20138
rect 2128 20106 2160 20138
rect 2200 20106 2232 20138
rect 2272 20106 2304 20138
rect 2344 20106 2376 20138
rect 2416 20106 2448 20138
rect 2488 20106 2520 20138
rect 2560 20106 2592 20138
rect 2632 20106 2664 20138
rect 2704 20106 2736 20138
rect 2776 20106 2808 20138
rect 2848 20106 2880 20138
rect 2920 20106 2952 20138
rect 2992 20106 3024 20138
rect 3064 20106 3096 20138
rect 3136 20106 3168 20138
rect 3208 20106 3240 20138
rect 3280 20106 3312 20138
rect 3352 20106 3384 20138
rect 3424 20106 3456 20138
rect 3496 20106 3528 20138
rect 3568 20106 3600 20138
rect 3640 20106 3672 20138
rect 3712 20106 3744 20138
rect 3784 20106 3816 20138
rect 3856 20106 3888 20138
rect 112 20034 144 20066
rect 184 20034 216 20066
rect 256 20034 288 20066
rect 328 20034 360 20066
rect 400 20034 432 20066
rect 472 20034 504 20066
rect 544 20034 576 20066
rect 616 20034 648 20066
rect 688 20034 720 20066
rect 760 20034 792 20066
rect 832 20034 864 20066
rect 904 20034 936 20066
rect 976 20034 1008 20066
rect 1048 20034 1080 20066
rect 1120 20034 1152 20066
rect 1192 20034 1224 20066
rect 1264 20034 1296 20066
rect 1336 20034 1368 20066
rect 1408 20034 1440 20066
rect 1480 20034 1512 20066
rect 1552 20034 1584 20066
rect 1624 20034 1656 20066
rect 1696 20034 1728 20066
rect 1768 20034 1800 20066
rect 1840 20034 1872 20066
rect 1912 20034 1944 20066
rect 1984 20034 2016 20066
rect 2056 20034 2088 20066
rect 2128 20034 2160 20066
rect 2200 20034 2232 20066
rect 2272 20034 2304 20066
rect 2344 20034 2376 20066
rect 2416 20034 2448 20066
rect 2488 20034 2520 20066
rect 2560 20034 2592 20066
rect 2632 20034 2664 20066
rect 2704 20034 2736 20066
rect 2776 20034 2808 20066
rect 2848 20034 2880 20066
rect 2920 20034 2952 20066
rect 2992 20034 3024 20066
rect 3064 20034 3096 20066
rect 3136 20034 3168 20066
rect 3208 20034 3240 20066
rect 3280 20034 3312 20066
rect 3352 20034 3384 20066
rect 3424 20034 3456 20066
rect 3496 20034 3528 20066
rect 3568 20034 3600 20066
rect 3640 20034 3672 20066
rect 3712 20034 3744 20066
rect 3784 20034 3816 20066
rect 3856 20034 3888 20066
rect 112 19962 144 19994
rect 184 19962 216 19994
rect 256 19962 288 19994
rect 328 19962 360 19994
rect 400 19962 432 19994
rect 472 19962 504 19994
rect 544 19962 576 19994
rect 616 19962 648 19994
rect 688 19962 720 19994
rect 760 19962 792 19994
rect 832 19962 864 19994
rect 904 19962 936 19994
rect 976 19962 1008 19994
rect 1048 19962 1080 19994
rect 1120 19962 1152 19994
rect 1192 19962 1224 19994
rect 1264 19962 1296 19994
rect 1336 19962 1368 19994
rect 1408 19962 1440 19994
rect 1480 19962 1512 19994
rect 1552 19962 1584 19994
rect 1624 19962 1656 19994
rect 1696 19962 1728 19994
rect 1768 19962 1800 19994
rect 1840 19962 1872 19994
rect 1912 19962 1944 19994
rect 1984 19962 2016 19994
rect 2056 19962 2088 19994
rect 2128 19962 2160 19994
rect 2200 19962 2232 19994
rect 2272 19962 2304 19994
rect 2344 19962 2376 19994
rect 2416 19962 2448 19994
rect 2488 19962 2520 19994
rect 2560 19962 2592 19994
rect 2632 19962 2664 19994
rect 2704 19962 2736 19994
rect 2776 19962 2808 19994
rect 2848 19962 2880 19994
rect 2920 19962 2952 19994
rect 2992 19962 3024 19994
rect 3064 19962 3096 19994
rect 3136 19962 3168 19994
rect 3208 19962 3240 19994
rect 3280 19962 3312 19994
rect 3352 19962 3384 19994
rect 3424 19962 3456 19994
rect 3496 19962 3528 19994
rect 3568 19962 3600 19994
rect 3640 19962 3672 19994
rect 3712 19962 3744 19994
rect 3784 19962 3816 19994
rect 3856 19962 3888 19994
rect 112 19890 144 19922
rect 184 19890 216 19922
rect 256 19890 288 19922
rect 328 19890 360 19922
rect 400 19890 432 19922
rect 472 19890 504 19922
rect 544 19890 576 19922
rect 616 19890 648 19922
rect 688 19890 720 19922
rect 760 19890 792 19922
rect 832 19890 864 19922
rect 904 19890 936 19922
rect 976 19890 1008 19922
rect 1048 19890 1080 19922
rect 1120 19890 1152 19922
rect 1192 19890 1224 19922
rect 1264 19890 1296 19922
rect 1336 19890 1368 19922
rect 1408 19890 1440 19922
rect 1480 19890 1512 19922
rect 1552 19890 1584 19922
rect 1624 19890 1656 19922
rect 1696 19890 1728 19922
rect 1768 19890 1800 19922
rect 1840 19890 1872 19922
rect 1912 19890 1944 19922
rect 1984 19890 2016 19922
rect 2056 19890 2088 19922
rect 2128 19890 2160 19922
rect 2200 19890 2232 19922
rect 2272 19890 2304 19922
rect 2344 19890 2376 19922
rect 2416 19890 2448 19922
rect 2488 19890 2520 19922
rect 2560 19890 2592 19922
rect 2632 19890 2664 19922
rect 2704 19890 2736 19922
rect 2776 19890 2808 19922
rect 2848 19890 2880 19922
rect 2920 19890 2952 19922
rect 2992 19890 3024 19922
rect 3064 19890 3096 19922
rect 3136 19890 3168 19922
rect 3208 19890 3240 19922
rect 3280 19890 3312 19922
rect 3352 19890 3384 19922
rect 3424 19890 3456 19922
rect 3496 19890 3528 19922
rect 3568 19890 3600 19922
rect 3640 19890 3672 19922
rect 3712 19890 3744 19922
rect 3784 19890 3816 19922
rect 3856 19890 3888 19922
rect 112 19818 144 19850
rect 184 19818 216 19850
rect 256 19818 288 19850
rect 328 19818 360 19850
rect 400 19818 432 19850
rect 472 19818 504 19850
rect 544 19818 576 19850
rect 616 19818 648 19850
rect 688 19818 720 19850
rect 760 19818 792 19850
rect 832 19818 864 19850
rect 904 19818 936 19850
rect 976 19818 1008 19850
rect 1048 19818 1080 19850
rect 1120 19818 1152 19850
rect 1192 19818 1224 19850
rect 1264 19818 1296 19850
rect 1336 19818 1368 19850
rect 1408 19818 1440 19850
rect 1480 19818 1512 19850
rect 1552 19818 1584 19850
rect 1624 19818 1656 19850
rect 1696 19818 1728 19850
rect 1768 19818 1800 19850
rect 1840 19818 1872 19850
rect 1912 19818 1944 19850
rect 1984 19818 2016 19850
rect 2056 19818 2088 19850
rect 2128 19818 2160 19850
rect 2200 19818 2232 19850
rect 2272 19818 2304 19850
rect 2344 19818 2376 19850
rect 2416 19818 2448 19850
rect 2488 19818 2520 19850
rect 2560 19818 2592 19850
rect 2632 19818 2664 19850
rect 2704 19818 2736 19850
rect 2776 19818 2808 19850
rect 2848 19818 2880 19850
rect 2920 19818 2952 19850
rect 2992 19818 3024 19850
rect 3064 19818 3096 19850
rect 3136 19818 3168 19850
rect 3208 19818 3240 19850
rect 3280 19818 3312 19850
rect 3352 19818 3384 19850
rect 3424 19818 3456 19850
rect 3496 19818 3528 19850
rect 3568 19818 3600 19850
rect 3640 19818 3672 19850
rect 3712 19818 3744 19850
rect 3784 19818 3816 19850
rect 3856 19818 3888 19850
rect 112 19746 144 19778
rect 184 19746 216 19778
rect 256 19746 288 19778
rect 328 19746 360 19778
rect 400 19746 432 19778
rect 472 19746 504 19778
rect 544 19746 576 19778
rect 616 19746 648 19778
rect 688 19746 720 19778
rect 760 19746 792 19778
rect 832 19746 864 19778
rect 904 19746 936 19778
rect 976 19746 1008 19778
rect 1048 19746 1080 19778
rect 1120 19746 1152 19778
rect 1192 19746 1224 19778
rect 1264 19746 1296 19778
rect 1336 19746 1368 19778
rect 1408 19746 1440 19778
rect 1480 19746 1512 19778
rect 1552 19746 1584 19778
rect 1624 19746 1656 19778
rect 1696 19746 1728 19778
rect 1768 19746 1800 19778
rect 1840 19746 1872 19778
rect 1912 19746 1944 19778
rect 1984 19746 2016 19778
rect 2056 19746 2088 19778
rect 2128 19746 2160 19778
rect 2200 19746 2232 19778
rect 2272 19746 2304 19778
rect 2344 19746 2376 19778
rect 2416 19746 2448 19778
rect 2488 19746 2520 19778
rect 2560 19746 2592 19778
rect 2632 19746 2664 19778
rect 2704 19746 2736 19778
rect 2776 19746 2808 19778
rect 2848 19746 2880 19778
rect 2920 19746 2952 19778
rect 2992 19746 3024 19778
rect 3064 19746 3096 19778
rect 3136 19746 3168 19778
rect 3208 19746 3240 19778
rect 3280 19746 3312 19778
rect 3352 19746 3384 19778
rect 3424 19746 3456 19778
rect 3496 19746 3528 19778
rect 3568 19746 3600 19778
rect 3640 19746 3672 19778
rect 3712 19746 3744 19778
rect 3784 19746 3816 19778
rect 3856 19746 3888 19778
rect 112 19674 144 19706
rect 184 19674 216 19706
rect 256 19674 288 19706
rect 328 19674 360 19706
rect 400 19674 432 19706
rect 472 19674 504 19706
rect 544 19674 576 19706
rect 616 19674 648 19706
rect 688 19674 720 19706
rect 760 19674 792 19706
rect 832 19674 864 19706
rect 904 19674 936 19706
rect 976 19674 1008 19706
rect 1048 19674 1080 19706
rect 1120 19674 1152 19706
rect 1192 19674 1224 19706
rect 1264 19674 1296 19706
rect 1336 19674 1368 19706
rect 1408 19674 1440 19706
rect 1480 19674 1512 19706
rect 1552 19674 1584 19706
rect 1624 19674 1656 19706
rect 1696 19674 1728 19706
rect 1768 19674 1800 19706
rect 1840 19674 1872 19706
rect 1912 19674 1944 19706
rect 1984 19674 2016 19706
rect 2056 19674 2088 19706
rect 2128 19674 2160 19706
rect 2200 19674 2232 19706
rect 2272 19674 2304 19706
rect 2344 19674 2376 19706
rect 2416 19674 2448 19706
rect 2488 19674 2520 19706
rect 2560 19674 2592 19706
rect 2632 19674 2664 19706
rect 2704 19674 2736 19706
rect 2776 19674 2808 19706
rect 2848 19674 2880 19706
rect 2920 19674 2952 19706
rect 2992 19674 3024 19706
rect 3064 19674 3096 19706
rect 3136 19674 3168 19706
rect 3208 19674 3240 19706
rect 3280 19674 3312 19706
rect 3352 19674 3384 19706
rect 3424 19674 3456 19706
rect 3496 19674 3528 19706
rect 3568 19674 3600 19706
rect 3640 19674 3672 19706
rect 3712 19674 3744 19706
rect 3784 19674 3816 19706
rect 3856 19674 3888 19706
rect 112 19602 144 19634
rect 184 19602 216 19634
rect 256 19602 288 19634
rect 328 19602 360 19634
rect 400 19602 432 19634
rect 472 19602 504 19634
rect 544 19602 576 19634
rect 616 19602 648 19634
rect 688 19602 720 19634
rect 760 19602 792 19634
rect 832 19602 864 19634
rect 904 19602 936 19634
rect 976 19602 1008 19634
rect 1048 19602 1080 19634
rect 1120 19602 1152 19634
rect 1192 19602 1224 19634
rect 1264 19602 1296 19634
rect 1336 19602 1368 19634
rect 1408 19602 1440 19634
rect 1480 19602 1512 19634
rect 1552 19602 1584 19634
rect 1624 19602 1656 19634
rect 1696 19602 1728 19634
rect 1768 19602 1800 19634
rect 1840 19602 1872 19634
rect 1912 19602 1944 19634
rect 1984 19602 2016 19634
rect 2056 19602 2088 19634
rect 2128 19602 2160 19634
rect 2200 19602 2232 19634
rect 2272 19602 2304 19634
rect 2344 19602 2376 19634
rect 2416 19602 2448 19634
rect 2488 19602 2520 19634
rect 2560 19602 2592 19634
rect 2632 19602 2664 19634
rect 2704 19602 2736 19634
rect 2776 19602 2808 19634
rect 2848 19602 2880 19634
rect 2920 19602 2952 19634
rect 2992 19602 3024 19634
rect 3064 19602 3096 19634
rect 3136 19602 3168 19634
rect 3208 19602 3240 19634
rect 3280 19602 3312 19634
rect 3352 19602 3384 19634
rect 3424 19602 3456 19634
rect 3496 19602 3528 19634
rect 3568 19602 3600 19634
rect 3640 19602 3672 19634
rect 3712 19602 3744 19634
rect 3784 19602 3816 19634
rect 3856 19602 3888 19634
rect 112 19530 144 19562
rect 184 19530 216 19562
rect 256 19530 288 19562
rect 328 19530 360 19562
rect 400 19530 432 19562
rect 472 19530 504 19562
rect 544 19530 576 19562
rect 616 19530 648 19562
rect 688 19530 720 19562
rect 760 19530 792 19562
rect 832 19530 864 19562
rect 904 19530 936 19562
rect 976 19530 1008 19562
rect 1048 19530 1080 19562
rect 1120 19530 1152 19562
rect 1192 19530 1224 19562
rect 1264 19530 1296 19562
rect 1336 19530 1368 19562
rect 1408 19530 1440 19562
rect 1480 19530 1512 19562
rect 1552 19530 1584 19562
rect 1624 19530 1656 19562
rect 1696 19530 1728 19562
rect 1768 19530 1800 19562
rect 1840 19530 1872 19562
rect 1912 19530 1944 19562
rect 1984 19530 2016 19562
rect 2056 19530 2088 19562
rect 2128 19530 2160 19562
rect 2200 19530 2232 19562
rect 2272 19530 2304 19562
rect 2344 19530 2376 19562
rect 2416 19530 2448 19562
rect 2488 19530 2520 19562
rect 2560 19530 2592 19562
rect 2632 19530 2664 19562
rect 2704 19530 2736 19562
rect 2776 19530 2808 19562
rect 2848 19530 2880 19562
rect 2920 19530 2952 19562
rect 2992 19530 3024 19562
rect 3064 19530 3096 19562
rect 3136 19530 3168 19562
rect 3208 19530 3240 19562
rect 3280 19530 3312 19562
rect 3352 19530 3384 19562
rect 3424 19530 3456 19562
rect 3496 19530 3528 19562
rect 3568 19530 3600 19562
rect 3640 19530 3672 19562
rect 3712 19530 3744 19562
rect 3784 19530 3816 19562
rect 3856 19530 3888 19562
rect 112 19458 144 19490
rect 184 19458 216 19490
rect 256 19458 288 19490
rect 328 19458 360 19490
rect 400 19458 432 19490
rect 472 19458 504 19490
rect 544 19458 576 19490
rect 616 19458 648 19490
rect 688 19458 720 19490
rect 760 19458 792 19490
rect 832 19458 864 19490
rect 904 19458 936 19490
rect 976 19458 1008 19490
rect 1048 19458 1080 19490
rect 1120 19458 1152 19490
rect 1192 19458 1224 19490
rect 1264 19458 1296 19490
rect 1336 19458 1368 19490
rect 1408 19458 1440 19490
rect 1480 19458 1512 19490
rect 1552 19458 1584 19490
rect 1624 19458 1656 19490
rect 1696 19458 1728 19490
rect 1768 19458 1800 19490
rect 1840 19458 1872 19490
rect 1912 19458 1944 19490
rect 1984 19458 2016 19490
rect 2056 19458 2088 19490
rect 2128 19458 2160 19490
rect 2200 19458 2232 19490
rect 2272 19458 2304 19490
rect 2344 19458 2376 19490
rect 2416 19458 2448 19490
rect 2488 19458 2520 19490
rect 2560 19458 2592 19490
rect 2632 19458 2664 19490
rect 2704 19458 2736 19490
rect 2776 19458 2808 19490
rect 2848 19458 2880 19490
rect 2920 19458 2952 19490
rect 2992 19458 3024 19490
rect 3064 19458 3096 19490
rect 3136 19458 3168 19490
rect 3208 19458 3240 19490
rect 3280 19458 3312 19490
rect 3352 19458 3384 19490
rect 3424 19458 3456 19490
rect 3496 19458 3528 19490
rect 3568 19458 3600 19490
rect 3640 19458 3672 19490
rect 3712 19458 3744 19490
rect 3784 19458 3816 19490
rect 3856 19458 3888 19490
rect 112 19386 144 19418
rect 184 19386 216 19418
rect 256 19386 288 19418
rect 328 19386 360 19418
rect 400 19386 432 19418
rect 472 19386 504 19418
rect 544 19386 576 19418
rect 616 19386 648 19418
rect 688 19386 720 19418
rect 760 19386 792 19418
rect 832 19386 864 19418
rect 904 19386 936 19418
rect 976 19386 1008 19418
rect 1048 19386 1080 19418
rect 1120 19386 1152 19418
rect 1192 19386 1224 19418
rect 1264 19386 1296 19418
rect 1336 19386 1368 19418
rect 1408 19386 1440 19418
rect 1480 19386 1512 19418
rect 1552 19386 1584 19418
rect 1624 19386 1656 19418
rect 1696 19386 1728 19418
rect 1768 19386 1800 19418
rect 1840 19386 1872 19418
rect 1912 19386 1944 19418
rect 1984 19386 2016 19418
rect 2056 19386 2088 19418
rect 2128 19386 2160 19418
rect 2200 19386 2232 19418
rect 2272 19386 2304 19418
rect 2344 19386 2376 19418
rect 2416 19386 2448 19418
rect 2488 19386 2520 19418
rect 2560 19386 2592 19418
rect 2632 19386 2664 19418
rect 2704 19386 2736 19418
rect 2776 19386 2808 19418
rect 2848 19386 2880 19418
rect 2920 19386 2952 19418
rect 2992 19386 3024 19418
rect 3064 19386 3096 19418
rect 3136 19386 3168 19418
rect 3208 19386 3240 19418
rect 3280 19386 3312 19418
rect 3352 19386 3384 19418
rect 3424 19386 3456 19418
rect 3496 19386 3528 19418
rect 3568 19386 3600 19418
rect 3640 19386 3672 19418
rect 3712 19386 3744 19418
rect 3784 19386 3816 19418
rect 3856 19386 3888 19418
rect 112 19314 144 19346
rect 184 19314 216 19346
rect 256 19314 288 19346
rect 328 19314 360 19346
rect 400 19314 432 19346
rect 472 19314 504 19346
rect 544 19314 576 19346
rect 616 19314 648 19346
rect 688 19314 720 19346
rect 760 19314 792 19346
rect 832 19314 864 19346
rect 904 19314 936 19346
rect 976 19314 1008 19346
rect 1048 19314 1080 19346
rect 1120 19314 1152 19346
rect 1192 19314 1224 19346
rect 1264 19314 1296 19346
rect 1336 19314 1368 19346
rect 1408 19314 1440 19346
rect 1480 19314 1512 19346
rect 1552 19314 1584 19346
rect 1624 19314 1656 19346
rect 1696 19314 1728 19346
rect 1768 19314 1800 19346
rect 1840 19314 1872 19346
rect 1912 19314 1944 19346
rect 1984 19314 2016 19346
rect 2056 19314 2088 19346
rect 2128 19314 2160 19346
rect 2200 19314 2232 19346
rect 2272 19314 2304 19346
rect 2344 19314 2376 19346
rect 2416 19314 2448 19346
rect 2488 19314 2520 19346
rect 2560 19314 2592 19346
rect 2632 19314 2664 19346
rect 2704 19314 2736 19346
rect 2776 19314 2808 19346
rect 2848 19314 2880 19346
rect 2920 19314 2952 19346
rect 2992 19314 3024 19346
rect 3064 19314 3096 19346
rect 3136 19314 3168 19346
rect 3208 19314 3240 19346
rect 3280 19314 3312 19346
rect 3352 19314 3384 19346
rect 3424 19314 3456 19346
rect 3496 19314 3528 19346
rect 3568 19314 3600 19346
rect 3640 19314 3672 19346
rect 3712 19314 3744 19346
rect 3784 19314 3816 19346
rect 3856 19314 3888 19346
rect 112 19242 144 19274
rect 184 19242 216 19274
rect 256 19242 288 19274
rect 328 19242 360 19274
rect 400 19242 432 19274
rect 472 19242 504 19274
rect 544 19242 576 19274
rect 616 19242 648 19274
rect 688 19242 720 19274
rect 760 19242 792 19274
rect 832 19242 864 19274
rect 904 19242 936 19274
rect 976 19242 1008 19274
rect 1048 19242 1080 19274
rect 1120 19242 1152 19274
rect 1192 19242 1224 19274
rect 1264 19242 1296 19274
rect 1336 19242 1368 19274
rect 1408 19242 1440 19274
rect 1480 19242 1512 19274
rect 1552 19242 1584 19274
rect 1624 19242 1656 19274
rect 1696 19242 1728 19274
rect 1768 19242 1800 19274
rect 1840 19242 1872 19274
rect 1912 19242 1944 19274
rect 1984 19242 2016 19274
rect 2056 19242 2088 19274
rect 2128 19242 2160 19274
rect 2200 19242 2232 19274
rect 2272 19242 2304 19274
rect 2344 19242 2376 19274
rect 2416 19242 2448 19274
rect 2488 19242 2520 19274
rect 2560 19242 2592 19274
rect 2632 19242 2664 19274
rect 2704 19242 2736 19274
rect 2776 19242 2808 19274
rect 2848 19242 2880 19274
rect 2920 19242 2952 19274
rect 2992 19242 3024 19274
rect 3064 19242 3096 19274
rect 3136 19242 3168 19274
rect 3208 19242 3240 19274
rect 3280 19242 3312 19274
rect 3352 19242 3384 19274
rect 3424 19242 3456 19274
rect 3496 19242 3528 19274
rect 3568 19242 3600 19274
rect 3640 19242 3672 19274
rect 3712 19242 3744 19274
rect 3784 19242 3816 19274
rect 3856 19242 3888 19274
rect 112 19170 144 19202
rect 184 19170 216 19202
rect 256 19170 288 19202
rect 328 19170 360 19202
rect 400 19170 432 19202
rect 472 19170 504 19202
rect 544 19170 576 19202
rect 616 19170 648 19202
rect 688 19170 720 19202
rect 760 19170 792 19202
rect 832 19170 864 19202
rect 904 19170 936 19202
rect 976 19170 1008 19202
rect 1048 19170 1080 19202
rect 1120 19170 1152 19202
rect 1192 19170 1224 19202
rect 1264 19170 1296 19202
rect 1336 19170 1368 19202
rect 1408 19170 1440 19202
rect 1480 19170 1512 19202
rect 1552 19170 1584 19202
rect 1624 19170 1656 19202
rect 1696 19170 1728 19202
rect 1768 19170 1800 19202
rect 1840 19170 1872 19202
rect 1912 19170 1944 19202
rect 1984 19170 2016 19202
rect 2056 19170 2088 19202
rect 2128 19170 2160 19202
rect 2200 19170 2232 19202
rect 2272 19170 2304 19202
rect 2344 19170 2376 19202
rect 2416 19170 2448 19202
rect 2488 19170 2520 19202
rect 2560 19170 2592 19202
rect 2632 19170 2664 19202
rect 2704 19170 2736 19202
rect 2776 19170 2808 19202
rect 2848 19170 2880 19202
rect 2920 19170 2952 19202
rect 2992 19170 3024 19202
rect 3064 19170 3096 19202
rect 3136 19170 3168 19202
rect 3208 19170 3240 19202
rect 3280 19170 3312 19202
rect 3352 19170 3384 19202
rect 3424 19170 3456 19202
rect 3496 19170 3528 19202
rect 3568 19170 3600 19202
rect 3640 19170 3672 19202
rect 3712 19170 3744 19202
rect 3784 19170 3816 19202
rect 3856 19170 3888 19202
rect 112 19098 144 19130
rect 184 19098 216 19130
rect 256 19098 288 19130
rect 328 19098 360 19130
rect 400 19098 432 19130
rect 472 19098 504 19130
rect 544 19098 576 19130
rect 616 19098 648 19130
rect 688 19098 720 19130
rect 760 19098 792 19130
rect 832 19098 864 19130
rect 904 19098 936 19130
rect 976 19098 1008 19130
rect 1048 19098 1080 19130
rect 1120 19098 1152 19130
rect 1192 19098 1224 19130
rect 1264 19098 1296 19130
rect 1336 19098 1368 19130
rect 1408 19098 1440 19130
rect 1480 19098 1512 19130
rect 1552 19098 1584 19130
rect 1624 19098 1656 19130
rect 1696 19098 1728 19130
rect 1768 19098 1800 19130
rect 1840 19098 1872 19130
rect 1912 19098 1944 19130
rect 1984 19098 2016 19130
rect 2056 19098 2088 19130
rect 2128 19098 2160 19130
rect 2200 19098 2232 19130
rect 2272 19098 2304 19130
rect 2344 19098 2376 19130
rect 2416 19098 2448 19130
rect 2488 19098 2520 19130
rect 2560 19098 2592 19130
rect 2632 19098 2664 19130
rect 2704 19098 2736 19130
rect 2776 19098 2808 19130
rect 2848 19098 2880 19130
rect 2920 19098 2952 19130
rect 2992 19098 3024 19130
rect 3064 19098 3096 19130
rect 3136 19098 3168 19130
rect 3208 19098 3240 19130
rect 3280 19098 3312 19130
rect 3352 19098 3384 19130
rect 3424 19098 3456 19130
rect 3496 19098 3528 19130
rect 3568 19098 3600 19130
rect 3640 19098 3672 19130
rect 3712 19098 3744 19130
rect 3784 19098 3816 19130
rect 3856 19098 3888 19130
rect 112 19026 144 19058
rect 184 19026 216 19058
rect 256 19026 288 19058
rect 328 19026 360 19058
rect 400 19026 432 19058
rect 472 19026 504 19058
rect 544 19026 576 19058
rect 616 19026 648 19058
rect 688 19026 720 19058
rect 760 19026 792 19058
rect 832 19026 864 19058
rect 904 19026 936 19058
rect 976 19026 1008 19058
rect 1048 19026 1080 19058
rect 1120 19026 1152 19058
rect 1192 19026 1224 19058
rect 1264 19026 1296 19058
rect 1336 19026 1368 19058
rect 1408 19026 1440 19058
rect 1480 19026 1512 19058
rect 1552 19026 1584 19058
rect 1624 19026 1656 19058
rect 1696 19026 1728 19058
rect 1768 19026 1800 19058
rect 1840 19026 1872 19058
rect 1912 19026 1944 19058
rect 1984 19026 2016 19058
rect 2056 19026 2088 19058
rect 2128 19026 2160 19058
rect 2200 19026 2232 19058
rect 2272 19026 2304 19058
rect 2344 19026 2376 19058
rect 2416 19026 2448 19058
rect 2488 19026 2520 19058
rect 2560 19026 2592 19058
rect 2632 19026 2664 19058
rect 2704 19026 2736 19058
rect 2776 19026 2808 19058
rect 2848 19026 2880 19058
rect 2920 19026 2952 19058
rect 2992 19026 3024 19058
rect 3064 19026 3096 19058
rect 3136 19026 3168 19058
rect 3208 19026 3240 19058
rect 3280 19026 3312 19058
rect 3352 19026 3384 19058
rect 3424 19026 3456 19058
rect 3496 19026 3528 19058
rect 3568 19026 3600 19058
rect 3640 19026 3672 19058
rect 3712 19026 3744 19058
rect 3784 19026 3816 19058
rect 3856 19026 3888 19058
rect 112 18954 144 18986
rect 184 18954 216 18986
rect 256 18954 288 18986
rect 328 18954 360 18986
rect 400 18954 432 18986
rect 472 18954 504 18986
rect 544 18954 576 18986
rect 616 18954 648 18986
rect 688 18954 720 18986
rect 760 18954 792 18986
rect 832 18954 864 18986
rect 904 18954 936 18986
rect 976 18954 1008 18986
rect 1048 18954 1080 18986
rect 1120 18954 1152 18986
rect 1192 18954 1224 18986
rect 1264 18954 1296 18986
rect 1336 18954 1368 18986
rect 1408 18954 1440 18986
rect 1480 18954 1512 18986
rect 1552 18954 1584 18986
rect 1624 18954 1656 18986
rect 1696 18954 1728 18986
rect 1768 18954 1800 18986
rect 1840 18954 1872 18986
rect 1912 18954 1944 18986
rect 1984 18954 2016 18986
rect 2056 18954 2088 18986
rect 2128 18954 2160 18986
rect 2200 18954 2232 18986
rect 2272 18954 2304 18986
rect 2344 18954 2376 18986
rect 2416 18954 2448 18986
rect 2488 18954 2520 18986
rect 2560 18954 2592 18986
rect 2632 18954 2664 18986
rect 2704 18954 2736 18986
rect 2776 18954 2808 18986
rect 2848 18954 2880 18986
rect 2920 18954 2952 18986
rect 2992 18954 3024 18986
rect 3064 18954 3096 18986
rect 3136 18954 3168 18986
rect 3208 18954 3240 18986
rect 3280 18954 3312 18986
rect 3352 18954 3384 18986
rect 3424 18954 3456 18986
rect 3496 18954 3528 18986
rect 3568 18954 3600 18986
rect 3640 18954 3672 18986
rect 3712 18954 3744 18986
rect 3784 18954 3816 18986
rect 3856 18954 3888 18986
rect 112 18882 144 18914
rect 184 18882 216 18914
rect 256 18882 288 18914
rect 328 18882 360 18914
rect 400 18882 432 18914
rect 472 18882 504 18914
rect 544 18882 576 18914
rect 616 18882 648 18914
rect 688 18882 720 18914
rect 760 18882 792 18914
rect 832 18882 864 18914
rect 904 18882 936 18914
rect 976 18882 1008 18914
rect 1048 18882 1080 18914
rect 1120 18882 1152 18914
rect 1192 18882 1224 18914
rect 1264 18882 1296 18914
rect 1336 18882 1368 18914
rect 1408 18882 1440 18914
rect 1480 18882 1512 18914
rect 1552 18882 1584 18914
rect 1624 18882 1656 18914
rect 1696 18882 1728 18914
rect 1768 18882 1800 18914
rect 1840 18882 1872 18914
rect 1912 18882 1944 18914
rect 1984 18882 2016 18914
rect 2056 18882 2088 18914
rect 2128 18882 2160 18914
rect 2200 18882 2232 18914
rect 2272 18882 2304 18914
rect 2344 18882 2376 18914
rect 2416 18882 2448 18914
rect 2488 18882 2520 18914
rect 2560 18882 2592 18914
rect 2632 18882 2664 18914
rect 2704 18882 2736 18914
rect 2776 18882 2808 18914
rect 2848 18882 2880 18914
rect 2920 18882 2952 18914
rect 2992 18882 3024 18914
rect 3064 18882 3096 18914
rect 3136 18882 3168 18914
rect 3208 18882 3240 18914
rect 3280 18882 3312 18914
rect 3352 18882 3384 18914
rect 3424 18882 3456 18914
rect 3496 18882 3528 18914
rect 3568 18882 3600 18914
rect 3640 18882 3672 18914
rect 3712 18882 3744 18914
rect 3784 18882 3816 18914
rect 3856 18882 3888 18914
rect 112 18810 144 18842
rect 184 18810 216 18842
rect 256 18810 288 18842
rect 328 18810 360 18842
rect 400 18810 432 18842
rect 472 18810 504 18842
rect 544 18810 576 18842
rect 616 18810 648 18842
rect 688 18810 720 18842
rect 760 18810 792 18842
rect 832 18810 864 18842
rect 904 18810 936 18842
rect 976 18810 1008 18842
rect 1048 18810 1080 18842
rect 1120 18810 1152 18842
rect 1192 18810 1224 18842
rect 1264 18810 1296 18842
rect 1336 18810 1368 18842
rect 1408 18810 1440 18842
rect 1480 18810 1512 18842
rect 1552 18810 1584 18842
rect 1624 18810 1656 18842
rect 1696 18810 1728 18842
rect 1768 18810 1800 18842
rect 1840 18810 1872 18842
rect 1912 18810 1944 18842
rect 1984 18810 2016 18842
rect 2056 18810 2088 18842
rect 2128 18810 2160 18842
rect 2200 18810 2232 18842
rect 2272 18810 2304 18842
rect 2344 18810 2376 18842
rect 2416 18810 2448 18842
rect 2488 18810 2520 18842
rect 2560 18810 2592 18842
rect 2632 18810 2664 18842
rect 2704 18810 2736 18842
rect 2776 18810 2808 18842
rect 2848 18810 2880 18842
rect 2920 18810 2952 18842
rect 2992 18810 3024 18842
rect 3064 18810 3096 18842
rect 3136 18810 3168 18842
rect 3208 18810 3240 18842
rect 3280 18810 3312 18842
rect 3352 18810 3384 18842
rect 3424 18810 3456 18842
rect 3496 18810 3528 18842
rect 3568 18810 3600 18842
rect 3640 18810 3672 18842
rect 3712 18810 3744 18842
rect 3784 18810 3816 18842
rect 3856 18810 3888 18842
rect 112 18738 144 18770
rect 184 18738 216 18770
rect 256 18738 288 18770
rect 328 18738 360 18770
rect 400 18738 432 18770
rect 472 18738 504 18770
rect 544 18738 576 18770
rect 616 18738 648 18770
rect 688 18738 720 18770
rect 760 18738 792 18770
rect 832 18738 864 18770
rect 904 18738 936 18770
rect 976 18738 1008 18770
rect 1048 18738 1080 18770
rect 1120 18738 1152 18770
rect 1192 18738 1224 18770
rect 1264 18738 1296 18770
rect 1336 18738 1368 18770
rect 1408 18738 1440 18770
rect 1480 18738 1512 18770
rect 1552 18738 1584 18770
rect 1624 18738 1656 18770
rect 1696 18738 1728 18770
rect 1768 18738 1800 18770
rect 1840 18738 1872 18770
rect 1912 18738 1944 18770
rect 1984 18738 2016 18770
rect 2056 18738 2088 18770
rect 2128 18738 2160 18770
rect 2200 18738 2232 18770
rect 2272 18738 2304 18770
rect 2344 18738 2376 18770
rect 2416 18738 2448 18770
rect 2488 18738 2520 18770
rect 2560 18738 2592 18770
rect 2632 18738 2664 18770
rect 2704 18738 2736 18770
rect 2776 18738 2808 18770
rect 2848 18738 2880 18770
rect 2920 18738 2952 18770
rect 2992 18738 3024 18770
rect 3064 18738 3096 18770
rect 3136 18738 3168 18770
rect 3208 18738 3240 18770
rect 3280 18738 3312 18770
rect 3352 18738 3384 18770
rect 3424 18738 3456 18770
rect 3496 18738 3528 18770
rect 3568 18738 3600 18770
rect 3640 18738 3672 18770
rect 3712 18738 3744 18770
rect 3784 18738 3816 18770
rect 3856 18738 3888 18770
rect 112 18666 144 18698
rect 184 18666 216 18698
rect 256 18666 288 18698
rect 328 18666 360 18698
rect 400 18666 432 18698
rect 472 18666 504 18698
rect 544 18666 576 18698
rect 616 18666 648 18698
rect 688 18666 720 18698
rect 760 18666 792 18698
rect 832 18666 864 18698
rect 904 18666 936 18698
rect 976 18666 1008 18698
rect 1048 18666 1080 18698
rect 1120 18666 1152 18698
rect 1192 18666 1224 18698
rect 1264 18666 1296 18698
rect 1336 18666 1368 18698
rect 1408 18666 1440 18698
rect 1480 18666 1512 18698
rect 1552 18666 1584 18698
rect 1624 18666 1656 18698
rect 1696 18666 1728 18698
rect 1768 18666 1800 18698
rect 1840 18666 1872 18698
rect 1912 18666 1944 18698
rect 1984 18666 2016 18698
rect 2056 18666 2088 18698
rect 2128 18666 2160 18698
rect 2200 18666 2232 18698
rect 2272 18666 2304 18698
rect 2344 18666 2376 18698
rect 2416 18666 2448 18698
rect 2488 18666 2520 18698
rect 2560 18666 2592 18698
rect 2632 18666 2664 18698
rect 2704 18666 2736 18698
rect 2776 18666 2808 18698
rect 2848 18666 2880 18698
rect 2920 18666 2952 18698
rect 2992 18666 3024 18698
rect 3064 18666 3096 18698
rect 3136 18666 3168 18698
rect 3208 18666 3240 18698
rect 3280 18666 3312 18698
rect 3352 18666 3384 18698
rect 3424 18666 3456 18698
rect 3496 18666 3528 18698
rect 3568 18666 3600 18698
rect 3640 18666 3672 18698
rect 3712 18666 3744 18698
rect 3784 18666 3816 18698
rect 3856 18666 3888 18698
rect 112 18594 144 18626
rect 184 18594 216 18626
rect 256 18594 288 18626
rect 328 18594 360 18626
rect 400 18594 432 18626
rect 472 18594 504 18626
rect 544 18594 576 18626
rect 616 18594 648 18626
rect 688 18594 720 18626
rect 760 18594 792 18626
rect 832 18594 864 18626
rect 904 18594 936 18626
rect 976 18594 1008 18626
rect 1048 18594 1080 18626
rect 1120 18594 1152 18626
rect 1192 18594 1224 18626
rect 1264 18594 1296 18626
rect 1336 18594 1368 18626
rect 1408 18594 1440 18626
rect 1480 18594 1512 18626
rect 1552 18594 1584 18626
rect 1624 18594 1656 18626
rect 1696 18594 1728 18626
rect 1768 18594 1800 18626
rect 1840 18594 1872 18626
rect 1912 18594 1944 18626
rect 1984 18594 2016 18626
rect 2056 18594 2088 18626
rect 2128 18594 2160 18626
rect 2200 18594 2232 18626
rect 2272 18594 2304 18626
rect 2344 18594 2376 18626
rect 2416 18594 2448 18626
rect 2488 18594 2520 18626
rect 2560 18594 2592 18626
rect 2632 18594 2664 18626
rect 2704 18594 2736 18626
rect 2776 18594 2808 18626
rect 2848 18594 2880 18626
rect 2920 18594 2952 18626
rect 2992 18594 3024 18626
rect 3064 18594 3096 18626
rect 3136 18594 3168 18626
rect 3208 18594 3240 18626
rect 3280 18594 3312 18626
rect 3352 18594 3384 18626
rect 3424 18594 3456 18626
rect 3496 18594 3528 18626
rect 3568 18594 3600 18626
rect 3640 18594 3672 18626
rect 3712 18594 3744 18626
rect 3784 18594 3816 18626
rect 3856 18594 3888 18626
rect 112 18522 144 18554
rect 184 18522 216 18554
rect 256 18522 288 18554
rect 328 18522 360 18554
rect 400 18522 432 18554
rect 472 18522 504 18554
rect 544 18522 576 18554
rect 616 18522 648 18554
rect 688 18522 720 18554
rect 760 18522 792 18554
rect 832 18522 864 18554
rect 904 18522 936 18554
rect 976 18522 1008 18554
rect 1048 18522 1080 18554
rect 1120 18522 1152 18554
rect 1192 18522 1224 18554
rect 1264 18522 1296 18554
rect 1336 18522 1368 18554
rect 1408 18522 1440 18554
rect 1480 18522 1512 18554
rect 1552 18522 1584 18554
rect 1624 18522 1656 18554
rect 1696 18522 1728 18554
rect 1768 18522 1800 18554
rect 1840 18522 1872 18554
rect 1912 18522 1944 18554
rect 1984 18522 2016 18554
rect 2056 18522 2088 18554
rect 2128 18522 2160 18554
rect 2200 18522 2232 18554
rect 2272 18522 2304 18554
rect 2344 18522 2376 18554
rect 2416 18522 2448 18554
rect 2488 18522 2520 18554
rect 2560 18522 2592 18554
rect 2632 18522 2664 18554
rect 2704 18522 2736 18554
rect 2776 18522 2808 18554
rect 2848 18522 2880 18554
rect 2920 18522 2952 18554
rect 2992 18522 3024 18554
rect 3064 18522 3096 18554
rect 3136 18522 3168 18554
rect 3208 18522 3240 18554
rect 3280 18522 3312 18554
rect 3352 18522 3384 18554
rect 3424 18522 3456 18554
rect 3496 18522 3528 18554
rect 3568 18522 3600 18554
rect 3640 18522 3672 18554
rect 3712 18522 3744 18554
rect 3784 18522 3816 18554
rect 3856 18522 3888 18554
rect 112 18450 144 18482
rect 184 18450 216 18482
rect 256 18450 288 18482
rect 328 18450 360 18482
rect 400 18450 432 18482
rect 472 18450 504 18482
rect 544 18450 576 18482
rect 616 18450 648 18482
rect 688 18450 720 18482
rect 760 18450 792 18482
rect 832 18450 864 18482
rect 904 18450 936 18482
rect 976 18450 1008 18482
rect 1048 18450 1080 18482
rect 1120 18450 1152 18482
rect 1192 18450 1224 18482
rect 1264 18450 1296 18482
rect 1336 18450 1368 18482
rect 1408 18450 1440 18482
rect 1480 18450 1512 18482
rect 1552 18450 1584 18482
rect 1624 18450 1656 18482
rect 1696 18450 1728 18482
rect 1768 18450 1800 18482
rect 1840 18450 1872 18482
rect 1912 18450 1944 18482
rect 1984 18450 2016 18482
rect 2056 18450 2088 18482
rect 2128 18450 2160 18482
rect 2200 18450 2232 18482
rect 2272 18450 2304 18482
rect 2344 18450 2376 18482
rect 2416 18450 2448 18482
rect 2488 18450 2520 18482
rect 2560 18450 2592 18482
rect 2632 18450 2664 18482
rect 2704 18450 2736 18482
rect 2776 18450 2808 18482
rect 2848 18450 2880 18482
rect 2920 18450 2952 18482
rect 2992 18450 3024 18482
rect 3064 18450 3096 18482
rect 3136 18450 3168 18482
rect 3208 18450 3240 18482
rect 3280 18450 3312 18482
rect 3352 18450 3384 18482
rect 3424 18450 3456 18482
rect 3496 18450 3528 18482
rect 3568 18450 3600 18482
rect 3640 18450 3672 18482
rect 3712 18450 3744 18482
rect 3784 18450 3816 18482
rect 3856 18450 3888 18482
rect 112 18378 144 18410
rect 184 18378 216 18410
rect 256 18378 288 18410
rect 328 18378 360 18410
rect 400 18378 432 18410
rect 472 18378 504 18410
rect 544 18378 576 18410
rect 616 18378 648 18410
rect 688 18378 720 18410
rect 760 18378 792 18410
rect 832 18378 864 18410
rect 904 18378 936 18410
rect 976 18378 1008 18410
rect 1048 18378 1080 18410
rect 1120 18378 1152 18410
rect 1192 18378 1224 18410
rect 1264 18378 1296 18410
rect 1336 18378 1368 18410
rect 1408 18378 1440 18410
rect 1480 18378 1512 18410
rect 1552 18378 1584 18410
rect 1624 18378 1656 18410
rect 1696 18378 1728 18410
rect 1768 18378 1800 18410
rect 1840 18378 1872 18410
rect 1912 18378 1944 18410
rect 1984 18378 2016 18410
rect 2056 18378 2088 18410
rect 2128 18378 2160 18410
rect 2200 18378 2232 18410
rect 2272 18378 2304 18410
rect 2344 18378 2376 18410
rect 2416 18378 2448 18410
rect 2488 18378 2520 18410
rect 2560 18378 2592 18410
rect 2632 18378 2664 18410
rect 2704 18378 2736 18410
rect 2776 18378 2808 18410
rect 2848 18378 2880 18410
rect 2920 18378 2952 18410
rect 2992 18378 3024 18410
rect 3064 18378 3096 18410
rect 3136 18378 3168 18410
rect 3208 18378 3240 18410
rect 3280 18378 3312 18410
rect 3352 18378 3384 18410
rect 3424 18378 3456 18410
rect 3496 18378 3528 18410
rect 3568 18378 3600 18410
rect 3640 18378 3672 18410
rect 3712 18378 3744 18410
rect 3784 18378 3816 18410
rect 3856 18378 3888 18410
rect 112 18306 144 18338
rect 184 18306 216 18338
rect 256 18306 288 18338
rect 328 18306 360 18338
rect 400 18306 432 18338
rect 472 18306 504 18338
rect 544 18306 576 18338
rect 616 18306 648 18338
rect 688 18306 720 18338
rect 760 18306 792 18338
rect 832 18306 864 18338
rect 904 18306 936 18338
rect 976 18306 1008 18338
rect 1048 18306 1080 18338
rect 1120 18306 1152 18338
rect 1192 18306 1224 18338
rect 1264 18306 1296 18338
rect 1336 18306 1368 18338
rect 1408 18306 1440 18338
rect 1480 18306 1512 18338
rect 1552 18306 1584 18338
rect 1624 18306 1656 18338
rect 1696 18306 1728 18338
rect 1768 18306 1800 18338
rect 1840 18306 1872 18338
rect 1912 18306 1944 18338
rect 1984 18306 2016 18338
rect 2056 18306 2088 18338
rect 2128 18306 2160 18338
rect 2200 18306 2232 18338
rect 2272 18306 2304 18338
rect 2344 18306 2376 18338
rect 2416 18306 2448 18338
rect 2488 18306 2520 18338
rect 2560 18306 2592 18338
rect 2632 18306 2664 18338
rect 2704 18306 2736 18338
rect 2776 18306 2808 18338
rect 2848 18306 2880 18338
rect 2920 18306 2952 18338
rect 2992 18306 3024 18338
rect 3064 18306 3096 18338
rect 3136 18306 3168 18338
rect 3208 18306 3240 18338
rect 3280 18306 3312 18338
rect 3352 18306 3384 18338
rect 3424 18306 3456 18338
rect 3496 18306 3528 18338
rect 3568 18306 3600 18338
rect 3640 18306 3672 18338
rect 3712 18306 3744 18338
rect 3784 18306 3816 18338
rect 3856 18306 3888 18338
rect 112 18234 144 18266
rect 184 18234 216 18266
rect 256 18234 288 18266
rect 328 18234 360 18266
rect 400 18234 432 18266
rect 472 18234 504 18266
rect 544 18234 576 18266
rect 616 18234 648 18266
rect 688 18234 720 18266
rect 760 18234 792 18266
rect 832 18234 864 18266
rect 904 18234 936 18266
rect 976 18234 1008 18266
rect 1048 18234 1080 18266
rect 1120 18234 1152 18266
rect 1192 18234 1224 18266
rect 1264 18234 1296 18266
rect 1336 18234 1368 18266
rect 1408 18234 1440 18266
rect 1480 18234 1512 18266
rect 1552 18234 1584 18266
rect 1624 18234 1656 18266
rect 1696 18234 1728 18266
rect 1768 18234 1800 18266
rect 1840 18234 1872 18266
rect 1912 18234 1944 18266
rect 1984 18234 2016 18266
rect 2056 18234 2088 18266
rect 2128 18234 2160 18266
rect 2200 18234 2232 18266
rect 2272 18234 2304 18266
rect 2344 18234 2376 18266
rect 2416 18234 2448 18266
rect 2488 18234 2520 18266
rect 2560 18234 2592 18266
rect 2632 18234 2664 18266
rect 2704 18234 2736 18266
rect 2776 18234 2808 18266
rect 2848 18234 2880 18266
rect 2920 18234 2952 18266
rect 2992 18234 3024 18266
rect 3064 18234 3096 18266
rect 3136 18234 3168 18266
rect 3208 18234 3240 18266
rect 3280 18234 3312 18266
rect 3352 18234 3384 18266
rect 3424 18234 3456 18266
rect 3496 18234 3528 18266
rect 3568 18234 3600 18266
rect 3640 18234 3672 18266
rect 3712 18234 3744 18266
rect 3784 18234 3816 18266
rect 3856 18234 3888 18266
rect 112 18162 144 18194
rect 184 18162 216 18194
rect 256 18162 288 18194
rect 328 18162 360 18194
rect 400 18162 432 18194
rect 472 18162 504 18194
rect 544 18162 576 18194
rect 616 18162 648 18194
rect 688 18162 720 18194
rect 760 18162 792 18194
rect 832 18162 864 18194
rect 904 18162 936 18194
rect 976 18162 1008 18194
rect 1048 18162 1080 18194
rect 1120 18162 1152 18194
rect 1192 18162 1224 18194
rect 1264 18162 1296 18194
rect 1336 18162 1368 18194
rect 1408 18162 1440 18194
rect 1480 18162 1512 18194
rect 1552 18162 1584 18194
rect 1624 18162 1656 18194
rect 1696 18162 1728 18194
rect 1768 18162 1800 18194
rect 1840 18162 1872 18194
rect 1912 18162 1944 18194
rect 1984 18162 2016 18194
rect 2056 18162 2088 18194
rect 2128 18162 2160 18194
rect 2200 18162 2232 18194
rect 2272 18162 2304 18194
rect 2344 18162 2376 18194
rect 2416 18162 2448 18194
rect 2488 18162 2520 18194
rect 2560 18162 2592 18194
rect 2632 18162 2664 18194
rect 2704 18162 2736 18194
rect 2776 18162 2808 18194
rect 2848 18162 2880 18194
rect 2920 18162 2952 18194
rect 2992 18162 3024 18194
rect 3064 18162 3096 18194
rect 3136 18162 3168 18194
rect 3208 18162 3240 18194
rect 3280 18162 3312 18194
rect 3352 18162 3384 18194
rect 3424 18162 3456 18194
rect 3496 18162 3528 18194
rect 3568 18162 3600 18194
rect 3640 18162 3672 18194
rect 3712 18162 3744 18194
rect 3784 18162 3816 18194
rect 3856 18162 3888 18194
rect 184 17816 216 17848
rect 256 17816 288 17848
rect 328 17816 360 17848
rect 400 17816 432 17848
rect 472 17816 504 17848
rect 544 17816 576 17848
rect 616 17816 648 17848
rect 688 17816 720 17848
rect 760 17816 792 17848
rect 832 17816 864 17848
rect 904 17816 936 17848
rect 976 17816 1008 17848
rect 1048 17816 1080 17848
rect 1120 17816 1152 17848
rect 1192 17816 1224 17848
rect 1264 17816 1296 17848
rect 1336 17816 1368 17848
rect 1408 17816 1440 17848
rect 1480 17816 1512 17848
rect 1552 17816 1584 17848
rect 1624 17816 1656 17848
rect 1696 17816 1728 17848
rect 1768 17816 1800 17848
rect 1840 17816 1872 17848
rect 1912 17816 1944 17848
rect 1984 17816 2016 17848
rect 2056 17816 2088 17848
rect 2128 17816 2160 17848
rect 2200 17816 2232 17848
rect 2272 17816 2304 17848
rect 2344 17816 2376 17848
rect 2416 17816 2448 17848
rect 2488 17816 2520 17848
rect 2560 17816 2592 17848
rect 2632 17816 2664 17848
rect 2704 17816 2736 17848
rect 2776 17816 2808 17848
rect 2848 17816 2880 17848
rect 2920 17816 2952 17848
rect 2992 17816 3024 17848
rect 3064 17816 3096 17848
rect 3136 17816 3168 17848
rect 3208 17816 3240 17848
rect 3280 17816 3312 17848
rect 3352 17816 3384 17848
rect 3424 17816 3456 17848
rect 3496 17816 3528 17848
rect 3568 17816 3600 17848
rect 3640 17816 3672 17848
rect 3712 17816 3744 17848
rect 3784 17816 3816 17848
rect 3856 17816 3888 17848
rect 112 17744 144 17776
rect 184 17744 216 17776
rect 256 17744 288 17776
rect 328 17744 360 17776
rect 400 17744 432 17776
rect 472 17744 504 17776
rect 544 17744 576 17776
rect 616 17744 648 17776
rect 688 17744 720 17776
rect 760 17744 792 17776
rect 832 17744 864 17776
rect 904 17744 936 17776
rect 976 17744 1008 17776
rect 1048 17744 1080 17776
rect 1120 17744 1152 17776
rect 1192 17744 1224 17776
rect 1264 17744 1296 17776
rect 1336 17744 1368 17776
rect 1408 17744 1440 17776
rect 1480 17744 1512 17776
rect 1552 17744 1584 17776
rect 1624 17744 1656 17776
rect 1696 17744 1728 17776
rect 1768 17744 1800 17776
rect 1840 17744 1872 17776
rect 1912 17744 1944 17776
rect 1984 17744 2016 17776
rect 2056 17744 2088 17776
rect 2128 17744 2160 17776
rect 2200 17744 2232 17776
rect 2272 17744 2304 17776
rect 2344 17744 2376 17776
rect 2416 17744 2448 17776
rect 2488 17744 2520 17776
rect 2560 17744 2592 17776
rect 2632 17744 2664 17776
rect 2704 17744 2736 17776
rect 2776 17744 2808 17776
rect 2848 17744 2880 17776
rect 2920 17744 2952 17776
rect 2992 17744 3024 17776
rect 3064 17744 3096 17776
rect 3136 17744 3168 17776
rect 3208 17744 3240 17776
rect 3280 17744 3312 17776
rect 3352 17744 3384 17776
rect 3424 17744 3456 17776
rect 3496 17744 3528 17776
rect 3568 17744 3600 17776
rect 3640 17744 3672 17776
rect 3712 17744 3744 17776
rect 3784 17744 3816 17776
rect 3856 17744 3888 17776
rect 112 17672 144 17704
rect 184 17672 216 17704
rect 256 17672 288 17704
rect 328 17672 360 17704
rect 400 17672 432 17704
rect 472 17672 504 17704
rect 544 17672 576 17704
rect 616 17672 648 17704
rect 688 17672 720 17704
rect 760 17672 792 17704
rect 832 17672 864 17704
rect 904 17672 936 17704
rect 976 17672 1008 17704
rect 1048 17672 1080 17704
rect 1120 17672 1152 17704
rect 1192 17672 1224 17704
rect 1264 17672 1296 17704
rect 1336 17672 1368 17704
rect 1408 17672 1440 17704
rect 1480 17672 1512 17704
rect 1552 17672 1584 17704
rect 1624 17672 1656 17704
rect 1696 17672 1728 17704
rect 1768 17672 1800 17704
rect 1840 17672 1872 17704
rect 1912 17672 1944 17704
rect 1984 17672 2016 17704
rect 2056 17672 2088 17704
rect 2128 17672 2160 17704
rect 2200 17672 2232 17704
rect 2272 17672 2304 17704
rect 2344 17672 2376 17704
rect 2416 17672 2448 17704
rect 2488 17672 2520 17704
rect 2560 17672 2592 17704
rect 2632 17672 2664 17704
rect 2704 17672 2736 17704
rect 2776 17672 2808 17704
rect 2848 17672 2880 17704
rect 2920 17672 2952 17704
rect 2992 17672 3024 17704
rect 3064 17672 3096 17704
rect 3136 17672 3168 17704
rect 3208 17672 3240 17704
rect 3280 17672 3312 17704
rect 3352 17672 3384 17704
rect 3424 17672 3456 17704
rect 3496 17672 3528 17704
rect 3568 17672 3600 17704
rect 3640 17672 3672 17704
rect 3712 17672 3744 17704
rect 3784 17672 3816 17704
rect 3856 17672 3888 17704
rect 112 17600 144 17632
rect 184 17600 216 17632
rect 256 17600 288 17632
rect 328 17600 360 17632
rect 400 17600 432 17632
rect 472 17600 504 17632
rect 544 17600 576 17632
rect 616 17600 648 17632
rect 688 17600 720 17632
rect 760 17600 792 17632
rect 832 17600 864 17632
rect 904 17600 936 17632
rect 976 17600 1008 17632
rect 1048 17600 1080 17632
rect 1120 17600 1152 17632
rect 1192 17600 1224 17632
rect 1264 17600 1296 17632
rect 1336 17600 1368 17632
rect 1408 17600 1440 17632
rect 1480 17600 1512 17632
rect 1552 17600 1584 17632
rect 1624 17600 1656 17632
rect 1696 17600 1728 17632
rect 1768 17600 1800 17632
rect 1840 17600 1872 17632
rect 1912 17600 1944 17632
rect 1984 17600 2016 17632
rect 2056 17600 2088 17632
rect 2128 17600 2160 17632
rect 2200 17600 2232 17632
rect 2272 17600 2304 17632
rect 2344 17600 2376 17632
rect 2416 17600 2448 17632
rect 2488 17600 2520 17632
rect 2560 17600 2592 17632
rect 2632 17600 2664 17632
rect 2704 17600 2736 17632
rect 2776 17600 2808 17632
rect 2848 17600 2880 17632
rect 2920 17600 2952 17632
rect 2992 17600 3024 17632
rect 3064 17600 3096 17632
rect 3136 17600 3168 17632
rect 3208 17600 3240 17632
rect 3280 17600 3312 17632
rect 3352 17600 3384 17632
rect 3424 17600 3456 17632
rect 3496 17600 3528 17632
rect 3568 17600 3600 17632
rect 3640 17600 3672 17632
rect 3712 17600 3744 17632
rect 3784 17600 3816 17632
rect 3856 17600 3888 17632
rect 112 17528 144 17560
rect 184 17528 216 17560
rect 256 17528 288 17560
rect 328 17528 360 17560
rect 400 17528 432 17560
rect 472 17528 504 17560
rect 544 17528 576 17560
rect 616 17528 648 17560
rect 688 17528 720 17560
rect 760 17528 792 17560
rect 832 17528 864 17560
rect 904 17528 936 17560
rect 976 17528 1008 17560
rect 1048 17528 1080 17560
rect 1120 17528 1152 17560
rect 1192 17528 1224 17560
rect 1264 17528 1296 17560
rect 1336 17528 1368 17560
rect 1408 17528 1440 17560
rect 1480 17528 1512 17560
rect 1552 17528 1584 17560
rect 1624 17528 1656 17560
rect 1696 17528 1728 17560
rect 1768 17528 1800 17560
rect 1840 17528 1872 17560
rect 1912 17528 1944 17560
rect 1984 17528 2016 17560
rect 2056 17528 2088 17560
rect 2128 17528 2160 17560
rect 2200 17528 2232 17560
rect 2272 17528 2304 17560
rect 2344 17528 2376 17560
rect 2416 17528 2448 17560
rect 2488 17528 2520 17560
rect 2560 17528 2592 17560
rect 2632 17528 2664 17560
rect 2704 17528 2736 17560
rect 2776 17528 2808 17560
rect 2848 17528 2880 17560
rect 2920 17528 2952 17560
rect 2992 17528 3024 17560
rect 3064 17528 3096 17560
rect 3136 17528 3168 17560
rect 3208 17528 3240 17560
rect 3280 17528 3312 17560
rect 3352 17528 3384 17560
rect 3424 17528 3456 17560
rect 3496 17528 3528 17560
rect 3568 17528 3600 17560
rect 3640 17528 3672 17560
rect 3712 17528 3744 17560
rect 3784 17528 3816 17560
rect 3856 17528 3888 17560
rect 112 17456 144 17488
rect 184 17456 216 17488
rect 256 17456 288 17488
rect 328 17456 360 17488
rect 400 17456 432 17488
rect 472 17456 504 17488
rect 544 17456 576 17488
rect 616 17456 648 17488
rect 688 17456 720 17488
rect 760 17456 792 17488
rect 832 17456 864 17488
rect 904 17456 936 17488
rect 976 17456 1008 17488
rect 1048 17456 1080 17488
rect 1120 17456 1152 17488
rect 1192 17456 1224 17488
rect 1264 17456 1296 17488
rect 1336 17456 1368 17488
rect 1408 17456 1440 17488
rect 1480 17456 1512 17488
rect 1552 17456 1584 17488
rect 1624 17456 1656 17488
rect 1696 17456 1728 17488
rect 1768 17456 1800 17488
rect 1840 17456 1872 17488
rect 1912 17456 1944 17488
rect 1984 17456 2016 17488
rect 2056 17456 2088 17488
rect 2128 17456 2160 17488
rect 2200 17456 2232 17488
rect 2272 17456 2304 17488
rect 2344 17456 2376 17488
rect 2416 17456 2448 17488
rect 2488 17456 2520 17488
rect 2560 17456 2592 17488
rect 2632 17456 2664 17488
rect 2704 17456 2736 17488
rect 2776 17456 2808 17488
rect 2848 17456 2880 17488
rect 2920 17456 2952 17488
rect 2992 17456 3024 17488
rect 3064 17456 3096 17488
rect 3136 17456 3168 17488
rect 3208 17456 3240 17488
rect 3280 17456 3312 17488
rect 3352 17456 3384 17488
rect 3424 17456 3456 17488
rect 3496 17456 3528 17488
rect 3568 17456 3600 17488
rect 3640 17456 3672 17488
rect 3712 17456 3744 17488
rect 3784 17456 3816 17488
rect 3856 17456 3888 17488
rect 112 17384 144 17416
rect 184 17384 216 17416
rect 256 17384 288 17416
rect 328 17384 360 17416
rect 400 17384 432 17416
rect 472 17384 504 17416
rect 544 17384 576 17416
rect 616 17384 648 17416
rect 688 17384 720 17416
rect 760 17384 792 17416
rect 832 17384 864 17416
rect 904 17384 936 17416
rect 976 17384 1008 17416
rect 1048 17384 1080 17416
rect 1120 17384 1152 17416
rect 1192 17384 1224 17416
rect 1264 17384 1296 17416
rect 1336 17384 1368 17416
rect 1408 17384 1440 17416
rect 1480 17384 1512 17416
rect 1552 17384 1584 17416
rect 1624 17384 1656 17416
rect 1696 17384 1728 17416
rect 1768 17384 1800 17416
rect 1840 17384 1872 17416
rect 1912 17384 1944 17416
rect 1984 17384 2016 17416
rect 2056 17384 2088 17416
rect 2128 17384 2160 17416
rect 2200 17384 2232 17416
rect 2272 17384 2304 17416
rect 2344 17384 2376 17416
rect 2416 17384 2448 17416
rect 2488 17384 2520 17416
rect 2560 17384 2592 17416
rect 2632 17384 2664 17416
rect 2704 17384 2736 17416
rect 2776 17384 2808 17416
rect 2848 17384 2880 17416
rect 2920 17384 2952 17416
rect 2992 17384 3024 17416
rect 3064 17384 3096 17416
rect 3136 17384 3168 17416
rect 3208 17384 3240 17416
rect 3280 17384 3312 17416
rect 3352 17384 3384 17416
rect 3424 17384 3456 17416
rect 3496 17384 3528 17416
rect 3568 17384 3600 17416
rect 3640 17384 3672 17416
rect 3712 17384 3744 17416
rect 3784 17384 3816 17416
rect 3856 17384 3888 17416
rect 112 17312 144 17344
rect 184 17312 216 17344
rect 256 17312 288 17344
rect 328 17312 360 17344
rect 400 17312 432 17344
rect 472 17312 504 17344
rect 544 17312 576 17344
rect 616 17312 648 17344
rect 688 17312 720 17344
rect 760 17312 792 17344
rect 832 17312 864 17344
rect 904 17312 936 17344
rect 976 17312 1008 17344
rect 1048 17312 1080 17344
rect 1120 17312 1152 17344
rect 1192 17312 1224 17344
rect 1264 17312 1296 17344
rect 1336 17312 1368 17344
rect 1408 17312 1440 17344
rect 1480 17312 1512 17344
rect 1552 17312 1584 17344
rect 1624 17312 1656 17344
rect 1696 17312 1728 17344
rect 1768 17312 1800 17344
rect 1840 17312 1872 17344
rect 1912 17312 1944 17344
rect 1984 17312 2016 17344
rect 2056 17312 2088 17344
rect 2128 17312 2160 17344
rect 2200 17312 2232 17344
rect 2272 17312 2304 17344
rect 2344 17312 2376 17344
rect 2416 17312 2448 17344
rect 2488 17312 2520 17344
rect 2560 17312 2592 17344
rect 2632 17312 2664 17344
rect 2704 17312 2736 17344
rect 2776 17312 2808 17344
rect 2848 17312 2880 17344
rect 2920 17312 2952 17344
rect 2992 17312 3024 17344
rect 3064 17312 3096 17344
rect 3136 17312 3168 17344
rect 3208 17312 3240 17344
rect 3280 17312 3312 17344
rect 3352 17312 3384 17344
rect 3424 17312 3456 17344
rect 3496 17312 3528 17344
rect 3568 17312 3600 17344
rect 3640 17312 3672 17344
rect 3712 17312 3744 17344
rect 3784 17312 3816 17344
rect 3856 17312 3888 17344
rect 112 17240 144 17272
rect 184 17240 216 17272
rect 256 17240 288 17272
rect 328 17240 360 17272
rect 400 17240 432 17272
rect 472 17240 504 17272
rect 544 17240 576 17272
rect 616 17240 648 17272
rect 688 17240 720 17272
rect 760 17240 792 17272
rect 832 17240 864 17272
rect 904 17240 936 17272
rect 976 17240 1008 17272
rect 1048 17240 1080 17272
rect 1120 17240 1152 17272
rect 1192 17240 1224 17272
rect 1264 17240 1296 17272
rect 1336 17240 1368 17272
rect 1408 17240 1440 17272
rect 1480 17240 1512 17272
rect 1552 17240 1584 17272
rect 1624 17240 1656 17272
rect 1696 17240 1728 17272
rect 1768 17240 1800 17272
rect 1840 17240 1872 17272
rect 1912 17240 1944 17272
rect 1984 17240 2016 17272
rect 2056 17240 2088 17272
rect 2128 17240 2160 17272
rect 2200 17240 2232 17272
rect 2272 17240 2304 17272
rect 2344 17240 2376 17272
rect 2416 17240 2448 17272
rect 2488 17240 2520 17272
rect 2560 17240 2592 17272
rect 2632 17240 2664 17272
rect 2704 17240 2736 17272
rect 2776 17240 2808 17272
rect 2848 17240 2880 17272
rect 2920 17240 2952 17272
rect 2992 17240 3024 17272
rect 3064 17240 3096 17272
rect 3136 17240 3168 17272
rect 3208 17240 3240 17272
rect 3280 17240 3312 17272
rect 3352 17240 3384 17272
rect 3424 17240 3456 17272
rect 3496 17240 3528 17272
rect 3568 17240 3600 17272
rect 3640 17240 3672 17272
rect 3712 17240 3744 17272
rect 3784 17240 3816 17272
rect 3856 17240 3888 17272
rect 112 17168 144 17200
rect 184 17168 216 17200
rect 256 17168 288 17200
rect 328 17168 360 17200
rect 400 17168 432 17200
rect 472 17168 504 17200
rect 544 17168 576 17200
rect 616 17168 648 17200
rect 688 17168 720 17200
rect 760 17168 792 17200
rect 832 17168 864 17200
rect 904 17168 936 17200
rect 976 17168 1008 17200
rect 1048 17168 1080 17200
rect 1120 17168 1152 17200
rect 1192 17168 1224 17200
rect 1264 17168 1296 17200
rect 1336 17168 1368 17200
rect 1408 17168 1440 17200
rect 1480 17168 1512 17200
rect 1552 17168 1584 17200
rect 1624 17168 1656 17200
rect 1696 17168 1728 17200
rect 1768 17168 1800 17200
rect 1840 17168 1872 17200
rect 1912 17168 1944 17200
rect 1984 17168 2016 17200
rect 2056 17168 2088 17200
rect 2128 17168 2160 17200
rect 2200 17168 2232 17200
rect 2272 17168 2304 17200
rect 2344 17168 2376 17200
rect 2416 17168 2448 17200
rect 2488 17168 2520 17200
rect 2560 17168 2592 17200
rect 2632 17168 2664 17200
rect 2704 17168 2736 17200
rect 2776 17168 2808 17200
rect 2848 17168 2880 17200
rect 2920 17168 2952 17200
rect 2992 17168 3024 17200
rect 3064 17168 3096 17200
rect 3136 17168 3168 17200
rect 3208 17168 3240 17200
rect 3280 17168 3312 17200
rect 3352 17168 3384 17200
rect 3424 17168 3456 17200
rect 3496 17168 3528 17200
rect 3568 17168 3600 17200
rect 3640 17168 3672 17200
rect 3712 17168 3744 17200
rect 3784 17168 3816 17200
rect 3856 17168 3888 17200
rect 112 17096 144 17128
rect 184 17096 216 17128
rect 256 17096 288 17128
rect 328 17096 360 17128
rect 400 17096 432 17128
rect 472 17096 504 17128
rect 544 17096 576 17128
rect 616 17096 648 17128
rect 688 17096 720 17128
rect 760 17096 792 17128
rect 832 17096 864 17128
rect 904 17096 936 17128
rect 976 17096 1008 17128
rect 1048 17096 1080 17128
rect 1120 17096 1152 17128
rect 1192 17096 1224 17128
rect 1264 17096 1296 17128
rect 1336 17096 1368 17128
rect 1408 17096 1440 17128
rect 1480 17096 1512 17128
rect 1552 17096 1584 17128
rect 1624 17096 1656 17128
rect 1696 17096 1728 17128
rect 1768 17096 1800 17128
rect 1840 17096 1872 17128
rect 1912 17096 1944 17128
rect 1984 17096 2016 17128
rect 2056 17096 2088 17128
rect 2128 17096 2160 17128
rect 2200 17096 2232 17128
rect 2272 17096 2304 17128
rect 2344 17096 2376 17128
rect 2416 17096 2448 17128
rect 2488 17096 2520 17128
rect 2560 17096 2592 17128
rect 2632 17096 2664 17128
rect 2704 17096 2736 17128
rect 2776 17096 2808 17128
rect 2848 17096 2880 17128
rect 2920 17096 2952 17128
rect 2992 17096 3024 17128
rect 3064 17096 3096 17128
rect 3136 17096 3168 17128
rect 3208 17096 3240 17128
rect 3280 17096 3312 17128
rect 3352 17096 3384 17128
rect 3424 17096 3456 17128
rect 3496 17096 3528 17128
rect 3568 17096 3600 17128
rect 3640 17096 3672 17128
rect 3712 17096 3744 17128
rect 3784 17096 3816 17128
rect 3856 17096 3888 17128
rect 112 17024 144 17056
rect 184 17024 216 17056
rect 256 17024 288 17056
rect 328 17024 360 17056
rect 400 17024 432 17056
rect 472 17024 504 17056
rect 544 17024 576 17056
rect 616 17024 648 17056
rect 688 17024 720 17056
rect 760 17024 792 17056
rect 832 17024 864 17056
rect 904 17024 936 17056
rect 976 17024 1008 17056
rect 1048 17024 1080 17056
rect 1120 17024 1152 17056
rect 1192 17024 1224 17056
rect 1264 17024 1296 17056
rect 1336 17024 1368 17056
rect 1408 17024 1440 17056
rect 1480 17024 1512 17056
rect 1552 17024 1584 17056
rect 1624 17024 1656 17056
rect 1696 17024 1728 17056
rect 1768 17024 1800 17056
rect 1840 17024 1872 17056
rect 1912 17024 1944 17056
rect 1984 17024 2016 17056
rect 2056 17024 2088 17056
rect 2128 17024 2160 17056
rect 2200 17024 2232 17056
rect 2272 17024 2304 17056
rect 2344 17024 2376 17056
rect 2416 17024 2448 17056
rect 2488 17024 2520 17056
rect 2560 17024 2592 17056
rect 2632 17024 2664 17056
rect 2704 17024 2736 17056
rect 2776 17024 2808 17056
rect 2848 17024 2880 17056
rect 2920 17024 2952 17056
rect 2992 17024 3024 17056
rect 3064 17024 3096 17056
rect 3136 17024 3168 17056
rect 3208 17024 3240 17056
rect 3280 17024 3312 17056
rect 3352 17024 3384 17056
rect 3424 17024 3456 17056
rect 3496 17024 3528 17056
rect 3568 17024 3600 17056
rect 3640 17024 3672 17056
rect 3712 17024 3744 17056
rect 3784 17024 3816 17056
rect 3856 17024 3888 17056
rect 112 16952 144 16984
rect 184 16952 216 16984
rect 256 16952 288 16984
rect 328 16952 360 16984
rect 400 16952 432 16984
rect 472 16952 504 16984
rect 544 16952 576 16984
rect 616 16952 648 16984
rect 688 16952 720 16984
rect 760 16952 792 16984
rect 832 16952 864 16984
rect 904 16952 936 16984
rect 976 16952 1008 16984
rect 1048 16952 1080 16984
rect 1120 16952 1152 16984
rect 1192 16952 1224 16984
rect 1264 16952 1296 16984
rect 1336 16952 1368 16984
rect 1408 16952 1440 16984
rect 1480 16952 1512 16984
rect 1552 16952 1584 16984
rect 1624 16952 1656 16984
rect 1696 16952 1728 16984
rect 1768 16952 1800 16984
rect 1840 16952 1872 16984
rect 1912 16952 1944 16984
rect 1984 16952 2016 16984
rect 2056 16952 2088 16984
rect 2128 16952 2160 16984
rect 2200 16952 2232 16984
rect 2272 16952 2304 16984
rect 2344 16952 2376 16984
rect 2416 16952 2448 16984
rect 2488 16952 2520 16984
rect 2560 16952 2592 16984
rect 2632 16952 2664 16984
rect 2704 16952 2736 16984
rect 2776 16952 2808 16984
rect 2848 16952 2880 16984
rect 2920 16952 2952 16984
rect 2992 16952 3024 16984
rect 3064 16952 3096 16984
rect 3136 16952 3168 16984
rect 3208 16952 3240 16984
rect 3280 16952 3312 16984
rect 3352 16952 3384 16984
rect 3424 16952 3456 16984
rect 3496 16952 3528 16984
rect 3568 16952 3600 16984
rect 3640 16952 3672 16984
rect 3712 16952 3744 16984
rect 3784 16952 3816 16984
rect 3856 16952 3888 16984
rect 112 16880 144 16912
rect 184 16880 216 16912
rect 256 16880 288 16912
rect 328 16880 360 16912
rect 400 16880 432 16912
rect 472 16880 504 16912
rect 544 16880 576 16912
rect 616 16880 648 16912
rect 688 16880 720 16912
rect 760 16880 792 16912
rect 832 16880 864 16912
rect 904 16880 936 16912
rect 976 16880 1008 16912
rect 1048 16880 1080 16912
rect 1120 16880 1152 16912
rect 1192 16880 1224 16912
rect 1264 16880 1296 16912
rect 1336 16880 1368 16912
rect 1408 16880 1440 16912
rect 1480 16880 1512 16912
rect 1552 16880 1584 16912
rect 1624 16880 1656 16912
rect 1696 16880 1728 16912
rect 1768 16880 1800 16912
rect 1840 16880 1872 16912
rect 1912 16880 1944 16912
rect 1984 16880 2016 16912
rect 2056 16880 2088 16912
rect 2128 16880 2160 16912
rect 2200 16880 2232 16912
rect 2272 16880 2304 16912
rect 2344 16880 2376 16912
rect 2416 16880 2448 16912
rect 2488 16880 2520 16912
rect 2560 16880 2592 16912
rect 2632 16880 2664 16912
rect 2704 16880 2736 16912
rect 2776 16880 2808 16912
rect 2848 16880 2880 16912
rect 2920 16880 2952 16912
rect 2992 16880 3024 16912
rect 3064 16880 3096 16912
rect 3136 16880 3168 16912
rect 3208 16880 3240 16912
rect 3280 16880 3312 16912
rect 3352 16880 3384 16912
rect 3424 16880 3456 16912
rect 3496 16880 3528 16912
rect 3568 16880 3600 16912
rect 3640 16880 3672 16912
rect 3712 16880 3744 16912
rect 3784 16880 3816 16912
rect 3856 16880 3888 16912
rect 112 16808 144 16840
rect 184 16808 216 16840
rect 256 16808 288 16840
rect 328 16808 360 16840
rect 400 16808 432 16840
rect 472 16808 504 16840
rect 544 16808 576 16840
rect 616 16808 648 16840
rect 688 16808 720 16840
rect 760 16808 792 16840
rect 832 16808 864 16840
rect 904 16808 936 16840
rect 976 16808 1008 16840
rect 1048 16808 1080 16840
rect 1120 16808 1152 16840
rect 1192 16808 1224 16840
rect 1264 16808 1296 16840
rect 1336 16808 1368 16840
rect 1408 16808 1440 16840
rect 1480 16808 1512 16840
rect 1552 16808 1584 16840
rect 1624 16808 1656 16840
rect 1696 16808 1728 16840
rect 1768 16808 1800 16840
rect 1840 16808 1872 16840
rect 1912 16808 1944 16840
rect 1984 16808 2016 16840
rect 2056 16808 2088 16840
rect 2128 16808 2160 16840
rect 2200 16808 2232 16840
rect 2272 16808 2304 16840
rect 2344 16808 2376 16840
rect 2416 16808 2448 16840
rect 2488 16808 2520 16840
rect 2560 16808 2592 16840
rect 2632 16808 2664 16840
rect 2704 16808 2736 16840
rect 2776 16808 2808 16840
rect 2848 16808 2880 16840
rect 2920 16808 2952 16840
rect 2992 16808 3024 16840
rect 3064 16808 3096 16840
rect 3136 16808 3168 16840
rect 3208 16808 3240 16840
rect 3280 16808 3312 16840
rect 3352 16808 3384 16840
rect 3424 16808 3456 16840
rect 3496 16808 3528 16840
rect 3568 16808 3600 16840
rect 3640 16808 3672 16840
rect 3712 16808 3744 16840
rect 3784 16808 3816 16840
rect 3856 16808 3888 16840
rect 112 16736 144 16768
rect 184 16736 216 16768
rect 256 16736 288 16768
rect 328 16736 360 16768
rect 400 16736 432 16768
rect 472 16736 504 16768
rect 544 16736 576 16768
rect 616 16736 648 16768
rect 688 16736 720 16768
rect 760 16736 792 16768
rect 832 16736 864 16768
rect 904 16736 936 16768
rect 976 16736 1008 16768
rect 1048 16736 1080 16768
rect 1120 16736 1152 16768
rect 1192 16736 1224 16768
rect 1264 16736 1296 16768
rect 1336 16736 1368 16768
rect 1408 16736 1440 16768
rect 1480 16736 1512 16768
rect 1552 16736 1584 16768
rect 1624 16736 1656 16768
rect 1696 16736 1728 16768
rect 1768 16736 1800 16768
rect 1840 16736 1872 16768
rect 1912 16736 1944 16768
rect 1984 16736 2016 16768
rect 2056 16736 2088 16768
rect 2128 16736 2160 16768
rect 2200 16736 2232 16768
rect 2272 16736 2304 16768
rect 2344 16736 2376 16768
rect 2416 16736 2448 16768
rect 2488 16736 2520 16768
rect 2560 16736 2592 16768
rect 2632 16736 2664 16768
rect 2704 16736 2736 16768
rect 2776 16736 2808 16768
rect 2848 16736 2880 16768
rect 2920 16736 2952 16768
rect 2992 16736 3024 16768
rect 3064 16736 3096 16768
rect 3136 16736 3168 16768
rect 3208 16736 3240 16768
rect 3280 16736 3312 16768
rect 3352 16736 3384 16768
rect 3424 16736 3456 16768
rect 3496 16736 3528 16768
rect 3568 16736 3600 16768
rect 3640 16736 3672 16768
rect 3712 16736 3744 16768
rect 3784 16736 3816 16768
rect 3856 16736 3888 16768
rect 112 16664 144 16696
rect 184 16664 216 16696
rect 256 16664 288 16696
rect 328 16664 360 16696
rect 400 16664 432 16696
rect 472 16664 504 16696
rect 544 16664 576 16696
rect 616 16664 648 16696
rect 688 16664 720 16696
rect 760 16664 792 16696
rect 832 16664 864 16696
rect 904 16664 936 16696
rect 976 16664 1008 16696
rect 1048 16664 1080 16696
rect 1120 16664 1152 16696
rect 1192 16664 1224 16696
rect 1264 16664 1296 16696
rect 1336 16664 1368 16696
rect 1408 16664 1440 16696
rect 1480 16664 1512 16696
rect 1552 16664 1584 16696
rect 1624 16664 1656 16696
rect 1696 16664 1728 16696
rect 1768 16664 1800 16696
rect 1840 16664 1872 16696
rect 1912 16664 1944 16696
rect 1984 16664 2016 16696
rect 2056 16664 2088 16696
rect 2128 16664 2160 16696
rect 2200 16664 2232 16696
rect 2272 16664 2304 16696
rect 2344 16664 2376 16696
rect 2416 16664 2448 16696
rect 2488 16664 2520 16696
rect 2560 16664 2592 16696
rect 2632 16664 2664 16696
rect 2704 16664 2736 16696
rect 2776 16664 2808 16696
rect 2848 16664 2880 16696
rect 2920 16664 2952 16696
rect 2992 16664 3024 16696
rect 3064 16664 3096 16696
rect 3136 16664 3168 16696
rect 3208 16664 3240 16696
rect 3280 16664 3312 16696
rect 3352 16664 3384 16696
rect 3424 16664 3456 16696
rect 3496 16664 3528 16696
rect 3568 16664 3600 16696
rect 3640 16664 3672 16696
rect 3712 16664 3744 16696
rect 3784 16664 3816 16696
rect 3856 16664 3888 16696
rect 112 16592 144 16624
rect 184 16592 216 16624
rect 256 16592 288 16624
rect 328 16592 360 16624
rect 400 16592 432 16624
rect 472 16592 504 16624
rect 544 16592 576 16624
rect 616 16592 648 16624
rect 688 16592 720 16624
rect 760 16592 792 16624
rect 832 16592 864 16624
rect 904 16592 936 16624
rect 976 16592 1008 16624
rect 1048 16592 1080 16624
rect 1120 16592 1152 16624
rect 1192 16592 1224 16624
rect 1264 16592 1296 16624
rect 1336 16592 1368 16624
rect 1408 16592 1440 16624
rect 1480 16592 1512 16624
rect 1552 16592 1584 16624
rect 1624 16592 1656 16624
rect 1696 16592 1728 16624
rect 1768 16592 1800 16624
rect 1840 16592 1872 16624
rect 1912 16592 1944 16624
rect 1984 16592 2016 16624
rect 2056 16592 2088 16624
rect 2128 16592 2160 16624
rect 2200 16592 2232 16624
rect 2272 16592 2304 16624
rect 2344 16592 2376 16624
rect 2416 16592 2448 16624
rect 2488 16592 2520 16624
rect 2560 16592 2592 16624
rect 2632 16592 2664 16624
rect 2704 16592 2736 16624
rect 2776 16592 2808 16624
rect 2848 16592 2880 16624
rect 2920 16592 2952 16624
rect 2992 16592 3024 16624
rect 3064 16592 3096 16624
rect 3136 16592 3168 16624
rect 3208 16592 3240 16624
rect 3280 16592 3312 16624
rect 3352 16592 3384 16624
rect 3424 16592 3456 16624
rect 3496 16592 3528 16624
rect 3568 16592 3600 16624
rect 3640 16592 3672 16624
rect 3712 16592 3744 16624
rect 3784 16592 3816 16624
rect 3856 16592 3888 16624
rect 112 16520 144 16552
rect 184 16520 216 16552
rect 256 16520 288 16552
rect 328 16520 360 16552
rect 400 16520 432 16552
rect 472 16520 504 16552
rect 544 16520 576 16552
rect 616 16520 648 16552
rect 688 16520 720 16552
rect 760 16520 792 16552
rect 832 16520 864 16552
rect 904 16520 936 16552
rect 976 16520 1008 16552
rect 1048 16520 1080 16552
rect 1120 16520 1152 16552
rect 1192 16520 1224 16552
rect 1264 16520 1296 16552
rect 1336 16520 1368 16552
rect 1408 16520 1440 16552
rect 1480 16520 1512 16552
rect 1552 16520 1584 16552
rect 1624 16520 1656 16552
rect 1696 16520 1728 16552
rect 1768 16520 1800 16552
rect 1840 16520 1872 16552
rect 1912 16520 1944 16552
rect 1984 16520 2016 16552
rect 2056 16520 2088 16552
rect 2128 16520 2160 16552
rect 2200 16520 2232 16552
rect 2272 16520 2304 16552
rect 2344 16520 2376 16552
rect 2416 16520 2448 16552
rect 2488 16520 2520 16552
rect 2560 16520 2592 16552
rect 2632 16520 2664 16552
rect 2704 16520 2736 16552
rect 2776 16520 2808 16552
rect 2848 16520 2880 16552
rect 2920 16520 2952 16552
rect 2992 16520 3024 16552
rect 3064 16520 3096 16552
rect 3136 16520 3168 16552
rect 3208 16520 3240 16552
rect 3280 16520 3312 16552
rect 3352 16520 3384 16552
rect 3424 16520 3456 16552
rect 3496 16520 3528 16552
rect 3568 16520 3600 16552
rect 3640 16520 3672 16552
rect 3712 16520 3744 16552
rect 3784 16520 3816 16552
rect 3856 16520 3888 16552
rect 112 16448 144 16480
rect 184 16448 216 16480
rect 256 16448 288 16480
rect 328 16448 360 16480
rect 400 16448 432 16480
rect 472 16448 504 16480
rect 544 16448 576 16480
rect 616 16448 648 16480
rect 688 16448 720 16480
rect 760 16448 792 16480
rect 832 16448 864 16480
rect 904 16448 936 16480
rect 976 16448 1008 16480
rect 1048 16448 1080 16480
rect 1120 16448 1152 16480
rect 1192 16448 1224 16480
rect 1264 16448 1296 16480
rect 1336 16448 1368 16480
rect 1408 16448 1440 16480
rect 1480 16448 1512 16480
rect 1552 16448 1584 16480
rect 1624 16448 1656 16480
rect 1696 16448 1728 16480
rect 1768 16448 1800 16480
rect 1840 16448 1872 16480
rect 1912 16448 1944 16480
rect 1984 16448 2016 16480
rect 2056 16448 2088 16480
rect 2128 16448 2160 16480
rect 2200 16448 2232 16480
rect 2272 16448 2304 16480
rect 2344 16448 2376 16480
rect 2416 16448 2448 16480
rect 2488 16448 2520 16480
rect 2560 16448 2592 16480
rect 2632 16448 2664 16480
rect 2704 16448 2736 16480
rect 2776 16448 2808 16480
rect 2848 16448 2880 16480
rect 2920 16448 2952 16480
rect 2992 16448 3024 16480
rect 3064 16448 3096 16480
rect 3136 16448 3168 16480
rect 3208 16448 3240 16480
rect 3280 16448 3312 16480
rect 3352 16448 3384 16480
rect 3424 16448 3456 16480
rect 3496 16448 3528 16480
rect 3568 16448 3600 16480
rect 3640 16448 3672 16480
rect 3712 16448 3744 16480
rect 3784 16448 3816 16480
rect 3856 16448 3888 16480
rect 112 16376 144 16408
rect 184 16376 216 16408
rect 256 16376 288 16408
rect 328 16376 360 16408
rect 400 16376 432 16408
rect 472 16376 504 16408
rect 544 16376 576 16408
rect 616 16376 648 16408
rect 688 16376 720 16408
rect 760 16376 792 16408
rect 832 16376 864 16408
rect 904 16376 936 16408
rect 976 16376 1008 16408
rect 1048 16376 1080 16408
rect 1120 16376 1152 16408
rect 1192 16376 1224 16408
rect 1264 16376 1296 16408
rect 1336 16376 1368 16408
rect 1408 16376 1440 16408
rect 1480 16376 1512 16408
rect 1552 16376 1584 16408
rect 1624 16376 1656 16408
rect 1696 16376 1728 16408
rect 1768 16376 1800 16408
rect 1840 16376 1872 16408
rect 1912 16376 1944 16408
rect 1984 16376 2016 16408
rect 2056 16376 2088 16408
rect 2128 16376 2160 16408
rect 2200 16376 2232 16408
rect 2272 16376 2304 16408
rect 2344 16376 2376 16408
rect 2416 16376 2448 16408
rect 2488 16376 2520 16408
rect 2560 16376 2592 16408
rect 2632 16376 2664 16408
rect 2704 16376 2736 16408
rect 2776 16376 2808 16408
rect 2848 16376 2880 16408
rect 2920 16376 2952 16408
rect 2992 16376 3024 16408
rect 3064 16376 3096 16408
rect 3136 16376 3168 16408
rect 3208 16376 3240 16408
rect 3280 16376 3312 16408
rect 3352 16376 3384 16408
rect 3424 16376 3456 16408
rect 3496 16376 3528 16408
rect 3568 16376 3600 16408
rect 3640 16376 3672 16408
rect 3712 16376 3744 16408
rect 3784 16376 3816 16408
rect 3856 16376 3888 16408
rect 112 16304 144 16336
rect 184 16304 216 16336
rect 256 16304 288 16336
rect 328 16304 360 16336
rect 400 16304 432 16336
rect 472 16304 504 16336
rect 544 16304 576 16336
rect 616 16304 648 16336
rect 688 16304 720 16336
rect 760 16304 792 16336
rect 832 16304 864 16336
rect 904 16304 936 16336
rect 976 16304 1008 16336
rect 1048 16304 1080 16336
rect 1120 16304 1152 16336
rect 1192 16304 1224 16336
rect 1264 16304 1296 16336
rect 1336 16304 1368 16336
rect 1408 16304 1440 16336
rect 1480 16304 1512 16336
rect 1552 16304 1584 16336
rect 1624 16304 1656 16336
rect 1696 16304 1728 16336
rect 1768 16304 1800 16336
rect 1840 16304 1872 16336
rect 1912 16304 1944 16336
rect 1984 16304 2016 16336
rect 2056 16304 2088 16336
rect 2128 16304 2160 16336
rect 2200 16304 2232 16336
rect 2272 16304 2304 16336
rect 2344 16304 2376 16336
rect 2416 16304 2448 16336
rect 2488 16304 2520 16336
rect 2560 16304 2592 16336
rect 2632 16304 2664 16336
rect 2704 16304 2736 16336
rect 2776 16304 2808 16336
rect 2848 16304 2880 16336
rect 2920 16304 2952 16336
rect 2992 16304 3024 16336
rect 3064 16304 3096 16336
rect 3136 16304 3168 16336
rect 3208 16304 3240 16336
rect 3280 16304 3312 16336
rect 3352 16304 3384 16336
rect 3424 16304 3456 16336
rect 3496 16304 3528 16336
rect 3568 16304 3600 16336
rect 3640 16304 3672 16336
rect 3712 16304 3744 16336
rect 3784 16304 3816 16336
rect 3856 16304 3888 16336
rect 112 16232 144 16264
rect 184 16232 216 16264
rect 256 16232 288 16264
rect 328 16232 360 16264
rect 400 16232 432 16264
rect 472 16232 504 16264
rect 544 16232 576 16264
rect 616 16232 648 16264
rect 688 16232 720 16264
rect 760 16232 792 16264
rect 832 16232 864 16264
rect 904 16232 936 16264
rect 976 16232 1008 16264
rect 1048 16232 1080 16264
rect 1120 16232 1152 16264
rect 1192 16232 1224 16264
rect 1264 16232 1296 16264
rect 1336 16232 1368 16264
rect 1408 16232 1440 16264
rect 1480 16232 1512 16264
rect 1552 16232 1584 16264
rect 1624 16232 1656 16264
rect 1696 16232 1728 16264
rect 1768 16232 1800 16264
rect 1840 16232 1872 16264
rect 1912 16232 1944 16264
rect 1984 16232 2016 16264
rect 2056 16232 2088 16264
rect 2128 16232 2160 16264
rect 2200 16232 2232 16264
rect 2272 16232 2304 16264
rect 2344 16232 2376 16264
rect 2416 16232 2448 16264
rect 2488 16232 2520 16264
rect 2560 16232 2592 16264
rect 2632 16232 2664 16264
rect 2704 16232 2736 16264
rect 2776 16232 2808 16264
rect 2848 16232 2880 16264
rect 2920 16232 2952 16264
rect 2992 16232 3024 16264
rect 3064 16232 3096 16264
rect 3136 16232 3168 16264
rect 3208 16232 3240 16264
rect 3280 16232 3312 16264
rect 3352 16232 3384 16264
rect 3424 16232 3456 16264
rect 3496 16232 3528 16264
rect 3568 16232 3600 16264
rect 3640 16232 3672 16264
rect 3712 16232 3744 16264
rect 3784 16232 3816 16264
rect 3856 16232 3888 16264
rect 112 16160 144 16192
rect 184 16160 216 16192
rect 256 16160 288 16192
rect 328 16160 360 16192
rect 400 16160 432 16192
rect 472 16160 504 16192
rect 544 16160 576 16192
rect 616 16160 648 16192
rect 688 16160 720 16192
rect 760 16160 792 16192
rect 832 16160 864 16192
rect 904 16160 936 16192
rect 976 16160 1008 16192
rect 1048 16160 1080 16192
rect 1120 16160 1152 16192
rect 1192 16160 1224 16192
rect 1264 16160 1296 16192
rect 1336 16160 1368 16192
rect 1408 16160 1440 16192
rect 1480 16160 1512 16192
rect 1552 16160 1584 16192
rect 1624 16160 1656 16192
rect 1696 16160 1728 16192
rect 1768 16160 1800 16192
rect 1840 16160 1872 16192
rect 1912 16160 1944 16192
rect 1984 16160 2016 16192
rect 2056 16160 2088 16192
rect 2128 16160 2160 16192
rect 2200 16160 2232 16192
rect 2272 16160 2304 16192
rect 2344 16160 2376 16192
rect 2416 16160 2448 16192
rect 2488 16160 2520 16192
rect 2560 16160 2592 16192
rect 2632 16160 2664 16192
rect 2704 16160 2736 16192
rect 2776 16160 2808 16192
rect 2848 16160 2880 16192
rect 2920 16160 2952 16192
rect 2992 16160 3024 16192
rect 3064 16160 3096 16192
rect 3136 16160 3168 16192
rect 3208 16160 3240 16192
rect 3280 16160 3312 16192
rect 3352 16160 3384 16192
rect 3424 16160 3456 16192
rect 3496 16160 3528 16192
rect 3568 16160 3600 16192
rect 3640 16160 3672 16192
rect 3712 16160 3744 16192
rect 3784 16160 3816 16192
rect 3856 16160 3888 16192
rect 112 16088 144 16120
rect 184 16088 216 16120
rect 256 16088 288 16120
rect 328 16088 360 16120
rect 400 16088 432 16120
rect 472 16088 504 16120
rect 544 16088 576 16120
rect 616 16088 648 16120
rect 688 16088 720 16120
rect 760 16088 792 16120
rect 832 16088 864 16120
rect 904 16088 936 16120
rect 976 16088 1008 16120
rect 1048 16088 1080 16120
rect 1120 16088 1152 16120
rect 1192 16088 1224 16120
rect 1264 16088 1296 16120
rect 1336 16088 1368 16120
rect 1408 16088 1440 16120
rect 1480 16088 1512 16120
rect 1552 16088 1584 16120
rect 1624 16088 1656 16120
rect 1696 16088 1728 16120
rect 1768 16088 1800 16120
rect 1840 16088 1872 16120
rect 1912 16088 1944 16120
rect 1984 16088 2016 16120
rect 2056 16088 2088 16120
rect 2128 16088 2160 16120
rect 2200 16088 2232 16120
rect 2272 16088 2304 16120
rect 2344 16088 2376 16120
rect 2416 16088 2448 16120
rect 2488 16088 2520 16120
rect 2560 16088 2592 16120
rect 2632 16088 2664 16120
rect 2704 16088 2736 16120
rect 2776 16088 2808 16120
rect 2848 16088 2880 16120
rect 2920 16088 2952 16120
rect 2992 16088 3024 16120
rect 3064 16088 3096 16120
rect 3136 16088 3168 16120
rect 3208 16088 3240 16120
rect 3280 16088 3312 16120
rect 3352 16088 3384 16120
rect 3424 16088 3456 16120
rect 3496 16088 3528 16120
rect 3568 16088 3600 16120
rect 3640 16088 3672 16120
rect 3712 16088 3744 16120
rect 3784 16088 3816 16120
rect 3856 16088 3888 16120
rect 112 16016 144 16048
rect 184 16016 216 16048
rect 256 16016 288 16048
rect 328 16016 360 16048
rect 400 16016 432 16048
rect 472 16016 504 16048
rect 544 16016 576 16048
rect 616 16016 648 16048
rect 688 16016 720 16048
rect 760 16016 792 16048
rect 832 16016 864 16048
rect 904 16016 936 16048
rect 976 16016 1008 16048
rect 1048 16016 1080 16048
rect 1120 16016 1152 16048
rect 1192 16016 1224 16048
rect 1264 16016 1296 16048
rect 1336 16016 1368 16048
rect 1408 16016 1440 16048
rect 1480 16016 1512 16048
rect 1552 16016 1584 16048
rect 1624 16016 1656 16048
rect 1696 16016 1728 16048
rect 1768 16016 1800 16048
rect 1840 16016 1872 16048
rect 1912 16016 1944 16048
rect 1984 16016 2016 16048
rect 2056 16016 2088 16048
rect 2128 16016 2160 16048
rect 2200 16016 2232 16048
rect 2272 16016 2304 16048
rect 2344 16016 2376 16048
rect 2416 16016 2448 16048
rect 2488 16016 2520 16048
rect 2560 16016 2592 16048
rect 2632 16016 2664 16048
rect 2704 16016 2736 16048
rect 2776 16016 2808 16048
rect 2848 16016 2880 16048
rect 2920 16016 2952 16048
rect 2992 16016 3024 16048
rect 3064 16016 3096 16048
rect 3136 16016 3168 16048
rect 3208 16016 3240 16048
rect 3280 16016 3312 16048
rect 3352 16016 3384 16048
rect 3424 16016 3456 16048
rect 3496 16016 3528 16048
rect 3568 16016 3600 16048
rect 3640 16016 3672 16048
rect 3712 16016 3744 16048
rect 3784 16016 3816 16048
rect 3856 16016 3888 16048
rect 112 15944 144 15976
rect 184 15944 216 15976
rect 256 15944 288 15976
rect 328 15944 360 15976
rect 400 15944 432 15976
rect 472 15944 504 15976
rect 544 15944 576 15976
rect 616 15944 648 15976
rect 688 15944 720 15976
rect 760 15944 792 15976
rect 832 15944 864 15976
rect 904 15944 936 15976
rect 976 15944 1008 15976
rect 1048 15944 1080 15976
rect 1120 15944 1152 15976
rect 1192 15944 1224 15976
rect 1264 15944 1296 15976
rect 1336 15944 1368 15976
rect 1408 15944 1440 15976
rect 1480 15944 1512 15976
rect 1552 15944 1584 15976
rect 1624 15944 1656 15976
rect 1696 15944 1728 15976
rect 1768 15944 1800 15976
rect 1840 15944 1872 15976
rect 1912 15944 1944 15976
rect 1984 15944 2016 15976
rect 2056 15944 2088 15976
rect 2128 15944 2160 15976
rect 2200 15944 2232 15976
rect 2272 15944 2304 15976
rect 2344 15944 2376 15976
rect 2416 15944 2448 15976
rect 2488 15944 2520 15976
rect 2560 15944 2592 15976
rect 2632 15944 2664 15976
rect 2704 15944 2736 15976
rect 2776 15944 2808 15976
rect 2848 15944 2880 15976
rect 2920 15944 2952 15976
rect 2992 15944 3024 15976
rect 3064 15944 3096 15976
rect 3136 15944 3168 15976
rect 3208 15944 3240 15976
rect 3280 15944 3312 15976
rect 3352 15944 3384 15976
rect 3424 15944 3456 15976
rect 3496 15944 3528 15976
rect 3568 15944 3600 15976
rect 3640 15944 3672 15976
rect 3712 15944 3744 15976
rect 3784 15944 3816 15976
rect 3856 15944 3888 15976
rect 112 15872 144 15904
rect 184 15872 216 15904
rect 256 15872 288 15904
rect 328 15872 360 15904
rect 400 15872 432 15904
rect 472 15872 504 15904
rect 544 15872 576 15904
rect 616 15872 648 15904
rect 688 15872 720 15904
rect 760 15872 792 15904
rect 832 15872 864 15904
rect 904 15872 936 15904
rect 976 15872 1008 15904
rect 1048 15872 1080 15904
rect 1120 15872 1152 15904
rect 1192 15872 1224 15904
rect 1264 15872 1296 15904
rect 1336 15872 1368 15904
rect 1408 15872 1440 15904
rect 1480 15872 1512 15904
rect 1552 15872 1584 15904
rect 1624 15872 1656 15904
rect 1696 15872 1728 15904
rect 1768 15872 1800 15904
rect 1840 15872 1872 15904
rect 1912 15872 1944 15904
rect 1984 15872 2016 15904
rect 2056 15872 2088 15904
rect 2128 15872 2160 15904
rect 2200 15872 2232 15904
rect 2272 15872 2304 15904
rect 2344 15872 2376 15904
rect 2416 15872 2448 15904
rect 2488 15872 2520 15904
rect 2560 15872 2592 15904
rect 2632 15872 2664 15904
rect 2704 15872 2736 15904
rect 2776 15872 2808 15904
rect 2848 15872 2880 15904
rect 2920 15872 2952 15904
rect 2992 15872 3024 15904
rect 3064 15872 3096 15904
rect 3136 15872 3168 15904
rect 3208 15872 3240 15904
rect 3280 15872 3312 15904
rect 3352 15872 3384 15904
rect 3424 15872 3456 15904
rect 3496 15872 3528 15904
rect 3568 15872 3600 15904
rect 3640 15872 3672 15904
rect 3712 15872 3744 15904
rect 3784 15872 3816 15904
rect 3856 15872 3888 15904
rect 112 15800 144 15832
rect 184 15800 216 15832
rect 256 15800 288 15832
rect 328 15800 360 15832
rect 400 15800 432 15832
rect 472 15800 504 15832
rect 544 15800 576 15832
rect 616 15800 648 15832
rect 688 15800 720 15832
rect 760 15800 792 15832
rect 832 15800 864 15832
rect 904 15800 936 15832
rect 976 15800 1008 15832
rect 1048 15800 1080 15832
rect 1120 15800 1152 15832
rect 1192 15800 1224 15832
rect 1264 15800 1296 15832
rect 1336 15800 1368 15832
rect 1408 15800 1440 15832
rect 1480 15800 1512 15832
rect 1552 15800 1584 15832
rect 1624 15800 1656 15832
rect 1696 15800 1728 15832
rect 1768 15800 1800 15832
rect 1840 15800 1872 15832
rect 1912 15800 1944 15832
rect 1984 15800 2016 15832
rect 2056 15800 2088 15832
rect 2128 15800 2160 15832
rect 2200 15800 2232 15832
rect 2272 15800 2304 15832
rect 2344 15800 2376 15832
rect 2416 15800 2448 15832
rect 2488 15800 2520 15832
rect 2560 15800 2592 15832
rect 2632 15800 2664 15832
rect 2704 15800 2736 15832
rect 2776 15800 2808 15832
rect 2848 15800 2880 15832
rect 2920 15800 2952 15832
rect 2992 15800 3024 15832
rect 3064 15800 3096 15832
rect 3136 15800 3168 15832
rect 3208 15800 3240 15832
rect 3280 15800 3312 15832
rect 3352 15800 3384 15832
rect 3424 15800 3456 15832
rect 3496 15800 3528 15832
rect 3568 15800 3600 15832
rect 3640 15800 3672 15832
rect 3712 15800 3744 15832
rect 3784 15800 3816 15832
rect 3856 15800 3888 15832
rect 112 15728 144 15760
rect 184 15728 216 15760
rect 256 15728 288 15760
rect 328 15728 360 15760
rect 400 15728 432 15760
rect 472 15728 504 15760
rect 544 15728 576 15760
rect 616 15728 648 15760
rect 688 15728 720 15760
rect 760 15728 792 15760
rect 832 15728 864 15760
rect 904 15728 936 15760
rect 976 15728 1008 15760
rect 1048 15728 1080 15760
rect 1120 15728 1152 15760
rect 1192 15728 1224 15760
rect 1264 15728 1296 15760
rect 1336 15728 1368 15760
rect 1408 15728 1440 15760
rect 1480 15728 1512 15760
rect 1552 15728 1584 15760
rect 1624 15728 1656 15760
rect 1696 15728 1728 15760
rect 1768 15728 1800 15760
rect 1840 15728 1872 15760
rect 1912 15728 1944 15760
rect 1984 15728 2016 15760
rect 2056 15728 2088 15760
rect 2128 15728 2160 15760
rect 2200 15728 2232 15760
rect 2272 15728 2304 15760
rect 2344 15728 2376 15760
rect 2416 15728 2448 15760
rect 2488 15728 2520 15760
rect 2560 15728 2592 15760
rect 2632 15728 2664 15760
rect 2704 15728 2736 15760
rect 2776 15728 2808 15760
rect 2848 15728 2880 15760
rect 2920 15728 2952 15760
rect 2992 15728 3024 15760
rect 3064 15728 3096 15760
rect 3136 15728 3168 15760
rect 3208 15728 3240 15760
rect 3280 15728 3312 15760
rect 3352 15728 3384 15760
rect 3424 15728 3456 15760
rect 3496 15728 3528 15760
rect 3568 15728 3600 15760
rect 3640 15728 3672 15760
rect 3712 15728 3744 15760
rect 3784 15728 3816 15760
rect 3856 15728 3888 15760
rect 112 15656 144 15688
rect 184 15656 216 15688
rect 256 15656 288 15688
rect 328 15656 360 15688
rect 400 15656 432 15688
rect 472 15656 504 15688
rect 544 15656 576 15688
rect 616 15656 648 15688
rect 688 15656 720 15688
rect 760 15656 792 15688
rect 832 15656 864 15688
rect 904 15656 936 15688
rect 976 15656 1008 15688
rect 1048 15656 1080 15688
rect 1120 15656 1152 15688
rect 1192 15656 1224 15688
rect 1264 15656 1296 15688
rect 1336 15656 1368 15688
rect 1408 15656 1440 15688
rect 1480 15656 1512 15688
rect 1552 15656 1584 15688
rect 1624 15656 1656 15688
rect 1696 15656 1728 15688
rect 1768 15656 1800 15688
rect 1840 15656 1872 15688
rect 1912 15656 1944 15688
rect 1984 15656 2016 15688
rect 2056 15656 2088 15688
rect 2128 15656 2160 15688
rect 2200 15656 2232 15688
rect 2272 15656 2304 15688
rect 2344 15656 2376 15688
rect 2416 15656 2448 15688
rect 2488 15656 2520 15688
rect 2560 15656 2592 15688
rect 2632 15656 2664 15688
rect 2704 15656 2736 15688
rect 2776 15656 2808 15688
rect 2848 15656 2880 15688
rect 2920 15656 2952 15688
rect 2992 15656 3024 15688
rect 3064 15656 3096 15688
rect 3136 15656 3168 15688
rect 3208 15656 3240 15688
rect 3280 15656 3312 15688
rect 3352 15656 3384 15688
rect 3424 15656 3456 15688
rect 3496 15656 3528 15688
rect 3568 15656 3600 15688
rect 3640 15656 3672 15688
rect 3712 15656 3744 15688
rect 3784 15656 3816 15688
rect 3856 15656 3888 15688
rect 112 15584 144 15616
rect 184 15584 216 15616
rect 256 15584 288 15616
rect 328 15584 360 15616
rect 400 15584 432 15616
rect 472 15584 504 15616
rect 544 15584 576 15616
rect 616 15584 648 15616
rect 688 15584 720 15616
rect 760 15584 792 15616
rect 832 15584 864 15616
rect 904 15584 936 15616
rect 976 15584 1008 15616
rect 1048 15584 1080 15616
rect 1120 15584 1152 15616
rect 1192 15584 1224 15616
rect 1264 15584 1296 15616
rect 1336 15584 1368 15616
rect 1408 15584 1440 15616
rect 1480 15584 1512 15616
rect 1552 15584 1584 15616
rect 1624 15584 1656 15616
rect 1696 15584 1728 15616
rect 1768 15584 1800 15616
rect 1840 15584 1872 15616
rect 1912 15584 1944 15616
rect 1984 15584 2016 15616
rect 2056 15584 2088 15616
rect 2128 15584 2160 15616
rect 2200 15584 2232 15616
rect 2272 15584 2304 15616
rect 2344 15584 2376 15616
rect 2416 15584 2448 15616
rect 2488 15584 2520 15616
rect 2560 15584 2592 15616
rect 2632 15584 2664 15616
rect 2704 15584 2736 15616
rect 2776 15584 2808 15616
rect 2848 15584 2880 15616
rect 2920 15584 2952 15616
rect 2992 15584 3024 15616
rect 3064 15584 3096 15616
rect 3136 15584 3168 15616
rect 3208 15584 3240 15616
rect 3280 15584 3312 15616
rect 3352 15584 3384 15616
rect 3424 15584 3456 15616
rect 3496 15584 3528 15616
rect 3568 15584 3600 15616
rect 3640 15584 3672 15616
rect 3712 15584 3744 15616
rect 3784 15584 3816 15616
rect 3856 15584 3888 15616
rect 112 15512 144 15544
rect 184 15512 216 15544
rect 256 15512 288 15544
rect 328 15512 360 15544
rect 400 15512 432 15544
rect 472 15512 504 15544
rect 544 15512 576 15544
rect 616 15512 648 15544
rect 688 15512 720 15544
rect 760 15512 792 15544
rect 832 15512 864 15544
rect 904 15512 936 15544
rect 976 15512 1008 15544
rect 1048 15512 1080 15544
rect 1120 15512 1152 15544
rect 1192 15512 1224 15544
rect 1264 15512 1296 15544
rect 1336 15512 1368 15544
rect 1408 15512 1440 15544
rect 1480 15512 1512 15544
rect 1552 15512 1584 15544
rect 1624 15512 1656 15544
rect 1696 15512 1728 15544
rect 1768 15512 1800 15544
rect 1840 15512 1872 15544
rect 1912 15512 1944 15544
rect 1984 15512 2016 15544
rect 2056 15512 2088 15544
rect 2128 15512 2160 15544
rect 2200 15512 2232 15544
rect 2272 15512 2304 15544
rect 2344 15512 2376 15544
rect 2416 15512 2448 15544
rect 2488 15512 2520 15544
rect 2560 15512 2592 15544
rect 2632 15512 2664 15544
rect 2704 15512 2736 15544
rect 2776 15512 2808 15544
rect 2848 15512 2880 15544
rect 2920 15512 2952 15544
rect 2992 15512 3024 15544
rect 3064 15512 3096 15544
rect 3136 15512 3168 15544
rect 3208 15512 3240 15544
rect 3280 15512 3312 15544
rect 3352 15512 3384 15544
rect 3424 15512 3456 15544
rect 3496 15512 3528 15544
rect 3568 15512 3600 15544
rect 3640 15512 3672 15544
rect 3712 15512 3744 15544
rect 3784 15512 3816 15544
rect 3856 15512 3888 15544
rect 112 15440 144 15472
rect 184 15440 216 15472
rect 256 15440 288 15472
rect 328 15440 360 15472
rect 400 15440 432 15472
rect 472 15440 504 15472
rect 544 15440 576 15472
rect 616 15440 648 15472
rect 688 15440 720 15472
rect 760 15440 792 15472
rect 832 15440 864 15472
rect 904 15440 936 15472
rect 976 15440 1008 15472
rect 1048 15440 1080 15472
rect 1120 15440 1152 15472
rect 1192 15440 1224 15472
rect 1264 15440 1296 15472
rect 1336 15440 1368 15472
rect 1408 15440 1440 15472
rect 1480 15440 1512 15472
rect 1552 15440 1584 15472
rect 1624 15440 1656 15472
rect 1696 15440 1728 15472
rect 1768 15440 1800 15472
rect 1840 15440 1872 15472
rect 1912 15440 1944 15472
rect 1984 15440 2016 15472
rect 2056 15440 2088 15472
rect 2128 15440 2160 15472
rect 2200 15440 2232 15472
rect 2272 15440 2304 15472
rect 2344 15440 2376 15472
rect 2416 15440 2448 15472
rect 2488 15440 2520 15472
rect 2560 15440 2592 15472
rect 2632 15440 2664 15472
rect 2704 15440 2736 15472
rect 2776 15440 2808 15472
rect 2848 15440 2880 15472
rect 2920 15440 2952 15472
rect 2992 15440 3024 15472
rect 3064 15440 3096 15472
rect 3136 15440 3168 15472
rect 3208 15440 3240 15472
rect 3280 15440 3312 15472
rect 3352 15440 3384 15472
rect 3424 15440 3456 15472
rect 3496 15440 3528 15472
rect 3568 15440 3600 15472
rect 3640 15440 3672 15472
rect 3712 15440 3744 15472
rect 3784 15440 3816 15472
rect 3856 15440 3888 15472
rect 112 15368 144 15400
rect 184 15368 216 15400
rect 256 15368 288 15400
rect 328 15368 360 15400
rect 400 15368 432 15400
rect 472 15368 504 15400
rect 544 15368 576 15400
rect 616 15368 648 15400
rect 688 15368 720 15400
rect 760 15368 792 15400
rect 832 15368 864 15400
rect 904 15368 936 15400
rect 976 15368 1008 15400
rect 1048 15368 1080 15400
rect 1120 15368 1152 15400
rect 1192 15368 1224 15400
rect 1264 15368 1296 15400
rect 1336 15368 1368 15400
rect 1408 15368 1440 15400
rect 1480 15368 1512 15400
rect 1552 15368 1584 15400
rect 1624 15368 1656 15400
rect 1696 15368 1728 15400
rect 1768 15368 1800 15400
rect 1840 15368 1872 15400
rect 1912 15368 1944 15400
rect 1984 15368 2016 15400
rect 2056 15368 2088 15400
rect 2128 15368 2160 15400
rect 2200 15368 2232 15400
rect 2272 15368 2304 15400
rect 2344 15368 2376 15400
rect 2416 15368 2448 15400
rect 2488 15368 2520 15400
rect 2560 15368 2592 15400
rect 2632 15368 2664 15400
rect 2704 15368 2736 15400
rect 2776 15368 2808 15400
rect 2848 15368 2880 15400
rect 2920 15368 2952 15400
rect 2992 15368 3024 15400
rect 3064 15368 3096 15400
rect 3136 15368 3168 15400
rect 3208 15368 3240 15400
rect 3280 15368 3312 15400
rect 3352 15368 3384 15400
rect 3424 15368 3456 15400
rect 3496 15368 3528 15400
rect 3568 15368 3600 15400
rect 3640 15368 3672 15400
rect 3712 15368 3744 15400
rect 3784 15368 3816 15400
rect 3856 15368 3888 15400
rect 112 15296 144 15328
rect 184 15296 216 15328
rect 256 15296 288 15328
rect 328 15296 360 15328
rect 400 15296 432 15328
rect 472 15296 504 15328
rect 544 15296 576 15328
rect 616 15296 648 15328
rect 688 15296 720 15328
rect 760 15296 792 15328
rect 832 15296 864 15328
rect 904 15296 936 15328
rect 976 15296 1008 15328
rect 1048 15296 1080 15328
rect 1120 15296 1152 15328
rect 1192 15296 1224 15328
rect 1264 15296 1296 15328
rect 1336 15296 1368 15328
rect 1408 15296 1440 15328
rect 1480 15296 1512 15328
rect 1552 15296 1584 15328
rect 1624 15296 1656 15328
rect 1696 15296 1728 15328
rect 1768 15296 1800 15328
rect 1840 15296 1872 15328
rect 1912 15296 1944 15328
rect 1984 15296 2016 15328
rect 2056 15296 2088 15328
rect 2128 15296 2160 15328
rect 2200 15296 2232 15328
rect 2272 15296 2304 15328
rect 2344 15296 2376 15328
rect 2416 15296 2448 15328
rect 2488 15296 2520 15328
rect 2560 15296 2592 15328
rect 2632 15296 2664 15328
rect 2704 15296 2736 15328
rect 2776 15296 2808 15328
rect 2848 15296 2880 15328
rect 2920 15296 2952 15328
rect 2992 15296 3024 15328
rect 3064 15296 3096 15328
rect 3136 15296 3168 15328
rect 3208 15296 3240 15328
rect 3280 15296 3312 15328
rect 3352 15296 3384 15328
rect 3424 15296 3456 15328
rect 3496 15296 3528 15328
rect 3568 15296 3600 15328
rect 3640 15296 3672 15328
rect 3712 15296 3744 15328
rect 3784 15296 3816 15328
rect 3856 15296 3888 15328
rect 112 15224 144 15256
rect 184 15224 216 15256
rect 256 15224 288 15256
rect 328 15224 360 15256
rect 400 15224 432 15256
rect 472 15224 504 15256
rect 544 15224 576 15256
rect 616 15224 648 15256
rect 688 15224 720 15256
rect 760 15224 792 15256
rect 832 15224 864 15256
rect 904 15224 936 15256
rect 976 15224 1008 15256
rect 1048 15224 1080 15256
rect 1120 15224 1152 15256
rect 1192 15224 1224 15256
rect 1264 15224 1296 15256
rect 1336 15224 1368 15256
rect 1408 15224 1440 15256
rect 1480 15224 1512 15256
rect 1552 15224 1584 15256
rect 1624 15224 1656 15256
rect 1696 15224 1728 15256
rect 1768 15224 1800 15256
rect 1840 15224 1872 15256
rect 1912 15224 1944 15256
rect 1984 15224 2016 15256
rect 2056 15224 2088 15256
rect 2128 15224 2160 15256
rect 2200 15224 2232 15256
rect 2272 15224 2304 15256
rect 2344 15224 2376 15256
rect 2416 15224 2448 15256
rect 2488 15224 2520 15256
rect 2560 15224 2592 15256
rect 2632 15224 2664 15256
rect 2704 15224 2736 15256
rect 2776 15224 2808 15256
rect 2848 15224 2880 15256
rect 2920 15224 2952 15256
rect 2992 15224 3024 15256
rect 3064 15224 3096 15256
rect 3136 15224 3168 15256
rect 3208 15224 3240 15256
rect 3280 15224 3312 15256
rect 3352 15224 3384 15256
rect 3424 15224 3456 15256
rect 3496 15224 3528 15256
rect 3568 15224 3600 15256
rect 3640 15224 3672 15256
rect 3712 15224 3744 15256
rect 3784 15224 3816 15256
rect 3856 15224 3888 15256
rect 112 15152 144 15184
rect 184 15152 216 15184
rect 256 15152 288 15184
rect 328 15152 360 15184
rect 400 15152 432 15184
rect 472 15152 504 15184
rect 544 15152 576 15184
rect 616 15152 648 15184
rect 688 15152 720 15184
rect 760 15152 792 15184
rect 832 15152 864 15184
rect 904 15152 936 15184
rect 976 15152 1008 15184
rect 1048 15152 1080 15184
rect 1120 15152 1152 15184
rect 1192 15152 1224 15184
rect 1264 15152 1296 15184
rect 1336 15152 1368 15184
rect 1408 15152 1440 15184
rect 1480 15152 1512 15184
rect 1552 15152 1584 15184
rect 1624 15152 1656 15184
rect 1696 15152 1728 15184
rect 1768 15152 1800 15184
rect 1840 15152 1872 15184
rect 1912 15152 1944 15184
rect 1984 15152 2016 15184
rect 2056 15152 2088 15184
rect 2128 15152 2160 15184
rect 2200 15152 2232 15184
rect 2272 15152 2304 15184
rect 2344 15152 2376 15184
rect 2416 15152 2448 15184
rect 2488 15152 2520 15184
rect 2560 15152 2592 15184
rect 2632 15152 2664 15184
rect 2704 15152 2736 15184
rect 2776 15152 2808 15184
rect 2848 15152 2880 15184
rect 2920 15152 2952 15184
rect 2992 15152 3024 15184
rect 3064 15152 3096 15184
rect 3136 15152 3168 15184
rect 3208 15152 3240 15184
rect 3280 15152 3312 15184
rect 3352 15152 3384 15184
rect 3424 15152 3456 15184
rect 3496 15152 3528 15184
rect 3568 15152 3600 15184
rect 3640 15152 3672 15184
rect 3712 15152 3744 15184
rect 3784 15152 3816 15184
rect 3856 15152 3888 15184
rect 112 15080 144 15112
rect 184 15080 216 15112
rect 256 15080 288 15112
rect 328 15080 360 15112
rect 400 15080 432 15112
rect 472 15080 504 15112
rect 544 15080 576 15112
rect 616 15080 648 15112
rect 688 15080 720 15112
rect 760 15080 792 15112
rect 832 15080 864 15112
rect 904 15080 936 15112
rect 976 15080 1008 15112
rect 1048 15080 1080 15112
rect 1120 15080 1152 15112
rect 1192 15080 1224 15112
rect 1264 15080 1296 15112
rect 1336 15080 1368 15112
rect 1408 15080 1440 15112
rect 1480 15080 1512 15112
rect 1552 15080 1584 15112
rect 1624 15080 1656 15112
rect 1696 15080 1728 15112
rect 1768 15080 1800 15112
rect 1840 15080 1872 15112
rect 1912 15080 1944 15112
rect 1984 15080 2016 15112
rect 2056 15080 2088 15112
rect 2128 15080 2160 15112
rect 2200 15080 2232 15112
rect 2272 15080 2304 15112
rect 2344 15080 2376 15112
rect 2416 15080 2448 15112
rect 2488 15080 2520 15112
rect 2560 15080 2592 15112
rect 2632 15080 2664 15112
rect 2704 15080 2736 15112
rect 2776 15080 2808 15112
rect 2848 15080 2880 15112
rect 2920 15080 2952 15112
rect 2992 15080 3024 15112
rect 3064 15080 3096 15112
rect 3136 15080 3168 15112
rect 3208 15080 3240 15112
rect 3280 15080 3312 15112
rect 3352 15080 3384 15112
rect 3424 15080 3456 15112
rect 3496 15080 3528 15112
rect 3568 15080 3600 15112
rect 3640 15080 3672 15112
rect 3712 15080 3744 15112
rect 3784 15080 3816 15112
rect 3856 15080 3888 15112
rect 112 15008 144 15040
rect 184 15008 216 15040
rect 256 15008 288 15040
rect 328 15008 360 15040
rect 400 15008 432 15040
rect 472 15008 504 15040
rect 544 15008 576 15040
rect 616 15008 648 15040
rect 688 15008 720 15040
rect 760 15008 792 15040
rect 832 15008 864 15040
rect 904 15008 936 15040
rect 976 15008 1008 15040
rect 1048 15008 1080 15040
rect 1120 15008 1152 15040
rect 1192 15008 1224 15040
rect 1264 15008 1296 15040
rect 1336 15008 1368 15040
rect 1408 15008 1440 15040
rect 1480 15008 1512 15040
rect 1552 15008 1584 15040
rect 1624 15008 1656 15040
rect 1696 15008 1728 15040
rect 1768 15008 1800 15040
rect 1840 15008 1872 15040
rect 1912 15008 1944 15040
rect 1984 15008 2016 15040
rect 2056 15008 2088 15040
rect 2128 15008 2160 15040
rect 2200 15008 2232 15040
rect 2272 15008 2304 15040
rect 2344 15008 2376 15040
rect 2416 15008 2448 15040
rect 2488 15008 2520 15040
rect 2560 15008 2592 15040
rect 2632 15008 2664 15040
rect 2704 15008 2736 15040
rect 2776 15008 2808 15040
rect 2848 15008 2880 15040
rect 2920 15008 2952 15040
rect 2992 15008 3024 15040
rect 3064 15008 3096 15040
rect 3136 15008 3168 15040
rect 3208 15008 3240 15040
rect 3280 15008 3312 15040
rect 3352 15008 3384 15040
rect 3424 15008 3456 15040
rect 3496 15008 3528 15040
rect 3568 15008 3600 15040
rect 3640 15008 3672 15040
rect 3712 15008 3744 15040
rect 3784 15008 3816 15040
rect 3856 15008 3888 15040
rect 112 14936 144 14968
rect 184 14936 216 14968
rect 256 14936 288 14968
rect 328 14936 360 14968
rect 400 14936 432 14968
rect 472 14936 504 14968
rect 544 14936 576 14968
rect 616 14936 648 14968
rect 688 14936 720 14968
rect 760 14936 792 14968
rect 832 14936 864 14968
rect 904 14936 936 14968
rect 976 14936 1008 14968
rect 1048 14936 1080 14968
rect 1120 14936 1152 14968
rect 1192 14936 1224 14968
rect 1264 14936 1296 14968
rect 1336 14936 1368 14968
rect 1408 14936 1440 14968
rect 1480 14936 1512 14968
rect 1552 14936 1584 14968
rect 1624 14936 1656 14968
rect 1696 14936 1728 14968
rect 1768 14936 1800 14968
rect 1840 14936 1872 14968
rect 1912 14936 1944 14968
rect 1984 14936 2016 14968
rect 2056 14936 2088 14968
rect 2128 14936 2160 14968
rect 2200 14936 2232 14968
rect 2272 14936 2304 14968
rect 2344 14936 2376 14968
rect 2416 14936 2448 14968
rect 2488 14936 2520 14968
rect 2560 14936 2592 14968
rect 2632 14936 2664 14968
rect 2704 14936 2736 14968
rect 2776 14936 2808 14968
rect 2848 14936 2880 14968
rect 2920 14936 2952 14968
rect 2992 14936 3024 14968
rect 3064 14936 3096 14968
rect 3136 14936 3168 14968
rect 3208 14936 3240 14968
rect 3280 14936 3312 14968
rect 3352 14936 3384 14968
rect 3424 14936 3456 14968
rect 3496 14936 3528 14968
rect 3568 14936 3600 14968
rect 3640 14936 3672 14968
rect 3712 14936 3744 14968
rect 3784 14936 3816 14968
rect 3856 14936 3888 14968
rect 112 14864 144 14896
rect 184 14864 216 14896
rect 256 14864 288 14896
rect 328 14864 360 14896
rect 400 14864 432 14896
rect 472 14864 504 14896
rect 544 14864 576 14896
rect 616 14864 648 14896
rect 688 14864 720 14896
rect 760 14864 792 14896
rect 832 14864 864 14896
rect 904 14864 936 14896
rect 976 14864 1008 14896
rect 1048 14864 1080 14896
rect 1120 14864 1152 14896
rect 1192 14864 1224 14896
rect 1264 14864 1296 14896
rect 1336 14864 1368 14896
rect 1408 14864 1440 14896
rect 1480 14864 1512 14896
rect 1552 14864 1584 14896
rect 1624 14864 1656 14896
rect 1696 14864 1728 14896
rect 1768 14864 1800 14896
rect 1840 14864 1872 14896
rect 1912 14864 1944 14896
rect 1984 14864 2016 14896
rect 2056 14864 2088 14896
rect 2128 14864 2160 14896
rect 2200 14864 2232 14896
rect 2272 14864 2304 14896
rect 2344 14864 2376 14896
rect 2416 14864 2448 14896
rect 2488 14864 2520 14896
rect 2560 14864 2592 14896
rect 2632 14864 2664 14896
rect 2704 14864 2736 14896
rect 2776 14864 2808 14896
rect 2848 14864 2880 14896
rect 2920 14864 2952 14896
rect 2992 14864 3024 14896
rect 3064 14864 3096 14896
rect 3136 14864 3168 14896
rect 3208 14864 3240 14896
rect 3280 14864 3312 14896
rect 3352 14864 3384 14896
rect 3424 14864 3456 14896
rect 3496 14864 3528 14896
rect 3568 14864 3600 14896
rect 3640 14864 3672 14896
rect 3712 14864 3744 14896
rect 3784 14864 3816 14896
rect 3856 14864 3888 14896
rect 112 14792 144 14824
rect 184 14792 216 14824
rect 256 14792 288 14824
rect 328 14792 360 14824
rect 400 14792 432 14824
rect 472 14792 504 14824
rect 544 14792 576 14824
rect 616 14792 648 14824
rect 688 14792 720 14824
rect 760 14792 792 14824
rect 832 14792 864 14824
rect 904 14792 936 14824
rect 976 14792 1008 14824
rect 1048 14792 1080 14824
rect 1120 14792 1152 14824
rect 1192 14792 1224 14824
rect 1264 14792 1296 14824
rect 1336 14792 1368 14824
rect 1408 14792 1440 14824
rect 1480 14792 1512 14824
rect 1552 14792 1584 14824
rect 1624 14792 1656 14824
rect 1696 14792 1728 14824
rect 1768 14792 1800 14824
rect 1840 14792 1872 14824
rect 1912 14792 1944 14824
rect 1984 14792 2016 14824
rect 2056 14792 2088 14824
rect 2128 14792 2160 14824
rect 2200 14792 2232 14824
rect 2272 14792 2304 14824
rect 2344 14792 2376 14824
rect 2416 14792 2448 14824
rect 2488 14792 2520 14824
rect 2560 14792 2592 14824
rect 2632 14792 2664 14824
rect 2704 14792 2736 14824
rect 2776 14792 2808 14824
rect 2848 14792 2880 14824
rect 2920 14792 2952 14824
rect 2992 14792 3024 14824
rect 3064 14792 3096 14824
rect 3136 14792 3168 14824
rect 3208 14792 3240 14824
rect 3280 14792 3312 14824
rect 3352 14792 3384 14824
rect 3424 14792 3456 14824
rect 3496 14792 3528 14824
rect 3568 14792 3600 14824
rect 3640 14792 3672 14824
rect 3712 14792 3744 14824
rect 3784 14792 3816 14824
rect 3856 14792 3888 14824
rect 112 14720 144 14752
rect 184 14720 216 14752
rect 256 14720 288 14752
rect 328 14720 360 14752
rect 400 14720 432 14752
rect 472 14720 504 14752
rect 544 14720 576 14752
rect 616 14720 648 14752
rect 688 14720 720 14752
rect 760 14720 792 14752
rect 832 14720 864 14752
rect 904 14720 936 14752
rect 976 14720 1008 14752
rect 1048 14720 1080 14752
rect 1120 14720 1152 14752
rect 1192 14720 1224 14752
rect 1264 14720 1296 14752
rect 1336 14720 1368 14752
rect 1408 14720 1440 14752
rect 1480 14720 1512 14752
rect 1552 14720 1584 14752
rect 1624 14720 1656 14752
rect 1696 14720 1728 14752
rect 1768 14720 1800 14752
rect 1840 14720 1872 14752
rect 1912 14720 1944 14752
rect 1984 14720 2016 14752
rect 2056 14720 2088 14752
rect 2128 14720 2160 14752
rect 2200 14720 2232 14752
rect 2272 14720 2304 14752
rect 2344 14720 2376 14752
rect 2416 14720 2448 14752
rect 2488 14720 2520 14752
rect 2560 14720 2592 14752
rect 2632 14720 2664 14752
rect 2704 14720 2736 14752
rect 2776 14720 2808 14752
rect 2848 14720 2880 14752
rect 2920 14720 2952 14752
rect 2992 14720 3024 14752
rect 3064 14720 3096 14752
rect 3136 14720 3168 14752
rect 3208 14720 3240 14752
rect 3280 14720 3312 14752
rect 3352 14720 3384 14752
rect 3424 14720 3456 14752
rect 3496 14720 3528 14752
rect 3568 14720 3600 14752
rect 3640 14720 3672 14752
rect 3712 14720 3744 14752
rect 3784 14720 3816 14752
rect 3856 14720 3888 14752
rect 112 14648 144 14680
rect 184 14648 216 14680
rect 256 14648 288 14680
rect 328 14648 360 14680
rect 400 14648 432 14680
rect 472 14648 504 14680
rect 544 14648 576 14680
rect 616 14648 648 14680
rect 688 14648 720 14680
rect 760 14648 792 14680
rect 832 14648 864 14680
rect 904 14648 936 14680
rect 976 14648 1008 14680
rect 1048 14648 1080 14680
rect 1120 14648 1152 14680
rect 1192 14648 1224 14680
rect 1264 14648 1296 14680
rect 1336 14648 1368 14680
rect 1408 14648 1440 14680
rect 1480 14648 1512 14680
rect 1552 14648 1584 14680
rect 1624 14648 1656 14680
rect 1696 14648 1728 14680
rect 1768 14648 1800 14680
rect 1840 14648 1872 14680
rect 1912 14648 1944 14680
rect 1984 14648 2016 14680
rect 2056 14648 2088 14680
rect 2128 14648 2160 14680
rect 2200 14648 2232 14680
rect 2272 14648 2304 14680
rect 2344 14648 2376 14680
rect 2416 14648 2448 14680
rect 2488 14648 2520 14680
rect 2560 14648 2592 14680
rect 2632 14648 2664 14680
rect 2704 14648 2736 14680
rect 2776 14648 2808 14680
rect 2848 14648 2880 14680
rect 2920 14648 2952 14680
rect 2992 14648 3024 14680
rect 3064 14648 3096 14680
rect 3136 14648 3168 14680
rect 3208 14648 3240 14680
rect 3280 14648 3312 14680
rect 3352 14648 3384 14680
rect 3424 14648 3456 14680
rect 3496 14648 3528 14680
rect 3568 14648 3600 14680
rect 3640 14648 3672 14680
rect 3712 14648 3744 14680
rect 3784 14648 3816 14680
rect 3856 14648 3888 14680
rect 112 14576 144 14608
rect 184 14576 216 14608
rect 256 14576 288 14608
rect 328 14576 360 14608
rect 400 14576 432 14608
rect 472 14576 504 14608
rect 544 14576 576 14608
rect 616 14576 648 14608
rect 688 14576 720 14608
rect 760 14576 792 14608
rect 832 14576 864 14608
rect 904 14576 936 14608
rect 976 14576 1008 14608
rect 1048 14576 1080 14608
rect 1120 14576 1152 14608
rect 1192 14576 1224 14608
rect 1264 14576 1296 14608
rect 1336 14576 1368 14608
rect 1408 14576 1440 14608
rect 1480 14576 1512 14608
rect 1552 14576 1584 14608
rect 1624 14576 1656 14608
rect 1696 14576 1728 14608
rect 1768 14576 1800 14608
rect 1840 14576 1872 14608
rect 1912 14576 1944 14608
rect 1984 14576 2016 14608
rect 2056 14576 2088 14608
rect 2128 14576 2160 14608
rect 2200 14576 2232 14608
rect 2272 14576 2304 14608
rect 2344 14576 2376 14608
rect 2416 14576 2448 14608
rect 2488 14576 2520 14608
rect 2560 14576 2592 14608
rect 2632 14576 2664 14608
rect 2704 14576 2736 14608
rect 2776 14576 2808 14608
rect 2848 14576 2880 14608
rect 2920 14576 2952 14608
rect 2992 14576 3024 14608
rect 3064 14576 3096 14608
rect 3136 14576 3168 14608
rect 3208 14576 3240 14608
rect 3280 14576 3312 14608
rect 3352 14576 3384 14608
rect 3424 14576 3456 14608
rect 3496 14576 3528 14608
rect 3568 14576 3600 14608
rect 3640 14576 3672 14608
rect 3712 14576 3744 14608
rect 3784 14576 3816 14608
rect 3856 14576 3888 14608
rect 112 14504 144 14536
rect 184 14504 216 14536
rect 256 14504 288 14536
rect 328 14504 360 14536
rect 400 14504 432 14536
rect 472 14504 504 14536
rect 544 14504 576 14536
rect 616 14504 648 14536
rect 688 14504 720 14536
rect 760 14504 792 14536
rect 832 14504 864 14536
rect 904 14504 936 14536
rect 976 14504 1008 14536
rect 1048 14504 1080 14536
rect 1120 14504 1152 14536
rect 1192 14504 1224 14536
rect 1264 14504 1296 14536
rect 1336 14504 1368 14536
rect 1408 14504 1440 14536
rect 1480 14504 1512 14536
rect 1552 14504 1584 14536
rect 1624 14504 1656 14536
rect 1696 14504 1728 14536
rect 1768 14504 1800 14536
rect 1840 14504 1872 14536
rect 1912 14504 1944 14536
rect 1984 14504 2016 14536
rect 2056 14504 2088 14536
rect 2128 14504 2160 14536
rect 2200 14504 2232 14536
rect 2272 14504 2304 14536
rect 2344 14504 2376 14536
rect 2416 14504 2448 14536
rect 2488 14504 2520 14536
rect 2560 14504 2592 14536
rect 2632 14504 2664 14536
rect 2704 14504 2736 14536
rect 2776 14504 2808 14536
rect 2848 14504 2880 14536
rect 2920 14504 2952 14536
rect 2992 14504 3024 14536
rect 3064 14504 3096 14536
rect 3136 14504 3168 14536
rect 3208 14504 3240 14536
rect 3280 14504 3312 14536
rect 3352 14504 3384 14536
rect 3424 14504 3456 14536
rect 3496 14504 3528 14536
rect 3568 14504 3600 14536
rect 3640 14504 3672 14536
rect 3712 14504 3744 14536
rect 3784 14504 3816 14536
rect 3856 14504 3888 14536
rect 112 14432 144 14464
rect 184 14432 216 14464
rect 256 14432 288 14464
rect 328 14432 360 14464
rect 400 14432 432 14464
rect 472 14432 504 14464
rect 544 14432 576 14464
rect 616 14432 648 14464
rect 688 14432 720 14464
rect 760 14432 792 14464
rect 832 14432 864 14464
rect 904 14432 936 14464
rect 976 14432 1008 14464
rect 1048 14432 1080 14464
rect 1120 14432 1152 14464
rect 1192 14432 1224 14464
rect 1264 14432 1296 14464
rect 1336 14432 1368 14464
rect 1408 14432 1440 14464
rect 1480 14432 1512 14464
rect 1552 14432 1584 14464
rect 1624 14432 1656 14464
rect 1696 14432 1728 14464
rect 1768 14432 1800 14464
rect 1840 14432 1872 14464
rect 1912 14432 1944 14464
rect 1984 14432 2016 14464
rect 2056 14432 2088 14464
rect 2128 14432 2160 14464
rect 2200 14432 2232 14464
rect 2272 14432 2304 14464
rect 2344 14432 2376 14464
rect 2416 14432 2448 14464
rect 2488 14432 2520 14464
rect 2560 14432 2592 14464
rect 2632 14432 2664 14464
rect 2704 14432 2736 14464
rect 2776 14432 2808 14464
rect 2848 14432 2880 14464
rect 2920 14432 2952 14464
rect 2992 14432 3024 14464
rect 3064 14432 3096 14464
rect 3136 14432 3168 14464
rect 3208 14432 3240 14464
rect 3280 14432 3312 14464
rect 3352 14432 3384 14464
rect 3424 14432 3456 14464
rect 3496 14432 3528 14464
rect 3568 14432 3600 14464
rect 3640 14432 3672 14464
rect 3712 14432 3744 14464
rect 3784 14432 3816 14464
rect 3856 14432 3888 14464
rect 112 14360 144 14392
rect 184 14360 216 14392
rect 256 14360 288 14392
rect 328 14360 360 14392
rect 400 14360 432 14392
rect 472 14360 504 14392
rect 544 14360 576 14392
rect 616 14360 648 14392
rect 688 14360 720 14392
rect 760 14360 792 14392
rect 832 14360 864 14392
rect 904 14360 936 14392
rect 976 14360 1008 14392
rect 1048 14360 1080 14392
rect 1120 14360 1152 14392
rect 1192 14360 1224 14392
rect 1264 14360 1296 14392
rect 1336 14360 1368 14392
rect 1408 14360 1440 14392
rect 1480 14360 1512 14392
rect 1552 14360 1584 14392
rect 1624 14360 1656 14392
rect 1696 14360 1728 14392
rect 1768 14360 1800 14392
rect 1840 14360 1872 14392
rect 1912 14360 1944 14392
rect 1984 14360 2016 14392
rect 2056 14360 2088 14392
rect 2128 14360 2160 14392
rect 2200 14360 2232 14392
rect 2272 14360 2304 14392
rect 2344 14360 2376 14392
rect 2416 14360 2448 14392
rect 2488 14360 2520 14392
rect 2560 14360 2592 14392
rect 2632 14360 2664 14392
rect 2704 14360 2736 14392
rect 2776 14360 2808 14392
rect 2848 14360 2880 14392
rect 2920 14360 2952 14392
rect 2992 14360 3024 14392
rect 3064 14360 3096 14392
rect 3136 14360 3168 14392
rect 3208 14360 3240 14392
rect 3280 14360 3312 14392
rect 3352 14360 3384 14392
rect 3424 14360 3456 14392
rect 3496 14360 3528 14392
rect 3568 14360 3600 14392
rect 3640 14360 3672 14392
rect 3712 14360 3744 14392
rect 3784 14360 3816 14392
rect 3856 14360 3888 14392
rect 112 14288 144 14320
rect 184 14288 216 14320
rect 256 14288 288 14320
rect 328 14288 360 14320
rect 400 14288 432 14320
rect 472 14288 504 14320
rect 544 14288 576 14320
rect 616 14288 648 14320
rect 688 14288 720 14320
rect 760 14288 792 14320
rect 832 14288 864 14320
rect 904 14288 936 14320
rect 976 14288 1008 14320
rect 1048 14288 1080 14320
rect 1120 14288 1152 14320
rect 1192 14288 1224 14320
rect 1264 14288 1296 14320
rect 1336 14288 1368 14320
rect 1408 14288 1440 14320
rect 1480 14288 1512 14320
rect 1552 14288 1584 14320
rect 1624 14288 1656 14320
rect 1696 14288 1728 14320
rect 1768 14288 1800 14320
rect 1840 14288 1872 14320
rect 1912 14288 1944 14320
rect 1984 14288 2016 14320
rect 2056 14288 2088 14320
rect 2128 14288 2160 14320
rect 2200 14288 2232 14320
rect 2272 14288 2304 14320
rect 2344 14288 2376 14320
rect 2416 14288 2448 14320
rect 2488 14288 2520 14320
rect 2560 14288 2592 14320
rect 2632 14288 2664 14320
rect 2704 14288 2736 14320
rect 2776 14288 2808 14320
rect 2848 14288 2880 14320
rect 2920 14288 2952 14320
rect 2992 14288 3024 14320
rect 3064 14288 3096 14320
rect 3136 14288 3168 14320
rect 3208 14288 3240 14320
rect 3280 14288 3312 14320
rect 3352 14288 3384 14320
rect 3424 14288 3456 14320
rect 3496 14288 3528 14320
rect 3568 14288 3600 14320
rect 3640 14288 3672 14320
rect 3712 14288 3744 14320
rect 3784 14288 3816 14320
rect 3856 14288 3888 14320
rect 112 14216 144 14248
rect 184 14216 216 14248
rect 256 14216 288 14248
rect 328 14216 360 14248
rect 400 14216 432 14248
rect 472 14216 504 14248
rect 544 14216 576 14248
rect 616 14216 648 14248
rect 688 14216 720 14248
rect 760 14216 792 14248
rect 832 14216 864 14248
rect 904 14216 936 14248
rect 976 14216 1008 14248
rect 1048 14216 1080 14248
rect 1120 14216 1152 14248
rect 1192 14216 1224 14248
rect 1264 14216 1296 14248
rect 1336 14216 1368 14248
rect 1408 14216 1440 14248
rect 1480 14216 1512 14248
rect 1552 14216 1584 14248
rect 1624 14216 1656 14248
rect 1696 14216 1728 14248
rect 1768 14216 1800 14248
rect 1840 14216 1872 14248
rect 1912 14216 1944 14248
rect 1984 14216 2016 14248
rect 2056 14216 2088 14248
rect 2128 14216 2160 14248
rect 2200 14216 2232 14248
rect 2272 14216 2304 14248
rect 2344 14216 2376 14248
rect 2416 14216 2448 14248
rect 2488 14216 2520 14248
rect 2560 14216 2592 14248
rect 2632 14216 2664 14248
rect 2704 14216 2736 14248
rect 2776 14216 2808 14248
rect 2848 14216 2880 14248
rect 2920 14216 2952 14248
rect 2992 14216 3024 14248
rect 3064 14216 3096 14248
rect 3136 14216 3168 14248
rect 3208 14216 3240 14248
rect 3280 14216 3312 14248
rect 3352 14216 3384 14248
rect 3424 14216 3456 14248
rect 3496 14216 3528 14248
rect 3568 14216 3600 14248
rect 3640 14216 3672 14248
rect 3712 14216 3744 14248
rect 3784 14216 3816 14248
rect 3856 14216 3888 14248
rect 112 14144 144 14176
rect 184 14144 216 14176
rect 256 14144 288 14176
rect 328 14144 360 14176
rect 400 14144 432 14176
rect 472 14144 504 14176
rect 544 14144 576 14176
rect 616 14144 648 14176
rect 688 14144 720 14176
rect 760 14144 792 14176
rect 832 14144 864 14176
rect 904 14144 936 14176
rect 976 14144 1008 14176
rect 1048 14144 1080 14176
rect 1120 14144 1152 14176
rect 1192 14144 1224 14176
rect 1264 14144 1296 14176
rect 1336 14144 1368 14176
rect 1408 14144 1440 14176
rect 1480 14144 1512 14176
rect 1552 14144 1584 14176
rect 1624 14144 1656 14176
rect 1696 14144 1728 14176
rect 1768 14144 1800 14176
rect 1840 14144 1872 14176
rect 1912 14144 1944 14176
rect 1984 14144 2016 14176
rect 2056 14144 2088 14176
rect 2128 14144 2160 14176
rect 2200 14144 2232 14176
rect 2272 14144 2304 14176
rect 2344 14144 2376 14176
rect 2416 14144 2448 14176
rect 2488 14144 2520 14176
rect 2560 14144 2592 14176
rect 2632 14144 2664 14176
rect 2704 14144 2736 14176
rect 2776 14144 2808 14176
rect 2848 14144 2880 14176
rect 2920 14144 2952 14176
rect 2992 14144 3024 14176
rect 3064 14144 3096 14176
rect 3136 14144 3168 14176
rect 3208 14144 3240 14176
rect 3280 14144 3312 14176
rect 3352 14144 3384 14176
rect 3424 14144 3456 14176
rect 3496 14144 3528 14176
rect 3568 14144 3600 14176
rect 3640 14144 3672 14176
rect 3712 14144 3744 14176
rect 3784 14144 3816 14176
rect 3856 14144 3888 14176
rect 112 14072 144 14104
rect 184 14072 216 14104
rect 256 14072 288 14104
rect 328 14072 360 14104
rect 400 14072 432 14104
rect 472 14072 504 14104
rect 544 14072 576 14104
rect 616 14072 648 14104
rect 688 14072 720 14104
rect 760 14072 792 14104
rect 832 14072 864 14104
rect 904 14072 936 14104
rect 976 14072 1008 14104
rect 1048 14072 1080 14104
rect 1120 14072 1152 14104
rect 1192 14072 1224 14104
rect 1264 14072 1296 14104
rect 1336 14072 1368 14104
rect 1408 14072 1440 14104
rect 1480 14072 1512 14104
rect 1552 14072 1584 14104
rect 1624 14072 1656 14104
rect 1696 14072 1728 14104
rect 1768 14072 1800 14104
rect 1840 14072 1872 14104
rect 1912 14072 1944 14104
rect 1984 14072 2016 14104
rect 2056 14072 2088 14104
rect 2128 14072 2160 14104
rect 2200 14072 2232 14104
rect 2272 14072 2304 14104
rect 2344 14072 2376 14104
rect 2416 14072 2448 14104
rect 2488 14072 2520 14104
rect 2560 14072 2592 14104
rect 2632 14072 2664 14104
rect 2704 14072 2736 14104
rect 2776 14072 2808 14104
rect 2848 14072 2880 14104
rect 2920 14072 2952 14104
rect 2992 14072 3024 14104
rect 3064 14072 3096 14104
rect 3136 14072 3168 14104
rect 3208 14072 3240 14104
rect 3280 14072 3312 14104
rect 3352 14072 3384 14104
rect 3424 14072 3456 14104
rect 3496 14072 3528 14104
rect 3568 14072 3600 14104
rect 3640 14072 3672 14104
rect 3712 14072 3744 14104
rect 3784 14072 3816 14104
rect 3856 14072 3888 14104
rect 112 14000 144 14032
rect 184 14000 216 14032
rect 256 14000 288 14032
rect 328 14000 360 14032
rect 400 14000 432 14032
rect 472 14000 504 14032
rect 544 14000 576 14032
rect 616 14000 648 14032
rect 688 14000 720 14032
rect 760 14000 792 14032
rect 832 14000 864 14032
rect 904 14000 936 14032
rect 976 14000 1008 14032
rect 1048 14000 1080 14032
rect 1120 14000 1152 14032
rect 1192 14000 1224 14032
rect 1264 14000 1296 14032
rect 1336 14000 1368 14032
rect 1408 14000 1440 14032
rect 1480 14000 1512 14032
rect 1552 14000 1584 14032
rect 1624 14000 1656 14032
rect 1696 14000 1728 14032
rect 1768 14000 1800 14032
rect 1840 14000 1872 14032
rect 1912 14000 1944 14032
rect 1984 14000 2016 14032
rect 2056 14000 2088 14032
rect 2128 14000 2160 14032
rect 2200 14000 2232 14032
rect 2272 14000 2304 14032
rect 2344 14000 2376 14032
rect 2416 14000 2448 14032
rect 2488 14000 2520 14032
rect 2560 14000 2592 14032
rect 2632 14000 2664 14032
rect 2704 14000 2736 14032
rect 2776 14000 2808 14032
rect 2848 14000 2880 14032
rect 2920 14000 2952 14032
rect 2992 14000 3024 14032
rect 3064 14000 3096 14032
rect 3136 14000 3168 14032
rect 3208 14000 3240 14032
rect 3280 14000 3312 14032
rect 3352 14000 3384 14032
rect 3424 14000 3456 14032
rect 3496 14000 3528 14032
rect 3568 14000 3600 14032
rect 3640 14000 3672 14032
rect 3712 14000 3744 14032
rect 3784 14000 3816 14032
rect 3856 14000 3888 14032
rect 112 13928 144 13960
rect 184 13928 216 13960
rect 256 13928 288 13960
rect 328 13928 360 13960
rect 400 13928 432 13960
rect 472 13928 504 13960
rect 544 13928 576 13960
rect 616 13928 648 13960
rect 688 13928 720 13960
rect 760 13928 792 13960
rect 832 13928 864 13960
rect 904 13928 936 13960
rect 976 13928 1008 13960
rect 1048 13928 1080 13960
rect 1120 13928 1152 13960
rect 1192 13928 1224 13960
rect 1264 13928 1296 13960
rect 1336 13928 1368 13960
rect 1408 13928 1440 13960
rect 1480 13928 1512 13960
rect 1552 13928 1584 13960
rect 1624 13928 1656 13960
rect 1696 13928 1728 13960
rect 1768 13928 1800 13960
rect 1840 13928 1872 13960
rect 1912 13928 1944 13960
rect 1984 13928 2016 13960
rect 2056 13928 2088 13960
rect 2128 13928 2160 13960
rect 2200 13928 2232 13960
rect 2272 13928 2304 13960
rect 2344 13928 2376 13960
rect 2416 13928 2448 13960
rect 2488 13928 2520 13960
rect 2560 13928 2592 13960
rect 2632 13928 2664 13960
rect 2704 13928 2736 13960
rect 2776 13928 2808 13960
rect 2848 13928 2880 13960
rect 2920 13928 2952 13960
rect 2992 13928 3024 13960
rect 3064 13928 3096 13960
rect 3136 13928 3168 13960
rect 3208 13928 3240 13960
rect 3280 13928 3312 13960
rect 3352 13928 3384 13960
rect 3424 13928 3456 13960
rect 3496 13928 3528 13960
rect 3568 13928 3600 13960
rect 3640 13928 3672 13960
rect 3712 13928 3744 13960
rect 3784 13928 3816 13960
rect 3856 13928 3888 13960
rect 112 13856 144 13888
rect 184 13856 216 13888
rect 256 13856 288 13888
rect 328 13856 360 13888
rect 400 13856 432 13888
rect 472 13856 504 13888
rect 544 13856 576 13888
rect 616 13856 648 13888
rect 688 13856 720 13888
rect 760 13856 792 13888
rect 832 13856 864 13888
rect 904 13856 936 13888
rect 976 13856 1008 13888
rect 1048 13856 1080 13888
rect 1120 13856 1152 13888
rect 1192 13856 1224 13888
rect 1264 13856 1296 13888
rect 1336 13856 1368 13888
rect 1408 13856 1440 13888
rect 1480 13856 1512 13888
rect 1552 13856 1584 13888
rect 1624 13856 1656 13888
rect 1696 13856 1728 13888
rect 1768 13856 1800 13888
rect 1840 13856 1872 13888
rect 1912 13856 1944 13888
rect 1984 13856 2016 13888
rect 2056 13856 2088 13888
rect 2128 13856 2160 13888
rect 2200 13856 2232 13888
rect 2272 13856 2304 13888
rect 2344 13856 2376 13888
rect 2416 13856 2448 13888
rect 2488 13856 2520 13888
rect 2560 13856 2592 13888
rect 2632 13856 2664 13888
rect 2704 13856 2736 13888
rect 2776 13856 2808 13888
rect 2848 13856 2880 13888
rect 2920 13856 2952 13888
rect 2992 13856 3024 13888
rect 3064 13856 3096 13888
rect 3136 13856 3168 13888
rect 3208 13856 3240 13888
rect 3280 13856 3312 13888
rect 3352 13856 3384 13888
rect 3424 13856 3456 13888
rect 3496 13856 3528 13888
rect 3568 13856 3600 13888
rect 3640 13856 3672 13888
rect 3712 13856 3744 13888
rect 3784 13856 3816 13888
rect 3856 13856 3888 13888
rect 112 13784 144 13816
rect 184 13784 216 13816
rect 256 13784 288 13816
rect 328 13784 360 13816
rect 400 13784 432 13816
rect 472 13784 504 13816
rect 544 13784 576 13816
rect 616 13784 648 13816
rect 688 13784 720 13816
rect 760 13784 792 13816
rect 832 13784 864 13816
rect 904 13784 936 13816
rect 976 13784 1008 13816
rect 1048 13784 1080 13816
rect 1120 13784 1152 13816
rect 1192 13784 1224 13816
rect 1264 13784 1296 13816
rect 1336 13784 1368 13816
rect 1408 13784 1440 13816
rect 1480 13784 1512 13816
rect 1552 13784 1584 13816
rect 1624 13784 1656 13816
rect 1696 13784 1728 13816
rect 1768 13784 1800 13816
rect 1840 13784 1872 13816
rect 1912 13784 1944 13816
rect 1984 13784 2016 13816
rect 2056 13784 2088 13816
rect 2128 13784 2160 13816
rect 2200 13784 2232 13816
rect 2272 13784 2304 13816
rect 2344 13784 2376 13816
rect 2416 13784 2448 13816
rect 2488 13784 2520 13816
rect 2560 13784 2592 13816
rect 2632 13784 2664 13816
rect 2704 13784 2736 13816
rect 2776 13784 2808 13816
rect 2848 13784 2880 13816
rect 2920 13784 2952 13816
rect 2992 13784 3024 13816
rect 3064 13784 3096 13816
rect 3136 13784 3168 13816
rect 3208 13784 3240 13816
rect 3280 13784 3312 13816
rect 3352 13784 3384 13816
rect 3424 13784 3456 13816
rect 3496 13784 3528 13816
rect 3568 13784 3600 13816
rect 3640 13784 3672 13816
rect 3712 13784 3744 13816
rect 3784 13784 3816 13816
rect 3856 13784 3888 13816
rect 112 13712 144 13744
rect 184 13712 216 13744
rect 256 13712 288 13744
rect 328 13712 360 13744
rect 400 13712 432 13744
rect 472 13712 504 13744
rect 544 13712 576 13744
rect 616 13712 648 13744
rect 688 13712 720 13744
rect 760 13712 792 13744
rect 832 13712 864 13744
rect 904 13712 936 13744
rect 976 13712 1008 13744
rect 1048 13712 1080 13744
rect 1120 13712 1152 13744
rect 1192 13712 1224 13744
rect 1264 13712 1296 13744
rect 1336 13712 1368 13744
rect 1408 13712 1440 13744
rect 1480 13712 1512 13744
rect 1552 13712 1584 13744
rect 1624 13712 1656 13744
rect 1696 13712 1728 13744
rect 1768 13712 1800 13744
rect 1840 13712 1872 13744
rect 1912 13712 1944 13744
rect 1984 13712 2016 13744
rect 2056 13712 2088 13744
rect 2128 13712 2160 13744
rect 2200 13712 2232 13744
rect 2272 13712 2304 13744
rect 2344 13712 2376 13744
rect 2416 13712 2448 13744
rect 2488 13712 2520 13744
rect 2560 13712 2592 13744
rect 2632 13712 2664 13744
rect 2704 13712 2736 13744
rect 2776 13712 2808 13744
rect 2848 13712 2880 13744
rect 2920 13712 2952 13744
rect 2992 13712 3024 13744
rect 3064 13712 3096 13744
rect 3136 13712 3168 13744
rect 3208 13712 3240 13744
rect 3280 13712 3312 13744
rect 3352 13712 3384 13744
rect 3424 13712 3456 13744
rect 3496 13712 3528 13744
rect 3568 13712 3600 13744
rect 3640 13712 3672 13744
rect 3712 13712 3744 13744
rect 3784 13712 3816 13744
rect 3856 13712 3888 13744
rect 112 13640 144 13672
rect 184 13640 216 13672
rect 256 13640 288 13672
rect 328 13640 360 13672
rect 400 13640 432 13672
rect 472 13640 504 13672
rect 544 13640 576 13672
rect 616 13640 648 13672
rect 688 13640 720 13672
rect 760 13640 792 13672
rect 832 13640 864 13672
rect 904 13640 936 13672
rect 976 13640 1008 13672
rect 1048 13640 1080 13672
rect 1120 13640 1152 13672
rect 1192 13640 1224 13672
rect 1264 13640 1296 13672
rect 1336 13640 1368 13672
rect 1408 13640 1440 13672
rect 1480 13640 1512 13672
rect 1552 13640 1584 13672
rect 1624 13640 1656 13672
rect 1696 13640 1728 13672
rect 1768 13640 1800 13672
rect 1840 13640 1872 13672
rect 1912 13640 1944 13672
rect 1984 13640 2016 13672
rect 2056 13640 2088 13672
rect 2128 13640 2160 13672
rect 2200 13640 2232 13672
rect 2272 13640 2304 13672
rect 2344 13640 2376 13672
rect 2416 13640 2448 13672
rect 2488 13640 2520 13672
rect 2560 13640 2592 13672
rect 2632 13640 2664 13672
rect 2704 13640 2736 13672
rect 2776 13640 2808 13672
rect 2848 13640 2880 13672
rect 2920 13640 2952 13672
rect 2992 13640 3024 13672
rect 3064 13640 3096 13672
rect 3136 13640 3168 13672
rect 3208 13640 3240 13672
rect 3280 13640 3312 13672
rect 3352 13640 3384 13672
rect 3424 13640 3456 13672
rect 3496 13640 3528 13672
rect 3568 13640 3600 13672
rect 3640 13640 3672 13672
rect 3712 13640 3744 13672
rect 3784 13640 3816 13672
rect 3856 13640 3888 13672
rect 112 13568 144 13600
rect 184 13568 216 13600
rect 256 13568 288 13600
rect 328 13568 360 13600
rect 400 13568 432 13600
rect 472 13568 504 13600
rect 544 13568 576 13600
rect 616 13568 648 13600
rect 688 13568 720 13600
rect 760 13568 792 13600
rect 832 13568 864 13600
rect 904 13568 936 13600
rect 976 13568 1008 13600
rect 1048 13568 1080 13600
rect 1120 13568 1152 13600
rect 1192 13568 1224 13600
rect 1264 13568 1296 13600
rect 1336 13568 1368 13600
rect 1408 13568 1440 13600
rect 1480 13568 1512 13600
rect 1552 13568 1584 13600
rect 1624 13568 1656 13600
rect 1696 13568 1728 13600
rect 1768 13568 1800 13600
rect 1840 13568 1872 13600
rect 1912 13568 1944 13600
rect 1984 13568 2016 13600
rect 2056 13568 2088 13600
rect 2128 13568 2160 13600
rect 2200 13568 2232 13600
rect 2272 13568 2304 13600
rect 2344 13568 2376 13600
rect 2416 13568 2448 13600
rect 2488 13568 2520 13600
rect 2560 13568 2592 13600
rect 2632 13568 2664 13600
rect 2704 13568 2736 13600
rect 2776 13568 2808 13600
rect 2848 13568 2880 13600
rect 2920 13568 2952 13600
rect 2992 13568 3024 13600
rect 3064 13568 3096 13600
rect 3136 13568 3168 13600
rect 3208 13568 3240 13600
rect 3280 13568 3312 13600
rect 3352 13568 3384 13600
rect 3424 13568 3456 13600
rect 3496 13568 3528 13600
rect 3568 13568 3600 13600
rect 3640 13568 3672 13600
rect 3712 13568 3744 13600
rect 3784 13568 3816 13600
rect 3856 13568 3888 13600
rect 112 13496 144 13528
rect 184 13496 216 13528
rect 256 13496 288 13528
rect 328 13496 360 13528
rect 400 13496 432 13528
rect 472 13496 504 13528
rect 544 13496 576 13528
rect 616 13496 648 13528
rect 688 13496 720 13528
rect 760 13496 792 13528
rect 832 13496 864 13528
rect 904 13496 936 13528
rect 976 13496 1008 13528
rect 1048 13496 1080 13528
rect 1120 13496 1152 13528
rect 1192 13496 1224 13528
rect 1264 13496 1296 13528
rect 1336 13496 1368 13528
rect 1408 13496 1440 13528
rect 1480 13496 1512 13528
rect 1552 13496 1584 13528
rect 1624 13496 1656 13528
rect 1696 13496 1728 13528
rect 1768 13496 1800 13528
rect 1840 13496 1872 13528
rect 1912 13496 1944 13528
rect 1984 13496 2016 13528
rect 2056 13496 2088 13528
rect 2128 13496 2160 13528
rect 2200 13496 2232 13528
rect 2272 13496 2304 13528
rect 2344 13496 2376 13528
rect 2416 13496 2448 13528
rect 2488 13496 2520 13528
rect 2560 13496 2592 13528
rect 2632 13496 2664 13528
rect 2704 13496 2736 13528
rect 2776 13496 2808 13528
rect 2848 13496 2880 13528
rect 2920 13496 2952 13528
rect 2992 13496 3024 13528
rect 3064 13496 3096 13528
rect 3136 13496 3168 13528
rect 3208 13496 3240 13528
rect 3280 13496 3312 13528
rect 3352 13496 3384 13528
rect 3424 13496 3456 13528
rect 3496 13496 3528 13528
rect 3568 13496 3600 13528
rect 3640 13496 3672 13528
rect 3712 13496 3744 13528
rect 3784 13496 3816 13528
rect 3856 13496 3888 13528
rect 112 13424 144 13456
rect 184 13424 216 13456
rect 256 13424 288 13456
rect 328 13424 360 13456
rect 400 13424 432 13456
rect 472 13424 504 13456
rect 544 13424 576 13456
rect 616 13424 648 13456
rect 688 13424 720 13456
rect 760 13424 792 13456
rect 832 13424 864 13456
rect 904 13424 936 13456
rect 976 13424 1008 13456
rect 1048 13424 1080 13456
rect 1120 13424 1152 13456
rect 1192 13424 1224 13456
rect 1264 13424 1296 13456
rect 1336 13424 1368 13456
rect 1408 13424 1440 13456
rect 1480 13424 1512 13456
rect 1552 13424 1584 13456
rect 1624 13424 1656 13456
rect 1696 13424 1728 13456
rect 1768 13424 1800 13456
rect 1840 13424 1872 13456
rect 1912 13424 1944 13456
rect 1984 13424 2016 13456
rect 2056 13424 2088 13456
rect 2128 13424 2160 13456
rect 2200 13424 2232 13456
rect 2272 13424 2304 13456
rect 2344 13424 2376 13456
rect 2416 13424 2448 13456
rect 2488 13424 2520 13456
rect 2560 13424 2592 13456
rect 2632 13424 2664 13456
rect 2704 13424 2736 13456
rect 2776 13424 2808 13456
rect 2848 13424 2880 13456
rect 2920 13424 2952 13456
rect 2992 13424 3024 13456
rect 3064 13424 3096 13456
rect 3136 13424 3168 13456
rect 3208 13424 3240 13456
rect 3280 13424 3312 13456
rect 3352 13424 3384 13456
rect 3424 13424 3456 13456
rect 3496 13424 3528 13456
rect 3568 13424 3600 13456
rect 3640 13424 3672 13456
rect 3712 13424 3744 13456
rect 3784 13424 3816 13456
rect 3856 13424 3888 13456
rect 112 13352 144 13384
rect 184 13352 216 13384
rect 256 13352 288 13384
rect 328 13352 360 13384
rect 400 13352 432 13384
rect 472 13352 504 13384
rect 544 13352 576 13384
rect 616 13352 648 13384
rect 688 13352 720 13384
rect 760 13352 792 13384
rect 832 13352 864 13384
rect 904 13352 936 13384
rect 976 13352 1008 13384
rect 1048 13352 1080 13384
rect 1120 13352 1152 13384
rect 1192 13352 1224 13384
rect 1264 13352 1296 13384
rect 1336 13352 1368 13384
rect 1408 13352 1440 13384
rect 1480 13352 1512 13384
rect 1552 13352 1584 13384
rect 1624 13352 1656 13384
rect 1696 13352 1728 13384
rect 1768 13352 1800 13384
rect 1840 13352 1872 13384
rect 1912 13352 1944 13384
rect 1984 13352 2016 13384
rect 2056 13352 2088 13384
rect 2128 13352 2160 13384
rect 2200 13352 2232 13384
rect 2272 13352 2304 13384
rect 2344 13352 2376 13384
rect 2416 13352 2448 13384
rect 2488 13352 2520 13384
rect 2560 13352 2592 13384
rect 2632 13352 2664 13384
rect 2704 13352 2736 13384
rect 2776 13352 2808 13384
rect 2848 13352 2880 13384
rect 2920 13352 2952 13384
rect 2992 13352 3024 13384
rect 3064 13352 3096 13384
rect 3136 13352 3168 13384
rect 3208 13352 3240 13384
rect 3280 13352 3312 13384
rect 3352 13352 3384 13384
rect 3424 13352 3456 13384
rect 3496 13352 3528 13384
rect 3568 13352 3600 13384
rect 3640 13352 3672 13384
rect 3712 13352 3744 13384
rect 3784 13352 3816 13384
rect 3856 13352 3888 13384
rect 112 13280 144 13312
rect 184 13280 216 13312
rect 256 13280 288 13312
rect 328 13280 360 13312
rect 400 13280 432 13312
rect 472 13280 504 13312
rect 544 13280 576 13312
rect 616 13280 648 13312
rect 688 13280 720 13312
rect 760 13280 792 13312
rect 832 13280 864 13312
rect 904 13280 936 13312
rect 976 13280 1008 13312
rect 1048 13280 1080 13312
rect 1120 13280 1152 13312
rect 1192 13280 1224 13312
rect 1264 13280 1296 13312
rect 1336 13280 1368 13312
rect 1408 13280 1440 13312
rect 1480 13280 1512 13312
rect 1552 13280 1584 13312
rect 1624 13280 1656 13312
rect 1696 13280 1728 13312
rect 1768 13280 1800 13312
rect 1840 13280 1872 13312
rect 1912 13280 1944 13312
rect 1984 13280 2016 13312
rect 2056 13280 2088 13312
rect 2128 13280 2160 13312
rect 2200 13280 2232 13312
rect 2272 13280 2304 13312
rect 2344 13280 2376 13312
rect 2416 13280 2448 13312
rect 2488 13280 2520 13312
rect 2560 13280 2592 13312
rect 2632 13280 2664 13312
rect 2704 13280 2736 13312
rect 2776 13280 2808 13312
rect 2848 13280 2880 13312
rect 2920 13280 2952 13312
rect 2992 13280 3024 13312
rect 3064 13280 3096 13312
rect 3136 13280 3168 13312
rect 3208 13280 3240 13312
rect 3280 13280 3312 13312
rect 3352 13280 3384 13312
rect 3424 13280 3456 13312
rect 3496 13280 3528 13312
rect 3568 13280 3600 13312
rect 3640 13280 3672 13312
rect 3712 13280 3744 13312
rect 3784 13280 3816 13312
rect 3856 13280 3888 13312
rect 112 13208 144 13240
rect 184 13208 216 13240
rect 256 13208 288 13240
rect 328 13208 360 13240
rect 400 13208 432 13240
rect 472 13208 504 13240
rect 544 13208 576 13240
rect 616 13208 648 13240
rect 688 13208 720 13240
rect 760 13208 792 13240
rect 832 13208 864 13240
rect 904 13208 936 13240
rect 976 13208 1008 13240
rect 1048 13208 1080 13240
rect 1120 13208 1152 13240
rect 1192 13208 1224 13240
rect 1264 13208 1296 13240
rect 1336 13208 1368 13240
rect 1408 13208 1440 13240
rect 1480 13208 1512 13240
rect 1552 13208 1584 13240
rect 1624 13208 1656 13240
rect 1696 13208 1728 13240
rect 1768 13208 1800 13240
rect 1840 13208 1872 13240
rect 1912 13208 1944 13240
rect 1984 13208 2016 13240
rect 2056 13208 2088 13240
rect 2128 13208 2160 13240
rect 2200 13208 2232 13240
rect 2272 13208 2304 13240
rect 2344 13208 2376 13240
rect 2416 13208 2448 13240
rect 2488 13208 2520 13240
rect 2560 13208 2592 13240
rect 2632 13208 2664 13240
rect 2704 13208 2736 13240
rect 2776 13208 2808 13240
rect 2848 13208 2880 13240
rect 2920 13208 2952 13240
rect 2992 13208 3024 13240
rect 3064 13208 3096 13240
rect 3136 13208 3168 13240
rect 3208 13208 3240 13240
rect 3280 13208 3312 13240
rect 3352 13208 3384 13240
rect 3424 13208 3456 13240
rect 3496 13208 3528 13240
rect 3568 13208 3600 13240
rect 3640 13208 3672 13240
rect 3712 13208 3744 13240
rect 3784 13208 3816 13240
rect 3856 13208 3888 13240
rect 112 13136 144 13168
rect 184 13136 216 13168
rect 256 13136 288 13168
rect 328 13136 360 13168
rect 400 13136 432 13168
rect 472 13136 504 13168
rect 544 13136 576 13168
rect 616 13136 648 13168
rect 688 13136 720 13168
rect 760 13136 792 13168
rect 832 13136 864 13168
rect 904 13136 936 13168
rect 976 13136 1008 13168
rect 1048 13136 1080 13168
rect 1120 13136 1152 13168
rect 1192 13136 1224 13168
rect 1264 13136 1296 13168
rect 1336 13136 1368 13168
rect 1408 13136 1440 13168
rect 1480 13136 1512 13168
rect 1552 13136 1584 13168
rect 1624 13136 1656 13168
rect 1696 13136 1728 13168
rect 1768 13136 1800 13168
rect 1840 13136 1872 13168
rect 1912 13136 1944 13168
rect 1984 13136 2016 13168
rect 2056 13136 2088 13168
rect 2128 13136 2160 13168
rect 2200 13136 2232 13168
rect 2272 13136 2304 13168
rect 2344 13136 2376 13168
rect 2416 13136 2448 13168
rect 2488 13136 2520 13168
rect 2560 13136 2592 13168
rect 2632 13136 2664 13168
rect 2704 13136 2736 13168
rect 2776 13136 2808 13168
rect 2848 13136 2880 13168
rect 2920 13136 2952 13168
rect 2992 13136 3024 13168
rect 3064 13136 3096 13168
rect 3136 13136 3168 13168
rect 3208 13136 3240 13168
rect 3280 13136 3312 13168
rect 3352 13136 3384 13168
rect 3424 13136 3456 13168
rect 3496 13136 3528 13168
rect 3568 13136 3600 13168
rect 3640 13136 3672 13168
rect 3712 13136 3744 13168
rect 3784 13136 3816 13168
rect 3856 13136 3888 13168
rect 112 13064 144 13096
rect 184 13064 216 13096
rect 256 13064 288 13096
rect 328 13064 360 13096
rect 400 13064 432 13096
rect 472 13064 504 13096
rect 544 13064 576 13096
rect 616 13064 648 13096
rect 688 13064 720 13096
rect 760 13064 792 13096
rect 832 13064 864 13096
rect 904 13064 936 13096
rect 976 13064 1008 13096
rect 1048 13064 1080 13096
rect 1120 13064 1152 13096
rect 1192 13064 1224 13096
rect 1264 13064 1296 13096
rect 1336 13064 1368 13096
rect 1408 13064 1440 13096
rect 1480 13064 1512 13096
rect 1552 13064 1584 13096
rect 1624 13064 1656 13096
rect 1696 13064 1728 13096
rect 1768 13064 1800 13096
rect 1840 13064 1872 13096
rect 1912 13064 1944 13096
rect 1984 13064 2016 13096
rect 2056 13064 2088 13096
rect 2128 13064 2160 13096
rect 2200 13064 2232 13096
rect 2272 13064 2304 13096
rect 2344 13064 2376 13096
rect 2416 13064 2448 13096
rect 2488 13064 2520 13096
rect 2560 13064 2592 13096
rect 2632 13064 2664 13096
rect 2704 13064 2736 13096
rect 2776 13064 2808 13096
rect 2848 13064 2880 13096
rect 2920 13064 2952 13096
rect 2992 13064 3024 13096
rect 3064 13064 3096 13096
rect 3136 13064 3168 13096
rect 3208 13064 3240 13096
rect 3280 13064 3312 13096
rect 3352 13064 3384 13096
rect 3424 13064 3456 13096
rect 3496 13064 3528 13096
rect 3568 13064 3600 13096
rect 3640 13064 3672 13096
rect 3712 13064 3744 13096
rect 3784 13064 3816 13096
rect 3856 13064 3888 13096
rect 50 31416 3950 31430
rect 50 31384 112 31416
rect 144 31384 184 31416
rect 216 31384 256 31416
rect 288 31384 328 31416
rect 360 31384 400 31416
rect 432 31384 472 31416
rect 504 31384 544 31416
rect 576 31384 616 31416
rect 648 31384 688 31416
rect 720 31384 760 31416
rect 792 31384 832 31416
rect 864 31384 904 31416
rect 936 31384 976 31416
rect 1008 31384 1048 31416
rect 1080 31384 1120 31416
rect 1152 31384 1192 31416
rect 1224 31384 1264 31416
rect 1296 31384 1336 31416
rect 1368 31384 1408 31416
rect 1440 31384 1480 31416
rect 1512 31384 1552 31416
rect 1584 31384 1624 31416
rect 1656 31384 1696 31416
rect 1728 31384 1768 31416
rect 1800 31384 1840 31416
rect 1872 31384 1912 31416
rect 1944 31384 1984 31416
rect 2016 31384 2056 31416
rect 2088 31384 2128 31416
rect 2160 31384 2200 31416
rect 2232 31384 2272 31416
rect 2304 31384 2344 31416
rect 2376 31384 2416 31416
rect 2448 31384 2488 31416
rect 2520 31384 2560 31416
rect 2592 31384 2632 31416
rect 2664 31384 2704 31416
rect 2736 31384 2776 31416
rect 2808 31384 2848 31416
rect 2880 31384 2920 31416
rect 2952 31384 2992 31416
rect 3024 31384 3064 31416
rect 3096 31384 3136 31416
rect 3168 31384 3208 31416
rect 3240 31384 3280 31416
rect 3312 31384 3352 31416
rect 3384 31384 3424 31416
rect 3456 31384 3496 31416
rect 3528 31384 3568 31416
rect 3600 31384 3640 31416
rect 3672 31384 3712 31416
rect 3744 31384 3784 31416
rect 3816 31384 3856 31416
rect 3888 31384 3950 31416
rect 50 31370 3950 31384
rect 50 27971 3950 28034
rect 50 27939 112 27971
rect 144 27939 184 27971
rect 216 27939 256 27971
rect 288 27939 328 27971
rect 360 27939 400 27971
rect 432 27939 472 27971
rect 504 27939 544 27971
rect 576 27939 616 27971
rect 648 27939 688 27971
rect 720 27939 760 27971
rect 792 27939 832 27971
rect 864 27939 904 27971
rect 936 27939 976 27971
rect 1008 27939 1048 27971
rect 1080 27939 1120 27971
rect 1152 27939 1192 27971
rect 1224 27939 1264 27971
rect 1296 27939 1336 27971
rect 1368 27939 1408 27971
rect 1440 27939 1480 27971
rect 1512 27939 1552 27971
rect 1584 27939 1624 27971
rect 1656 27939 1696 27971
rect 1728 27939 1768 27971
rect 1800 27939 1840 27971
rect 1872 27939 1912 27971
rect 1944 27939 1984 27971
rect 2016 27939 2056 27971
rect 2088 27939 2128 27971
rect 2160 27939 2200 27971
rect 2232 27939 2272 27971
rect 2304 27939 2344 27971
rect 2376 27939 2416 27971
rect 2448 27939 2488 27971
rect 2520 27939 2560 27971
rect 2592 27939 2632 27971
rect 2664 27939 2704 27971
rect 2736 27939 2776 27971
rect 2808 27939 2848 27971
rect 2880 27939 2920 27971
rect 2952 27939 2992 27971
rect 3024 27939 3064 27971
rect 3096 27939 3136 27971
rect 3168 27939 3208 27971
rect 3240 27939 3280 27971
rect 3312 27939 3352 27971
rect 3384 27939 3424 27971
rect 3456 27939 3496 27971
rect 3528 27939 3568 27971
rect 3600 27939 3640 27971
rect 3672 27939 3712 27971
rect 3744 27939 3784 27971
rect 3816 27939 3856 27971
rect 3888 27939 3950 27971
rect 50 27899 3950 27939
rect 50 27867 112 27899
rect 144 27867 184 27899
rect 216 27867 256 27899
rect 288 27867 328 27899
rect 360 27867 400 27899
rect 432 27867 472 27899
rect 504 27867 544 27899
rect 576 27867 616 27899
rect 648 27867 688 27899
rect 720 27867 760 27899
rect 792 27867 832 27899
rect 864 27867 904 27899
rect 936 27867 976 27899
rect 1008 27867 1048 27899
rect 1080 27867 1120 27899
rect 1152 27867 1192 27899
rect 1224 27867 1264 27899
rect 1296 27867 1336 27899
rect 1368 27867 1408 27899
rect 1440 27867 1480 27899
rect 1512 27867 1552 27899
rect 1584 27867 1624 27899
rect 1656 27867 1696 27899
rect 1728 27867 1768 27899
rect 1800 27867 1840 27899
rect 1872 27867 1912 27899
rect 1944 27867 1984 27899
rect 2016 27867 2056 27899
rect 2088 27867 2128 27899
rect 2160 27867 2200 27899
rect 2232 27867 2272 27899
rect 2304 27867 2344 27899
rect 2376 27867 2416 27899
rect 2448 27867 2488 27899
rect 2520 27867 2560 27899
rect 2592 27867 2632 27899
rect 2664 27867 2704 27899
rect 2736 27867 2776 27899
rect 2808 27867 2848 27899
rect 2880 27867 2920 27899
rect 2952 27867 2992 27899
rect 3024 27867 3064 27899
rect 3096 27867 3136 27899
rect 3168 27867 3208 27899
rect 3240 27867 3280 27899
rect 3312 27867 3352 27899
rect 3384 27867 3424 27899
rect 3456 27867 3496 27899
rect 3528 27867 3568 27899
rect 3600 27867 3640 27899
rect 3672 27867 3712 27899
rect 3744 27867 3784 27899
rect 3816 27867 3856 27899
rect 3888 27867 3950 27899
rect 50 27827 3950 27867
rect 50 27795 112 27827
rect 144 27795 184 27827
rect 216 27795 256 27827
rect 288 27795 328 27827
rect 360 27795 400 27827
rect 432 27795 472 27827
rect 504 27795 544 27827
rect 576 27795 616 27827
rect 648 27795 688 27827
rect 720 27795 760 27827
rect 792 27795 832 27827
rect 864 27795 904 27827
rect 936 27795 976 27827
rect 1008 27795 1048 27827
rect 1080 27795 1120 27827
rect 1152 27795 1192 27827
rect 1224 27795 1264 27827
rect 1296 27795 1336 27827
rect 1368 27795 1408 27827
rect 1440 27795 1480 27827
rect 1512 27795 1552 27827
rect 1584 27795 1624 27827
rect 1656 27795 1696 27827
rect 1728 27795 1768 27827
rect 1800 27795 1840 27827
rect 1872 27795 1912 27827
rect 1944 27795 1984 27827
rect 2016 27795 2056 27827
rect 2088 27795 2128 27827
rect 2160 27795 2200 27827
rect 2232 27795 2272 27827
rect 2304 27795 2344 27827
rect 2376 27795 2416 27827
rect 2448 27795 2488 27827
rect 2520 27795 2560 27827
rect 2592 27795 2632 27827
rect 2664 27795 2704 27827
rect 2736 27795 2776 27827
rect 2808 27795 2848 27827
rect 2880 27795 2920 27827
rect 2952 27795 2992 27827
rect 3024 27795 3064 27827
rect 3096 27795 3136 27827
rect 3168 27795 3208 27827
rect 3240 27795 3280 27827
rect 3312 27795 3352 27827
rect 3384 27795 3424 27827
rect 3456 27795 3496 27827
rect 3528 27795 3568 27827
rect 3600 27795 3640 27827
rect 3672 27795 3712 27827
rect 3744 27795 3784 27827
rect 3816 27795 3856 27827
rect 3888 27795 3950 27827
rect 50 27755 3950 27795
rect 50 27723 112 27755
rect 144 27723 184 27755
rect 216 27723 256 27755
rect 288 27723 328 27755
rect 360 27723 400 27755
rect 432 27723 472 27755
rect 504 27723 544 27755
rect 576 27723 616 27755
rect 648 27723 688 27755
rect 720 27723 760 27755
rect 792 27723 832 27755
rect 864 27723 904 27755
rect 936 27723 976 27755
rect 1008 27723 1048 27755
rect 1080 27723 1120 27755
rect 1152 27723 1192 27755
rect 1224 27723 1264 27755
rect 1296 27723 1336 27755
rect 1368 27723 1408 27755
rect 1440 27723 1480 27755
rect 1512 27723 1552 27755
rect 1584 27723 1624 27755
rect 1656 27723 1696 27755
rect 1728 27723 1768 27755
rect 1800 27723 1840 27755
rect 1872 27723 1912 27755
rect 1944 27723 1984 27755
rect 2016 27723 2056 27755
rect 2088 27723 2128 27755
rect 2160 27723 2200 27755
rect 2232 27723 2272 27755
rect 2304 27723 2344 27755
rect 2376 27723 2416 27755
rect 2448 27723 2488 27755
rect 2520 27723 2560 27755
rect 2592 27723 2632 27755
rect 2664 27723 2704 27755
rect 2736 27723 2776 27755
rect 2808 27723 2848 27755
rect 2880 27723 2920 27755
rect 2952 27723 2992 27755
rect 3024 27723 3064 27755
rect 3096 27723 3136 27755
rect 3168 27723 3208 27755
rect 3240 27723 3280 27755
rect 3312 27723 3352 27755
rect 3384 27723 3424 27755
rect 3456 27723 3496 27755
rect 3528 27723 3568 27755
rect 3600 27723 3640 27755
rect 3672 27723 3712 27755
rect 3744 27723 3784 27755
rect 3816 27723 3856 27755
rect 3888 27723 3950 27755
rect 50 27683 3950 27723
rect 50 27651 112 27683
rect 144 27651 184 27683
rect 216 27651 256 27683
rect 288 27651 328 27683
rect 360 27651 400 27683
rect 432 27651 472 27683
rect 504 27651 544 27683
rect 576 27651 616 27683
rect 648 27651 688 27683
rect 720 27651 760 27683
rect 792 27651 832 27683
rect 864 27651 904 27683
rect 936 27651 976 27683
rect 1008 27651 1048 27683
rect 1080 27651 1120 27683
rect 1152 27651 1192 27683
rect 1224 27651 1264 27683
rect 1296 27651 1336 27683
rect 1368 27651 1408 27683
rect 1440 27651 1480 27683
rect 1512 27651 1552 27683
rect 1584 27651 1624 27683
rect 1656 27651 1696 27683
rect 1728 27651 1768 27683
rect 1800 27651 1840 27683
rect 1872 27651 1912 27683
rect 1944 27651 1984 27683
rect 2016 27651 2056 27683
rect 2088 27651 2128 27683
rect 2160 27651 2200 27683
rect 2232 27651 2272 27683
rect 2304 27651 2344 27683
rect 2376 27651 2416 27683
rect 2448 27651 2488 27683
rect 2520 27651 2560 27683
rect 2592 27651 2632 27683
rect 2664 27651 2704 27683
rect 2736 27651 2776 27683
rect 2808 27651 2848 27683
rect 2880 27651 2920 27683
rect 2952 27651 2992 27683
rect 3024 27651 3064 27683
rect 3096 27651 3136 27683
rect 3168 27651 3208 27683
rect 3240 27651 3280 27683
rect 3312 27651 3352 27683
rect 3384 27651 3424 27683
rect 3456 27651 3496 27683
rect 3528 27651 3568 27683
rect 3600 27651 3640 27683
rect 3672 27651 3712 27683
rect 3744 27651 3784 27683
rect 3816 27651 3856 27683
rect 3888 27651 3950 27683
rect 50 27611 3950 27651
rect 50 27579 112 27611
rect 144 27579 184 27611
rect 216 27579 256 27611
rect 288 27579 328 27611
rect 360 27579 400 27611
rect 432 27579 472 27611
rect 504 27579 544 27611
rect 576 27579 616 27611
rect 648 27579 688 27611
rect 720 27579 760 27611
rect 792 27579 832 27611
rect 864 27579 904 27611
rect 936 27579 976 27611
rect 1008 27579 1048 27611
rect 1080 27579 1120 27611
rect 1152 27579 1192 27611
rect 1224 27579 1264 27611
rect 1296 27579 1336 27611
rect 1368 27579 1408 27611
rect 1440 27579 1480 27611
rect 1512 27579 1552 27611
rect 1584 27579 1624 27611
rect 1656 27579 1696 27611
rect 1728 27579 1768 27611
rect 1800 27579 1840 27611
rect 1872 27579 1912 27611
rect 1944 27579 1984 27611
rect 2016 27579 2056 27611
rect 2088 27579 2128 27611
rect 2160 27579 2200 27611
rect 2232 27579 2272 27611
rect 2304 27579 2344 27611
rect 2376 27579 2416 27611
rect 2448 27579 2488 27611
rect 2520 27579 2560 27611
rect 2592 27579 2632 27611
rect 2664 27579 2704 27611
rect 2736 27579 2776 27611
rect 2808 27579 2848 27611
rect 2880 27579 2920 27611
rect 2952 27579 2992 27611
rect 3024 27579 3064 27611
rect 3096 27579 3136 27611
rect 3168 27579 3208 27611
rect 3240 27579 3280 27611
rect 3312 27579 3352 27611
rect 3384 27579 3424 27611
rect 3456 27579 3496 27611
rect 3528 27579 3568 27611
rect 3600 27579 3640 27611
rect 3672 27579 3712 27611
rect 3744 27579 3784 27611
rect 3816 27579 3856 27611
rect 3888 27579 3950 27611
rect 50 27539 3950 27579
rect 50 27507 112 27539
rect 144 27507 184 27539
rect 216 27507 256 27539
rect 288 27507 328 27539
rect 360 27507 400 27539
rect 432 27507 472 27539
rect 504 27507 544 27539
rect 576 27507 616 27539
rect 648 27507 688 27539
rect 720 27507 760 27539
rect 792 27507 832 27539
rect 864 27507 904 27539
rect 936 27507 976 27539
rect 1008 27507 1048 27539
rect 1080 27507 1120 27539
rect 1152 27507 1192 27539
rect 1224 27507 1264 27539
rect 1296 27507 1336 27539
rect 1368 27507 1408 27539
rect 1440 27507 1480 27539
rect 1512 27507 1552 27539
rect 1584 27507 1624 27539
rect 1656 27507 1696 27539
rect 1728 27507 1768 27539
rect 1800 27507 1840 27539
rect 1872 27507 1912 27539
rect 1944 27507 1984 27539
rect 2016 27507 2056 27539
rect 2088 27507 2128 27539
rect 2160 27507 2200 27539
rect 2232 27507 2272 27539
rect 2304 27507 2344 27539
rect 2376 27507 2416 27539
rect 2448 27507 2488 27539
rect 2520 27507 2560 27539
rect 2592 27507 2632 27539
rect 2664 27507 2704 27539
rect 2736 27507 2776 27539
rect 2808 27507 2848 27539
rect 2880 27507 2920 27539
rect 2952 27507 2992 27539
rect 3024 27507 3064 27539
rect 3096 27507 3136 27539
rect 3168 27507 3208 27539
rect 3240 27507 3280 27539
rect 3312 27507 3352 27539
rect 3384 27507 3424 27539
rect 3456 27507 3496 27539
rect 3528 27507 3568 27539
rect 3600 27507 3640 27539
rect 3672 27507 3712 27539
rect 3744 27507 3784 27539
rect 3816 27507 3856 27539
rect 3888 27507 3950 27539
rect 50 27467 3950 27507
rect 50 27435 112 27467
rect 144 27435 184 27467
rect 216 27435 256 27467
rect 288 27435 328 27467
rect 360 27435 400 27467
rect 432 27435 472 27467
rect 504 27435 544 27467
rect 576 27435 616 27467
rect 648 27435 688 27467
rect 720 27435 760 27467
rect 792 27435 832 27467
rect 864 27435 904 27467
rect 936 27435 976 27467
rect 1008 27435 1048 27467
rect 1080 27435 1120 27467
rect 1152 27435 1192 27467
rect 1224 27435 1264 27467
rect 1296 27435 1336 27467
rect 1368 27435 1408 27467
rect 1440 27435 1480 27467
rect 1512 27435 1552 27467
rect 1584 27435 1624 27467
rect 1656 27435 1696 27467
rect 1728 27435 1768 27467
rect 1800 27435 1840 27467
rect 1872 27435 1912 27467
rect 1944 27435 1984 27467
rect 2016 27435 2056 27467
rect 2088 27435 2128 27467
rect 2160 27435 2200 27467
rect 2232 27435 2272 27467
rect 2304 27435 2344 27467
rect 2376 27435 2416 27467
rect 2448 27435 2488 27467
rect 2520 27435 2560 27467
rect 2592 27435 2632 27467
rect 2664 27435 2704 27467
rect 2736 27435 2776 27467
rect 2808 27435 2848 27467
rect 2880 27435 2920 27467
rect 2952 27435 2992 27467
rect 3024 27435 3064 27467
rect 3096 27435 3136 27467
rect 3168 27435 3208 27467
rect 3240 27435 3280 27467
rect 3312 27435 3352 27467
rect 3384 27435 3424 27467
rect 3456 27435 3496 27467
rect 3528 27435 3568 27467
rect 3600 27435 3640 27467
rect 3672 27435 3712 27467
rect 3744 27435 3784 27467
rect 3816 27435 3856 27467
rect 3888 27435 3950 27467
rect 50 27395 3950 27435
rect 50 27363 112 27395
rect 144 27363 184 27395
rect 216 27363 256 27395
rect 288 27363 328 27395
rect 360 27363 400 27395
rect 432 27363 472 27395
rect 504 27363 544 27395
rect 576 27363 616 27395
rect 648 27363 688 27395
rect 720 27363 760 27395
rect 792 27363 832 27395
rect 864 27363 904 27395
rect 936 27363 976 27395
rect 1008 27363 1048 27395
rect 1080 27363 1120 27395
rect 1152 27363 1192 27395
rect 1224 27363 1264 27395
rect 1296 27363 1336 27395
rect 1368 27363 1408 27395
rect 1440 27363 1480 27395
rect 1512 27363 1552 27395
rect 1584 27363 1624 27395
rect 1656 27363 1696 27395
rect 1728 27363 1768 27395
rect 1800 27363 1840 27395
rect 1872 27363 1912 27395
rect 1944 27363 1984 27395
rect 2016 27363 2056 27395
rect 2088 27363 2128 27395
rect 2160 27363 2200 27395
rect 2232 27363 2272 27395
rect 2304 27363 2344 27395
rect 2376 27363 2416 27395
rect 2448 27363 2488 27395
rect 2520 27363 2560 27395
rect 2592 27363 2632 27395
rect 2664 27363 2704 27395
rect 2736 27363 2776 27395
rect 2808 27363 2848 27395
rect 2880 27363 2920 27395
rect 2952 27363 2992 27395
rect 3024 27363 3064 27395
rect 3096 27363 3136 27395
rect 3168 27363 3208 27395
rect 3240 27363 3280 27395
rect 3312 27363 3352 27395
rect 3384 27363 3424 27395
rect 3456 27363 3496 27395
rect 3528 27363 3568 27395
rect 3600 27363 3640 27395
rect 3672 27363 3712 27395
rect 3744 27363 3784 27395
rect 3816 27363 3856 27395
rect 3888 27363 3950 27395
rect 50 27323 3950 27363
rect 50 27291 112 27323
rect 144 27291 184 27323
rect 216 27291 256 27323
rect 288 27291 328 27323
rect 360 27291 400 27323
rect 432 27291 472 27323
rect 504 27291 544 27323
rect 576 27291 616 27323
rect 648 27291 688 27323
rect 720 27291 760 27323
rect 792 27291 832 27323
rect 864 27291 904 27323
rect 936 27291 976 27323
rect 1008 27291 1048 27323
rect 1080 27291 1120 27323
rect 1152 27291 1192 27323
rect 1224 27291 1264 27323
rect 1296 27291 1336 27323
rect 1368 27291 1408 27323
rect 1440 27291 1480 27323
rect 1512 27291 1552 27323
rect 1584 27291 1624 27323
rect 1656 27291 1696 27323
rect 1728 27291 1768 27323
rect 1800 27291 1840 27323
rect 1872 27291 1912 27323
rect 1944 27291 1984 27323
rect 2016 27291 2056 27323
rect 2088 27291 2128 27323
rect 2160 27291 2200 27323
rect 2232 27291 2272 27323
rect 2304 27291 2344 27323
rect 2376 27291 2416 27323
rect 2448 27291 2488 27323
rect 2520 27291 2560 27323
rect 2592 27291 2632 27323
rect 2664 27291 2704 27323
rect 2736 27291 2776 27323
rect 2808 27291 2848 27323
rect 2880 27291 2920 27323
rect 2952 27291 2992 27323
rect 3024 27291 3064 27323
rect 3096 27291 3136 27323
rect 3168 27291 3208 27323
rect 3240 27291 3280 27323
rect 3312 27291 3352 27323
rect 3384 27291 3424 27323
rect 3456 27291 3496 27323
rect 3528 27291 3568 27323
rect 3600 27291 3640 27323
rect 3672 27291 3712 27323
rect 3744 27291 3784 27323
rect 3816 27291 3856 27323
rect 3888 27291 3950 27323
rect 50 27251 3950 27291
rect 50 27219 112 27251
rect 144 27219 184 27251
rect 216 27219 256 27251
rect 288 27219 328 27251
rect 360 27219 400 27251
rect 432 27219 472 27251
rect 504 27219 544 27251
rect 576 27219 616 27251
rect 648 27219 688 27251
rect 720 27219 760 27251
rect 792 27219 832 27251
rect 864 27219 904 27251
rect 936 27219 976 27251
rect 1008 27219 1048 27251
rect 1080 27219 1120 27251
rect 1152 27219 1192 27251
rect 1224 27219 1264 27251
rect 1296 27219 1336 27251
rect 1368 27219 1408 27251
rect 1440 27219 1480 27251
rect 1512 27219 1552 27251
rect 1584 27219 1624 27251
rect 1656 27219 1696 27251
rect 1728 27219 1768 27251
rect 1800 27219 1840 27251
rect 1872 27219 1912 27251
rect 1944 27219 1984 27251
rect 2016 27219 2056 27251
rect 2088 27219 2128 27251
rect 2160 27219 2200 27251
rect 2232 27219 2272 27251
rect 2304 27219 2344 27251
rect 2376 27219 2416 27251
rect 2448 27219 2488 27251
rect 2520 27219 2560 27251
rect 2592 27219 2632 27251
rect 2664 27219 2704 27251
rect 2736 27219 2776 27251
rect 2808 27219 2848 27251
rect 2880 27219 2920 27251
rect 2952 27219 2992 27251
rect 3024 27219 3064 27251
rect 3096 27219 3136 27251
rect 3168 27219 3208 27251
rect 3240 27219 3280 27251
rect 3312 27219 3352 27251
rect 3384 27219 3424 27251
rect 3456 27219 3496 27251
rect 3528 27219 3568 27251
rect 3600 27219 3640 27251
rect 3672 27219 3712 27251
rect 3744 27219 3784 27251
rect 3816 27219 3856 27251
rect 3888 27219 3950 27251
rect 50 27179 3950 27219
rect 50 27147 112 27179
rect 144 27147 184 27179
rect 216 27147 256 27179
rect 288 27147 328 27179
rect 360 27147 400 27179
rect 432 27147 472 27179
rect 504 27147 544 27179
rect 576 27147 616 27179
rect 648 27147 688 27179
rect 720 27147 760 27179
rect 792 27147 832 27179
rect 864 27147 904 27179
rect 936 27147 976 27179
rect 1008 27147 1048 27179
rect 1080 27147 1120 27179
rect 1152 27147 1192 27179
rect 1224 27147 1264 27179
rect 1296 27147 1336 27179
rect 1368 27147 1408 27179
rect 1440 27147 1480 27179
rect 1512 27147 1552 27179
rect 1584 27147 1624 27179
rect 1656 27147 1696 27179
rect 1728 27147 1768 27179
rect 1800 27147 1840 27179
rect 1872 27147 1912 27179
rect 1944 27147 1984 27179
rect 2016 27147 2056 27179
rect 2088 27147 2128 27179
rect 2160 27147 2200 27179
rect 2232 27147 2272 27179
rect 2304 27147 2344 27179
rect 2376 27147 2416 27179
rect 2448 27147 2488 27179
rect 2520 27147 2560 27179
rect 2592 27147 2632 27179
rect 2664 27147 2704 27179
rect 2736 27147 2776 27179
rect 2808 27147 2848 27179
rect 2880 27147 2920 27179
rect 2952 27147 2992 27179
rect 3024 27147 3064 27179
rect 3096 27147 3136 27179
rect 3168 27147 3208 27179
rect 3240 27147 3280 27179
rect 3312 27147 3352 27179
rect 3384 27147 3424 27179
rect 3456 27147 3496 27179
rect 3528 27147 3568 27179
rect 3600 27147 3640 27179
rect 3672 27147 3712 27179
rect 3744 27147 3784 27179
rect 3816 27147 3856 27179
rect 3888 27147 3950 27179
rect 50 27107 3950 27147
rect 50 27075 112 27107
rect 144 27075 184 27107
rect 216 27075 256 27107
rect 288 27075 328 27107
rect 360 27075 400 27107
rect 432 27075 472 27107
rect 504 27075 544 27107
rect 576 27075 616 27107
rect 648 27075 688 27107
rect 720 27075 760 27107
rect 792 27075 832 27107
rect 864 27075 904 27107
rect 936 27075 976 27107
rect 1008 27075 1048 27107
rect 1080 27075 1120 27107
rect 1152 27075 1192 27107
rect 1224 27075 1264 27107
rect 1296 27075 1336 27107
rect 1368 27075 1408 27107
rect 1440 27075 1480 27107
rect 1512 27075 1552 27107
rect 1584 27075 1624 27107
rect 1656 27075 1696 27107
rect 1728 27075 1768 27107
rect 1800 27075 1840 27107
rect 1872 27075 1912 27107
rect 1944 27075 1984 27107
rect 2016 27075 2056 27107
rect 2088 27075 2128 27107
rect 2160 27075 2200 27107
rect 2232 27075 2272 27107
rect 2304 27075 2344 27107
rect 2376 27075 2416 27107
rect 2448 27075 2488 27107
rect 2520 27075 2560 27107
rect 2592 27075 2632 27107
rect 2664 27075 2704 27107
rect 2736 27075 2776 27107
rect 2808 27075 2848 27107
rect 2880 27075 2920 27107
rect 2952 27075 2992 27107
rect 3024 27075 3064 27107
rect 3096 27075 3136 27107
rect 3168 27075 3208 27107
rect 3240 27075 3280 27107
rect 3312 27075 3352 27107
rect 3384 27075 3424 27107
rect 3456 27075 3496 27107
rect 3528 27075 3568 27107
rect 3600 27075 3640 27107
rect 3672 27075 3712 27107
rect 3744 27075 3784 27107
rect 3816 27075 3856 27107
rect 3888 27075 3950 27107
rect 50 27035 3950 27075
rect 50 27003 112 27035
rect 144 27003 184 27035
rect 216 27003 256 27035
rect 288 27003 328 27035
rect 360 27003 400 27035
rect 432 27003 472 27035
rect 504 27003 544 27035
rect 576 27003 616 27035
rect 648 27003 688 27035
rect 720 27003 760 27035
rect 792 27003 832 27035
rect 864 27003 904 27035
rect 936 27003 976 27035
rect 1008 27003 1048 27035
rect 1080 27003 1120 27035
rect 1152 27003 1192 27035
rect 1224 27003 1264 27035
rect 1296 27003 1336 27035
rect 1368 27003 1408 27035
rect 1440 27003 1480 27035
rect 1512 27003 1552 27035
rect 1584 27003 1624 27035
rect 1656 27003 1696 27035
rect 1728 27003 1768 27035
rect 1800 27003 1840 27035
rect 1872 27003 1912 27035
rect 1944 27003 1984 27035
rect 2016 27003 2056 27035
rect 2088 27003 2128 27035
rect 2160 27003 2200 27035
rect 2232 27003 2272 27035
rect 2304 27003 2344 27035
rect 2376 27003 2416 27035
rect 2448 27003 2488 27035
rect 2520 27003 2560 27035
rect 2592 27003 2632 27035
rect 2664 27003 2704 27035
rect 2736 27003 2776 27035
rect 2808 27003 2848 27035
rect 2880 27003 2920 27035
rect 2952 27003 2992 27035
rect 3024 27003 3064 27035
rect 3096 27003 3136 27035
rect 3168 27003 3208 27035
rect 3240 27003 3280 27035
rect 3312 27003 3352 27035
rect 3384 27003 3424 27035
rect 3456 27003 3496 27035
rect 3528 27003 3568 27035
rect 3600 27003 3640 27035
rect 3672 27003 3712 27035
rect 3744 27003 3784 27035
rect 3816 27003 3856 27035
rect 3888 27003 3950 27035
rect 50 26963 3950 27003
rect 50 26931 112 26963
rect 144 26931 184 26963
rect 216 26931 256 26963
rect 288 26931 328 26963
rect 360 26931 400 26963
rect 432 26931 472 26963
rect 504 26931 544 26963
rect 576 26931 616 26963
rect 648 26931 688 26963
rect 720 26931 760 26963
rect 792 26931 832 26963
rect 864 26931 904 26963
rect 936 26931 976 26963
rect 1008 26931 1048 26963
rect 1080 26931 1120 26963
rect 1152 26931 1192 26963
rect 1224 26931 1264 26963
rect 1296 26931 1336 26963
rect 1368 26931 1408 26963
rect 1440 26931 1480 26963
rect 1512 26931 1552 26963
rect 1584 26931 1624 26963
rect 1656 26931 1696 26963
rect 1728 26931 1768 26963
rect 1800 26931 1840 26963
rect 1872 26931 1912 26963
rect 1944 26931 1984 26963
rect 2016 26931 2056 26963
rect 2088 26931 2128 26963
rect 2160 26931 2200 26963
rect 2232 26931 2272 26963
rect 2304 26931 2344 26963
rect 2376 26931 2416 26963
rect 2448 26931 2488 26963
rect 2520 26931 2560 26963
rect 2592 26931 2632 26963
rect 2664 26931 2704 26963
rect 2736 26931 2776 26963
rect 2808 26931 2848 26963
rect 2880 26931 2920 26963
rect 2952 26931 2992 26963
rect 3024 26931 3064 26963
rect 3096 26931 3136 26963
rect 3168 26931 3208 26963
rect 3240 26931 3280 26963
rect 3312 26931 3352 26963
rect 3384 26931 3424 26963
rect 3456 26931 3496 26963
rect 3528 26931 3568 26963
rect 3600 26931 3640 26963
rect 3672 26931 3712 26963
rect 3744 26931 3784 26963
rect 3816 26931 3856 26963
rect 3888 26931 3950 26963
rect 50 26891 3950 26931
rect 50 26859 112 26891
rect 144 26859 184 26891
rect 216 26859 256 26891
rect 288 26859 328 26891
rect 360 26859 400 26891
rect 432 26859 472 26891
rect 504 26859 544 26891
rect 576 26859 616 26891
rect 648 26859 688 26891
rect 720 26859 760 26891
rect 792 26859 832 26891
rect 864 26859 904 26891
rect 936 26859 976 26891
rect 1008 26859 1048 26891
rect 1080 26859 1120 26891
rect 1152 26859 1192 26891
rect 1224 26859 1264 26891
rect 1296 26859 1336 26891
rect 1368 26859 1408 26891
rect 1440 26859 1480 26891
rect 1512 26859 1552 26891
rect 1584 26859 1624 26891
rect 1656 26859 1696 26891
rect 1728 26859 1768 26891
rect 1800 26859 1840 26891
rect 1872 26859 1912 26891
rect 1944 26859 1984 26891
rect 2016 26859 2056 26891
rect 2088 26859 2128 26891
rect 2160 26859 2200 26891
rect 2232 26859 2272 26891
rect 2304 26859 2344 26891
rect 2376 26859 2416 26891
rect 2448 26859 2488 26891
rect 2520 26859 2560 26891
rect 2592 26859 2632 26891
rect 2664 26859 2704 26891
rect 2736 26859 2776 26891
rect 2808 26859 2848 26891
rect 2880 26859 2920 26891
rect 2952 26859 2992 26891
rect 3024 26859 3064 26891
rect 3096 26859 3136 26891
rect 3168 26859 3208 26891
rect 3240 26859 3280 26891
rect 3312 26859 3352 26891
rect 3384 26859 3424 26891
rect 3456 26859 3496 26891
rect 3528 26859 3568 26891
rect 3600 26859 3640 26891
rect 3672 26859 3712 26891
rect 3744 26859 3784 26891
rect 3816 26859 3856 26891
rect 3888 26859 3950 26891
rect 50 26819 3950 26859
rect 50 26787 112 26819
rect 144 26787 184 26819
rect 216 26787 256 26819
rect 288 26787 328 26819
rect 360 26787 400 26819
rect 432 26787 472 26819
rect 504 26787 544 26819
rect 576 26787 616 26819
rect 648 26787 688 26819
rect 720 26787 760 26819
rect 792 26787 832 26819
rect 864 26787 904 26819
rect 936 26787 976 26819
rect 1008 26787 1048 26819
rect 1080 26787 1120 26819
rect 1152 26787 1192 26819
rect 1224 26787 1264 26819
rect 1296 26787 1336 26819
rect 1368 26787 1408 26819
rect 1440 26787 1480 26819
rect 1512 26787 1552 26819
rect 1584 26787 1624 26819
rect 1656 26787 1696 26819
rect 1728 26787 1768 26819
rect 1800 26787 1840 26819
rect 1872 26787 1912 26819
rect 1944 26787 1984 26819
rect 2016 26787 2056 26819
rect 2088 26787 2128 26819
rect 2160 26787 2200 26819
rect 2232 26787 2272 26819
rect 2304 26787 2344 26819
rect 2376 26787 2416 26819
rect 2448 26787 2488 26819
rect 2520 26787 2560 26819
rect 2592 26787 2632 26819
rect 2664 26787 2704 26819
rect 2736 26787 2776 26819
rect 2808 26787 2848 26819
rect 2880 26787 2920 26819
rect 2952 26787 2992 26819
rect 3024 26787 3064 26819
rect 3096 26787 3136 26819
rect 3168 26787 3208 26819
rect 3240 26787 3280 26819
rect 3312 26787 3352 26819
rect 3384 26787 3424 26819
rect 3456 26787 3496 26819
rect 3528 26787 3568 26819
rect 3600 26787 3640 26819
rect 3672 26787 3712 26819
rect 3744 26787 3784 26819
rect 3816 26787 3856 26819
rect 3888 26787 3950 26819
rect 50 26747 3950 26787
rect 50 26715 112 26747
rect 144 26715 184 26747
rect 216 26715 256 26747
rect 288 26715 328 26747
rect 360 26715 400 26747
rect 432 26715 472 26747
rect 504 26715 544 26747
rect 576 26715 616 26747
rect 648 26715 688 26747
rect 720 26715 760 26747
rect 792 26715 832 26747
rect 864 26715 904 26747
rect 936 26715 976 26747
rect 1008 26715 1048 26747
rect 1080 26715 1120 26747
rect 1152 26715 1192 26747
rect 1224 26715 1264 26747
rect 1296 26715 1336 26747
rect 1368 26715 1408 26747
rect 1440 26715 1480 26747
rect 1512 26715 1552 26747
rect 1584 26715 1624 26747
rect 1656 26715 1696 26747
rect 1728 26715 1768 26747
rect 1800 26715 1840 26747
rect 1872 26715 1912 26747
rect 1944 26715 1984 26747
rect 2016 26715 2056 26747
rect 2088 26715 2128 26747
rect 2160 26715 2200 26747
rect 2232 26715 2272 26747
rect 2304 26715 2344 26747
rect 2376 26715 2416 26747
rect 2448 26715 2488 26747
rect 2520 26715 2560 26747
rect 2592 26715 2632 26747
rect 2664 26715 2704 26747
rect 2736 26715 2776 26747
rect 2808 26715 2848 26747
rect 2880 26715 2920 26747
rect 2952 26715 2992 26747
rect 3024 26715 3064 26747
rect 3096 26715 3136 26747
rect 3168 26715 3208 26747
rect 3240 26715 3280 26747
rect 3312 26715 3352 26747
rect 3384 26715 3424 26747
rect 3456 26715 3496 26747
rect 3528 26715 3568 26747
rect 3600 26715 3640 26747
rect 3672 26715 3712 26747
rect 3744 26715 3784 26747
rect 3816 26715 3856 26747
rect 3888 26715 3950 26747
rect 50 26675 3950 26715
rect 50 26643 112 26675
rect 144 26643 184 26675
rect 216 26643 256 26675
rect 288 26643 328 26675
rect 360 26643 400 26675
rect 432 26643 472 26675
rect 504 26643 544 26675
rect 576 26643 616 26675
rect 648 26643 688 26675
rect 720 26643 760 26675
rect 792 26643 832 26675
rect 864 26643 904 26675
rect 936 26643 976 26675
rect 1008 26643 1048 26675
rect 1080 26643 1120 26675
rect 1152 26643 1192 26675
rect 1224 26643 1264 26675
rect 1296 26643 1336 26675
rect 1368 26643 1408 26675
rect 1440 26643 1480 26675
rect 1512 26643 1552 26675
rect 1584 26643 1624 26675
rect 1656 26643 1696 26675
rect 1728 26643 1768 26675
rect 1800 26643 1840 26675
rect 1872 26643 1912 26675
rect 1944 26643 1984 26675
rect 2016 26643 2056 26675
rect 2088 26643 2128 26675
rect 2160 26643 2200 26675
rect 2232 26643 2272 26675
rect 2304 26643 2344 26675
rect 2376 26643 2416 26675
rect 2448 26643 2488 26675
rect 2520 26643 2560 26675
rect 2592 26643 2632 26675
rect 2664 26643 2704 26675
rect 2736 26643 2776 26675
rect 2808 26643 2848 26675
rect 2880 26643 2920 26675
rect 2952 26643 2992 26675
rect 3024 26643 3064 26675
rect 3096 26643 3136 26675
rect 3168 26643 3208 26675
rect 3240 26643 3280 26675
rect 3312 26643 3352 26675
rect 3384 26643 3424 26675
rect 3456 26643 3496 26675
rect 3528 26643 3568 26675
rect 3600 26643 3640 26675
rect 3672 26643 3712 26675
rect 3744 26643 3784 26675
rect 3816 26643 3856 26675
rect 3888 26643 3950 26675
rect 50 26603 3950 26643
rect 50 26571 112 26603
rect 144 26571 184 26603
rect 216 26571 256 26603
rect 288 26571 328 26603
rect 360 26571 400 26603
rect 432 26571 472 26603
rect 504 26571 544 26603
rect 576 26571 616 26603
rect 648 26571 688 26603
rect 720 26571 760 26603
rect 792 26571 832 26603
rect 864 26571 904 26603
rect 936 26571 976 26603
rect 1008 26571 1048 26603
rect 1080 26571 1120 26603
rect 1152 26571 1192 26603
rect 1224 26571 1264 26603
rect 1296 26571 1336 26603
rect 1368 26571 1408 26603
rect 1440 26571 1480 26603
rect 1512 26571 1552 26603
rect 1584 26571 1624 26603
rect 1656 26571 1696 26603
rect 1728 26571 1768 26603
rect 1800 26571 1840 26603
rect 1872 26571 1912 26603
rect 1944 26571 1984 26603
rect 2016 26571 2056 26603
rect 2088 26571 2128 26603
rect 2160 26571 2200 26603
rect 2232 26571 2272 26603
rect 2304 26571 2344 26603
rect 2376 26571 2416 26603
rect 2448 26571 2488 26603
rect 2520 26571 2560 26603
rect 2592 26571 2632 26603
rect 2664 26571 2704 26603
rect 2736 26571 2776 26603
rect 2808 26571 2848 26603
rect 2880 26571 2920 26603
rect 2952 26571 2992 26603
rect 3024 26571 3064 26603
rect 3096 26571 3136 26603
rect 3168 26571 3208 26603
rect 3240 26571 3280 26603
rect 3312 26571 3352 26603
rect 3384 26571 3424 26603
rect 3456 26571 3496 26603
rect 3528 26571 3568 26603
rect 3600 26571 3640 26603
rect 3672 26571 3712 26603
rect 3744 26571 3784 26603
rect 3816 26571 3856 26603
rect 3888 26571 3950 26603
rect 50 26531 3950 26571
rect 50 26499 112 26531
rect 144 26499 184 26531
rect 216 26499 256 26531
rect 288 26499 328 26531
rect 360 26499 400 26531
rect 432 26499 472 26531
rect 504 26499 544 26531
rect 576 26499 616 26531
rect 648 26499 688 26531
rect 720 26499 760 26531
rect 792 26499 832 26531
rect 864 26499 904 26531
rect 936 26499 976 26531
rect 1008 26499 1048 26531
rect 1080 26499 1120 26531
rect 1152 26499 1192 26531
rect 1224 26499 1264 26531
rect 1296 26499 1336 26531
rect 1368 26499 1408 26531
rect 1440 26499 1480 26531
rect 1512 26499 1552 26531
rect 1584 26499 1624 26531
rect 1656 26499 1696 26531
rect 1728 26499 1768 26531
rect 1800 26499 1840 26531
rect 1872 26499 1912 26531
rect 1944 26499 1984 26531
rect 2016 26499 2056 26531
rect 2088 26499 2128 26531
rect 2160 26499 2200 26531
rect 2232 26499 2272 26531
rect 2304 26499 2344 26531
rect 2376 26499 2416 26531
rect 2448 26499 2488 26531
rect 2520 26499 2560 26531
rect 2592 26499 2632 26531
rect 2664 26499 2704 26531
rect 2736 26499 2776 26531
rect 2808 26499 2848 26531
rect 2880 26499 2920 26531
rect 2952 26499 2992 26531
rect 3024 26499 3064 26531
rect 3096 26499 3136 26531
rect 3168 26499 3208 26531
rect 3240 26499 3280 26531
rect 3312 26499 3352 26531
rect 3384 26499 3424 26531
rect 3456 26499 3496 26531
rect 3528 26499 3568 26531
rect 3600 26499 3640 26531
rect 3672 26499 3712 26531
rect 3744 26499 3784 26531
rect 3816 26499 3856 26531
rect 3888 26499 3950 26531
rect 50 26459 3950 26499
rect 50 26427 112 26459
rect 144 26427 184 26459
rect 216 26427 256 26459
rect 288 26427 328 26459
rect 360 26427 400 26459
rect 432 26427 472 26459
rect 504 26427 544 26459
rect 576 26427 616 26459
rect 648 26427 688 26459
rect 720 26427 760 26459
rect 792 26427 832 26459
rect 864 26427 904 26459
rect 936 26427 976 26459
rect 1008 26427 1048 26459
rect 1080 26427 1120 26459
rect 1152 26427 1192 26459
rect 1224 26427 1264 26459
rect 1296 26427 1336 26459
rect 1368 26427 1408 26459
rect 1440 26427 1480 26459
rect 1512 26427 1552 26459
rect 1584 26427 1624 26459
rect 1656 26427 1696 26459
rect 1728 26427 1768 26459
rect 1800 26427 1840 26459
rect 1872 26427 1912 26459
rect 1944 26427 1984 26459
rect 2016 26427 2056 26459
rect 2088 26427 2128 26459
rect 2160 26427 2200 26459
rect 2232 26427 2272 26459
rect 2304 26427 2344 26459
rect 2376 26427 2416 26459
rect 2448 26427 2488 26459
rect 2520 26427 2560 26459
rect 2592 26427 2632 26459
rect 2664 26427 2704 26459
rect 2736 26427 2776 26459
rect 2808 26427 2848 26459
rect 2880 26427 2920 26459
rect 2952 26427 2992 26459
rect 3024 26427 3064 26459
rect 3096 26427 3136 26459
rect 3168 26427 3208 26459
rect 3240 26427 3280 26459
rect 3312 26427 3352 26459
rect 3384 26427 3424 26459
rect 3456 26427 3496 26459
rect 3528 26427 3568 26459
rect 3600 26427 3640 26459
rect 3672 26427 3712 26459
rect 3744 26427 3784 26459
rect 3816 26427 3856 26459
rect 3888 26427 3950 26459
rect 50 26387 3950 26427
rect 50 26355 112 26387
rect 144 26355 184 26387
rect 216 26355 256 26387
rect 288 26355 328 26387
rect 360 26355 400 26387
rect 432 26355 472 26387
rect 504 26355 544 26387
rect 576 26355 616 26387
rect 648 26355 688 26387
rect 720 26355 760 26387
rect 792 26355 832 26387
rect 864 26355 904 26387
rect 936 26355 976 26387
rect 1008 26355 1048 26387
rect 1080 26355 1120 26387
rect 1152 26355 1192 26387
rect 1224 26355 1264 26387
rect 1296 26355 1336 26387
rect 1368 26355 1408 26387
rect 1440 26355 1480 26387
rect 1512 26355 1552 26387
rect 1584 26355 1624 26387
rect 1656 26355 1696 26387
rect 1728 26355 1768 26387
rect 1800 26355 1840 26387
rect 1872 26355 1912 26387
rect 1944 26355 1984 26387
rect 2016 26355 2056 26387
rect 2088 26355 2128 26387
rect 2160 26355 2200 26387
rect 2232 26355 2272 26387
rect 2304 26355 2344 26387
rect 2376 26355 2416 26387
rect 2448 26355 2488 26387
rect 2520 26355 2560 26387
rect 2592 26355 2632 26387
rect 2664 26355 2704 26387
rect 2736 26355 2776 26387
rect 2808 26355 2848 26387
rect 2880 26355 2920 26387
rect 2952 26355 2992 26387
rect 3024 26355 3064 26387
rect 3096 26355 3136 26387
rect 3168 26355 3208 26387
rect 3240 26355 3280 26387
rect 3312 26355 3352 26387
rect 3384 26355 3424 26387
rect 3456 26355 3496 26387
rect 3528 26355 3568 26387
rect 3600 26355 3640 26387
rect 3672 26355 3712 26387
rect 3744 26355 3784 26387
rect 3816 26355 3856 26387
rect 3888 26355 3950 26387
rect 50 26315 3950 26355
rect 50 26283 112 26315
rect 144 26283 184 26315
rect 216 26283 256 26315
rect 288 26283 328 26315
rect 360 26283 400 26315
rect 432 26283 472 26315
rect 504 26283 544 26315
rect 576 26283 616 26315
rect 648 26283 688 26315
rect 720 26283 760 26315
rect 792 26283 832 26315
rect 864 26283 904 26315
rect 936 26283 976 26315
rect 1008 26283 1048 26315
rect 1080 26283 1120 26315
rect 1152 26283 1192 26315
rect 1224 26283 1264 26315
rect 1296 26283 1336 26315
rect 1368 26283 1408 26315
rect 1440 26283 1480 26315
rect 1512 26283 1552 26315
rect 1584 26283 1624 26315
rect 1656 26283 1696 26315
rect 1728 26283 1768 26315
rect 1800 26283 1840 26315
rect 1872 26283 1912 26315
rect 1944 26283 1984 26315
rect 2016 26283 2056 26315
rect 2088 26283 2128 26315
rect 2160 26283 2200 26315
rect 2232 26283 2272 26315
rect 2304 26283 2344 26315
rect 2376 26283 2416 26315
rect 2448 26283 2488 26315
rect 2520 26283 2560 26315
rect 2592 26283 2632 26315
rect 2664 26283 2704 26315
rect 2736 26283 2776 26315
rect 2808 26283 2848 26315
rect 2880 26283 2920 26315
rect 2952 26283 2992 26315
rect 3024 26283 3064 26315
rect 3096 26283 3136 26315
rect 3168 26283 3208 26315
rect 3240 26283 3280 26315
rect 3312 26283 3352 26315
rect 3384 26283 3424 26315
rect 3456 26283 3496 26315
rect 3528 26283 3568 26315
rect 3600 26283 3640 26315
rect 3672 26283 3712 26315
rect 3744 26283 3784 26315
rect 3816 26283 3856 26315
rect 3888 26283 3950 26315
rect 50 26243 3950 26283
rect 50 26211 112 26243
rect 144 26211 184 26243
rect 216 26211 256 26243
rect 288 26211 328 26243
rect 360 26211 400 26243
rect 432 26211 472 26243
rect 504 26211 544 26243
rect 576 26211 616 26243
rect 648 26211 688 26243
rect 720 26211 760 26243
rect 792 26211 832 26243
rect 864 26211 904 26243
rect 936 26211 976 26243
rect 1008 26211 1048 26243
rect 1080 26211 1120 26243
rect 1152 26211 1192 26243
rect 1224 26211 1264 26243
rect 1296 26211 1336 26243
rect 1368 26211 1408 26243
rect 1440 26211 1480 26243
rect 1512 26211 1552 26243
rect 1584 26211 1624 26243
rect 1656 26211 1696 26243
rect 1728 26211 1768 26243
rect 1800 26211 1840 26243
rect 1872 26211 1912 26243
rect 1944 26211 1984 26243
rect 2016 26211 2056 26243
rect 2088 26211 2128 26243
rect 2160 26211 2200 26243
rect 2232 26211 2272 26243
rect 2304 26211 2344 26243
rect 2376 26211 2416 26243
rect 2448 26211 2488 26243
rect 2520 26211 2560 26243
rect 2592 26211 2632 26243
rect 2664 26211 2704 26243
rect 2736 26211 2776 26243
rect 2808 26211 2848 26243
rect 2880 26211 2920 26243
rect 2952 26211 2992 26243
rect 3024 26211 3064 26243
rect 3096 26211 3136 26243
rect 3168 26211 3208 26243
rect 3240 26211 3280 26243
rect 3312 26211 3352 26243
rect 3384 26211 3424 26243
rect 3456 26211 3496 26243
rect 3528 26211 3568 26243
rect 3600 26211 3640 26243
rect 3672 26211 3712 26243
rect 3744 26211 3784 26243
rect 3816 26211 3856 26243
rect 3888 26211 3950 26243
rect 50 26171 3950 26211
rect 50 26139 112 26171
rect 144 26139 184 26171
rect 216 26139 256 26171
rect 288 26139 328 26171
rect 360 26139 400 26171
rect 432 26139 472 26171
rect 504 26139 544 26171
rect 576 26139 616 26171
rect 648 26139 688 26171
rect 720 26139 760 26171
rect 792 26139 832 26171
rect 864 26139 904 26171
rect 936 26139 976 26171
rect 1008 26139 1048 26171
rect 1080 26139 1120 26171
rect 1152 26139 1192 26171
rect 1224 26139 1264 26171
rect 1296 26139 1336 26171
rect 1368 26139 1408 26171
rect 1440 26139 1480 26171
rect 1512 26139 1552 26171
rect 1584 26139 1624 26171
rect 1656 26139 1696 26171
rect 1728 26139 1768 26171
rect 1800 26139 1840 26171
rect 1872 26139 1912 26171
rect 1944 26139 1984 26171
rect 2016 26139 2056 26171
rect 2088 26139 2128 26171
rect 2160 26139 2200 26171
rect 2232 26139 2272 26171
rect 2304 26139 2344 26171
rect 2376 26139 2416 26171
rect 2448 26139 2488 26171
rect 2520 26139 2560 26171
rect 2592 26139 2632 26171
rect 2664 26139 2704 26171
rect 2736 26139 2776 26171
rect 2808 26139 2848 26171
rect 2880 26139 2920 26171
rect 2952 26139 2992 26171
rect 3024 26139 3064 26171
rect 3096 26139 3136 26171
rect 3168 26139 3208 26171
rect 3240 26139 3280 26171
rect 3312 26139 3352 26171
rect 3384 26139 3424 26171
rect 3456 26139 3496 26171
rect 3528 26139 3568 26171
rect 3600 26139 3640 26171
rect 3672 26139 3712 26171
rect 3744 26139 3784 26171
rect 3816 26139 3856 26171
rect 3888 26139 3950 26171
rect 50 26099 3950 26139
rect 50 26067 112 26099
rect 144 26067 184 26099
rect 216 26067 256 26099
rect 288 26067 328 26099
rect 360 26067 400 26099
rect 432 26067 472 26099
rect 504 26067 544 26099
rect 576 26067 616 26099
rect 648 26067 688 26099
rect 720 26067 760 26099
rect 792 26067 832 26099
rect 864 26067 904 26099
rect 936 26067 976 26099
rect 1008 26067 1048 26099
rect 1080 26067 1120 26099
rect 1152 26067 1192 26099
rect 1224 26067 1264 26099
rect 1296 26067 1336 26099
rect 1368 26067 1408 26099
rect 1440 26067 1480 26099
rect 1512 26067 1552 26099
rect 1584 26067 1624 26099
rect 1656 26067 1696 26099
rect 1728 26067 1768 26099
rect 1800 26067 1840 26099
rect 1872 26067 1912 26099
rect 1944 26067 1984 26099
rect 2016 26067 2056 26099
rect 2088 26067 2128 26099
rect 2160 26067 2200 26099
rect 2232 26067 2272 26099
rect 2304 26067 2344 26099
rect 2376 26067 2416 26099
rect 2448 26067 2488 26099
rect 2520 26067 2560 26099
rect 2592 26067 2632 26099
rect 2664 26067 2704 26099
rect 2736 26067 2776 26099
rect 2808 26067 2848 26099
rect 2880 26067 2920 26099
rect 2952 26067 2992 26099
rect 3024 26067 3064 26099
rect 3096 26067 3136 26099
rect 3168 26067 3208 26099
rect 3240 26067 3280 26099
rect 3312 26067 3352 26099
rect 3384 26067 3424 26099
rect 3456 26067 3496 26099
rect 3528 26067 3568 26099
rect 3600 26067 3640 26099
rect 3672 26067 3712 26099
rect 3744 26067 3784 26099
rect 3816 26067 3856 26099
rect 3888 26067 3950 26099
rect 50 26027 3950 26067
rect 50 25995 112 26027
rect 144 25995 184 26027
rect 216 25995 256 26027
rect 288 25995 328 26027
rect 360 25995 400 26027
rect 432 25995 472 26027
rect 504 25995 544 26027
rect 576 25995 616 26027
rect 648 25995 688 26027
rect 720 25995 760 26027
rect 792 25995 832 26027
rect 864 25995 904 26027
rect 936 25995 976 26027
rect 1008 25995 1048 26027
rect 1080 25995 1120 26027
rect 1152 25995 1192 26027
rect 1224 25995 1264 26027
rect 1296 25995 1336 26027
rect 1368 25995 1408 26027
rect 1440 25995 1480 26027
rect 1512 25995 1552 26027
rect 1584 25995 1624 26027
rect 1656 25995 1696 26027
rect 1728 25995 1768 26027
rect 1800 25995 1840 26027
rect 1872 25995 1912 26027
rect 1944 25995 1984 26027
rect 2016 25995 2056 26027
rect 2088 25995 2128 26027
rect 2160 25995 2200 26027
rect 2232 25995 2272 26027
rect 2304 25995 2344 26027
rect 2376 25995 2416 26027
rect 2448 25995 2488 26027
rect 2520 25995 2560 26027
rect 2592 25995 2632 26027
rect 2664 25995 2704 26027
rect 2736 25995 2776 26027
rect 2808 25995 2848 26027
rect 2880 25995 2920 26027
rect 2952 25995 2992 26027
rect 3024 25995 3064 26027
rect 3096 25995 3136 26027
rect 3168 25995 3208 26027
rect 3240 25995 3280 26027
rect 3312 25995 3352 26027
rect 3384 25995 3424 26027
rect 3456 25995 3496 26027
rect 3528 25995 3568 26027
rect 3600 25995 3640 26027
rect 3672 25995 3712 26027
rect 3744 25995 3784 26027
rect 3816 25995 3856 26027
rect 3888 25995 3950 26027
rect 50 25955 3950 25995
rect 50 25923 112 25955
rect 144 25923 184 25955
rect 216 25923 256 25955
rect 288 25923 328 25955
rect 360 25923 400 25955
rect 432 25923 472 25955
rect 504 25923 544 25955
rect 576 25923 616 25955
rect 648 25923 688 25955
rect 720 25923 760 25955
rect 792 25923 832 25955
rect 864 25923 904 25955
rect 936 25923 976 25955
rect 1008 25923 1048 25955
rect 1080 25923 1120 25955
rect 1152 25923 1192 25955
rect 1224 25923 1264 25955
rect 1296 25923 1336 25955
rect 1368 25923 1408 25955
rect 1440 25923 1480 25955
rect 1512 25923 1552 25955
rect 1584 25923 1624 25955
rect 1656 25923 1696 25955
rect 1728 25923 1768 25955
rect 1800 25923 1840 25955
rect 1872 25923 1912 25955
rect 1944 25923 1984 25955
rect 2016 25923 2056 25955
rect 2088 25923 2128 25955
rect 2160 25923 2200 25955
rect 2232 25923 2272 25955
rect 2304 25923 2344 25955
rect 2376 25923 2416 25955
rect 2448 25923 2488 25955
rect 2520 25923 2560 25955
rect 2592 25923 2632 25955
rect 2664 25923 2704 25955
rect 2736 25923 2776 25955
rect 2808 25923 2848 25955
rect 2880 25923 2920 25955
rect 2952 25923 2992 25955
rect 3024 25923 3064 25955
rect 3096 25923 3136 25955
rect 3168 25923 3208 25955
rect 3240 25923 3280 25955
rect 3312 25923 3352 25955
rect 3384 25923 3424 25955
rect 3456 25923 3496 25955
rect 3528 25923 3568 25955
rect 3600 25923 3640 25955
rect 3672 25923 3712 25955
rect 3744 25923 3784 25955
rect 3816 25923 3856 25955
rect 3888 25923 3950 25955
rect 50 25883 3950 25923
rect 50 25851 112 25883
rect 144 25851 184 25883
rect 216 25851 256 25883
rect 288 25851 328 25883
rect 360 25851 400 25883
rect 432 25851 472 25883
rect 504 25851 544 25883
rect 576 25851 616 25883
rect 648 25851 688 25883
rect 720 25851 760 25883
rect 792 25851 832 25883
rect 864 25851 904 25883
rect 936 25851 976 25883
rect 1008 25851 1048 25883
rect 1080 25851 1120 25883
rect 1152 25851 1192 25883
rect 1224 25851 1264 25883
rect 1296 25851 1336 25883
rect 1368 25851 1408 25883
rect 1440 25851 1480 25883
rect 1512 25851 1552 25883
rect 1584 25851 1624 25883
rect 1656 25851 1696 25883
rect 1728 25851 1768 25883
rect 1800 25851 1840 25883
rect 1872 25851 1912 25883
rect 1944 25851 1984 25883
rect 2016 25851 2056 25883
rect 2088 25851 2128 25883
rect 2160 25851 2200 25883
rect 2232 25851 2272 25883
rect 2304 25851 2344 25883
rect 2376 25851 2416 25883
rect 2448 25851 2488 25883
rect 2520 25851 2560 25883
rect 2592 25851 2632 25883
rect 2664 25851 2704 25883
rect 2736 25851 2776 25883
rect 2808 25851 2848 25883
rect 2880 25851 2920 25883
rect 2952 25851 2992 25883
rect 3024 25851 3064 25883
rect 3096 25851 3136 25883
rect 3168 25851 3208 25883
rect 3240 25851 3280 25883
rect 3312 25851 3352 25883
rect 3384 25851 3424 25883
rect 3456 25851 3496 25883
rect 3528 25851 3568 25883
rect 3600 25851 3640 25883
rect 3672 25851 3712 25883
rect 3744 25851 3784 25883
rect 3816 25851 3856 25883
rect 3888 25851 3950 25883
rect 50 25811 3950 25851
rect 50 25779 112 25811
rect 144 25779 184 25811
rect 216 25779 256 25811
rect 288 25779 328 25811
rect 360 25779 400 25811
rect 432 25779 472 25811
rect 504 25779 544 25811
rect 576 25779 616 25811
rect 648 25779 688 25811
rect 720 25779 760 25811
rect 792 25779 832 25811
rect 864 25779 904 25811
rect 936 25779 976 25811
rect 1008 25779 1048 25811
rect 1080 25779 1120 25811
rect 1152 25779 1192 25811
rect 1224 25779 1264 25811
rect 1296 25779 1336 25811
rect 1368 25779 1408 25811
rect 1440 25779 1480 25811
rect 1512 25779 1552 25811
rect 1584 25779 1624 25811
rect 1656 25779 1696 25811
rect 1728 25779 1768 25811
rect 1800 25779 1840 25811
rect 1872 25779 1912 25811
rect 1944 25779 1984 25811
rect 2016 25779 2056 25811
rect 2088 25779 2128 25811
rect 2160 25779 2200 25811
rect 2232 25779 2272 25811
rect 2304 25779 2344 25811
rect 2376 25779 2416 25811
rect 2448 25779 2488 25811
rect 2520 25779 2560 25811
rect 2592 25779 2632 25811
rect 2664 25779 2704 25811
rect 2736 25779 2776 25811
rect 2808 25779 2848 25811
rect 2880 25779 2920 25811
rect 2952 25779 2992 25811
rect 3024 25779 3064 25811
rect 3096 25779 3136 25811
rect 3168 25779 3208 25811
rect 3240 25779 3280 25811
rect 3312 25779 3352 25811
rect 3384 25779 3424 25811
rect 3456 25779 3496 25811
rect 3528 25779 3568 25811
rect 3600 25779 3640 25811
rect 3672 25779 3712 25811
rect 3744 25779 3784 25811
rect 3816 25779 3856 25811
rect 3888 25779 3950 25811
rect 50 25739 3950 25779
rect 50 25707 112 25739
rect 144 25707 184 25739
rect 216 25707 256 25739
rect 288 25707 328 25739
rect 360 25707 400 25739
rect 432 25707 472 25739
rect 504 25707 544 25739
rect 576 25707 616 25739
rect 648 25707 688 25739
rect 720 25707 760 25739
rect 792 25707 832 25739
rect 864 25707 904 25739
rect 936 25707 976 25739
rect 1008 25707 1048 25739
rect 1080 25707 1120 25739
rect 1152 25707 1192 25739
rect 1224 25707 1264 25739
rect 1296 25707 1336 25739
rect 1368 25707 1408 25739
rect 1440 25707 1480 25739
rect 1512 25707 1552 25739
rect 1584 25707 1624 25739
rect 1656 25707 1696 25739
rect 1728 25707 1768 25739
rect 1800 25707 1840 25739
rect 1872 25707 1912 25739
rect 1944 25707 1984 25739
rect 2016 25707 2056 25739
rect 2088 25707 2128 25739
rect 2160 25707 2200 25739
rect 2232 25707 2272 25739
rect 2304 25707 2344 25739
rect 2376 25707 2416 25739
rect 2448 25707 2488 25739
rect 2520 25707 2560 25739
rect 2592 25707 2632 25739
rect 2664 25707 2704 25739
rect 2736 25707 2776 25739
rect 2808 25707 2848 25739
rect 2880 25707 2920 25739
rect 2952 25707 2992 25739
rect 3024 25707 3064 25739
rect 3096 25707 3136 25739
rect 3168 25707 3208 25739
rect 3240 25707 3280 25739
rect 3312 25707 3352 25739
rect 3384 25707 3424 25739
rect 3456 25707 3496 25739
rect 3528 25707 3568 25739
rect 3600 25707 3640 25739
rect 3672 25707 3712 25739
rect 3744 25707 3784 25739
rect 3816 25707 3856 25739
rect 3888 25707 3950 25739
rect 50 25667 3950 25707
rect 50 25635 112 25667
rect 144 25635 184 25667
rect 216 25635 256 25667
rect 288 25635 328 25667
rect 360 25635 400 25667
rect 432 25635 472 25667
rect 504 25635 544 25667
rect 576 25635 616 25667
rect 648 25635 688 25667
rect 720 25635 760 25667
rect 792 25635 832 25667
rect 864 25635 904 25667
rect 936 25635 976 25667
rect 1008 25635 1048 25667
rect 1080 25635 1120 25667
rect 1152 25635 1192 25667
rect 1224 25635 1264 25667
rect 1296 25635 1336 25667
rect 1368 25635 1408 25667
rect 1440 25635 1480 25667
rect 1512 25635 1552 25667
rect 1584 25635 1624 25667
rect 1656 25635 1696 25667
rect 1728 25635 1768 25667
rect 1800 25635 1840 25667
rect 1872 25635 1912 25667
rect 1944 25635 1984 25667
rect 2016 25635 2056 25667
rect 2088 25635 2128 25667
rect 2160 25635 2200 25667
rect 2232 25635 2272 25667
rect 2304 25635 2344 25667
rect 2376 25635 2416 25667
rect 2448 25635 2488 25667
rect 2520 25635 2560 25667
rect 2592 25635 2632 25667
rect 2664 25635 2704 25667
rect 2736 25635 2776 25667
rect 2808 25635 2848 25667
rect 2880 25635 2920 25667
rect 2952 25635 2992 25667
rect 3024 25635 3064 25667
rect 3096 25635 3136 25667
rect 3168 25635 3208 25667
rect 3240 25635 3280 25667
rect 3312 25635 3352 25667
rect 3384 25635 3424 25667
rect 3456 25635 3496 25667
rect 3528 25635 3568 25667
rect 3600 25635 3640 25667
rect 3672 25635 3712 25667
rect 3744 25635 3784 25667
rect 3816 25635 3856 25667
rect 3888 25635 3950 25667
rect 50 25595 3950 25635
rect 50 25563 112 25595
rect 144 25563 184 25595
rect 216 25563 256 25595
rect 288 25563 328 25595
rect 360 25563 400 25595
rect 432 25563 472 25595
rect 504 25563 544 25595
rect 576 25563 616 25595
rect 648 25563 688 25595
rect 720 25563 760 25595
rect 792 25563 832 25595
rect 864 25563 904 25595
rect 936 25563 976 25595
rect 1008 25563 1048 25595
rect 1080 25563 1120 25595
rect 1152 25563 1192 25595
rect 1224 25563 1264 25595
rect 1296 25563 1336 25595
rect 1368 25563 1408 25595
rect 1440 25563 1480 25595
rect 1512 25563 1552 25595
rect 1584 25563 1624 25595
rect 1656 25563 1696 25595
rect 1728 25563 1768 25595
rect 1800 25563 1840 25595
rect 1872 25563 1912 25595
rect 1944 25563 1984 25595
rect 2016 25563 2056 25595
rect 2088 25563 2128 25595
rect 2160 25563 2200 25595
rect 2232 25563 2272 25595
rect 2304 25563 2344 25595
rect 2376 25563 2416 25595
rect 2448 25563 2488 25595
rect 2520 25563 2560 25595
rect 2592 25563 2632 25595
rect 2664 25563 2704 25595
rect 2736 25563 2776 25595
rect 2808 25563 2848 25595
rect 2880 25563 2920 25595
rect 2952 25563 2992 25595
rect 3024 25563 3064 25595
rect 3096 25563 3136 25595
rect 3168 25563 3208 25595
rect 3240 25563 3280 25595
rect 3312 25563 3352 25595
rect 3384 25563 3424 25595
rect 3456 25563 3496 25595
rect 3528 25563 3568 25595
rect 3600 25563 3640 25595
rect 3672 25563 3712 25595
rect 3744 25563 3784 25595
rect 3816 25563 3856 25595
rect 3888 25563 3950 25595
rect 50 25523 3950 25563
rect 50 25491 112 25523
rect 144 25491 184 25523
rect 216 25491 256 25523
rect 288 25491 328 25523
rect 360 25491 400 25523
rect 432 25491 472 25523
rect 504 25491 544 25523
rect 576 25491 616 25523
rect 648 25491 688 25523
rect 720 25491 760 25523
rect 792 25491 832 25523
rect 864 25491 904 25523
rect 936 25491 976 25523
rect 1008 25491 1048 25523
rect 1080 25491 1120 25523
rect 1152 25491 1192 25523
rect 1224 25491 1264 25523
rect 1296 25491 1336 25523
rect 1368 25491 1408 25523
rect 1440 25491 1480 25523
rect 1512 25491 1552 25523
rect 1584 25491 1624 25523
rect 1656 25491 1696 25523
rect 1728 25491 1768 25523
rect 1800 25491 1840 25523
rect 1872 25491 1912 25523
rect 1944 25491 1984 25523
rect 2016 25491 2056 25523
rect 2088 25491 2128 25523
rect 2160 25491 2200 25523
rect 2232 25491 2272 25523
rect 2304 25491 2344 25523
rect 2376 25491 2416 25523
rect 2448 25491 2488 25523
rect 2520 25491 2560 25523
rect 2592 25491 2632 25523
rect 2664 25491 2704 25523
rect 2736 25491 2776 25523
rect 2808 25491 2848 25523
rect 2880 25491 2920 25523
rect 2952 25491 2992 25523
rect 3024 25491 3064 25523
rect 3096 25491 3136 25523
rect 3168 25491 3208 25523
rect 3240 25491 3280 25523
rect 3312 25491 3352 25523
rect 3384 25491 3424 25523
rect 3456 25491 3496 25523
rect 3528 25491 3568 25523
rect 3600 25491 3640 25523
rect 3672 25491 3712 25523
rect 3744 25491 3784 25523
rect 3816 25491 3856 25523
rect 3888 25491 3950 25523
rect 50 25451 3950 25491
rect 50 25419 112 25451
rect 144 25419 184 25451
rect 216 25419 256 25451
rect 288 25419 328 25451
rect 360 25419 400 25451
rect 432 25419 472 25451
rect 504 25419 544 25451
rect 576 25419 616 25451
rect 648 25419 688 25451
rect 720 25419 760 25451
rect 792 25419 832 25451
rect 864 25419 904 25451
rect 936 25419 976 25451
rect 1008 25419 1048 25451
rect 1080 25419 1120 25451
rect 1152 25419 1192 25451
rect 1224 25419 1264 25451
rect 1296 25419 1336 25451
rect 1368 25419 1408 25451
rect 1440 25419 1480 25451
rect 1512 25419 1552 25451
rect 1584 25419 1624 25451
rect 1656 25419 1696 25451
rect 1728 25419 1768 25451
rect 1800 25419 1840 25451
rect 1872 25419 1912 25451
rect 1944 25419 1984 25451
rect 2016 25419 2056 25451
rect 2088 25419 2128 25451
rect 2160 25419 2200 25451
rect 2232 25419 2272 25451
rect 2304 25419 2344 25451
rect 2376 25419 2416 25451
rect 2448 25419 2488 25451
rect 2520 25419 2560 25451
rect 2592 25419 2632 25451
rect 2664 25419 2704 25451
rect 2736 25419 2776 25451
rect 2808 25419 2848 25451
rect 2880 25419 2920 25451
rect 2952 25419 2992 25451
rect 3024 25419 3064 25451
rect 3096 25419 3136 25451
rect 3168 25419 3208 25451
rect 3240 25419 3280 25451
rect 3312 25419 3352 25451
rect 3384 25419 3424 25451
rect 3456 25419 3496 25451
rect 3528 25419 3568 25451
rect 3600 25419 3640 25451
rect 3672 25419 3712 25451
rect 3744 25419 3784 25451
rect 3816 25419 3856 25451
rect 3888 25419 3950 25451
rect 50 25379 3950 25419
rect 50 25347 112 25379
rect 144 25347 184 25379
rect 216 25347 256 25379
rect 288 25347 328 25379
rect 360 25347 400 25379
rect 432 25347 472 25379
rect 504 25347 544 25379
rect 576 25347 616 25379
rect 648 25347 688 25379
rect 720 25347 760 25379
rect 792 25347 832 25379
rect 864 25347 904 25379
rect 936 25347 976 25379
rect 1008 25347 1048 25379
rect 1080 25347 1120 25379
rect 1152 25347 1192 25379
rect 1224 25347 1264 25379
rect 1296 25347 1336 25379
rect 1368 25347 1408 25379
rect 1440 25347 1480 25379
rect 1512 25347 1552 25379
rect 1584 25347 1624 25379
rect 1656 25347 1696 25379
rect 1728 25347 1768 25379
rect 1800 25347 1840 25379
rect 1872 25347 1912 25379
rect 1944 25347 1984 25379
rect 2016 25347 2056 25379
rect 2088 25347 2128 25379
rect 2160 25347 2200 25379
rect 2232 25347 2272 25379
rect 2304 25347 2344 25379
rect 2376 25347 2416 25379
rect 2448 25347 2488 25379
rect 2520 25347 2560 25379
rect 2592 25347 2632 25379
rect 2664 25347 2704 25379
rect 2736 25347 2776 25379
rect 2808 25347 2848 25379
rect 2880 25347 2920 25379
rect 2952 25347 2992 25379
rect 3024 25347 3064 25379
rect 3096 25347 3136 25379
rect 3168 25347 3208 25379
rect 3240 25347 3280 25379
rect 3312 25347 3352 25379
rect 3384 25347 3424 25379
rect 3456 25347 3496 25379
rect 3528 25347 3568 25379
rect 3600 25347 3640 25379
rect 3672 25347 3712 25379
rect 3744 25347 3784 25379
rect 3816 25347 3856 25379
rect 3888 25347 3950 25379
rect 50 25307 3950 25347
rect 50 25275 112 25307
rect 144 25275 184 25307
rect 216 25275 256 25307
rect 288 25275 328 25307
rect 360 25275 400 25307
rect 432 25275 472 25307
rect 504 25275 544 25307
rect 576 25275 616 25307
rect 648 25275 688 25307
rect 720 25275 760 25307
rect 792 25275 832 25307
rect 864 25275 904 25307
rect 936 25275 976 25307
rect 1008 25275 1048 25307
rect 1080 25275 1120 25307
rect 1152 25275 1192 25307
rect 1224 25275 1264 25307
rect 1296 25275 1336 25307
rect 1368 25275 1408 25307
rect 1440 25275 1480 25307
rect 1512 25275 1552 25307
rect 1584 25275 1624 25307
rect 1656 25275 1696 25307
rect 1728 25275 1768 25307
rect 1800 25275 1840 25307
rect 1872 25275 1912 25307
rect 1944 25275 1984 25307
rect 2016 25275 2056 25307
rect 2088 25275 2128 25307
rect 2160 25275 2200 25307
rect 2232 25275 2272 25307
rect 2304 25275 2344 25307
rect 2376 25275 2416 25307
rect 2448 25275 2488 25307
rect 2520 25275 2560 25307
rect 2592 25275 2632 25307
rect 2664 25275 2704 25307
rect 2736 25275 2776 25307
rect 2808 25275 2848 25307
rect 2880 25275 2920 25307
rect 2952 25275 2992 25307
rect 3024 25275 3064 25307
rect 3096 25275 3136 25307
rect 3168 25275 3208 25307
rect 3240 25275 3280 25307
rect 3312 25275 3352 25307
rect 3384 25275 3424 25307
rect 3456 25275 3496 25307
rect 3528 25275 3568 25307
rect 3600 25275 3640 25307
rect 3672 25275 3712 25307
rect 3744 25275 3784 25307
rect 3816 25275 3856 25307
rect 3888 25275 3950 25307
rect 50 25235 3950 25275
rect 50 25203 112 25235
rect 144 25203 184 25235
rect 216 25203 256 25235
rect 288 25203 328 25235
rect 360 25203 400 25235
rect 432 25203 472 25235
rect 504 25203 544 25235
rect 576 25203 616 25235
rect 648 25203 688 25235
rect 720 25203 760 25235
rect 792 25203 832 25235
rect 864 25203 904 25235
rect 936 25203 976 25235
rect 1008 25203 1048 25235
rect 1080 25203 1120 25235
rect 1152 25203 1192 25235
rect 1224 25203 1264 25235
rect 1296 25203 1336 25235
rect 1368 25203 1408 25235
rect 1440 25203 1480 25235
rect 1512 25203 1552 25235
rect 1584 25203 1624 25235
rect 1656 25203 1696 25235
rect 1728 25203 1768 25235
rect 1800 25203 1840 25235
rect 1872 25203 1912 25235
rect 1944 25203 1984 25235
rect 2016 25203 2056 25235
rect 2088 25203 2128 25235
rect 2160 25203 2200 25235
rect 2232 25203 2272 25235
rect 2304 25203 2344 25235
rect 2376 25203 2416 25235
rect 2448 25203 2488 25235
rect 2520 25203 2560 25235
rect 2592 25203 2632 25235
rect 2664 25203 2704 25235
rect 2736 25203 2776 25235
rect 2808 25203 2848 25235
rect 2880 25203 2920 25235
rect 2952 25203 2992 25235
rect 3024 25203 3064 25235
rect 3096 25203 3136 25235
rect 3168 25203 3208 25235
rect 3240 25203 3280 25235
rect 3312 25203 3352 25235
rect 3384 25203 3424 25235
rect 3456 25203 3496 25235
rect 3528 25203 3568 25235
rect 3600 25203 3640 25235
rect 3672 25203 3712 25235
rect 3744 25203 3784 25235
rect 3816 25203 3856 25235
rect 3888 25203 3950 25235
rect 50 25163 3950 25203
rect 50 25131 112 25163
rect 144 25131 184 25163
rect 216 25131 256 25163
rect 288 25131 328 25163
rect 360 25131 400 25163
rect 432 25131 472 25163
rect 504 25131 544 25163
rect 576 25131 616 25163
rect 648 25131 688 25163
rect 720 25131 760 25163
rect 792 25131 832 25163
rect 864 25131 904 25163
rect 936 25131 976 25163
rect 1008 25131 1048 25163
rect 1080 25131 1120 25163
rect 1152 25131 1192 25163
rect 1224 25131 1264 25163
rect 1296 25131 1336 25163
rect 1368 25131 1408 25163
rect 1440 25131 1480 25163
rect 1512 25131 1552 25163
rect 1584 25131 1624 25163
rect 1656 25131 1696 25163
rect 1728 25131 1768 25163
rect 1800 25131 1840 25163
rect 1872 25131 1912 25163
rect 1944 25131 1984 25163
rect 2016 25131 2056 25163
rect 2088 25131 2128 25163
rect 2160 25131 2200 25163
rect 2232 25131 2272 25163
rect 2304 25131 2344 25163
rect 2376 25131 2416 25163
rect 2448 25131 2488 25163
rect 2520 25131 2560 25163
rect 2592 25131 2632 25163
rect 2664 25131 2704 25163
rect 2736 25131 2776 25163
rect 2808 25131 2848 25163
rect 2880 25131 2920 25163
rect 2952 25131 2992 25163
rect 3024 25131 3064 25163
rect 3096 25131 3136 25163
rect 3168 25131 3208 25163
rect 3240 25131 3280 25163
rect 3312 25131 3352 25163
rect 3384 25131 3424 25163
rect 3456 25131 3496 25163
rect 3528 25131 3568 25163
rect 3600 25131 3640 25163
rect 3672 25131 3712 25163
rect 3744 25131 3784 25163
rect 3816 25131 3856 25163
rect 3888 25131 3950 25163
rect 50 25091 3950 25131
rect 50 25059 112 25091
rect 144 25059 184 25091
rect 216 25059 256 25091
rect 288 25059 328 25091
rect 360 25059 400 25091
rect 432 25059 472 25091
rect 504 25059 544 25091
rect 576 25059 616 25091
rect 648 25059 688 25091
rect 720 25059 760 25091
rect 792 25059 832 25091
rect 864 25059 904 25091
rect 936 25059 976 25091
rect 1008 25059 1048 25091
rect 1080 25059 1120 25091
rect 1152 25059 1192 25091
rect 1224 25059 1264 25091
rect 1296 25059 1336 25091
rect 1368 25059 1408 25091
rect 1440 25059 1480 25091
rect 1512 25059 1552 25091
rect 1584 25059 1624 25091
rect 1656 25059 1696 25091
rect 1728 25059 1768 25091
rect 1800 25059 1840 25091
rect 1872 25059 1912 25091
rect 1944 25059 1984 25091
rect 2016 25059 2056 25091
rect 2088 25059 2128 25091
rect 2160 25059 2200 25091
rect 2232 25059 2272 25091
rect 2304 25059 2344 25091
rect 2376 25059 2416 25091
rect 2448 25059 2488 25091
rect 2520 25059 2560 25091
rect 2592 25059 2632 25091
rect 2664 25059 2704 25091
rect 2736 25059 2776 25091
rect 2808 25059 2848 25091
rect 2880 25059 2920 25091
rect 2952 25059 2992 25091
rect 3024 25059 3064 25091
rect 3096 25059 3136 25091
rect 3168 25059 3208 25091
rect 3240 25059 3280 25091
rect 3312 25059 3352 25091
rect 3384 25059 3424 25091
rect 3456 25059 3496 25091
rect 3528 25059 3568 25091
rect 3600 25059 3640 25091
rect 3672 25059 3712 25091
rect 3744 25059 3784 25091
rect 3816 25059 3856 25091
rect 3888 25059 3950 25091
rect 50 25019 3950 25059
rect 50 24987 112 25019
rect 144 24987 184 25019
rect 216 24987 256 25019
rect 288 24987 328 25019
rect 360 24987 400 25019
rect 432 24987 472 25019
rect 504 24987 544 25019
rect 576 24987 616 25019
rect 648 24987 688 25019
rect 720 24987 760 25019
rect 792 24987 832 25019
rect 864 24987 904 25019
rect 936 24987 976 25019
rect 1008 24987 1048 25019
rect 1080 24987 1120 25019
rect 1152 24987 1192 25019
rect 1224 24987 1264 25019
rect 1296 24987 1336 25019
rect 1368 24987 1408 25019
rect 1440 24987 1480 25019
rect 1512 24987 1552 25019
rect 1584 24987 1624 25019
rect 1656 24987 1696 25019
rect 1728 24987 1768 25019
rect 1800 24987 1840 25019
rect 1872 24987 1912 25019
rect 1944 24987 1984 25019
rect 2016 24987 2056 25019
rect 2088 24987 2128 25019
rect 2160 24987 2200 25019
rect 2232 24987 2272 25019
rect 2304 24987 2344 25019
rect 2376 24987 2416 25019
rect 2448 24987 2488 25019
rect 2520 24987 2560 25019
rect 2592 24987 2632 25019
rect 2664 24987 2704 25019
rect 2736 24987 2776 25019
rect 2808 24987 2848 25019
rect 2880 24987 2920 25019
rect 2952 24987 2992 25019
rect 3024 24987 3064 25019
rect 3096 24987 3136 25019
rect 3168 24987 3208 25019
rect 3240 24987 3280 25019
rect 3312 24987 3352 25019
rect 3384 24987 3424 25019
rect 3456 24987 3496 25019
rect 3528 24987 3568 25019
rect 3600 24987 3640 25019
rect 3672 24987 3712 25019
rect 3744 24987 3784 25019
rect 3816 24987 3856 25019
rect 3888 24987 3950 25019
rect 50 24947 3950 24987
rect 50 24915 112 24947
rect 144 24915 184 24947
rect 216 24915 256 24947
rect 288 24915 328 24947
rect 360 24915 400 24947
rect 432 24915 472 24947
rect 504 24915 544 24947
rect 576 24915 616 24947
rect 648 24915 688 24947
rect 720 24915 760 24947
rect 792 24915 832 24947
rect 864 24915 904 24947
rect 936 24915 976 24947
rect 1008 24915 1048 24947
rect 1080 24915 1120 24947
rect 1152 24915 1192 24947
rect 1224 24915 1264 24947
rect 1296 24915 1336 24947
rect 1368 24915 1408 24947
rect 1440 24915 1480 24947
rect 1512 24915 1552 24947
rect 1584 24915 1624 24947
rect 1656 24915 1696 24947
rect 1728 24915 1768 24947
rect 1800 24915 1840 24947
rect 1872 24915 1912 24947
rect 1944 24915 1984 24947
rect 2016 24915 2056 24947
rect 2088 24915 2128 24947
rect 2160 24915 2200 24947
rect 2232 24915 2272 24947
rect 2304 24915 2344 24947
rect 2376 24915 2416 24947
rect 2448 24915 2488 24947
rect 2520 24915 2560 24947
rect 2592 24915 2632 24947
rect 2664 24915 2704 24947
rect 2736 24915 2776 24947
rect 2808 24915 2848 24947
rect 2880 24915 2920 24947
rect 2952 24915 2992 24947
rect 3024 24915 3064 24947
rect 3096 24915 3136 24947
rect 3168 24915 3208 24947
rect 3240 24915 3280 24947
rect 3312 24915 3352 24947
rect 3384 24915 3424 24947
rect 3456 24915 3496 24947
rect 3528 24915 3568 24947
rect 3600 24915 3640 24947
rect 3672 24915 3712 24947
rect 3744 24915 3784 24947
rect 3816 24915 3856 24947
rect 3888 24915 3950 24947
rect 50 24875 3950 24915
rect 50 24843 112 24875
rect 144 24843 184 24875
rect 216 24843 256 24875
rect 288 24843 328 24875
rect 360 24843 400 24875
rect 432 24843 472 24875
rect 504 24843 544 24875
rect 576 24843 616 24875
rect 648 24843 688 24875
rect 720 24843 760 24875
rect 792 24843 832 24875
rect 864 24843 904 24875
rect 936 24843 976 24875
rect 1008 24843 1048 24875
rect 1080 24843 1120 24875
rect 1152 24843 1192 24875
rect 1224 24843 1264 24875
rect 1296 24843 1336 24875
rect 1368 24843 1408 24875
rect 1440 24843 1480 24875
rect 1512 24843 1552 24875
rect 1584 24843 1624 24875
rect 1656 24843 1696 24875
rect 1728 24843 1768 24875
rect 1800 24843 1840 24875
rect 1872 24843 1912 24875
rect 1944 24843 1984 24875
rect 2016 24843 2056 24875
rect 2088 24843 2128 24875
rect 2160 24843 2200 24875
rect 2232 24843 2272 24875
rect 2304 24843 2344 24875
rect 2376 24843 2416 24875
rect 2448 24843 2488 24875
rect 2520 24843 2560 24875
rect 2592 24843 2632 24875
rect 2664 24843 2704 24875
rect 2736 24843 2776 24875
rect 2808 24843 2848 24875
rect 2880 24843 2920 24875
rect 2952 24843 2992 24875
rect 3024 24843 3064 24875
rect 3096 24843 3136 24875
rect 3168 24843 3208 24875
rect 3240 24843 3280 24875
rect 3312 24843 3352 24875
rect 3384 24843 3424 24875
rect 3456 24843 3496 24875
rect 3528 24843 3568 24875
rect 3600 24843 3640 24875
rect 3672 24843 3712 24875
rect 3744 24843 3784 24875
rect 3816 24843 3856 24875
rect 3888 24843 3950 24875
rect 50 24803 3950 24843
rect 50 24771 112 24803
rect 144 24771 184 24803
rect 216 24771 256 24803
rect 288 24771 328 24803
rect 360 24771 400 24803
rect 432 24771 472 24803
rect 504 24771 544 24803
rect 576 24771 616 24803
rect 648 24771 688 24803
rect 720 24771 760 24803
rect 792 24771 832 24803
rect 864 24771 904 24803
rect 936 24771 976 24803
rect 1008 24771 1048 24803
rect 1080 24771 1120 24803
rect 1152 24771 1192 24803
rect 1224 24771 1264 24803
rect 1296 24771 1336 24803
rect 1368 24771 1408 24803
rect 1440 24771 1480 24803
rect 1512 24771 1552 24803
rect 1584 24771 1624 24803
rect 1656 24771 1696 24803
rect 1728 24771 1768 24803
rect 1800 24771 1840 24803
rect 1872 24771 1912 24803
rect 1944 24771 1984 24803
rect 2016 24771 2056 24803
rect 2088 24771 2128 24803
rect 2160 24771 2200 24803
rect 2232 24771 2272 24803
rect 2304 24771 2344 24803
rect 2376 24771 2416 24803
rect 2448 24771 2488 24803
rect 2520 24771 2560 24803
rect 2592 24771 2632 24803
rect 2664 24771 2704 24803
rect 2736 24771 2776 24803
rect 2808 24771 2848 24803
rect 2880 24771 2920 24803
rect 2952 24771 2992 24803
rect 3024 24771 3064 24803
rect 3096 24771 3136 24803
rect 3168 24771 3208 24803
rect 3240 24771 3280 24803
rect 3312 24771 3352 24803
rect 3384 24771 3424 24803
rect 3456 24771 3496 24803
rect 3528 24771 3568 24803
rect 3600 24771 3640 24803
rect 3672 24771 3712 24803
rect 3744 24771 3784 24803
rect 3816 24771 3856 24803
rect 3888 24771 3950 24803
rect 50 24731 3950 24771
rect 50 24699 112 24731
rect 144 24699 184 24731
rect 216 24699 256 24731
rect 288 24699 328 24731
rect 360 24699 400 24731
rect 432 24699 472 24731
rect 504 24699 544 24731
rect 576 24699 616 24731
rect 648 24699 688 24731
rect 720 24699 760 24731
rect 792 24699 832 24731
rect 864 24699 904 24731
rect 936 24699 976 24731
rect 1008 24699 1048 24731
rect 1080 24699 1120 24731
rect 1152 24699 1192 24731
rect 1224 24699 1264 24731
rect 1296 24699 1336 24731
rect 1368 24699 1408 24731
rect 1440 24699 1480 24731
rect 1512 24699 1552 24731
rect 1584 24699 1624 24731
rect 1656 24699 1696 24731
rect 1728 24699 1768 24731
rect 1800 24699 1840 24731
rect 1872 24699 1912 24731
rect 1944 24699 1984 24731
rect 2016 24699 2056 24731
rect 2088 24699 2128 24731
rect 2160 24699 2200 24731
rect 2232 24699 2272 24731
rect 2304 24699 2344 24731
rect 2376 24699 2416 24731
rect 2448 24699 2488 24731
rect 2520 24699 2560 24731
rect 2592 24699 2632 24731
rect 2664 24699 2704 24731
rect 2736 24699 2776 24731
rect 2808 24699 2848 24731
rect 2880 24699 2920 24731
rect 2952 24699 2992 24731
rect 3024 24699 3064 24731
rect 3096 24699 3136 24731
rect 3168 24699 3208 24731
rect 3240 24699 3280 24731
rect 3312 24699 3352 24731
rect 3384 24699 3424 24731
rect 3456 24699 3496 24731
rect 3528 24699 3568 24731
rect 3600 24699 3640 24731
rect 3672 24699 3712 24731
rect 3744 24699 3784 24731
rect 3816 24699 3856 24731
rect 3888 24699 3950 24731
rect 50 24659 3950 24699
rect 50 24627 112 24659
rect 144 24627 184 24659
rect 216 24627 256 24659
rect 288 24627 328 24659
rect 360 24627 400 24659
rect 432 24627 472 24659
rect 504 24627 544 24659
rect 576 24627 616 24659
rect 648 24627 688 24659
rect 720 24627 760 24659
rect 792 24627 832 24659
rect 864 24627 904 24659
rect 936 24627 976 24659
rect 1008 24627 1048 24659
rect 1080 24627 1120 24659
rect 1152 24627 1192 24659
rect 1224 24627 1264 24659
rect 1296 24627 1336 24659
rect 1368 24627 1408 24659
rect 1440 24627 1480 24659
rect 1512 24627 1552 24659
rect 1584 24627 1624 24659
rect 1656 24627 1696 24659
rect 1728 24627 1768 24659
rect 1800 24627 1840 24659
rect 1872 24627 1912 24659
rect 1944 24627 1984 24659
rect 2016 24627 2056 24659
rect 2088 24627 2128 24659
rect 2160 24627 2200 24659
rect 2232 24627 2272 24659
rect 2304 24627 2344 24659
rect 2376 24627 2416 24659
rect 2448 24627 2488 24659
rect 2520 24627 2560 24659
rect 2592 24627 2632 24659
rect 2664 24627 2704 24659
rect 2736 24627 2776 24659
rect 2808 24627 2848 24659
rect 2880 24627 2920 24659
rect 2952 24627 2992 24659
rect 3024 24627 3064 24659
rect 3096 24627 3136 24659
rect 3168 24627 3208 24659
rect 3240 24627 3280 24659
rect 3312 24627 3352 24659
rect 3384 24627 3424 24659
rect 3456 24627 3496 24659
rect 3528 24627 3568 24659
rect 3600 24627 3640 24659
rect 3672 24627 3712 24659
rect 3744 24627 3784 24659
rect 3816 24627 3856 24659
rect 3888 24627 3950 24659
rect 50 24587 3950 24627
rect 50 24555 112 24587
rect 144 24555 184 24587
rect 216 24555 256 24587
rect 288 24555 328 24587
rect 360 24555 400 24587
rect 432 24555 472 24587
rect 504 24555 544 24587
rect 576 24555 616 24587
rect 648 24555 688 24587
rect 720 24555 760 24587
rect 792 24555 832 24587
rect 864 24555 904 24587
rect 936 24555 976 24587
rect 1008 24555 1048 24587
rect 1080 24555 1120 24587
rect 1152 24555 1192 24587
rect 1224 24555 1264 24587
rect 1296 24555 1336 24587
rect 1368 24555 1408 24587
rect 1440 24555 1480 24587
rect 1512 24555 1552 24587
rect 1584 24555 1624 24587
rect 1656 24555 1696 24587
rect 1728 24555 1768 24587
rect 1800 24555 1840 24587
rect 1872 24555 1912 24587
rect 1944 24555 1984 24587
rect 2016 24555 2056 24587
rect 2088 24555 2128 24587
rect 2160 24555 2200 24587
rect 2232 24555 2272 24587
rect 2304 24555 2344 24587
rect 2376 24555 2416 24587
rect 2448 24555 2488 24587
rect 2520 24555 2560 24587
rect 2592 24555 2632 24587
rect 2664 24555 2704 24587
rect 2736 24555 2776 24587
rect 2808 24555 2848 24587
rect 2880 24555 2920 24587
rect 2952 24555 2992 24587
rect 3024 24555 3064 24587
rect 3096 24555 3136 24587
rect 3168 24555 3208 24587
rect 3240 24555 3280 24587
rect 3312 24555 3352 24587
rect 3384 24555 3424 24587
rect 3456 24555 3496 24587
rect 3528 24555 3568 24587
rect 3600 24555 3640 24587
rect 3672 24555 3712 24587
rect 3744 24555 3784 24587
rect 3816 24555 3856 24587
rect 3888 24555 3950 24587
rect 50 24515 3950 24555
rect 50 24483 112 24515
rect 144 24483 184 24515
rect 216 24483 256 24515
rect 288 24483 328 24515
rect 360 24483 400 24515
rect 432 24483 472 24515
rect 504 24483 544 24515
rect 576 24483 616 24515
rect 648 24483 688 24515
rect 720 24483 760 24515
rect 792 24483 832 24515
rect 864 24483 904 24515
rect 936 24483 976 24515
rect 1008 24483 1048 24515
rect 1080 24483 1120 24515
rect 1152 24483 1192 24515
rect 1224 24483 1264 24515
rect 1296 24483 1336 24515
rect 1368 24483 1408 24515
rect 1440 24483 1480 24515
rect 1512 24483 1552 24515
rect 1584 24483 1624 24515
rect 1656 24483 1696 24515
rect 1728 24483 1768 24515
rect 1800 24483 1840 24515
rect 1872 24483 1912 24515
rect 1944 24483 1984 24515
rect 2016 24483 2056 24515
rect 2088 24483 2128 24515
rect 2160 24483 2200 24515
rect 2232 24483 2272 24515
rect 2304 24483 2344 24515
rect 2376 24483 2416 24515
rect 2448 24483 2488 24515
rect 2520 24483 2560 24515
rect 2592 24483 2632 24515
rect 2664 24483 2704 24515
rect 2736 24483 2776 24515
rect 2808 24483 2848 24515
rect 2880 24483 2920 24515
rect 2952 24483 2992 24515
rect 3024 24483 3064 24515
rect 3096 24483 3136 24515
rect 3168 24483 3208 24515
rect 3240 24483 3280 24515
rect 3312 24483 3352 24515
rect 3384 24483 3424 24515
rect 3456 24483 3496 24515
rect 3528 24483 3568 24515
rect 3600 24483 3640 24515
rect 3672 24483 3712 24515
rect 3744 24483 3784 24515
rect 3816 24483 3856 24515
rect 3888 24483 3950 24515
rect 50 24443 3950 24483
rect 50 24411 112 24443
rect 144 24411 184 24443
rect 216 24411 256 24443
rect 288 24411 328 24443
rect 360 24411 400 24443
rect 432 24411 472 24443
rect 504 24411 544 24443
rect 576 24411 616 24443
rect 648 24411 688 24443
rect 720 24411 760 24443
rect 792 24411 832 24443
rect 864 24411 904 24443
rect 936 24411 976 24443
rect 1008 24411 1048 24443
rect 1080 24411 1120 24443
rect 1152 24411 1192 24443
rect 1224 24411 1264 24443
rect 1296 24411 1336 24443
rect 1368 24411 1408 24443
rect 1440 24411 1480 24443
rect 1512 24411 1552 24443
rect 1584 24411 1624 24443
rect 1656 24411 1696 24443
rect 1728 24411 1768 24443
rect 1800 24411 1840 24443
rect 1872 24411 1912 24443
rect 1944 24411 1984 24443
rect 2016 24411 2056 24443
rect 2088 24411 2128 24443
rect 2160 24411 2200 24443
rect 2232 24411 2272 24443
rect 2304 24411 2344 24443
rect 2376 24411 2416 24443
rect 2448 24411 2488 24443
rect 2520 24411 2560 24443
rect 2592 24411 2632 24443
rect 2664 24411 2704 24443
rect 2736 24411 2776 24443
rect 2808 24411 2848 24443
rect 2880 24411 2920 24443
rect 2952 24411 2992 24443
rect 3024 24411 3064 24443
rect 3096 24411 3136 24443
rect 3168 24411 3208 24443
rect 3240 24411 3280 24443
rect 3312 24411 3352 24443
rect 3384 24411 3424 24443
rect 3456 24411 3496 24443
rect 3528 24411 3568 24443
rect 3600 24411 3640 24443
rect 3672 24411 3712 24443
rect 3744 24411 3784 24443
rect 3816 24411 3856 24443
rect 3888 24411 3950 24443
rect 50 24371 3950 24411
rect 50 24339 112 24371
rect 144 24339 184 24371
rect 216 24339 256 24371
rect 288 24339 328 24371
rect 360 24339 400 24371
rect 432 24339 472 24371
rect 504 24339 544 24371
rect 576 24339 616 24371
rect 648 24339 688 24371
rect 720 24339 760 24371
rect 792 24339 832 24371
rect 864 24339 904 24371
rect 936 24339 976 24371
rect 1008 24339 1048 24371
rect 1080 24339 1120 24371
rect 1152 24339 1192 24371
rect 1224 24339 1264 24371
rect 1296 24339 1336 24371
rect 1368 24339 1408 24371
rect 1440 24339 1480 24371
rect 1512 24339 1552 24371
rect 1584 24339 1624 24371
rect 1656 24339 1696 24371
rect 1728 24339 1768 24371
rect 1800 24339 1840 24371
rect 1872 24339 1912 24371
rect 1944 24339 1984 24371
rect 2016 24339 2056 24371
rect 2088 24339 2128 24371
rect 2160 24339 2200 24371
rect 2232 24339 2272 24371
rect 2304 24339 2344 24371
rect 2376 24339 2416 24371
rect 2448 24339 2488 24371
rect 2520 24339 2560 24371
rect 2592 24339 2632 24371
rect 2664 24339 2704 24371
rect 2736 24339 2776 24371
rect 2808 24339 2848 24371
rect 2880 24339 2920 24371
rect 2952 24339 2992 24371
rect 3024 24339 3064 24371
rect 3096 24339 3136 24371
rect 3168 24339 3208 24371
rect 3240 24339 3280 24371
rect 3312 24339 3352 24371
rect 3384 24339 3424 24371
rect 3456 24339 3496 24371
rect 3528 24339 3568 24371
rect 3600 24339 3640 24371
rect 3672 24339 3712 24371
rect 3744 24339 3784 24371
rect 3816 24339 3856 24371
rect 3888 24339 3950 24371
rect 50 24299 3950 24339
rect 50 24267 112 24299
rect 144 24267 184 24299
rect 216 24267 256 24299
rect 288 24267 328 24299
rect 360 24267 400 24299
rect 432 24267 472 24299
rect 504 24267 544 24299
rect 576 24267 616 24299
rect 648 24267 688 24299
rect 720 24267 760 24299
rect 792 24267 832 24299
rect 864 24267 904 24299
rect 936 24267 976 24299
rect 1008 24267 1048 24299
rect 1080 24267 1120 24299
rect 1152 24267 1192 24299
rect 1224 24267 1264 24299
rect 1296 24267 1336 24299
rect 1368 24267 1408 24299
rect 1440 24267 1480 24299
rect 1512 24267 1552 24299
rect 1584 24267 1624 24299
rect 1656 24267 1696 24299
rect 1728 24267 1768 24299
rect 1800 24267 1840 24299
rect 1872 24267 1912 24299
rect 1944 24267 1984 24299
rect 2016 24267 2056 24299
rect 2088 24267 2128 24299
rect 2160 24267 2200 24299
rect 2232 24267 2272 24299
rect 2304 24267 2344 24299
rect 2376 24267 2416 24299
rect 2448 24267 2488 24299
rect 2520 24267 2560 24299
rect 2592 24267 2632 24299
rect 2664 24267 2704 24299
rect 2736 24267 2776 24299
rect 2808 24267 2848 24299
rect 2880 24267 2920 24299
rect 2952 24267 2992 24299
rect 3024 24267 3064 24299
rect 3096 24267 3136 24299
rect 3168 24267 3208 24299
rect 3240 24267 3280 24299
rect 3312 24267 3352 24299
rect 3384 24267 3424 24299
rect 3456 24267 3496 24299
rect 3528 24267 3568 24299
rect 3600 24267 3640 24299
rect 3672 24267 3712 24299
rect 3744 24267 3784 24299
rect 3816 24267 3856 24299
rect 3888 24267 3950 24299
rect 50 24227 3950 24267
rect 50 24195 112 24227
rect 144 24195 184 24227
rect 216 24195 256 24227
rect 288 24195 328 24227
rect 360 24195 400 24227
rect 432 24195 472 24227
rect 504 24195 544 24227
rect 576 24195 616 24227
rect 648 24195 688 24227
rect 720 24195 760 24227
rect 792 24195 832 24227
rect 864 24195 904 24227
rect 936 24195 976 24227
rect 1008 24195 1048 24227
rect 1080 24195 1120 24227
rect 1152 24195 1192 24227
rect 1224 24195 1264 24227
rect 1296 24195 1336 24227
rect 1368 24195 1408 24227
rect 1440 24195 1480 24227
rect 1512 24195 1552 24227
rect 1584 24195 1624 24227
rect 1656 24195 1696 24227
rect 1728 24195 1768 24227
rect 1800 24195 1840 24227
rect 1872 24195 1912 24227
rect 1944 24195 1984 24227
rect 2016 24195 2056 24227
rect 2088 24195 2128 24227
rect 2160 24195 2200 24227
rect 2232 24195 2272 24227
rect 2304 24195 2344 24227
rect 2376 24195 2416 24227
rect 2448 24195 2488 24227
rect 2520 24195 2560 24227
rect 2592 24195 2632 24227
rect 2664 24195 2704 24227
rect 2736 24195 2776 24227
rect 2808 24195 2848 24227
rect 2880 24195 2920 24227
rect 2952 24195 2992 24227
rect 3024 24195 3064 24227
rect 3096 24195 3136 24227
rect 3168 24195 3208 24227
rect 3240 24195 3280 24227
rect 3312 24195 3352 24227
rect 3384 24195 3424 24227
rect 3456 24195 3496 24227
rect 3528 24195 3568 24227
rect 3600 24195 3640 24227
rect 3672 24195 3712 24227
rect 3744 24195 3784 24227
rect 3816 24195 3856 24227
rect 3888 24195 3950 24227
rect 50 24155 3950 24195
rect 50 24123 112 24155
rect 144 24123 184 24155
rect 216 24123 256 24155
rect 288 24123 328 24155
rect 360 24123 400 24155
rect 432 24123 472 24155
rect 504 24123 544 24155
rect 576 24123 616 24155
rect 648 24123 688 24155
rect 720 24123 760 24155
rect 792 24123 832 24155
rect 864 24123 904 24155
rect 936 24123 976 24155
rect 1008 24123 1048 24155
rect 1080 24123 1120 24155
rect 1152 24123 1192 24155
rect 1224 24123 1264 24155
rect 1296 24123 1336 24155
rect 1368 24123 1408 24155
rect 1440 24123 1480 24155
rect 1512 24123 1552 24155
rect 1584 24123 1624 24155
rect 1656 24123 1696 24155
rect 1728 24123 1768 24155
rect 1800 24123 1840 24155
rect 1872 24123 1912 24155
rect 1944 24123 1984 24155
rect 2016 24123 2056 24155
rect 2088 24123 2128 24155
rect 2160 24123 2200 24155
rect 2232 24123 2272 24155
rect 2304 24123 2344 24155
rect 2376 24123 2416 24155
rect 2448 24123 2488 24155
rect 2520 24123 2560 24155
rect 2592 24123 2632 24155
rect 2664 24123 2704 24155
rect 2736 24123 2776 24155
rect 2808 24123 2848 24155
rect 2880 24123 2920 24155
rect 2952 24123 2992 24155
rect 3024 24123 3064 24155
rect 3096 24123 3136 24155
rect 3168 24123 3208 24155
rect 3240 24123 3280 24155
rect 3312 24123 3352 24155
rect 3384 24123 3424 24155
rect 3456 24123 3496 24155
rect 3528 24123 3568 24155
rect 3600 24123 3640 24155
rect 3672 24123 3712 24155
rect 3744 24123 3784 24155
rect 3816 24123 3856 24155
rect 3888 24123 3950 24155
rect 50 24083 3950 24123
rect 50 24051 112 24083
rect 144 24051 184 24083
rect 216 24051 256 24083
rect 288 24051 328 24083
rect 360 24051 400 24083
rect 432 24051 472 24083
rect 504 24051 544 24083
rect 576 24051 616 24083
rect 648 24051 688 24083
rect 720 24051 760 24083
rect 792 24051 832 24083
rect 864 24051 904 24083
rect 936 24051 976 24083
rect 1008 24051 1048 24083
rect 1080 24051 1120 24083
rect 1152 24051 1192 24083
rect 1224 24051 1264 24083
rect 1296 24051 1336 24083
rect 1368 24051 1408 24083
rect 1440 24051 1480 24083
rect 1512 24051 1552 24083
rect 1584 24051 1624 24083
rect 1656 24051 1696 24083
rect 1728 24051 1768 24083
rect 1800 24051 1840 24083
rect 1872 24051 1912 24083
rect 1944 24051 1984 24083
rect 2016 24051 2056 24083
rect 2088 24051 2128 24083
rect 2160 24051 2200 24083
rect 2232 24051 2272 24083
rect 2304 24051 2344 24083
rect 2376 24051 2416 24083
rect 2448 24051 2488 24083
rect 2520 24051 2560 24083
rect 2592 24051 2632 24083
rect 2664 24051 2704 24083
rect 2736 24051 2776 24083
rect 2808 24051 2848 24083
rect 2880 24051 2920 24083
rect 2952 24051 2992 24083
rect 3024 24051 3064 24083
rect 3096 24051 3136 24083
rect 3168 24051 3208 24083
rect 3240 24051 3280 24083
rect 3312 24051 3352 24083
rect 3384 24051 3424 24083
rect 3456 24051 3496 24083
rect 3528 24051 3568 24083
rect 3600 24051 3640 24083
rect 3672 24051 3712 24083
rect 3744 24051 3784 24083
rect 3816 24051 3856 24083
rect 3888 24051 3950 24083
rect 50 24011 3950 24051
rect 50 23979 112 24011
rect 144 23979 184 24011
rect 216 23979 256 24011
rect 288 23979 328 24011
rect 360 23979 400 24011
rect 432 23979 472 24011
rect 504 23979 544 24011
rect 576 23979 616 24011
rect 648 23979 688 24011
rect 720 23979 760 24011
rect 792 23979 832 24011
rect 864 23979 904 24011
rect 936 23979 976 24011
rect 1008 23979 1048 24011
rect 1080 23979 1120 24011
rect 1152 23979 1192 24011
rect 1224 23979 1264 24011
rect 1296 23979 1336 24011
rect 1368 23979 1408 24011
rect 1440 23979 1480 24011
rect 1512 23979 1552 24011
rect 1584 23979 1624 24011
rect 1656 23979 1696 24011
rect 1728 23979 1768 24011
rect 1800 23979 1840 24011
rect 1872 23979 1912 24011
rect 1944 23979 1984 24011
rect 2016 23979 2056 24011
rect 2088 23979 2128 24011
rect 2160 23979 2200 24011
rect 2232 23979 2272 24011
rect 2304 23979 2344 24011
rect 2376 23979 2416 24011
rect 2448 23979 2488 24011
rect 2520 23979 2560 24011
rect 2592 23979 2632 24011
rect 2664 23979 2704 24011
rect 2736 23979 2776 24011
rect 2808 23979 2848 24011
rect 2880 23979 2920 24011
rect 2952 23979 2992 24011
rect 3024 23979 3064 24011
rect 3096 23979 3136 24011
rect 3168 23979 3208 24011
rect 3240 23979 3280 24011
rect 3312 23979 3352 24011
rect 3384 23979 3424 24011
rect 3456 23979 3496 24011
rect 3528 23979 3568 24011
rect 3600 23979 3640 24011
rect 3672 23979 3712 24011
rect 3744 23979 3784 24011
rect 3816 23979 3856 24011
rect 3888 23979 3950 24011
rect 50 23939 3950 23979
rect 50 23907 112 23939
rect 144 23907 184 23939
rect 216 23907 256 23939
rect 288 23907 328 23939
rect 360 23907 400 23939
rect 432 23907 472 23939
rect 504 23907 544 23939
rect 576 23907 616 23939
rect 648 23907 688 23939
rect 720 23907 760 23939
rect 792 23907 832 23939
rect 864 23907 904 23939
rect 936 23907 976 23939
rect 1008 23907 1048 23939
rect 1080 23907 1120 23939
rect 1152 23907 1192 23939
rect 1224 23907 1264 23939
rect 1296 23907 1336 23939
rect 1368 23907 1408 23939
rect 1440 23907 1480 23939
rect 1512 23907 1552 23939
rect 1584 23907 1624 23939
rect 1656 23907 1696 23939
rect 1728 23907 1768 23939
rect 1800 23907 1840 23939
rect 1872 23907 1912 23939
rect 1944 23907 1984 23939
rect 2016 23907 2056 23939
rect 2088 23907 2128 23939
rect 2160 23907 2200 23939
rect 2232 23907 2272 23939
rect 2304 23907 2344 23939
rect 2376 23907 2416 23939
rect 2448 23907 2488 23939
rect 2520 23907 2560 23939
rect 2592 23907 2632 23939
rect 2664 23907 2704 23939
rect 2736 23907 2776 23939
rect 2808 23907 2848 23939
rect 2880 23907 2920 23939
rect 2952 23907 2992 23939
rect 3024 23907 3064 23939
rect 3096 23907 3136 23939
rect 3168 23907 3208 23939
rect 3240 23907 3280 23939
rect 3312 23907 3352 23939
rect 3384 23907 3424 23939
rect 3456 23907 3496 23939
rect 3528 23907 3568 23939
rect 3600 23907 3640 23939
rect 3672 23907 3712 23939
rect 3744 23907 3784 23939
rect 3816 23907 3856 23939
rect 3888 23907 3950 23939
rect 50 23867 3950 23907
rect 50 23835 112 23867
rect 144 23835 184 23867
rect 216 23835 256 23867
rect 288 23835 328 23867
rect 360 23835 400 23867
rect 432 23835 472 23867
rect 504 23835 544 23867
rect 576 23835 616 23867
rect 648 23835 688 23867
rect 720 23835 760 23867
rect 792 23835 832 23867
rect 864 23835 904 23867
rect 936 23835 976 23867
rect 1008 23835 1048 23867
rect 1080 23835 1120 23867
rect 1152 23835 1192 23867
rect 1224 23835 1264 23867
rect 1296 23835 1336 23867
rect 1368 23835 1408 23867
rect 1440 23835 1480 23867
rect 1512 23835 1552 23867
rect 1584 23835 1624 23867
rect 1656 23835 1696 23867
rect 1728 23835 1768 23867
rect 1800 23835 1840 23867
rect 1872 23835 1912 23867
rect 1944 23835 1984 23867
rect 2016 23835 2056 23867
rect 2088 23835 2128 23867
rect 2160 23835 2200 23867
rect 2232 23835 2272 23867
rect 2304 23835 2344 23867
rect 2376 23835 2416 23867
rect 2448 23835 2488 23867
rect 2520 23835 2560 23867
rect 2592 23835 2632 23867
rect 2664 23835 2704 23867
rect 2736 23835 2776 23867
rect 2808 23835 2848 23867
rect 2880 23835 2920 23867
rect 2952 23835 2992 23867
rect 3024 23835 3064 23867
rect 3096 23835 3136 23867
rect 3168 23835 3208 23867
rect 3240 23835 3280 23867
rect 3312 23835 3352 23867
rect 3384 23835 3424 23867
rect 3456 23835 3496 23867
rect 3528 23835 3568 23867
rect 3600 23835 3640 23867
rect 3672 23835 3712 23867
rect 3744 23835 3784 23867
rect 3816 23835 3856 23867
rect 3888 23835 3950 23867
rect 50 23795 3950 23835
rect 50 23763 112 23795
rect 144 23763 184 23795
rect 216 23763 256 23795
rect 288 23763 328 23795
rect 360 23763 400 23795
rect 432 23763 472 23795
rect 504 23763 544 23795
rect 576 23763 616 23795
rect 648 23763 688 23795
rect 720 23763 760 23795
rect 792 23763 832 23795
rect 864 23763 904 23795
rect 936 23763 976 23795
rect 1008 23763 1048 23795
rect 1080 23763 1120 23795
rect 1152 23763 1192 23795
rect 1224 23763 1264 23795
rect 1296 23763 1336 23795
rect 1368 23763 1408 23795
rect 1440 23763 1480 23795
rect 1512 23763 1552 23795
rect 1584 23763 1624 23795
rect 1656 23763 1696 23795
rect 1728 23763 1768 23795
rect 1800 23763 1840 23795
rect 1872 23763 1912 23795
rect 1944 23763 1984 23795
rect 2016 23763 2056 23795
rect 2088 23763 2128 23795
rect 2160 23763 2200 23795
rect 2232 23763 2272 23795
rect 2304 23763 2344 23795
rect 2376 23763 2416 23795
rect 2448 23763 2488 23795
rect 2520 23763 2560 23795
rect 2592 23763 2632 23795
rect 2664 23763 2704 23795
rect 2736 23763 2776 23795
rect 2808 23763 2848 23795
rect 2880 23763 2920 23795
rect 2952 23763 2992 23795
rect 3024 23763 3064 23795
rect 3096 23763 3136 23795
rect 3168 23763 3208 23795
rect 3240 23763 3280 23795
rect 3312 23763 3352 23795
rect 3384 23763 3424 23795
rect 3456 23763 3496 23795
rect 3528 23763 3568 23795
rect 3600 23763 3640 23795
rect 3672 23763 3712 23795
rect 3744 23763 3784 23795
rect 3816 23763 3856 23795
rect 3888 23763 3950 23795
rect 50 23723 3950 23763
rect 50 23691 112 23723
rect 144 23691 184 23723
rect 216 23691 256 23723
rect 288 23691 328 23723
rect 360 23691 400 23723
rect 432 23691 472 23723
rect 504 23691 544 23723
rect 576 23691 616 23723
rect 648 23691 688 23723
rect 720 23691 760 23723
rect 792 23691 832 23723
rect 864 23691 904 23723
rect 936 23691 976 23723
rect 1008 23691 1048 23723
rect 1080 23691 1120 23723
rect 1152 23691 1192 23723
rect 1224 23691 1264 23723
rect 1296 23691 1336 23723
rect 1368 23691 1408 23723
rect 1440 23691 1480 23723
rect 1512 23691 1552 23723
rect 1584 23691 1624 23723
rect 1656 23691 1696 23723
rect 1728 23691 1768 23723
rect 1800 23691 1840 23723
rect 1872 23691 1912 23723
rect 1944 23691 1984 23723
rect 2016 23691 2056 23723
rect 2088 23691 2128 23723
rect 2160 23691 2200 23723
rect 2232 23691 2272 23723
rect 2304 23691 2344 23723
rect 2376 23691 2416 23723
rect 2448 23691 2488 23723
rect 2520 23691 2560 23723
rect 2592 23691 2632 23723
rect 2664 23691 2704 23723
rect 2736 23691 2776 23723
rect 2808 23691 2848 23723
rect 2880 23691 2920 23723
rect 2952 23691 2992 23723
rect 3024 23691 3064 23723
rect 3096 23691 3136 23723
rect 3168 23691 3208 23723
rect 3240 23691 3280 23723
rect 3312 23691 3352 23723
rect 3384 23691 3424 23723
rect 3456 23691 3496 23723
rect 3528 23691 3568 23723
rect 3600 23691 3640 23723
rect 3672 23691 3712 23723
rect 3744 23691 3784 23723
rect 3816 23691 3856 23723
rect 3888 23691 3950 23723
rect 50 23651 3950 23691
rect 50 23619 112 23651
rect 144 23619 184 23651
rect 216 23619 256 23651
rect 288 23619 328 23651
rect 360 23619 400 23651
rect 432 23619 472 23651
rect 504 23619 544 23651
rect 576 23619 616 23651
rect 648 23619 688 23651
rect 720 23619 760 23651
rect 792 23619 832 23651
rect 864 23619 904 23651
rect 936 23619 976 23651
rect 1008 23619 1048 23651
rect 1080 23619 1120 23651
rect 1152 23619 1192 23651
rect 1224 23619 1264 23651
rect 1296 23619 1336 23651
rect 1368 23619 1408 23651
rect 1440 23619 1480 23651
rect 1512 23619 1552 23651
rect 1584 23619 1624 23651
rect 1656 23619 1696 23651
rect 1728 23619 1768 23651
rect 1800 23619 1840 23651
rect 1872 23619 1912 23651
rect 1944 23619 1984 23651
rect 2016 23619 2056 23651
rect 2088 23619 2128 23651
rect 2160 23619 2200 23651
rect 2232 23619 2272 23651
rect 2304 23619 2344 23651
rect 2376 23619 2416 23651
rect 2448 23619 2488 23651
rect 2520 23619 2560 23651
rect 2592 23619 2632 23651
rect 2664 23619 2704 23651
rect 2736 23619 2776 23651
rect 2808 23619 2848 23651
rect 2880 23619 2920 23651
rect 2952 23619 2992 23651
rect 3024 23619 3064 23651
rect 3096 23619 3136 23651
rect 3168 23619 3208 23651
rect 3240 23619 3280 23651
rect 3312 23619 3352 23651
rect 3384 23619 3424 23651
rect 3456 23619 3496 23651
rect 3528 23619 3568 23651
rect 3600 23619 3640 23651
rect 3672 23619 3712 23651
rect 3744 23619 3784 23651
rect 3816 23619 3856 23651
rect 3888 23619 3950 23651
rect 50 23579 3950 23619
rect 50 23547 112 23579
rect 144 23547 184 23579
rect 216 23547 256 23579
rect 288 23547 328 23579
rect 360 23547 400 23579
rect 432 23547 472 23579
rect 504 23547 544 23579
rect 576 23547 616 23579
rect 648 23547 688 23579
rect 720 23547 760 23579
rect 792 23547 832 23579
rect 864 23547 904 23579
rect 936 23547 976 23579
rect 1008 23547 1048 23579
rect 1080 23547 1120 23579
rect 1152 23547 1192 23579
rect 1224 23547 1264 23579
rect 1296 23547 1336 23579
rect 1368 23547 1408 23579
rect 1440 23547 1480 23579
rect 1512 23547 1552 23579
rect 1584 23547 1624 23579
rect 1656 23547 1696 23579
rect 1728 23547 1768 23579
rect 1800 23547 1840 23579
rect 1872 23547 1912 23579
rect 1944 23547 1984 23579
rect 2016 23547 2056 23579
rect 2088 23547 2128 23579
rect 2160 23547 2200 23579
rect 2232 23547 2272 23579
rect 2304 23547 2344 23579
rect 2376 23547 2416 23579
rect 2448 23547 2488 23579
rect 2520 23547 2560 23579
rect 2592 23547 2632 23579
rect 2664 23547 2704 23579
rect 2736 23547 2776 23579
rect 2808 23547 2848 23579
rect 2880 23547 2920 23579
rect 2952 23547 2992 23579
rect 3024 23547 3064 23579
rect 3096 23547 3136 23579
rect 3168 23547 3208 23579
rect 3240 23547 3280 23579
rect 3312 23547 3352 23579
rect 3384 23547 3424 23579
rect 3456 23547 3496 23579
rect 3528 23547 3568 23579
rect 3600 23547 3640 23579
rect 3672 23547 3712 23579
rect 3744 23547 3784 23579
rect 3816 23547 3856 23579
rect 3888 23547 3950 23579
rect 50 23507 3950 23547
rect 50 23475 112 23507
rect 144 23475 184 23507
rect 216 23475 256 23507
rect 288 23475 328 23507
rect 360 23475 400 23507
rect 432 23475 472 23507
rect 504 23475 544 23507
rect 576 23475 616 23507
rect 648 23475 688 23507
rect 720 23475 760 23507
rect 792 23475 832 23507
rect 864 23475 904 23507
rect 936 23475 976 23507
rect 1008 23475 1048 23507
rect 1080 23475 1120 23507
rect 1152 23475 1192 23507
rect 1224 23475 1264 23507
rect 1296 23475 1336 23507
rect 1368 23475 1408 23507
rect 1440 23475 1480 23507
rect 1512 23475 1552 23507
rect 1584 23475 1624 23507
rect 1656 23475 1696 23507
rect 1728 23475 1768 23507
rect 1800 23475 1840 23507
rect 1872 23475 1912 23507
rect 1944 23475 1984 23507
rect 2016 23475 2056 23507
rect 2088 23475 2128 23507
rect 2160 23475 2200 23507
rect 2232 23475 2272 23507
rect 2304 23475 2344 23507
rect 2376 23475 2416 23507
rect 2448 23475 2488 23507
rect 2520 23475 2560 23507
rect 2592 23475 2632 23507
rect 2664 23475 2704 23507
rect 2736 23475 2776 23507
rect 2808 23475 2848 23507
rect 2880 23475 2920 23507
rect 2952 23475 2992 23507
rect 3024 23475 3064 23507
rect 3096 23475 3136 23507
rect 3168 23475 3208 23507
rect 3240 23475 3280 23507
rect 3312 23475 3352 23507
rect 3384 23475 3424 23507
rect 3456 23475 3496 23507
rect 3528 23475 3568 23507
rect 3600 23475 3640 23507
rect 3672 23475 3712 23507
rect 3744 23475 3784 23507
rect 3816 23475 3856 23507
rect 3888 23475 3950 23507
rect 50 23435 3950 23475
rect 50 23403 112 23435
rect 144 23403 184 23435
rect 216 23403 256 23435
rect 288 23403 328 23435
rect 360 23403 400 23435
rect 432 23403 472 23435
rect 504 23403 544 23435
rect 576 23403 616 23435
rect 648 23403 688 23435
rect 720 23403 760 23435
rect 792 23403 832 23435
rect 864 23403 904 23435
rect 936 23403 976 23435
rect 1008 23403 1048 23435
rect 1080 23403 1120 23435
rect 1152 23403 1192 23435
rect 1224 23403 1264 23435
rect 1296 23403 1336 23435
rect 1368 23403 1408 23435
rect 1440 23403 1480 23435
rect 1512 23403 1552 23435
rect 1584 23403 1624 23435
rect 1656 23403 1696 23435
rect 1728 23403 1768 23435
rect 1800 23403 1840 23435
rect 1872 23403 1912 23435
rect 1944 23403 1984 23435
rect 2016 23403 2056 23435
rect 2088 23403 2128 23435
rect 2160 23403 2200 23435
rect 2232 23403 2272 23435
rect 2304 23403 2344 23435
rect 2376 23403 2416 23435
rect 2448 23403 2488 23435
rect 2520 23403 2560 23435
rect 2592 23403 2632 23435
rect 2664 23403 2704 23435
rect 2736 23403 2776 23435
rect 2808 23403 2848 23435
rect 2880 23403 2920 23435
rect 2952 23403 2992 23435
rect 3024 23403 3064 23435
rect 3096 23403 3136 23435
rect 3168 23403 3208 23435
rect 3240 23403 3280 23435
rect 3312 23403 3352 23435
rect 3384 23403 3424 23435
rect 3456 23403 3496 23435
rect 3528 23403 3568 23435
rect 3600 23403 3640 23435
rect 3672 23403 3712 23435
rect 3744 23403 3784 23435
rect 3816 23403 3856 23435
rect 3888 23403 3950 23435
rect 50 23363 3950 23403
rect 50 23331 112 23363
rect 144 23331 184 23363
rect 216 23331 256 23363
rect 288 23331 328 23363
rect 360 23331 400 23363
rect 432 23331 472 23363
rect 504 23331 544 23363
rect 576 23331 616 23363
rect 648 23331 688 23363
rect 720 23331 760 23363
rect 792 23331 832 23363
rect 864 23331 904 23363
rect 936 23331 976 23363
rect 1008 23331 1048 23363
rect 1080 23331 1120 23363
rect 1152 23331 1192 23363
rect 1224 23331 1264 23363
rect 1296 23331 1336 23363
rect 1368 23331 1408 23363
rect 1440 23331 1480 23363
rect 1512 23331 1552 23363
rect 1584 23331 1624 23363
rect 1656 23331 1696 23363
rect 1728 23331 1768 23363
rect 1800 23331 1840 23363
rect 1872 23331 1912 23363
rect 1944 23331 1984 23363
rect 2016 23331 2056 23363
rect 2088 23331 2128 23363
rect 2160 23331 2200 23363
rect 2232 23331 2272 23363
rect 2304 23331 2344 23363
rect 2376 23331 2416 23363
rect 2448 23331 2488 23363
rect 2520 23331 2560 23363
rect 2592 23331 2632 23363
rect 2664 23331 2704 23363
rect 2736 23331 2776 23363
rect 2808 23331 2848 23363
rect 2880 23331 2920 23363
rect 2952 23331 2992 23363
rect 3024 23331 3064 23363
rect 3096 23331 3136 23363
rect 3168 23331 3208 23363
rect 3240 23331 3280 23363
rect 3312 23331 3352 23363
rect 3384 23331 3424 23363
rect 3456 23331 3496 23363
rect 3528 23331 3568 23363
rect 3600 23331 3640 23363
rect 3672 23331 3712 23363
rect 3744 23331 3784 23363
rect 3816 23331 3856 23363
rect 3888 23331 3950 23363
rect 50 23291 3950 23331
rect 50 23259 112 23291
rect 144 23259 184 23291
rect 216 23259 256 23291
rect 288 23259 328 23291
rect 360 23259 400 23291
rect 432 23259 472 23291
rect 504 23259 544 23291
rect 576 23259 616 23291
rect 648 23259 688 23291
rect 720 23259 760 23291
rect 792 23259 832 23291
rect 864 23259 904 23291
rect 936 23259 976 23291
rect 1008 23259 1048 23291
rect 1080 23259 1120 23291
rect 1152 23259 1192 23291
rect 1224 23259 1264 23291
rect 1296 23259 1336 23291
rect 1368 23259 1408 23291
rect 1440 23259 1480 23291
rect 1512 23259 1552 23291
rect 1584 23259 1624 23291
rect 1656 23259 1696 23291
rect 1728 23259 1768 23291
rect 1800 23259 1840 23291
rect 1872 23259 1912 23291
rect 1944 23259 1984 23291
rect 2016 23259 2056 23291
rect 2088 23259 2128 23291
rect 2160 23259 2200 23291
rect 2232 23259 2272 23291
rect 2304 23259 2344 23291
rect 2376 23259 2416 23291
rect 2448 23259 2488 23291
rect 2520 23259 2560 23291
rect 2592 23259 2632 23291
rect 2664 23259 2704 23291
rect 2736 23259 2776 23291
rect 2808 23259 2848 23291
rect 2880 23259 2920 23291
rect 2952 23259 2992 23291
rect 3024 23259 3064 23291
rect 3096 23259 3136 23291
rect 3168 23259 3208 23291
rect 3240 23259 3280 23291
rect 3312 23259 3352 23291
rect 3384 23259 3424 23291
rect 3456 23259 3496 23291
rect 3528 23259 3568 23291
rect 3600 23259 3640 23291
rect 3672 23259 3712 23291
rect 3744 23259 3784 23291
rect 3816 23259 3856 23291
rect 3888 23259 3950 23291
rect 50 23219 3950 23259
rect 50 23187 112 23219
rect 144 23187 184 23219
rect 216 23187 256 23219
rect 288 23187 328 23219
rect 360 23187 400 23219
rect 432 23187 472 23219
rect 504 23187 544 23219
rect 576 23187 616 23219
rect 648 23187 688 23219
rect 720 23187 760 23219
rect 792 23187 832 23219
rect 864 23187 904 23219
rect 936 23187 976 23219
rect 1008 23187 1048 23219
rect 1080 23187 1120 23219
rect 1152 23187 1192 23219
rect 1224 23187 1264 23219
rect 1296 23187 1336 23219
rect 1368 23187 1408 23219
rect 1440 23187 1480 23219
rect 1512 23187 1552 23219
rect 1584 23187 1624 23219
rect 1656 23187 1696 23219
rect 1728 23187 1768 23219
rect 1800 23187 1840 23219
rect 1872 23187 1912 23219
rect 1944 23187 1984 23219
rect 2016 23187 2056 23219
rect 2088 23187 2128 23219
rect 2160 23187 2200 23219
rect 2232 23187 2272 23219
rect 2304 23187 2344 23219
rect 2376 23187 2416 23219
rect 2448 23187 2488 23219
rect 2520 23187 2560 23219
rect 2592 23187 2632 23219
rect 2664 23187 2704 23219
rect 2736 23187 2776 23219
rect 2808 23187 2848 23219
rect 2880 23187 2920 23219
rect 2952 23187 2992 23219
rect 3024 23187 3064 23219
rect 3096 23187 3136 23219
rect 3168 23187 3208 23219
rect 3240 23187 3280 23219
rect 3312 23187 3352 23219
rect 3384 23187 3424 23219
rect 3456 23187 3496 23219
rect 3528 23187 3568 23219
rect 3600 23187 3640 23219
rect 3672 23187 3712 23219
rect 3744 23187 3784 23219
rect 3816 23187 3856 23219
rect 3888 23187 3950 23219
rect 50 23124 3950 23187
rect 50 22874 3950 22924
rect 50 22842 112 22874
rect 144 22842 184 22874
rect 216 22842 256 22874
rect 288 22842 328 22874
rect 360 22842 400 22874
rect 432 22842 472 22874
rect 504 22842 544 22874
rect 576 22842 616 22874
rect 648 22842 688 22874
rect 720 22842 760 22874
rect 792 22842 832 22874
rect 864 22842 904 22874
rect 936 22842 976 22874
rect 1008 22842 1048 22874
rect 1080 22842 1120 22874
rect 1152 22842 1192 22874
rect 1224 22842 1264 22874
rect 1296 22842 1336 22874
rect 1368 22842 1408 22874
rect 1440 22842 1480 22874
rect 1512 22842 1552 22874
rect 1584 22842 1624 22874
rect 1656 22842 1696 22874
rect 1728 22842 1768 22874
rect 1800 22842 1840 22874
rect 1872 22842 1912 22874
rect 1944 22842 1984 22874
rect 2016 22842 2056 22874
rect 2088 22842 2128 22874
rect 2160 22842 2200 22874
rect 2232 22842 2272 22874
rect 2304 22842 2344 22874
rect 2376 22842 2416 22874
rect 2448 22842 2488 22874
rect 2520 22842 2560 22874
rect 2592 22842 2632 22874
rect 2664 22842 2704 22874
rect 2736 22842 2776 22874
rect 2808 22842 2848 22874
rect 2880 22842 2920 22874
rect 2952 22842 2992 22874
rect 3024 22842 3064 22874
rect 3096 22842 3136 22874
rect 3168 22842 3208 22874
rect 3240 22842 3280 22874
rect 3312 22842 3352 22874
rect 3384 22842 3424 22874
rect 3456 22842 3496 22874
rect 3528 22842 3568 22874
rect 3600 22842 3640 22874
rect 3672 22842 3712 22874
rect 3744 22842 3784 22874
rect 3816 22842 3856 22874
rect 3888 22842 3950 22874
rect 50 22802 3950 22842
rect 50 22770 112 22802
rect 144 22770 184 22802
rect 216 22770 256 22802
rect 288 22770 328 22802
rect 360 22770 400 22802
rect 432 22770 472 22802
rect 504 22770 544 22802
rect 576 22770 616 22802
rect 648 22770 688 22802
rect 720 22770 760 22802
rect 792 22770 832 22802
rect 864 22770 904 22802
rect 936 22770 976 22802
rect 1008 22770 1048 22802
rect 1080 22770 1120 22802
rect 1152 22770 1192 22802
rect 1224 22770 1264 22802
rect 1296 22770 1336 22802
rect 1368 22770 1408 22802
rect 1440 22770 1480 22802
rect 1512 22770 1552 22802
rect 1584 22770 1624 22802
rect 1656 22770 1696 22802
rect 1728 22770 1768 22802
rect 1800 22770 1840 22802
rect 1872 22770 1912 22802
rect 1944 22770 1984 22802
rect 2016 22770 2056 22802
rect 2088 22770 2128 22802
rect 2160 22770 2200 22802
rect 2232 22770 2272 22802
rect 2304 22770 2344 22802
rect 2376 22770 2416 22802
rect 2448 22770 2488 22802
rect 2520 22770 2560 22802
rect 2592 22770 2632 22802
rect 2664 22770 2704 22802
rect 2736 22770 2776 22802
rect 2808 22770 2848 22802
rect 2880 22770 2920 22802
rect 2952 22770 2992 22802
rect 3024 22770 3064 22802
rect 3096 22770 3136 22802
rect 3168 22770 3208 22802
rect 3240 22770 3280 22802
rect 3312 22770 3352 22802
rect 3384 22770 3424 22802
rect 3456 22770 3496 22802
rect 3528 22770 3568 22802
rect 3600 22770 3640 22802
rect 3672 22770 3712 22802
rect 3744 22770 3784 22802
rect 3816 22770 3856 22802
rect 3888 22770 3950 22802
rect 50 22730 3950 22770
rect 50 22698 112 22730
rect 144 22698 184 22730
rect 216 22698 256 22730
rect 288 22698 328 22730
rect 360 22698 400 22730
rect 432 22698 472 22730
rect 504 22698 544 22730
rect 576 22698 616 22730
rect 648 22698 688 22730
rect 720 22698 760 22730
rect 792 22698 832 22730
rect 864 22698 904 22730
rect 936 22698 976 22730
rect 1008 22698 1048 22730
rect 1080 22698 1120 22730
rect 1152 22698 1192 22730
rect 1224 22698 1264 22730
rect 1296 22698 1336 22730
rect 1368 22698 1408 22730
rect 1440 22698 1480 22730
rect 1512 22698 1552 22730
rect 1584 22698 1624 22730
rect 1656 22698 1696 22730
rect 1728 22698 1768 22730
rect 1800 22698 1840 22730
rect 1872 22698 1912 22730
rect 1944 22698 1984 22730
rect 2016 22698 2056 22730
rect 2088 22698 2128 22730
rect 2160 22698 2200 22730
rect 2232 22698 2272 22730
rect 2304 22698 2344 22730
rect 2376 22698 2416 22730
rect 2448 22698 2488 22730
rect 2520 22698 2560 22730
rect 2592 22698 2632 22730
rect 2664 22698 2704 22730
rect 2736 22698 2776 22730
rect 2808 22698 2848 22730
rect 2880 22698 2920 22730
rect 2952 22698 2992 22730
rect 3024 22698 3064 22730
rect 3096 22698 3136 22730
rect 3168 22698 3208 22730
rect 3240 22698 3280 22730
rect 3312 22698 3352 22730
rect 3384 22698 3424 22730
rect 3456 22698 3496 22730
rect 3528 22698 3568 22730
rect 3600 22698 3640 22730
rect 3672 22698 3712 22730
rect 3744 22698 3784 22730
rect 3816 22698 3856 22730
rect 3888 22698 3950 22730
rect 50 22658 3950 22698
rect 50 22626 112 22658
rect 144 22626 184 22658
rect 216 22626 256 22658
rect 288 22626 328 22658
rect 360 22626 400 22658
rect 432 22626 472 22658
rect 504 22626 544 22658
rect 576 22626 616 22658
rect 648 22626 688 22658
rect 720 22626 760 22658
rect 792 22626 832 22658
rect 864 22626 904 22658
rect 936 22626 976 22658
rect 1008 22626 1048 22658
rect 1080 22626 1120 22658
rect 1152 22626 1192 22658
rect 1224 22626 1264 22658
rect 1296 22626 1336 22658
rect 1368 22626 1408 22658
rect 1440 22626 1480 22658
rect 1512 22626 1552 22658
rect 1584 22626 1624 22658
rect 1656 22626 1696 22658
rect 1728 22626 1768 22658
rect 1800 22626 1840 22658
rect 1872 22626 1912 22658
rect 1944 22626 1984 22658
rect 2016 22626 2056 22658
rect 2088 22626 2128 22658
rect 2160 22626 2200 22658
rect 2232 22626 2272 22658
rect 2304 22626 2344 22658
rect 2376 22626 2416 22658
rect 2448 22626 2488 22658
rect 2520 22626 2560 22658
rect 2592 22626 2632 22658
rect 2664 22626 2704 22658
rect 2736 22626 2776 22658
rect 2808 22626 2848 22658
rect 2880 22626 2920 22658
rect 2952 22626 2992 22658
rect 3024 22626 3064 22658
rect 3096 22626 3136 22658
rect 3168 22626 3208 22658
rect 3240 22626 3280 22658
rect 3312 22626 3352 22658
rect 3384 22626 3424 22658
rect 3456 22626 3496 22658
rect 3528 22626 3568 22658
rect 3600 22626 3640 22658
rect 3672 22626 3712 22658
rect 3744 22626 3784 22658
rect 3816 22626 3856 22658
rect 3888 22626 3950 22658
rect 50 22586 3950 22626
rect 50 22554 112 22586
rect 144 22554 184 22586
rect 216 22554 256 22586
rect 288 22554 328 22586
rect 360 22554 400 22586
rect 432 22554 472 22586
rect 504 22554 544 22586
rect 576 22554 616 22586
rect 648 22554 688 22586
rect 720 22554 760 22586
rect 792 22554 832 22586
rect 864 22554 904 22586
rect 936 22554 976 22586
rect 1008 22554 1048 22586
rect 1080 22554 1120 22586
rect 1152 22554 1192 22586
rect 1224 22554 1264 22586
rect 1296 22554 1336 22586
rect 1368 22554 1408 22586
rect 1440 22554 1480 22586
rect 1512 22554 1552 22586
rect 1584 22554 1624 22586
rect 1656 22554 1696 22586
rect 1728 22554 1768 22586
rect 1800 22554 1840 22586
rect 1872 22554 1912 22586
rect 1944 22554 1984 22586
rect 2016 22554 2056 22586
rect 2088 22554 2128 22586
rect 2160 22554 2200 22586
rect 2232 22554 2272 22586
rect 2304 22554 2344 22586
rect 2376 22554 2416 22586
rect 2448 22554 2488 22586
rect 2520 22554 2560 22586
rect 2592 22554 2632 22586
rect 2664 22554 2704 22586
rect 2736 22554 2776 22586
rect 2808 22554 2848 22586
rect 2880 22554 2920 22586
rect 2952 22554 2992 22586
rect 3024 22554 3064 22586
rect 3096 22554 3136 22586
rect 3168 22554 3208 22586
rect 3240 22554 3280 22586
rect 3312 22554 3352 22586
rect 3384 22554 3424 22586
rect 3456 22554 3496 22586
rect 3528 22554 3568 22586
rect 3600 22554 3640 22586
rect 3672 22554 3712 22586
rect 3744 22554 3784 22586
rect 3816 22554 3856 22586
rect 3888 22554 3950 22586
rect 50 22514 3950 22554
rect 50 22482 112 22514
rect 144 22482 184 22514
rect 216 22482 256 22514
rect 288 22482 328 22514
rect 360 22482 400 22514
rect 432 22482 472 22514
rect 504 22482 544 22514
rect 576 22482 616 22514
rect 648 22482 688 22514
rect 720 22482 760 22514
rect 792 22482 832 22514
rect 864 22482 904 22514
rect 936 22482 976 22514
rect 1008 22482 1048 22514
rect 1080 22482 1120 22514
rect 1152 22482 1192 22514
rect 1224 22482 1264 22514
rect 1296 22482 1336 22514
rect 1368 22482 1408 22514
rect 1440 22482 1480 22514
rect 1512 22482 1552 22514
rect 1584 22482 1624 22514
rect 1656 22482 1696 22514
rect 1728 22482 1768 22514
rect 1800 22482 1840 22514
rect 1872 22482 1912 22514
rect 1944 22482 1984 22514
rect 2016 22482 2056 22514
rect 2088 22482 2128 22514
rect 2160 22482 2200 22514
rect 2232 22482 2272 22514
rect 2304 22482 2344 22514
rect 2376 22482 2416 22514
rect 2448 22482 2488 22514
rect 2520 22482 2560 22514
rect 2592 22482 2632 22514
rect 2664 22482 2704 22514
rect 2736 22482 2776 22514
rect 2808 22482 2848 22514
rect 2880 22482 2920 22514
rect 2952 22482 2992 22514
rect 3024 22482 3064 22514
rect 3096 22482 3136 22514
rect 3168 22482 3208 22514
rect 3240 22482 3280 22514
rect 3312 22482 3352 22514
rect 3384 22482 3424 22514
rect 3456 22482 3496 22514
rect 3528 22482 3568 22514
rect 3600 22482 3640 22514
rect 3672 22482 3712 22514
rect 3744 22482 3784 22514
rect 3816 22482 3856 22514
rect 3888 22482 3950 22514
rect 50 22442 3950 22482
rect 50 22410 112 22442
rect 144 22410 184 22442
rect 216 22410 256 22442
rect 288 22410 328 22442
rect 360 22410 400 22442
rect 432 22410 472 22442
rect 504 22410 544 22442
rect 576 22410 616 22442
rect 648 22410 688 22442
rect 720 22410 760 22442
rect 792 22410 832 22442
rect 864 22410 904 22442
rect 936 22410 976 22442
rect 1008 22410 1048 22442
rect 1080 22410 1120 22442
rect 1152 22410 1192 22442
rect 1224 22410 1264 22442
rect 1296 22410 1336 22442
rect 1368 22410 1408 22442
rect 1440 22410 1480 22442
rect 1512 22410 1552 22442
rect 1584 22410 1624 22442
rect 1656 22410 1696 22442
rect 1728 22410 1768 22442
rect 1800 22410 1840 22442
rect 1872 22410 1912 22442
rect 1944 22410 1984 22442
rect 2016 22410 2056 22442
rect 2088 22410 2128 22442
rect 2160 22410 2200 22442
rect 2232 22410 2272 22442
rect 2304 22410 2344 22442
rect 2376 22410 2416 22442
rect 2448 22410 2488 22442
rect 2520 22410 2560 22442
rect 2592 22410 2632 22442
rect 2664 22410 2704 22442
rect 2736 22410 2776 22442
rect 2808 22410 2848 22442
rect 2880 22410 2920 22442
rect 2952 22410 2992 22442
rect 3024 22410 3064 22442
rect 3096 22410 3136 22442
rect 3168 22410 3208 22442
rect 3240 22410 3280 22442
rect 3312 22410 3352 22442
rect 3384 22410 3424 22442
rect 3456 22410 3496 22442
rect 3528 22410 3568 22442
rect 3600 22410 3640 22442
rect 3672 22410 3712 22442
rect 3744 22410 3784 22442
rect 3816 22410 3856 22442
rect 3888 22410 3950 22442
rect 50 22370 3950 22410
rect 50 22338 112 22370
rect 144 22338 184 22370
rect 216 22338 256 22370
rect 288 22338 328 22370
rect 360 22338 400 22370
rect 432 22338 472 22370
rect 504 22338 544 22370
rect 576 22338 616 22370
rect 648 22338 688 22370
rect 720 22338 760 22370
rect 792 22338 832 22370
rect 864 22338 904 22370
rect 936 22338 976 22370
rect 1008 22338 1048 22370
rect 1080 22338 1120 22370
rect 1152 22338 1192 22370
rect 1224 22338 1264 22370
rect 1296 22338 1336 22370
rect 1368 22338 1408 22370
rect 1440 22338 1480 22370
rect 1512 22338 1552 22370
rect 1584 22338 1624 22370
rect 1656 22338 1696 22370
rect 1728 22338 1768 22370
rect 1800 22338 1840 22370
rect 1872 22338 1912 22370
rect 1944 22338 1984 22370
rect 2016 22338 2056 22370
rect 2088 22338 2128 22370
rect 2160 22338 2200 22370
rect 2232 22338 2272 22370
rect 2304 22338 2344 22370
rect 2376 22338 2416 22370
rect 2448 22338 2488 22370
rect 2520 22338 2560 22370
rect 2592 22338 2632 22370
rect 2664 22338 2704 22370
rect 2736 22338 2776 22370
rect 2808 22338 2848 22370
rect 2880 22338 2920 22370
rect 2952 22338 2992 22370
rect 3024 22338 3064 22370
rect 3096 22338 3136 22370
rect 3168 22338 3208 22370
rect 3240 22338 3280 22370
rect 3312 22338 3352 22370
rect 3384 22338 3424 22370
rect 3456 22338 3496 22370
rect 3528 22338 3568 22370
rect 3600 22338 3640 22370
rect 3672 22338 3712 22370
rect 3744 22338 3784 22370
rect 3816 22338 3856 22370
rect 3888 22338 3950 22370
rect 50 22298 3950 22338
rect 50 22266 112 22298
rect 144 22266 184 22298
rect 216 22266 256 22298
rect 288 22266 328 22298
rect 360 22266 400 22298
rect 432 22266 472 22298
rect 504 22266 544 22298
rect 576 22266 616 22298
rect 648 22266 688 22298
rect 720 22266 760 22298
rect 792 22266 832 22298
rect 864 22266 904 22298
rect 936 22266 976 22298
rect 1008 22266 1048 22298
rect 1080 22266 1120 22298
rect 1152 22266 1192 22298
rect 1224 22266 1264 22298
rect 1296 22266 1336 22298
rect 1368 22266 1408 22298
rect 1440 22266 1480 22298
rect 1512 22266 1552 22298
rect 1584 22266 1624 22298
rect 1656 22266 1696 22298
rect 1728 22266 1768 22298
rect 1800 22266 1840 22298
rect 1872 22266 1912 22298
rect 1944 22266 1984 22298
rect 2016 22266 2056 22298
rect 2088 22266 2128 22298
rect 2160 22266 2200 22298
rect 2232 22266 2272 22298
rect 2304 22266 2344 22298
rect 2376 22266 2416 22298
rect 2448 22266 2488 22298
rect 2520 22266 2560 22298
rect 2592 22266 2632 22298
rect 2664 22266 2704 22298
rect 2736 22266 2776 22298
rect 2808 22266 2848 22298
rect 2880 22266 2920 22298
rect 2952 22266 2992 22298
rect 3024 22266 3064 22298
rect 3096 22266 3136 22298
rect 3168 22266 3208 22298
rect 3240 22266 3280 22298
rect 3312 22266 3352 22298
rect 3384 22266 3424 22298
rect 3456 22266 3496 22298
rect 3528 22266 3568 22298
rect 3600 22266 3640 22298
rect 3672 22266 3712 22298
rect 3744 22266 3784 22298
rect 3816 22266 3856 22298
rect 3888 22266 3950 22298
rect 50 22226 3950 22266
rect 50 22194 112 22226
rect 144 22194 184 22226
rect 216 22194 256 22226
rect 288 22194 328 22226
rect 360 22194 400 22226
rect 432 22194 472 22226
rect 504 22194 544 22226
rect 576 22194 616 22226
rect 648 22194 688 22226
rect 720 22194 760 22226
rect 792 22194 832 22226
rect 864 22194 904 22226
rect 936 22194 976 22226
rect 1008 22194 1048 22226
rect 1080 22194 1120 22226
rect 1152 22194 1192 22226
rect 1224 22194 1264 22226
rect 1296 22194 1336 22226
rect 1368 22194 1408 22226
rect 1440 22194 1480 22226
rect 1512 22194 1552 22226
rect 1584 22194 1624 22226
rect 1656 22194 1696 22226
rect 1728 22194 1768 22226
rect 1800 22194 1840 22226
rect 1872 22194 1912 22226
rect 1944 22194 1984 22226
rect 2016 22194 2056 22226
rect 2088 22194 2128 22226
rect 2160 22194 2200 22226
rect 2232 22194 2272 22226
rect 2304 22194 2344 22226
rect 2376 22194 2416 22226
rect 2448 22194 2488 22226
rect 2520 22194 2560 22226
rect 2592 22194 2632 22226
rect 2664 22194 2704 22226
rect 2736 22194 2776 22226
rect 2808 22194 2848 22226
rect 2880 22194 2920 22226
rect 2952 22194 2992 22226
rect 3024 22194 3064 22226
rect 3096 22194 3136 22226
rect 3168 22194 3208 22226
rect 3240 22194 3280 22226
rect 3312 22194 3352 22226
rect 3384 22194 3424 22226
rect 3456 22194 3496 22226
rect 3528 22194 3568 22226
rect 3600 22194 3640 22226
rect 3672 22194 3712 22226
rect 3744 22194 3784 22226
rect 3816 22194 3856 22226
rect 3888 22194 3950 22226
rect 50 22154 3950 22194
rect 50 22122 112 22154
rect 144 22122 184 22154
rect 216 22122 256 22154
rect 288 22122 328 22154
rect 360 22122 400 22154
rect 432 22122 472 22154
rect 504 22122 544 22154
rect 576 22122 616 22154
rect 648 22122 688 22154
rect 720 22122 760 22154
rect 792 22122 832 22154
rect 864 22122 904 22154
rect 936 22122 976 22154
rect 1008 22122 1048 22154
rect 1080 22122 1120 22154
rect 1152 22122 1192 22154
rect 1224 22122 1264 22154
rect 1296 22122 1336 22154
rect 1368 22122 1408 22154
rect 1440 22122 1480 22154
rect 1512 22122 1552 22154
rect 1584 22122 1624 22154
rect 1656 22122 1696 22154
rect 1728 22122 1768 22154
rect 1800 22122 1840 22154
rect 1872 22122 1912 22154
rect 1944 22122 1984 22154
rect 2016 22122 2056 22154
rect 2088 22122 2128 22154
rect 2160 22122 2200 22154
rect 2232 22122 2272 22154
rect 2304 22122 2344 22154
rect 2376 22122 2416 22154
rect 2448 22122 2488 22154
rect 2520 22122 2560 22154
rect 2592 22122 2632 22154
rect 2664 22122 2704 22154
rect 2736 22122 2776 22154
rect 2808 22122 2848 22154
rect 2880 22122 2920 22154
rect 2952 22122 2992 22154
rect 3024 22122 3064 22154
rect 3096 22122 3136 22154
rect 3168 22122 3208 22154
rect 3240 22122 3280 22154
rect 3312 22122 3352 22154
rect 3384 22122 3424 22154
rect 3456 22122 3496 22154
rect 3528 22122 3568 22154
rect 3600 22122 3640 22154
rect 3672 22122 3712 22154
rect 3744 22122 3784 22154
rect 3816 22122 3856 22154
rect 3888 22122 3950 22154
rect 50 22082 3950 22122
rect 50 22050 112 22082
rect 144 22050 184 22082
rect 216 22050 256 22082
rect 288 22050 328 22082
rect 360 22050 400 22082
rect 432 22050 472 22082
rect 504 22050 544 22082
rect 576 22050 616 22082
rect 648 22050 688 22082
rect 720 22050 760 22082
rect 792 22050 832 22082
rect 864 22050 904 22082
rect 936 22050 976 22082
rect 1008 22050 1048 22082
rect 1080 22050 1120 22082
rect 1152 22050 1192 22082
rect 1224 22050 1264 22082
rect 1296 22050 1336 22082
rect 1368 22050 1408 22082
rect 1440 22050 1480 22082
rect 1512 22050 1552 22082
rect 1584 22050 1624 22082
rect 1656 22050 1696 22082
rect 1728 22050 1768 22082
rect 1800 22050 1840 22082
rect 1872 22050 1912 22082
rect 1944 22050 1984 22082
rect 2016 22050 2056 22082
rect 2088 22050 2128 22082
rect 2160 22050 2200 22082
rect 2232 22050 2272 22082
rect 2304 22050 2344 22082
rect 2376 22050 2416 22082
rect 2448 22050 2488 22082
rect 2520 22050 2560 22082
rect 2592 22050 2632 22082
rect 2664 22050 2704 22082
rect 2736 22050 2776 22082
rect 2808 22050 2848 22082
rect 2880 22050 2920 22082
rect 2952 22050 2992 22082
rect 3024 22050 3064 22082
rect 3096 22050 3136 22082
rect 3168 22050 3208 22082
rect 3240 22050 3280 22082
rect 3312 22050 3352 22082
rect 3384 22050 3424 22082
rect 3456 22050 3496 22082
rect 3528 22050 3568 22082
rect 3600 22050 3640 22082
rect 3672 22050 3712 22082
rect 3744 22050 3784 22082
rect 3816 22050 3856 22082
rect 3888 22050 3950 22082
rect 50 22010 3950 22050
rect 50 21978 112 22010
rect 144 21978 184 22010
rect 216 21978 256 22010
rect 288 21978 328 22010
rect 360 21978 400 22010
rect 432 21978 472 22010
rect 504 21978 544 22010
rect 576 21978 616 22010
rect 648 21978 688 22010
rect 720 21978 760 22010
rect 792 21978 832 22010
rect 864 21978 904 22010
rect 936 21978 976 22010
rect 1008 21978 1048 22010
rect 1080 21978 1120 22010
rect 1152 21978 1192 22010
rect 1224 21978 1264 22010
rect 1296 21978 1336 22010
rect 1368 21978 1408 22010
rect 1440 21978 1480 22010
rect 1512 21978 1552 22010
rect 1584 21978 1624 22010
rect 1656 21978 1696 22010
rect 1728 21978 1768 22010
rect 1800 21978 1840 22010
rect 1872 21978 1912 22010
rect 1944 21978 1984 22010
rect 2016 21978 2056 22010
rect 2088 21978 2128 22010
rect 2160 21978 2200 22010
rect 2232 21978 2272 22010
rect 2304 21978 2344 22010
rect 2376 21978 2416 22010
rect 2448 21978 2488 22010
rect 2520 21978 2560 22010
rect 2592 21978 2632 22010
rect 2664 21978 2704 22010
rect 2736 21978 2776 22010
rect 2808 21978 2848 22010
rect 2880 21978 2920 22010
rect 2952 21978 2992 22010
rect 3024 21978 3064 22010
rect 3096 21978 3136 22010
rect 3168 21978 3208 22010
rect 3240 21978 3280 22010
rect 3312 21978 3352 22010
rect 3384 21978 3424 22010
rect 3456 21978 3496 22010
rect 3528 21978 3568 22010
rect 3600 21978 3640 22010
rect 3672 21978 3712 22010
rect 3744 21978 3784 22010
rect 3816 21978 3856 22010
rect 3888 21978 3950 22010
rect 50 21938 3950 21978
rect 50 21906 112 21938
rect 144 21906 184 21938
rect 216 21906 256 21938
rect 288 21906 328 21938
rect 360 21906 400 21938
rect 432 21906 472 21938
rect 504 21906 544 21938
rect 576 21906 616 21938
rect 648 21906 688 21938
rect 720 21906 760 21938
rect 792 21906 832 21938
rect 864 21906 904 21938
rect 936 21906 976 21938
rect 1008 21906 1048 21938
rect 1080 21906 1120 21938
rect 1152 21906 1192 21938
rect 1224 21906 1264 21938
rect 1296 21906 1336 21938
rect 1368 21906 1408 21938
rect 1440 21906 1480 21938
rect 1512 21906 1552 21938
rect 1584 21906 1624 21938
rect 1656 21906 1696 21938
rect 1728 21906 1768 21938
rect 1800 21906 1840 21938
rect 1872 21906 1912 21938
rect 1944 21906 1984 21938
rect 2016 21906 2056 21938
rect 2088 21906 2128 21938
rect 2160 21906 2200 21938
rect 2232 21906 2272 21938
rect 2304 21906 2344 21938
rect 2376 21906 2416 21938
rect 2448 21906 2488 21938
rect 2520 21906 2560 21938
rect 2592 21906 2632 21938
rect 2664 21906 2704 21938
rect 2736 21906 2776 21938
rect 2808 21906 2848 21938
rect 2880 21906 2920 21938
rect 2952 21906 2992 21938
rect 3024 21906 3064 21938
rect 3096 21906 3136 21938
rect 3168 21906 3208 21938
rect 3240 21906 3280 21938
rect 3312 21906 3352 21938
rect 3384 21906 3424 21938
rect 3456 21906 3496 21938
rect 3528 21906 3568 21938
rect 3600 21906 3640 21938
rect 3672 21906 3712 21938
rect 3744 21906 3784 21938
rect 3816 21906 3856 21938
rect 3888 21906 3950 21938
rect 50 21866 3950 21906
rect 50 21834 112 21866
rect 144 21834 184 21866
rect 216 21834 256 21866
rect 288 21834 328 21866
rect 360 21834 400 21866
rect 432 21834 472 21866
rect 504 21834 544 21866
rect 576 21834 616 21866
rect 648 21834 688 21866
rect 720 21834 760 21866
rect 792 21834 832 21866
rect 864 21834 904 21866
rect 936 21834 976 21866
rect 1008 21834 1048 21866
rect 1080 21834 1120 21866
rect 1152 21834 1192 21866
rect 1224 21834 1264 21866
rect 1296 21834 1336 21866
rect 1368 21834 1408 21866
rect 1440 21834 1480 21866
rect 1512 21834 1552 21866
rect 1584 21834 1624 21866
rect 1656 21834 1696 21866
rect 1728 21834 1768 21866
rect 1800 21834 1840 21866
rect 1872 21834 1912 21866
rect 1944 21834 1984 21866
rect 2016 21834 2056 21866
rect 2088 21834 2128 21866
rect 2160 21834 2200 21866
rect 2232 21834 2272 21866
rect 2304 21834 2344 21866
rect 2376 21834 2416 21866
rect 2448 21834 2488 21866
rect 2520 21834 2560 21866
rect 2592 21834 2632 21866
rect 2664 21834 2704 21866
rect 2736 21834 2776 21866
rect 2808 21834 2848 21866
rect 2880 21834 2920 21866
rect 2952 21834 2992 21866
rect 3024 21834 3064 21866
rect 3096 21834 3136 21866
rect 3168 21834 3208 21866
rect 3240 21834 3280 21866
rect 3312 21834 3352 21866
rect 3384 21834 3424 21866
rect 3456 21834 3496 21866
rect 3528 21834 3568 21866
rect 3600 21834 3640 21866
rect 3672 21834 3712 21866
rect 3744 21834 3784 21866
rect 3816 21834 3856 21866
rect 3888 21834 3950 21866
rect 50 21794 3950 21834
rect 50 21762 112 21794
rect 144 21762 184 21794
rect 216 21762 256 21794
rect 288 21762 328 21794
rect 360 21762 400 21794
rect 432 21762 472 21794
rect 504 21762 544 21794
rect 576 21762 616 21794
rect 648 21762 688 21794
rect 720 21762 760 21794
rect 792 21762 832 21794
rect 864 21762 904 21794
rect 936 21762 976 21794
rect 1008 21762 1048 21794
rect 1080 21762 1120 21794
rect 1152 21762 1192 21794
rect 1224 21762 1264 21794
rect 1296 21762 1336 21794
rect 1368 21762 1408 21794
rect 1440 21762 1480 21794
rect 1512 21762 1552 21794
rect 1584 21762 1624 21794
rect 1656 21762 1696 21794
rect 1728 21762 1768 21794
rect 1800 21762 1840 21794
rect 1872 21762 1912 21794
rect 1944 21762 1984 21794
rect 2016 21762 2056 21794
rect 2088 21762 2128 21794
rect 2160 21762 2200 21794
rect 2232 21762 2272 21794
rect 2304 21762 2344 21794
rect 2376 21762 2416 21794
rect 2448 21762 2488 21794
rect 2520 21762 2560 21794
rect 2592 21762 2632 21794
rect 2664 21762 2704 21794
rect 2736 21762 2776 21794
rect 2808 21762 2848 21794
rect 2880 21762 2920 21794
rect 2952 21762 2992 21794
rect 3024 21762 3064 21794
rect 3096 21762 3136 21794
rect 3168 21762 3208 21794
rect 3240 21762 3280 21794
rect 3312 21762 3352 21794
rect 3384 21762 3424 21794
rect 3456 21762 3496 21794
rect 3528 21762 3568 21794
rect 3600 21762 3640 21794
rect 3672 21762 3712 21794
rect 3744 21762 3784 21794
rect 3816 21762 3856 21794
rect 3888 21762 3950 21794
rect 50 21722 3950 21762
rect 50 21690 112 21722
rect 144 21690 184 21722
rect 216 21690 256 21722
rect 288 21690 328 21722
rect 360 21690 400 21722
rect 432 21690 472 21722
rect 504 21690 544 21722
rect 576 21690 616 21722
rect 648 21690 688 21722
rect 720 21690 760 21722
rect 792 21690 832 21722
rect 864 21690 904 21722
rect 936 21690 976 21722
rect 1008 21690 1048 21722
rect 1080 21690 1120 21722
rect 1152 21690 1192 21722
rect 1224 21690 1264 21722
rect 1296 21690 1336 21722
rect 1368 21690 1408 21722
rect 1440 21690 1480 21722
rect 1512 21690 1552 21722
rect 1584 21690 1624 21722
rect 1656 21690 1696 21722
rect 1728 21690 1768 21722
rect 1800 21690 1840 21722
rect 1872 21690 1912 21722
rect 1944 21690 1984 21722
rect 2016 21690 2056 21722
rect 2088 21690 2128 21722
rect 2160 21690 2200 21722
rect 2232 21690 2272 21722
rect 2304 21690 2344 21722
rect 2376 21690 2416 21722
rect 2448 21690 2488 21722
rect 2520 21690 2560 21722
rect 2592 21690 2632 21722
rect 2664 21690 2704 21722
rect 2736 21690 2776 21722
rect 2808 21690 2848 21722
rect 2880 21690 2920 21722
rect 2952 21690 2992 21722
rect 3024 21690 3064 21722
rect 3096 21690 3136 21722
rect 3168 21690 3208 21722
rect 3240 21690 3280 21722
rect 3312 21690 3352 21722
rect 3384 21690 3424 21722
rect 3456 21690 3496 21722
rect 3528 21690 3568 21722
rect 3600 21690 3640 21722
rect 3672 21690 3712 21722
rect 3744 21690 3784 21722
rect 3816 21690 3856 21722
rect 3888 21690 3950 21722
rect 50 21650 3950 21690
rect 50 21618 112 21650
rect 144 21618 184 21650
rect 216 21618 256 21650
rect 288 21618 328 21650
rect 360 21618 400 21650
rect 432 21618 472 21650
rect 504 21618 544 21650
rect 576 21618 616 21650
rect 648 21618 688 21650
rect 720 21618 760 21650
rect 792 21618 832 21650
rect 864 21618 904 21650
rect 936 21618 976 21650
rect 1008 21618 1048 21650
rect 1080 21618 1120 21650
rect 1152 21618 1192 21650
rect 1224 21618 1264 21650
rect 1296 21618 1336 21650
rect 1368 21618 1408 21650
rect 1440 21618 1480 21650
rect 1512 21618 1552 21650
rect 1584 21618 1624 21650
rect 1656 21618 1696 21650
rect 1728 21618 1768 21650
rect 1800 21618 1840 21650
rect 1872 21618 1912 21650
rect 1944 21618 1984 21650
rect 2016 21618 2056 21650
rect 2088 21618 2128 21650
rect 2160 21618 2200 21650
rect 2232 21618 2272 21650
rect 2304 21618 2344 21650
rect 2376 21618 2416 21650
rect 2448 21618 2488 21650
rect 2520 21618 2560 21650
rect 2592 21618 2632 21650
rect 2664 21618 2704 21650
rect 2736 21618 2776 21650
rect 2808 21618 2848 21650
rect 2880 21618 2920 21650
rect 2952 21618 2992 21650
rect 3024 21618 3064 21650
rect 3096 21618 3136 21650
rect 3168 21618 3208 21650
rect 3240 21618 3280 21650
rect 3312 21618 3352 21650
rect 3384 21618 3424 21650
rect 3456 21618 3496 21650
rect 3528 21618 3568 21650
rect 3600 21618 3640 21650
rect 3672 21618 3712 21650
rect 3744 21618 3784 21650
rect 3816 21618 3856 21650
rect 3888 21618 3950 21650
rect 50 21578 3950 21618
rect 50 21546 112 21578
rect 144 21546 184 21578
rect 216 21546 256 21578
rect 288 21546 328 21578
rect 360 21546 400 21578
rect 432 21546 472 21578
rect 504 21546 544 21578
rect 576 21546 616 21578
rect 648 21546 688 21578
rect 720 21546 760 21578
rect 792 21546 832 21578
rect 864 21546 904 21578
rect 936 21546 976 21578
rect 1008 21546 1048 21578
rect 1080 21546 1120 21578
rect 1152 21546 1192 21578
rect 1224 21546 1264 21578
rect 1296 21546 1336 21578
rect 1368 21546 1408 21578
rect 1440 21546 1480 21578
rect 1512 21546 1552 21578
rect 1584 21546 1624 21578
rect 1656 21546 1696 21578
rect 1728 21546 1768 21578
rect 1800 21546 1840 21578
rect 1872 21546 1912 21578
rect 1944 21546 1984 21578
rect 2016 21546 2056 21578
rect 2088 21546 2128 21578
rect 2160 21546 2200 21578
rect 2232 21546 2272 21578
rect 2304 21546 2344 21578
rect 2376 21546 2416 21578
rect 2448 21546 2488 21578
rect 2520 21546 2560 21578
rect 2592 21546 2632 21578
rect 2664 21546 2704 21578
rect 2736 21546 2776 21578
rect 2808 21546 2848 21578
rect 2880 21546 2920 21578
rect 2952 21546 2992 21578
rect 3024 21546 3064 21578
rect 3096 21546 3136 21578
rect 3168 21546 3208 21578
rect 3240 21546 3280 21578
rect 3312 21546 3352 21578
rect 3384 21546 3424 21578
rect 3456 21546 3496 21578
rect 3528 21546 3568 21578
rect 3600 21546 3640 21578
rect 3672 21546 3712 21578
rect 3744 21546 3784 21578
rect 3816 21546 3856 21578
rect 3888 21546 3950 21578
rect 50 21506 3950 21546
rect 50 21474 112 21506
rect 144 21474 184 21506
rect 216 21474 256 21506
rect 288 21474 328 21506
rect 360 21474 400 21506
rect 432 21474 472 21506
rect 504 21474 544 21506
rect 576 21474 616 21506
rect 648 21474 688 21506
rect 720 21474 760 21506
rect 792 21474 832 21506
rect 864 21474 904 21506
rect 936 21474 976 21506
rect 1008 21474 1048 21506
rect 1080 21474 1120 21506
rect 1152 21474 1192 21506
rect 1224 21474 1264 21506
rect 1296 21474 1336 21506
rect 1368 21474 1408 21506
rect 1440 21474 1480 21506
rect 1512 21474 1552 21506
rect 1584 21474 1624 21506
rect 1656 21474 1696 21506
rect 1728 21474 1768 21506
rect 1800 21474 1840 21506
rect 1872 21474 1912 21506
rect 1944 21474 1984 21506
rect 2016 21474 2056 21506
rect 2088 21474 2128 21506
rect 2160 21474 2200 21506
rect 2232 21474 2272 21506
rect 2304 21474 2344 21506
rect 2376 21474 2416 21506
rect 2448 21474 2488 21506
rect 2520 21474 2560 21506
rect 2592 21474 2632 21506
rect 2664 21474 2704 21506
rect 2736 21474 2776 21506
rect 2808 21474 2848 21506
rect 2880 21474 2920 21506
rect 2952 21474 2992 21506
rect 3024 21474 3064 21506
rect 3096 21474 3136 21506
rect 3168 21474 3208 21506
rect 3240 21474 3280 21506
rect 3312 21474 3352 21506
rect 3384 21474 3424 21506
rect 3456 21474 3496 21506
rect 3528 21474 3568 21506
rect 3600 21474 3640 21506
rect 3672 21474 3712 21506
rect 3744 21474 3784 21506
rect 3816 21474 3856 21506
rect 3888 21474 3950 21506
rect 50 21434 3950 21474
rect 50 21402 112 21434
rect 144 21402 184 21434
rect 216 21402 256 21434
rect 288 21402 328 21434
rect 360 21402 400 21434
rect 432 21402 472 21434
rect 504 21402 544 21434
rect 576 21402 616 21434
rect 648 21402 688 21434
rect 720 21402 760 21434
rect 792 21402 832 21434
rect 864 21402 904 21434
rect 936 21402 976 21434
rect 1008 21402 1048 21434
rect 1080 21402 1120 21434
rect 1152 21402 1192 21434
rect 1224 21402 1264 21434
rect 1296 21402 1336 21434
rect 1368 21402 1408 21434
rect 1440 21402 1480 21434
rect 1512 21402 1552 21434
rect 1584 21402 1624 21434
rect 1656 21402 1696 21434
rect 1728 21402 1768 21434
rect 1800 21402 1840 21434
rect 1872 21402 1912 21434
rect 1944 21402 1984 21434
rect 2016 21402 2056 21434
rect 2088 21402 2128 21434
rect 2160 21402 2200 21434
rect 2232 21402 2272 21434
rect 2304 21402 2344 21434
rect 2376 21402 2416 21434
rect 2448 21402 2488 21434
rect 2520 21402 2560 21434
rect 2592 21402 2632 21434
rect 2664 21402 2704 21434
rect 2736 21402 2776 21434
rect 2808 21402 2848 21434
rect 2880 21402 2920 21434
rect 2952 21402 2992 21434
rect 3024 21402 3064 21434
rect 3096 21402 3136 21434
rect 3168 21402 3208 21434
rect 3240 21402 3280 21434
rect 3312 21402 3352 21434
rect 3384 21402 3424 21434
rect 3456 21402 3496 21434
rect 3528 21402 3568 21434
rect 3600 21402 3640 21434
rect 3672 21402 3712 21434
rect 3744 21402 3784 21434
rect 3816 21402 3856 21434
rect 3888 21402 3950 21434
rect 50 21362 3950 21402
rect 50 21330 112 21362
rect 144 21330 184 21362
rect 216 21330 256 21362
rect 288 21330 328 21362
rect 360 21330 400 21362
rect 432 21330 472 21362
rect 504 21330 544 21362
rect 576 21330 616 21362
rect 648 21330 688 21362
rect 720 21330 760 21362
rect 792 21330 832 21362
rect 864 21330 904 21362
rect 936 21330 976 21362
rect 1008 21330 1048 21362
rect 1080 21330 1120 21362
rect 1152 21330 1192 21362
rect 1224 21330 1264 21362
rect 1296 21330 1336 21362
rect 1368 21330 1408 21362
rect 1440 21330 1480 21362
rect 1512 21330 1552 21362
rect 1584 21330 1624 21362
rect 1656 21330 1696 21362
rect 1728 21330 1768 21362
rect 1800 21330 1840 21362
rect 1872 21330 1912 21362
rect 1944 21330 1984 21362
rect 2016 21330 2056 21362
rect 2088 21330 2128 21362
rect 2160 21330 2200 21362
rect 2232 21330 2272 21362
rect 2304 21330 2344 21362
rect 2376 21330 2416 21362
rect 2448 21330 2488 21362
rect 2520 21330 2560 21362
rect 2592 21330 2632 21362
rect 2664 21330 2704 21362
rect 2736 21330 2776 21362
rect 2808 21330 2848 21362
rect 2880 21330 2920 21362
rect 2952 21330 2992 21362
rect 3024 21330 3064 21362
rect 3096 21330 3136 21362
rect 3168 21330 3208 21362
rect 3240 21330 3280 21362
rect 3312 21330 3352 21362
rect 3384 21330 3424 21362
rect 3456 21330 3496 21362
rect 3528 21330 3568 21362
rect 3600 21330 3640 21362
rect 3672 21330 3712 21362
rect 3744 21330 3784 21362
rect 3816 21330 3856 21362
rect 3888 21330 3950 21362
rect 50 21290 3950 21330
rect 50 21258 112 21290
rect 144 21258 184 21290
rect 216 21258 256 21290
rect 288 21258 328 21290
rect 360 21258 400 21290
rect 432 21258 472 21290
rect 504 21258 544 21290
rect 576 21258 616 21290
rect 648 21258 688 21290
rect 720 21258 760 21290
rect 792 21258 832 21290
rect 864 21258 904 21290
rect 936 21258 976 21290
rect 1008 21258 1048 21290
rect 1080 21258 1120 21290
rect 1152 21258 1192 21290
rect 1224 21258 1264 21290
rect 1296 21258 1336 21290
rect 1368 21258 1408 21290
rect 1440 21258 1480 21290
rect 1512 21258 1552 21290
rect 1584 21258 1624 21290
rect 1656 21258 1696 21290
rect 1728 21258 1768 21290
rect 1800 21258 1840 21290
rect 1872 21258 1912 21290
rect 1944 21258 1984 21290
rect 2016 21258 2056 21290
rect 2088 21258 2128 21290
rect 2160 21258 2200 21290
rect 2232 21258 2272 21290
rect 2304 21258 2344 21290
rect 2376 21258 2416 21290
rect 2448 21258 2488 21290
rect 2520 21258 2560 21290
rect 2592 21258 2632 21290
rect 2664 21258 2704 21290
rect 2736 21258 2776 21290
rect 2808 21258 2848 21290
rect 2880 21258 2920 21290
rect 2952 21258 2992 21290
rect 3024 21258 3064 21290
rect 3096 21258 3136 21290
rect 3168 21258 3208 21290
rect 3240 21258 3280 21290
rect 3312 21258 3352 21290
rect 3384 21258 3424 21290
rect 3456 21258 3496 21290
rect 3528 21258 3568 21290
rect 3600 21258 3640 21290
rect 3672 21258 3712 21290
rect 3744 21258 3784 21290
rect 3816 21258 3856 21290
rect 3888 21258 3950 21290
rect 50 21218 3950 21258
rect 50 21186 112 21218
rect 144 21186 184 21218
rect 216 21186 256 21218
rect 288 21186 328 21218
rect 360 21186 400 21218
rect 432 21186 472 21218
rect 504 21186 544 21218
rect 576 21186 616 21218
rect 648 21186 688 21218
rect 720 21186 760 21218
rect 792 21186 832 21218
rect 864 21186 904 21218
rect 936 21186 976 21218
rect 1008 21186 1048 21218
rect 1080 21186 1120 21218
rect 1152 21186 1192 21218
rect 1224 21186 1264 21218
rect 1296 21186 1336 21218
rect 1368 21186 1408 21218
rect 1440 21186 1480 21218
rect 1512 21186 1552 21218
rect 1584 21186 1624 21218
rect 1656 21186 1696 21218
rect 1728 21186 1768 21218
rect 1800 21186 1840 21218
rect 1872 21186 1912 21218
rect 1944 21186 1984 21218
rect 2016 21186 2056 21218
rect 2088 21186 2128 21218
rect 2160 21186 2200 21218
rect 2232 21186 2272 21218
rect 2304 21186 2344 21218
rect 2376 21186 2416 21218
rect 2448 21186 2488 21218
rect 2520 21186 2560 21218
rect 2592 21186 2632 21218
rect 2664 21186 2704 21218
rect 2736 21186 2776 21218
rect 2808 21186 2848 21218
rect 2880 21186 2920 21218
rect 2952 21186 2992 21218
rect 3024 21186 3064 21218
rect 3096 21186 3136 21218
rect 3168 21186 3208 21218
rect 3240 21186 3280 21218
rect 3312 21186 3352 21218
rect 3384 21186 3424 21218
rect 3456 21186 3496 21218
rect 3528 21186 3568 21218
rect 3600 21186 3640 21218
rect 3672 21186 3712 21218
rect 3744 21186 3784 21218
rect 3816 21186 3856 21218
rect 3888 21186 3950 21218
rect 50 21146 3950 21186
rect 50 21114 112 21146
rect 144 21114 184 21146
rect 216 21114 256 21146
rect 288 21114 328 21146
rect 360 21114 400 21146
rect 432 21114 472 21146
rect 504 21114 544 21146
rect 576 21114 616 21146
rect 648 21114 688 21146
rect 720 21114 760 21146
rect 792 21114 832 21146
rect 864 21114 904 21146
rect 936 21114 976 21146
rect 1008 21114 1048 21146
rect 1080 21114 1120 21146
rect 1152 21114 1192 21146
rect 1224 21114 1264 21146
rect 1296 21114 1336 21146
rect 1368 21114 1408 21146
rect 1440 21114 1480 21146
rect 1512 21114 1552 21146
rect 1584 21114 1624 21146
rect 1656 21114 1696 21146
rect 1728 21114 1768 21146
rect 1800 21114 1840 21146
rect 1872 21114 1912 21146
rect 1944 21114 1984 21146
rect 2016 21114 2056 21146
rect 2088 21114 2128 21146
rect 2160 21114 2200 21146
rect 2232 21114 2272 21146
rect 2304 21114 2344 21146
rect 2376 21114 2416 21146
rect 2448 21114 2488 21146
rect 2520 21114 2560 21146
rect 2592 21114 2632 21146
rect 2664 21114 2704 21146
rect 2736 21114 2776 21146
rect 2808 21114 2848 21146
rect 2880 21114 2920 21146
rect 2952 21114 2992 21146
rect 3024 21114 3064 21146
rect 3096 21114 3136 21146
rect 3168 21114 3208 21146
rect 3240 21114 3280 21146
rect 3312 21114 3352 21146
rect 3384 21114 3424 21146
rect 3456 21114 3496 21146
rect 3528 21114 3568 21146
rect 3600 21114 3640 21146
rect 3672 21114 3712 21146
rect 3744 21114 3784 21146
rect 3816 21114 3856 21146
rect 3888 21114 3950 21146
rect 50 21074 3950 21114
rect 50 21042 112 21074
rect 144 21042 184 21074
rect 216 21042 256 21074
rect 288 21042 328 21074
rect 360 21042 400 21074
rect 432 21042 472 21074
rect 504 21042 544 21074
rect 576 21042 616 21074
rect 648 21042 688 21074
rect 720 21042 760 21074
rect 792 21042 832 21074
rect 864 21042 904 21074
rect 936 21042 976 21074
rect 1008 21042 1048 21074
rect 1080 21042 1120 21074
rect 1152 21042 1192 21074
rect 1224 21042 1264 21074
rect 1296 21042 1336 21074
rect 1368 21042 1408 21074
rect 1440 21042 1480 21074
rect 1512 21042 1552 21074
rect 1584 21042 1624 21074
rect 1656 21042 1696 21074
rect 1728 21042 1768 21074
rect 1800 21042 1840 21074
rect 1872 21042 1912 21074
rect 1944 21042 1984 21074
rect 2016 21042 2056 21074
rect 2088 21042 2128 21074
rect 2160 21042 2200 21074
rect 2232 21042 2272 21074
rect 2304 21042 2344 21074
rect 2376 21042 2416 21074
rect 2448 21042 2488 21074
rect 2520 21042 2560 21074
rect 2592 21042 2632 21074
rect 2664 21042 2704 21074
rect 2736 21042 2776 21074
rect 2808 21042 2848 21074
rect 2880 21042 2920 21074
rect 2952 21042 2992 21074
rect 3024 21042 3064 21074
rect 3096 21042 3136 21074
rect 3168 21042 3208 21074
rect 3240 21042 3280 21074
rect 3312 21042 3352 21074
rect 3384 21042 3424 21074
rect 3456 21042 3496 21074
rect 3528 21042 3568 21074
rect 3600 21042 3640 21074
rect 3672 21042 3712 21074
rect 3744 21042 3784 21074
rect 3816 21042 3856 21074
rect 3888 21042 3950 21074
rect 50 21002 3950 21042
rect 50 20970 112 21002
rect 144 20970 184 21002
rect 216 20970 256 21002
rect 288 20970 328 21002
rect 360 20970 400 21002
rect 432 20970 472 21002
rect 504 20970 544 21002
rect 576 20970 616 21002
rect 648 20970 688 21002
rect 720 20970 760 21002
rect 792 20970 832 21002
rect 864 20970 904 21002
rect 936 20970 976 21002
rect 1008 20970 1048 21002
rect 1080 20970 1120 21002
rect 1152 20970 1192 21002
rect 1224 20970 1264 21002
rect 1296 20970 1336 21002
rect 1368 20970 1408 21002
rect 1440 20970 1480 21002
rect 1512 20970 1552 21002
rect 1584 20970 1624 21002
rect 1656 20970 1696 21002
rect 1728 20970 1768 21002
rect 1800 20970 1840 21002
rect 1872 20970 1912 21002
rect 1944 20970 1984 21002
rect 2016 20970 2056 21002
rect 2088 20970 2128 21002
rect 2160 20970 2200 21002
rect 2232 20970 2272 21002
rect 2304 20970 2344 21002
rect 2376 20970 2416 21002
rect 2448 20970 2488 21002
rect 2520 20970 2560 21002
rect 2592 20970 2632 21002
rect 2664 20970 2704 21002
rect 2736 20970 2776 21002
rect 2808 20970 2848 21002
rect 2880 20970 2920 21002
rect 2952 20970 2992 21002
rect 3024 20970 3064 21002
rect 3096 20970 3136 21002
rect 3168 20970 3208 21002
rect 3240 20970 3280 21002
rect 3312 20970 3352 21002
rect 3384 20970 3424 21002
rect 3456 20970 3496 21002
rect 3528 20970 3568 21002
rect 3600 20970 3640 21002
rect 3672 20970 3712 21002
rect 3744 20970 3784 21002
rect 3816 20970 3856 21002
rect 3888 20970 3950 21002
rect 50 20930 3950 20970
rect 50 20898 112 20930
rect 144 20898 184 20930
rect 216 20898 256 20930
rect 288 20898 328 20930
rect 360 20898 400 20930
rect 432 20898 472 20930
rect 504 20898 544 20930
rect 576 20898 616 20930
rect 648 20898 688 20930
rect 720 20898 760 20930
rect 792 20898 832 20930
rect 864 20898 904 20930
rect 936 20898 976 20930
rect 1008 20898 1048 20930
rect 1080 20898 1120 20930
rect 1152 20898 1192 20930
rect 1224 20898 1264 20930
rect 1296 20898 1336 20930
rect 1368 20898 1408 20930
rect 1440 20898 1480 20930
rect 1512 20898 1552 20930
rect 1584 20898 1624 20930
rect 1656 20898 1696 20930
rect 1728 20898 1768 20930
rect 1800 20898 1840 20930
rect 1872 20898 1912 20930
rect 1944 20898 1984 20930
rect 2016 20898 2056 20930
rect 2088 20898 2128 20930
rect 2160 20898 2200 20930
rect 2232 20898 2272 20930
rect 2304 20898 2344 20930
rect 2376 20898 2416 20930
rect 2448 20898 2488 20930
rect 2520 20898 2560 20930
rect 2592 20898 2632 20930
rect 2664 20898 2704 20930
rect 2736 20898 2776 20930
rect 2808 20898 2848 20930
rect 2880 20898 2920 20930
rect 2952 20898 2992 20930
rect 3024 20898 3064 20930
rect 3096 20898 3136 20930
rect 3168 20898 3208 20930
rect 3240 20898 3280 20930
rect 3312 20898 3352 20930
rect 3384 20898 3424 20930
rect 3456 20898 3496 20930
rect 3528 20898 3568 20930
rect 3600 20898 3640 20930
rect 3672 20898 3712 20930
rect 3744 20898 3784 20930
rect 3816 20898 3856 20930
rect 3888 20898 3950 20930
rect 50 20858 3950 20898
rect 50 20826 112 20858
rect 144 20826 184 20858
rect 216 20826 256 20858
rect 288 20826 328 20858
rect 360 20826 400 20858
rect 432 20826 472 20858
rect 504 20826 544 20858
rect 576 20826 616 20858
rect 648 20826 688 20858
rect 720 20826 760 20858
rect 792 20826 832 20858
rect 864 20826 904 20858
rect 936 20826 976 20858
rect 1008 20826 1048 20858
rect 1080 20826 1120 20858
rect 1152 20826 1192 20858
rect 1224 20826 1264 20858
rect 1296 20826 1336 20858
rect 1368 20826 1408 20858
rect 1440 20826 1480 20858
rect 1512 20826 1552 20858
rect 1584 20826 1624 20858
rect 1656 20826 1696 20858
rect 1728 20826 1768 20858
rect 1800 20826 1840 20858
rect 1872 20826 1912 20858
rect 1944 20826 1984 20858
rect 2016 20826 2056 20858
rect 2088 20826 2128 20858
rect 2160 20826 2200 20858
rect 2232 20826 2272 20858
rect 2304 20826 2344 20858
rect 2376 20826 2416 20858
rect 2448 20826 2488 20858
rect 2520 20826 2560 20858
rect 2592 20826 2632 20858
rect 2664 20826 2704 20858
rect 2736 20826 2776 20858
rect 2808 20826 2848 20858
rect 2880 20826 2920 20858
rect 2952 20826 2992 20858
rect 3024 20826 3064 20858
rect 3096 20826 3136 20858
rect 3168 20826 3208 20858
rect 3240 20826 3280 20858
rect 3312 20826 3352 20858
rect 3384 20826 3424 20858
rect 3456 20826 3496 20858
rect 3528 20826 3568 20858
rect 3600 20826 3640 20858
rect 3672 20826 3712 20858
rect 3744 20826 3784 20858
rect 3816 20826 3856 20858
rect 3888 20826 3950 20858
rect 50 20786 3950 20826
rect 50 20754 112 20786
rect 144 20754 184 20786
rect 216 20754 256 20786
rect 288 20754 328 20786
rect 360 20754 400 20786
rect 432 20754 472 20786
rect 504 20754 544 20786
rect 576 20754 616 20786
rect 648 20754 688 20786
rect 720 20754 760 20786
rect 792 20754 832 20786
rect 864 20754 904 20786
rect 936 20754 976 20786
rect 1008 20754 1048 20786
rect 1080 20754 1120 20786
rect 1152 20754 1192 20786
rect 1224 20754 1264 20786
rect 1296 20754 1336 20786
rect 1368 20754 1408 20786
rect 1440 20754 1480 20786
rect 1512 20754 1552 20786
rect 1584 20754 1624 20786
rect 1656 20754 1696 20786
rect 1728 20754 1768 20786
rect 1800 20754 1840 20786
rect 1872 20754 1912 20786
rect 1944 20754 1984 20786
rect 2016 20754 2056 20786
rect 2088 20754 2128 20786
rect 2160 20754 2200 20786
rect 2232 20754 2272 20786
rect 2304 20754 2344 20786
rect 2376 20754 2416 20786
rect 2448 20754 2488 20786
rect 2520 20754 2560 20786
rect 2592 20754 2632 20786
rect 2664 20754 2704 20786
rect 2736 20754 2776 20786
rect 2808 20754 2848 20786
rect 2880 20754 2920 20786
rect 2952 20754 2992 20786
rect 3024 20754 3064 20786
rect 3096 20754 3136 20786
rect 3168 20754 3208 20786
rect 3240 20754 3280 20786
rect 3312 20754 3352 20786
rect 3384 20754 3424 20786
rect 3456 20754 3496 20786
rect 3528 20754 3568 20786
rect 3600 20754 3640 20786
rect 3672 20754 3712 20786
rect 3744 20754 3784 20786
rect 3816 20754 3856 20786
rect 3888 20754 3950 20786
rect 50 20714 3950 20754
rect 50 20682 112 20714
rect 144 20682 184 20714
rect 216 20682 256 20714
rect 288 20682 328 20714
rect 360 20682 400 20714
rect 432 20682 472 20714
rect 504 20682 544 20714
rect 576 20682 616 20714
rect 648 20682 688 20714
rect 720 20682 760 20714
rect 792 20682 832 20714
rect 864 20682 904 20714
rect 936 20682 976 20714
rect 1008 20682 1048 20714
rect 1080 20682 1120 20714
rect 1152 20682 1192 20714
rect 1224 20682 1264 20714
rect 1296 20682 1336 20714
rect 1368 20682 1408 20714
rect 1440 20682 1480 20714
rect 1512 20682 1552 20714
rect 1584 20682 1624 20714
rect 1656 20682 1696 20714
rect 1728 20682 1768 20714
rect 1800 20682 1840 20714
rect 1872 20682 1912 20714
rect 1944 20682 1984 20714
rect 2016 20682 2056 20714
rect 2088 20682 2128 20714
rect 2160 20682 2200 20714
rect 2232 20682 2272 20714
rect 2304 20682 2344 20714
rect 2376 20682 2416 20714
rect 2448 20682 2488 20714
rect 2520 20682 2560 20714
rect 2592 20682 2632 20714
rect 2664 20682 2704 20714
rect 2736 20682 2776 20714
rect 2808 20682 2848 20714
rect 2880 20682 2920 20714
rect 2952 20682 2992 20714
rect 3024 20682 3064 20714
rect 3096 20682 3136 20714
rect 3168 20682 3208 20714
rect 3240 20682 3280 20714
rect 3312 20682 3352 20714
rect 3384 20682 3424 20714
rect 3456 20682 3496 20714
rect 3528 20682 3568 20714
rect 3600 20682 3640 20714
rect 3672 20682 3712 20714
rect 3744 20682 3784 20714
rect 3816 20682 3856 20714
rect 3888 20682 3950 20714
rect 50 20642 3950 20682
rect 50 20610 112 20642
rect 144 20610 184 20642
rect 216 20610 256 20642
rect 288 20610 328 20642
rect 360 20610 400 20642
rect 432 20610 472 20642
rect 504 20610 544 20642
rect 576 20610 616 20642
rect 648 20610 688 20642
rect 720 20610 760 20642
rect 792 20610 832 20642
rect 864 20610 904 20642
rect 936 20610 976 20642
rect 1008 20610 1048 20642
rect 1080 20610 1120 20642
rect 1152 20610 1192 20642
rect 1224 20610 1264 20642
rect 1296 20610 1336 20642
rect 1368 20610 1408 20642
rect 1440 20610 1480 20642
rect 1512 20610 1552 20642
rect 1584 20610 1624 20642
rect 1656 20610 1696 20642
rect 1728 20610 1768 20642
rect 1800 20610 1840 20642
rect 1872 20610 1912 20642
rect 1944 20610 1984 20642
rect 2016 20610 2056 20642
rect 2088 20610 2128 20642
rect 2160 20610 2200 20642
rect 2232 20610 2272 20642
rect 2304 20610 2344 20642
rect 2376 20610 2416 20642
rect 2448 20610 2488 20642
rect 2520 20610 2560 20642
rect 2592 20610 2632 20642
rect 2664 20610 2704 20642
rect 2736 20610 2776 20642
rect 2808 20610 2848 20642
rect 2880 20610 2920 20642
rect 2952 20610 2992 20642
rect 3024 20610 3064 20642
rect 3096 20610 3136 20642
rect 3168 20610 3208 20642
rect 3240 20610 3280 20642
rect 3312 20610 3352 20642
rect 3384 20610 3424 20642
rect 3456 20610 3496 20642
rect 3528 20610 3568 20642
rect 3600 20610 3640 20642
rect 3672 20610 3712 20642
rect 3744 20610 3784 20642
rect 3816 20610 3856 20642
rect 3888 20610 3950 20642
rect 50 20570 3950 20610
rect 50 20538 112 20570
rect 144 20538 184 20570
rect 216 20538 256 20570
rect 288 20538 328 20570
rect 360 20538 400 20570
rect 432 20538 472 20570
rect 504 20538 544 20570
rect 576 20538 616 20570
rect 648 20538 688 20570
rect 720 20538 760 20570
rect 792 20538 832 20570
rect 864 20538 904 20570
rect 936 20538 976 20570
rect 1008 20538 1048 20570
rect 1080 20538 1120 20570
rect 1152 20538 1192 20570
rect 1224 20538 1264 20570
rect 1296 20538 1336 20570
rect 1368 20538 1408 20570
rect 1440 20538 1480 20570
rect 1512 20538 1552 20570
rect 1584 20538 1624 20570
rect 1656 20538 1696 20570
rect 1728 20538 1768 20570
rect 1800 20538 1840 20570
rect 1872 20538 1912 20570
rect 1944 20538 1984 20570
rect 2016 20538 2056 20570
rect 2088 20538 2128 20570
rect 2160 20538 2200 20570
rect 2232 20538 2272 20570
rect 2304 20538 2344 20570
rect 2376 20538 2416 20570
rect 2448 20538 2488 20570
rect 2520 20538 2560 20570
rect 2592 20538 2632 20570
rect 2664 20538 2704 20570
rect 2736 20538 2776 20570
rect 2808 20538 2848 20570
rect 2880 20538 2920 20570
rect 2952 20538 2992 20570
rect 3024 20538 3064 20570
rect 3096 20538 3136 20570
rect 3168 20538 3208 20570
rect 3240 20538 3280 20570
rect 3312 20538 3352 20570
rect 3384 20538 3424 20570
rect 3456 20538 3496 20570
rect 3528 20538 3568 20570
rect 3600 20538 3640 20570
rect 3672 20538 3712 20570
rect 3744 20538 3784 20570
rect 3816 20538 3856 20570
rect 3888 20538 3950 20570
rect 50 20498 3950 20538
rect 50 20466 112 20498
rect 144 20466 184 20498
rect 216 20466 256 20498
rect 288 20466 328 20498
rect 360 20466 400 20498
rect 432 20466 472 20498
rect 504 20466 544 20498
rect 576 20466 616 20498
rect 648 20466 688 20498
rect 720 20466 760 20498
rect 792 20466 832 20498
rect 864 20466 904 20498
rect 936 20466 976 20498
rect 1008 20466 1048 20498
rect 1080 20466 1120 20498
rect 1152 20466 1192 20498
rect 1224 20466 1264 20498
rect 1296 20466 1336 20498
rect 1368 20466 1408 20498
rect 1440 20466 1480 20498
rect 1512 20466 1552 20498
rect 1584 20466 1624 20498
rect 1656 20466 1696 20498
rect 1728 20466 1768 20498
rect 1800 20466 1840 20498
rect 1872 20466 1912 20498
rect 1944 20466 1984 20498
rect 2016 20466 2056 20498
rect 2088 20466 2128 20498
rect 2160 20466 2200 20498
rect 2232 20466 2272 20498
rect 2304 20466 2344 20498
rect 2376 20466 2416 20498
rect 2448 20466 2488 20498
rect 2520 20466 2560 20498
rect 2592 20466 2632 20498
rect 2664 20466 2704 20498
rect 2736 20466 2776 20498
rect 2808 20466 2848 20498
rect 2880 20466 2920 20498
rect 2952 20466 2992 20498
rect 3024 20466 3064 20498
rect 3096 20466 3136 20498
rect 3168 20466 3208 20498
rect 3240 20466 3280 20498
rect 3312 20466 3352 20498
rect 3384 20466 3424 20498
rect 3456 20466 3496 20498
rect 3528 20466 3568 20498
rect 3600 20466 3640 20498
rect 3672 20466 3712 20498
rect 3744 20466 3784 20498
rect 3816 20466 3856 20498
rect 3888 20466 3950 20498
rect 50 20426 3950 20466
rect 50 20394 112 20426
rect 144 20394 184 20426
rect 216 20394 256 20426
rect 288 20394 328 20426
rect 360 20394 400 20426
rect 432 20394 472 20426
rect 504 20394 544 20426
rect 576 20394 616 20426
rect 648 20394 688 20426
rect 720 20394 760 20426
rect 792 20394 832 20426
rect 864 20394 904 20426
rect 936 20394 976 20426
rect 1008 20394 1048 20426
rect 1080 20394 1120 20426
rect 1152 20394 1192 20426
rect 1224 20394 1264 20426
rect 1296 20394 1336 20426
rect 1368 20394 1408 20426
rect 1440 20394 1480 20426
rect 1512 20394 1552 20426
rect 1584 20394 1624 20426
rect 1656 20394 1696 20426
rect 1728 20394 1768 20426
rect 1800 20394 1840 20426
rect 1872 20394 1912 20426
rect 1944 20394 1984 20426
rect 2016 20394 2056 20426
rect 2088 20394 2128 20426
rect 2160 20394 2200 20426
rect 2232 20394 2272 20426
rect 2304 20394 2344 20426
rect 2376 20394 2416 20426
rect 2448 20394 2488 20426
rect 2520 20394 2560 20426
rect 2592 20394 2632 20426
rect 2664 20394 2704 20426
rect 2736 20394 2776 20426
rect 2808 20394 2848 20426
rect 2880 20394 2920 20426
rect 2952 20394 2992 20426
rect 3024 20394 3064 20426
rect 3096 20394 3136 20426
rect 3168 20394 3208 20426
rect 3240 20394 3280 20426
rect 3312 20394 3352 20426
rect 3384 20394 3424 20426
rect 3456 20394 3496 20426
rect 3528 20394 3568 20426
rect 3600 20394 3640 20426
rect 3672 20394 3712 20426
rect 3744 20394 3784 20426
rect 3816 20394 3856 20426
rect 3888 20394 3950 20426
rect 50 20354 3950 20394
rect 50 20322 112 20354
rect 144 20322 184 20354
rect 216 20322 256 20354
rect 288 20322 328 20354
rect 360 20322 400 20354
rect 432 20322 472 20354
rect 504 20322 544 20354
rect 576 20322 616 20354
rect 648 20322 688 20354
rect 720 20322 760 20354
rect 792 20322 832 20354
rect 864 20322 904 20354
rect 936 20322 976 20354
rect 1008 20322 1048 20354
rect 1080 20322 1120 20354
rect 1152 20322 1192 20354
rect 1224 20322 1264 20354
rect 1296 20322 1336 20354
rect 1368 20322 1408 20354
rect 1440 20322 1480 20354
rect 1512 20322 1552 20354
rect 1584 20322 1624 20354
rect 1656 20322 1696 20354
rect 1728 20322 1768 20354
rect 1800 20322 1840 20354
rect 1872 20322 1912 20354
rect 1944 20322 1984 20354
rect 2016 20322 2056 20354
rect 2088 20322 2128 20354
rect 2160 20322 2200 20354
rect 2232 20322 2272 20354
rect 2304 20322 2344 20354
rect 2376 20322 2416 20354
rect 2448 20322 2488 20354
rect 2520 20322 2560 20354
rect 2592 20322 2632 20354
rect 2664 20322 2704 20354
rect 2736 20322 2776 20354
rect 2808 20322 2848 20354
rect 2880 20322 2920 20354
rect 2952 20322 2992 20354
rect 3024 20322 3064 20354
rect 3096 20322 3136 20354
rect 3168 20322 3208 20354
rect 3240 20322 3280 20354
rect 3312 20322 3352 20354
rect 3384 20322 3424 20354
rect 3456 20322 3496 20354
rect 3528 20322 3568 20354
rect 3600 20322 3640 20354
rect 3672 20322 3712 20354
rect 3744 20322 3784 20354
rect 3816 20322 3856 20354
rect 3888 20322 3950 20354
rect 50 20282 3950 20322
rect 50 20250 112 20282
rect 144 20250 184 20282
rect 216 20250 256 20282
rect 288 20250 328 20282
rect 360 20250 400 20282
rect 432 20250 472 20282
rect 504 20250 544 20282
rect 576 20250 616 20282
rect 648 20250 688 20282
rect 720 20250 760 20282
rect 792 20250 832 20282
rect 864 20250 904 20282
rect 936 20250 976 20282
rect 1008 20250 1048 20282
rect 1080 20250 1120 20282
rect 1152 20250 1192 20282
rect 1224 20250 1264 20282
rect 1296 20250 1336 20282
rect 1368 20250 1408 20282
rect 1440 20250 1480 20282
rect 1512 20250 1552 20282
rect 1584 20250 1624 20282
rect 1656 20250 1696 20282
rect 1728 20250 1768 20282
rect 1800 20250 1840 20282
rect 1872 20250 1912 20282
rect 1944 20250 1984 20282
rect 2016 20250 2056 20282
rect 2088 20250 2128 20282
rect 2160 20250 2200 20282
rect 2232 20250 2272 20282
rect 2304 20250 2344 20282
rect 2376 20250 2416 20282
rect 2448 20250 2488 20282
rect 2520 20250 2560 20282
rect 2592 20250 2632 20282
rect 2664 20250 2704 20282
rect 2736 20250 2776 20282
rect 2808 20250 2848 20282
rect 2880 20250 2920 20282
rect 2952 20250 2992 20282
rect 3024 20250 3064 20282
rect 3096 20250 3136 20282
rect 3168 20250 3208 20282
rect 3240 20250 3280 20282
rect 3312 20250 3352 20282
rect 3384 20250 3424 20282
rect 3456 20250 3496 20282
rect 3528 20250 3568 20282
rect 3600 20250 3640 20282
rect 3672 20250 3712 20282
rect 3744 20250 3784 20282
rect 3816 20250 3856 20282
rect 3888 20250 3950 20282
rect 50 20210 3950 20250
rect 50 20178 112 20210
rect 144 20178 184 20210
rect 216 20178 256 20210
rect 288 20178 328 20210
rect 360 20178 400 20210
rect 432 20178 472 20210
rect 504 20178 544 20210
rect 576 20178 616 20210
rect 648 20178 688 20210
rect 720 20178 760 20210
rect 792 20178 832 20210
rect 864 20178 904 20210
rect 936 20178 976 20210
rect 1008 20178 1048 20210
rect 1080 20178 1120 20210
rect 1152 20178 1192 20210
rect 1224 20178 1264 20210
rect 1296 20178 1336 20210
rect 1368 20178 1408 20210
rect 1440 20178 1480 20210
rect 1512 20178 1552 20210
rect 1584 20178 1624 20210
rect 1656 20178 1696 20210
rect 1728 20178 1768 20210
rect 1800 20178 1840 20210
rect 1872 20178 1912 20210
rect 1944 20178 1984 20210
rect 2016 20178 2056 20210
rect 2088 20178 2128 20210
rect 2160 20178 2200 20210
rect 2232 20178 2272 20210
rect 2304 20178 2344 20210
rect 2376 20178 2416 20210
rect 2448 20178 2488 20210
rect 2520 20178 2560 20210
rect 2592 20178 2632 20210
rect 2664 20178 2704 20210
rect 2736 20178 2776 20210
rect 2808 20178 2848 20210
rect 2880 20178 2920 20210
rect 2952 20178 2992 20210
rect 3024 20178 3064 20210
rect 3096 20178 3136 20210
rect 3168 20178 3208 20210
rect 3240 20178 3280 20210
rect 3312 20178 3352 20210
rect 3384 20178 3424 20210
rect 3456 20178 3496 20210
rect 3528 20178 3568 20210
rect 3600 20178 3640 20210
rect 3672 20178 3712 20210
rect 3744 20178 3784 20210
rect 3816 20178 3856 20210
rect 3888 20178 3950 20210
rect 50 20138 3950 20178
rect 50 20106 112 20138
rect 144 20106 184 20138
rect 216 20106 256 20138
rect 288 20106 328 20138
rect 360 20106 400 20138
rect 432 20106 472 20138
rect 504 20106 544 20138
rect 576 20106 616 20138
rect 648 20106 688 20138
rect 720 20106 760 20138
rect 792 20106 832 20138
rect 864 20106 904 20138
rect 936 20106 976 20138
rect 1008 20106 1048 20138
rect 1080 20106 1120 20138
rect 1152 20106 1192 20138
rect 1224 20106 1264 20138
rect 1296 20106 1336 20138
rect 1368 20106 1408 20138
rect 1440 20106 1480 20138
rect 1512 20106 1552 20138
rect 1584 20106 1624 20138
rect 1656 20106 1696 20138
rect 1728 20106 1768 20138
rect 1800 20106 1840 20138
rect 1872 20106 1912 20138
rect 1944 20106 1984 20138
rect 2016 20106 2056 20138
rect 2088 20106 2128 20138
rect 2160 20106 2200 20138
rect 2232 20106 2272 20138
rect 2304 20106 2344 20138
rect 2376 20106 2416 20138
rect 2448 20106 2488 20138
rect 2520 20106 2560 20138
rect 2592 20106 2632 20138
rect 2664 20106 2704 20138
rect 2736 20106 2776 20138
rect 2808 20106 2848 20138
rect 2880 20106 2920 20138
rect 2952 20106 2992 20138
rect 3024 20106 3064 20138
rect 3096 20106 3136 20138
rect 3168 20106 3208 20138
rect 3240 20106 3280 20138
rect 3312 20106 3352 20138
rect 3384 20106 3424 20138
rect 3456 20106 3496 20138
rect 3528 20106 3568 20138
rect 3600 20106 3640 20138
rect 3672 20106 3712 20138
rect 3744 20106 3784 20138
rect 3816 20106 3856 20138
rect 3888 20106 3950 20138
rect 50 20066 3950 20106
rect 50 20034 112 20066
rect 144 20034 184 20066
rect 216 20034 256 20066
rect 288 20034 328 20066
rect 360 20034 400 20066
rect 432 20034 472 20066
rect 504 20034 544 20066
rect 576 20034 616 20066
rect 648 20034 688 20066
rect 720 20034 760 20066
rect 792 20034 832 20066
rect 864 20034 904 20066
rect 936 20034 976 20066
rect 1008 20034 1048 20066
rect 1080 20034 1120 20066
rect 1152 20034 1192 20066
rect 1224 20034 1264 20066
rect 1296 20034 1336 20066
rect 1368 20034 1408 20066
rect 1440 20034 1480 20066
rect 1512 20034 1552 20066
rect 1584 20034 1624 20066
rect 1656 20034 1696 20066
rect 1728 20034 1768 20066
rect 1800 20034 1840 20066
rect 1872 20034 1912 20066
rect 1944 20034 1984 20066
rect 2016 20034 2056 20066
rect 2088 20034 2128 20066
rect 2160 20034 2200 20066
rect 2232 20034 2272 20066
rect 2304 20034 2344 20066
rect 2376 20034 2416 20066
rect 2448 20034 2488 20066
rect 2520 20034 2560 20066
rect 2592 20034 2632 20066
rect 2664 20034 2704 20066
rect 2736 20034 2776 20066
rect 2808 20034 2848 20066
rect 2880 20034 2920 20066
rect 2952 20034 2992 20066
rect 3024 20034 3064 20066
rect 3096 20034 3136 20066
rect 3168 20034 3208 20066
rect 3240 20034 3280 20066
rect 3312 20034 3352 20066
rect 3384 20034 3424 20066
rect 3456 20034 3496 20066
rect 3528 20034 3568 20066
rect 3600 20034 3640 20066
rect 3672 20034 3712 20066
rect 3744 20034 3784 20066
rect 3816 20034 3856 20066
rect 3888 20034 3950 20066
rect 50 19994 3950 20034
rect 50 19962 112 19994
rect 144 19962 184 19994
rect 216 19962 256 19994
rect 288 19962 328 19994
rect 360 19962 400 19994
rect 432 19962 472 19994
rect 504 19962 544 19994
rect 576 19962 616 19994
rect 648 19962 688 19994
rect 720 19962 760 19994
rect 792 19962 832 19994
rect 864 19962 904 19994
rect 936 19962 976 19994
rect 1008 19962 1048 19994
rect 1080 19962 1120 19994
rect 1152 19962 1192 19994
rect 1224 19962 1264 19994
rect 1296 19962 1336 19994
rect 1368 19962 1408 19994
rect 1440 19962 1480 19994
rect 1512 19962 1552 19994
rect 1584 19962 1624 19994
rect 1656 19962 1696 19994
rect 1728 19962 1768 19994
rect 1800 19962 1840 19994
rect 1872 19962 1912 19994
rect 1944 19962 1984 19994
rect 2016 19962 2056 19994
rect 2088 19962 2128 19994
rect 2160 19962 2200 19994
rect 2232 19962 2272 19994
rect 2304 19962 2344 19994
rect 2376 19962 2416 19994
rect 2448 19962 2488 19994
rect 2520 19962 2560 19994
rect 2592 19962 2632 19994
rect 2664 19962 2704 19994
rect 2736 19962 2776 19994
rect 2808 19962 2848 19994
rect 2880 19962 2920 19994
rect 2952 19962 2992 19994
rect 3024 19962 3064 19994
rect 3096 19962 3136 19994
rect 3168 19962 3208 19994
rect 3240 19962 3280 19994
rect 3312 19962 3352 19994
rect 3384 19962 3424 19994
rect 3456 19962 3496 19994
rect 3528 19962 3568 19994
rect 3600 19962 3640 19994
rect 3672 19962 3712 19994
rect 3744 19962 3784 19994
rect 3816 19962 3856 19994
rect 3888 19962 3950 19994
rect 50 19922 3950 19962
rect 50 19890 112 19922
rect 144 19890 184 19922
rect 216 19890 256 19922
rect 288 19890 328 19922
rect 360 19890 400 19922
rect 432 19890 472 19922
rect 504 19890 544 19922
rect 576 19890 616 19922
rect 648 19890 688 19922
rect 720 19890 760 19922
rect 792 19890 832 19922
rect 864 19890 904 19922
rect 936 19890 976 19922
rect 1008 19890 1048 19922
rect 1080 19890 1120 19922
rect 1152 19890 1192 19922
rect 1224 19890 1264 19922
rect 1296 19890 1336 19922
rect 1368 19890 1408 19922
rect 1440 19890 1480 19922
rect 1512 19890 1552 19922
rect 1584 19890 1624 19922
rect 1656 19890 1696 19922
rect 1728 19890 1768 19922
rect 1800 19890 1840 19922
rect 1872 19890 1912 19922
rect 1944 19890 1984 19922
rect 2016 19890 2056 19922
rect 2088 19890 2128 19922
rect 2160 19890 2200 19922
rect 2232 19890 2272 19922
rect 2304 19890 2344 19922
rect 2376 19890 2416 19922
rect 2448 19890 2488 19922
rect 2520 19890 2560 19922
rect 2592 19890 2632 19922
rect 2664 19890 2704 19922
rect 2736 19890 2776 19922
rect 2808 19890 2848 19922
rect 2880 19890 2920 19922
rect 2952 19890 2992 19922
rect 3024 19890 3064 19922
rect 3096 19890 3136 19922
rect 3168 19890 3208 19922
rect 3240 19890 3280 19922
rect 3312 19890 3352 19922
rect 3384 19890 3424 19922
rect 3456 19890 3496 19922
rect 3528 19890 3568 19922
rect 3600 19890 3640 19922
rect 3672 19890 3712 19922
rect 3744 19890 3784 19922
rect 3816 19890 3856 19922
rect 3888 19890 3950 19922
rect 50 19850 3950 19890
rect 50 19818 112 19850
rect 144 19818 184 19850
rect 216 19818 256 19850
rect 288 19818 328 19850
rect 360 19818 400 19850
rect 432 19818 472 19850
rect 504 19818 544 19850
rect 576 19818 616 19850
rect 648 19818 688 19850
rect 720 19818 760 19850
rect 792 19818 832 19850
rect 864 19818 904 19850
rect 936 19818 976 19850
rect 1008 19818 1048 19850
rect 1080 19818 1120 19850
rect 1152 19818 1192 19850
rect 1224 19818 1264 19850
rect 1296 19818 1336 19850
rect 1368 19818 1408 19850
rect 1440 19818 1480 19850
rect 1512 19818 1552 19850
rect 1584 19818 1624 19850
rect 1656 19818 1696 19850
rect 1728 19818 1768 19850
rect 1800 19818 1840 19850
rect 1872 19818 1912 19850
rect 1944 19818 1984 19850
rect 2016 19818 2056 19850
rect 2088 19818 2128 19850
rect 2160 19818 2200 19850
rect 2232 19818 2272 19850
rect 2304 19818 2344 19850
rect 2376 19818 2416 19850
rect 2448 19818 2488 19850
rect 2520 19818 2560 19850
rect 2592 19818 2632 19850
rect 2664 19818 2704 19850
rect 2736 19818 2776 19850
rect 2808 19818 2848 19850
rect 2880 19818 2920 19850
rect 2952 19818 2992 19850
rect 3024 19818 3064 19850
rect 3096 19818 3136 19850
rect 3168 19818 3208 19850
rect 3240 19818 3280 19850
rect 3312 19818 3352 19850
rect 3384 19818 3424 19850
rect 3456 19818 3496 19850
rect 3528 19818 3568 19850
rect 3600 19818 3640 19850
rect 3672 19818 3712 19850
rect 3744 19818 3784 19850
rect 3816 19818 3856 19850
rect 3888 19818 3950 19850
rect 50 19778 3950 19818
rect 50 19746 112 19778
rect 144 19746 184 19778
rect 216 19746 256 19778
rect 288 19746 328 19778
rect 360 19746 400 19778
rect 432 19746 472 19778
rect 504 19746 544 19778
rect 576 19746 616 19778
rect 648 19746 688 19778
rect 720 19746 760 19778
rect 792 19746 832 19778
rect 864 19746 904 19778
rect 936 19746 976 19778
rect 1008 19746 1048 19778
rect 1080 19746 1120 19778
rect 1152 19746 1192 19778
rect 1224 19746 1264 19778
rect 1296 19746 1336 19778
rect 1368 19746 1408 19778
rect 1440 19746 1480 19778
rect 1512 19746 1552 19778
rect 1584 19746 1624 19778
rect 1656 19746 1696 19778
rect 1728 19746 1768 19778
rect 1800 19746 1840 19778
rect 1872 19746 1912 19778
rect 1944 19746 1984 19778
rect 2016 19746 2056 19778
rect 2088 19746 2128 19778
rect 2160 19746 2200 19778
rect 2232 19746 2272 19778
rect 2304 19746 2344 19778
rect 2376 19746 2416 19778
rect 2448 19746 2488 19778
rect 2520 19746 2560 19778
rect 2592 19746 2632 19778
rect 2664 19746 2704 19778
rect 2736 19746 2776 19778
rect 2808 19746 2848 19778
rect 2880 19746 2920 19778
rect 2952 19746 2992 19778
rect 3024 19746 3064 19778
rect 3096 19746 3136 19778
rect 3168 19746 3208 19778
rect 3240 19746 3280 19778
rect 3312 19746 3352 19778
rect 3384 19746 3424 19778
rect 3456 19746 3496 19778
rect 3528 19746 3568 19778
rect 3600 19746 3640 19778
rect 3672 19746 3712 19778
rect 3744 19746 3784 19778
rect 3816 19746 3856 19778
rect 3888 19746 3950 19778
rect 50 19706 3950 19746
rect 50 19674 112 19706
rect 144 19674 184 19706
rect 216 19674 256 19706
rect 288 19674 328 19706
rect 360 19674 400 19706
rect 432 19674 472 19706
rect 504 19674 544 19706
rect 576 19674 616 19706
rect 648 19674 688 19706
rect 720 19674 760 19706
rect 792 19674 832 19706
rect 864 19674 904 19706
rect 936 19674 976 19706
rect 1008 19674 1048 19706
rect 1080 19674 1120 19706
rect 1152 19674 1192 19706
rect 1224 19674 1264 19706
rect 1296 19674 1336 19706
rect 1368 19674 1408 19706
rect 1440 19674 1480 19706
rect 1512 19674 1552 19706
rect 1584 19674 1624 19706
rect 1656 19674 1696 19706
rect 1728 19674 1768 19706
rect 1800 19674 1840 19706
rect 1872 19674 1912 19706
rect 1944 19674 1984 19706
rect 2016 19674 2056 19706
rect 2088 19674 2128 19706
rect 2160 19674 2200 19706
rect 2232 19674 2272 19706
rect 2304 19674 2344 19706
rect 2376 19674 2416 19706
rect 2448 19674 2488 19706
rect 2520 19674 2560 19706
rect 2592 19674 2632 19706
rect 2664 19674 2704 19706
rect 2736 19674 2776 19706
rect 2808 19674 2848 19706
rect 2880 19674 2920 19706
rect 2952 19674 2992 19706
rect 3024 19674 3064 19706
rect 3096 19674 3136 19706
rect 3168 19674 3208 19706
rect 3240 19674 3280 19706
rect 3312 19674 3352 19706
rect 3384 19674 3424 19706
rect 3456 19674 3496 19706
rect 3528 19674 3568 19706
rect 3600 19674 3640 19706
rect 3672 19674 3712 19706
rect 3744 19674 3784 19706
rect 3816 19674 3856 19706
rect 3888 19674 3950 19706
rect 50 19634 3950 19674
rect 50 19602 112 19634
rect 144 19602 184 19634
rect 216 19602 256 19634
rect 288 19602 328 19634
rect 360 19602 400 19634
rect 432 19602 472 19634
rect 504 19602 544 19634
rect 576 19602 616 19634
rect 648 19602 688 19634
rect 720 19602 760 19634
rect 792 19602 832 19634
rect 864 19602 904 19634
rect 936 19602 976 19634
rect 1008 19602 1048 19634
rect 1080 19602 1120 19634
rect 1152 19602 1192 19634
rect 1224 19602 1264 19634
rect 1296 19602 1336 19634
rect 1368 19602 1408 19634
rect 1440 19602 1480 19634
rect 1512 19602 1552 19634
rect 1584 19602 1624 19634
rect 1656 19602 1696 19634
rect 1728 19602 1768 19634
rect 1800 19602 1840 19634
rect 1872 19602 1912 19634
rect 1944 19602 1984 19634
rect 2016 19602 2056 19634
rect 2088 19602 2128 19634
rect 2160 19602 2200 19634
rect 2232 19602 2272 19634
rect 2304 19602 2344 19634
rect 2376 19602 2416 19634
rect 2448 19602 2488 19634
rect 2520 19602 2560 19634
rect 2592 19602 2632 19634
rect 2664 19602 2704 19634
rect 2736 19602 2776 19634
rect 2808 19602 2848 19634
rect 2880 19602 2920 19634
rect 2952 19602 2992 19634
rect 3024 19602 3064 19634
rect 3096 19602 3136 19634
rect 3168 19602 3208 19634
rect 3240 19602 3280 19634
rect 3312 19602 3352 19634
rect 3384 19602 3424 19634
rect 3456 19602 3496 19634
rect 3528 19602 3568 19634
rect 3600 19602 3640 19634
rect 3672 19602 3712 19634
rect 3744 19602 3784 19634
rect 3816 19602 3856 19634
rect 3888 19602 3950 19634
rect 50 19562 3950 19602
rect 50 19530 112 19562
rect 144 19530 184 19562
rect 216 19530 256 19562
rect 288 19530 328 19562
rect 360 19530 400 19562
rect 432 19530 472 19562
rect 504 19530 544 19562
rect 576 19530 616 19562
rect 648 19530 688 19562
rect 720 19530 760 19562
rect 792 19530 832 19562
rect 864 19530 904 19562
rect 936 19530 976 19562
rect 1008 19530 1048 19562
rect 1080 19530 1120 19562
rect 1152 19530 1192 19562
rect 1224 19530 1264 19562
rect 1296 19530 1336 19562
rect 1368 19530 1408 19562
rect 1440 19530 1480 19562
rect 1512 19530 1552 19562
rect 1584 19530 1624 19562
rect 1656 19530 1696 19562
rect 1728 19530 1768 19562
rect 1800 19530 1840 19562
rect 1872 19530 1912 19562
rect 1944 19530 1984 19562
rect 2016 19530 2056 19562
rect 2088 19530 2128 19562
rect 2160 19530 2200 19562
rect 2232 19530 2272 19562
rect 2304 19530 2344 19562
rect 2376 19530 2416 19562
rect 2448 19530 2488 19562
rect 2520 19530 2560 19562
rect 2592 19530 2632 19562
rect 2664 19530 2704 19562
rect 2736 19530 2776 19562
rect 2808 19530 2848 19562
rect 2880 19530 2920 19562
rect 2952 19530 2992 19562
rect 3024 19530 3064 19562
rect 3096 19530 3136 19562
rect 3168 19530 3208 19562
rect 3240 19530 3280 19562
rect 3312 19530 3352 19562
rect 3384 19530 3424 19562
rect 3456 19530 3496 19562
rect 3528 19530 3568 19562
rect 3600 19530 3640 19562
rect 3672 19530 3712 19562
rect 3744 19530 3784 19562
rect 3816 19530 3856 19562
rect 3888 19530 3950 19562
rect 50 19490 3950 19530
rect 50 19458 112 19490
rect 144 19458 184 19490
rect 216 19458 256 19490
rect 288 19458 328 19490
rect 360 19458 400 19490
rect 432 19458 472 19490
rect 504 19458 544 19490
rect 576 19458 616 19490
rect 648 19458 688 19490
rect 720 19458 760 19490
rect 792 19458 832 19490
rect 864 19458 904 19490
rect 936 19458 976 19490
rect 1008 19458 1048 19490
rect 1080 19458 1120 19490
rect 1152 19458 1192 19490
rect 1224 19458 1264 19490
rect 1296 19458 1336 19490
rect 1368 19458 1408 19490
rect 1440 19458 1480 19490
rect 1512 19458 1552 19490
rect 1584 19458 1624 19490
rect 1656 19458 1696 19490
rect 1728 19458 1768 19490
rect 1800 19458 1840 19490
rect 1872 19458 1912 19490
rect 1944 19458 1984 19490
rect 2016 19458 2056 19490
rect 2088 19458 2128 19490
rect 2160 19458 2200 19490
rect 2232 19458 2272 19490
rect 2304 19458 2344 19490
rect 2376 19458 2416 19490
rect 2448 19458 2488 19490
rect 2520 19458 2560 19490
rect 2592 19458 2632 19490
rect 2664 19458 2704 19490
rect 2736 19458 2776 19490
rect 2808 19458 2848 19490
rect 2880 19458 2920 19490
rect 2952 19458 2992 19490
rect 3024 19458 3064 19490
rect 3096 19458 3136 19490
rect 3168 19458 3208 19490
rect 3240 19458 3280 19490
rect 3312 19458 3352 19490
rect 3384 19458 3424 19490
rect 3456 19458 3496 19490
rect 3528 19458 3568 19490
rect 3600 19458 3640 19490
rect 3672 19458 3712 19490
rect 3744 19458 3784 19490
rect 3816 19458 3856 19490
rect 3888 19458 3950 19490
rect 50 19418 3950 19458
rect 50 19386 112 19418
rect 144 19386 184 19418
rect 216 19386 256 19418
rect 288 19386 328 19418
rect 360 19386 400 19418
rect 432 19386 472 19418
rect 504 19386 544 19418
rect 576 19386 616 19418
rect 648 19386 688 19418
rect 720 19386 760 19418
rect 792 19386 832 19418
rect 864 19386 904 19418
rect 936 19386 976 19418
rect 1008 19386 1048 19418
rect 1080 19386 1120 19418
rect 1152 19386 1192 19418
rect 1224 19386 1264 19418
rect 1296 19386 1336 19418
rect 1368 19386 1408 19418
rect 1440 19386 1480 19418
rect 1512 19386 1552 19418
rect 1584 19386 1624 19418
rect 1656 19386 1696 19418
rect 1728 19386 1768 19418
rect 1800 19386 1840 19418
rect 1872 19386 1912 19418
rect 1944 19386 1984 19418
rect 2016 19386 2056 19418
rect 2088 19386 2128 19418
rect 2160 19386 2200 19418
rect 2232 19386 2272 19418
rect 2304 19386 2344 19418
rect 2376 19386 2416 19418
rect 2448 19386 2488 19418
rect 2520 19386 2560 19418
rect 2592 19386 2632 19418
rect 2664 19386 2704 19418
rect 2736 19386 2776 19418
rect 2808 19386 2848 19418
rect 2880 19386 2920 19418
rect 2952 19386 2992 19418
rect 3024 19386 3064 19418
rect 3096 19386 3136 19418
rect 3168 19386 3208 19418
rect 3240 19386 3280 19418
rect 3312 19386 3352 19418
rect 3384 19386 3424 19418
rect 3456 19386 3496 19418
rect 3528 19386 3568 19418
rect 3600 19386 3640 19418
rect 3672 19386 3712 19418
rect 3744 19386 3784 19418
rect 3816 19386 3856 19418
rect 3888 19386 3950 19418
rect 50 19346 3950 19386
rect 50 19314 112 19346
rect 144 19314 184 19346
rect 216 19314 256 19346
rect 288 19314 328 19346
rect 360 19314 400 19346
rect 432 19314 472 19346
rect 504 19314 544 19346
rect 576 19314 616 19346
rect 648 19314 688 19346
rect 720 19314 760 19346
rect 792 19314 832 19346
rect 864 19314 904 19346
rect 936 19314 976 19346
rect 1008 19314 1048 19346
rect 1080 19314 1120 19346
rect 1152 19314 1192 19346
rect 1224 19314 1264 19346
rect 1296 19314 1336 19346
rect 1368 19314 1408 19346
rect 1440 19314 1480 19346
rect 1512 19314 1552 19346
rect 1584 19314 1624 19346
rect 1656 19314 1696 19346
rect 1728 19314 1768 19346
rect 1800 19314 1840 19346
rect 1872 19314 1912 19346
rect 1944 19314 1984 19346
rect 2016 19314 2056 19346
rect 2088 19314 2128 19346
rect 2160 19314 2200 19346
rect 2232 19314 2272 19346
rect 2304 19314 2344 19346
rect 2376 19314 2416 19346
rect 2448 19314 2488 19346
rect 2520 19314 2560 19346
rect 2592 19314 2632 19346
rect 2664 19314 2704 19346
rect 2736 19314 2776 19346
rect 2808 19314 2848 19346
rect 2880 19314 2920 19346
rect 2952 19314 2992 19346
rect 3024 19314 3064 19346
rect 3096 19314 3136 19346
rect 3168 19314 3208 19346
rect 3240 19314 3280 19346
rect 3312 19314 3352 19346
rect 3384 19314 3424 19346
rect 3456 19314 3496 19346
rect 3528 19314 3568 19346
rect 3600 19314 3640 19346
rect 3672 19314 3712 19346
rect 3744 19314 3784 19346
rect 3816 19314 3856 19346
rect 3888 19314 3950 19346
rect 50 19274 3950 19314
rect 50 19242 112 19274
rect 144 19242 184 19274
rect 216 19242 256 19274
rect 288 19242 328 19274
rect 360 19242 400 19274
rect 432 19242 472 19274
rect 504 19242 544 19274
rect 576 19242 616 19274
rect 648 19242 688 19274
rect 720 19242 760 19274
rect 792 19242 832 19274
rect 864 19242 904 19274
rect 936 19242 976 19274
rect 1008 19242 1048 19274
rect 1080 19242 1120 19274
rect 1152 19242 1192 19274
rect 1224 19242 1264 19274
rect 1296 19242 1336 19274
rect 1368 19242 1408 19274
rect 1440 19242 1480 19274
rect 1512 19242 1552 19274
rect 1584 19242 1624 19274
rect 1656 19242 1696 19274
rect 1728 19242 1768 19274
rect 1800 19242 1840 19274
rect 1872 19242 1912 19274
rect 1944 19242 1984 19274
rect 2016 19242 2056 19274
rect 2088 19242 2128 19274
rect 2160 19242 2200 19274
rect 2232 19242 2272 19274
rect 2304 19242 2344 19274
rect 2376 19242 2416 19274
rect 2448 19242 2488 19274
rect 2520 19242 2560 19274
rect 2592 19242 2632 19274
rect 2664 19242 2704 19274
rect 2736 19242 2776 19274
rect 2808 19242 2848 19274
rect 2880 19242 2920 19274
rect 2952 19242 2992 19274
rect 3024 19242 3064 19274
rect 3096 19242 3136 19274
rect 3168 19242 3208 19274
rect 3240 19242 3280 19274
rect 3312 19242 3352 19274
rect 3384 19242 3424 19274
rect 3456 19242 3496 19274
rect 3528 19242 3568 19274
rect 3600 19242 3640 19274
rect 3672 19242 3712 19274
rect 3744 19242 3784 19274
rect 3816 19242 3856 19274
rect 3888 19242 3950 19274
rect 50 19202 3950 19242
rect 50 19170 112 19202
rect 144 19170 184 19202
rect 216 19170 256 19202
rect 288 19170 328 19202
rect 360 19170 400 19202
rect 432 19170 472 19202
rect 504 19170 544 19202
rect 576 19170 616 19202
rect 648 19170 688 19202
rect 720 19170 760 19202
rect 792 19170 832 19202
rect 864 19170 904 19202
rect 936 19170 976 19202
rect 1008 19170 1048 19202
rect 1080 19170 1120 19202
rect 1152 19170 1192 19202
rect 1224 19170 1264 19202
rect 1296 19170 1336 19202
rect 1368 19170 1408 19202
rect 1440 19170 1480 19202
rect 1512 19170 1552 19202
rect 1584 19170 1624 19202
rect 1656 19170 1696 19202
rect 1728 19170 1768 19202
rect 1800 19170 1840 19202
rect 1872 19170 1912 19202
rect 1944 19170 1984 19202
rect 2016 19170 2056 19202
rect 2088 19170 2128 19202
rect 2160 19170 2200 19202
rect 2232 19170 2272 19202
rect 2304 19170 2344 19202
rect 2376 19170 2416 19202
rect 2448 19170 2488 19202
rect 2520 19170 2560 19202
rect 2592 19170 2632 19202
rect 2664 19170 2704 19202
rect 2736 19170 2776 19202
rect 2808 19170 2848 19202
rect 2880 19170 2920 19202
rect 2952 19170 2992 19202
rect 3024 19170 3064 19202
rect 3096 19170 3136 19202
rect 3168 19170 3208 19202
rect 3240 19170 3280 19202
rect 3312 19170 3352 19202
rect 3384 19170 3424 19202
rect 3456 19170 3496 19202
rect 3528 19170 3568 19202
rect 3600 19170 3640 19202
rect 3672 19170 3712 19202
rect 3744 19170 3784 19202
rect 3816 19170 3856 19202
rect 3888 19170 3950 19202
rect 50 19130 3950 19170
rect 50 19098 112 19130
rect 144 19098 184 19130
rect 216 19098 256 19130
rect 288 19098 328 19130
rect 360 19098 400 19130
rect 432 19098 472 19130
rect 504 19098 544 19130
rect 576 19098 616 19130
rect 648 19098 688 19130
rect 720 19098 760 19130
rect 792 19098 832 19130
rect 864 19098 904 19130
rect 936 19098 976 19130
rect 1008 19098 1048 19130
rect 1080 19098 1120 19130
rect 1152 19098 1192 19130
rect 1224 19098 1264 19130
rect 1296 19098 1336 19130
rect 1368 19098 1408 19130
rect 1440 19098 1480 19130
rect 1512 19098 1552 19130
rect 1584 19098 1624 19130
rect 1656 19098 1696 19130
rect 1728 19098 1768 19130
rect 1800 19098 1840 19130
rect 1872 19098 1912 19130
rect 1944 19098 1984 19130
rect 2016 19098 2056 19130
rect 2088 19098 2128 19130
rect 2160 19098 2200 19130
rect 2232 19098 2272 19130
rect 2304 19098 2344 19130
rect 2376 19098 2416 19130
rect 2448 19098 2488 19130
rect 2520 19098 2560 19130
rect 2592 19098 2632 19130
rect 2664 19098 2704 19130
rect 2736 19098 2776 19130
rect 2808 19098 2848 19130
rect 2880 19098 2920 19130
rect 2952 19098 2992 19130
rect 3024 19098 3064 19130
rect 3096 19098 3136 19130
rect 3168 19098 3208 19130
rect 3240 19098 3280 19130
rect 3312 19098 3352 19130
rect 3384 19098 3424 19130
rect 3456 19098 3496 19130
rect 3528 19098 3568 19130
rect 3600 19098 3640 19130
rect 3672 19098 3712 19130
rect 3744 19098 3784 19130
rect 3816 19098 3856 19130
rect 3888 19098 3950 19130
rect 50 19058 3950 19098
rect 50 19026 112 19058
rect 144 19026 184 19058
rect 216 19026 256 19058
rect 288 19026 328 19058
rect 360 19026 400 19058
rect 432 19026 472 19058
rect 504 19026 544 19058
rect 576 19026 616 19058
rect 648 19026 688 19058
rect 720 19026 760 19058
rect 792 19026 832 19058
rect 864 19026 904 19058
rect 936 19026 976 19058
rect 1008 19026 1048 19058
rect 1080 19026 1120 19058
rect 1152 19026 1192 19058
rect 1224 19026 1264 19058
rect 1296 19026 1336 19058
rect 1368 19026 1408 19058
rect 1440 19026 1480 19058
rect 1512 19026 1552 19058
rect 1584 19026 1624 19058
rect 1656 19026 1696 19058
rect 1728 19026 1768 19058
rect 1800 19026 1840 19058
rect 1872 19026 1912 19058
rect 1944 19026 1984 19058
rect 2016 19026 2056 19058
rect 2088 19026 2128 19058
rect 2160 19026 2200 19058
rect 2232 19026 2272 19058
rect 2304 19026 2344 19058
rect 2376 19026 2416 19058
rect 2448 19026 2488 19058
rect 2520 19026 2560 19058
rect 2592 19026 2632 19058
rect 2664 19026 2704 19058
rect 2736 19026 2776 19058
rect 2808 19026 2848 19058
rect 2880 19026 2920 19058
rect 2952 19026 2992 19058
rect 3024 19026 3064 19058
rect 3096 19026 3136 19058
rect 3168 19026 3208 19058
rect 3240 19026 3280 19058
rect 3312 19026 3352 19058
rect 3384 19026 3424 19058
rect 3456 19026 3496 19058
rect 3528 19026 3568 19058
rect 3600 19026 3640 19058
rect 3672 19026 3712 19058
rect 3744 19026 3784 19058
rect 3816 19026 3856 19058
rect 3888 19026 3950 19058
rect 50 18986 3950 19026
rect 50 18954 112 18986
rect 144 18954 184 18986
rect 216 18954 256 18986
rect 288 18954 328 18986
rect 360 18954 400 18986
rect 432 18954 472 18986
rect 504 18954 544 18986
rect 576 18954 616 18986
rect 648 18954 688 18986
rect 720 18954 760 18986
rect 792 18954 832 18986
rect 864 18954 904 18986
rect 936 18954 976 18986
rect 1008 18954 1048 18986
rect 1080 18954 1120 18986
rect 1152 18954 1192 18986
rect 1224 18954 1264 18986
rect 1296 18954 1336 18986
rect 1368 18954 1408 18986
rect 1440 18954 1480 18986
rect 1512 18954 1552 18986
rect 1584 18954 1624 18986
rect 1656 18954 1696 18986
rect 1728 18954 1768 18986
rect 1800 18954 1840 18986
rect 1872 18954 1912 18986
rect 1944 18954 1984 18986
rect 2016 18954 2056 18986
rect 2088 18954 2128 18986
rect 2160 18954 2200 18986
rect 2232 18954 2272 18986
rect 2304 18954 2344 18986
rect 2376 18954 2416 18986
rect 2448 18954 2488 18986
rect 2520 18954 2560 18986
rect 2592 18954 2632 18986
rect 2664 18954 2704 18986
rect 2736 18954 2776 18986
rect 2808 18954 2848 18986
rect 2880 18954 2920 18986
rect 2952 18954 2992 18986
rect 3024 18954 3064 18986
rect 3096 18954 3136 18986
rect 3168 18954 3208 18986
rect 3240 18954 3280 18986
rect 3312 18954 3352 18986
rect 3384 18954 3424 18986
rect 3456 18954 3496 18986
rect 3528 18954 3568 18986
rect 3600 18954 3640 18986
rect 3672 18954 3712 18986
rect 3744 18954 3784 18986
rect 3816 18954 3856 18986
rect 3888 18954 3950 18986
rect 50 18914 3950 18954
rect 50 18882 112 18914
rect 144 18882 184 18914
rect 216 18882 256 18914
rect 288 18882 328 18914
rect 360 18882 400 18914
rect 432 18882 472 18914
rect 504 18882 544 18914
rect 576 18882 616 18914
rect 648 18882 688 18914
rect 720 18882 760 18914
rect 792 18882 832 18914
rect 864 18882 904 18914
rect 936 18882 976 18914
rect 1008 18882 1048 18914
rect 1080 18882 1120 18914
rect 1152 18882 1192 18914
rect 1224 18882 1264 18914
rect 1296 18882 1336 18914
rect 1368 18882 1408 18914
rect 1440 18882 1480 18914
rect 1512 18882 1552 18914
rect 1584 18882 1624 18914
rect 1656 18882 1696 18914
rect 1728 18882 1768 18914
rect 1800 18882 1840 18914
rect 1872 18882 1912 18914
rect 1944 18882 1984 18914
rect 2016 18882 2056 18914
rect 2088 18882 2128 18914
rect 2160 18882 2200 18914
rect 2232 18882 2272 18914
rect 2304 18882 2344 18914
rect 2376 18882 2416 18914
rect 2448 18882 2488 18914
rect 2520 18882 2560 18914
rect 2592 18882 2632 18914
rect 2664 18882 2704 18914
rect 2736 18882 2776 18914
rect 2808 18882 2848 18914
rect 2880 18882 2920 18914
rect 2952 18882 2992 18914
rect 3024 18882 3064 18914
rect 3096 18882 3136 18914
rect 3168 18882 3208 18914
rect 3240 18882 3280 18914
rect 3312 18882 3352 18914
rect 3384 18882 3424 18914
rect 3456 18882 3496 18914
rect 3528 18882 3568 18914
rect 3600 18882 3640 18914
rect 3672 18882 3712 18914
rect 3744 18882 3784 18914
rect 3816 18882 3856 18914
rect 3888 18882 3950 18914
rect 50 18842 3950 18882
rect 50 18810 112 18842
rect 144 18810 184 18842
rect 216 18810 256 18842
rect 288 18810 328 18842
rect 360 18810 400 18842
rect 432 18810 472 18842
rect 504 18810 544 18842
rect 576 18810 616 18842
rect 648 18810 688 18842
rect 720 18810 760 18842
rect 792 18810 832 18842
rect 864 18810 904 18842
rect 936 18810 976 18842
rect 1008 18810 1048 18842
rect 1080 18810 1120 18842
rect 1152 18810 1192 18842
rect 1224 18810 1264 18842
rect 1296 18810 1336 18842
rect 1368 18810 1408 18842
rect 1440 18810 1480 18842
rect 1512 18810 1552 18842
rect 1584 18810 1624 18842
rect 1656 18810 1696 18842
rect 1728 18810 1768 18842
rect 1800 18810 1840 18842
rect 1872 18810 1912 18842
rect 1944 18810 1984 18842
rect 2016 18810 2056 18842
rect 2088 18810 2128 18842
rect 2160 18810 2200 18842
rect 2232 18810 2272 18842
rect 2304 18810 2344 18842
rect 2376 18810 2416 18842
rect 2448 18810 2488 18842
rect 2520 18810 2560 18842
rect 2592 18810 2632 18842
rect 2664 18810 2704 18842
rect 2736 18810 2776 18842
rect 2808 18810 2848 18842
rect 2880 18810 2920 18842
rect 2952 18810 2992 18842
rect 3024 18810 3064 18842
rect 3096 18810 3136 18842
rect 3168 18810 3208 18842
rect 3240 18810 3280 18842
rect 3312 18810 3352 18842
rect 3384 18810 3424 18842
rect 3456 18810 3496 18842
rect 3528 18810 3568 18842
rect 3600 18810 3640 18842
rect 3672 18810 3712 18842
rect 3744 18810 3784 18842
rect 3816 18810 3856 18842
rect 3888 18810 3950 18842
rect 50 18770 3950 18810
rect 50 18738 112 18770
rect 144 18738 184 18770
rect 216 18738 256 18770
rect 288 18738 328 18770
rect 360 18738 400 18770
rect 432 18738 472 18770
rect 504 18738 544 18770
rect 576 18738 616 18770
rect 648 18738 688 18770
rect 720 18738 760 18770
rect 792 18738 832 18770
rect 864 18738 904 18770
rect 936 18738 976 18770
rect 1008 18738 1048 18770
rect 1080 18738 1120 18770
rect 1152 18738 1192 18770
rect 1224 18738 1264 18770
rect 1296 18738 1336 18770
rect 1368 18738 1408 18770
rect 1440 18738 1480 18770
rect 1512 18738 1552 18770
rect 1584 18738 1624 18770
rect 1656 18738 1696 18770
rect 1728 18738 1768 18770
rect 1800 18738 1840 18770
rect 1872 18738 1912 18770
rect 1944 18738 1984 18770
rect 2016 18738 2056 18770
rect 2088 18738 2128 18770
rect 2160 18738 2200 18770
rect 2232 18738 2272 18770
rect 2304 18738 2344 18770
rect 2376 18738 2416 18770
rect 2448 18738 2488 18770
rect 2520 18738 2560 18770
rect 2592 18738 2632 18770
rect 2664 18738 2704 18770
rect 2736 18738 2776 18770
rect 2808 18738 2848 18770
rect 2880 18738 2920 18770
rect 2952 18738 2992 18770
rect 3024 18738 3064 18770
rect 3096 18738 3136 18770
rect 3168 18738 3208 18770
rect 3240 18738 3280 18770
rect 3312 18738 3352 18770
rect 3384 18738 3424 18770
rect 3456 18738 3496 18770
rect 3528 18738 3568 18770
rect 3600 18738 3640 18770
rect 3672 18738 3712 18770
rect 3744 18738 3784 18770
rect 3816 18738 3856 18770
rect 3888 18738 3950 18770
rect 50 18698 3950 18738
rect 50 18666 112 18698
rect 144 18666 184 18698
rect 216 18666 256 18698
rect 288 18666 328 18698
rect 360 18666 400 18698
rect 432 18666 472 18698
rect 504 18666 544 18698
rect 576 18666 616 18698
rect 648 18666 688 18698
rect 720 18666 760 18698
rect 792 18666 832 18698
rect 864 18666 904 18698
rect 936 18666 976 18698
rect 1008 18666 1048 18698
rect 1080 18666 1120 18698
rect 1152 18666 1192 18698
rect 1224 18666 1264 18698
rect 1296 18666 1336 18698
rect 1368 18666 1408 18698
rect 1440 18666 1480 18698
rect 1512 18666 1552 18698
rect 1584 18666 1624 18698
rect 1656 18666 1696 18698
rect 1728 18666 1768 18698
rect 1800 18666 1840 18698
rect 1872 18666 1912 18698
rect 1944 18666 1984 18698
rect 2016 18666 2056 18698
rect 2088 18666 2128 18698
rect 2160 18666 2200 18698
rect 2232 18666 2272 18698
rect 2304 18666 2344 18698
rect 2376 18666 2416 18698
rect 2448 18666 2488 18698
rect 2520 18666 2560 18698
rect 2592 18666 2632 18698
rect 2664 18666 2704 18698
rect 2736 18666 2776 18698
rect 2808 18666 2848 18698
rect 2880 18666 2920 18698
rect 2952 18666 2992 18698
rect 3024 18666 3064 18698
rect 3096 18666 3136 18698
rect 3168 18666 3208 18698
rect 3240 18666 3280 18698
rect 3312 18666 3352 18698
rect 3384 18666 3424 18698
rect 3456 18666 3496 18698
rect 3528 18666 3568 18698
rect 3600 18666 3640 18698
rect 3672 18666 3712 18698
rect 3744 18666 3784 18698
rect 3816 18666 3856 18698
rect 3888 18666 3950 18698
rect 50 18626 3950 18666
rect 50 18594 112 18626
rect 144 18594 184 18626
rect 216 18594 256 18626
rect 288 18594 328 18626
rect 360 18594 400 18626
rect 432 18594 472 18626
rect 504 18594 544 18626
rect 576 18594 616 18626
rect 648 18594 688 18626
rect 720 18594 760 18626
rect 792 18594 832 18626
rect 864 18594 904 18626
rect 936 18594 976 18626
rect 1008 18594 1048 18626
rect 1080 18594 1120 18626
rect 1152 18594 1192 18626
rect 1224 18594 1264 18626
rect 1296 18594 1336 18626
rect 1368 18594 1408 18626
rect 1440 18594 1480 18626
rect 1512 18594 1552 18626
rect 1584 18594 1624 18626
rect 1656 18594 1696 18626
rect 1728 18594 1768 18626
rect 1800 18594 1840 18626
rect 1872 18594 1912 18626
rect 1944 18594 1984 18626
rect 2016 18594 2056 18626
rect 2088 18594 2128 18626
rect 2160 18594 2200 18626
rect 2232 18594 2272 18626
rect 2304 18594 2344 18626
rect 2376 18594 2416 18626
rect 2448 18594 2488 18626
rect 2520 18594 2560 18626
rect 2592 18594 2632 18626
rect 2664 18594 2704 18626
rect 2736 18594 2776 18626
rect 2808 18594 2848 18626
rect 2880 18594 2920 18626
rect 2952 18594 2992 18626
rect 3024 18594 3064 18626
rect 3096 18594 3136 18626
rect 3168 18594 3208 18626
rect 3240 18594 3280 18626
rect 3312 18594 3352 18626
rect 3384 18594 3424 18626
rect 3456 18594 3496 18626
rect 3528 18594 3568 18626
rect 3600 18594 3640 18626
rect 3672 18594 3712 18626
rect 3744 18594 3784 18626
rect 3816 18594 3856 18626
rect 3888 18594 3950 18626
rect 50 18554 3950 18594
rect 50 18522 112 18554
rect 144 18522 184 18554
rect 216 18522 256 18554
rect 288 18522 328 18554
rect 360 18522 400 18554
rect 432 18522 472 18554
rect 504 18522 544 18554
rect 576 18522 616 18554
rect 648 18522 688 18554
rect 720 18522 760 18554
rect 792 18522 832 18554
rect 864 18522 904 18554
rect 936 18522 976 18554
rect 1008 18522 1048 18554
rect 1080 18522 1120 18554
rect 1152 18522 1192 18554
rect 1224 18522 1264 18554
rect 1296 18522 1336 18554
rect 1368 18522 1408 18554
rect 1440 18522 1480 18554
rect 1512 18522 1552 18554
rect 1584 18522 1624 18554
rect 1656 18522 1696 18554
rect 1728 18522 1768 18554
rect 1800 18522 1840 18554
rect 1872 18522 1912 18554
rect 1944 18522 1984 18554
rect 2016 18522 2056 18554
rect 2088 18522 2128 18554
rect 2160 18522 2200 18554
rect 2232 18522 2272 18554
rect 2304 18522 2344 18554
rect 2376 18522 2416 18554
rect 2448 18522 2488 18554
rect 2520 18522 2560 18554
rect 2592 18522 2632 18554
rect 2664 18522 2704 18554
rect 2736 18522 2776 18554
rect 2808 18522 2848 18554
rect 2880 18522 2920 18554
rect 2952 18522 2992 18554
rect 3024 18522 3064 18554
rect 3096 18522 3136 18554
rect 3168 18522 3208 18554
rect 3240 18522 3280 18554
rect 3312 18522 3352 18554
rect 3384 18522 3424 18554
rect 3456 18522 3496 18554
rect 3528 18522 3568 18554
rect 3600 18522 3640 18554
rect 3672 18522 3712 18554
rect 3744 18522 3784 18554
rect 3816 18522 3856 18554
rect 3888 18522 3950 18554
rect 50 18482 3950 18522
rect 50 18450 112 18482
rect 144 18450 184 18482
rect 216 18450 256 18482
rect 288 18450 328 18482
rect 360 18450 400 18482
rect 432 18450 472 18482
rect 504 18450 544 18482
rect 576 18450 616 18482
rect 648 18450 688 18482
rect 720 18450 760 18482
rect 792 18450 832 18482
rect 864 18450 904 18482
rect 936 18450 976 18482
rect 1008 18450 1048 18482
rect 1080 18450 1120 18482
rect 1152 18450 1192 18482
rect 1224 18450 1264 18482
rect 1296 18450 1336 18482
rect 1368 18450 1408 18482
rect 1440 18450 1480 18482
rect 1512 18450 1552 18482
rect 1584 18450 1624 18482
rect 1656 18450 1696 18482
rect 1728 18450 1768 18482
rect 1800 18450 1840 18482
rect 1872 18450 1912 18482
rect 1944 18450 1984 18482
rect 2016 18450 2056 18482
rect 2088 18450 2128 18482
rect 2160 18450 2200 18482
rect 2232 18450 2272 18482
rect 2304 18450 2344 18482
rect 2376 18450 2416 18482
rect 2448 18450 2488 18482
rect 2520 18450 2560 18482
rect 2592 18450 2632 18482
rect 2664 18450 2704 18482
rect 2736 18450 2776 18482
rect 2808 18450 2848 18482
rect 2880 18450 2920 18482
rect 2952 18450 2992 18482
rect 3024 18450 3064 18482
rect 3096 18450 3136 18482
rect 3168 18450 3208 18482
rect 3240 18450 3280 18482
rect 3312 18450 3352 18482
rect 3384 18450 3424 18482
rect 3456 18450 3496 18482
rect 3528 18450 3568 18482
rect 3600 18450 3640 18482
rect 3672 18450 3712 18482
rect 3744 18450 3784 18482
rect 3816 18450 3856 18482
rect 3888 18450 3950 18482
rect 50 18410 3950 18450
rect 50 18378 112 18410
rect 144 18378 184 18410
rect 216 18378 256 18410
rect 288 18378 328 18410
rect 360 18378 400 18410
rect 432 18378 472 18410
rect 504 18378 544 18410
rect 576 18378 616 18410
rect 648 18378 688 18410
rect 720 18378 760 18410
rect 792 18378 832 18410
rect 864 18378 904 18410
rect 936 18378 976 18410
rect 1008 18378 1048 18410
rect 1080 18378 1120 18410
rect 1152 18378 1192 18410
rect 1224 18378 1264 18410
rect 1296 18378 1336 18410
rect 1368 18378 1408 18410
rect 1440 18378 1480 18410
rect 1512 18378 1552 18410
rect 1584 18378 1624 18410
rect 1656 18378 1696 18410
rect 1728 18378 1768 18410
rect 1800 18378 1840 18410
rect 1872 18378 1912 18410
rect 1944 18378 1984 18410
rect 2016 18378 2056 18410
rect 2088 18378 2128 18410
rect 2160 18378 2200 18410
rect 2232 18378 2272 18410
rect 2304 18378 2344 18410
rect 2376 18378 2416 18410
rect 2448 18378 2488 18410
rect 2520 18378 2560 18410
rect 2592 18378 2632 18410
rect 2664 18378 2704 18410
rect 2736 18378 2776 18410
rect 2808 18378 2848 18410
rect 2880 18378 2920 18410
rect 2952 18378 2992 18410
rect 3024 18378 3064 18410
rect 3096 18378 3136 18410
rect 3168 18378 3208 18410
rect 3240 18378 3280 18410
rect 3312 18378 3352 18410
rect 3384 18378 3424 18410
rect 3456 18378 3496 18410
rect 3528 18378 3568 18410
rect 3600 18378 3640 18410
rect 3672 18378 3712 18410
rect 3744 18378 3784 18410
rect 3816 18378 3856 18410
rect 3888 18378 3950 18410
rect 50 18338 3950 18378
rect 50 18306 112 18338
rect 144 18306 184 18338
rect 216 18306 256 18338
rect 288 18306 328 18338
rect 360 18306 400 18338
rect 432 18306 472 18338
rect 504 18306 544 18338
rect 576 18306 616 18338
rect 648 18306 688 18338
rect 720 18306 760 18338
rect 792 18306 832 18338
rect 864 18306 904 18338
rect 936 18306 976 18338
rect 1008 18306 1048 18338
rect 1080 18306 1120 18338
rect 1152 18306 1192 18338
rect 1224 18306 1264 18338
rect 1296 18306 1336 18338
rect 1368 18306 1408 18338
rect 1440 18306 1480 18338
rect 1512 18306 1552 18338
rect 1584 18306 1624 18338
rect 1656 18306 1696 18338
rect 1728 18306 1768 18338
rect 1800 18306 1840 18338
rect 1872 18306 1912 18338
rect 1944 18306 1984 18338
rect 2016 18306 2056 18338
rect 2088 18306 2128 18338
rect 2160 18306 2200 18338
rect 2232 18306 2272 18338
rect 2304 18306 2344 18338
rect 2376 18306 2416 18338
rect 2448 18306 2488 18338
rect 2520 18306 2560 18338
rect 2592 18306 2632 18338
rect 2664 18306 2704 18338
rect 2736 18306 2776 18338
rect 2808 18306 2848 18338
rect 2880 18306 2920 18338
rect 2952 18306 2992 18338
rect 3024 18306 3064 18338
rect 3096 18306 3136 18338
rect 3168 18306 3208 18338
rect 3240 18306 3280 18338
rect 3312 18306 3352 18338
rect 3384 18306 3424 18338
rect 3456 18306 3496 18338
rect 3528 18306 3568 18338
rect 3600 18306 3640 18338
rect 3672 18306 3712 18338
rect 3744 18306 3784 18338
rect 3816 18306 3856 18338
rect 3888 18306 3950 18338
rect 50 18266 3950 18306
rect 50 18234 112 18266
rect 144 18234 184 18266
rect 216 18234 256 18266
rect 288 18234 328 18266
rect 360 18234 400 18266
rect 432 18234 472 18266
rect 504 18234 544 18266
rect 576 18234 616 18266
rect 648 18234 688 18266
rect 720 18234 760 18266
rect 792 18234 832 18266
rect 864 18234 904 18266
rect 936 18234 976 18266
rect 1008 18234 1048 18266
rect 1080 18234 1120 18266
rect 1152 18234 1192 18266
rect 1224 18234 1264 18266
rect 1296 18234 1336 18266
rect 1368 18234 1408 18266
rect 1440 18234 1480 18266
rect 1512 18234 1552 18266
rect 1584 18234 1624 18266
rect 1656 18234 1696 18266
rect 1728 18234 1768 18266
rect 1800 18234 1840 18266
rect 1872 18234 1912 18266
rect 1944 18234 1984 18266
rect 2016 18234 2056 18266
rect 2088 18234 2128 18266
rect 2160 18234 2200 18266
rect 2232 18234 2272 18266
rect 2304 18234 2344 18266
rect 2376 18234 2416 18266
rect 2448 18234 2488 18266
rect 2520 18234 2560 18266
rect 2592 18234 2632 18266
rect 2664 18234 2704 18266
rect 2736 18234 2776 18266
rect 2808 18234 2848 18266
rect 2880 18234 2920 18266
rect 2952 18234 2992 18266
rect 3024 18234 3064 18266
rect 3096 18234 3136 18266
rect 3168 18234 3208 18266
rect 3240 18234 3280 18266
rect 3312 18234 3352 18266
rect 3384 18234 3424 18266
rect 3456 18234 3496 18266
rect 3528 18234 3568 18266
rect 3600 18234 3640 18266
rect 3672 18234 3712 18266
rect 3744 18234 3784 18266
rect 3816 18234 3856 18266
rect 3888 18234 3950 18266
rect 50 18194 3950 18234
rect 50 18162 112 18194
rect 144 18162 184 18194
rect 216 18162 256 18194
rect 288 18162 328 18194
rect 360 18162 400 18194
rect 432 18162 472 18194
rect 504 18162 544 18194
rect 576 18162 616 18194
rect 648 18162 688 18194
rect 720 18162 760 18194
rect 792 18162 832 18194
rect 864 18162 904 18194
rect 936 18162 976 18194
rect 1008 18162 1048 18194
rect 1080 18162 1120 18194
rect 1152 18162 1192 18194
rect 1224 18162 1264 18194
rect 1296 18162 1336 18194
rect 1368 18162 1408 18194
rect 1440 18162 1480 18194
rect 1512 18162 1552 18194
rect 1584 18162 1624 18194
rect 1656 18162 1696 18194
rect 1728 18162 1768 18194
rect 1800 18162 1840 18194
rect 1872 18162 1912 18194
rect 1944 18162 1984 18194
rect 2016 18162 2056 18194
rect 2088 18162 2128 18194
rect 2160 18162 2200 18194
rect 2232 18162 2272 18194
rect 2304 18162 2344 18194
rect 2376 18162 2416 18194
rect 2448 18162 2488 18194
rect 2520 18162 2560 18194
rect 2592 18162 2632 18194
rect 2664 18162 2704 18194
rect 2736 18162 2776 18194
rect 2808 18162 2848 18194
rect 2880 18162 2920 18194
rect 2952 18162 2992 18194
rect 3024 18162 3064 18194
rect 3096 18162 3136 18194
rect 3168 18162 3208 18194
rect 3240 18162 3280 18194
rect 3312 18162 3352 18194
rect 3384 18162 3424 18194
rect 3456 18162 3496 18194
rect 3528 18162 3568 18194
rect 3600 18162 3640 18194
rect 3672 18162 3712 18194
rect 3744 18162 3784 18194
rect 3816 18162 3856 18194
rect 3888 18162 3950 18194
rect 50 18112 3950 18162
rect 50 17848 3950 17912
rect 50 17816 112 17848
rect 144 17816 184 17848
rect 216 17816 256 17848
rect 288 17816 328 17848
rect 360 17816 400 17848
rect 432 17816 472 17848
rect 504 17816 544 17848
rect 576 17816 616 17848
rect 648 17816 688 17848
rect 720 17816 760 17848
rect 792 17816 832 17848
rect 864 17816 904 17848
rect 936 17816 976 17848
rect 1008 17816 1048 17848
rect 1080 17816 1120 17848
rect 1152 17816 1192 17848
rect 1224 17816 1264 17848
rect 1296 17816 1336 17848
rect 1368 17816 1408 17848
rect 1440 17816 1480 17848
rect 1512 17816 1552 17848
rect 1584 17816 1624 17848
rect 1656 17816 1696 17848
rect 1728 17816 1768 17848
rect 1800 17816 1840 17848
rect 1872 17816 1912 17848
rect 1944 17816 1984 17848
rect 2016 17816 2056 17848
rect 2088 17816 2128 17848
rect 2160 17816 2200 17848
rect 2232 17816 2272 17848
rect 2304 17816 2344 17848
rect 2376 17816 2416 17848
rect 2448 17816 2488 17848
rect 2520 17816 2560 17848
rect 2592 17816 2632 17848
rect 2664 17816 2704 17848
rect 2736 17816 2776 17848
rect 2808 17816 2848 17848
rect 2880 17816 2920 17848
rect 2952 17816 2992 17848
rect 3024 17816 3064 17848
rect 3096 17816 3136 17848
rect 3168 17816 3208 17848
rect 3240 17816 3280 17848
rect 3312 17816 3352 17848
rect 3384 17816 3424 17848
rect 3456 17816 3496 17848
rect 3528 17816 3568 17848
rect 3600 17816 3640 17848
rect 3672 17816 3712 17848
rect 3744 17816 3784 17848
rect 3816 17816 3856 17848
rect 3888 17816 3950 17848
rect 50 17776 3950 17816
rect 50 17744 112 17776
rect 144 17744 184 17776
rect 216 17744 256 17776
rect 288 17744 328 17776
rect 360 17744 400 17776
rect 432 17744 472 17776
rect 504 17744 544 17776
rect 576 17744 616 17776
rect 648 17744 688 17776
rect 720 17744 760 17776
rect 792 17744 832 17776
rect 864 17744 904 17776
rect 936 17744 976 17776
rect 1008 17744 1048 17776
rect 1080 17744 1120 17776
rect 1152 17744 1192 17776
rect 1224 17744 1264 17776
rect 1296 17744 1336 17776
rect 1368 17744 1408 17776
rect 1440 17744 1480 17776
rect 1512 17744 1552 17776
rect 1584 17744 1624 17776
rect 1656 17744 1696 17776
rect 1728 17744 1768 17776
rect 1800 17744 1840 17776
rect 1872 17744 1912 17776
rect 1944 17744 1984 17776
rect 2016 17744 2056 17776
rect 2088 17744 2128 17776
rect 2160 17744 2200 17776
rect 2232 17744 2272 17776
rect 2304 17744 2344 17776
rect 2376 17744 2416 17776
rect 2448 17744 2488 17776
rect 2520 17744 2560 17776
rect 2592 17744 2632 17776
rect 2664 17744 2704 17776
rect 2736 17744 2776 17776
rect 2808 17744 2848 17776
rect 2880 17744 2920 17776
rect 2952 17744 2992 17776
rect 3024 17744 3064 17776
rect 3096 17744 3136 17776
rect 3168 17744 3208 17776
rect 3240 17744 3280 17776
rect 3312 17744 3352 17776
rect 3384 17744 3424 17776
rect 3456 17744 3496 17776
rect 3528 17744 3568 17776
rect 3600 17744 3640 17776
rect 3672 17744 3712 17776
rect 3744 17744 3784 17776
rect 3816 17744 3856 17776
rect 3888 17744 3950 17776
rect 50 17704 3950 17744
rect 50 17672 112 17704
rect 144 17672 184 17704
rect 216 17672 256 17704
rect 288 17672 328 17704
rect 360 17672 400 17704
rect 432 17672 472 17704
rect 504 17672 544 17704
rect 576 17672 616 17704
rect 648 17672 688 17704
rect 720 17672 760 17704
rect 792 17672 832 17704
rect 864 17672 904 17704
rect 936 17672 976 17704
rect 1008 17672 1048 17704
rect 1080 17672 1120 17704
rect 1152 17672 1192 17704
rect 1224 17672 1264 17704
rect 1296 17672 1336 17704
rect 1368 17672 1408 17704
rect 1440 17672 1480 17704
rect 1512 17672 1552 17704
rect 1584 17672 1624 17704
rect 1656 17672 1696 17704
rect 1728 17672 1768 17704
rect 1800 17672 1840 17704
rect 1872 17672 1912 17704
rect 1944 17672 1984 17704
rect 2016 17672 2056 17704
rect 2088 17672 2128 17704
rect 2160 17672 2200 17704
rect 2232 17672 2272 17704
rect 2304 17672 2344 17704
rect 2376 17672 2416 17704
rect 2448 17672 2488 17704
rect 2520 17672 2560 17704
rect 2592 17672 2632 17704
rect 2664 17672 2704 17704
rect 2736 17672 2776 17704
rect 2808 17672 2848 17704
rect 2880 17672 2920 17704
rect 2952 17672 2992 17704
rect 3024 17672 3064 17704
rect 3096 17672 3136 17704
rect 3168 17672 3208 17704
rect 3240 17672 3280 17704
rect 3312 17672 3352 17704
rect 3384 17672 3424 17704
rect 3456 17672 3496 17704
rect 3528 17672 3568 17704
rect 3600 17672 3640 17704
rect 3672 17672 3712 17704
rect 3744 17672 3784 17704
rect 3816 17672 3856 17704
rect 3888 17672 3950 17704
rect 50 17632 3950 17672
rect 50 17600 112 17632
rect 144 17600 184 17632
rect 216 17600 256 17632
rect 288 17600 328 17632
rect 360 17600 400 17632
rect 432 17600 472 17632
rect 504 17600 544 17632
rect 576 17600 616 17632
rect 648 17600 688 17632
rect 720 17600 760 17632
rect 792 17600 832 17632
rect 864 17600 904 17632
rect 936 17600 976 17632
rect 1008 17600 1048 17632
rect 1080 17600 1120 17632
rect 1152 17600 1192 17632
rect 1224 17600 1264 17632
rect 1296 17600 1336 17632
rect 1368 17600 1408 17632
rect 1440 17600 1480 17632
rect 1512 17600 1552 17632
rect 1584 17600 1624 17632
rect 1656 17600 1696 17632
rect 1728 17600 1768 17632
rect 1800 17600 1840 17632
rect 1872 17600 1912 17632
rect 1944 17600 1984 17632
rect 2016 17600 2056 17632
rect 2088 17600 2128 17632
rect 2160 17600 2200 17632
rect 2232 17600 2272 17632
rect 2304 17600 2344 17632
rect 2376 17600 2416 17632
rect 2448 17600 2488 17632
rect 2520 17600 2560 17632
rect 2592 17600 2632 17632
rect 2664 17600 2704 17632
rect 2736 17600 2776 17632
rect 2808 17600 2848 17632
rect 2880 17600 2920 17632
rect 2952 17600 2992 17632
rect 3024 17600 3064 17632
rect 3096 17600 3136 17632
rect 3168 17600 3208 17632
rect 3240 17600 3280 17632
rect 3312 17600 3352 17632
rect 3384 17600 3424 17632
rect 3456 17600 3496 17632
rect 3528 17600 3568 17632
rect 3600 17600 3640 17632
rect 3672 17600 3712 17632
rect 3744 17600 3784 17632
rect 3816 17600 3856 17632
rect 3888 17600 3950 17632
rect 50 17560 3950 17600
rect 50 17528 112 17560
rect 144 17528 184 17560
rect 216 17528 256 17560
rect 288 17528 328 17560
rect 360 17528 400 17560
rect 432 17528 472 17560
rect 504 17528 544 17560
rect 576 17528 616 17560
rect 648 17528 688 17560
rect 720 17528 760 17560
rect 792 17528 832 17560
rect 864 17528 904 17560
rect 936 17528 976 17560
rect 1008 17528 1048 17560
rect 1080 17528 1120 17560
rect 1152 17528 1192 17560
rect 1224 17528 1264 17560
rect 1296 17528 1336 17560
rect 1368 17528 1408 17560
rect 1440 17528 1480 17560
rect 1512 17528 1552 17560
rect 1584 17528 1624 17560
rect 1656 17528 1696 17560
rect 1728 17528 1768 17560
rect 1800 17528 1840 17560
rect 1872 17528 1912 17560
rect 1944 17528 1984 17560
rect 2016 17528 2056 17560
rect 2088 17528 2128 17560
rect 2160 17528 2200 17560
rect 2232 17528 2272 17560
rect 2304 17528 2344 17560
rect 2376 17528 2416 17560
rect 2448 17528 2488 17560
rect 2520 17528 2560 17560
rect 2592 17528 2632 17560
rect 2664 17528 2704 17560
rect 2736 17528 2776 17560
rect 2808 17528 2848 17560
rect 2880 17528 2920 17560
rect 2952 17528 2992 17560
rect 3024 17528 3064 17560
rect 3096 17528 3136 17560
rect 3168 17528 3208 17560
rect 3240 17528 3280 17560
rect 3312 17528 3352 17560
rect 3384 17528 3424 17560
rect 3456 17528 3496 17560
rect 3528 17528 3568 17560
rect 3600 17528 3640 17560
rect 3672 17528 3712 17560
rect 3744 17528 3784 17560
rect 3816 17528 3856 17560
rect 3888 17528 3950 17560
rect 50 17488 3950 17528
rect 50 17456 112 17488
rect 144 17456 184 17488
rect 216 17456 256 17488
rect 288 17456 328 17488
rect 360 17456 400 17488
rect 432 17456 472 17488
rect 504 17456 544 17488
rect 576 17456 616 17488
rect 648 17456 688 17488
rect 720 17456 760 17488
rect 792 17456 832 17488
rect 864 17456 904 17488
rect 936 17456 976 17488
rect 1008 17456 1048 17488
rect 1080 17456 1120 17488
rect 1152 17456 1192 17488
rect 1224 17456 1264 17488
rect 1296 17456 1336 17488
rect 1368 17456 1408 17488
rect 1440 17456 1480 17488
rect 1512 17456 1552 17488
rect 1584 17456 1624 17488
rect 1656 17456 1696 17488
rect 1728 17456 1768 17488
rect 1800 17456 1840 17488
rect 1872 17456 1912 17488
rect 1944 17456 1984 17488
rect 2016 17456 2056 17488
rect 2088 17456 2128 17488
rect 2160 17456 2200 17488
rect 2232 17456 2272 17488
rect 2304 17456 2344 17488
rect 2376 17456 2416 17488
rect 2448 17456 2488 17488
rect 2520 17456 2560 17488
rect 2592 17456 2632 17488
rect 2664 17456 2704 17488
rect 2736 17456 2776 17488
rect 2808 17456 2848 17488
rect 2880 17456 2920 17488
rect 2952 17456 2992 17488
rect 3024 17456 3064 17488
rect 3096 17456 3136 17488
rect 3168 17456 3208 17488
rect 3240 17456 3280 17488
rect 3312 17456 3352 17488
rect 3384 17456 3424 17488
rect 3456 17456 3496 17488
rect 3528 17456 3568 17488
rect 3600 17456 3640 17488
rect 3672 17456 3712 17488
rect 3744 17456 3784 17488
rect 3816 17456 3856 17488
rect 3888 17456 3950 17488
rect 50 17416 3950 17456
rect 50 17384 112 17416
rect 144 17384 184 17416
rect 216 17384 256 17416
rect 288 17384 328 17416
rect 360 17384 400 17416
rect 432 17384 472 17416
rect 504 17384 544 17416
rect 576 17384 616 17416
rect 648 17384 688 17416
rect 720 17384 760 17416
rect 792 17384 832 17416
rect 864 17384 904 17416
rect 936 17384 976 17416
rect 1008 17384 1048 17416
rect 1080 17384 1120 17416
rect 1152 17384 1192 17416
rect 1224 17384 1264 17416
rect 1296 17384 1336 17416
rect 1368 17384 1408 17416
rect 1440 17384 1480 17416
rect 1512 17384 1552 17416
rect 1584 17384 1624 17416
rect 1656 17384 1696 17416
rect 1728 17384 1768 17416
rect 1800 17384 1840 17416
rect 1872 17384 1912 17416
rect 1944 17384 1984 17416
rect 2016 17384 2056 17416
rect 2088 17384 2128 17416
rect 2160 17384 2200 17416
rect 2232 17384 2272 17416
rect 2304 17384 2344 17416
rect 2376 17384 2416 17416
rect 2448 17384 2488 17416
rect 2520 17384 2560 17416
rect 2592 17384 2632 17416
rect 2664 17384 2704 17416
rect 2736 17384 2776 17416
rect 2808 17384 2848 17416
rect 2880 17384 2920 17416
rect 2952 17384 2992 17416
rect 3024 17384 3064 17416
rect 3096 17384 3136 17416
rect 3168 17384 3208 17416
rect 3240 17384 3280 17416
rect 3312 17384 3352 17416
rect 3384 17384 3424 17416
rect 3456 17384 3496 17416
rect 3528 17384 3568 17416
rect 3600 17384 3640 17416
rect 3672 17384 3712 17416
rect 3744 17384 3784 17416
rect 3816 17384 3856 17416
rect 3888 17384 3950 17416
rect 50 17344 3950 17384
rect 50 17312 112 17344
rect 144 17312 184 17344
rect 216 17312 256 17344
rect 288 17312 328 17344
rect 360 17312 400 17344
rect 432 17312 472 17344
rect 504 17312 544 17344
rect 576 17312 616 17344
rect 648 17312 688 17344
rect 720 17312 760 17344
rect 792 17312 832 17344
rect 864 17312 904 17344
rect 936 17312 976 17344
rect 1008 17312 1048 17344
rect 1080 17312 1120 17344
rect 1152 17312 1192 17344
rect 1224 17312 1264 17344
rect 1296 17312 1336 17344
rect 1368 17312 1408 17344
rect 1440 17312 1480 17344
rect 1512 17312 1552 17344
rect 1584 17312 1624 17344
rect 1656 17312 1696 17344
rect 1728 17312 1768 17344
rect 1800 17312 1840 17344
rect 1872 17312 1912 17344
rect 1944 17312 1984 17344
rect 2016 17312 2056 17344
rect 2088 17312 2128 17344
rect 2160 17312 2200 17344
rect 2232 17312 2272 17344
rect 2304 17312 2344 17344
rect 2376 17312 2416 17344
rect 2448 17312 2488 17344
rect 2520 17312 2560 17344
rect 2592 17312 2632 17344
rect 2664 17312 2704 17344
rect 2736 17312 2776 17344
rect 2808 17312 2848 17344
rect 2880 17312 2920 17344
rect 2952 17312 2992 17344
rect 3024 17312 3064 17344
rect 3096 17312 3136 17344
rect 3168 17312 3208 17344
rect 3240 17312 3280 17344
rect 3312 17312 3352 17344
rect 3384 17312 3424 17344
rect 3456 17312 3496 17344
rect 3528 17312 3568 17344
rect 3600 17312 3640 17344
rect 3672 17312 3712 17344
rect 3744 17312 3784 17344
rect 3816 17312 3856 17344
rect 3888 17312 3950 17344
rect 50 17272 3950 17312
rect 50 17240 112 17272
rect 144 17240 184 17272
rect 216 17240 256 17272
rect 288 17240 328 17272
rect 360 17240 400 17272
rect 432 17240 472 17272
rect 504 17240 544 17272
rect 576 17240 616 17272
rect 648 17240 688 17272
rect 720 17240 760 17272
rect 792 17240 832 17272
rect 864 17240 904 17272
rect 936 17240 976 17272
rect 1008 17240 1048 17272
rect 1080 17240 1120 17272
rect 1152 17240 1192 17272
rect 1224 17240 1264 17272
rect 1296 17240 1336 17272
rect 1368 17240 1408 17272
rect 1440 17240 1480 17272
rect 1512 17240 1552 17272
rect 1584 17240 1624 17272
rect 1656 17240 1696 17272
rect 1728 17240 1768 17272
rect 1800 17240 1840 17272
rect 1872 17240 1912 17272
rect 1944 17240 1984 17272
rect 2016 17240 2056 17272
rect 2088 17240 2128 17272
rect 2160 17240 2200 17272
rect 2232 17240 2272 17272
rect 2304 17240 2344 17272
rect 2376 17240 2416 17272
rect 2448 17240 2488 17272
rect 2520 17240 2560 17272
rect 2592 17240 2632 17272
rect 2664 17240 2704 17272
rect 2736 17240 2776 17272
rect 2808 17240 2848 17272
rect 2880 17240 2920 17272
rect 2952 17240 2992 17272
rect 3024 17240 3064 17272
rect 3096 17240 3136 17272
rect 3168 17240 3208 17272
rect 3240 17240 3280 17272
rect 3312 17240 3352 17272
rect 3384 17240 3424 17272
rect 3456 17240 3496 17272
rect 3528 17240 3568 17272
rect 3600 17240 3640 17272
rect 3672 17240 3712 17272
rect 3744 17240 3784 17272
rect 3816 17240 3856 17272
rect 3888 17240 3950 17272
rect 50 17200 3950 17240
rect 50 17168 112 17200
rect 144 17168 184 17200
rect 216 17168 256 17200
rect 288 17168 328 17200
rect 360 17168 400 17200
rect 432 17168 472 17200
rect 504 17168 544 17200
rect 576 17168 616 17200
rect 648 17168 688 17200
rect 720 17168 760 17200
rect 792 17168 832 17200
rect 864 17168 904 17200
rect 936 17168 976 17200
rect 1008 17168 1048 17200
rect 1080 17168 1120 17200
rect 1152 17168 1192 17200
rect 1224 17168 1264 17200
rect 1296 17168 1336 17200
rect 1368 17168 1408 17200
rect 1440 17168 1480 17200
rect 1512 17168 1552 17200
rect 1584 17168 1624 17200
rect 1656 17168 1696 17200
rect 1728 17168 1768 17200
rect 1800 17168 1840 17200
rect 1872 17168 1912 17200
rect 1944 17168 1984 17200
rect 2016 17168 2056 17200
rect 2088 17168 2128 17200
rect 2160 17168 2200 17200
rect 2232 17168 2272 17200
rect 2304 17168 2344 17200
rect 2376 17168 2416 17200
rect 2448 17168 2488 17200
rect 2520 17168 2560 17200
rect 2592 17168 2632 17200
rect 2664 17168 2704 17200
rect 2736 17168 2776 17200
rect 2808 17168 2848 17200
rect 2880 17168 2920 17200
rect 2952 17168 2992 17200
rect 3024 17168 3064 17200
rect 3096 17168 3136 17200
rect 3168 17168 3208 17200
rect 3240 17168 3280 17200
rect 3312 17168 3352 17200
rect 3384 17168 3424 17200
rect 3456 17168 3496 17200
rect 3528 17168 3568 17200
rect 3600 17168 3640 17200
rect 3672 17168 3712 17200
rect 3744 17168 3784 17200
rect 3816 17168 3856 17200
rect 3888 17168 3950 17200
rect 50 17128 3950 17168
rect 50 17096 112 17128
rect 144 17096 184 17128
rect 216 17096 256 17128
rect 288 17096 328 17128
rect 360 17096 400 17128
rect 432 17096 472 17128
rect 504 17096 544 17128
rect 576 17096 616 17128
rect 648 17096 688 17128
rect 720 17096 760 17128
rect 792 17096 832 17128
rect 864 17096 904 17128
rect 936 17096 976 17128
rect 1008 17096 1048 17128
rect 1080 17096 1120 17128
rect 1152 17096 1192 17128
rect 1224 17096 1264 17128
rect 1296 17096 1336 17128
rect 1368 17096 1408 17128
rect 1440 17096 1480 17128
rect 1512 17096 1552 17128
rect 1584 17096 1624 17128
rect 1656 17096 1696 17128
rect 1728 17096 1768 17128
rect 1800 17096 1840 17128
rect 1872 17096 1912 17128
rect 1944 17096 1984 17128
rect 2016 17096 2056 17128
rect 2088 17096 2128 17128
rect 2160 17096 2200 17128
rect 2232 17096 2272 17128
rect 2304 17096 2344 17128
rect 2376 17096 2416 17128
rect 2448 17096 2488 17128
rect 2520 17096 2560 17128
rect 2592 17096 2632 17128
rect 2664 17096 2704 17128
rect 2736 17096 2776 17128
rect 2808 17096 2848 17128
rect 2880 17096 2920 17128
rect 2952 17096 2992 17128
rect 3024 17096 3064 17128
rect 3096 17096 3136 17128
rect 3168 17096 3208 17128
rect 3240 17096 3280 17128
rect 3312 17096 3352 17128
rect 3384 17096 3424 17128
rect 3456 17096 3496 17128
rect 3528 17096 3568 17128
rect 3600 17096 3640 17128
rect 3672 17096 3712 17128
rect 3744 17096 3784 17128
rect 3816 17096 3856 17128
rect 3888 17096 3950 17128
rect 50 17056 3950 17096
rect 50 17024 112 17056
rect 144 17024 184 17056
rect 216 17024 256 17056
rect 288 17024 328 17056
rect 360 17024 400 17056
rect 432 17024 472 17056
rect 504 17024 544 17056
rect 576 17024 616 17056
rect 648 17024 688 17056
rect 720 17024 760 17056
rect 792 17024 832 17056
rect 864 17024 904 17056
rect 936 17024 976 17056
rect 1008 17024 1048 17056
rect 1080 17024 1120 17056
rect 1152 17024 1192 17056
rect 1224 17024 1264 17056
rect 1296 17024 1336 17056
rect 1368 17024 1408 17056
rect 1440 17024 1480 17056
rect 1512 17024 1552 17056
rect 1584 17024 1624 17056
rect 1656 17024 1696 17056
rect 1728 17024 1768 17056
rect 1800 17024 1840 17056
rect 1872 17024 1912 17056
rect 1944 17024 1984 17056
rect 2016 17024 2056 17056
rect 2088 17024 2128 17056
rect 2160 17024 2200 17056
rect 2232 17024 2272 17056
rect 2304 17024 2344 17056
rect 2376 17024 2416 17056
rect 2448 17024 2488 17056
rect 2520 17024 2560 17056
rect 2592 17024 2632 17056
rect 2664 17024 2704 17056
rect 2736 17024 2776 17056
rect 2808 17024 2848 17056
rect 2880 17024 2920 17056
rect 2952 17024 2992 17056
rect 3024 17024 3064 17056
rect 3096 17024 3136 17056
rect 3168 17024 3208 17056
rect 3240 17024 3280 17056
rect 3312 17024 3352 17056
rect 3384 17024 3424 17056
rect 3456 17024 3496 17056
rect 3528 17024 3568 17056
rect 3600 17024 3640 17056
rect 3672 17024 3712 17056
rect 3744 17024 3784 17056
rect 3816 17024 3856 17056
rect 3888 17024 3950 17056
rect 50 16984 3950 17024
rect 50 16952 112 16984
rect 144 16952 184 16984
rect 216 16952 256 16984
rect 288 16952 328 16984
rect 360 16952 400 16984
rect 432 16952 472 16984
rect 504 16952 544 16984
rect 576 16952 616 16984
rect 648 16952 688 16984
rect 720 16952 760 16984
rect 792 16952 832 16984
rect 864 16952 904 16984
rect 936 16952 976 16984
rect 1008 16952 1048 16984
rect 1080 16952 1120 16984
rect 1152 16952 1192 16984
rect 1224 16952 1264 16984
rect 1296 16952 1336 16984
rect 1368 16952 1408 16984
rect 1440 16952 1480 16984
rect 1512 16952 1552 16984
rect 1584 16952 1624 16984
rect 1656 16952 1696 16984
rect 1728 16952 1768 16984
rect 1800 16952 1840 16984
rect 1872 16952 1912 16984
rect 1944 16952 1984 16984
rect 2016 16952 2056 16984
rect 2088 16952 2128 16984
rect 2160 16952 2200 16984
rect 2232 16952 2272 16984
rect 2304 16952 2344 16984
rect 2376 16952 2416 16984
rect 2448 16952 2488 16984
rect 2520 16952 2560 16984
rect 2592 16952 2632 16984
rect 2664 16952 2704 16984
rect 2736 16952 2776 16984
rect 2808 16952 2848 16984
rect 2880 16952 2920 16984
rect 2952 16952 2992 16984
rect 3024 16952 3064 16984
rect 3096 16952 3136 16984
rect 3168 16952 3208 16984
rect 3240 16952 3280 16984
rect 3312 16952 3352 16984
rect 3384 16952 3424 16984
rect 3456 16952 3496 16984
rect 3528 16952 3568 16984
rect 3600 16952 3640 16984
rect 3672 16952 3712 16984
rect 3744 16952 3784 16984
rect 3816 16952 3856 16984
rect 3888 16952 3950 16984
rect 50 16912 3950 16952
rect 50 16880 112 16912
rect 144 16880 184 16912
rect 216 16880 256 16912
rect 288 16880 328 16912
rect 360 16880 400 16912
rect 432 16880 472 16912
rect 504 16880 544 16912
rect 576 16880 616 16912
rect 648 16880 688 16912
rect 720 16880 760 16912
rect 792 16880 832 16912
rect 864 16880 904 16912
rect 936 16880 976 16912
rect 1008 16880 1048 16912
rect 1080 16880 1120 16912
rect 1152 16880 1192 16912
rect 1224 16880 1264 16912
rect 1296 16880 1336 16912
rect 1368 16880 1408 16912
rect 1440 16880 1480 16912
rect 1512 16880 1552 16912
rect 1584 16880 1624 16912
rect 1656 16880 1696 16912
rect 1728 16880 1768 16912
rect 1800 16880 1840 16912
rect 1872 16880 1912 16912
rect 1944 16880 1984 16912
rect 2016 16880 2056 16912
rect 2088 16880 2128 16912
rect 2160 16880 2200 16912
rect 2232 16880 2272 16912
rect 2304 16880 2344 16912
rect 2376 16880 2416 16912
rect 2448 16880 2488 16912
rect 2520 16880 2560 16912
rect 2592 16880 2632 16912
rect 2664 16880 2704 16912
rect 2736 16880 2776 16912
rect 2808 16880 2848 16912
rect 2880 16880 2920 16912
rect 2952 16880 2992 16912
rect 3024 16880 3064 16912
rect 3096 16880 3136 16912
rect 3168 16880 3208 16912
rect 3240 16880 3280 16912
rect 3312 16880 3352 16912
rect 3384 16880 3424 16912
rect 3456 16880 3496 16912
rect 3528 16880 3568 16912
rect 3600 16880 3640 16912
rect 3672 16880 3712 16912
rect 3744 16880 3784 16912
rect 3816 16880 3856 16912
rect 3888 16880 3950 16912
rect 50 16840 3950 16880
rect 50 16808 112 16840
rect 144 16808 184 16840
rect 216 16808 256 16840
rect 288 16808 328 16840
rect 360 16808 400 16840
rect 432 16808 472 16840
rect 504 16808 544 16840
rect 576 16808 616 16840
rect 648 16808 688 16840
rect 720 16808 760 16840
rect 792 16808 832 16840
rect 864 16808 904 16840
rect 936 16808 976 16840
rect 1008 16808 1048 16840
rect 1080 16808 1120 16840
rect 1152 16808 1192 16840
rect 1224 16808 1264 16840
rect 1296 16808 1336 16840
rect 1368 16808 1408 16840
rect 1440 16808 1480 16840
rect 1512 16808 1552 16840
rect 1584 16808 1624 16840
rect 1656 16808 1696 16840
rect 1728 16808 1768 16840
rect 1800 16808 1840 16840
rect 1872 16808 1912 16840
rect 1944 16808 1984 16840
rect 2016 16808 2056 16840
rect 2088 16808 2128 16840
rect 2160 16808 2200 16840
rect 2232 16808 2272 16840
rect 2304 16808 2344 16840
rect 2376 16808 2416 16840
rect 2448 16808 2488 16840
rect 2520 16808 2560 16840
rect 2592 16808 2632 16840
rect 2664 16808 2704 16840
rect 2736 16808 2776 16840
rect 2808 16808 2848 16840
rect 2880 16808 2920 16840
rect 2952 16808 2992 16840
rect 3024 16808 3064 16840
rect 3096 16808 3136 16840
rect 3168 16808 3208 16840
rect 3240 16808 3280 16840
rect 3312 16808 3352 16840
rect 3384 16808 3424 16840
rect 3456 16808 3496 16840
rect 3528 16808 3568 16840
rect 3600 16808 3640 16840
rect 3672 16808 3712 16840
rect 3744 16808 3784 16840
rect 3816 16808 3856 16840
rect 3888 16808 3950 16840
rect 50 16768 3950 16808
rect 50 16736 112 16768
rect 144 16736 184 16768
rect 216 16736 256 16768
rect 288 16736 328 16768
rect 360 16736 400 16768
rect 432 16736 472 16768
rect 504 16736 544 16768
rect 576 16736 616 16768
rect 648 16736 688 16768
rect 720 16736 760 16768
rect 792 16736 832 16768
rect 864 16736 904 16768
rect 936 16736 976 16768
rect 1008 16736 1048 16768
rect 1080 16736 1120 16768
rect 1152 16736 1192 16768
rect 1224 16736 1264 16768
rect 1296 16736 1336 16768
rect 1368 16736 1408 16768
rect 1440 16736 1480 16768
rect 1512 16736 1552 16768
rect 1584 16736 1624 16768
rect 1656 16736 1696 16768
rect 1728 16736 1768 16768
rect 1800 16736 1840 16768
rect 1872 16736 1912 16768
rect 1944 16736 1984 16768
rect 2016 16736 2056 16768
rect 2088 16736 2128 16768
rect 2160 16736 2200 16768
rect 2232 16736 2272 16768
rect 2304 16736 2344 16768
rect 2376 16736 2416 16768
rect 2448 16736 2488 16768
rect 2520 16736 2560 16768
rect 2592 16736 2632 16768
rect 2664 16736 2704 16768
rect 2736 16736 2776 16768
rect 2808 16736 2848 16768
rect 2880 16736 2920 16768
rect 2952 16736 2992 16768
rect 3024 16736 3064 16768
rect 3096 16736 3136 16768
rect 3168 16736 3208 16768
rect 3240 16736 3280 16768
rect 3312 16736 3352 16768
rect 3384 16736 3424 16768
rect 3456 16736 3496 16768
rect 3528 16736 3568 16768
rect 3600 16736 3640 16768
rect 3672 16736 3712 16768
rect 3744 16736 3784 16768
rect 3816 16736 3856 16768
rect 3888 16736 3950 16768
rect 50 16696 3950 16736
rect 50 16664 112 16696
rect 144 16664 184 16696
rect 216 16664 256 16696
rect 288 16664 328 16696
rect 360 16664 400 16696
rect 432 16664 472 16696
rect 504 16664 544 16696
rect 576 16664 616 16696
rect 648 16664 688 16696
rect 720 16664 760 16696
rect 792 16664 832 16696
rect 864 16664 904 16696
rect 936 16664 976 16696
rect 1008 16664 1048 16696
rect 1080 16664 1120 16696
rect 1152 16664 1192 16696
rect 1224 16664 1264 16696
rect 1296 16664 1336 16696
rect 1368 16664 1408 16696
rect 1440 16664 1480 16696
rect 1512 16664 1552 16696
rect 1584 16664 1624 16696
rect 1656 16664 1696 16696
rect 1728 16664 1768 16696
rect 1800 16664 1840 16696
rect 1872 16664 1912 16696
rect 1944 16664 1984 16696
rect 2016 16664 2056 16696
rect 2088 16664 2128 16696
rect 2160 16664 2200 16696
rect 2232 16664 2272 16696
rect 2304 16664 2344 16696
rect 2376 16664 2416 16696
rect 2448 16664 2488 16696
rect 2520 16664 2560 16696
rect 2592 16664 2632 16696
rect 2664 16664 2704 16696
rect 2736 16664 2776 16696
rect 2808 16664 2848 16696
rect 2880 16664 2920 16696
rect 2952 16664 2992 16696
rect 3024 16664 3064 16696
rect 3096 16664 3136 16696
rect 3168 16664 3208 16696
rect 3240 16664 3280 16696
rect 3312 16664 3352 16696
rect 3384 16664 3424 16696
rect 3456 16664 3496 16696
rect 3528 16664 3568 16696
rect 3600 16664 3640 16696
rect 3672 16664 3712 16696
rect 3744 16664 3784 16696
rect 3816 16664 3856 16696
rect 3888 16664 3950 16696
rect 50 16624 3950 16664
rect 50 16592 112 16624
rect 144 16592 184 16624
rect 216 16592 256 16624
rect 288 16592 328 16624
rect 360 16592 400 16624
rect 432 16592 472 16624
rect 504 16592 544 16624
rect 576 16592 616 16624
rect 648 16592 688 16624
rect 720 16592 760 16624
rect 792 16592 832 16624
rect 864 16592 904 16624
rect 936 16592 976 16624
rect 1008 16592 1048 16624
rect 1080 16592 1120 16624
rect 1152 16592 1192 16624
rect 1224 16592 1264 16624
rect 1296 16592 1336 16624
rect 1368 16592 1408 16624
rect 1440 16592 1480 16624
rect 1512 16592 1552 16624
rect 1584 16592 1624 16624
rect 1656 16592 1696 16624
rect 1728 16592 1768 16624
rect 1800 16592 1840 16624
rect 1872 16592 1912 16624
rect 1944 16592 1984 16624
rect 2016 16592 2056 16624
rect 2088 16592 2128 16624
rect 2160 16592 2200 16624
rect 2232 16592 2272 16624
rect 2304 16592 2344 16624
rect 2376 16592 2416 16624
rect 2448 16592 2488 16624
rect 2520 16592 2560 16624
rect 2592 16592 2632 16624
rect 2664 16592 2704 16624
rect 2736 16592 2776 16624
rect 2808 16592 2848 16624
rect 2880 16592 2920 16624
rect 2952 16592 2992 16624
rect 3024 16592 3064 16624
rect 3096 16592 3136 16624
rect 3168 16592 3208 16624
rect 3240 16592 3280 16624
rect 3312 16592 3352 16624
rect 3384 16592 3424 16624
rect 3456 16592 3496 16624
rect 3528 16592 3568 16624
rect 3600 16592 3640 16624
rect 3672 16592 3712 16624
rect 3744 16592 3784 16624
rect 3816 16592 3856 16624
rect 3888 16592 3950 16624
rect 50 16552 3950 16592
rect 50 16520 112 16552
rect 144 16520 184 16552
rect 216 16520 256 16552
rect 288 16520 328 16552
rect 360 16520 400 16552
rect 432 16520 472 16552
rect 504 16520 544 16552
rect 576 16520 616 16552
rect 648 16520 688 16552
rect 720 16520 760 16552
rect 792 16520 832 16552
rect 864 16520 904 16552
rect 936 16520 976 16552
rect 1008 16520 1048 16552
rect 1080 16520 1120 16552
rect 1152 16520 1192 16552
rect 1224 16520 1264 16552
rect 1296 16520 1336 16552
rect 1368 16520 1408 16552
rect 1440 16520 1480 16552
rect 1512 16520 1552 16552
rect 1584 16520 1624 16552
rect 1656 16520 1696 16552
rect 1728 16520 1768 16552
rect 1800 16520 1840 16552
rect 1872 16520 1912 16552
rect 1944 16520 1984 16552
rect 2016 16520 2056 16552
rect 2088 16520 2128 16552
rect 2160 16520 2200 16552
rect 2232 16520 2272 16552
rect 2304 16520 2344 16552
rect 2376 16520 2416 16552
rect 2448 16520 2488 16552
rect 2520 16520 2560 16552
rect 2592 16520 2632 16552
rect 2664 16520 2704 16552
rect 2736 16520 2776 16552
rect 2808 16520 2848 16552
rect 2880 16520 2920 16552
rect 2952 16520 2992 16552
rect 3024 16520 3064 16552
rect 3096 16520 3136 16552
rect 3168 16520 3208 16552
rect 3240 16520 3280 16552
rect 3312 16520 3352 16552
rect 3384 16520 3424 16552
rect 3456 16520 3496 16552
rect 3528 16520 3568 16552
rect 3600 16520 3640 16552
rect 3672 16520 3712 16552
rect 3744 16520 3784 16552
rect 3816 16520 3856 16552
rect 3888 16520 3950 16552
rect 50 16480 3950 16520
rect 50 16448 112 16480
rect 144 16448 184 16480
rect 216 16448 256 16480
rect 288 16448 328 16480
rect 360 16448 400 16480
rect 432 16448 472 16480
rect 504 16448 544 16480
rect 576 16448 616 16480
rect 648 16448 688 16480
rect 720 16448 760 16480
rect 792 16448 832 16480
rect 864 16448 904 16480
rect 936 16448 976 16480
rect 1008 16448 1048 16480
rect 1080 16448 1120 16480
rect 1152 16448 1192 16480
rect 1224 16448 1264 16480
rect 1296 16448 1336 16480
rect 1368 16448 1408 16480
rect 1440 16448 1480 16480
rect 1512 16448 1552 16480
rect 1584 16448 1624 16480
rect 1656 16448 1696 16480
rect 1728 16448 1768 16480
rect 1800 16448 1840 16480
rect 1872 16448 1912 16480
rect 1944 16448 1984 16480
rect 2016 16448 2056 16480
rect 2088 16448 2128 16480
rect 2160 16448 2200 16480
rect 2232 16448 2272 16480
rect 2304 16448 2344 16480
rect 2376 16448 2416 16480
rect 2448 16448 2488 16480
rect 2520 16448 2560 16480
rect 2592 16448 2632 16480
rect 2664 16448 2704 16480
rect 2736 16448 2776 16480
rect 2808 16448 2848 16480
rect 2880 16448 2920 16480
rect 2952 16448 2992 16480
rect 3024 16448 3064 16480
rect 3096 16448 3136 16480
rect 3168 16448 3208 16480
rect 3240 16448 3280 16480
rect 3312 16448 3352 16480
rect 3384 16448 3424 16480
rect 3456 16448 3496 16480
rect 3528 16448 3568 16480
rect 3600 16448 3640 16480
rect 3672 16448 3712 16480
rect 3744 16448 3784 16480
rect 3816 16448 3856 16480
rect 3888 16448 3950 16480
rect 50 16408 3950 16448
rect 50 16376 112 16408
rect 144 16376 184 16408
rect 216 16376 256 16408
rect 288 16376 328 16408
rect 360 16376 400 16408
rect 432 16376 472 16408
rect 504 16376 544 16408
rect 576 16376 616 16408
rect 648 16376 688 16408
rect 720 16376 760 16408
rect 792 16376 832 16408
rect 864 16376 904 16408
rect 936 16376 976 16408
rect 1008 16376 1048 16408
rect 1080 16376 1120 16408
rect 1152 16376 1192 16408
rect 1224 16376 1264 16408
rect 1296 16376 1336 16408
rect 1368 16376 1408 16408
rect 1440 16376 1480 16408
rect 1512 16376 1552 16408
rect 1584 16376 1624 16408
rect 1656 16376 1696 16408
rect 1728 16376 1768 16408
rect 1800 16376 1840 16408
rect 1872 16376 1912 16408
rect 1944 16376 1984 16408
rect 2016 16376 2056 16408
rect 2088 16376 2128 16408
rect 2160 16376 2200 16408
rect 2232 16376 2272 16408
rect 2304 16376 2344 16408
rect 2376 16376 2416 16408
rect 2448 16376 2488 16408
rect 2520 16376 2560 16408
rect 2592 16376 2632 16408
rect 2664 16376 2704 16408
rect 2736 16376 2776 16408
rect 2808 16376 2848 16408
rect 2880 16376 2920 16408
rect 2952 16376 2992 16408
rect 3024 16376 3064 16408
rect 3096 16376 3136 16408
rect 3168 16376 3208 16408
rect 3240 16376 3280 16408
rect 3312 16376 3352 16408
rect 3384 16376 3424 16408
rect 3456 16376 3496 16408
rect 3528 16376 3568 16408
rect 3600 16376 3640 16408
rect 3672 16376 3712 16408
rect 3744 16376 3784 16408
rect 3816 16376 3856 16408
rect 3888 16376 3950 16408
rect 50 16336 3950 16376
rect 50 16304 112 16336
rect 144 16304 184 16336
rect 216 16304 256 16336
rect 288 16304 328 16336
rect 360 16304 400 16336
rect 432 16304 472 16336
rect 504 16304 544 16336
rect 576 16304 616 16336
rect 648 16304 688 16336
rect 720 16304 760 16336
rect 792 16304 832 16336
rect 864 16304 904 16336
rect 936 16304 976 16336
rect 1008 16304 1048 16336
rect 1080 16304 1120 16336
rect 1152 16304 1192 16336
rect 1224 16304 1264 16336
rect 1296 16304 1336 16336
rect 1368 16304 1408 16336
rect 1440 16304 1480 16336
rect 1512 16304 1552 16336
rect 1584 16304 1624 16336
rect 1656 16304 1696 16336
rect 1728 16304 1768 16336
rect 1800 16304 1840 16336
rect 1872 16304 1912 16336
rect 1944 16304 1984 16336
rect 2016 16304 2056 16336
rect 2088 16304 2128 16336
rect 2160 16304 2200 16336
rect 2232 16304 2272 16336
rect 2304 16304 2344 16336
rect 2376 16304 2416 16336
rect 2448 16304 2488 16336
rect 2520 16304 2560 16336
rect 2592 16304 2632 16336
rect 2664 16304 2704 16336
rect 2736 16304 2776 16336
rect 2808 16304 2848 16336
rect 2880 16304 2920 16336
rect 2952 16304 2992 16336
rect 3024 16304 3064 16336
rect 3096 16304 3136 16336
rect 3168 16304 3208 16336
rect 3240 16304 3280 16336
rect 3312 16304 3352 16336
rect 3384 16304 3424 16336
rect 3456 16304 3496 16336
rect 3528 16304 3568 16336
rect 3600 16304 3640 16336
rect 3672 16304 3712 16336
rect 3744 16304 3784 16336
rect 3816 16304 3856 16336
rect 3888 16304 3950 16336
rect 50 16264 3950 16304
rect 50 16232 112 16264
rect 144 16232 184 16264
rect 216 16232 256 16264
rect 288 16232 328 16264
rect 360 16232 400 16264
rect 432 16232 472 16264
rect 504 16232 544 16264
rect 576 16232 616 16264
rect 648 16232 688 16264
rect 720 16232 760 16264
rect 792 16232 832 16264
rect 864 16232 904 16264
rect 936 16232 976 16264
rect 1008 16232 1048 16264
rect 1080 16232 1120 16264
rect 1152 16232 1192 16264
rect 1224 16232 1264 16264
rect 1296 16232 1336 16264
rect 1368 16232 1408 16264
rect 1440 16232 1480 16264
rect 1512 16232 1552 16264
rect 1584 16232 1624 16264
rect 1656 16232 1696 16264
rect 1728 16232 1768 16264
rect 1800 16232 1840 16264
rect 1872 16232 1912 16264
rect 1944 16232 1984 16264
rect 2016 16232 2056 16264
rect 2088 16232 2128 16264
rect 2160 16232 2200 16264
rect 2232 16232 2272 16264
rect 2304 16232 2344 16264
rect 2376 16232 2416 16264
rect 2448 16232 2488 16264
rect 2520 16232 2560 16264
rect 2592 16232 2632 16264
rect 2664 16232 2704 16264
rect 2736 16232 2776 16264
rect 2808 16232 2848 16264
rect 2880 16232 2920 16264
rect 2952 16232 2992 16264
rect 3024 16232 3064 16264
rect 3096 16232 3136 16264
rect 3168 16232 3208 16264
rect 3240 16232 3280 16264
rect 3312 16232 3352 16264
rect 3384 16232 3424 16264
rect 3456 16232 3496 16264
rect 3528 16232 3568 16264
rect 3600 16232 3640 16264
rect 3672 16232 3712 16264
rect 3744 16232 3784 16264
rect 3816 16232 3856 16264
rect 3888 16232 3950 16264
rect 50 16192 3950 16232
rect 50 16160 112 16192
rect 144 16160 184 16192
rect 216 16160 256 16192
rect 288 16160 328 16192
rect 360 16160 400 16192
rect 432 16160 472 16192
rect 504 16160 544 16192
rect 576 16160 616 16192
rect 648 16160 688 16192
rect 720 16160 760 16192
rect 792 16160 832 16192
rect 864 16160 904 16192
rect 936 16160 976 16192
rect 1008 16160 1048 16192
rect 1080 16160 1120 16192
rect 1152 16160 1192 16192
rect 1224 16160 1264 16192
rect 1296 16160 1336 16192
rect 1368 16160 1408 16192
rect 1440 16160 1480 16192
rect 1512 16160 1552 16192
rect 1584 16160 1624 16192
rect 1656 16160 1696 16192
rect 1728 16160 1768 16192
rect 1800 16160 1840 16192
rect 1872 16160 1912 16192
rect 1944 16160 1984 16192
rect 2016 16160 2056 16192
rect 2088 16160 2128 16192
rect 2160 16160 2200 16192
rect 2232 16160 2272 16192
rect 2304 16160 2344 16192
rect 2376 16160 2416 16192
rect 2448 16160 2488 16192
rect 2520 16160 2560 16192
rect 2592 16160 2632 16192
rect 2664 16160 2704 16192
rect 2736 16160 2776 16192
rect 2808 16160 2848 16192
rect 2880 16160 2920 16192
rect 2952 16160 2992 16192
rect 3024 16160 3064 16192
rect 3096 16160 3136 16192
rect 3168 16160 3208 16192
rect 3240 16160 3280 16192
rect 3312 16160 3352 16192
rect 3384 16160 3424 16192
rect 3456 16160 3496 16192
rect 3528 16160 3568 16192
rect 3600 16160 3640 16192
rect 3672 16160 3712 16192
rect 3744 16160 3784 16192
rect 3816 16160 3856 16192
rect 3888 16160 3950 16192
rect 50 16120 3950 16160
rect 50 16088 112 16120
rect 144 16088 184 16120
rect 216 16088 256 16120
rect 288 16088 328 16120
rect 360 16088 400 16120
rect 432 16088 472 16120
rect 504 16088 544 16120
rect 576 16088 616 16120
rect 648 16088 688 16120
rect 720 16088 760 16120
rect 792 16088 832 16120
rect 864 16088 904 16120
rect 936 16088 976 16120
rect 1008 16088 1048 16120
rect 1080 16088 1120 16120
rect 1152 16088 1192 16120
rect 1224 16088 1264 16120
rect 1296 16088 1336 16120
rect 1368 16088 1408 16120
rect 1440 16088 1480 16120
rect 1512 16088 1552 16120
rect 1584 16088 1624 16120
rect 1656 16088 1696 16120
rect 1728 16088 1768 16120
rect 1800 16088 1840 16120
rect 1872 16088 1912 16120
rect 1944 16088 1984 16120
rect 2016 16088 2056 16120
rect 2088 16088 2128 16120
rect 2160 16088 2200 16120
rect 2232 16088 2272 16120
rect 2304 16088 2344 16120
rect 2376 16088 2416 16120
rect 2448 16088 2488 16120
rect 2520 16088 2560 16120
rect 2592 16088 2632 16120
rect 2664 16088 2704 16120
rect 2736 16088 2776 16120
rect 2808 16088 2848 16120
rect 2880 16088 2920 16120
rect 2952 16088 2992 16120
rect 3024 16088 3064 16120
rect 3096 16088 3136 16120
rect 3168 16088 3208 16120
rect 3240 16088 3280 16120
rect 3312 16088 3352 16120
rect 3384 16088 3424 16120
rect 3456 16088 3496 16120
rect 3528 16088 3568 16120
rect 3600 16088 3640 16120
rect 3672 16088 3712 16120
rect 3744 16088 3784 16120
rect 3816 16088 3856 16120
rect 3888 16088 3950 16120
rect 50 16048 3950 16088
rect 50 16016 112 16048
rect 144 16016 184 16048
rect 216 16016 256 16048
rect 288 16016 328 16048
rect 360 16016 400 16048
rect 432 16016 472 16048
rect 504 16016 544 16048
rect 576 16016 616 16048
rect 648 16016 688 16048
rect 720 16016 760 16048
rect 792 16016 832 16048
rect 864 16016 904 16048
rect 936 16016 976 16048
rect 1008 16016 1048 16048
rect 1080 16016 1120 16048
rect 1152 16016 1192 16048
rect 1224 16016 1264 16048
rect 1296 16016 1336 16048
rect 1368 16016 1408 16048
rect 1440 16016 1480 16048
rect 1512 16016 1552 16048
rect 1584 16016 1624 16048
rect 1656 16016 1696 16048
rect 1728 16016 1768 16048
rect 1800 16016 1840 16048
rect 1872 16016 1912 16048
rect 1944 16016 1984 16048
rect 2016 16016 2056 16048
rect 2088 16016 2128 16048
rect 2160 16016 2200 16048
rect 2232 16016 2272 16048
rect 2304 16016 2344 16048
rect 2376 16016 2416 16048
rect 2448 16016 2488 16048
rect 2520 16016 2560 16048
rect 2592 16016 2632 16048
rect 2664 16016 2704 16048
rect 2736 16016 2776 16048
rect 2808 16016 2848 16048
rect 2880 16016 2920 16048
rect 2952 16016 2992 16048
rect 3024 16016 3064 16048
rect 3096 16016 3136 16048
rect 3168 16016 3208 16048
rect 3240 16016 3280 16048
rect 3312 16016 3352 16048
rect 3384 16016 3424 16048
rect 3456 16016 3496 16048
rect 3528 16016 3568 16048
rect 3600 16016 3640 16048
rect 3672 16016 3712 16048
rect 3744 16016 3784 16048
rect 3816 16016 3856 16048
rect 3888 16016 3950 16048
rect 50 15976 3950 16016
rect 50 15944 112 15976
rect 144 15944 184 15976
rect 216 15944 256 15976
rect 288 15944 328 15976
rect 360 15944 400 15976
rect 432 15944 472 15976
rect 504 15944 544 15976
rect 576 15944 616 15976
rect 648 15944 688 15976
rect 720 15944 760 15976
rect 792 15944 832 15976
rect 864 15944 904 15976
rect 936 15944 976 15976
rect 1008 15944 1048 15976
rect 1080 15944 1120 15976
rect 1152 15944 1192 15976
rect 1224 15944 1264 15976
rect 1296 15944 1336 15976
rect 1368 15944 1408 15976
rect 1440 15944 1480 15976
rect 1512 15944 1552 15976
rect 1584 15944 1624 15976
rect 1656 15944 1696 15976
rect 1728 15944 1768 15976
rect 1800 15944 1840 15976
rect 1872 15944 1912 15976
rect 1944 15944 1984 15976
rect 2016 15944 2056 15976
rect 2088 15944 2128 15976
rect 2160 15944 2200 15976
rect 2232 15944 2272 15976
rect 2304 15944 2344 15976
rect 2376 15944 2416 15976
rect 2448 15944 2488 15976
rect 2520 15944 2560 15976
rect 2592 15944 2632 15976
rect 2664 15944 2704 15976
rect 2736 15944 2776 15976
rect 2808 15944 2848 15976
rect 2880 15944 2920 15976
rect 2952 15944 2992 15976
rect 3024 15944 3064 15976
rect 3096 15944 3136 15976
rect 3168 15944 3208 15976
rect 3240 15944 3280 15976
rect 3312 15944 3352 15976
rect 3384 15944 3424 15976
rect 3456 15944 3496 15976
rect 3528 15944 3568 15976
rect 3600 15944 3640 15976
rect 3672 15944 3712 15976
rect 3744 15944 3784 15976
rect 3816 15944 3856 15976
rect 3888 15944 3950 15976
rect 50 15904 3950 15944
rect 50 15872 112 15904
rect 144 15872 184 15904
rect 216 15872 256 15904
rect 288 15872 328 15904
rect 360 15872 400 15904
rect 432 15872 472 15904
rect 504 15872 544 15904
rect 576 15872 616 15904
rect 648 15872 688 15904
rect 720 15872 760 15904
rect 792 15872 832 15904
rect 864 15872 904 15904
rect 936 15872 976 15904
rect 1008 15872 1048 15904
rect 1080 15872 1120 15904
rect 1152 15872 1192 15904
rect 1224 15872 1264 15904
rect 1296 15872 1336 15904
rect 1368 15872 1408 15904
rect 1440 15872 1480 15904
rect 1512 15872 1552 15904
rect 1584 15872 1624 15904
rect 1656 15872 1696 15904
rect 1728 15872 1768 15904
rect 1800 15872 1840 15904
rect 1872 15872 1912 15904
rect 1944 15872 1984 15904
rect 2016 15872 2056 15904
rect 2088 15872 2128 15904
rect 2160 15872 2200 15904
rect 2232 15872 2272 15904
rect 2304 15872 2344 15904
rect 2376 15872 2416 15904
rect 2448 15872 2488 15904
rect 2520 15872 2560 15904
rect 2592 15872 2632 15904
rect 2664 15872 2704 15904
rect 2736 15872 2776 15904
rect 2808 15872 2848 15904
rect 2880 15872 2920 15904
rect 2952 15872 2992 15904
rect 3024 15872 3064 15904
rect 3096 15872 3136 15904
rect 3168 15872 3208 15904
rect 3240 15872 3280 15904
rect 3312 15872 3352 15904
rect 3384 15872 3424 15904
rect 3456 15872 3496 15904
rect 3528 15872 3568 15904
rect 3600 15872 3640 15904
rect 3672 15872 3712 15904
rect 3744 15872 3784 15904
rect 3816 15872 3856 15904
rect 3888 15872 3950 15904
rect 50 15832 3950 15872
rect 50 15800 112 15832
rect 144 15800 184 15832
rect 216 15800 256 15832
rect 288 15800 328 15832
rect 360 15800 400 15832
rect 432 15800 472 15832
rect 504 15800 544 15832
rect 576 15800 616 15832
rect 648 15800 688 15832
rect 720 15800 760 15832
rect 792 15800 832 15832
rect 864 15800 904 15832
rect 936 15800 976 15832
rect 1008 15800 1048 15832
rect 1080 15800 1120 15832
rect 1152 15800 1192 15832
rect 1224 15800 1264 15832
rect 1296 15800 1336 15832
rect 1368 15800 1408 15832
rect 1440 15800 1480 15832
rect 1512 15800 1552 15832
rect 1584 15800 1624 15832
rect 1656 15800 1696 15832
rect 1728 15800 1768 15832
rect 1800 15800 1840 15832
rect 1872 15800 1912 15832
rect 1944 15800 1984 15832
rect 2016 15800 2056 15832
rect 2088 15800 2128 15832
rect 2160 15800 2200 15832
rect 2232 15800 2272 15832
rect 2304 15800 2344 15832
rect 2376 15800 2416 15832
rect 2448 15800 2488 15832
rect 2520 15800 2560 15832
rect 2592 15800 2632 15832
rect 2664 15800 2704 15832
rect 2736 15800 2776 15832
rect 2808 15800 2848 15832
rect 2880 15800 2920 15832
rect 2952 15800 2992 15832
rect 3024 15800 3064 15832
rect 3096 15800 3136 15832
rect 3168 15800 3208 15832
rect 3240 15800 3280 15832
rect 3312 15800 3352 15832
rect 3384 15800 3424 15832
rect 3456 15800 3496 15832
rect 3528 15800 3568 15832
rect 3600 15800 3640 15832
rect 3672 15800 3712 15832
rect 3744 15800 3784 15832
rect 3816 15800 3856 15832
rect 3888 15800 3950 15832
rect 50 15760 3950 15800
rect 50 15728 112 15760
rect 144 15728 184 15760
rect 216 15728 256 15760
rect 288 15728 328 15760
rect 360 15728 400 15760
rect 432 15728 472 15760
rect 504 15728 544 15760
rect 576 15728 616 15760
rect 648 15728 688 15760
rect 720 15728 760 15760
rect 792 15728 832 15760
rect 864 15728 904 15760
rect 936 15728 976 15760
rect 1008 15728 1048 15760
rect 1080 15728 1120 15760
rect 1152 15728 1192 15760
rect 1224 15728 1264 15760
rect 1296 15728 1336 15760
rect 1368 15728 1408 15760
rect 1440 15728 1480 15760
rect 1512 15728 1552 15760
rect 1584 15728 1624 15760
rect 1656 15728 1696 15760
rect 1728 15728 1768 15760
rect 1800 15728 1840 15760
rect 1872 15728 1912 15760
rect 1944 15728 1984 15760
rect 2016 15728 2056 15760
rect 2088 15728 2128 15760
rect 2160 15728 2200 15760
rect 2232 15728 2272 15760
rect 2304 15728 2344 15760
rect 2376 15728 2416 15760
rect 2448 15728 2488 15760
rect 2520 15728 2560 15760
rect 2592 15728 2632 15760
rect 2664 15728 2704 15760
rect 2736 15728 2776 15760
rect 2808 15728 2848 15760
rect 2880 15728 2920 15760
rect 2952 15728 2992 15760
rect 3024 15728 3064 15760
rect 3096 15728 3136 15760
rect 3168 15728 3208 15760
rect 3240 15728 3280 15760
rect 3312 15728 3352 15760
rect 3384 15728 3424 15760
rect 3456 15728 3496 15760
rect 3528 15728 3568 15760
rect 3600 15728 3640 15760
rect 3672 15728 3712 15760
rect 3744 15728 3784 15760
rect 3816 15728 3856 15760
rect 3888 15728 3950 15760
rect 50 15688 3950 15728
rect 50 15656 112 15688
rect 144 15656 184 15688
rect 216 15656 256 15688
rect 288 15656 328 15688
rect 360 15656 400 15688
rect 432 15656 472 15688
rect 504 15656 544 15688
rect 576 15656 616 15688
rect 648 15656 688 15688
rect 720 15656 760 15688
rect 792 15656 832 15688
rect 864 15656 904 15688
rect 936 15656 976 15688
rect 1008 15656 1048 15688
rect 1080 15656 1120 15688
rect 1152 15656 1192 15688
rect 1224 15656 1264 15688
rect 1296 15656 1336 15688
rect 1368 15656 1408 15688
rect 1440 15656 1480 15688
rect 1512 15656 1552 15688
rect 1584 15656 1624 15688
rect 1656 15656 1696 15688
rect 1728 15656 1768 15688
rect 1800 15656 1840 15688
rect 1872 15656 1912 15688
rect 1944 15656 1984 15688
rect 2016 15656 2056 15688
rect 2088 15656 2128 15688
rect 2160 15656 2200 15688
rect 2232 15656 2272 15688
rect 2304 15656 2344 15688
rect 2376 15656 2416 15688
rect 2448 15656 2488 15688
rect 2520 15656 2560 15688
rect 2592 15656 2632 15688
rect 2664 15656 2704 15688
rect 2736 15656 2776 15688
rect 2808 15656 2848 15688
rect 2880 15656 2920 15688
rect 2952 15656 2992 15688
rect 3024 15656 3064 15688
rect 3096 15656 3136 15688
rect 3168 15656 3208 15688
rect 3240 15656 3280 15688
rect 3312 15656 3352 15688
rect 3384 15656 3424 15688
rect 3456 15656 3496 15688
rect 3528 15656 3568 15688
rect 3600 15656 3640 15688
rect 3672 15656 3712 15688
rect 3744 15656 3784 15688
rect 3816 15656 3856 15688
rect 3888 15656 3950 15688
rect 50 15616 3950 15656
rect 50 15584 112 15616
rect 144 15584 184 15616
rect 216 15584 256 15616
rect 288 15584 328 15616
rect 360 15584 400 15616
rect 432 15584 472 15616
rect 504 15584 544 15616
rect 576 15584 616 15616
rect 648 15584 688 15616
rect 720 15584 760 15616
rect 792 15584 832 15616
rect 864 15584 904 15616
rect 936 15584 976 15616
rect 1008 15584 1048 15616
rect 1080 15584 1120 15616
rect 1152 15584 1192 15616
rect 1224 15584 1264 15616
rect 1296 15584 1336 15616
rect 1368 15584 1408 15616
rect 1440 15584 1480 15616
rect 1512 15584 1552 15616
rect 1584 15584 1624 15616
rect 1656 15584 1696 15616
rect 1728 15584 1768 15616
rect 1800 15584 1840 15616
rect 1872 15584 1912 15616
rect 1944 15584 1984 15616
rect 2016 15584 2056 15616
rect 2088 15584 2128 15616
rect 2160 15584 2200 15616
rect 2232 15584 2272 15616
rect 2304 15584 2344 15616
rect 2376 15584 2416 15616
rect 2448 15584 2488 15616
rect 2520 15584 2560 15616
rect 2592 15584 2632 15616
rect 2664 15584 2704 15616
rect 2736 15584 2776 15616
rect 2808 15584 2848 15616
rect 2880 15584 2920 15616
rect 2952 15584 2992 15616
rect 3024 15584 3064 15616
rect 3096 15584 3136 15616
rect 3168 15584 3208 15616
rect 3240 15584 3280 15616
rect 3312 15584 3352 15616
rect 3384 15584 3424 15616
rect 3456 15584 3496 15616
rect 3528 15584 3568 15616
rect 3600 15584 3640 15616
rect 3672 15584 3712 15616
rect 3744 15584 3784 15616
rect 3816 15584 3856 15616
rect 3888 15584 3950 15616
rect 50 15544 3950 15584
rect 50 15512 112 15544
rect 144 15512 184 15544
rect 216 15512 256 15544
rect 288 15512 328 15544
rect 360 15512 400 15544
rect 432 15512 472 15544
rect 504 15512 544 15544
rect 576 15512 616 15544
rect 648 15512 688 15544
rect 720 15512 760 15544
rect 792 15512 832 15544
rect 864 15512 904 15544
rect 936 15512 976 15544
rect 1008 15512 1048 15544
rect 1080 15512 1120 15544
rect 1152 15512 1192 15544
rect 1224 15512 1264 15544
rect 1296 15512 1336 15544
rect 1368 15512 1408 15544
rect 1440 15512 1480 15544
rect 1512 15512 1552 15544
rect 1584 15512 1624 15544
rect 1656 15512 1696 15544
rect 1728 15512 1768 15544
rect 1800 15512 1840 15544
rect 1872 15512 1912 15544
rect 1944 15512 1984 15544
rect 2016 15512 2056 15544
rect 2088 15512 2128 15544
rect 2160 15512 2200 15544
rect 2232 15512 2272 15544
rect 2304 15512 2344 15544
rect 2376 15512 2416 15544
rect 2448 15512 2488 15544
rect 2520 15512 2560 15544
rect 2592 15512 2632 15544
rect 2664 15512 2704 15544
rect 2736 15512 2776 15544
rect 2808 15512 2848 15544
rect 2880 15512 2920 15544
rect 2952 15512 2992 15544
rect 3024 15512 3064 15544
rect 3096 15512 3136 15544
rect 3168 15512 3208 15544
rect 3240 15512 3280 15544
rect 3312 15512 3352 15544
rect 3384 15512 3424 15544
rect 3456 15512 3496 15544
rect 3528 15512 3568 15544
rect 3600 15512 3640 15544
rect 3672 15512 3712 15544
rect 3744 15512 3784 15544
rect 3816 15512 3856 15544
rect 3888 15512 3950 15544
rect 50 15472 3950 15512
rect 50 15440 112 15472
rect 144 15440 184 15472
rect 216 15440 256 15472
rect 288 15440 328 15472
rect 360 15440 400 15472
rect 432 15440 472 15472
rect 504 15440 544 15472
rect 576 15440 616 15472
rect 648 15440 688 15472
rect 720 15440 760 15472
rect 792 15440 832 15472
rect 864 15440 904 15472
rect 936 15440 976 15472
rect 1008 15440 1048 15472
rect 1080 15440 1120 15472
rect 1152 15440 1192 15472
rect 1224 15440 1264 15472
rect 1296 15440 1336 15472
rect 1368 15440 1408 15472
rect 1440 15440 1480 15472
rect 1512 15440 1552 15472
rect 1584 15440 1624 15472
rect 1656 15440 1696 15472
rect 1728 15440 1768 15472
rect 1800 15440 1840 15472
rect 1872 15440 1912 15472
rect 1944 15440 1984 15472
rect 2016 15440 2056 15472
rect 2088 15440 2128 15472
rect 2160 15440 2200 15472
rect 2232 15440 2272 15472
rect 2304 15440 2344 15472
rect 2376 15440 2416 15472
rect 2448 15440 2488 15472
rect 2520 15440 2560 15472
rect 2592 15440 2632 15472
rect 2664 15440 2704 15472
rect 2736 15440 2776 15472
rect 2808 15440 2848 15472
rect 2880 15440 2920 15472
rect 2952 15440 2992 15472
rect 3024 15440 3064 15472
rect 3096 15440 3136 15472
rect 3168 15440 3208 15472
rect 3240 15440 3280 15472
rect 3312 15440 3352 15472
rect 3384 15440 3424 15472
rect 3456 15440 3496 15472
rect 3528 15440 3568 15472
rect 3600 15440 3640 15472
rect 3672 15440 3712 15472
rect 3744 15440 3784 15472
rect 3816 15440 3856 15472
rect 3888 15440 3950 15472
rect 50 15400 3950 15440
rect 50 15368 112 15400
rect 144 15368 184 15400
rect 216 15368 256 15400
rect 288 15368 328 15400
rect 360 15368 400 15400
rect 432 15368 472 15400
rect 504 15368 544 15400
rect 576 15368 616 15400
rect 648 15368 688 15400
rect 720 15368 760 15400
rect 792 15368 832 15400
rect 864 15368 904 15400
rect 936 15368 976 15400
rect 1008 15368 1048 15400
rect 1080 15368 1120 15400
rect 1152 15368 1192 15400
rect 1224 15368 1264 15400
rect 1296 15368 1336 15400
rect 1368 15368 1408 15400
rect 1440 15368 1480 15400
rect 1512 15368 1552 15400
rect 1584 15368 1624 15400
rect 1656 15368 1696 15400
rect 1728 15368 1768 15400
rect 1800 15368 1840 15400
rect 1872 15368 1912 15400
rect 1944 15368 1984 15400
rect 2016 15368 2056 15400
rect 2088 15368 2128 15400
rect 2160 15368 2200 15400
rect 2232 15368 2272 15400
rect 2304 15368 2344 15400
rect 2376 15368 2416 15400
rect 2448 15368 2488 15400
rect 2520 15368 2560 15400
rect 2592 15368 2632 15400
rect 2664 15368 2704 15400
rect 2736 15368 2776 15400
rect 2808 15368 2848 15400
rect 2880 15368 2920 15400
rect 2952 15368 2992 15400
rect 3024 15368 3064 15400
rect 3096 15368 3136 15400
rect 3168 15368 3208 15400
rect 3240 15368 3280 15400
rect 3312 15368 3352 15400
rect 3384 15368 3424 15400
rect 3456 15368 3496 15400
rect 3528 15368 3568 15400
rect 3600 15368 3640 15400
rect 3672 15368 3712 15400
rect 3744 15368 3784 15400
rect 3816 15368 3856 15400
rect 3888 15368 3950 15400
rect 50 15328 3950 15368
rect 50 15296 112 15328
rect 144 15296 184 15328
rect 216 15296 256 15328
rect 288 15296 328 15328
rect 360 15296 400 15328
rect 432 15296 472 15328
rect 504 15296 544 15328
rect 576 15296 616 15328
rect 648 15296 688 15328
rect 720 15296 760 15328
rect 792 15296 832 15328
rect 864 15296 904 15328
rect 936 15296 976 15328
rect 1008 15296 1048 15328
rect 1080 15296 1120 15328
rect 1152 15296 1192 15328
rect 1224 15296 1264 15328
rect 1296 15296 1336 15328
rect 1368 15296 1408 15328
rect 1440 15296 1480 15328
rect 1512 15296 1552 15328
rect 1584 15296 1624 15328
rect 1656 15296 1696 15328
rect 1728 15296 1768 15328
rect 1800 15296 1840 15328
rect 1872 15296 1912 15328
rect 1944 15296 1984 15328
rect 2016 15296 2056 15328
rect 2088 15296 2128 15328
rect 2160 15296 2200 15328
rect 2232 15296 2272 15328
rect 2304 15296 2344 15328
rect 2376 15296 2416 15328
rect 2448 15296 2488 15328
rect 2520 15296 2560 15328
rect 2592 15296 2632 15328
rect 2664 15296 2704 15328
rect 2736 15296 2776 15328
rect 2808 15296 2848 15328
rect 2880 15296 2920 15328
rect 2952 15296 2992 15328
rect 3024 15296 3064 15328
rect 3096 15296 3136 15328
rect 3168 15296 3208 15328
rect 3240 15296 3280 15328
rect 3312 15296 3352 15328
rect 3384 15296 3424 15328
rect 3456 15296 3496 15328
rect 3528 15296 3568 15328
rect 3600 15296 3640 15328
rect 3672 15296 3712 15328
rect 3744 15296 3784 15328
rect 3816 15296 3856 15328
rect 3888 15296 3950 15328
rect 50 15256 3950 15296
rect 50 15224 112 15256
rect 144 15224 184 15256
rect 216 15224 256 15256
rect 288 15224 328 15256
rect 360 15224 400 15256
rect 432 15224 472 15256
rect 504 15224 544 15256
rect 576 15224 616 15256
rect 648 15224 688 15256
rect 720 15224 760 15256
rect 792 15224 832 15256
rect 864 15224 904 15256
rect 936 15224 976 15256
rect 1008 15224 1048 15256
rect 1080 15224 1120 15256
rect 1152 15224 1192 15256
rect 1224 15224 1264 15256
rect 1296 15224 1336 15256
rect 1368 15224 1408 15256
rect 1440 15224 1480 15256
rect 1512 15224 1552 15256
rect 1584 15224 1624 15256
rect 1656 15224 1696 15256
rect 1728 15224 1768 15256
rect 1800 15224 1840 15256
rect 1872 15224 1912 15256
rect 1944 15224 1984 15256
rect 2016 15224 2056 15256
rect 2088 15224 2128 15256
rect 2160 15224 2200 15256
rect 2232 15224 2272 15256
rect 2304 15224 2344 15256
rect 2376 15224 2416 15256
rect 2448 15224 2488 15256
rect 2520 15224 2560 15256
rect 2592 15224 2632 15256
rect 2664 15224 2704 15256
rect 2736 15224 2776 15256
rect 2808 15224 2848 15256
rect 2880 15224 2920 15256
rect 2952 15224 2992 15256
rect 3024 15224 3064 15256
rect 3096 15224 3136 15256
rect 3168 15224 3208 15256
rect 3240 15224 3280 15256
rect 3312 15224 3352 15256
rect 3384 15224 3424 15256
rect 3456 15224 3496 15256
rect 3528 15224 3568 15256
rect 3600 15224 3640 15256
rect 3672 15224 3712 15256
rect 3744 15224 3784 15256
rect 3816 15224 3856 15256
rect 3888 15224 3950 15256
rect 50 15184 3950 15224
rect 50 15152 112 15184
rect 144 15152 184 15184
rect 216 15152 256 15184
rect 288 15152 328 15184
rect 360 15152 400 15184
rect 432 15152 472 15184
rect 504 15152 544 15184
rect 576 15152 616 15184
rect 648 15152 688 15184
rect 720 15152 760 15184
rect 792 15152 832 15184
rect 864 15152 904 15184
rect 936 15152 976 15184
rect 1008 15152 1048 15184
rect 1080 15152 1120 15184
rect 1152 15152 1192 15184
rect 1224 15152 1264 15184
rect 1296 15152 1336 15184
rect 1368 15152 1408 15184
rect 1440 15152 1480 15184
rect 1512 15152 1552 15184
rect 1584 15152 1624 15184
rect 1656 15152 1696 15184
rect 1728 15152 1768 15184
rect 1800 15152 1840 15184
rect 1872 15152 1912 15184
rect 1944 15152 1984 15184
rect 2016 15152 2056 15184
rect 2088 15152 2128 15184
rect 2160 15152 2200 15184
rect 2232 15152 2272 15184
rect 2304 15152 2344 15184
rect 2376 15152 2416 15184
rect 2448 15152 2488 15184
rect 2520 15152 2560 15184
rect 2592 15152 2632 15184
rect 2664 15152 2704 15184
rect 2736 15152 2776 15184
rect 2808 15152 2848 15184
rect 2880 15152 2920 15184
rect 2952 15152 2992 15184
rect 3024 15152 3064 15184
rect 3096 15152 3136 15184
rect 3168 15152 3208 15184
rect 3240 15152 3280 15184
rect 3312 15152 3352 15184
rect 3384 15152 3424 15184
rect 3456 15152 3496 15184
rect 3528 15152 3568 15184
rect 3600 15152 3640 15184
rect 3672 15152 3712 15184
rect 3744 15152 3784 15184
rect 3816 15152 3856 15184
rect 3888 15152 3950 15184
rect 50 15112 3950 15152
rect 50 15080 112 15112
rect 144 15080 184 15112
rect 216 15080 256 15112
rect 288 15080 328 15112
rect 360 15080 400 15112
rect 432 15080 472 15112
rect 504 15080 544 15112
rect 576 15080 616 15112
rect 648 15080 688 15112
rect 720 15080 760 15112
rect 792 15080 832 15112
rect 864 15080 904 15112
rect 936 15080 976 15112
rect 1008 15080 1048 15112
rect 1080 15080 1120 15112
rect 1152 15080 1192 15112
rect 1224 15080 1264 15112
rect 1296 15080 1336 15112
rect 1368 15080 1408 15112
rect 1440 15080 1480 15112
rect 1512 15080 1552 15112
rect 1584 15080 1624 15112
rect 1656 15080 1696 15112
rect 1728 15080 1768 15112
rect 1800 15080 1840 15112
rect 1872 15080 1912 15112
rect 1944 15080 1984 15112
rect 2016 15080 2056 15112
rect 2088 15080 2128 15112
rect 2160 15080 2200 15112
rect 2232 15080 2272 15112
rect 2304 15080 2344 15112
rect 2376 15080 2416 15112
rect 2448 15080 2488 15112
rect 2520 15080 2560 15112
rect 2592 15080 2632 15112
rect 2664 15080 2704 15112
rect 2736 15080 2776 15112
rect 2808 15080 2848 15112
rect 2880 15080 2920 15112
rect 2952 15080 2992 15112
rect 3024 15080 3064 15112
rect 3096 15080 3136 15112
rect 3168 15080 3208 15112
rect 3240 15080 3280 15112
rect 3312 15080 3352 15112
rect 3384 15080 3424 15112
rect 3456 15080 3496 15112
rect 3528 15080 3568 15112
rect 3600 15080 3640 15112
rect 3672 15080 3712 15112
rect 3744 15080 3784 15112
rect 3816 15080 3856 15112
rect 3888 15080 3950 15112
rect 50 15040 3950 15080
rect 50 15008 112 15040
rect 144 15008 184 15040
rect 216 15008 256 15040
rect 288 15008 328 15040
rect 360 15008 400 15040
rect 432 15008 472 15040
rect 504 15008 544 15040
rect 576 15008 616 15040
rect 648 15008 688 15040
rect 720 15008 760 15040
rect 792 15008 832 15040
rect 864 15008 904 15040
rect 936 15008 976 15040
rect 1008 15008 1048 15040
rect 1080 15008 1120 15040
rect 1152 15008 1192 15040
rect 1224 15008 1264 15040
rect 1296 15008 1336 15040
rect 1368 15008 1408 15040
rect 1440 15008 1480 15040
rect 1512 15008 1552 15040
rect 1584 15008 1624 15040
rect 1656 15008 1696 15040
rect 1728 15008 1768 15040
rect 1800 15008 1840 15040
rect 1872 15008 1912 15040
rect 1944 15008 1984 15040
rect 2016 15008 2056 15040
rect 2088 15008 2128 15040
rect 2160 15008 2200 15040
rect 2232 15008 2272 15040
rect 2304 15008 2344 15040
rect 2376 15008 2416 15040
rect 2448 15008 2488 15040
rect 2520 15008 2560 15040
rect 2592 15008 2632 15040
rect 2664 15008 2704 15040
rect 2736 15008 2776 15040
rect 2808 15008 2848 15040
rect 2880 15008 2920 15040
rect 2952 15008 2992 15040
rect 3024 15008 3064 15040
rect 3096 15008 3136 15040
rect 3168 15008 3208 15040
rect 3240 15008 3280 15040
rect 3312 15008 3352 15040
rect 3384 15008 3424 15040
rect 3456 15008 3496 15040
rect 3528 15008 3568 15040
rect 3600 15008 3640 15040
rect 3672 15008 3712 15040
rect 3744 15008 3784 15040
rect 3816 15008 3856 15040
rect 3888 15008 3950 15040
rect 50 14968 3950 15008
rect 50 14936 112 14968
rect 144 14936 184 14968
rect 216 14936 256 14968
rect 288 14936 328 14968
rect 360 14936 400 14968
rect 432 14936 472 14968
rect 504 14936 544 14968
rect 576 14936 616 14968
rect 648 14936 688 14968
rect 720 14936 760 14968
rect 792 14936 832 14968
rect 864 14936 904 14968
rect 936 14936 976 14968
rect 1008 14936 1048 14968
rect 1080 14936 1120 14968
rect 1152 14936 1192 14968
rect 1224 14936 1264 14968
rect 1296 14936 1336 14968
rect 1368 14936 1408 14968
rect 1440 14936 1480 14968
rect 1512 14936 1552 14968
rect 1584 14936 1624 14968
rect 1656 14936 1696 14968
rect 1728 14936 1768 14968
rect 1800 14936 1840 14968
rect 1872 14936 1912 14968
rect 1944 14936 1984 14968
rect 2016 14936 2056 14968
rect 2088 14936 2128 14968
rect 2160 14936 2200 14968
rect 2232 14936 2272 14968
rect 2304 14936 2344 14968
rect 2376 14936 2416 14968
rect 2448 14936 2488 14968
rect 2520 14936 2560 14968
rect 2592 14936 2632 14968
rect 2664 14936 2704 14968
rect 2736 14936 2776 14968
rect 2808 14936 2848 14968
rect 2880 14936 2920 14968
rect 2952 14936 2992 14968
rect 3024 14936 3064 14968
rect 3096 14936 3136 14968
rect 3168 14936 3208 14968
rect 3240 14936 3280 14968
rect 3312 14936 3352 14968
rect 3384 14936 3424 14968
rect 3456 14936 3496 14968
rect 3528 14936 3568 14968
rect 3600 14936 3640 14968
rect 3672 14936 3712 14968
rect 3744 14936 3784 14968
rect 3816 14936 3856 14968
rect 3888 14936 3950 14968
rect 50 14896 3950 14936
rect 50 14864 112 14896
rect 144 14864 184 14896
rect 216 14864 256 14896
rect 288 14864 328 14896
rect 360 14864 400 14896
rect 432 14864 472 14896
rect 504 14864 544 14896
rect 576 14864 616 14896
rect 648 14864 688 14896
rect 720 14864 760 14896
rect 792 14864 832 14896
rect 864 14864 904 14896
rect 936 14864 976 14896
rect 1008 14864 1048 14896
rect 1080 14864 1120 14896
rect 1152 14864 1192 14896
rect 1224 14864 1264 14896
rect 1296 14864 1336 14896
rect 1368 14864 1408 14896
rect 1440 14864 1480 14896
rect 1512 14864 1552 14896
rect 1584 14864 1624 14896
rect 1656 14864 1696 14896
rect 1728 14864 1768 14896
rect 1800 14864 1840 14896
rect 1872 14864 1912 14896
rect 1944 14864 1984 14896
rect 2016 14864 2056 14896
rect 2088 14864 2128 14896
rect 2160 14864 2200 14896
rect 2232 14864 2272 14896
rect 2304 14864 2344 14896
rect 2376 14864 2416 14896
rect 2448 14864 2488 14896
rect 2520 14864 2560 14896
rect 2592 14864 2632 14896
rect 2664 14864 2704 14896
rect 2736 14864 2776 14896
rect 2808 14864 2848 14896
rect 2880 14864 2920 14896
rect 2952 14864 2992 14896
rect 3024 14864 3064 14896
rect 3096 14864 3136 14896
rect 3168 14864 3208 14896
rect 3240 14864 3280 14896
rect 3312 14864 3352 14896
rect 3384 14864 3424 14896
rect 3456 14864 3496 14896
rect 3528 14864 3568 14896
rect 3600 14864 3640 14896
rect 3672 14864 3712 14896
rect 3744 14864 3784 14896
rect 3816 14864 3856 14896
rect 3888 14864 3950 14896
rect 50 14824 3950 14864
rect 50 14792 112 14824
rect 144 14792 184 14824
rect 216 14792 256 14824
rect 288 14792 328 14824
rect 360 14792 400 14824
rect 432 14792 472 14824
rect 504 14792 544 14824
rect 576 14792 616 14824
rect 648 14792 688 14824
rect 720 14792 760 14824
rect 792 14792 832 14824
rect 864 14792 904 14824
rect 936 14792 976 14824
rect 1008 14792 1048 14824
rect 1080 14792 1120 14824
rect 1152 14792 1192 14824
rect 1224 14792 1264 14824
rect 1296 14792 1336 14824
rect 1368 14792 1408 14824
rect 1440 14792 1480 14824
rect 1512 14792 1552 14824
rect 1584 14792 1624 14824
rect 1656 14792 1696 14824
rect 1728 14792 1768 14824
rect 1800 14792 1840 14824
rect 1872 14792 1912 14824
rect 1944 14792 1984 14824
rect 2016 14792 2056 14824
rect 2088 14792 2128 14824
rect 2160 14792 2200 14824
rect 2232 14792 2272 14824
rect 2304 14792 2344 14824
rect 2376 14792 2416 14824
rect 2448 14792 2488 14824
rect 2520 14792 2560 14824
rect 2592 14792 2632 14824
rect 2664 14792 2704 14824
rect 2736 14792 2776 14824
rect 2808 14792 2848 14824
rect 2880 14792 2920 14824
rect 2952 14792 2992 14824
rect 3024 14792 3064 14824
rect 3096 14792 3136 14824
rect 3168 14792 3208 14824
rect 3240 14792 3280 14824
rect 3312 14792 3352 14824
rect 3384 14792 3424 14824
rect 3456 14792 3496 14824
rect 3528 14792 3568 14824
rect 3600 14792 3640 14824
rect 3672 14792 3712 14824
rect 3744 14792 3784 14824
rect 3816 14792 3856 14824
rect 3888 14792 3950 14824
rect 50 14752 3950 14792
rect 50 14720 112 14752
rect 144 14720 184 14752
rect 216 14720 256 14752
rect 288 14720 328 14752
rect 360 14720 400 14752
rect 432 14720 472 14752
rect 504 14720 544 14752
rect 576 14720 616 14752
rect 648 14720 688 14752
rect 720 14720 760 14752
rect 792 14720 832 14752
rect 864 14720 904 14752
rect 936 14720 976 14752
rect 1008 14720 1048 14752
rect 1080 14720 1120 14752
rect 1152 14720 1192 14752
rect 1224 14720 1264 14752
rect 1296 14720 1336 14752
rect 1368 14720 1408 14752
rect 1440 14720 1480 14752
rect 1512 14720 1552 14752
rect 1584 14720 1624 14752
rect 1656 14720 1696 14752
rect 1728 14720 1768 14752
rect 1800 14720 1840 14752
rect 1872 14720 1912 14752
rect 1944 14720 1984 14752
rect 2016 14720 2056 14752
rect 2088 14720 2128 14752
rect 2160 14720 2200 14752
rect 2232 14720 2272 14752
rect 2304 14720 2344 14752
rect 2376 14720 2416 14752
rect 2448 14720 2488 14752
rect 2520 14720 2560 14752
rect 2592 14720 2632 14752
rect 2664 14720 2704 14752
rect 2736 14720 2776 14752
rect 2808 14720 2848 14752
rect 2880 14720 2920 14752
rect 2952 14720 2992 14752
rect 3024 14720 3064 14752
rect 3096 14720 3136 14752
rect 3168 14720 3208 14752
rect 3240 14720 3280 14752
rect 3312 14720 3352 14752
rect 3384 14720 3424 14752
rect 3456 14720 3496 14752
rect 3528 14720 3568 14752
rect 3600 14720 3640 14752
rect 3672 14720 3712 14752
rect 3744 14720 3784 14752
rect 3816 14720 3856 14752
rect 3888 14720 3950 14752
rect 50 14680 3950 14720
rect 50 14648 112 14680
rect 144 14648 184 14680
rect 216 14648 256 14680
rect 288 14648 328 14680
rect 360 14648 400 14680
rect 432 14648 472 14680
rect 504 14648 544 14680
rect 576 14648 616 14680
rect 648 14648 688 14680
rect 720 14648 760 14680
rect 792 14648 832 14680
rect 864 14648 904 14680
rect 936 14648 976 14680
rect 1008 14648 1048 14680
rect 1080 14648 1120 14680
rect 1152 14648 1192 14680
rect 1224 14648 1264 14680
rect 1296 14648 1336 14680
rect 1368 14648 1408 14680
rect 1440 14648 1480 14680
rect 1512 14648 1552 14680
rect 1584 14648 1624 14680
rect 1656 14648 1696 14680
rect 1728 14648 1768 14680
rect 1800 14648 1840 14680
rect 1872 14648 1912 14680
rect 1944 14648 1984 14680
rect 2016 14648 2056 14680
rect 2088 14648 2128 14680
rect 2160 14648 2200 14680
rect 2232 14648 2272 14680
rect 2304 14648 2344 14680
rect 2376 14648 2416 14680
rect 2448 14648 2488 14680
rect 2520 14648 2560 14680
rect 2592 14648 2632 14680
rect 2664 14648 2704 14680
rect 2736 14648 2776 14680
rect 2808 14648 2848 14680
rect 2880 14648 2920 14680
rect 2952 14648 2992 14680
rect 3024 14648 3064 14680
rect 3096 14648 3136 14680
rect 3168 14648 3208 14680
rect 3240 14648 3280 14680
rect 3312 14648 3352 14680
rect 3384 14648 3424 14680
rect 3456 14648 3496 14680
rect 3528 14648 3568 14680
rect 3600 14648 3640 14680
rect 3672 14648 3712 14680
rect 3744 14648 3784 14680
rect 3816 14648 3856 14680
rect 3888 14648 3950 14680
rect 50 14608 3950 14648
rect 50 14576 112 14608
rect 144 14576 184 14608
rect 216 14576 256 14608
rect 288 14576 328 14608
rect 360 14576 400 14608
rect 432 14576 472 14608
rect 504 14576 544 14608
rect 576 14576 616 14608
rect 648 14576 688 14608
rect 720 14576 760 14608
rect 792 14576 832 14608
rect 864 14576 904 14608
rect 936 14576 976 14608
rect 1008 14576 1048 14608
rect 1080 14576 1120 14608
rect 1152 14576 1192 14608
rect 1224 14576 1264 14608
rect 1296 14576 1336 14608
rect 1368 14576 1408 14608
rect 1440 14576 1480 14608
rect 1512 14576 1552 14608
rect 1584 14576 1624 14608
rect 1656 14576 1696 14608
rect 1728 14576 1768 14608
rect 1800 14576 1840 14608
rect 1872 14576 1912 14608
rect 1944 14576 1984 14608
rect 2016 14576 2056 14608
rect 2088 14576 2128 14608
rect 2160 14576 2200 14608
rect 2232 14576 2272 14608
rect 2304 14576 2344 14608
rect 2376 14576 2416 14608
rect 2448 14576 2488 14608
rect 2520 14576 2560 14608
rect 2592 14576 2632 14608
rect 2664 14576 2704 14608
rect 2736 14576 2776 14608
rect 2808 14576 2848 14608
rect 2880 14576 2920 14608
rect 2952 14576 2992 14608
rect 3024 14576 3064 14608
rect 3096 14576 3136 14608
rect 3168 14576 3208 14608
rect 3240 14576 3280 14608
rect 3312 14576 3352 14608
rect 3384 14576 3424 14608
rect 3456 14576 3496 14608
rect 3528 14576 3568 14608
rect 3600 14576 3640 14608
rect 3672 14576 3712 14608
rect 3744 14576 3784 14608
rect 3816 14576 3856 14608
rect 3888 14576 3950 14608
rect 50 14536 3950 14576
rect 50 14504 112 14536
rect 144 14504 184 14536
rect 216 14504 256 14536
rect 288 14504 328 14536
rect 360 14504 400 14536
rect 432 14504 472 14536
rect 504 14504 544 14536
rect 576 14504 616 14536
rect 648 14504 688 14536
rect 720 14504 760 14536
rect 792 14504 832 14536
rect 864 14504 904 14536
rect 936 14504 976 14536
rect 1008 14504 1048 14536
rect 1080 14504 1120 14536
rect 1152 14504 1192 14536
rect 1224 14504 1264 14536
rect 1296 14504 1336 14536
rect 1368 14504 1408 14536
rect 1440 14504 1480 14536
rect 1512 14504 1552 14536
rect 1584 14504 1624 14536
rect 1656 14504 1696 14536
rect 1728 14504 1768 14536
rect 1800 14504 1840 14536
rect 1872 14504 1912 14536
rect 1944 14504 1984 14536
rect 2016 14504 2056 14536
rect 2088 14504 2128 14536
rect 2160 14504 2200 14536
rect 2232 14504 2272 14536
rect 2304 14504 2344 14536
rect 2376 14504 2416 14536
rect 2448 14504 2488 14536
rect 2520 14504 2560 14536
rect 2592 14504 2632 14536
rect 2664 14504 2704 14536
rect 2736 14504 2776 14536
rect 2808 14504 2848 14536
rect 2880 14504 2920 14536
rect 2952 14504 2992 14536
rect 3024 14504 3064 14536
rect 3096 14504 3136 14536
rect 3168 14504 3208 14536
rect 3240 14504 3280 14536
rect 3312 14504 3352 14536
rect 3384 14504 3424 14536
rect 3456 14504 3496 14536
rect 3528 14504 3568 14536
rect 3600 14504 3640 14536
rect 3672 14504 3712 14536
rect 3744 14504 3784 14536
rect 3816 14504 3856 14536
rect 3888 14504 3950 14536
rect 50 14464 3950 14504
rect 50 14432 112 14464
rect 144 14432 184 14464
rect 216 14432 256 14464
rect 288 14432 328 14464
rect 360 14432 400 14464
rect 432 14432 472 14464
rect 504 14432 544 14464
rect 576 14432 616 14464
rect 648 14432 688 14464
rect 720 14432 760 14464
rect 792 14432 832 14464
rect 864 14432 904 14464
rect 936 14432 976 14464
rect 1008 14432 1048 14464
rect 1080 14432 1120 14464
rect 1152 14432 1192 14464
rect 1224 14432 1264 14464
rect 1296 14432 1336 14464
rect 1368 14432 1408 14464
rect 1440 14432 1480 14464
rect 1512 14432 1552 14464
rect 1584 14432 1624 14464
rect 1656 14432 1696 14464
rect 1728 14432 1768 14464
rect 1800 14432 1840 14464
rect 1872 14432 1912 14464
rect 1944 14432 1984 14464
rect 2016 14432 2056 14464
rect 2088 14432 2128 14464
rect 2160 14432 2200 14464
rect 2232 14432 2272 14464
rect 2304 14432 2344 14464
rect 2376 14432 2416 14464
rect 2448 14432 2488 14464
rect 2520 14432 2560 14464
rect 2592 14432 2632 14464
rect 2664 14432 2704 14464
rect 2736 14432 2776 14464
rect 2808 14432 2848 14464
rect 2880 14432 2920 14464
rect 2952 14432 2992 14464
rect 3024 14432 3064 14464
rect 3096 14432 3136 14464
rect 3168 14432 3208 14464
rect 3240 14432 3280 14464
rect 3312 14432 3352 14464
rect 3384 14432 3424 14464
rect 3456 14432 3496 14464
rect 3528 14432 3568 14464
rect 3600 14432 3640 14464
rect 3672 14432 3712 14464
rect 3744 14432 3784 14464
rect 3816 14432 3856 14464
rect 3888 14432 3950 14464
rect 50 14392 3950 14432
rect 50 14360 112 14392
rect 144 14360 184 14392
rect 216 14360 256 14392
rect 288 14360 328 14392
rect 360 14360 400 14392
rect 432 14360 472 14392
rect 504 14360 544 14392
rect 576 14360 616 14392
rect 648 14360 688 14392
rect 720 14360 760 14392
rect 792 14360 832 14392
rect 864 14360 904 14392
rect 936 14360 976 14392
rect 1008 14360 1048 14392
rect 1080 14360 1120 14392
rect 1152 14360 1192 14392
rect 1224 14360 1264 14392
rect 1296 14360 1336 14392
rect 1368 14360 1408 14392
rect 1440 14360 1480 14392
rect 1512 14360 1552 14392
rect 1584 14360 1624 14392
rect 1656 14360 1696 14392
rect 1728 14360 1768 14392
rect 1800 14360 1840 14392
rect 1872 14360 1912 14392
rect 1944 14360 1984 14392
rect 2016 14360 2056 14392
rect 2088 14360 2128 14392
rect 2160 14360 2200 14392
rect 2232 14360 2272 14392
rect 2304 14360 2344 14392
rect 2376 14360 2416 14392
rect 2448 14360 2488 14392
rect 2520 14360 2560 14392
rect 2592 14360 2632 14392
rect 2664 14360 2704 14392
rect 2736 14360 2776 14392
rect 2808 14360 2848 14392
rect 2880 14360 2920 14392
rect 2952 14360 2992 14392
rect 3024 14360 3064 14392
rect 3096 14360 3136 14392
rect 3168 14360 3208 14392
rect 3240 14360 3280 14392
rect 3312 14360 3352 14392
rect 3384 14360 3424 14392
rect 3456 14360 3496 14392
rect 3528 14360 3568 14392
rect 3600 14360 3640 14392
rect 3672 14360 3712 14392
rect 3744 14360 3784 14392
rect 3816 14360 3856 14392
rect 3888 14360 3950 14392
rect 50 14320 3950 14360
rect 50 14288 112 14320
rect 144 14288 184 14320
rect 216 14288 256 14320
rect 288 14288 328 14320
rect 360 14288 400 14320
rect 432 14288 472 14320
rect 504 14288 544 14320
rect 576 14288 616 14320
rect 648 14288 688 14320
rect 720 14288 760 14320
rect 792 14288 832 14320
rect 864 14288 904 14320
rect 936 14288 976 14320
rect 1008 14288 1048 14320
rect 1080 14288 1120 14320
rect 1152 14288 1192 14320
rect 1224 14288 1264 14320
rect 1296 14288 1336 14320
rect 1368 14288 1408 14320
rect 1440 14288 1480 14320
rect 1512 14288 1552 14320
rect 1584 14288 1624 14320
rect 1656 14288 1696 14320
rect 1728 14288 1768 14320
rect 1800 14288 1840 14320
rect 1872 14288 1912 14320
rect 1944 14288 1984 14320
rect 2016 14288 2056 14320
rect 2088 14288 2128 14320
rect 2160 14288 2200 14320
rect 2232 14288 2272 14320
rect 2304 14288 2344 14320
rect 2376 14288 2416 14320
rect 2448 14288 2488 14320
rect 2520 14288 2560 14320
rect 2592 14288 2632 14320
rect 2664 14288 2704 14320
rect 2736 14288 2776 14320
rect 2808 14288 2848 14320
rect 2880 14288 2920 14320
rect 2952 14288 2992 14320
rect 3024 14288 3064 14320
rect 3096 14288 3136 14320
rect 3168 14288 3208 14320
rect 3240 14288 3280 14320
rect 3312 14288 3352 14320
rect 3384 14288 3424 14320
rect 3456 14288 3496 14320
rect 3528 14288 3568 14320
rect 3600 14288 3640 14320
rect 3672 14288 3712 14320
rect 3744 14288 3784 14320
rect 3816 14288 3856 14320
rect 3888 14288 3950 14320
rect 50 14248 3950 14288
rect 50 14216 112 14248
rect 144 14216 184 14248
rect 216 14216 256 14248
rect 288 14216 328 14248
rect 360 14216 400 14248
rect 432 14216 472 14248
rect 504 14216 544 14248
rect 576 14216 616 14248
rect 648 14216 688 14248
rect 720 14216 760 14248
rect 792 14216 832 14248
rect 864 14216 904 14248
rect 936 14216 976 14248
rect 1008 14216 1048 14248
rect 1080 14216 1120 14248
rect 1152 14216 1192 14248
rect 1224 14216 1264 14248
rect 1296 14216 1336 14248
rect 1368 14216 1408 14248
rect 1440 14216 1480 14248
rect 1512 14216 1552 14248
rect 1584 14216 1624 14248
rect 1656 14216 1696 14248
rect 1728 14216 1768 14248
rect 1800 14216 1840 14248
rect 1872 14216 1912 14248
rect 1944 14216 1984 14248
rect 2016 14216 2056 14248
rect 2088 14216 2128 14248
rect 2160 14216 2200 14248
rect 2232 14216 2272 14248
rect 2304 14216 2344 14248
rect 2376 14216 2416 14248
rect 2448 14216 2488 14248
rect 2520 14216 2560 14248
rect 2592 14216 2632 14248
rect 2664 14216 2704 14248
rect 2736 14216 2776 14248
rect 2808 14216 2848 14248
rect 2880 14216 2920 14248
rect 2952 14216 2992 14248
rect 3024 14216 3064 14248
rect 3096 14216 3136 14248
rect 3168 14216 3208 14248
rect 3240 14216 3280 14248
rect 3312 14216 3352 14248
rect 3384 14216 3424 14248
rect 3456 14216 3496 14248
rect 3528 14216 3568 14248
rect 3600 14216 3640 14248
rect 3672 14216 3712 14248
rect 3744 14216 3784 14248
rect 3816 14216 3856 14248
rect 3888 14216 3950 14248
rect 50 14176 3950 14216
rect 50 14144 112 14176
rect 144 14144 184 14176
rect 216 14144 256 14176
rect 288 14144 328 14176
rect 360 14144 400 14176
rect 432 14144 472 14176
rect 504 14144 544 14176
rect 576 14144 616 14176
rect 648 14144 688 14176
rect 720 14144 760 14176
rect 792 14144 832 14176
rect 864 14144 904 14176
rect 936 14144 976 14176
rect 1008 14144 1048 14176
rect 1080 14144 1120 14176
rect 1152 14144 1192 14176
rect 1224 14144 1264 14176
rect 1296 14144 1336 14176
rect 1368 14144 1408 14176
rect 1440 14144 1480 14176
rect 1512 14144 1552 14176
rect 1584 14144 1624 14176
rect 1656 14144 1696 14176
rect 1728 14144 1768 14176
rect 1800 14144 1840 14176
rect 1872 14144 1912 14176
rect 1944 14144 1984 14176
rect 2016 14144 2056 14176
rect 2088 14144 2128 14176
rect 2160 14144 2200 14176
rect 2232 14144 2272 14176
rect 2304 14144 2344 14176
rect 2376 14144 2416 14176
rect 2448 14144 2488 14176
rect 2520 14144 2560 14176
rect 2592 14144 2632 14176
rect 2664 14144 2704 14176
rect 2736 14144 2776 14176
rect 2808 14144 2848 14176
rect 2880 14144 2920 14176
rect 2952 14144 2992 14176
rect 3024 14144 3064 14176
rect 3096 14144 3136 14176
rect 3168 14144 3208 14176
rect 3240 14144 3280 14176
rect 3312 14144 3352 14176
rect 3384 14144 3424 14176
rect 3456 14144 3496 14176
rect 3528 14144 3568 14176
rect 3600 14144 3640 14176
rect 3672 14144 3712 14176
rect 3744 14144 3784 14176
rect 3816 14144 3856 14176
rect 3888 14144 3950 14176
rect 50 14104 3950 14144
rect 50 14072 112 14104
rect 144 14072 184 14104
rect 216 14072 256 14104
rect 288 14072 328 14104
rect 360 14072 400 14104
rect 432 14072 472 14104
rect 504 14072 544 14104
rect 576 14072 616 14104
rect 648 14072 688 14104
rect 720 14072 760 14104
rect 792 14072 832 14104
rect 864 14072 904 14104
rect 936 14072 976 14104
rect 1008 14072 1048 14104
rect 1080 14072 1120 14104
rect 1152 14072 1192 14104
rect 1224 14072 1264 14104
rect 1296 14072 1336 14104
rect 1368 14072 1408 14104
rect 1440 14072 1480 14104
rect 1512 14072 1552 14104
rect 1584 14072 1624 14104
rect 1656 14072 1696 14104
rect 1728 14072 1768 14104
rect 1800 14072 1840 14104
rect 1872 14072 1912 14104
rect 1944 14072 1984 14104
rect 2016 14072 2056 14104
rect 2088 14072 2128 14104
rect 2160 14072 2200 14104
rect 2232 14072 2272 14104
rect 2304 14072 2344 14104
rect 2376 14072 2416 14104
rect 2448 14072 2488 14104
rect 2520 14072 2560 14104
rect 2592 14072 2632 14104
rect 2664 14072 2704 14104
rect 2736 14072 2776 14104
rect 2808 14072 2848 14104
rect 2880 14072 2920 14104
rect 2952 14072 2992 14104
rect 3024 14072 3064 14104
rect 3096 14072 3136 14104
rect 3168 14072 3208 14104
rect 3240 14072 3280 14104
rect 3312 14072 3352 14104
rect 3384 14072 3424 14104
rect 3456 14072 3496 14104
rect 3528 14072 3568 14104
rect 3600 14072 3640 14104
rect 3672 14072 3712 14104
rect 3744 14072 3784 14104
rect 3816 14072 3856 14104
rect 3888 14072 3950 14104
rect 50 14032 3950 14072
rect 50 14000 112 14032
rect 144 14000 184 14032
rect 216 14000 256 14032
rect 288 14000 328 14032
rect 360 14000 400 14032
rect 432 14000 472 14032
rect 504 14000 544 14032
rect 576 14000 616 14032
rect 648 14000 688 14032
rect 720 14000 760 14032
rect 792 14000 832 14032
rect 864 14000 904 14032
rect 936 14000 976 14032
rect 1008 14000 1048 14032
rect 1080 14000 1120 14032
rect 1152 14000 1192 14032
rect 1224 14000 1264 14032
rect 1296 14000 1336 14032
rect 1368 14000 1408 14032
rect 1440 14000 1480 14032
rect 1512 14000 1552 14032
rect 1584 14000 1624 14032
rect 1656 14000 1696 14032
rect 1728 14000 1768 14032
rect 1800 14000 1840 14032
rect 1872 14000 1912 14032
rect 1944 14000 1984 14032
rect 2016 14000 2056 14032
rect 2088 14000 2128 14032
rect 2160 14000 2200 14032
rect 2232 14000 2272 14032
rect 2304 14000 2344 14032
rect 2376 14000 2416 14032
rect 2448 14000 2488 14032
rect 2520 14000 2560 14032
rect 2592 14000 2632 14032
rect 2664 14000 2704 14032
rect 2736 14000 2776 14032
rect 2808 14000 2848 14032
rect 2880 14000 2920 14032
rect 2952 14000 2992 14032
rect 3024 14000 3064 14032
rect 3096 14000 3136 14032
rect 3168 14000 3208 14032
rect 3240 14000 3280 14032
rect 3312 14000 3352 14032
rect 3384 14000 3424 14032
rect 3456 14000 3496 14032
rect 3528 14000 3568 14032
rect 3600 14000 3640 14032
rect 3672 14000 3712 14032
rect 3744 14000 3784 14032
rect 3816 14000 3856 14032
rect 3888 14000 3950 14032
rect 50 13960 3950 14000
rect 50 13928 112 13960
rect 144 13928 184 13960
rect 216 13928 256 13960
rect 288 13928 328 13960
rect 360 13928 400 13960
rect 432 13928 472 13960
rect 504 13928 544 13960
rect 576 13928 616 13960
rect 648 13928 688 13960
rect 720 13928 760 13960
rect 792 13928 832 13960
rect 864 13928 904 13960
rect 936 13928 976 13960
rect 1008 13928 1048 13960
rect 1080 13928 1120 13960
rect 1152 13928 1192 13960
rect 1224 13928 1264 13960
rect 1296 13928 1336 13960
rect 1368 13928 1408 13960
rect 1440 13928 1480 13960
rect 1512 13928 1552 13960
rect 1584 13928 1624 13960
rect 1656 13928 1696 13960
rect 1728 13928 1768 13960
rect 1800 13928 1840 13960
rect 1872 13928 1912 13960
rect 1944 13928 1984 13960
rect 2016 13928 2056 13960
rect 2088 13928 2128 13960
rect 2160 13928 2200 13960
rect 2232 13928 2272 13960
rect 2304 13928 2344 13960
rect 2376 13928 2416 13960
rect 2448 13928 2488 13960
rect 2520 13928 2560 13960
rect 2592 13928 2632 13960
rect 2664 13928 2704 13960
rect 2736 13928 2776 13960
rect 2808 13928 2848 13960
rect 2880 13928 2920 13960
rect 2952 13928 2992 13960
rect 3024 13928 3064 13960
rect 3096 13928 3136 13960
rect 3168 13928 3208 13960
rect 3240 13928 3280 13960
rect 3312 13928 3352 13960
rect 3384 13928 3424 13960
rect 3456 13928 3496 13960
rect 3528 13928 3568 13960
rect 3600 13928 3640 13960
rect 3672 13928 3712 13960
rect 3744 13928 3784 13960
rect 3816 13928 3856 13960
rect 3888 13928 3950 13960
rect 50 13888 3950 13928
rect 50 13856 112 13888
rect 144 13856 184 13888
rect 216 13856 256 13888
rect 288 13856 328 13888
rect 360 13856 400 13888
rect 432 13856 472 13888
rect 504 13856 544 13888
rect 576 13856 616 13888
rect 648 13856 688 13888
rect 720 13856 760 13888
rect 792 13856 832 13888
rect 864 13856 904 13888
rect 936 13856 976 13888
rect 1008 13856 1048 13888
rect 1080 13856 1120 13888
rect 1152 13856 1192 13888
rect 1224 13856 1264 13888
rect 1296 13856 1336 13888
rect 1368 13856 1408 13888
rect 1440 13856 1480 13888
rect 1512 13856 1552 13888
rect 1584 13856 1624 13888
rect 1656 13856 1696 13888
rect 1728 13856 1768 13888
rect 1800 13856 1840 13888
rect 1872 13856 1912 13888
rect 1944 13856 1984 13888
rect 2016 13856 2056 13888
rect 2088 13856 2128 13888
rect 2160 13856 2200 13888
rect 2232 13856 2272 13888
rect 2304 13856 2344 13888
rect 2376 13856 2416 13888
rect 2448 13856 2488 13888
rect 2520 13856 2560 13888
rect 2592 13856 2632 13888
rect 2664 13856 2704 13888
rect 2736 13856 2776 13888
rect 2808 13856 2848 13888
rect 2880 13856 2920 13888
rect 2952 13856 2992 13888
rect 3024 13856 3064 13888
rect 3096 13856 3136 13888
rect 3168 13856 3208 13888
rect 3240 13856 3280 13888
rect 3312 13856 3352 13888
rect 3384 13856 3424 13888
rect 3456 13856 3496 13888
rect 3528 13856 3568 13888
rect 3600 13856 3640 13888
rect 3672 13856 3712 13888
rect 3744 13856 3784 13888
rect 3816 13856 3856 13888
rect 3888 13856 3950 13888
rect 50 13816 3950 13856
rect 50 13784 112 13816
rect 144 13784 184 13816
rect 216 13784 256 13816
rect 288 13784 328 13816
rect 360 13784 400 13816
rect 432 13784 472 13816
rect 504 13784 544 13816
rect 576 13784 616 13816
rect 648 13784 688 13816
rect 720 13784 760 13816
rect 792 13784 832 13816
rect 864 13784 904 13816
rect 936 13784 976 13816
rect 1008 13784 1048 13816
rect 1080 13784 1120 13816
rect 1152 13784 1192 13816
rect 1224 13784 1264 13816
rect 1296 13784 1336 13816
rect 1368 13784 1408 13816
rect 1440 13784 1480 13816
rect 1512 13784 1552 13816
rect 1584 13784 1624 13816
rect 1656 13784 1696 13816
rect 1728 13784 1768 13816
rect 1800 13784 1840 13816
rect 1872 13784 1912 13816
rect 1944 13784 1984 13816
rect 2016 13784 2056 13816
rect 2088 13784 2128 13816
rect 2160 13784 2200 13816
rect 2232 13784 2272 13816
rect 2304 13784 2344 13816
rect 2376 13784 2416 13816
rect 2448 13784 2488 13816
rect 2520 13784 2560 13816
rect 2592 13784 2632 13816
rect 2664 13784 2704 13816
rect 2736 13784 2776 13816
rect 2808 13784 2848 13816
rect 2880 13784 2920 13816
rect 2952 13784 2992 13816
rect 3024 13784 3064 13816
rect 3096 13784 3136 13816
rect 3168 13784 3208 13816
rect 3240 13784 3280 13816
rect 3312 13784 3352 13816
rect 3384 13784 3424 13816
rect 3456 13784 3496 13816
rect 3528 13784 3568 13816
rect 3600 13784 3640 13816
rect 3672 13784 3712 13816
rect 3744 13784 3784 13816
rect 3816 13784 3856 13816
rect 3888 13784 3950 13816
rect 50 13744 3950 13784
rect 50 13712 112 13744
rect 144 13712 184 13744
rect 216 13712 256 13744
rect 288 13712 328 13744
rect 360 13712 400 13744
rect 432 13712 472 13744
rect 504 13712 544 13744
rect 576 13712 616 13744
rect 648 13712 688 13744
rect 720 13712 760 13744
rect 792 13712 832 13744
rect 864 13712 904 13744
rect 936 13712 976 13744
rect 1008 13712 1048 13744
rect 1080 13712 1120 13744
rect 1152 13712 1192 13744
rect 1224 13712 1264 13744
rect 1296 13712 1336 13744
rect 1368 13712 1408 13744
rect 1440 13712 1480 13744
rect 1512 13712 1552 13744
rect 1584 13712 1624 13744
rect 1656 13712 1696 13744
rect 1728 13712 1768 13744
rect 1800 13712 1840 13744
rect 1872 13712 1912 13744
rect 1944 13712 1984 13744
rect 2016 13712 2056 13744
rect 2088 13712 2128 13744
rect 2160 13712 2200 13744
rect 2232 13712 2272 13744
rect 2304 13712 2344 13744
rect 2376 13712 2416 13744
rect 2448 13712 2488 13744
rect 2520 13712 2560 13744
rect 2592 13712 2632 13744
rect 2664 13712 2704 13744
rect 2736 13712 2776 13744
rect 2808 13712 2848 13744
rect 2880 13712 2920 13744
rect 2952 13712 2992 13744
rect 3024 13712 3064 13744
rect 3096 13712 3136 13744
rect 3168 13712 3208 13744
rect 3240 13712 3280 13744
rect 3312 13712 3352 13744
rect 3384 13712 3424 13744
rect 3456 13712 3496 13744
rect 3528 13712 3568 13744
rect 3600 13712 3640 13744
rect 3672 13712 3712 13744
rect 3744 13712 3784 13744
rect 3816 13712 3856 13744
rect 3888 13712 3950 13744
rect 50 13672 3950 13712
rect 50 13640 112 13672
rect 144 13640 184 13672
rect 216 13640 256 13672
rect 288 13640 328 13672
rect 360 13640 400 13672
rect 432 13640 472 13672
rect 504 13640 544 13672
rect 576 13640 616 13672
rect 648 13640 688 13672
rect 720 13640 760 13672
rect 792 13640 832 13672
rect 864 13640 904 13672
rect 936 13640 976 13672
rect 1008 13640 1048 13672
rect 1080 13640 1120 13672
rect 1152 13640 1192 13672
rect 1224 13640 1264 13672
rect 1296 13640 1336 13672
rect 1368 13640 1408 13672
rect 1440 13640 1480 13672
rect 1512 13640 1552 13672
rect 1584 13640 1624 13672
rect 1656 13640 1696 13672
rect 1728 13640 1768 13672
rect 1800 13640 1840 13672
rect 1872 13640 1912 13672
rect 1944 13640 1984 13672
rect 2016 13640 2056 13672
rect 2088 13640 2128 13672
rect 2160 13640 2200 13672
rect 2232 13640 2272 13672
rect 2304 13640 2344 13672
rect 2376 13640 2416 13672
rect 2448 13640 2488 13672
rect 2520 13640 2560 13672
rect 2592 13640 2632 13672
rect 2664 13640 2704 13672
rect 2736 13640 2776 13672
rect 2808 13640 2848 13672
rect 2880 13640 2920 13672
rect 2952 13640 2992 13672
rect 3024 13640 3064 13672
rect 3096 13640 3136 13672
rect 3168 13640 3208 13672
rect 3240 13640 3280 13672
rect 3312 13640 3352 13672
rect 3384 13640 3424 13672
rect 3456 13640 3496 13672
rect 3528 13640 3568 13672
rect 3600 13640 3640 13672
rect 3672 13640 3712 13672
rect 3744 13640 3784 13672
rect 3816 13640 3856 13672
rect 3888 13640 3950 13672
rect 50 13600 3950 13640
rect 50 13568 112 13600
rect 144 13568 184 13600
rect 216 13568 256 13600
rect 288 13568 328 13600
rect 360 13568 400 13600
rect 432 13568 472 13600
rect 504 13568 544 13600
rect 576 13568 616 13600
rect 648 13568 688 13600
rect 720 13568 760 13600
rect 792 13568 832 13600
rect 864 13568 904 13600
rect 936 13568 976 13600
rect 1008 13568 1048 13600
rect 1080 13568 1120 13600
rect 1152 13568 1192 13600
rect 1224 13568 1264 13600
rect 1296 13568 1336 13600
rect 1368 13568 1408 13600
rect 1440 13568 1480 13600
rect 1512 13568 1552 13600
rect 1584 13568 1624 13600
rect 1656 13568 1696 13600
rect 1728 13568 1768 13600
rect 1800 13568 1840 13600
rect 1872 13568 1912 13600
rect 1944 13568 1984 13600
rect 2016 13568 2056 13600
rect 2088 13568 2128 13600
rect 2160 13568 2200 13600
rect 2232 13568 2272 13600
rect 2304 13568 2344 13600
rect 2376 13568 2416 13600
rect 2448 13568 2488 13600
rect 2520 13568 2560 13600
rect 2592 13568 2632 13600
rect 2664 13568 2704 13600
rect 2736 13568 2776 13600
rect 2808 13568 2848 13600
rect 2880 13568 2920 13600
rect 2952 13568 2992 13600
rect 3024 13568 3064 13600
rect 3096 13568 3136 13600
rect 3168 13568 3208 13600
rect 3240 13568 3280 13600
rect 3312 13568 3352 13600
rect 3384 13568 3424 13600
rect 3456 13568 3496 13600
rect 3528 13568 3568 13600
rect 3600 13568 3640 13600
rect 3672 13568 3712 13600
rect 3744 13568 3784 13600
rect 3816 13568 3856 13600
rect 3888 13568 3950 13600
rect 50 13528 3950 13568
rect 50 13496 112 13528
rect 144 13496 184 13528
rect 216 13496 256 13528
rect 288 13496 328 13528
rect 360 13496 400 13528
rect 432 13496 472 13528
rect 504 13496 544 13528
rect 576 13496 616 13528
rect 648 13496 688 13528
rect 720 13496 760 13528
rect 792 13496 832 13528
rect 864 13496 904 13528
rect 936 13496 976 13528
rect 1008 13496 1048 13528
rect 1080 13496 1120 13528
rect 1152 13496 1192 13528
rect 1224 13496 1264 13528
rect 1296 13496 1336 13528
rect 1368 13496 1408 13528
rect 1440 13496 1480 13528
rect 1512 13496 1552 13528
rect 1584 13496 1624 13528
rect 1656 13496 1696 13528
rect 1728 13496 1768 13528
rect 1800 13496 1840 13528
rect 1872 13496 1912 13528
rect 1944 13496 1984 13528
rect 2016 13496 2056 13528
rect 2088 13496 2128 13528
rect 2160 13496 2200 13528
rect 2232 13496 2272 13528
rect 2304 13496 2344 13528
rect 2376 13496 2416 13528
rect 2448 13496 2488 13528
rect 2520 13496 2560 13528
rect 2592 13496 2632 13528
rect 2664 13496 2704 13528
rect 2736 13496 2776 13528
rect 2808 13496 2848 13528
rect 2880 13496 2920 13528
rect 2952 13496 2992 13528
rect 3024 13496 3064 13528
rect 3096 13496 3136 13528
rect 3168 13496 3208 13528
rect 3240 13496 3280 13528
rect 3312 13496 3352 13528
rect 3384 13496 3424 13528
rect 3456 13496 3496 13528
rect 3528 13496 3568 13528
rect 3600 13496 3640 13528
rect 3672 13496 3712 13528
rect 3744 13496 3784 13528
rect 3816 13496 3856 13528
rect 3888 13496 3950 13528
rect 50 13456 3950 13496
rect 50 13424 112 13456
rect 144 13424 184 13456
rect 216 13424 256 13456
rect 288 13424 328 13456
rect 360 13424 400 13456
rect 432 13424 472 13456
rect 504 13424 544 13456
rect 576 13424 616 13456
rect 648 13424 688 13456
rect 720 13424 760 13456
rect 792 13424 832 13456
rect 864 13424 904 13456
rect 936 13424 976 13456
rect 1008 13424 1048 13456
rect 1080 13424 1120 13456
rect 1152 13424 1192 13456
rect 1224 13424 1264 13456
rect 1296 13424 1336 13456
rect 1368 13424 1408 13456
rect 1440 13424 1480 13456
rect 1512 13424 1552 13456
rect 1584 13424 1624 13456
rect 1656 13424 1696 13456
rect 1728 13424 1768 13456
rect 1800 13424 1840 13456
rect 1872 13424 1912 13456
rect 1944 13424 1984 13456
rect 2016 13424 2056 13456
rect 2088 13424 2128 13456
rect 2160 13424 2200 13456
rect 2232 13424 2272 13456
rect 2304 13424 2344 13456
rect 2376 13424 2416 13456
rect 2448 13424 2488 13456
rect 2520 13424 2560 13456
rect 2592 13424 2632 13456
rect 2664 13424 2704 13456
rect 2736 13424 2776 13456
rect 2808 13424 2848 13456
rect 2880 13424 2920 13456
rect 2952 13424 2992 13456
rect 3024 13424 3064 13456
rect 3096 13424 3136 13456
rect 3168 13424 3208 13456
rect 3240 13424 3280 13456
rect 3312 13424 3352 13456
rect 3384 13424 3424 13456
rect 3456 13424 3496 13456
rect 3528 13424 3568 13456
rect 3600 13424 3640 13456
rect 3672 13424 3712 13456
rect 3744 13424 3784 13456
rect 3816 13424 3856 13456
rect 3888 13424 3950 13456
rect 50 13384 3950 13424
rect 50 13352 112 13384
rect 144 13352 184 13384
rect 216 13352 256 13384
rect 288 13352 328 13384
rect 360 13352 400 13384
rect 432 13352 472 13384
rect 504 13352 544 13384
rect 576 13352 616 13384
rect 648 13352 688 13384
rect 720 13352 760 13384
rect 792 13352 832 13384
rect 864 13352 904 13384
rect 936 13352 976 13384
rect 1008 13352 1048 13384
rect 1080 13352 1120 13384
rect 1152 13352 1192 13384
rect 1224 13352 1264 13384
rect 1296 13352 1336 13384
rect 1368 13352 1408 13384
rect 1440 13352 1480 13384
rect 1512 13352 1552 13384
rect 1584 13352 1624 13384
rect 1656 13352 1696 13384
rect 1728 13352 1768 13384
rect 1800 13352 1840 13384
rect 1872 13352 1912 13384
rect 1944 13352 1984 13384
rect 2016 13352 2056 13384
rect 2088 13352 2128 13384
rect 2160 13352 2200 13384
rect 2232 13352 2272 13384
rect 2304 13352 2344 13384
rect 2376 13352 2416 13384
rect 2448 13352 2488 13384
rect 2520 13352 2560 13384
rect 2592 13352 2632 13384
rect 2664 13352 2704 13384
rect 2736 13352 2776 13384
rect 2808 13352 2848 13384
rect 2880 13352 2920 13384
rect 2952 13352 2992 13384
rect 3024 13352 3064 13384
rect 3096 13352 3136 13384
rect 3168 13352 3208 13384
rect 3240 13352 3280 13384
rect 3312 13352 3352 13384
rect 3384 13352 3424 13384
rect 3456 13352 3496 13384
rect 3528 13352 3568 13384
rect 3600 13352 3640 13384
rect 3672 13352 3712 13384
rect 3744 13352 3784 13384
rect 3816 13352 3856 13384
rect 3888 13352 3950 13384
rect 50 13312 3950 13352
rect 50 13280 112 13312
rect 144 13280 184 13312
rect 216 13280 256 13312
rect 288 13280 328 13312
rect 360 13280 400 13312
rect 432 13280 472 13312
rect 504 13280 544 13312
rect 576 13280 616 13312
rect 648 13280 688 13312
rect 720 13280 760 13312
rect 792 13280 832 13312
rect 864 13280 904 13312
rect 936 13280 976 13312
rect 1008 13280 1048 13312
rect 1080 13280 1120 13312
rect 1152 13280 1192 13312
rect 1224 13280 1264 13312
rect 1296 13280 1336 13312
rect 1368 13280 1408 13312
rect 1440 13280 1480 13312
rect 1512 13280 1552 13312
rect 1584 13280 1624 13312
rect 1656 13280 1696 13312
rect 1728 13280 1768 13312
rect 1800 13280 1840 13312
rect 1872 13280 1912 13312
rect 1944 13280 1984 13312
rect 2016 13280 2056 13312
rect 2088 13280 2128 13312
rect 2160 13280 2200 13312
rect 2232 13280 2272 13312
rect 2304 13280 2344 13312
rect 2376 13280 2416 13312
rect 2448 13280 2488 13312
rect 2520 13280 2560 13312
rect 2592 13280 2632 13312
rect 2664 13280 2704 13312
rect 2736 13280 2776 13312
rect 2808 13280 2848 13312
rect 2880 13280 2920 13312
rect 2952 13280 2992 13312
rect 3024 13280 3064 13312
rect 3096 13280 3136 13312
rect 3168 13280 3208 13312
rect 3240 13280 3280 13312
rect 3312 13280 3352 13312
rect 3384 13280 3424 13312
rect 3456 13280 3496 13312
rect 3528 13280 3568 13312
rect 3600 13280 3640 13312
rect 3672 13280 3712 13312
rect 3744 13280 3784 13312
rect 3816 13280 3856 13312
rect 3888 13280 3950 13312
rect 50 13240 3950 13280
rect 50 13208 112 13240
rect 144 13208 184 13240
rect 216 13208 256 13240
rect 288 13208 328 13240
rect 360 13208 400 13240
rect 432 13208 472 13240
rect 504 13208 544 13240
rect 576 13208 616 13240
rect 648 13208 688 13240
rect 720 13208 760 13240
rect 792 13208 832 13240
rect 864 13208 904 13240
rect 936 13208 976 13240
rect 1008 13208 1048 13240
rect 1080 13208 1120 13240
rect 1152 13208 1192 13240
rect 1224 13208 1264 13240
rect 1296 13208 1336 13240
rect 1368 13208 1408 13240
rect 1440 13208 1480 13240
rect 1512 13208 1552 13240
rect 1584 13208 1624 13240
rect 1656 13208 1696 13240
rect 1728 13208 1768 13240
rect 1800 13208 1840 13240
rect 1872 13208 1912 13240
rect 1944 13208 1984 13240
rect 2016 13208 2056 13240
rect 2088 13208 2128 13240
rect 2160 13208 2200 13240
rect 2232 13208 2272 13240
rect 2304 13208 2344 13240
rect 2376 13208 2416 13240
rect 2448 13208 2488 13240
rect 2520 13208 2560 13240
rect 2592 13208 2632 13240
rect 2664 13208 2704 13240
rect 2736 13208 2776 13240
rect 2808 13208 2848 13240
rect 2880 13208 2920 13240
rect 2952 13208 2992 13240
rect 3024 13208 3064 13240
rect 3096 13208 3136 13240
rect 3168 13208 3208 13240
rect 3240 13208 3280 13240
rect 3312 13208 3352 13240
rect 3384 13208 3424 13240
rect 3456 13208 3496 13240
rect 3528 13208 3568 13240
rect 3600 13208 3640 13240
rect 3672 13208 3712 13240
rect 3744 13208 3784 13240
rect 3816 13208 3856 13240
rect 3888 13208 3950 13240
rect 50 13168 3950 13208
rect 50 13136 112 13168
rect 144 13136 184 13168
rect 216 13136 256 13168
rect 288 13136 328 13168
rect 360 13136 400 13168
rect 432 13136 472 13168
rect 504 13136 544 13168
rect 576 13136 616 13168
rect 648 13136 688 13168
rect 720 13136 760 13168
rect 792 13136 832 13168
rect 864 13136 904 13168
rect 936 13136 976 13168
rect 1008 13136 1048 13168
rect 1080 13136 1120 13168
rect 1152 13136 1192 13168
rect 1224 13136 1264 13168
rect 1296 13136 1336 13168
rect 1368 13136 1408 13168
rect 1440 13136 1480 13168
rect 1512 13136 1552 13168
rect 1584 13136 1624 13168
rect 1656 13136 1696 13168
rect 1728 13136 1768 13168
rect 1800 13136 1840 13168
rect 1872 13136 1912 13168
rect 1944 13136 1984 13168
rect 2016 13136 2056 13168
rect 2088 13136 2128 13168
rect 2160 13136 2200 13168
rect 2232 13136 2272 13168
rect 2304 13136 2344 13168
rect 2376 13136 2416 13168
rect 2448 13136 2488 13168
rect 2520 13136 2560 13168
rect 2592 13136 2632 13168
rect 2664 13136 2704 13168
rect 2736 13136 2776 13168
rect 2808 13136 2848 13168
rect 2880 13136 2920 13168
rect 2952 13136 2992 13168
rect 3024 13136 3064 13168
rect 3096 13136 3136 13168
rect 3168 13136 3208 13168
rect 3240 13136 3280 13168
rect 3312 13136 3352 13168
rect 3384 13136 3424 13168
rect 3456 13136 3496 13168
rect 3528 13136 3568 13168
rect 3600 13136 3640 13168
rect 3672 13136 3712 13168
rect 3744 13136 3784 13168
rect 3816 13136 3856 13168
rect 3888 13136 3950 13168
rect 50 13096 3950 13136
rect 50 13064 112 13096
rect 144 13064 184 13096
rect 216 13064 256 13096
rect 288 13064 328 13096
rect 360 13064 400 13096
rect 432 13064 472 13096
rect 504 13064 544 13096
rect 576 13064 616 13096
rect 648 13064 688 13096
rect 720 13064 760 13096
rect 792 13064 832 13096
rect 864 13064 904 13096
rect 936 13064 976 13096
rect 1008 13064 1048 13096
rect 1080 13064 1120 13096
rect 1152 13064 1192 13096
rect 1224 13064 1264 13096
rect 1296 13064 1336 13096
rect 1368 13064 1408 13096
rect 1440 13064 1480 13096
rect 1512 13064 1552 13096
rect 1584 13064 1624 13096
rect 1656 13064 1696 13096
rect 1728 13064 1768 13096
rect 1800 13064 1840 13096
rect 1872 13064 1912 13096
rect 1944 13064 1984 13096
rect 2016 13064 2056 13096
rect 2088 13064 2128 13096
rect 2160 13064 2200 13096
rect 2232 13064 2272 13096
rect 2304 13064 2344 13096
rect 2376 13064 2416 13096
rect 2448 13064 2488 13096
rect 2520 13064 2560 13096
rect 2592 13064 2632 13096
rect 2664 13064 2704 13096
rect 2736 13064 2776 13096
rect 2808 13064 2848 13096
rect 2880 13064 2920 13096
rect 2952 13064 2992 13096
rect 3024 13064 3064 13096
rect 3096 13064 3136 13096
rect 3168 13064 3208 13096
rect 3240 13064 3280 13096
rect 3312 13064 3352 13096
rect 3384 13064 3424 13096
rect 3456 13064 3496 13096
rect 3528 13064 3568 13096
rect 3600 13064 3640 13096
rect 3672 13064 3712 13096
rect 3744 13064 3784 13096
rect 3816 13064 3856 13096
rect 3888 13064 3950 13096
rect 50 13000 3950 13064
<< nsubdiff >>
rect 184 33384 216 33416
rect 256 33384 288 33416
rect 328 33384 360 33416
rect 400 33384 432 33416
rect 472 33384 504 33416
rect 544 33384 576 33416
rect 616 33384 648 33416
rect 688 33384 720 33416
rect 760 33384 792 33416
rect 832 33384 864 33416
rect 904 33384 936 33416
rect 976 33384 1008 33416
rect 1048 33384 1080 33416
rect 1120 33384 1152 33416
rect 1192 33384 1224 33416
rect 1264 33384 1296 33416
rect 1336 33384 1368 33416
rect 1408 33384 1440 33416
rect 1480 33384 1512 33416
rect 1552 33384 1584 33416
rect 1624 33384 1656 33416
rect 1696 33384 1728 33416
rect 1768 33384 1800 33416
rect 1840 33384 1872 33416
rect 1912 33384 1944 33416
rect 1984 33384 2016 33416
rect 2056 33384 2088 33416
rect 2128 33384 2160 33416
rect 2200 33384 2232 33416
rect 2272 33384 2304 33416
rect 2344 33384 2376 33416
rect 2416 33384 2448 33416
rect 2488 33384 2520 33416
rect 2560 33384 2592 33416
rect 2632 33384 2664 33416
rect 2704 33384 2736 33416
rect 2776 33384 2808 33416
rect 2848 33384 2880 33416
rect 2920 33384 2952 33416
rect 2992 33384 3024 33416
rect 3064 33384 3096 33416
rect 3136 33384 3168 33416
rect 3208 33384 3240 33416
rect 3280 33384 3312 33416
rect 3352 33384 3384 33416
rect 3424 33384 3456 33416
rect 3496 33384 3528 33416
rect 3568 33384 3600 33416
rect 3640 33384 3672 33416
rect 3712 33384 3744 33416
rect 3784 33384 3816 33416
rect 3856 33384 3888 33416
rect 184 29684 216 29716
rect 256 29684 288 29716
rect 328 29684 360 29716
rect 400 29684 432 29716
rect 472 29684 504 29716
rect 544 29684 576 29716
rect 616 29684 648 29716
rect 688 29684 720 29716
rect 760 29684 792 29716
rect 832 29684 864 29716
rect 904 29684 936 29716
rect 976 29684 1008 29716
rect 1048 29684 1080 29716
rect 1120 29684 1152 29716
rect 1192 29684 1224 29716
rect 1264 29684 1296 29716
rect 1336 29684 1368 29716
rect 1408 29684 1440 29716
rect 1480 29684 1512 29716
rect 1552 29684 1584 29716
rect 1624 29684 1656 29716
rect 1696 29684 1728 29716
rect 1768 29684 1800 29716
rect 1840 29684 1872 29716
rect 1912 29684 1944 29716
rect 1984 29684 2016 29716
rect 2056 29684 2088 29716
rect 2128 29684 2160 29716
rect 2200 29684 2232 29716
rect 2272 29684 2304 29716
rect 2344 29684 2376 29716
rect 2416 29684 2448 29716
rect 2488 29684 2520 29716
rect 2560 29684 2592 29716
rect 2632 29684 2664 29716
rect 2704 29684 2736 29716
rect 2776 29684 2808 29716
rect 2848 29684 2880 29716
rect 2920 29684 2952 29716
rect 2992 29684 3024 29716
rect 3064 29684 3096 29716
rect 3136 29684 3168 29716
rect 3208 29684 3240 29716
rect 3280 29684 3312 29716
rect 3352 29684 3384 29716
rect 3424 29684 3456 29716
rect 3496 29684 3528 29716
rect 3568 29684 3600 29716
rect 3640 29684 3672 29716
rect 3712 29684 3744 29716
rect 3784 29684 3816 29716
rect 3856 29684 3888 29716
rect 112 12112 144 12144
rect 184 12112 216 12144
rect 256 12112 288 12144
rect 328 12112 360 12144
rect 400 12112 432 12144
rect 472 12112 504 12144
rect 544 12112 576 12144
rect 616 12112 648 12144
rect 688 12112 720 12144
rect 760 12112 792 12144
rect 832 12112 864 12144
rect 904 12112 936 12144
rect 976 12112 1008 12144
rect 1048 12112 1080 12144
rect 1120 12112 1152 12144
rect 1192 12112 1224 12144
rect 1264 12112 1296 12144
rect 1336 12112 1368 12144
rect 1408 12112 1440 12144
rect 1480 12112 1512 12144
rect 1552 12112 1584 12144
rect 1624 12112 1656 12144
rect 1696 12112 1728 12144
rect 1768 12112 1800 12144
rect 1840 12112 1872 12144
rect 1912 12112 1944 12144
rect 1984 12112 2016 12144
rect 2056 12112 2088 12144
rect 2128 12112 2160 12144
rect 2200 12112 2232 12144
rect 2272 12112 2304 12144
rect 2344 12112 2376 12144
rect 2416 12112 2448 12144
rect 2488 12112 2520 12144
rect 2560 12112 2592 12144
rect 2632 12112 2664 12144
rect 2704 12112 2736 12144
rect 2776 12112 2808 12144
rect 2848 12112 2880 12144
rect 2920 12112 2952 12144
rect 2992 12112 3024 12144
rect 3064 12112 3096 12144
rect 3136 12112 3168 12144
rect 3208 12112 3240 12144
rect 3280 12112 3312 12144
rect 3352 12112 3384 12144
rect 3424 12112 3456 12144
rect 3496 12112 3528 12144
rect 3568 12112 3600 12144
rect 3640 12112 3672 12144
rect 3712 12112 3744 12144
rect 3784 12112 3816 12144
rect 3856 12112 3888 12144
rect 3928 12112 3960 12144
rect 40 12040 72 12072
rect 112 12040 144 12072
rect 184 12040 216 12072
rect 256 12040 288 12072
rect 328 12040 360 12072
rect 400 12040 432 12072
rect 472 12040 504 12072
rect 544 12040 576 12072
rect 616 12040 648 12072
rect 688 12040 720 12072
rect 760 12040 792 12072
rect 832 12040 864 12072
rect 904 12040 936 12072
rect 976 12040 1008 12072
rect 1048 12040 1080 12072
rect 1120 12040 1152 12072
rect 1192 12040 1224 12072
rect 1264 12040 1296 12072
rect 1336 12040 1368 12072
rect 1408 12040 1440 12072
rect 1480 12040 1512 12072
rect 1552 12040 1584 12072
rect 1624 12040 1656 12072
rect 1696 12040 1728 12072
rect 1768 12040 1800 12072
rect 1840 12040 1872 12072
rect 1912 12040 1944 12072
rect 1984 12040 2016 12072
rect 2056 12040 2088 12072
rect 2128 12040 2160 12072
rect 2200 12040 2232 12072
rect 2272 12040 2304 12072
rect 2344 12040 2376 12072
rect 2416 12040 2448 12072
rect 2488 12040 2520 12072
rect 2560 12040 2592 12072
rect 2632 12040 2664 12072
rect 2704 12040 2736 12072
rect 2776 12040 2808 12072
rect 2848 12040 2880 12072
rect 2920 12040 2952 12072
rect 2992 12040 3024 12072
rect 3064 12040 3096 12072
rect 3136 12040 3168 12072
rect 3208 12040 3240 12072
rect 3280 12040 3312 12072
rect 3352 12040 3384 12072
rect 3424 12040 3456 12072
rect 3496 12040 3528 12072
rect 3568 12040 3600 12072
rect 3640 12040 3672 12072
rect 3712 12040 3744 12072
rect 3784 12040 3816 12072
rect 3856 12040 3888 12072
rect 3928 12040 3960 12072
rect 40 11968 72 12000
rect 112 11968 144 12000
rect 184 11968 216 12000
rect 256 11968 288 12000
rect 328 11968 360 12000
rect 400 11968 432 12000
rect 472 11968 504 12000
rect 544 11968 576 12000
rect 616 11968 648 12000
rect 688 11968 720 12000
rect 760 11968 792 12000
rect 832 11968 864 12000
rect 904 11968 936 12000
rect 976 11968 1008 12000
rect 1048 11968 1080 12000
rect 1120 11968 1152 12000
rect 1192 11968 1224 12000
rect 1264 11968 1296 12000
rect 1336 11968 1368 12000
rect 1408 11968 1440 12000
rect 1480 11968 1512 12000
rect 1552 11968 1584 12000
rect 1624 11968 1656 12000
rect 1696 11968 1728 12000
rect 1768 11968 1800 12000
rect 1840 11968 1872 12000
rect 1912 11968 1944 12000
rect 1984 11968 2016 12000
rect 2056 11968 2088 12000
rect 2128 11968 2160 12000
rect 2200 11968 2232 12000
rect 2272 11968 2304 12000
rect 2344 11968 2376 12000
rect 2416 11968 2448 12000
rect 2488 11968 2520 12000
rect 2560 11968 2592 12000
rect 2632 11968 2664 12000
rect 2704 11968 2736 12000
rect 2776 11968 2808 12000
rect 2848 11968 2880 12000
rect 2920 11968 2952 12000
rect 2992 11968 3024 12000
rect 3064 11968 3096 12000
rect 3136 11968 3168 12000
rect 3208 11968 3240 12000
rect 3280 11968 3312 12000
rect 3352 11968 3384 12000
rect 3424 11968 3456 12000
rect 3496 11968 3528 12000
rect 3568 11968 3600 12000
rect 3640 11968 3672 12000
rect 3712 11968 3744 12000
rect 3784 11968 3816 12000
rect 3856 11968 3888 12000
rect 3928 11968 3960 12000
rect 40 11896 72 11928
rect 112 11896 144 11928
rect 184 11896 216 11928
rect 256 11896 288 11928
rect 328 11896 360 11928
rect 400 11896 432 11928
rect 472 11896 504 11928
rect 544 11896 576 11928
rect 616 11896 648 11928
rect 688 11896 720 11928
rect 760 11896 792 11928
rect 832 11896 864 11928
rect 904 11896 936 11928
rect 976 11896 1008 11928
rect 1048 11896 1080 11928
rect 1120 11896 1152 11928
rect 1192 11896 1224 11928
rect 1264 11896 1296 11928
rect 1336 11896 1368 11928
rect 1408 11896 1440 11928
rect 1480 11896 1512 11928
rect 1552 11896 1584 11928
rect 1624 11896 1656 11928
rect 1696 11896 1728 11928
rect 1768 11896 1800 11928
rect 1840 11896 1872 11928
rect 1912 11896 1944 11928
rect 1984 11896 2016 11928
rect 2056 11896 2088 11928
rect 2128 11896 2160 11928
rect 2200 11896 2232 11928
rect 2272 11896 2304 11928
rect 2344 11896 2376 11928
rect 2416 11896 2448 11928
rect 2488 11896 2520 11928
rect 2560 11896 2592 11928
rect 2632 11896 2664 11928
rect 2704 11896 2736 11928
rect 2776 11896 2808 11928
rect 2848 11896 2880 11928
rect 2920 11896 2952 11928
rect 2992 11896 3024 11928
rect 3064 11896 3096 11928
rect 3136 11896 3168 11928
rect 3208 11896 3240 11928
rect 3280 11896 3312 11928
rect 3352 11896 3384 11928
rect 3424 11896 3456 11928
rect 3496 11896 3528 11928
rect 3568 11896 3600 11928
rect 3640 11896 3672 11928
rect 3712 11896 3744 11928
rect 3784 11896 3816 11928
rect 3856 11896 3888 11928
rect 3928 11896 3960 11928
rect 40 11824 72 11856
rect 112 11824 144 11856
rect 184 11824 216 11856
rect 256 11824 288 11856
rect 328 11824 360 11856
rect 400 11824 432 11856
rect 472 11824 504 11856
rect 544 11824 576 11856
rect 616 11824 648 11856
rect 688 11824 720 11856
rect 760 11824 792 11856
rect 832 11824 864 11856
rect 904 11824 936 11856
rect 976 11824 1008 11856
rect 1048 11824 1080 11856
rect 1120 11824 1152 11856
rect 1192 11824 1224 11856
rect 1264 11824 1296 11856
rect 1336 11824 1368 11856
rect 1408 11824 1440 11856
rect 1480 11824 1512 11856
rect 1552 11824 1584 11856
rect 1624 11824 1656 11856
rect 1696 11824 1728 11856
rect 1768 11824 1800 11856
rect 1840 11824 1872 11856
rect 1912 11824 1944 11856
rect 1984 11824 2016 11856
rect 2056 11824 2088 11856
rect 2128 11824 2160 11856
rect 2200 11824 2232 11856
rect 2272 11824 2304 11856
rect 2344 11824 2376 11856
rect 2416 11824 2448 11856
rect 2488 11824 2520 11856
rect 2560 11824 2592 11856
rect 2632 11824 2664 11856
rect 2704 11824 2736 11856
rect 2776 11824 2808 11856
rect 2848 11824 2880 11856
rect 2920 11824 2952 11856
rect 2992 11824 3024 11856
rect 3064 11824 3096 11856
rect 3136 11824 3168 11856
rect 3208 11824 3240 11856
rect 3280 11824 3312 11856
rect 3352 11824 3384 11856
rect 3424 11824 3456 11856
rect 3496 11824 3528 11856
rect 3568 11824 3600 11856
rect 3640 11824 3672 11856
rect 3712 11824 3744 11856
rect 3784 11824 3816 11856
rect 3856 11824 3888 11856
rect 3928 11824 3960 11856
rect 40 11752 72 11784
rect 112 11752 144 11784
rect 184 11752 216 11784
rect 256 11752 288 11784
rect 328 11752 360 11784
rect 400 11752 432 11784
rect 472 11752 504 11784
rect 544 11752 576 11784
rect 616 11752 648 11784
rect 688 11752 720 11784
rect 760 11752 792 11784
rect 832 11752 864 11784
rect 904 11752 936 11784
rect 976 11752 1008 11784
rect 1048 11752 1080 11784
rect 1120 11752 1152 11784
rect 1192 11752 1224 11784
rect 1264 11752 1296 11784
rect 1336 11752 1368 11784
rect 1408 11752 1440 11784
rect 1480 11752 1512 11784
rect 1552 11752 1584 11784
rect 1624 11752 1656 11784
rect 1696 11752 1728 11784
rect 1768 11752 1800 11784
rect 1840 11752 1872 11784
rect 1912 11752 1944 11784
rect 1984 11752 2016 11784
rect 2056 11752 2088 11784
rect 2128 11752 2160 11784
rect 2200 11752 2232 11784
rect 2272 11752 2304 11784
rect 2344 11752 2376 11784
rect 2416 11752 2448 11784
rect 2488 11752 2520 11784
rect 2560 11752 2592 11784
rect 2632 11752 2664 11784
rect 2704 11752 2736 11784
rect 2776 11752 2808 11784
rect 2848 11752 2880 11784
rect 2920 11752 2952 11784
rect 2992 11752 3024 11784
rect 3064 11752 3096 11784
rect 3136 11752 3168 11784
rect 3208 11752 3240 11784
rect 3280 11752 3312 11784
rect 3352 11752 3384 11784
rect 3424 11752 3456 11784
rect 3496 11752 3528 11784
rect 3568 11752 3600 11784
rect 3640 11752 3672 11784
rect 3712 11752 3744 11784
rect 3784 11752 3816 11784
rect 3856 11752 3888 11784
rect 3928 11752 3960 11784
rect 40 11680 72 11712
rect 112 11680 144 11712
rect 184 11680 216 11712
rect 256 11680 288 11712
rect 328 11680 360 11712
rect 400 11680 432 11712
rect 472 11680 504 11712
rect 544 11680 576 11712
rect 616 11680 648 11712
rect 688 11680 720 11712
rect 760 11680 792 11712
rect 832 11680 864 11712
rect 904 11680 936 11712
rect 976 11680 1008 11712
rect 1048 11680 1080 11712
rect 1120 11680 1152 11712
rect 1192 11680 1224 11712
rect 1264 11680 1296 11712
rect 1336 11680 1368 11712
rect 1408 11680 1440 11712
rect 1480 11680 1512 11712
rect 1552 11680 1584 11712
rect 1624 11680 1656 11712
rect 1696 11680 1728 11712
rect 1768 11680 1800 11712
rect 1840 11680 1872 11712
rect 1912 11680 1944 11712
rect 1984 11680 2016 11712
rect 2056 11680 2088 11712
rect 2128 11680 2160 11712
rect 2200 11680 2232 11712
rect 2272 11680 2304 11712
rect 2344 11680 2376 11712
rect 2416 11680 2448 11712
rect 2488 11680 2520 11712
rect 2560 11680 2592 11712
rect 2632 11680 2664 11712
rect 2704 11680 2736 11712
rect 2776 11680 2808 11712
rect 2848 11680 2880 11712
rect 2920 11680 2952 11712
rect 2992 11680 3024 11712
rect 3064 11680 3096 11712
rect 3136 11680 3168 11712
rect 3208 11680 3240 11712
rect 3280 11680 3312 11712
rect 3352 11680 3384 11712
rect 3424 11680 3456 11712
rect 3496 11680 3528 11712
rect 3568 11680 3600 11712
rect 3640 11680 3672 11712
rect 3712 11680 3744 11712
rect 3784 11680 3816 11712
rect 3856 11680 3888 11712
rect 3928 11680 3960 11712
rect 40 11608 72 11640
rect 112 11608 144 11640
rect 184 11608 216 11640
rect 256 11608 288 11640
rect 328 11608 360 11640
rect 400 11608 432 11640
rect 472 11608 504 11640
rect 544 11608 576 11640
rect 616 11608 648 11640
rect 688 11608 720 11640
rect 760 11608 792 11640
rect 832 11608 864 11640
rect 904 11608 936 11640
rect 976 11608 1008 11640
rect 1048 11608 1080 11640
rect 1120 11608 1152 11640
rect 1192 11608 1224 11640
rect 1264 11608 1296 11640
rect 1336 11608 1368 11640
rect 1408 11608 1440 11640
rect 1480 11608 1512 11640
rect 1552 11608 1584 11640
rect 1624 11608 1656 11640
rect 1696 11608 1728 11640
rect 1768 11608 1800 11640
rect 1840 11608 1872 11640
rect 1912 11608 1944 11640
rect 1984 11608 2016 11640
rect 2056 11608 2088 11640
rect 2128 11608 2160 11640
rect 2200 11608 2232 11640
rect 2272 11608 2304 11640
rect 2344 11608 2376 11640
rect 2416 11608 2448 11640
rect 2488 11608 2520 11640
rect 2560 11608 2592 11640
rect 2632 11608 2664 11640
rect 2704 11608 2736 11640
rect 2776 11608 2808 11640
rect 2848 11608 2880 11640
rect 2920 11608 2952 11640
rect 2992 11608 3024 11640
rect 3064 11608 3096 11640
rect 3136 11608 3168 11640
rect 3208 11608 3240 11640
rect 3280 11608 3312 11640
rect 3352 11608 3384 11640
rect 3424 11608 3456 11640
rect 3496 11608 3528 11640
rect 3568 11608 3600 11640
rect 3640 11608 3672 11640
rect 3712 11608 3744 11640
rect 3784 11608 3816 11640
rect 3856 11608 3888 11640
rect 3928 11608 3960 11640
rect 40 11536 72 11568
rect 112 11536 144 11568
rect 184 11536 216 11568
rect 256 11536 288 11568
rect 328 11536 360 11568
rect 400 11536 432 11568
rect 472 11536 504 11568
rect 544 11536 576 11568
rect 616 11536 648 11568
rect 688 11536 720 11568
rect 760 11536 792 11568
rect 832 11536 864 11568
rect 904 11536 936 11568
rect 976 11536 1008 11568
rect 1048 11536 1080 11568
rect 1120 11536 1152 11568
rect 1192 11536 1224 11568
rect 1264 11536 1296 11568
rect 1336 11536 1368 11568
rect 1408 11536 1440 11568
rect 1480 11536 1512 11568
rect 1552 11536 1584 11568
rect 1624 11536 1656 11568
rect 1696 11536 1728 11568
rect 1768 11536 1800 11568
rect 1840 11536 1872 11568
rect 1912 11536 1944 11568
rect 1984 11536 2016 11568
rect 2056 11536 2088 11568
rect 2128 11536 2160 11568
rect 2200 11536 2232 11568
rect 2272 11536 2304 11568
rect 2344 11536 2376 11568
rect 2416 11536 2448 11568
rect 2488 11536 2520 11568
rect 2560 11536 2592 11568
rect 2632 11536 2664 11568
rect 2704 11536 2736 11568
rect 2776 11536 2808 11568
rect 2848 11536 2880 11568
rect 2920 11536 2952 11568
rect 2992 11536 3024 11568
rect 3064 11536 3096 11568
rect 3136 11536 3168 11568
rect 3208 11536 3240 11568
rect 3280 11536 3312 11568
rect 3352 11536 3384 11568
rect 3424 11536 3456 11568
rect 3496 11536 3528 11568
rect 3568 11536 3600 11568
rect 3640 11536 3672 11568
rect 3712 11536 3744 11568
rect 3784 11536 3816 11568
rect 3856 11536 3888 11568
rect 3928 11536 3960 11568
rect 40 11464 72 11496
rect 112 11464 144 11496
rect 184 11464 216 11496
rect 256 11464 288 11496
rect 328 11464 360 11496
rect 400 11464 432 11496
rect 472 11464 504 11496
rect 544 11464 576 11496
rect 616 11464 648 11496
rect 688 11464 720 11496
rect 760 11464 792 11496
rect 832 11464 864 11496
rect 904 11464 936 11496
rect 976 11464 1008 11496
rect 1048 11464 1080 11496
rect 1120 11464 1152 11496
rect 1192 11464 1224 11496
rect 1264 11464 1296 11496
rect 1336 11464 1368 11496
rect 1408 11464 1440 11496
rect 1480 11464 1512 11496
rect 1552 11464 1584 11496
rect 1624 11464 1656 11496
rect 1696 11464 1728 11496
rect 1768 11464 1800 11496
rect 1840 11464 1872 11496
rect 1912 11464 1944 11496
rect 1984 11464 2016 11496
rect 2056 11464 2088 11496
rect 2128 11464 2160 11496
rect 2200 11464 2232 11496
rect 2272 11464 2304 11496
rect 2344 11464 2376 11496
rect 2416 11464 2448 11496
rect 2488 11464 2520 11496
rect 2560 11464 2592 11496
rect 2632 11464 2664 11496
rect 2704 11464 2736 11496
rect 2776 11464 2808 11496
rect 2848 11464 2880 11496
rect 2920 11464 2952 11496
rect 2992 11464 3024 11496
rect 3064 11464 3096 11496
rect 3136 11464 3168 11496
rect 3208 11464 3240 11496
rect 3280 11464 3312 11496
rect 3352 11464 3384 11496
rect 3424 11464 3456 11496
rect 3496 11464 3528 11496
rect 3568 11464 3600 11496
rect 3640 11464 3672 11496
rect 3712 11464 3744 11496
rect 3784 11464 3816 11496
rect 3856 11464 3888 11496
rect 3928 11464 3960 11496
rect 40 11392 72 11424
rect 112 11392 144 11424
rect 184 11392 216 11424
rect 256 11392 288 11424
rect 328 11392 360 11424
rect 400 11392 432 11424
rect 472 11392 504 11424
rect 544 11392 576 11424
rect 616 11392 648 11424
rect 688 11392 720 11424
rect 760 11392 792 11424
rect 832 11392 864 11424
rect 904 11392 936 11424
rect 976 11392 1008 11424
rect 1048 11392 1080 11424
rect 1120 11392 1152 11424
rect 1192 11392 1224 11424
rect 1264 11392 1296 11424
rect 1336 11392 1368 11424
rect 1408 11392 1440 11424
rect 1480 11392 1512 11424
rect 1552 11392 1584 11424
rect 1624 11392 1656 11424
rect 1696 11392 1728 11424
rect 1768 11392 1800 11424
rect 1840 11392 1872 11424
rect 1912 11392 1944 11424
rect 1984 11392 2016 11424
rect 2056 11392 2088 11424
rect 2128 11392 2160 11424
rect 2200 11392 2232 11424
rect 2272 11392 2304 11424
rect 2344 11392 2376 11424
rect 2416 11392 2448 11424
rect 2488 11392 2520 11424
rect 2560 11392 2592 11424
rect 2632 11392 2664 11424
rect 2704 11392 2736 11424
rect 2776 11392 2808 11424
rect 2848 11392 2880 11424
rect 2920 11392 2952 11424
rect 2992 11392 3024 11424
rect 3064 11392 3096 11424
rect 3136 11392 3168 11424
rect 3208 11392 3240 11424
rect 3280 11392 3312 11424
rect 3352 11392 3384 11424
rect 3424 11392 3456 11424
rect 3496 11392 3528 11424
rect 3568 11392 3600 11424
rect 3640 11392 3672 11424
rect 3712 11392 3744 11424
rect 3784 11392 3816 11424
rect 3856 11392 3888 11424
rect 3928 11392 3960 11424
rect 40 11320 72 11352
rect 112 11320 144 11352
rect 184 11320 216 11352
rect 256 11320 288 11352
rect 328 11320 360 11352
rect 400 11320 432 11352
rect 472 11320 504 11352
rect 544 11320 576 11352
rect 616 11320 648 11352
rect 688 11320 720 11352
rect 760 11320 792 11352
rect 832 11320 864 11352
rect 904 11320 936 11352
rect 976 11320 1008 11352
rect 1048 11320 1080 11352
rect 1120 11320 1152 11352
rect 1192 11320 1224 11352
rect 1264 11320 1296 11352
rect 1336 11320 1368 11352
rect 1408 11320 1440 11352
rect 1480 11320 1512 11352
rect 1552 11320 1584 11352
rect 1624 11320 1656 11352
rect 1696 11320 1728 11352
rect 1768 11320 1800 11352
rect 1840 11320 1872 11352
rect 1912 11320 1944 11352
rect 1984 11320 2016 11352
rect 2056 11320 2088 11352
rect 2128 11320 2160 11352
rect 2200 11320 2232 11352
rect 2272 11320 2304 11352
rect 2344 11320 2376 11352
rect 2416 11320 2448 11352
rect 2488 11320 2520 11352
rect 2560 11320 2592 11352
rect 2632 11320 2664 11352
rect 2704 11320 2736 11352
rect 2776 11320 2808 11352
rect 2848 11320 2880 11352
rect 2920 11320 2952 11352
rect 2992 11320 3024 11352
rect 3064 11320 3096 11352
rect 3136 11320 3168 11352
rect 3208 11320 3240 11352
rect 3280 11320 3312 11352
rect 3352 11320 3384 11352
rect 3424 11320 3456 11352
rect 3496 11320 3528 11352
rect 3568 11320 3600 11352
rect 3640 11320 3672 11352
rect 3712 11320 3744 11352
rect 3784 11320 3816 11352
rect 3856 11320 3888 11352
rect 3928 11320 3960 11352
rect 40 11248 72 11280
rect 112 11248 144 11280
rect 184 11248 216 11280
rect 256 11248 288 11280
rect 328 11248 360 11280
rect 400 11248 432 11280
rect 472 11248 504 11280
rect 544 11248 576 11280
rect 616 11248 648 11280
rect 688 11248 720 11280
rect 760 11248 792 11280
rect 832 11248 864 11280
rect 904 11248 936 11280
rect 976 11248 1008 11280
rect 1048 11248 1080 11280
rect 1120 11248 1152 11280
rect 1192 11248 1224 11280
rect 1264 11248 1296 11280
rect 1336 11248 1368 11280
rect 1408 11248 1440 11280
rect 1480 11248 1512 11280
rect 1552 11248 1584 11280
rect 1624 11248 1656 11280
rect 1696 11248 1728 11280
rect 1768 11248 1800 11280
rect 1840 11248 1872 11280
rect 1912 11248 1944 11280
rect 1984 11248 2016 11280
rect 2056 11248 2088 11280
rect 2128 11248 2160 11280
rect 2200 11248 2232 11280
rect 2272 11248 2304 11280
rect 2344 11248 2376 11280
rect 2416 11248 2448 11280
rect 2488 11248 2520 11280
rect 2560 11248 2592 11280
rect 2632 11248 2664 11280
rect 2704 11248 2736 11280
rect 2776 11248 2808 11280
rect 2848 11248 2880 11280
rect 2920 11248 2952 11280
rect 2992 11248 3024 11280
rect 3064 11248 3096 11280
rect 3136 11248 3168 11280
rect 3208 11248 3240 11280
rect 3280 11248 3312 11280
rect 3352 11248 3384 11280
rect 3424 11248 3456 11280
rect 3496 11248 3528 11280
rect 3568 11248 3600 11280
rect 3640 11248 3672 11280
rect 3712 11248 3744 11280
rect 3784 11248 3816 11280
rect 3856 11248 3888 11280
rect 3928 11248 3960 11280
rect 40 11176 72 11208
rect 112 11176 144 11208
rect 184 11176 216 11208
rect 256 11176 288 11208
rect 328 11176 360 11208
rect 400 11176 432 11208
rect 472 11176 504 11208
rect 544 11176 576 11208
rect 616 11176 648 11208
rect 688 11176 720 11208
rect 760 11176 792 11208
rect 832 11176 864 11208
rect 904 11176 936 11208
rect 976 11176 1008 11208
rect 1048 11176 1080 11208
rect 1120 11176 1152 11208
rect 1192 11176 1224 11208
rect 1264 11176 1296 11208
rect 1336 11176 1368 11208
rect 1408 11176 1440 11208
rect 1480 11176 1512 11208
rect 1552 11176 1584 11208
rect 1624 11176 1656 11208
rect 1696 11176 1728 11208
rect 1768 11176 1800 11208
rect 1840 11176 1872 11208
rect 1912 11176 1944 11208
rect 1984 11176 2016 11208
rect 2056 11176 2088 11208
rect 2128 11176 2160 11208
rect 2200 11176 2232 11208
rect 2272 11176 2304 11208
rect 2344 11176 2376 11208
rect 2416 11176 2448 11208
rect 2488 11176 2520 11208
rect 2560 11176 2592 11208
rect 2632 11176 2664 11208
rect 2704 11176 2736 11208
rect 2776 11176 2808 11208
rect 2848 11176 2880 11208
rect 2920 11176 2952 11208
rect 2992 11176 3024 11208
rect 3064 11176 3096 11208
rect 3136 11176 3168 11208
rect 3208 11176 3240 11208
rect 3280 11176 3312 11208
rect 3352 11176 3384 11208
rect 3424 11176 3456 11208
rect 3496 11176 3528 11208
rect 3568 11176 3600 11208
rect 3640 11176 3672 11208
rect 3712 11176 3744 11208
rect 3784 11176 3816 11208
rect 3856 11176 3888 11208
rect 3928 11176 3960 11208
rect 40 11104 72 11136
rect 112 11104 144 11136
rect 184 11104 216 11136
rect 256 11104 288 11136
rect 328 11104 360 11136
rect 400 11104 432 11136
rect 472 11104 504 11136
rect 544 11104 576 11136
rect 616 11104 648 11136
rect 688 11104 720 11136
rect 760 11104 792 11136
rect 832 11104 864 11136
rect 904 11104 936 11136
rect 976 11104 1008 11136
rect 1048 11104 1080 11136
rect 1120 11104 1152 11136
rect 1192 11104 1224 11136
rect 1264 11104 1296 11136
rect 1336 11104 1368 11136
rect 1408 11104 1440 11136
rect 1480 11104 1512 11136
rect 1552 11104 1584 11136
rect 1624 11104 1656 11136
rect 1696 11104 1728 11136
rect 1768 11104 1800 11136
rect 1840 11104 1872 11136
rect 1912 11104 1944 11136
rect 1984 11104 2016 11136
rect 2056 11104 2088 11136
rect 2128 11104 2160 11136
rect 2200 11104 2232 11136
rect 2272 11104 2304 11136
rect 2344 11104 2376 11136
rect 2416 11104 2448 11136
rect 2488 11104 2520 11136
rect 2560 11104 2592 11136
rect 2632 11104 2664 11136
rect 2704 11104 2736 11136
rect 2776 11104 2808 11136
rect 2848 11104 2880 11136
rect 2920 11104 2952 11136
rect 2992 11104 3024 11136
rect 3064 11104 3096 11136
rect 3136 11104 3168 11136
rect 3208 11104 3240 11136
rect 3280 11104 3312 11136
rect 3352 11104 3384 11136
rect 3424 11104 3456 11136
rect 3496 11104 3528 11136
rect 3568 11104 3600 11136
rect 3640 11104 3672 11136
rect 3712 11104 3744 11136
rect 3784 11104 3816 11136
rect 3856 11104 3888 11136
rect 3928 11104 3960 11136
rect 40 11032 72 11064
rect 112 11032 144 11064
rect 184 11032 216 11064
rect 256 11032 288 11064
rect 328 11032 360 11064
rect 400 11032 432 11064
rect 472 11032 504 11064
rect 544 11032 576 11064
rect 616 11032 648 11064
rect 688 11032 720 11064
rect 760 11032 792 11064
rect 832 11032 864 11064
rect 904 11032 936 11064
rect 976 11032 1008 11064
rect 1048 11032 1080 11064
rect 1120 11032 1152 11064
rect 1192 11032 1224 11064
rect 1264 11032 1296 11064
rect 1336 11032 1368 11064
rect 1408 11032 1440 11064
rect 1480 11032 1512 11064
rect 1552 11032 1584 11064
rect 1624 11032 1656 11064
rect 1696 11032 1728 11064
rect 1768 11032 1800 11064
rect 1840 11032 1872 11064
rect 1912 11032 1944 11064
rect 1984 11032 2016 11064
rect 2056 11032 2088 11064
rect 2128 11032 2160 11064
rect 2200 11032 2232 11064
rect 2272 11032 2304 11064
rect 2344 11032 2376 11064
rect 2416 11032 2448 11064
rect 2488 11032 2520 11064
rect 2560 11032 2592 11064
rect 2632 11032 2664 11064
rect 2704 11032 2736 11064
rect 2776 11032 2808 11064
rect 2848 11032 2880 11064
rect 2920 11032 2952 11064
rect 2992 11032 3024 11064
rect 3064 11032 3096 11064
rect 3136 11032 3168 11064
rect 3208 11032 3240 11064
rect 3280 11032 3312 11064
rect 3352 11032 3384 11064
rect 3424 11032 3456 11064
rect 3496 11032 3528 11064
rect 3568 11032 3600 11064
rect 3640 11032 3672 11064
rect 3712 11032 3744 11064
rect 3784 11032 3816 11064
rect 3856 11032 3888 11064
rect 3928 11032 3960 11064
rect 40 10960 72 10992
rect 112 10960 144 10992
rect 184 10960 216 10992
rect 256 10960 288 10992
rect 328 10960 360 10992
rect 400 10960 432 10992
rect 472 10960 504 10992
rect 544 10960 576 10992
rect 616 10960 648 10992
rect 688 10960 720 10992
rect 760 10960 792 10992
rect 832 10960 864 10992
rect 904 10960 936 10992
rect 976 10960 1008 10992
rect 1048 10960 1080 10992
rect 1120 10960 1152 10992
rect 1192 10960 1224 10992
rect 1264 10960 1296 10992
rect 1336 10960 1368 10992
rect 1408 10960 1440 10992
rect 1480 10960 1512 10992
rect 1552 10960 1584 10992
rect 1624 10960 1656 10992
rect 1696 10960 1728 10992
rect 1768 10960 1800 10992
rect 1840 10960 1872 10992
rect 1912 10960 1944 10992
rect 1984 10960 2016 10992
rect 2056 10960 2088 10992
rect 2128 10960 2160 10992
rect 2200 10960 2232 10992
rect 2272 10960 2304 10992
rect 2344 10960 2376 10992
rect 2416 10960 2448 10992
rect 2488 10960 2520 10992
rect 2560 10960 2592 10992
rect 2632 10960 2664 10992
rect 2704 10960 2736 10992
rect 2776 10960 2808 10992
rect 2848 10960 2880 10992
rect 2920 10960 2952 10992
rect 2992 10960 3024 10992
rect 3064 10960 3096 10992
rect 3136 10960 3168 10992
rect 3208 10960 3240 10992
rect 3280 10960 3312 10992
rect 3352 10960 3384 10992
rect 3424 10960 3456 10992
rect 3496 10960 3528 10992
rect 3568 10960 3600 10992
rect 3640 10960 3672 10992
rect 3712 10960 3744 10992
rect 3784 10960 3816 10992
rect 3856 10960 3888 10992
rect 3928 10960 3960 10992
rect 40 10888 72 10920
rect 112 10888 144 10920
rect 184 10888 216 10920
rect 256 10888 288 10920
rect 328 10888 360 10920
rect 400 10888 432 10920
rect 472 10888 504 10920
rect 544 10888 576 10920
rect 616 10888 648 10920
rect 688 10888 720 10920
rect 760 10888 792 10920
rect 832 10888 864 10920
rect 904 10888 936 10920
rect 976 10888 1008 10920
rect 1048 10888 1080 10920
rect 1120 10888 1152 10920
rect 1192 10888 1224 10920
rect 1264 10888 1296 10920
rect 1336 10888 1368 10920
rect 1408 10888 1440 10920
rect 1480 10888 1512 10920
rect 1552 10888 1584 10920
rect 1624 10888 1656 10920
rect 1696 10888 1728 10920
rect 1768 10888 1800 10920
rect 1840 10888 1872 10920
rect 1912 10888 1944 10920
rect 1984 10888 2016 10920
rect 2056 10888 2088 10920
rect 2128 10888 2160 10920
rect 2200 10888 2232 10920
rect 2272 10888 2304 10920
rect 2344 10888 2376 10920
rect 2416 10888 2448 10920
rect 2488 10888 2520 10920
rect 2560 10888 2592 10920
rect 2632 10888 2664 10920
rect 2704 10888 2736 10920
rect 2776 10888 2808 10920
rect 2848 10888 2880 10920
rect 2920 10888 2952 10920
rect 2992 10888 3024 10920
rect 3064 10888 3096 10920
rect 3136 10888 3168 10920
rect 3208 10888 3240 10920
rect 3280 10888 3312 10920
rect 3352 10888 3384 10920
rect 3424 10888 3456 10920
rect 3496 10888 3528 10920
rect 3568 10888 3600 10920
rect 3640 10888 3672 10920
rect 3712 10888 3744 10920
rect 3784 10888 3816 10920
rect 3856 10888 3888 10920
rect 3928 10888 3960 10920
rect 40 10816 72 10848
rect 112 10816 144 10848
rect 184 10816 216 10848
rect 256 10816 288 10848
rect 328 10816 360 10848
rect 400 10816 432 10848
rect 472 10816 504 10848
rect 544 10816 576 10848
rect 616 10816 648 10848
rect 688 10816 720 10848
rect 760 10816 792 10848
rect 832 10816 864 10848
rect 904 10816 936 10848
rect 976 10816 1008 10848
rect 1048 10816 1080 10848
rect 1120 10816 1152 10848
rect 1192 10816 1224 10848
rect 1264 10816 1296 10848
rect 1336 10816 1368 10848
rect 1408 10816 1440 10848
rect 1480 10816 1512 10848
rect 1552 10816 1584 10848
rect 1624 10816 1656 10848
rect 1696 10816 1728 10848
rect 1768 10816 1800 10848
rect 1840 10816 1872 10848
rect 1912 10816 1944 10848
rect 1984 10816 2016 10848
rect 2056 10816 2088 10848
rect 2128 10816 2160 10848
rect 2200 10816 2232 10848
rect 2272 10816 2304 10848
rect 2344 10816 2376 10848
rect 2416 10816 2448 10848
rect 2488 10816 2520 10848
rect 2560 10816 2592 10848
rect 2632 10816 2664 10848
rect 2704 10816 2736 10848
rect 2776 10816 2808 10848
rect 2848 10816 2880 10848
rect 2920 10816 2952 10848
rect 2992 10816 3024 10848
rect 3064 10816 3096 10848
rect 3136 10816 3168 10848
rect 3208 10816 3240 10848
rect 3280 10816 3312 10848
rect 3352 10816 3384 10848
rect 3424 10816 3456 10848
rect 3496 10816 3528 10848
rect 3568 10816 3600 10848
rect 3640 10816 3672 10848
rect 3712 10816 3744 10848
rect 3784 10816 3816 10848
rect 3856 10816 3888 10848
rect 3928 10816 3960 10848
rect 40 10744 72 10776
rect 112 10744 144 10776
rect 184 10744 216 10776
rect 256 10744 288 10776
rect 328 10744 360 10776
rect 400 10744 432 10776
rect 472 10744 504 10776
rect 544 10744 576 10776
rect 616 10744 648 10776
rect 688 10744 720 10776
rect 760 10744 792 10776
rect 832 10744 864 10776
rect 904 10744 936 10776
rect 976 10744 1008 10776
rect 1048 10744 1080 10776
rect 1120 10744 1152 10776
rect 1192 10744 1224 10776
rect 1264 10744 1296 10776
rect 1336 10744 1368 10776
rect 1408 10744 1440 10776
rect 1480 10744 1512 10776
rect 1552 10744 1584 10776
rect 1624 10744 1656 10776
rect 1696 10744 1728 10776
rect 1768 10744 1800 10776
rect 1840 10744 1872 10776
rect 1912 10744 1944 10776
rect 1984 10744 2016 10776
rect 2056 10744 2088 10776
rect 2128 10744 2160 10776
rect 2200 10744 2232 10776
rect 2272 10744 2304 10776
rect 2344 10744 2376 10776
rect 2416 10744 2448 10776
rect 2488 10744 2520 10776
rect 2560 10744 2592 10776
rect 2632 10744 2664 10776
rect 2704 10744 2736 10776
rect 2776 10744 2808 10776
rect 2848 10744 2880 10776
rect 2920 10744 2952 10776
rect 2992 10744 3024 10776
rect 3064 10744 3096 10776
rect 3136 10744 3168 10776
rect 3208 10744 3240 10776
rect 3280 10744 3312 10776
rect 3352 10744 3384 10776
rect 3424 10744 3456 10776
rect 3496 10744 3528 10776
rect 3568 10744 3600 10776
rect 3640 10744 3672 10776
rect 3712 10744 3744 10776
rect 3784 10744 3816 10776
rect 3856 10744 3888 10776
rect 3928 10744 3960 10776
rect 40 10672 72 10704
rect 112 10672 144 10704
rect 184 10672 216 10704
rect 256 10672 288 10704
rect 328 10672 360 10704
rect 400 10672 432 10704
rect 472 10672 504 10704
rect 544 10672 576 10704
rect 616 10672 648 10704
rect 688 10672 720 10704
rect 760 10672 792 10704
rect 832 10672 864 10704
rect 904 10672 936 10704
rect 976 10672 1008 10704
rect 1048 10672 1080 10704
rect 1120 10672 1152 10704
rect 1192 10672 1224 10704
rect 1264 10672 1296 10704
rect 1336 10672 1368 10704
rect 1408 10672 1440 10704
rect 1480 10672 1512 10704
rect 1552 10672 1584 10704
rect 1624 10672 1656 10704
rect 1696 10672 1728 10704
rect 1768 10672 1800 10704
rect 1840 10672 1872 10704
rect 1912 10672 1944 10704
rect 1984 10672 2016 10704
rect 2056 10672 2088 10704
rect 2128 10672 2160 10704
rect 2200 10672 2232 10704
rect 2272 10672 2304 10704
rect 2344 10672 2376 10704
rect 2416 10672 2448 10704
rect 2488 10672 2520 10704
rect 2560 10672 2592 10704
rect 2632 10672 2664 10704
rect 2704 10672 2736 10704
rect 2776 10672 2808 10704
rect 2848 10672 2880 10704
rect 2920 10672 2952 10704
rect 2992 10672 3024 10704
rect 3064 10672 3096 10704
rect 3136 10672 3168 10704
rect 3208 10672 3240 10704
rect 3280 10672 3312 10704
rect 3352 10672 3384 10704
rect 3424 10672 3456 10704
rect 3496 10672 3528 10704
rect 3568 10672 3600 10704
rect 3640 10672 3672 10704
rect 3712 10672 3744 10704
rect 3784 10672 3816 10704
rect 3856 10672 3888 10704
rect 3928 10672 3960 10704
rect 40 10600 72 10632
rect 112 10600 144 10632
rect 184 10600 216 10632
rect 256 10600 288 10632
rect 328 10600 360 10632
rect 400 10600 432 10632
rect 472 10600 504 10632
rect 544 10600 576 10632
rect 616 10600 648 10632
rect 688 10600 720 10632
rect 760 10600 792 10632
rect 832 10600 864 10632
rect 904 10600 936 10632
rect 976 10600 1008 10632
rect 1048 10600 1080 10632
rect 1120 10600 1152 10632
rect 1192 10600 1224 10632
rect 1264 10600 1296 10632
rect 1336 10600 1368 10632
rect 1408 10600 1440 10632
rect 1480 10600 1512 10632
rect 1552 10600 1584 10632
rect 1624 10600 1656 10632
rect 1696 10600 1728 10632
rect 1768 10600 1800 10632
rect 1840 10600 1872 10632
rect 1912 10600 1944 10632
rect 1984 10600 2016 10632
rect 2056 10600 2088 10632
rect 2128 10600 2160 10632
rect 2200 10600 2232 10632
rect 2272 10600 2304 10632
rect 2344 10600 2376 10632
rect 2416 10600 2448 10632
rect 2488 10600 2520 10632
rect 2560 10600 2592 10632
rect 2632 10600 2664 10632
rect 2704 10600 2736 10632
rect 2776 10600 2808 10632
rect 2848 10600 2880 10632
rect 2920 10600 2952 10632
rect 2992 10600 3024 10632
rect 3064 10600 3096 10632
rect 3136 10600 3168 10632
rect 3208 10600 3240 10632
rect 3280 10600 3312 10632
rect 3352 10600 3384 10632
rect 3424 10600 3456 10632
rect 3496 10600 3528 10632
rect 3568 10600 3600 10632
rect 3640 10600 3672 10632
rect 3712 10600 3744 10632
rect 3784 10600 3816 10632
rect 3856 10600 3888 10632
rect 3928 10600 3960 10632
rect 40 10528 72 10560
rect 112 10528 144 10560
rect 184 10528 216 10560
rect 256 10528 288 10560
rect 328 10528 360 10560
rect 400 10528 432 10560
rect 472 10528 504 10560
rect 544 10528 576 10560
rect 616 10528 648 10560
rect 688 10528 720 10560
rect 760 10528 792 10560
rect 832 10528 864 10560
rect 904 10528 936 10560
rect 976 10528 1008 10560
rect 1048 10528 1080 10560
rect 1120 10528 1152 10560
rect 1192 10528 1224 10560
rect 1264 10528 1296 10560
rect 1336 10528 1368 10560
rect 1408 10528 1440 10560
rect 1480 10528 1512 10560
rect 1552 10528 1584 10560
rect 1624 10528 1656 10560
rect 1696 10528 1728 10560
rect 1768 10528 1800 10560
rect 1840 10528 1872 10560
rect 1912 10528 1944 10560
rect 1984 10528 2016 10560
rect 2056 10528 2088 10560
rect 2128 10528 2160 10560
rect 2200 10528 2232 10560
rect 2272 10528 2304 10560
rect 2344 10528 2376 10560
rect 2416 10528 2448 10560
rect 2488 10528 2520 10560
rect 2560 10528 2592 10560
rect 2632 10528 2664 10560
rect 2704 10528 2736 10560
rect 2776 10528 2808 10560
rect 2848 10528 2880 10560
rect 2920 10528 2952 10560
rect 2992 10528 3024 10560
rect 3064 10528 3096 10560
rect 3136 10528 3168 10560
rect 3208 10528 3240 10560
rect 3280 10528 3312 10560
rect 3352 10528 3384 10560
rect 3424 10528 3456 10560
rect 3496 10528 3528 10560
rect 3568 10528 3600 10560
rect 3640 10528 3672 10560
rect 3712 10528 3744 10560
rect 3784 10528 3816 10560
rect 3856 10528 3888 10560
rect 3928 10528 3960 10560
rect 40 10456 72 10488
rect 112 10456 144 10488
rect 184 10456 216 10488
rect 256 10456 288 10488
rect 328 10456 360 10488
rect 400 10456 432 10488
rect 472 10456 504 10488
rect 544 10456 576 10488
rect 616 10456 648 10488
rect 688 10456 720 10488
rect 760 10456 792 10488
rect 832 10456 864 10488
rect 904 10456 936 10488
rect 976 10456 1008 10488
rect 1048 10456 1080 10488
rect 1120 10456 1152 10488
rect 1192 10456 1224 10488
rect 1264 10456 1296 10488
rect 1336 10456 1368 10488
rect 1408 10456 1440 10488
rect 1480 10456 1512 10488
rect 1552 10456 1584 10488
rect 1624 10456 1656 10488
rect 1696 10456 1728 10488
rect 1768 10456 1800 10488
rect 1840 10456 1872 10488
rect 1912 10456 1944 10488
rect 1984 10456 2016 10488
rect 2056 10456 2088 10488
rect 2128 10456 2160 10488
rect 2200 10456 2232 10488
rect 2272 10456 2304 10488
rect 2344 10456 2376 10488
rect 2416 10456 2448 10488
rect 2488 10456 2520 10488
rect 2560 10456 2592 10488
rect 2632 10456 2664 10488
rect 2704 10456 2736 10488
rect 2776 10456 2808 10488
rect 2848 10456 2880 10488
rect 2920 10456 2952 10488
rect 2992 10456 3024 10488
rect 3064 10456 3096 10488
rect 3136 10456 3168 10488
rect 3208 10456 3240 10488
rect 3280 10456 3312 10488
rect 3352 10456 3384 10488
rect 3424 10456 3456 10488
rect 3496 10456 3528 10488
rect 3568 10456 3600 10488
rect 3640 10456 3672 10488
rect 3712 10456 3744 10488
rect 3784 10456 3816 10488
rect 3856 10456 3888 10488
rect 3928 10456 3960 10488
rect 40 10384 72 10416
rect 112 10384 144 10416
rect 184 10384 216 10416
rect 256 10384 288 10416
rect 328 10384 360 10416
rect 400 10384 432 10416
rect 472 10384 504 10416
rect 544 10384 576 10416
rect 616 10384 648 10416
rect 688 10384 720 10416
rect 760 10384 792 10416
rect 832 10384 864 10416
rect 904 10384 936 10416
rect 976 10384 1008 10416
rect 1048 10384 1080 10416
rect 1120 10384 1152 10416
rect 1192 10384 1224 10416
rect 1264 10384 1296 10416
rect 1336 10384 1368 10416
rect 1408 10384 1440 10416
rect 1480 10384 1512 10416
rect 1552 10384 1584 10416
rect 1624 10384 1656 10416
rect 1696 10384 1728 10416
rect 1768 10384 1800 10416
rect 1840 10384 1872 10416
rect 1912 10384 1944 10416
rect 1984 10384 2016 10416
rect 2056 10384 2088 10416
rect 2128 10384 2160 10416
rect 2200 10384 2232 10416
rect 2272 10384 2304 10416
rect 2344 10384 2376 10416
rect 2416 10384 2448 10416
rect 2488 10384 2520 10416
rect 2560 10384 2592 10416
rect 2632 10384 2664 10416
rect 2704 10384 2736 10416
rect 2776 10384 2808 10416
rect 2848 10384 2880 10416
rect 2920 10384 2952 10416
rect 2992 10384 3024 10416
rect 3064 10384 3096 10416
rect 3136 10384 3168 10416
rect 3208 10384 3240 10416
rect 3280 10384 3312 10416
rect 3352 10384 3384 10416
rect 3424 10384 3456 10416
rect 3496 10384 3528 10416
rect 3568 10384 3600 10416
rect 3640 10384 3672 10416
rect 3712 10384 3744 10416
rect 3784 10384 3816 10416
rect 3856 10384 3888 10416
rect 3928 10384 3960 10416
rect 40 10312 72 10344
rect 112 10312 144 10344
rect 184 10312 216 10344
rect 256 10312 288 10344
rect 328 10312 360 10344
rect 400 10312 432 10344
rect 472 10312 504 10344
rect 544 10312 576 10344
rect 616 10312 648 10344
rect 688 10312 720 10344
rect 760 10312 792 10344
rect 832 10312 864 10344
rect 904 10312 936 10344
rect 976 10312 1008 10344
rect 1048 10312 1080 10344
rect 1120 10312 1152 10344
rect 1192 10312 1224 10344
rect 1264 10312 1296 10344
rect 1336 10312 1368 10344
rect 1408 10312 1440 10344
rect 1480 10312 1512 10344
rect 1552 10312 1584 10344
rect 1624 10312 1656 10344
rect 1696 10312 1728 10344
rect 1768 10312 1800 10344
rect 1840 10312 1872 10344
rect 1912 10312 1944 10344
rect 1984 10312 2016 10344
rect 2056 10312 2088 10344
rect 2128 10312 2160 10344
rect 2200 10312 2232 10344
rect 2272 10312 2304 10344
rect 2344 10312 2376 10344
rect 2416 10312 2448 10344
rect 2488 10312 2520 10344
rect 2560 10312 2592 10344
rect 2632 10312 2664 10344
rect 2704 10312 2736 10344
rect 2776 10312 2808 10344
rect 2848 10312 2880 10344
rect 2920 10312 2952 10344
rect 2992 10312 3024 10344
rect 3064 10312 3096 10344
rect 3136 10312 3168 10344
rect 3208 10312 3240 10344
rect 3280 10312 3312 10344
rect 3352 10312 3384 10344
rect 3424 10312 3456 10344
rect 3496 10312 3528 10344
rect 3568 10312 3600 10344
rect 3640 10312 3672 10344
rect 3712 10312 3744 10344
rect 3784 10312 3816 10344
rect 3856 10312 3888 10344
rect 3928 10312 3960 10344
rect 40 10240 72 10272
rect 112 10240 144 10272
rect 184 10240 216 10272
rect 256 10240 288 10272
rect 328 10240 360 10272
rect 400 10240 432 10272
rect 472 10240 504 10272
rect 544 10240 576 10272
rect 616 10240 648 10272
rect 688 10240 720 10272
rect 760 10240 792 10272
rect 832 10240 864 10272
rect 904 10240 936 10272
rect 976 10240 1008 10272
rect 1048 10240 1080 10272
rect 1120 10240 1152 10272
rect 1192 10240 1224 10272
rect 1264 10240 1296 10272
rect 1336 10240 1368 10272
rect 1408 10240 1440 10272
rect 1480 10240 1512 10272
rect 1552 10240 1584 10272
rect 1624 10240 1656 10272
rect 1696 10240 1728 10272
rect 1768 10240 1800 10272
rect 1840 10240 1872 10272
rect 1912 10240 1944 10272
rect 1984 10240 2016 10272
rect 2056 10240 2088 10272
rect 2128 10240 2160 10272
rect 2200 10240 2232 10272
rect 2272 10240 2304 10272
rect 2344 10240 2376 10272
rect 2416 10240 2448 10272
rect 2488 10240 2520 10272
rect 2560 10240 2592 10272
rect 2632 10240 2664 10272
rect 2704 10240 2736 10272
rect 2776 10240 2808 10272
rect 2848 10240 2880 10272
rect 2920 10240 2952 10272
rect 2992 10240 3024 10272
rect 3064 10240 3096 10272
rect 3136 10240 3168 10272
rect 3208 10240 3240 10272
rect 3280 10240 3312 10272
rect 3352 10240 3384 10272
rect 3424 10240 3456 10272
rect 3496 10240 3528 10272
rect 3568 10240 3600 10272
rect 3640 10240 3672 10272
rect 3712 10240 3744 10272
rect 3784 10240 3816 10272
rect 3856 10240 3888 10272
rect 3928 10240 3960 10272
rect 40 10168 72 10200
rect 112 10168 144 10200
rect 184 10168 216 10200
rect 256 10168 288 10200
rect 328 10168 360 10200
rect 400 10168 432 10200
rect 472 10168 504 10200
rect 544 10168 576 10200
rect 616 10168 648 10200
rect 688 10168 720 10200
rect 760 10168 792 10200
rect 832 10168 864 10200
rect 904 10168 936 10200
rect 976 10168 1008 10200
rect 1048 10168 1080 10200
rect 1120 10168 1152 10200
rect 1192 10168 1224 10200
rect 1264 10168 1296 10200
rect 1336 10168 1368 10200
rect 1408 10168 1440 10200
rect 1480 10168 1512 10200
rect 1552 10168 1584 10200
rect 1624 10168 1656 10200
rect 1696 10168 1728 10200
rect 1768 10168 1800 10200
rect 1840 10168 1872 10200
rect 1912 10168 1944 10200
rect 1984 10168 2016 10200
rect 2056 10168 2088 10200
rect 2128 10168 2160 10200
rect 2200 10168 2232 10200
rect 2272 10168 2304 10200
rect 2344 10168 2376 10200
rect 2416 10168 2448 10200
rect 2488 10168 2520 10200
rect 2560 10168 2592 10200
rect 2632 10168 2664 10200
rect 2704 10168 2736 10200
rect 2776 10168 2808 10200
rect 2848 10168 2880 10200
rect 2920 10168 2952 10200
rect 2992 10168 3024 10200
rect 3064 10168 3096 10200
rect 3136 10168 3168 10200
rect 3208 10168 3240 10200
rect 3280 10168 3312 10200
rect 3352 10168 3384 10200
rect 3424 10168 3456 10200
rect 3496 10168 3528 10200
rect 3568 10168 3600 10200
rect 3640 10168 3672 10200
rect 3712 10168 3744 10200
rect 3784 10168 3816 10200
rect 3856 10168 3888 10200
rect 3928 10168 3960 10200
rect 40 10096 72 10128
rect 112 10096 144 10128
rect 184 10096 216 10128
rect 256 10096 288 10128
rect 328 10096 360 10128
rect 400 10096 432 10128
rect 472 10096 504 10128
rect 544 10096 576 10128
rect 616 10096 648 10128
rect 688 10096 720 10128
rect 760 10096 792 10128
rect 832 10096 864 10128
rect 904 10096 936 10128
rect 976 10096 1008 10128
rect 1048 10096 1080 10128
rect 1120 10096 1152 10128
rect 1192 10096 1224 10128
rect 1264 10096 1296 10128
rect 1336 10096 1368 10128
rect 1408 10096 1440 10128
rect 1480 10096 1512 10128
rect 1552 10096 1584 10128
rect 1624 10096 1656 10128
rect 1696 10096 1728 10128
rect 1768 10096 1800 10128
rect 1840 10096 1872 10128
rect 1912 10096 1944 10128
rect 1984 10096 2016 10128
rect 2056 10096 2088 10128
rect 2128 10096 2160 10128
rect 2200 10096 2232 10128
rect 2272 10096 2304 10128
rect 2344 10096 2376 10128
rect 2416 10096 2448 10128
rect 2488 10096 2520 10128
rect 2560 10096 2592 10128
rect 2632 10096 2664 10128
rect 2704 10096 2736 10128
rect 2776 10096 2808 10128
rect 2848 10096 2880 10128
rect 2920 10096 2952 10128
rect 2992 10096 3024 10128
rect 3064 10096 3096 10128
rect 3136 10096 3168 10128
rect 3208 10096 3240 10128
rect 3280 10096 3312 10128
rect 3352 10096 3384 10128
rect 3424 10096 3456 10128
rect 3496 10096 3528 10128
rect 3568 10096 3600 10128
rect 3640 10096 3672 10128
rect 3712 10096 3744 10128
rect 3784 10096 3816 10128
rect 3856 10096 3888 10128
rect 3928 10096 3960 10128
rect 40 10024 72 10056
rect 112 10024 144 10056
rect 184 10024 216 10056
rect 256 10024 288 10056
rect 328 10024 360 10056
rect 400 10024 432 10056
rect 472 10024 504 10056
rect 544 10024 576 10056
rect 616 10024 648 10056
rect 688 10024 720 10056
rect 760 10024 792 10056
rect 832 10024 864 10056
rect 904 10024 936 10056
rect 976 10024 1008 10056
rect 1048 10024 1080 10056
rect 1120 10024 1152 10056
rect 1192 10024 1224 10056
rect 1264 10024 1296 10056
rect 1336 10024 1368 10056
rect 1408 10024 1440 10056
rect 1480 10024 1512 10056
rect 1552 10024 1584 10056
rect 1624 10024 1656 10056
rect 1696 10024 1728 10056
rect 1768 10024 1800 10056
rect 1840 10024 1872 10056
rect 1912 10024 1944 10056
rect 1984 10024 2016 10056
rect 2056 10024 2088 10056
rect 2128 10024 2160 10056
rect 2200 10024 2232 10056
rect 2272 10024 2304 10056
rect 2344 10024 2376 10056
rect 2416 10024 2448 10056
rect 2488 10024 2520 10056
rect 2560 10024 2592 10056
rect 2632 10024 2664 10056
rect 2704 10024 2736 10056
rect 2776 10024 2808 10056
rect 2848 10024 2880 10056
rect 2920 10024 2952 10056
rect 2992 10024 3024 10056
rect 3064 10024 3096 10056
rect 3136 10024 3168 10056
rect 3208 10024 3240 10056
rect 3280 10024 3312 10056
rect 3352 10024 3384 10056
rect 3424 10024 3456 10056
rect 3496 10024 3528 10056
rect 3568 10024 3600 10056
rect 3640 10024 3672 10056
rect 3712 10024 3744 10056
rect 3784 10024 3816 10056
rect 3856 10024 3888 10056
rect 3928 10024 3960 10056
rect 40 9952 72 9984
rect 112 9952 144 9984
rect 184 9952 216 9984
rect 256 9952 288 9984
rect 328 9952 360 9984
rect 400 9952 432 9984
rect 472 9952 504 9984
rect 544 9952 576 9984
rect 616 9952 648 9984
rect 688 9952 720 9984
rect 760 9952 792 9984
rect 832 9952 864 9984
rect 904 9952 936 9984
rect 976 9952 1008 9984
rect 1048 9952 1080 9984
rect 1120 9952 1152 9984
rect 1192 9952 1224 9984
rect 1264 9952 1296 9984
rect 1336 9952 1368 9984
rect 1408 9952 1440 9984
rect 1480 9952 1512 9984
rect 1552 9952 1584 9984
rect 1624 9952 1656 9984
rect 1696 9952 1728 9984
rect 1768 9952 1800 9984
rect 1840 9952 1872 9984
rect 1912 9952 1944 9984
rect 1984 9952 2016 9984
rect 2056 9952 2088 9984
rect 2128 9952 2160 9984
rect 2200 9952 2232 9984
rect 2272 9952 2304 9984
rect 2344 9952 2376 9984
rect 2416 9952 2448 9984
rect 2488 9952 2520 9984
rect 2560 9952 2592 9984
rect 2632 9952 2664 9984
rect 2704 9952 2736 9984
rect 2776 9952 2808 9984
rect 2848 9952 2880 9984
rect 2920 9952 2952 9984
rect 2992 9952 3024 9984
rect 3064 9952 3096 9984
rect 3136 9952 3168 9984
rect 3208 9952 3240 9984
rect 3280 9952 3312 9984
rect 3352 9952 3384 9984
rect 3424 9952 3456 9984
rect 3496 9952 3528 9984
rect 3568 9952 3600 9984
rect 3640 9952 3672 9984
rect 3712 9952 3744 9984
rect 3784 9952 3816 9984
rect 3856 9952 3888 9984
rect 3928 9952 3960 9984
rect 40 9880 72 9912
rect 112 9880 144 9912
rect 184 9880 216 9912
rect 256 9880 288 9912
rect 328 9880 360 9912
rect 400 9880 432 9912
rect 472 9880 504 9912
rect 544 9880 576 9912
rect 616 9880 648 9912
rect 688 9880 720 9912
rect 760 9880 792 9912
rect 832 9880 864 9912
rect 904 9880 936 9912
rect 976 9880 1008 9912
rect 1048 9880 1080 9912
rect 1120 9880 1152 9912
rect 1192 9880 1224 9912
rect 1264 9880 1296 9912
rect 1336 9880 1368 9912
rect 1408 9880 1440 9912
rect 1480 9880 1512 9912
rect 1552 9880 1584 9912
rect 1624 9880 1656 9912
rect 1696 9880 1728 9912
rect 1768 9880 1800 9912
rect 1840 9880 1872 9912
rect 1912 9880 1944 9912
rect 1984 9880 2016 9912
rect 2056 9880 2088 9912
rect 2128 9880 2160 9912
rect 2200 9880 2232 9912
rect 2272 9880 2304 9912
rect 2344 9880 2376 9912
rect 2416 9880 2448 9912
rect 2488 9880 2520 9912
rect 2560 9880 2592 9912
rect 2632 9880 2664 9912
rect 2704 9880 2736 9912
rect 2776 9880 2808 9912
rect 2848 9880 2880 9912
rect 2920 9880 2952 9912
rect 2992 9880 3024 9912
rect 3064 9880 3096 9912
rect 3136 9880 3168 9912
rect 3208 9880 3240 9912
rect 3280 9880 3312 9912
rect 3352 9880 3384 9912
rect 3424 9880 3456 9912
rect 3496 9880 3528 9912
rect 3568 9880 3600 9912
rect 3640 9880 3672 9912
rect 3712 9880 3744 9912
rect 3784 9880 3816 9912
rect 3856 9880 3888 9912
rect 3928 9880 3960 9912
rect 40 9808 72 9840
rect 112 9808 144 9840
rect 184 9808 216 9840
rect 256 9808 288 9840
rect 328 9808 360 9840
rect 400 9808 432 9840
rect 472 9808 504 9840
rect 544 9808 576 9840
rect 616 9808 648 9840
rect 688 9808 720 9840
rect 760 9808 792 9840
rect 832 9808 864 9840
rect 904 9808 936 9840
rect 976 9808 1008 9840
rect 1048 9808 1080 9840
rect 1120 9808 1152 9840
rect 1192 9808 1224 9840
rect 1264 9808 1296 9840
rect 1336 9808 1368 9840
rect 1408 9808 1440 9840
rect 1480 9808 1512 9840
rect 1552 9808 1584 9840
rect 1624 9808 1656 9840
rect 1696 9808 1728 9840
rect 1768 9808 1800 9840
rect 1840 9808 1872 9840
rect 1912 9808 1944 9840
rect 1984 9808 2016 9840
rect 2056 9808 2088 9840
rect 2128 9808 2160 9840
rect 2200 9808 2232 9840
rect 2272 9808 2304 9840
rect 2344 9808 2376 9840
rect 2416 9808 2448 9840
rect 2488 9808 2520 9840
rect 2560 9808 2592 9840
rect 2632 9808 2664 9840
rect 2704 9808 2736 9840
rect 2776 9808 2808 9840
rect 2848 9808 2880 9840
rect 2920 9808 2952 9840
rect 2992 9808 3024 9840
rect 3064 9808 3096 9840
rect 3136 9808 3168 9840
rect 3208 9808 3240 9840
rect 3280 9808 3312 9840
rect 3352 9808 3384 9840
rect 3424 9808 3456 9840
rect 3496 9808 3528 9840
rect 3568 9808 3600 9840
rect 3640 9808 3672 9840
rect 3712 9808 3744 9840
rect 3784 9808 3816 9840
rect 3856 9808 3888 9840
rect 3928 9808 3960 9840
rect 40 9736 72 9768
rect 112 9736 144 9768
rect 184 9736 216 9768
rect 256 9736 288 9768
rect 328 9736 360 9768
rect 400 9736 432 9768
rect 472 9736 504 9768
rect 544 9736 576 9768
rect 616 9736 648 9768
rect 688 9736 720 9768
rect 760 9736 792 9768
rect 832 9736 864 9768
rect 904 9736 936 9768
rect 976 9736 1008 9768
rect 1048 9736 1080 9768
rect 1120 9736 1152 9768
rect 1192 9736 1224 9768
rect 1264 9736 1296 9768
rect 1336 9736 1368 9768
rect 1408 9736 1440 9768
rect 1480 9736 1512 9768
rect 1552 9736 1584 9768
rect 1624 9736 1656 9768
rect 1696 9736 1728 9768
rect 1768 9736 1800 9768
rect 1840 9736 1872 9768
rect 1912 9736 1944 9768
rect 1984 9736 2016 9768
rect 2056 9736 2088 9768
rect 2128 9736 2160 9768
rect 2200 9736 2232 9768
rect 2272 9736 2304 9768
rect 2344 9736 2376 9768
rect 2416 9736 2448 9768
rect 2488 9736 2520 9768
rect 2560 9736 2592 9768
rect 2632 9736 2664 9768
rect 2704 9736 2736 9768
rect 2776 9736 2808 9768
rect 2848 9736 2880 9768
rect 2920 9736 2952 9768
rect 2992 9736 3024 9768
rect 3064 9736 3096 9768
rect 3136 9736 3168 9768
rect 3208 9736 3240 9768
rect 3280 9736 3312 9768
rect 3352 9736 3384 9768
rect 3424 9736 3456 9768
rect 3496 9736 3528 9768
rect 3568 9736 3600 9768
rect 3640 9736 3672 9768
rect 3712 9736 3744 9768
rect 3784 9736 3816 9768
rect 3856 9736 3888 9768
rect 3928 9736 3960 9768
rect 40 9664 72 9696
rect 112 9664 144 9696
rect 184 9664 216 9696
rect 256 9664 288 9696
rect 328 9664 360 9696
rect 400 9664 432 9696
rect 472 9664 504 9696
rect 544 9664 576 9696
rect 616 9664 648 9696
rect 688 9664 720 9696
rect 760 9664 792 9696
rect 832 9664 864 9696
rect 904 9664 936 9696
rect 976 9664 1008 9696
rect 1048 9664 1080 9696
rect 1120 9664 1152 9696
rect 1192 9664 1224 9696
rect 1264 9664 1296 9696
rect 1336 9664 1368 9696
rect 1408 9664 1440 9696
rect 1480 9664 1512 9696
rect 1552 9664 1584 9696
rect 1624 9664 1656 9696
rect 1696 9664 1728 9696
rect 1768 9664 1800 9696
rect 1840 9664 1872 9696
rect 1912 9664 1944 9696
rect 1984 9664 2016 9696
rect 2056 9664 2088 9696
rect 2128 9664 2160 9696
rect 2200 9664 2232 9696
rect 2272 9664 2304 9696
rect 2344 9664 2376 9696
rect 2416 9664 2448 9696
rect 2488 9664 2520 9696
rect 2560 9664 2592 9696
rect 2632 9664 2664 9696
rect 2704 9664 2736 9696
rect 2776 9664 2808 9696
rect 2848 9664 2880 9696
rect 2920 9664 2952 9696
rect 2992 9664 3024 9696
rect 3064 9664 3096 9696
rect 3136 9664 3168 9696
rect 3208 9664 3240 9696
rect 3280 9664 3312 9696
rect 3352 9664 3384 9696
rect 3424 9664 3456 9696
rect 3496 9664 3528 9696
rect 3568 9664 3600 9696
rect 3640 9664 3672 9696
rect 3712 9664 3744 9696
rect 3784 9664 3816 9696
rect 3856 9664 3888 9696
rect 3928 9664 3960 9696
rect 40 9592 72 9624
rect 112 9592 144 9624
rect 184 9592 216 9624
rect 256 9592 288 9624
rect 328 9592 360 9624
rect 400 9592 432 9624
rect 472 9592 504 9624
rect 544 9592 576 9624
rect 616 9592 648 9624
rect 688 9592 720 9624
rect 760 9592 792 9624
rect 832 9592 864 9624
rect 904 9592 936 9624
rect 976 9592 1008 9624
rect 1048 9592 1080 9624
rect 1120 9592 1152 9624
rect 1192 9592 1224 9624
rect 1264 9592 1296 9624
rect 1336 9592 1368 9624
rect 1408 9592 1440 9624
rect 1480 9592 1512 9624
rect 1552 9592 1584 9624
rect 1624 9592 1656 9624
rect 1696 9592 1728 9624
rect 1768 9592 1800 9624
rect 1840 9592 1872 9624
rect 1912 9592 1944 9624
rect 1984 9592 2016 9624
rect 2056 9592 2088 9624
rect 2128 9592 2160 9624
rect 2200 9592 2232 9624
rect 2272 9592 2304 9624
rect 2344 9592 2376 9624
rect 2416 9592 2448 9624
rect 2488 9592 2520 9624
rect 2560 9592 2592 9624
rect 2632 9592 2664 9624
rect 2704 9592 2736 9624
rect 2776 9592 2808 9624
rect 2848 9592 2880 9624
rect 2920 9592 2952 9624
rect 2992 9592 3024 9624
rect 3064 9592 3096 9624
rect 3136 9592 3168 9624
rect 3208 9592 3240 9624
rect 3280 9592 3312 9624
rect 3352 9592 3384 9624
rect 3424 9592 3456 9624
rect 3496 9592 3528 9624
rect 3568 9592 3600 9624
rect 3640 9592 3672 9624
rect 3712 9592 3744 9624
rect 3784 9592 3816 9624
rect 3856 9592 3888 9624
rect 3928 9592 3960 9624
rect 40 9520 72 9552
rect 112 9520 144 9552
rect 184 9520 216 9552
rect 256 9520 288 9552
rect 328 9520 360 9552
rect 400 9520 432 9552
rect 472 9520 504 9552
rect 544 9520 576 9552
rect 616 9520 648 9552
rect 688 9520 720 9552
rect 760 9520 792 9552
rect 832 9520 864 9552
rect 904 9520 936 9552
rect 976 9520 1008 9552
rect 1048 9520 1080 9552
rect 1120 9520 1152 9552
rect 1192 9520 1224 9552
rect 1264 9520 1296 9552
rect 1336 9520 1368 9552
rect 1408 9520 1440 9552
rect 1480 9520 1512 9552
rect 1552 9520 1584 9552
rect 1624 9520 1656 9552
rect 1696 9520 1728 9552
rect 1768 9520 1800 9552
rect 1840 9520 1872 9552
rect 1912 9520 1944 9552
rect 1984 9520 2016 9552
rect 2056 9520 2088 9552
rect 2128 9520 2160 9552
rect 2200 9520 2232 9552
rect 2272 9520 2304 9552
rect 2344 9520 2376 9552
rect 2416 9520 2448 9552
rect 2488 9520 2520 9552
rect 2560 9520 2592 9552
rect 2632 9520 2664 9552
rect 2704 9520 2736 9552
rect 2776 9520 2808 9552
rect 2848 9520 2880 9552
rect 2920 9520 2952 9552
rect 2992 9520 3024 9552
rect 3064 9520 3096 9552
rect 3136 9520 3168 9552
rect 3208 9520 3240 9552
rect 3280 9520 3312 9552
rect 3352 9520 3384 9552
rect 3424 9520 3456 9552
rect 3496 9520 3528 9552
rect 3568 9520 3600 9552
rect 3640 9520 3672 9552
rect 3712 9520 3744 9552
rect 3784 9520 3816 9552
rect 3856 9520 3888 9552
rect 3928 9520 3960 9552
rect 40 9448 72 9480
rect 112 9448 144 9480
rect 184 9448 216 9480
rect 256 9448 288 9480
rect 328 9448 360 9480
rect 400 9448 432 9480
rect 472 9448 504 9480
rect 544 9448 576 9480
rect 616 9448 648 9480
rect 688 9448 720 9480
rect 760 9448 792 9480
rect 832 9448 864 9480
rect 904 9448 936 9480
rect 976 9448 1008 9480
rect 1048 9448 1080 9480
rect 1120 9448 1152 9480
rect 1192 9448 1224 9480
rect 1264 9448 1296 9480
rect 1336 9448 1368 9480
rect 1408 9448 1440 9480
rect 1480 9448 1512 9480
rect 1552 9448 1584 9480
rect 1624 9448 1656 9480
rect 1696 9448 1728 9480
rect 1768 9448 1800 9480
rect 1840 9448 1872 9480
rect 1912 9448 1944 9480
rect 1984 9448 2016 9480
rect 2056 9448 2088 9480
rect 2128 9448 2160 9480
rect 2200 9448 2232 9480
rect 2272 9448 2304 9480
rect 2344 9448 2376 9480
rect 2416 9448 2448 9480
rect 2488 9448 2520 9480
rect 2560 9448 2592 9480
rect 2632 9448 2664 9480
rect 2704 9448 2736 9480
rect 2776 9448 2808 9480
rect 2848 9448 2880 9480
rect 2920 9448 2952 9480
rect 2992 9448 3024 9480
rect 3064 9448 3096 9480
rect 3136 9448 3168 9480
rect 3208 9448 3240 9480
rect 3280 9448 3312 9480
rect 3352 9448 3384 9480
rect 3424 9448 3456 9480
rect 3496 9448 3528 9480
rect 3568 9448 3600 9480
rect 3640 9448 3672 9480
rect 3712 9448 3744 9480
rect 3784 9448 3816 9480
rect 3856 9448 3888 9480
rect 3928 9448 3960 9480
rect 40 9376 72 9408
rect 112 9376 144 9408
rect 184 9376 216 9408
rect 256 9376 288 9408
rect 328 9376 360 9408
rect 400 9376 432 9408
rect 472 9376 504 9408
rect 544 9376 576 9408
rect 616 9376 648 9408
rect 688 9376 720 9408
rect 760 9376 792 9408
rect 832 9376 864 9408
rect 904 9376 936 9408
rect 976 9376 1008 9408
rect 1048 9376 1080 9408
rect 1120 9376 1152 9408
rect 1192 9376 1224 9408
rect 1264 9376 1296 9408
rect 1336 9376 1368 9408
rect 1408 9376 1440 9408
rect 1480 9376 1512 9408
rect 1552 9376 1584 9408
rect 1624 9376 1656 9408
rect 1696 9376 1728 9408
rect 1768 9376 1800 9408
rect 1840 9376 1872 9408
rect 1912 9376 1944 9408
rect 1984 9376 2016 9408
rect 2056 9376 2088 9408
rect 2128 9376 2160 9408
rect 2200 9376 2232 9408
rect 2272 9376 2304 9408
rect 2344 9376 2376 9408
rect 2416 9376 2448 9408
rect 2488 9376 2520 9408
rect 2560 9376 2592 9408
rect 2632 9376 2664 9408
rect 2704 9376 2736 9408
rect 2776 9376 2808 9408
rect 2848 9376 2880 9408
rect 2920 9376 2952 9408
rect 2992 9376 3024 9408
rect 3064 9376 3096 9408
rect 3136 9376 3168 9408
rect 3208 9376 3240 9408
rect 3280 9376 3312 9408
rect 3352 9376 3384 9408
rect 3424 9376 3456 9408
rect 3496 9376 3528 9408
rect 3568 9376 3600 9408
rect 3640 9376 3672 9408
rect 3712 9376 3744 9408
rect 3784 9376 3816 9408
rect 3856 9376 3888 9408
rect 3928 9376 3960 9408
rect 40 9304 72 9336
rect 112 9304 144 9336
rect 184 9304 216 9336
rect 256 9304 288 9336
rect 328 9304 360 9336
rect 400 9304 432 9336
rect 472 9304 504 9336
rect 544 9304 576 9336
rect 616 9304 648 9336
rect 688 9304 720 9336
rect 760 9304 792 9336
rect 832 9304 864 9336
rect 904 9304 936 9336
rect 976 9304 1008 9336
rect 1048 9304 1080 9336
rect 1120 9304 1152 9336
rect 1192 9304 1224 9336
rect 1264 9304 1296 9336
rect 1336 9304 1368 9336
rect 1408 9304 1440 9336
rect 1480 9304 1512 9336
rect 1552 9304 1584 9336
rect 1624 9304 1656 9336
rect 1696 9304 1728 9336
rect 1768 9304 1800 9336
rect 1840 9304 1872 9336
rect 1912 9304 1944 9336
rect 1984 9304 2016 9336
rect 2056 9304 2088 9336
rect 2128 9304 2160 9336
rect 2200 9304 2232 9336
rect 2272 9304 2304 9336
rect 2344 9304 2376 9336
rect 2416 9304 2448 9336
rect 2488 9304 2520 9336
rect 2560 9304 2592 9336
rect 2632 9304 2664 9336
rect 2704 9304 2736 9336
rect 2776 9304 2808 9336
rect 2848 9304 2880 9336
rect 2920 9304 2952 9336
rect 2992 9304 3024 9336
rect 3064 9304 3096 9336
rect 3136 9304 3168 9336
rect 3208 9304 3240 9336
rect 3280 9304 3312 9336
rect 3352 9304 3384 9336
rect 3424 9304 3456 9336
rect 3496 9304 3528 9336
rect 3568 9304 3600 9336
rect 3640 9304 3672 9336
rect 3712 9304 3744 9336
rect 3784 9304 3816 9336
rect 3856 9304 3888 9336
rect 3928 9304 3960 9336
rect 40 9232 72 9264
rect 112 9232 144 9264
rect 184 9232 216 9264
rect 256 9232 288 9264
rect 328 9232 360 9264
rect 400 9232 432 9264
rect 472 9232 504 9264
rect 544 9232 576 9264
rect 616 9232 648 9264
rect 688 9232 720 9264
rect 760 9232 792 9264
rect 832 9232 864 9264
rect 904 9232 936 9264
rect 976 9232 1008 9264
rect 1048 9232 1080 9264
rect 1120 9232 1152 9264
rect 1192 9232 1224 9264
rect 1264 9232 1296 9264
rect 1336 9232 1368 9264
rect 1408 9232 1440 9264
rect 1480 9232 1512 9264
rect 1552 9232 1584 9264
rect 1624 9232 1656 9264
rect 1696 9232 1728 9264
rect 1768 9232 1800 9264
rect 1840 9232 1872 9264
rect 1912 9232 1944 9264
rect 1984 9232 2016 9264
rect 2056 9232 2088 9264
rect 2128 9232 2160 9264
rect 2200 9232 2232 9264
rect 2272 9232 2304 9264
rect 2344 9232 2376 9264
rect 2416 9232 2448 9264
rect 2488 9232 2520 9264
rect 2560 9232 2592 9264
rect 2632 9232 2664 9264
rect 2704 9232 2736 9264
rect 2776 9232 2808 9264
rect 2848 9232 2880 9264
rect 2920 9232 2952 9264
rect 2992 9232 3024 9264
rect 3064 9232 3096 9264
rect 3136 9232 3168 9264
rect 3208 9232 3240 9264
rect 3280 9232 3312 9264
rect 3352 9232 3384 9264
rect 3424 9232 3456 9264
rect 3496 9232 3528 9264
rect 3568 9232 3600 9264
rect 3640 9232 3672 9264
rect 3712 9232 3744 9264
rect 3784 9232 3816 9264
rect 3856 9232 3888 9264
rect 3928 9232 3960 9264
rect 40 9160 72 9192
rect 112 9160 144 9192
rect 184 9160 216 9192
rect 256 9160 288 9192
rect 328 9160 360 9192
rect 400 9160 432 9192
rect 472 9160 504 9192
rect 544 9160 576 9192
rect 616 9160 648 9192
rect 688 9160 720 9192
rect 760 9160 792 9192
rect 832 9160 864 9192
rect 904 9160 936 9192
rect 976 9160 1008 9192
rect 1048 9160 1080 9192
rect 1120 9160 1152 9192
rect 1192 9160 1224 9192
rect 1264 9160 1296 9192
rect 1336 9160 1368 9192
rect 1408 9160 1440 9192
rect 1480 9160 1512 9192
rect 1552 9160 1584 9192
rect 1624 9160 1656 9192
rect 1696 9160 1728 9192
rect 1768 9160 1800 9192
rect 1840 9160 1872 9192
rect 1912 9160 1944 9192
rect 1984 9160 2016 9192
rect 2056 9160 2088 9192
rect 2128 9160 2160 9192
rect 2200 9160 2232 9192
rect 2272 9160 2304 9192
rect 2344 9160 2376 9192
rect 2416 9160 2448 9192
rect 2488 9160 2520 9192
rect 2560 9160 2592 9192
rect 2632 9160 2664 9192
rect 2704 9160 2736 9192
rect 2776 9160 2808 9192
rect 2848 9160 2880 9192
rect 2920 9160 2952 9192
rect 2992 9160 3024 9192
rect 3064 9160 3096 9192
rect 3136 9160 3168 9192
rect 3208 9160 3240 9192
rect 3280 9160 3312 9192
rect 3352 9160 3384 9192
rect 3424 9160 3456 9192
rect 3496 9160 3528 9192
rect 3568 9160 3600 9192
rect 3640 9160 3672 9192
rect 3712 9160 3744 9192
rect 3784 9160 3816 9192
rect 3856 9160 3888 9192
rect 3928 9160 3960 9192
rect 40 9088 72 9120
rect 112 9088 144 9120
rect 184 9088 216 9120
rect 256 9088 288 9120
rect 328 9088 360 9120
rect 400 9088 432 9120
rect 472 9088 504 9120
rect 544 9088 576 9120
rect 616 9088 648 9120
rect 688 9088 720 9120
rect 760 9088 792 9120
rect 832 9088 864 9120
rect 904 9088 936 9120
rect 976 9088 1008 9120
rect 1048 9088 1080 9120
rect 1120 9088 1152 9120
rect 1192 9088 1224 9120
rect 1264 9088 1296 9120
rect 1336 9088 1368 9120
rect 1408 9088 1440 9120
rect 1480 9088 1512 9120
rect 1552 9088 1584 9120
rect 1624 9088 1656 9120
rect 1696 9088 1728 9120
rect 1768 9088 1800 9120
rect 1840 9088 1872 9120
rect 1912 9088 1944 9120
rect 1984 9088 2016 9120
rect 2056 9088 2088 9120
rect 2128 9088 2160 9120
rect 2200 9088 2232 9120
rect 2272 9088 2304 9120
rect 2344 9088 2376 9120
rect 2416 9088 2448 9120
rect 2488 9088 2520 9120
rect 2560 9088 2592 9120
rect 2632 9088 2664 9120
rect 2704 9088 2736 9120
rect 2776 9088 2808 9120
rect 2848 9088 2880 9120
rect 2920 9088 2952 9120
rect 2992 9088 3024 9120
rect 3064 9088 3096 9120
rect 3136 9088 3168 9120
rect 3208 9088 3240 9120
rect 3280 9088 3312 9120
rect 3352 9088 3384 9120
rect 3424 9088 3456 9120
rect 3496 9088 3528 9120
rect 3568 9088 3600 9120
rect 3640 9088 3672 9120
rect 3712 9088 3744 9120
rect 3784 9088 3816 9120
rect 3856 9088 3888 9120
rect 3928 9088 3960 9120
rect 40 9016 72 9048
rect 112 9016 144 9048
rect 184 9016 216 9048
rect 256 9016 288 9048
rect 328 9016 360 9048
rect 400 9016 432 9048
rect 472 9016 504 9048
rect 544 9016 576 9048
rect 616 9016 648 9048
rect 688 9016 720 9048
rect 760 9016 792 9048
rect 832 9016 864 9048
rect 904 9016 936 9048
rect 976 9016 1008 9048
rect 1048 9016 1080 9048
rect 1120 9016 1152 9048
rect 1192 9016 1224 9048
rect 1264 9016 1296 9048
rect 1336 9016 1368 9048
rect 1408 9016 1440 9048
rect 1480 9016 1512 9048
rect 1552 9016 1584 9048
rect 1624 9016 1656 9048
rect 1696 9016 1728 9048
rect 1768 9016 1800 9048
rect 1840 9016 1872 9048
rect 1912 9016 1944 9048
rect 1984 9016 2016 9048
rect 2056 9016 2088 9048
rect 2128 9016 2160 9048
rect 2200 9016 2232 9048
rect 2272 9016 2304 9048
rect 2344 9016 2376 9048
rect 2416 9016 2448 9048
rect 2488 9016 2520 9048
rect 2560 9016 2592 9048
rect 2632 9016 2664 9048
rect 2704 9016 2736 9048
rect 2776 9016 2808 9048
rect 2848 9016 2880 9048
rect 2920 9016 2952 9048
rect 2992 9016 3024 9048
rect 3064 9016 3096 9048
rect 3136 9016 3168 9048
rect 3208 9016 3240 9048
rect 3280 9016 3312 9048
rect 3352 9016 3384 9048
rect 3424 9016 3456 9048
rect 3496 9016 3528 9048
rect 3568 9016 3600 9048
rect 3640 9016 3672 9048
rect 3712 9016 3744 9048
rect 3784 9016 3816 9048
rect 3856 9016 3888 9048
rect 3928 9016 3960 9048
rect 40 8944 72 8976
rect 112 8944 144 8976
rect 184 8944 216 8976
rect 256 8944 288 8976
rect 328 8944 360 8976
rect 400 8944 432 8976
rect 472 8944 504 8976
rect 544 8944 576 8976
rect 616 8944 648 8976
rect 688 8944 720 8976
rect 760 8944 792 8976
rect 832 8944 864 8976
rect 904 8944 936 8976
rect 976 8944 1008 8976
rect 1048 8944 1080 8976
rect 1120 8944 1152 8976
rect 1192 8944 1224 8976
rect 1264 8944 1296 8976
rect 1336 8944 1368 8976
rect 1408 8944 1440 8976
rect 1480 8944 1512 8976
rect 1552 8944 1584 8976
rect 1624 8944 1656 8976
rect 1696 8944 1728 8976
rect 1768 8944 1800 8976
rect 1840 8944 1872 8976
rect 1912 8944 1944 8976
rect 1984 8944 2016 8976
rect 2056 8944 2088 8976
rect 2128 8944 2160 8976
rect 2200 8944 2232 8976
rect 2272 8944 2304 8976
rect 2344 8944 2376 8976
rect 2416 8944 2448 8976
rect 2488 8944 2520 8976
rect 2560 8944 2592 8976
rect 2632 8944 2664 8976
rect 2704 8944 2736 8976
rect 2776 8944 2808 8976
rect 2848 8944 2880 8976
rect 2920 8944 2952 8976
rect 2992 8944 3024 8976
rect 3064 8944 3096 8976
rect 3136 8944 3168 8976
rect 3208 8944 3240 8976
rect 3280 8944 3312 8976
rect 3352 8944 3384 8976
rect 3424 8944 3456 8976
rect 3496 8944 3528 8976
rect 3568 8944 3600 8976
rect 3640 8944 3672 8976
rect 3712 8944 3744 8976
rect 3784 8944 3816 8976
rect 3856 8944 3888 8976
rect 3928 8944 3960 8976
rect 40 8872 72 8904
rect 112 8872 144 8904
rect 184 8872 216 8904
rect 256 8872 288 8904
rect 328 8872 360 8904
rect 400 8872 432 8904
rect 472 8872 504 8904
rect 544 8872 576 8904
rect 616 8872 648 8904
rect 688 8872 720 8904
rect 760 8872 792 8904
rect 832 8872 864 8904
rect 904 8872 936 8904
rect 976 8872 1008 8904
rect 1048 8872 1080 8904
rect 1120 8872 1152 8904
rect 1192 8872 1224 8904
rect 1264 8872 1296 8904
rect 1336 8872 1368 8904
rect 1408 8872 1440 8904
rect 1480 8872 1512 8904
rect 1552 8872 1584 8904
rect 1624 8872 1656 8904
rect 1696 8872 1728 8904
rect 1768 8872 1800 8904
rect 1840 8872 1872 8904
rect 1912 8872 1944 8904
rect 1984 8872 2016 8904
rect 2056 8872 2088 8904
rect 2128 8872 2160 8904
rect 2200 8872 2232 8904
rect 2272 8872 2304 8904
rect 2344 8872 2376 8904
rect 2416 8872 2448 8904
rect 2488 8872 2520 8904
rect 2560 8872 2592 8904
rect 2632 8872 2664 8904
rect 2704 8872 2736 8904
rect 2776 8872 2808 8904
rect 2848 8872 2880 8904
rect 2920 8872 2952 8904
rect 2992 8872 3024 8904
rect 3064 8872 3096 8904
rect 3136 8872 3168 8904
rect 3208 8872 3240 8904
rect 3280 8872 3312 8904
rect 3352 8872 3384 8904
rect 3424 8872 3456 8904
rect 3496 8872 3528 8904
rect 3568 8872 3600 8904
rect 3640 8872 3672 8904
rect 3712 8872 3744 8904
rect 3784 8872 3816 8904
rect 3856 8872 3888 8904
rect 3928 8872 3960 8904
rect 40 8800 72 8832
rect 112 8800 144 8832
rect 184 8800 216 8832
rect 256 8800 288 8832
rect 328 8800 360 8832
rect 400 8800 432 8832
rect 472 8800 504 8832
rect 544 8800 576 8832
rect 616 8800 648 8832
rect 688 8800 720 8832
rect 760 8800 792 8832
rect 832 8800 864 8832
rect 904 8800 936 8832
rect 976 8800 1008 8832
rect 1048 8800 1080 8832
rect 1120 8800 1152 8832
rect 1192 8800 1224 8832
rect 1264 8800 1296 8832
rect 1336 8800 1368 8832
rect 1408 8800 1440 8832
rect 1480 8800 1512 8832
rect 1552 8800 1584 8832
rect 1624 8800 1656 8832
rect 1696 8800 1728 8832
rect 1768 8800 1800 8832
rect 1840 8800 1872 8832
rect 1912 8800 1944 8832
rect 1984 8800 2016 8832
rect 2056 8800 2088 8832
rect 2128 8800 2160 8832
rect 2200 8800 2232 8832
rect 2272 8800 2304 8832
rect 2344 8800 2376 8832
rect 2416 8800 2448 8832
rect 2488 8800 2520 8832
rect 2560 8800 2592 8832
rect 2632 8800 2664 8832
rect 2704 8800 2736 8832
rect 2776 8800 2808 8832
rect 2848 8800 2880 8832
rect 2920 8800 2952 8832
rect 2992 8800 3024 8832
rect 3064 8800 3096 8832
rect 3136 8800 3168 8832
rect 3208 8800 3240 8832
rect 3280 8800 3312 8832
rect 3352 8800 3384 8832
rect 3424 8800 3456 8832
rect 3496 8800 3528 8832
rect 3568 8800 3600 8832
rect 3640 8800 3672 8832
rect 3712 8800 3744 8832
rect 3784 8800 3816 8832
rect 3856 8800 3888 8832
rect 3928 8800 3960 8832
rect 40 8728 72 8760
rect 112 8728 144 8760
rect 184 8728 216 8760
rect 256 8728 288 8760
rect 328 8728 360 8760
rect 400 8728 432 8760
rect 472 8728 504 8760
rect 544 8728 576 8760
rect 616 8728 648 8760
rect 688 8728 720 8760
rect 760 8728 792 8760
rect 832 8728 864 8760
rect 904 8728 936 8760
rect 976 8728 1008 8760
rect 1048 8728 1080 8760
rect 1120 8728 1152 8760
rect 1192 8728 1224 8760
rect 1264 8728 1296 8760
rect 1336 8728 1368 8760
rect 1408 8728 1440 8760
rect 1480 8728 1512 8760
rect 1552 8728 1584 8760
rect 1624 8728 1656 8760
rect 1696 8728 1728 8760
rect 1768 8728 1800 8760
rect 1840 8728 1872 8760
rect 1912 8728 1944 8760
rect 1984 8728 2016 8760
rect 2056 8728 2088 8760
rect 2128 8728 2160 8760
rect 2200 8728 2232 8760
rect 2272 8728 2304 8760
rect 2344 8728 2376 8760
rect 2416 8728 2448 8760
rect 2488 8728 2520 8760
rect 2560 8728 2592 8760
rect 2632 8728 2664 8760
rect 2704 8728 2736 8760
rect 2776 8728 2808 8760
rect 2848 8728 2880 8760
rect 2920 8728 2952 8760
rect 2992 8728 3024 8760
rect 3064 8728 3096 8760
rect 3136 8728 3168 8760
rect 3208 8728 3240 8760
rect 3280 8728 3312 8760
rect 3352 8728 3384 8760
rect 3424 8728 3456 8760
rect 3496 8728 3528 8760
rect 3568 8728 3600 8760
rect 3640 8728 3672 8760
rect 3712 8728 3744 8760
rect 3784 8728 3816 8760
rect 3856 8728 3888 8760
rect 3928 8728 3960 8760
rect 40 8656 72 8688
rect 112 8656 144 8688
rect 184 8656 216 8688
rect 256 8656 288 8688
rect 328 8656 360 8688
rect 400 8656 432 8688
rect 472 8656 504 8688
rect 544 8656 576 8688
rect 616 8656 648 8688
rect 688 8656 720 8688
rect 760 8656 792 8688
rect 832 8656 864 8688
rect 904 8656 936 8688
rect 976 8656 1008 8688
rect 1048 8656 1080 8688
rect 1120 8656 1152 8688
rect 1192 8656 1224 8688
rect 1264 8656 1296 8688
rect 1336 8656 1368 8688
rect 1408 8656 1440 8688
rect 1480 8656 1512 8688
rect 1552 8656 1584 8688
rect 1624 8656 1656 8688
rect 1696 8656 1728 8688
rect 1768 8656 1800 8688
rect 1840 8656 1872 8688
rect 1912 8656 1944 8688
rect 1984 8656 2016 8688
rect 2056 8656 2088 8688
rect 2128 8656 2160 8688
rect 2200 8656 2232 8688
rect 2272 8656 2304 8688
rect 2344 8656 2376 8688
rect 2416 8656 2448 8688
rect 2488 8656 2520 8688
rect 2560 8656 2592 8688
rect 2632 8656 2664 8688
rect 2704 8656 2736 8688
rect 2776 8656 2808 8688
rect 2848 8656 2880 8688
rect 2920 8656 2952 8688
rect 2992 8656 3024 8688
rect 3064 8656 3096 8688
rect 3136 8656 3168 8688
rect 3208 8656 3240 8688
rect 3280 8656 3312 8688
rect 3352 8656 3384 8688
rect 3424 8656 3456 8688
rect 3496 8656 3528 8688
rect 3568 8656 3600 8688
rect 3640 8656 3672 8688
rect 3712 8656 3744 8688
rect 3784 8656 3816 8688
rect 3856 8656 3888 8688
rect 3928 8656 3960 8688
rect 40 8584 72 8616
rect 112 8584 144 8616
rect 184 8584 216 8616
rect 256 8584 288 8616
rect 328 8584 360 8616
rect 400 8584 432 8616
rect 472 8584 504 8616
rect 544 8584 576 8616
rect 616 8584 648 8616
rect 688 8584 720 8616
rect 760 8584 792 8616
rect 832 8584 864 8616
rect 904 8584 936 8616
rect 976 8584 1008 8616
rect 1048 8584 1080 8616
rect 1120 8584 1152 8616
rect 1192 8584 1224 8616
rect 1264 8584 1296 8616
rect 1336 8584 1368 8616
rect 1408 8584 1440 8616
rect 1480 8584 1512 8616
rect 1552 8584 1584 8616
rect 1624 8584 1656 8616
rect 1696 8584 1728 8616
rect 1768 8584 1800 8616
rect 1840 8584 1872 8616
rect 1912 8584 1944 8616
rect 1984 8584 2016 8616
rect 2056 8584 2088 8616
rect 2128 8584 2160 8616
rect 2200 8584 2232 8616
rect 2272 8584 2304 8616
rect 2344 8584 2376 8616
rect 2416 8584 2448 8616
rect 2488 8584 2520 8616
rect 2560 8584 2592 8616
rect 2632 8584 2664 8616
rect 2704 8584 2736 8616
rect 2776 8584 2808 8616
rect 2848 8584 2880 8616
rect 2920 8584 2952 8616
rect 2992 8584 3024 8616
rect 3064 8584 3096 8616
rect 3136 8584 3168 8616
rect 3208 8584 3240 8616
rect 3280 8584 3312 8616
rect 3352 8584 3384 8616
rect 3424 8584 3456 8616
rect 3496 8584 3528 8616
rect 3568 8584 3600 8616
rect 3640 8584 3672 8616
rect 3712 8584 3744 8616
rect 3784 8584 3816 8616
rect 3856 8584 3888 8616
rect 3928 8584 3960 8616
rect 40 8512 72 8544
rect 112 8512 144 8544
rect 184 8512 216 8544
rect 256 8512 288 8544
rect 328 8512 360 8544
rect 400 8512 432 8544
rect 472 8512 504 8544
rect 544 8512 576 8544
rect 616 8512 648 8544
rect 688 8512 720 8544
rect 760 8512 792 8544
rect 832 8512 864 8544
rect 904 8512 936 8544
rect 976 8512 1008 8544
rect 1048 8512 1080 8544
rect 1120 8512 1152 8544
rect 1192 8512 1224 8544
rect 1264 8512 1296 8544
rect 1336 8512 1368 8544
rect 1408 8512 1440 8544
rect 1480 8512 1512 8544
rect 1552 8512 1584 8544
rect 1624 8512 1656 8544
rect 1696 8512 1728 8544
rect 1768 8512 1800 8544
rect 1840 8512 1872 8544
rect 1912 8512 1944 8544
rect 1984 8512 2016 8544
rect 2056 8512 2088 8544
rect 2128 8512 2160 8544
rect 2200 8512 2232 8544
rect 2272 8512 2304 8544
rect 2344 8512 2376 8544
rect 2416 8512 2448 8544
rect 2488 8512 2520 8544
rect 2560 8512 2592 8544
rect 2632 8512 2664 8544
rect 2704 8512 2736 8544
rect 2776 8512 2808 8544
rect 2848 8512 2880 8544
rect 2920 8512 2952 8544
rect 2992 8512 3024 8544
rect 3064 8512 3096 8544
rect 3136 8512 3168 8544
rect 3208 8512 3240 8544
rect 3280 8512 3312 8544
rect 3352 8512 3384 8544
rect 3424 8512 3456 8544
rect 3496 8512 3528 8544
rect 3568 8512 3600 8544
rect 3640 8512 3672 8544
rect 3712 8512 3744 8544
rect 3784 8512 3816 8544
rect 3856 8512 3888 8544
rect 3928 8512 3960 8544
rect 40 8440 72 8472
rect 112 8440 144 8472
rect 184 8440 216 8472
rect 256 8440 288 8472
rect 328 8440 360 8472
rect 400 8440 432 8472
rect 472 8440 504 8472
rect 544 8440 576 8472
rect 616 8440 648 8472
rect 688 8440 720 8472
rect 760 8440 792 8472
rect 832 8440 864 8472
rect 904 8440 936 8472
rect 976 8440 1008 8472
rect 1048 8440 1080 8472
rect 1120 8440 1152 8472
rect 1192 8440 1224 8472
rect 1264 8440 1296 8472
rect 1336 8440 1368 8472
rect 1408 8440 1440 8472
rect 1480 8440 1512 8472
rect 1552 8440 1584 8472
rect 1624 8440 1656 8472
rect 1696 8440 1728 8472
rect 1768 8440 1800 8472
rect 1840 8440 1872 8472
rect 1912 8440 1944 8472
rect 1984 8440 2016 8472
rect 2056 8440 2088 8472
rect 2128 8440 2160 8472
rect 2200 8440 2232 8472
rect 2272 8440 2304 8472
rect 2344 8440 2376 8472
rect 2416 8440 2448 8472
rect 2488 8440 2520 8472
rect 2560 8440 2592 8472
rect 2632 8440 2664 8472
rect 2704 8440 2736 8472
rect 2776 8440 2808 8472
rect 2848 8440 2880 8472
rect 2920 8440 2952 8472
rect 2992 8440 3024 8472
rect 3064 8440 3096 8472
rect 3136 8440 3168 8472
rect 3208 8440 3240 8472
rect 3280 8440 3312 8472
rect 3352 8440 3384 8472
rect 3424 8440 3456 8472
rect 3496 8440 3528 8472
rect 3568 8440 3600 8472
rect 3640 8440 3672 8472
rect 3712 8440 3744 8472
rect 3784 8440 3816 8472
rect 3856 8440 3888 8472
rect 3928 8440 3960 8472
rect 40 8368 72 8400
rect 112 8368 144 8400
rect 184 8368 216 8400
rect 256 8368 288 8400
rect 328 8368 360 8400
rect 400 8368 432 8400
rect 472 8368 504 8400
rect 544 8368 576 8400
rect 616 8368 648 8400
rect 688 8368 720 8400
rect 760 8368 792 8400
rect 832 8368 864 8400
rect 904 8368 936 8400
rect 976 8368 1008 8400
rect 1048 8368 1080 8400
rect 1120 8368 1152 8400
rect 1192 8368 1224 8400
rect 1264 8368 1296 8400
rect 1336 8368 1368 8400
rect 1408 8368 1440 8400
rect 1480 8368 1512 8400
rect 1552 8368 1584 8400
rect 1624 8368 1656 8400
rect 1696 8368 1728 8400
rect 1768 8368 1800 8400
rect 1840 8368 1872 8400
rect 1912 8368 1944 8400
rect 1984 8368 2016 8400
rect 2056 8368 2088 8400
rect 2128 8368 2160 8400
rect 2200 8368 2232 8400
rect 2272 8368 2304 8400
rect 2344 8368 2376 8400
rect 2416 8368 2448 8400
rect 2488 8368 2520 8400
rect 2560 8368 2592 8400
rect 2632 8368 2664 8400
rect 2704 8368 2736 8400
rect 2776 8368 2808 8400
rect 2848 8368 2880 8400
rect 2920 8368 2952 8400
rect 2992 8368 3024 8400
rect 3064 8368 3096 8400
rect 3136 8368 3168 8400
rect 3208 8368 3240 8400
rect 3280 8368 3312 8400
rect 3352 8368 3384 8400
rect 3424 8368 3456 8400
rect 3496 8368 3528 8400
rect 3568 8368 3600 8400
rect 3640 8368 3672 8400
rect 3712 8368 3744 8400
rect 3784 8368 3816 8400
rect 3856 8368 3888 8400
rect 3928 8368 3960 8400
rect 40 8296 72 8328
rect 112 8296 144 8328
rect 184 8296 216 8328
rect 256 8296 288 8328
rect 328 8296 360 8328
rect 400 8296 432 8328
rect 472 8296 504 8328
rect 544 8296 576 8328
rect 616 8296 648 8328
rect 688 8296 720 8328
rect 760 8296 792 8328
rect 832 8296 864 8328
rect 904 8296 936 8328
rect 976 8296 1008 8328
rect 1048 8296 1080 8328
rect 1120 8296 1152 8328
rect 1192 8296 1224 8328
rect 1264 8296 1296 8328
rect 1336 8296 1368 8328
rect 1408 8296 1440 8328
rect 1480 8296 1512 8328
rect 1552 8296 1584 8328
rect 1624 8296 1656 8328
rect 1696 8296 1728 8328
rect 1768 8296 1800 8328
rect 1840 8296 1872 8328
rect 1912 8296 1944 8328
rect 1984 8296 2016 8328
rect 2056 8296 2088 8328
rect 2128 8296 2160 8328
rect 2200 8296 2232 8328
rect 2272 8296 2304 8328
rect 2344 8296 2376 8328
rect 2416 8296 2448 8328
rect 2488 8296 2520 8328
rect 2560 8296 2592 8328
rect 2632 8296 2664 8328
rect 2704 8296 2736 8328
rect 2776 8296 2808 8328
rect 2848 8296 2880 8328
rect 2920 8296 2952 8328
rect 2992 8296 3024 8328
rect 3064 8296 3096 8328
rect 3136 8296 3168 8328
rect 3208 8296 3240 8328
rect 3280 8296 3312 8328
rect 3352 8296 3384 8328
rect 3424 8296 3456 8328
rect 3496 8296 3528 8328
rect 3568 8296 3600 8328
rect 3640 8296 3672 8328
rect 3712 8296 3744 8328
rect 3784 8296 3816 8328
rect 3856 8296 3888 8328
rect 3928 8296 3960 8328
rect 40 8224 72 8256
rect 112 8224 144 8256
rect 184 8224 216 8256
rect 256 8224 288 8256
rect 328 8224 360 8256
rect 400 8224 432 8256
rect 472 8224 504 8256
rect 544 8224 576 8256
rect 616 8224 648 8256
rect 688 8224 720 8256
rect 760 8224 792 8256
rect 832 8224 864 8256
rect 904 8224 936 8256
rect 976 8224 1008 8256
rect 1048 8224 1080 8256
rect 1120 8224 1152 8256
rect 1192 8224 1224 8256
rect 1264 8224 1296 8256
rect 1336 8224 1368 8256
rect 1408 8224 1440 8256
rect 1480 8224 1512 8256
rect 1552 8224 1584 8256
rect 1624 8224 1656 8256
rect 1696 8224 1728 8256
rect 1768 8224 1800 8256
rect 1840 8224 1872 8256
rect 1912 8224 1944 8256
rect 1984 8224 2016 8256
rect 2056 8224 2088 8256
rect 2128 8224 2160 8256
rect 2200 8224 2232 8256
rect 2272 8224 2304 8256
rect 2344 8224 2376 8256
rect 2416 8224 2448 8256
rect 2488 8224 2520 8256
rect 2560 8224 2592 8256
rect 2632 8224 2664 8256
rect 2704 8224 2736 8256
rect 2776 8224 2808 8256
rect 2848 8224 2880 8256
rect 2920 8224 2952 8256
rect 2992 8224 3024 8256
rect 3064 8224 3096 8256
rect 3136 8224 3168 8256
rect 3208 8224 3240 8256
rect 3280 8224 3312 8256
rect 3352 8224 3384 8256
rect 3424 8224 3456 8256
rect 3496 8224 3528 8256
rect 3568 8224 3600 8256
rect 3640 8224 3672 8256
rect 3712 8224 3744 8256
rect 3784 8224 3816 8256
rect 3856 8224 3888 8256
rect 3928 8224 3960 8256
rect 40 8152 72 8184
rect 112 8152 144 8184
rect 184 8152 216 8184
rect 256 8152 288 8184
rect 328 8152 360 8184
rect 400 8152 432 8184
rect 472 8152 504 8184
rect 544 8152 576 8184
rect 616 8152 648 8184
rect 688 8152 720 8184
rect 760 8152 792 8184
rect 832 8152 864 8184
rect 904 8152 936 8184
rect 976 8152 1008 8184
rect 1048 8152 1080 8184
rect 1120 8152 1152 8184
rect 1192 8152 1224 8184
rect 1264 8152 1296 8184
rect 1336 8152 1368 8184
rect 1408 8152 1440 8184
rect 1480 8152 1512 8184
rect 1552 8152 1584 8184
rect 1624 8152 1656 8184
rect 1696 8152 1728 8184
rect 1768 8152 1800 8184
rect 1840 8152 1872 8184
rect 1912 8152 1944 8184
rect 1984 8152 2016 8184
rect 2056 8152 2088 8184
rect 2128 8152 2160 8184
rect 2200 8152 2232 8184
rect 2272 8152 2304 8184
rect 2344 8152 2376 8184
rect 2416 8152 2448 8184
rect 2488 8152 2520 8184
rect 2560 8152 2592 8184
rect 2632 8152 2664 8184
rect 2704 8152 2736 8184
rect 2776 8152 2808 8184
rect 2848 8152 2880 8184
rect 2920 8152 2952 8184
rect 2992 8152 3024 8184
rect 3064 8152 3096 8184
rect 3136 8152 3168 8184
rect 3208 8152 3240 8184
rect 3280 8152 3312 8184
rect 3352 8152 3384 8184
rect 3424 8152 3456 8184
rect 3496 8152 3528 8184
rect 3568 8152 3600 8184
rect 3640 8152 3672 8184
rect 3712 8152 3744 8184
rect 3784 8152 3816 8184
rect 3856 8152 3888 8184
rect 3928 8152 3960 8184
rect 40 8080 72 8112
rect 112 8080 144 8112
rect 184 8080 216 8112
rect 256 8080 288 8112
rect 328 8080 360 8112
rect 400 8080 432 8112
rect 472 8080 504 8112
rect 544 8080 576 8112
rect 616 8080 648 8112
rect 688 8080 720 8112
rect 760 8080 792 8112
rect 832 8080 864 8112
rect 904 8080 936 8112
rect 976 8080 1008 8112
rect 1048 8080 1080 8112
rect 1120 8080 1152 8112
rect 1192 8080 1224 8112
rect 1264 8080 1296 8112
rect 1336 8080 1368 8112
rect 1408 8080 1440 8112
rect 1480 8080 1512 8112
rect 1552 8080 1584 8112
rect 1624 8080 1656 8112
rect 1696 8080 1728 8112
rect 1768 8080 1800 8112
rect 1840 8080 1872 8112
rect 1912 8080 1944 8112
rect 1984 8080 2016 8112
rect 2056 8080 2088 8112
rect 2128 8080 2160 8112
rect 2200 8080 2232 8112
rect 2272 8080 2304 8112
rect 2344 8080 2376 8112
rect 2416 8080 2448 8112
rect 2488 8080 2520 8112
rect 2560 8080 2592 8112
rect 2632 8080 2664 8112
rect 2704 8080 2736 8112
rect 2776 8080 2808 8112
rect 2848 8080 2880 8112
rect 2920 8080 2952 8112
rect 2992 8080 3024 8112
rect 3064 8080 3096 8112
rect 3136 8080 3168 8112
rect 3208 8080 3240 8112
rect 3280 8080 3312 8112
rect 3352 8080 3384 8112
rect 3424 8080 3456 8112
rect 3496 8080 3528 8112
rect 3568 8080 3600 8112
rect 3640 8080 3672 8112
rect 3712 8080 3744 8112
rect 3784 8080 3816 8112
rect 3856 8080 3888 8112
rect 3928 8080 3960 8112
rect 40 8008 72 8040
rect 112 8008 144 8040
rect 184 8008 216 8040
rect 256 8008 288 8040
rect 328 8008 360 8040
rect 400 8008 432 8040
rect 472 8008 504 8040
rect 544 8008 576 8040
rect 616 8008 648 8040
rect 688 8008 720 8040
rect 760 8008 792 8040
rect 832 8008 864 8040
rect 904 8008 936 8040
rect 976 8008 1008 8040
rect 1048 8008 1080 8040
rect 1120 8008 1152 8040
rect 1192 8008 1224 8040
rect 1264 8008 1296 8040
rect 1336 8008 1368 8040
rect 1408 8008 1440 8040
rect 1480 8008 1512 8040
rect 1552 8008 1584 8040
rect 1624 8008 1656 8040
rect 1696 8008 1728 8040
rect 1768 8008 1800 8040
rect 1840 8008 1872 8040
rect 1912 8008 1944 8040
rect 1984 8008 2016 8040
rect 2056 8008 2088 8040
rect 2128 8008 2160 8040
rect 2200 8008 2232 8040
rect 2272 8008 2304 8040
rect 2344 8008 2376 8040
rect 2416 8008 2448 8040
rect 2488 8008 2520 8040
rect 2560 8008 2592 8040
rect 2632 8008 2664 8040
rect 2704 8008 2736 8040
rect 2776 8008 2808 8040
rect 2848 8008 2880 8040
rect 2920 8008 2952 8040
rect 2992 8008 3024 8040
rect 3064 8008 3096 8040
rect 3136 8008 3168 8040
rect 3208 8008 3240 8040
rect 3280 8008 3312 8040
rect 3352 8008 3384 8040
rect 3424 8008 3456 8040
rect 3496 8008 3528 8040
rect 3568 8008 3600 8040
rect 3640 8008 3672 8040
rect 3712 8008 3744 8040
rect 3784 8008 3816 8040
rect 3856 8008 3888 8040
rect 3928 8008 3960 8040
rect 40 7936 72 7968
rect 112 7936 144 7968
rect 184 7936 216 7968
rect 256 7936 288 7968
rect 328 7936 360 7968
rect 400 7936 432 7968
rect 472 7936 504 7968
rect 544 7936 576 7968
rect 616 7936 648 7968
rect 688 7936 720 7968
rect 760 7936 792 7968
rect 832 7936 864 7968
rect 904 7936 936 7968
rect 976 7936 1008 7968
rect 1048 7936 1080 7968
rect 1120 7936 1152 7968
rect 1192 7936 1224 7968
rect 1264 7936 1296 7968
rect 1336 7936 1368 7968
rect 1408 7936 1440 7968
rect 1480 7936 1512 7968
rect 1552 7936 1584 7968
rect 1624 7936 1656 7968
rect 1696 7936 1728 7968
rect 1768 7936 1800 7968
rect 1840 7936 1872 7968
rect 1912 7936 1944 7968
rect 1984 7936 2016 7968
rect 2056 7936 2088 7968
rect 2128 7936 2160 7968
rect 2200 7936 2232 7968
rect 2272 7936 2304 7968
rect 2344 7936 2376 7968
rect 2416 7936 2448 7968
rect 2488 7936 2520 7968
rect 2560 7936 2592 7968
rect 2632 7936 2664 7968
rect 2704 7936 2736 7968
rect 2776 7936 2808 7968
rect 2848 7936 2880 7968
rect 2920 7936 2952 7968
rect 2992 7936 3024 7968
rect 3064 7936 3096 7968
rect 3136 7936 3168 7968
rect 3208 7936 3240 7968
rect 3280 7936 3312 7968
rect 3352 7936 3384 7968
rect 3424 7936 3456 7968
rect 3496 7936 3528 7968
rect 3568 7936 3600 7968
rect 3640 7936 3672 7968
rect 3712 7936 3744 7968
rect 3784 7936 3816 7968
rect 3856 7936 3888 7968
rect 3928 7936 3960 7968
rect 40 7864 72 7896
rect 112 7864 144 7896
rect 184 7864 216 7896
rect 256 7864 288 7896
rect 328 7864 360 7896
rect 400 7864 432 7896
rect 472 7864 504 7896
rect 544 7864 576 7896
rect 616 7864 648 7896
rect 688 7864 720 7896
rect 760 7864 792 7896
rect 832 7864 864 7896
rect 904 7864 936 7896
rect 976 7864 1008 7896
rect 1048 7864 1080 7896
rect 1120 7864 1152 7896
rect 1192 7864 1224 7896
rect 1264 7864 1296 7896
rect 1336 7864 1368 7896
rect 1408 7864 1440 7896
rect 1480 7864 1512 7896
rect 1552 7864 1584 7896
rect 1624 7864 1656 7896
rect 1696 7864 1728 7896
rect 1768 7864 1800 7896
rect 1840 7864 1872 7896
rect 1912 7864 1944 7896
rect 1984 7864 2016 7896
rect 2056 7864 2088 7896
rect 2128 7864 2160 7896
rect 2200 7864 2232 7896
rect 2272 7864 2304 7896
rect 2344 7864 2376 7896
rect 2416 7864 2448 7896
rect 2488 7864 2520 7896
rect 2560 7864 2592 7896
rect 2632 7864 2664 7896
rect 2704 7864 2736 7896
rect 2776 7864 2808 7896
rect 2848 7864 2880 7896
rect 2920 7864 2952 7896
rect 2992 7864 3024 7896
rect 3064 7864 3096 7896
rect 3136 7864 3168 7896
rect 3208 7864 3240 7896
rect 3280 7864 3312 7896
rect 3352 7864 3384 7896
rect 3424 7864 3456 7896
rect 3496 7864 3528 7896
rect 3568 7864 3600 7896
rect 3640 7864 3672 7896
rect 3712 7864 3744 7896
rect 3784 7864 3816 7896
rect 3856 7864 3888 7896
rect 3928 7864 3960 7896
rect 40 7792 72 7824
rect 112 7792 144 7824
rect 184 7792 216 7824
rect 256 7792 288 7824
rect 328 7792 360 7824
rect 400 7792 432 7824
rect 472 7792 504 7824
rect 544 7792 576 7824
rect 616 7792 648 7824
rect 688 7792 720 7824
rect 760 7792 792 7824
rect 832 7792 864 7824
rect 904 7792 936 7824
rect 976 7792 1008 7824
rect 1048 7792 1080 7824
rect 1120 7792 1152 7824
rect 1192 7792 1224 7824
rect 1264 7792 1296 7824
rect 1336 7792 1368 7824
rect 1408 7792 1440 7824
rect 1480 7792 1512 7824
rect 1552 7792 1584 7824
rect 1624 7792 1656 7824
rect 1696 7792 1728 7824
rect 1768 7792 1800 7824
rect 1840 7792 1872 7824
rect 1912 7792 1944 7824
rect 1984 7792 2016 7824
rect 2056 7792 2088 7824
rect 2128 7792 2160 7824
rect 2200 7792 2232 7824
rect 2272 7792 2304 7824
rect 2344 7792 2376 7824
rect 2416 7792 2448 7824
rect 2488 7792 2520 7824
rect 2560 7792 2592 7824
rect 2632 7792 2664 7824
rect 2704 7792 2736 7824
rect 2776 7792 2808 7824
rect 2848 7792 2880 7824
rect 2920 7792 2952 7824
rect 2992 7792 3024 7824
rect 3064 7792 3096 7824
rect 3136 7792 3168 7824
rect 3208 7792 3240 7824
rect 3280 7792 3312 7824
rect 3352 7792 3384 7824
rect 3424 7792 3456 7824
rect 3496 7792 3528 7824
rect 3568 7792 3600 7824
rect 3640 7792 3672 7824
rect 3712 7792 3744 7824
rect 3784 7792 3816 7824
rect 3856 7792 3888 7824
rect 3928 7792 3960 7824
rect 40 7720 72 7752
rect 112 7720 144 7752
rect 184 7720 216 7752
rect 256 7720 288 7752
rect 328 7720 360 7752
rect 400 7720 432 7752
rect 472 7720 504 7752
rect 544 7720 576 7752
rect 616 7720 648 7752
rect 688 7720 720 7752
rect 760 7720 792 7752
rect 832 7720 864 7752
rect 904 7720 936 7752
rect 976 7720 1008 7752
rect 1048 7720 1080 7752
rect 1120 7720 1152 7752
rect 1192 7720 1224 7752
rect 1264 7720 1296 7752
rect 1336 7720 1368 7752
rect 1408 7720 1440 7752
rect 1480 7720 1512 7752
rect 1552 7720 1584 7752
rect 1624 7720 1656 7752
rect 1696 7720 1728 7752
rect 1768 7720 1800 7752
rect 1840 7720 1872 7752
rect 1912 7720 1944 7752
rect 1984 7720 2016 7752
rect 2056 7720 2088 7752
rect 2128 7720 2160 7752
rect 2200 7720 2232 7752
rect 2272 7720 2304 7752
rect 2344 7720 2376 7752
rect 2416 7720 2448 7752
rect 2488 7720 2520 7752
rect 2560 7720 2592 7752
rect 2632 7720 2664 7752
rect 2704 7720 2736 7752
rect 2776 7720 2808 7752
rect 2848 7720 2880 7752
rect 2920 7720 2952 7752
rect 2992 7720 3024 7752
rect 3064 7720 3096 7752
rect 3136 7720 3168 7752
rect 3208 7720 3240 7752
rect 3280 7720 3312 7752
rect 3352 7720 3384 7752
rect 3424 7720 3456 7752
rect 3496 7720 3528 7752
rect 3568 7720 3600 7752
rect 3640 7720 3672 7752
rect 3712 7720 3744 7752
rect 3784 7720 3816 7752
rect 3856 7720 3888 7752
rect 3928 7720 3960 7752
rect 40 7648 72 7680
rect 112 7648 144 7680
rect 184 7648 216 7680
rect 256 7648 288 7680
rect 328 7648 360 7680
rect 400 7648 432 7680
rect 472 7648 504 7680
rect 544 7648 576 7680
rect 616 7648 648 7680
rect 688 7648 720 7680
rect 760 7648 792 7680
rect 832 7648 864 7680
rect 904 7648 936 7680
rect 976 7648 1008 7680
rect 1048 7648 1080 7680
rect 1120 7648 1152 7680
rect 1192 7648 1224 7680
rect 1264 7648 1296 7680
rect 1336 7648 1368 7680
rect 1408 7648 1440 7680
rect 1480 7648 1512 7680
rect 1552 7648 1584 7680
rect 1624 7648 1656 7680
rect 1696 7648 1728 7680
rect 1768 7648 1800 7680
rect 1840 7648 1872 7680
rect 1912 7648 1944 7680
rect 1984 7648 2016 7680
rect 2056 7648 2088 7680
rect 2128 7648 2160 7680
rect 2200 7648 2232 7680
rect 2272 7648 2304 7680
rect 2344 7648 2376 7680
rect 2416 7648 2448 7680
rect 2488 7648 2520 7680
rect 2560 7648 2592 7680
rect 2632 7648 2664 7680
rect 2704 7648 2736 7680
rect 2776 7648 2808 7680
rect 2848 7648 2880 7680
rect 2920 7648 2952 7680
rect 2992 7648 3024 7680
rect 3064 7648 3096 7680
rect 3136 7648 3168 7680
rect 3208 7648 3240 7680
rect 3280 7648 3312 7680
rect 3352 7648 3384 7680
rect 3424 7648 3456 7680
rect 3496 7648 3528 7680
rect 3568 7648 3600 7680
rect 3640 7648 3672 7680
rect 3712 7648 3744 7680
rect 3784 7648 3816 7680
rect 3856 7648 3888 7680
rect 3928 7648 3960 7680
rect 40 7576 72 7608
rect 112 7576 144 7608
rect 184 7576 216 7608
rect 256 7576 288 7608
rect 328 7576 360 7608
rect 400 7576 432 7608
rect 472 7576 504 7608
rect 544 7576 576 7608
rect 616 7576 648 7608
rect 688 7576 720 7608
rect 760 7576 792 7608
rect 832 7576 864 7608
rect 904 7576 936 7608
rect 976 7576 1008 7608
rect 1048 7576 1080 7608
rect 1120 7576 1152 7608
rect 1192 7576 1224 7608
rect 1264 7576 1296 7608
rect 1336 7576 1368 7608
rect 1408 7576 1440 7608
rect 1480 7576 1512 7608
rect 1552 7576 1584 7608
rect 1624 7576 1656 7608
rect 1696 7576 1728 7608
rect 1768 7576 1800 7608
rect 1840 7576 1872 7608
rect 1912 7576 1944 7608
rect 1984 7576 2016 7608
rect 2056 7576 2088 7608
rect 2128 7576 2160 7608
rect 2200 7576 2232 7608
rect 2272 7576 2304 7608
rect 2344 7576 2376 7608
rect 2416 7576 2448 7608
rect 2488 7576 2520 7608
rect 2560 7576 2592 7608
rect 2632 7576 2664 7608
rect 2704 7576 2736 7608
rect 2776 7576 2808 7608
rect 2848 7576 2880 7608
rect 2920 7576 2952 7608
rect 2992 7576 3024 7608
rect 3064 7576 3096 7608
rect 3136 7576 3168 7608
rect 3208 7576 3240 7608
rect 3280 7576 3312 7608
rect 3352 7576 3384 7608
rect 3424 7576 3456 7608
rect 3496 7576 3528 7608
rect 3568 7576 3600 7608
rect 3640 7576 3672 7608
rect 3712 7576 3744 7608
rect 3784 7576 3816 7608
rect 3856 7576 3888 7608
rect 3928 7576 3960 7608
rect 40 7504 72 7536
rect 112 7504 144 7536
rect 184 7504 216 7536
rect 256 7504 288 7536
rect 328 7504 360 7536
rect 400 7504 432 7536
rect 472 7504 504 7536
rect 544 7504 576 7536
rect 616 7504 648 7536
rect 688 7504 720 7536
rect 760 7504 792 7536
rect 832 7504 864 7536
rect 904 7504 936 7536
rect 976 7504 1008 7536
rect 1048 7504 1080 7536
rect 1120 7504 1152 7536
rect 1192 7504 1224 7536
rect 1264 7504 1296 7536
rect 1336 7504 1368 7536
rect 1408 7504 1440 7536
rect 1480 7504 1512 7536
rect 1552 7504 1584 7536
rect 1624 7504 1656 7536
rect 1696 7504 1728 7536
rect 1768 7504 1800 7536
rect 1840 7504 1872 7536
rect 1912 7504 1944 7536
rect 1984 7504 2016 7536
rect 2056 7504 2088 7536
rect 2128 7504 2160 7536
rect 2200 7504 2232 7536
rect 2272 7504 2304 7536
rect 2344 7504 2376 7536
rect 2416 7504 2448 7536
rect 2488 7504 2520 7536
rect 2560 7504 2592 7536
rect 2632 7504 2664 7536
rect 2704 7504 2736 7536
rect 2776 7504 2808 7536
rect 2848 7504 2880 7536
rect 2920 7504 2952 7536
rect 2992 7504 3024 7536
rect 3064 7504 3096 7536
rect 3136 7504 3168 7536
rect 3208 7504 3240 7536
rect 3280 7504 3312 7536
rect 3352 7504 3384 7536
rect 3424 7504 3456 7536
rect 3496 7504 3528 7536
rect 3568 7504 3600 7536
rect 3640 7504 3672 7536
rect 3712 7504 3744 7536
rect 3784 7504 3816 7536
rect 3856 7504 3888 7536
rect 3928 7504 3960 7536
rect 40 7432 72 7464
rect 112 7432 144 7464
rect 184 7432 216 7464
rect 256 7432 288 7464
rect 328 7432 360 7464
rect 400 7432 432 7464
rect 472 7432 504 7464
rect 544 7432 576 7464
rect 616 7432 648 7464
rect 688 7432 720 7464
rect 760 7432 792 7464
rect 832 7432 864 7464
rect 904 7432 936 7464
rect 976 7432 1008 7464
rect 1048 7432 1080 7464
rect 1120 7432 1152 7464
rect 1192 7432 1224 7464
rect 1264 7432 1296 7464
rect 1336 7432 1368 7464
rect 1408 7432 1440 7464
rect 1480 7432 1512 7464
rect 1552 7432 1584 7464
rect 1624 7432 1656 7464
rect 1696 7432 1728 7464
rect 1768 7432 1800 7464
rect 1840 7432 1872 7464
rect 1912 7432 1944 7464
rect 1984 7432 2016 7464
rect 2056 7432 2088 7464
rect 2128 7432 2160 7464
rect 2200 7432 2232 7464
rect 2272 7432 2304 7464
rect 2344 7432 2376 7464
rect 2416 7432 2448 7464
rect 2488 7432 2520 7464
rect 2560 7432 2592 7464
rect 2632 7432 2664 7464
rect 2704 7432 2736 7464
rect 2776 7432 2808 7464
rect 2848 7432 2880 7464
rect 2920 7432 2952 7464
rect 2992 7432 3024 7464
rect 3064 7432 3096 7464
rect 3136 7432 3168 7464
rect 3208 7432 3240 7464
rect 3280 7432 3312 7464
rect 3352 7432 3384 7464
rect 3424 7432 3456 7464
rect 3496 7432 3528 7464
rect 3568 7432 3600 7464
rect 3640 7432 3672 7464
rect 3712 7432 3744 7464
rect 3784 7432 3816 7464
rect 3856 7432 3888 7464
rect 3928 7432 3960 7464
rect 40 7360 72 7392
rect 112 7360 144 7392
rect 184 7360 216 7392
rect 256 7360 288 7392
rect 328 7360 360 7392
rect 400 7360 432 7392
rect 472 7360 504 7392
rect 544 7360 576 7392
rect 616 7360 648 7392
rect 688 7360 720 7392
rect 760 7360 792 7392
rect 832 7360 864 7392
rect 904 7360 936 7392
rect 976 7360 1008 7392
rect 1048 7360 1080 7392
rect 1120 7360 1152 7392
rect 1192 7360 1224 7392
rect 1264 7360 1296 7392
rect 1336 7360 1368 7392
rect 1408 7360 1440 7392
rect 1480 7360 1512 7392
rect 1552 7360 1584 7392
rect 1624 7360 1656 7392
rect 1696 7360 1728 7392
rect 1768 7360 1800 7392
rect 1840 7360 1872 7392
rect 1912 7360 1944 7392
rect 1984 7360 2016 7392
rect 2056 7360 2088 7392
rect 2128 7360 2160 7392
rect 2200 7360 2232 7392
rect 2272 7360 2304 7392
rect 2344 7360 2376 7392
rect 2416 7360 2448 7392
rect 2488 7360 2520 7392
rect 2560 7360 2592 7392
rect 2632 7360 2664 7392
rect 2704 7360 2736 7392
rect 2776 7360 2808 7392
rect 2848 7360 2880 7392
rect 2920 7360 2952 7392
rect 2992 7360 3024 7392
rect 3064 7360 3096 7392
rect 3136 7360 3168 7392
rect 3208 7360 3240 7392
rect 3280 7360 3312 7392
rect 3352 7360 3384 7392
rect 3424 7360 3456 7392
rect 3496 7360 3528 7392
rect 3568 7360 3600 7392
rect 3640 7360 3672 7392
rect 3712 7360 3744 7392
rect 3784 7360 3816 7392
rect 3856 7360 3888 7392
rect 3928 7360 3960 7392
rect 40 7288 72 7320
rect 112 7288 144 7320
rect 184 7288 216 7320
rect 256 7288 288 7320
rect 328 7288 360 7320
rect 400 7288 432 7320
rect 472 7288 504 7320
rect 544 7288 576 7320
rect 616 7288 648 7320
rect 688 7288 720 7320
rect 760 7288 792 7320
rect 832 7288 864 7320
rect 904 7288 936 7320
rect 976 7288 1008 7320
rect 1048 7288 1080 7320
rect 1120 7288 1152 7320
rect 1192 7288 1224 7320
rect 1264 7288 1296 7320
rect 1336 7288 1368 7320
rect 1408 7288 1440 7320
rect 1480 7288 1512 7320
rect 1552 7288 1584 7320
rect 1624 7288 1656 7320
rect 1696 7288 1728 7320
rect 1768 7288 1800 7320
rect 1840 7288 1872 7320
rect 1912 7288 1944 7320
rect 1984 7288 2016 7320
rect 2056 7288 2088 7320
rect 2128 7288 2160 7320
rect 2200 7288 2232 7320
rect 2272 7288 2304 7320
rect 2344 7288 2376 7320
rect 2416 7288 2448 7320
rect 2488 7288 2520 7320
rect 2560 7288 2592 7320
rect 2632 7288 2664 7320
rect 2704 7288 2736 7320
rect 2776 7288 2808 7320
rect 2848 7288 2880 7320
rect 2920 7288 2952 7320
rect 2992 7288 3024 7320
rect 3064 7288 3096 7320
rect 3136 7288 3168 7320
rect 3208 7288 3240 7320
rect 3280 7288 3312 7320
rect 3352 7288 3384 7320
rect 3424 7288 3456 7320
rect 3496 7288 3528 7320
rect 3568 7288 3600 7320
rect 3640 7288 3672 7320
rect 3712 7288 3744 7320
rect 3784 7288 3816 7320
rect 3856 7288 3888 7320
rect 3928 7288 3960 7320
rect 40 7216 72 7248
rect 112 7216 144 7248
rect 184 7216 216 7248
rect 256 7216 288 7248
rect 328 7216 360 7248
rect 400 7216 432 7248
rect 472 7216 504 7248
rect 544 7216 576 7248
rect 616 7216 648 7248
rect 688 7216 720 7248
rect 760 7216 792 7248
rect 832 7216 864 7248
rect 904 7216 936 7248
rect 976 7216 1008 7248
rect 1048 7216 1080 7248
rect 1120 7216 1152 7248
rect 1192 7216 1224 7248
rect 1264 7216 1296 7248
rect 1336 7216 1368 7248
rect 1408 7216 1440 7248
rect 1480 7216 1512 7248
rect 1552 7216 1584 7248
rect 1624 7216 1656 7248
rect 1696 7216 1728 7248
rect 1768 7216 1800 7248
rect 1840 7216 1872 7248
rect 1912 7216 1944 7248
rect 1984 7216 2016 7248
rect 2056 7216 2088 7248
rect 2128 7216 2160 7248
rect 2200 7216 2232 7248
rect 2272 7216 2304 7248
rect 2344 7216 2376 7248
rect 2416 7216 2448 7248
rect 2488 7216 2520 7248
rect 2560 7216 2592 7248
rect 2632 7216 2664 7248
rect 2704 7216 2736 7248
rect 2776 7216 2808 7248
rect 2848 7216 2880 7248
rect 2920 7216 2952 7248
rect 2992 7216 3024 7248
rect 3064 7216 3096 7248
rect 3136 7216 3168 7248
rect 3208 7216 3240 7248
rect 3280 7216 3312 7248
rect 3352 7216 3384 7248
rect 3424 7216 3456 7248
rect 3496 7216 3528 7248
rect 3568 7216 3600 7248
rect 3640 7216 3672 7248
rect 3712 7216 3744 7248
rect 3784 7216 3816 7248
rect 3856 7216 3888 7248
rect 3928 7216 3960 7248
rect 40 7144 72 7176
rect 112 7144 144 7176
rect 184 7144 216 7176
rect 256 7144 288 7176
rect 328 7144 360 7176
rect 400 7144 432 7176
rect 472 7144 504 7176
rect 544 7144 576 7176
rect 616 7144 648 7176
rect 688 7144 720 7176
rect 760 7144 792 7176
rect 832 7144 864 7176
rect 904 7144 936 7176
rect 976 7144 1008 7176
rect 1048 7144 1080 7176
rect 1120 7144 1152 7176
rect 1192 7144 1224 7176
rect 1264 7144 1296 7176
rect 1336 7144 1368 7176
rect 1408 7144 1440 7176
rect 1480 7144 1512 7176
rect 1552 7144 1584 7176
rect 1624 7144 1656 7176
rect 1696 7144 1728 7176
rect 1768 7144 1800 7176
rect 1840 7144 1872 7176
rect 1912 7144 1944 7176
rect 1984 7144 2016 7176
rect 2056 7144 2088 7176
rect 2128 7144 2160 7176
rect 2200 7144 2232 7176
rect 2272 7144 2304 7176
rect 2344 7144 2376 7176
rect 2416 7144 2448 7176
rect 2488 7144 2520 7176
rect 2560 7144 2592 7176
rect 2632 7144 2664 7176
rect 2704 7144 2736 7176
rect 2776 7144 2808 7176
rect 2848 7144 2880 7176
rect 2920 7144 2952 7176
rect 2992 7144 3024 7176
rect 3064 7144 3096 7176
rect 3136 7144 3168 7176
rect 3208 7144 3240 7176
rect 3280 7144 3312 7176
rect 3352 7144 3384 7176
rect 3424 7144 3456 7176
rect 3496 7144 3528 7176
rect 3568 7144 3600 7176
rect 3640 7144 3672 7176
rect 3712 7144 3744 7176
rect 3784 7144 3816 7176
rect 3856 7144 3888 7176
rect 3928 7144 3960 7176
rect 40 7072 72 7104
rect 112 7072 144 7104
rect 184 7072 216 7104
rect 256 7072 288 7104
rect 328 7072 360 7104
rect 400 7072 432 7104
rect 472 7072 504 7104
rect 544 7072 576 7104
rect 616 7072 648 7104
rect 688 7072 720 7104
rect 760 7072 792 7104
rect 832 7072 864 7104
rect 904 7072 936 7104
rect 976 7072 1008 7104
rect 1048 7072 1080 7104
rect 1120 7072 1152 7104
rect 1192 7072 1224 7104
rect 1264 7072 1296 7104
rect 1336 7072 1368 7104
rect 1408 7072 1440 7104
rect 1480 7072 1512 7104
rect 1552 7072 1584 7104
rect 1624 7072 1656 7104
rect 1696 7072 1728 7104
rect 1768 7072 1800 7104
rect 1840 7072 1872 7104
rect 1912 7072 1944 7104
rect 1984 7072 2016 7104
rect 2056 7072 2088 7104
rect 2128 7072 2160 7104
rect 2200 7072 2232 7104
rect 2272 7072 2304 7104
rect 2344 7072 2376 7104
rect 2416 7072 2448 7104
rect 2488 7072 2520 7104
rect 2560 7072 2592 7104
rect 2632 7072 2664 7104
rect 2704 7072 2736 7104
rect 2776 7072 2808 7104
rect 2848 7072 2880 7104
rect 2920 7072 2952 7104
rect 2992 7072 3024 7104
rect 3064 7072 3096 7104
rect 3136 7072 3168 7104
rect 3208 7072 3240 7104
rect 3280 7072 3312 7104
rect 3352 7072 3384 7104
rect 3424 7072 3456 7104
rect 3496 7072 3528 7104
rect 3568 7072 3600 7104
rect 3640 7072 3672 7104
rect 3712 7072 3744 7104
rect 3784 7072 3816 7104
rect 3856 7072 3888 7104
rect 3928 7072 3960 7104
rect 40 7000 72 7032
rect 112 7000 144 7032
rect 184 7000 216 7032
rect 256 7000 288 7032
rect 328 7000 360 7032
rect 400 7000 432 7032
rect 472 7000 504 7032
rect 544 7000 576 7032
rect 616 7000 648 7032
rect 688 7000 720 7032
rect 760 7000 792 7032
rect 832 7000 864 7032
rect 904 7000 936 7032
rect 976 7000 1008 7032
rect 1048 7000 1080 7032
rect 1120 7000 1152 7032
rect 1192 7000 1224 7032
rect 1264 7000 1296 7032
rect 1336 7000 1368 7032
rect 1408 7000 1440 7032
rect 1480 7000 1512 7032
rect 1552 7000 1584 7032
rect 1624 7000 1656 7032
rect 1696 7000 1728 7032
rect 1768 7000 1800 7032
rect 1840 7000 1872 7032
rect 1912 7000 1944 7032
rect 1984 7000 2016 7032
rect 2056 7000 2088 7032
rect 2128 7000 2160 7032
rect 2200 7000 2232 7032
rect 2272 7000 2304 7032
rect 2344 7000 2376 7032
rect 2416 7000 2448 7032
rect 2488 7000 2520 7032
rect 2560 7000 2592 7032
rect 2632 7000 2664 7032
rect 2704 7000 2736 7032
rect 2776 7000 2808 7032
rect 2848 7000 2880 7032
rect 2920 7000 2952 7032
rect 2992 7000 3024 7032
rect 3064 7000 3096 7032
rect 3136 7000 3168 7032
rect 3208 7000 3240 7032
rect 3280 7000 3312 7032
rect 3352 7000 3384 7032
rect 3424 7000 3456 7032
rect 3496 7000 3528 7032
rect 3568 7000 3600 7032
rect 3640 7000 3672 7032
rect 3712 7000 3744 7032
rect 3784 7000 3816 7032
rect 3856 7000 3888 7032
rect 3928 7000 3960 7032
rect 40 6928 72 6960
rect 112 6928 144 6960
rect 184 6928 216 6960
rect 256 6928 288 6960
rect 328 6928 360 6960
rect 400 6928 432 6960
rect 472 6928 504 6960
rect 544 6928 576 6960
rect 616 6928 648 6960
rect 688 6928 720 6960
rect 760 6928 792 6960
rect 832 6928 864 6960
rect 904 6928 936 6960
rect 976 6928 1008 6960
rect 1048 6928 1080 6960
rect 1120 6928 1152 6960
rect 1192 6928 1224 6960
rect 1264 6928 1296 6960
rect 1336 6928 1368 6960
rect 1408 6928 1440 6960
rect 1480 6928 1512 6960
rect 1552 6928 1584 6960
rect 1624 6928 1656 6960
rect 1696 6928 1728 6960
rect 1768 6928 1800 6960
rect 1840 6928 1872 6960
rect 1912 6928 1944 6960
rect 1984 6928 2016 6960
rect 2056 6928 2088 6960
rect 2128 6928 2160 6960
rect 2200 6928 2232 6960
rect 2272 6928 2304 6960
rect 2344 6928 2376 6960
rect 2416 6928 2448 6960
rect 2488 6928 2520 6960
rect 2560 6928 2592 6960
rect 2632 6928 2664 6960
rect 2704 6928 2736 6960
rect 2776 6928 2808 6960
rect 2848 6928 2880 6960
rect 2920 6928 2952 6960
rect 2992 6928 3024 6960
rect 3064 6928 3096 6960
rect 3136 6928 3168 6960
rect 3208 6928 3240 6960
rect 3280 6928 3312 6960
rect 3352 6928 3384 6960
rect 3424 6928 3456 6960
rect 3496 6928 3528 6960
rect 3568 6928 3600 6960
rect 3640 6928 3672 6960
rect 3712 6928 3744 6960
rect 3784 6928 3816 6960
rect 3856 6928 3888 6960
rect 3928 6928 3960 6960
rect 40 6856 72 6888
rect 112 6856 144 6888
rect 184 6856 216 6888
rect 256 6856 288 6888
rect 328 6856 360 6888
rect 400 6856 432 6888
rect 472 6856 504 6888
rect 544 6856 576 6888
rect 616 6856 648 6888
rect 688 6856 720 6888
rect 760 6856 792 6888
rect 832 6856 864 6888
rect 904 6856 936 6888
rect 976 6856 1008 6888
rect 1048 6856 1080 6888
rect 1120 6856 1152 6888
rect 1192 6856 1224 6888
rect 1264 6856 1296 6888
rect 1336 6856 1368 6888
rect 1408 6856 1440 6888
rect 1480 6856 1512 6888
rect 1552 6856 1584 6888
rect 1624 6856 1656 6888
rect 1696 6856 1728 6888
rect 1768 6856 1800 6888
rect 1840 6856 1872 6888
rect 1912 6856 1944 6888
rect 1984 6856 2016 6888
rect 2056 6856 2088 6888
rect 2128 6856 2160 6888
rect 2200 6856 2232 6888
rect 2272 6856 2304 6888
rect 2344 6856 2376 6888
rect 2416 6856 2448 6888
rect 2488 6856 2520 6888
rect 2560 6856 2592 6888
rect 2632 6856 2664 6888
rect 2704 6856 2736 6888
rect 2776 6856 2808 6888
rect 2848 6856 2880 6888
rect 2920 6856 2952 6888
rect 2992 6856 3024 6888
rect 3064 6856 3096 6888
rect 3136 6856 3168 6888
rect 3208 6856 3240 6888
rect 3280 6856 3312 6888
rect 3352 6856 3384 6888
rect 3424 6856 3456 6888
rect 3496 6856 3528 6888
rect 3568 6856 3600 6888
rect 3640 6856 3672 6888
rect 3712 6856 3744 6888
rect 3784 6856 3816 6888
rect 3856 6856 3888 6888
rect 3928 6856 3960 6888
rect 112 6512 144 6544
rect 184 6512 216 6544
rect 256 6512 288 6544
rect 328 6512 360 6544
rect 400 6512 432 6544
rect 472 6512 504 6544
rect 544 6512 576 6544
rect 616 6512 648 6544
rect 688 6512 720 6544
rect 760 6512 792 6544
rect 832 6512 864 6544
rect 904 6512 936 6544
rect 976 6512 1008 6544
rect 1048 6512 1080 6544
rect 1120 6512 1152 6544
rect 1192 6512 1224 6544
rect 1264 6512 1296 6544
rect 1336 6512 1368 6544
rect 1408 6512 1440 6544
rect 1480 6512 1512 6544
rect 1552 6512 1584 6544
rect 1624 6512 1656 6544
rect 1696 6512 1728 6544
rect 1768 6512 1800 6544
rect 1840 6512 1872 6544
rect 1912 6512 1944 6544
rect 1984 6512 2016 6544
rect 2056 6512 2088 6544
rect 2128 6512 2160 6544
rect 2200 6512 2232 6544
rect 2272 6512 2304 6544
rect 2344 6512 2376 6544
rect 2416 6512 2448 6544
rect 2488 6512 2520 6544
rect 2560 6512 2592 6544
rect 2632 6512 2664 6544
rect 2704 6512 2736 6544
rect 2776 6512 2808 6544
rect 2848 6512 2880 6544
rect 2920 6512 2952 6544
rect 2992 6512 3024 6544
rect 3064 6512 3096 6544
rect 3136 6512 3168 6544
rect 3208 6512 3240 6544
rect 3280 6512 3312 6544
rect 3352 6512 3384 6544
rect 3424 6512 3456 6544
rect 3496 6512 3528 6544
rect 3568 6512 3600 6544
rect 3640 6512 3672 6544
rect 3712 6512 3744 6544
rect 3784 6512 3816 6544
rect 3856 6512 3888 6544
rect 3928 6512 3960 6544
rect 40 6440 72 6472
rect 112 6440 144 6472
rect 184 6440 216 6472
rect 256 6440 288 6472
rect 328 6440 360 6472
rect 400 6440 432 6472
rect 472 6440 504 6472
rect 544 6440 576 6472
rect 616 6440 648 6472
rect 688 6440 720 6472
rect 760 6440 792 6472
rect 832 6440 864 6472
rect 904 6440 936 6472
rect 976 6440 1008 6472
rect 1048 6440 1080 6472
rect 1120 6440 1152 6472
rect 1192 6440 1224 6472
rect 1264 6440 1296 6472
rect 1336 6440 1368 6472
rect 1408 6440 1440 6472
rect 1480 6440 1512 6472
rect 1552 6440 1584 6472
rect 1624 6440 1656 6472
rect 1696 6440 1728 6472
rect 1768 6440 1800 6472
rect 1840 6440 1872 6472
rect 1912 6440 1944 6472
rect 1984 6440 2016 6472
rect 2056 6440 2088 6472
rect 2128 6440 2160 6472
rect 2200 6440 2232 6472
rect 2272 6440 2304 6472
rect 2344 6440 2376 6472
rect 2416 6440 2448 6472
rect 2488 6440 2520 6472
rect 2560 6440 2592 6472
rect 2632 6440 2664 6472
rect 2704 6440 2736 6472
rect 2776 6440 2808 6472
rect 2848 6440 2880 6472
rect 2920 6440 2952 6472
rect 2992 6440 3024 6472
rect 3064 6440 3096 6472
rect 3136 6440 3168 6472
rect 3208 6440 3240 6472
rect 3280 6440 3312 6472
rect 3352 6440 3384 6472
rect 3424 6440 3456 6472
rect 3496 6440 3528 6472
rect 3568 6440 3600 6472
rect 3640 6440 3672 6472
rect 3712 6440 3744 6472
rect 3784 6440 3816 6472
rect 3856 6440 3888 6472
rect 3928 6440 3960 6472
rect 40 6368 72 6400
rect 112 6368 144 6400
rect 184 6368 216 6400
rect 256 6368 288 6400
rect 328 6368 360 6400
rect 400 6368 432 6400
rect 472 6368 504 6400
rect 544 6368 576 6400
rect 616 6368 648 6400
rect 688 6368 720 6400
rect 760 6368 792 6400
rect 832 6368 864 6400
rect 904 6368 936 6400
rect 976 6368 1008 6400
rect 1048 6368 1080 6400
rect 1120 6368 1152 6400
rect 1192 6368 1224 6400
rect 1264 6368 1296 6400
rect 1336 6368 1368 6400
rect 1408 6368 1440 6400
rect 1480 6368 1512 6400
rect 1552 6368 1584 6400
rect 1624 6368 1656 6400
rect 1696 6368 1728 6400
rect 1768 6368 1800 6400
rect 1840 6368 1872 6400
rect 1912 6368 1944 6400
rect 1984 6368 2016 6400
rect 2056 6368 2088 6400
rect 2128 6368 2160 6400
rect 2200 6368 2232 6400
rect 2272 6368 2304 6400
rect 2344 6368 2376 6400
rect 2416 6368 2448 6400
rect 2488 6368 2520 6400
rect 2560 6368 2592 6400
rect 2632 6368 2664 6400
rect 2704 6368 2736 6400
rect 2776 6368 2808 6400
rect 2848 6368 2880 6400
rect 2920 6368 2952 6400
rect 2992 6368 3024 6400
rect 3064 6368 3096 6400
rect 3136 6368 3168 6400
rect 3208 6368 3240 6400
rect 3280 6368 3312 6400
rect 3352 6368 3384 6400
rect 3424 6368 3456 6400
rect 3496 6368 3528 6400
rect 3568 6368 3600 6400
rect 3640 6368 3672 6400
rect 3712 6368 3744 6400
rect 3784 6368 3816 6400
rect 3856 6368 3888 6400
rect 3928 6368 3960 6400
rect 40 6296 72 6328
rect 112 6296 144 6328
rect 184 6296 216 6328
rect 256 6296 288 6328
rect 328 6296 360 6328
rect 400 6296 432 6328
rect 472 6296 504 6328
rect 544 6296 576 6328
rect 616 6296 648 6328
rect 688 6296 720 6328
rect 760 6296 792 6328
rect 832 6296 864 6328
rect 904 6296 936 6328
rect 976 6296 1008 6328
rect 1048 6296 1080 6328
rect 1120 6296 1152 6328
rect 1192 6296 1224 6328
rect 1264 6296 1296 6328
rect 1336 6296 1368 6328
rect 1408 6296 1440 6328
rect 1480 6296 1512 6328
rect 1552 6296 1584 6328
rect 1624 6296 1656 6328
rect 1696 6296 1728 6328
rect 1768 6296 1800 6328
rect 1840 6296 1872 6328
rect 1912 6296 1944 6328
rect 1984 6296 2016 6328
rect 2056 6296 2088 6328
rect 2128 6296 2160 6328
rect 2200 6296 2232 6328
rect 2272 6296 2304 6328
rect 2344 6296 2376 6328
rect 2416 6296 2448 6328
rect 2488 6296 2520 6328
rect 2560 6296 2592 6328
rect 2632 6296 2664 6328
rect 2704 6296 2736 6328
rect 2776 6296 2808 6328
rect 2848 6296 2880 6328
rect 2920 6296 2952 6328
rect 2992 6296 3024 6328
rect 3064 6296 3096 6328
rect 3136 6296 3168 6328
rect 3208 6296 3240 6328
rect 3280 6296 3312 6328
rect 3352 6296 3384 6328
rect 3424 6296 3456 6328
rect 3496 6296 3528 6328
rect 3568 6296 3600 6328
rect 3640 6296 3672 6328
rect 3712 6296 3744 6328
rect 3784 6296 3816 6328
rect 3856 6296 3888 6328
rect 3928 6296 3960 6328
rect 40 6224 72 6256
rect 112 6224 144 6256
rect 184 6224 216 6256
rect 256 6224 288 6256
rect 328 6224 360 6256
rect 400 6224 432 6256
rect 472 6224 504 6256
rect 544 6224 576 6256
rect 616 6224 648 6256
rect 688 6224 720 6256
rect 760 6224 792 6256
rect 832 6224 864 6256
rect 904 6224 936 6256
rect 976 6224 1008 6256
rect 1048 6224 1080 6256
rect 1120 6224 1152 6256
rect 1192 6224 1224 6256
rect 1264 6224 1296 6256
rect 1336 6224 1368 6256
rect 1408 6224 1440 6256
rect 1480 6224 1512 6256
rect 1552 6224 1584 6256
rect 1624 6224 1656 6256
rect 1696 6224 1728 6256
rect 1768 6224 1800 6256
rect 1840 6224 1872 6256
rect 1912 6224 1944 6256
rect 1984 6224 2016 6256
rect 2056 6224 2088 6256
rect 2128 6224 2160 6256
rect 2200 6224 2232 6256
rect 2272 6224 2304 6256
rect 2344 6224 2376 6256
rect 2416 6224 2448 6256
rect 2488 6224 2520 6256
rect 2560 6224 2592 6256
rect 2632 6224 2664 6256
rect 2704 6224 2736 6256
rect 2776 6224 2808 6256
rect 2848 6224 2880 6256
rect 2920 6224 2952 6256
rect 2992 6224 3024 6256
rect 3064 6224 3096 6256
rect 3136 6224 3168 6256
rect 3208 6224 3240 6256
rect 3280 6224 3312 6256
rect 3352 6224 3384 6256
rect 3424 6224 3456 6256
rect 3496 6224 3528 6256
rect 3568 6224 3600 6256
rect 3640 6224 3672 6256
rect 3712 6224 3744 6256
rect 3784 6224 3816 6256
rect 3856 6224 3888 6256
rect 3928 6224 3960 6256
rect 40 6152 72 6184
rect 112 6152 144 6184
rect 184 6152 216 6184
rect 256 6152 288 6184
rect 328 6152 360 6184
rect 400 6152 432 6184
rect 472 6152 504 6184
rect 544 6152 576 6184
rect 616 6152 648 6184
rect 688 6152 720 6184
rect 760 6152 792 6184
rect 832 6152 864 6184
rect 904 6152 936 6184
rect 976 6152 1008 6184
rect 1048 6152 1080 6184
rect 1120 6152 1152 6184
rect 1192 6152 1224 6184
rect 1264 6152 1296 6184
rect 1336 6152 1368 6184
rect 1408 6152 1440 6184
rect 1480 6152 1512 6184
rect 1552 6152 1584 6184
rect 1624 6152 1656 6184
rect 1696 6152 1728 6184
rect 1768 6152 1800 6184
rect 1840 6152 1872 6184
rect 1912 6152 1944 6184
rect 1984 6152 2016 6184
rect 2056 6152 2088 6184
rect 2128 6152 2160 6184
rect 2200 6152 2232 6184
rect 2272 6152 2304 6184
rect 2344 6152 2376 6184
rect 2416 6152 2448 6184
rect 2488 6152 2520 6184
rect 2560 6152 2592 6184
rect 2632 6152 2664 6184
rect 2704 6152 2736 6184
rect 2776 6152 2808 6184
rect 2848 6152 2880 6184
rect 2920 6152 2952 6184
rect 2992 6152 3024 6184
rect 3064 6152 3096 6184
rect 3136 6152 3168 6184
rect 3208 6152 3240 6184
rect 3280 6152 3312 6184
rect 3352 6152 3384 6184
rect 3424 6152 3456 6184
rect 3496 6152 3528 6184
rect 3568 6152 3600 6184
rect 3640 6152 3672 6184
rect 3712 6152 3744 6184
rect 3784 6152 3816 6184
rect 3856 6152 3888 6184
rect 3928 6152 3960 6184
rect 40 6080 72 6112
rect 112 6080 144 6112
rect 184 6080 216 6112
rect 256 6080 288 6112
rect 328 6080 360 6112
rect 400 6080 432 6112
rect 472 6080 504 6112
rect 544 6080 576 6112
rect 616 6080 648 6112
rect 688 6080 720 6112
rect 760 6080 792 6112
rect 832 6080 864 6112
rect 904 6080 936 6112
rect 976 6080 1008 6112
rect 1048 6080 1080 6112
rect 1120 6080 1152 6112
rect 1192 6080 1224 6112
rect 1264 6080 1296 6112
rect 1336 6080 1368 6112
rect 1408 6080 1440 6112
rect 1480 6080 1512 6112
rect 1552 6080 1584 6112
rect 1624 6080 1656 6112
rect 1696 6080 1728 6112
rect 1768 6080 1800 6112
rect 1840 6080 1872 6112
rect 1912 6080 1944 6112
rect 1984 6080 2016 6112
rect 2056 6080 2088 6112
rect 2128 6080 2160 6112
rect 2200 6080 2232 6112
rect 2272 6080 2304 6112
rect 2344 6080 2376 6112
rect 2416 6080 2448 6112
rect 2488 6080 2520 6112
rect 2560 6080 2592 6112
rect 2632 6080 2664 6112
rect 2704 6080 2736 6112
rect 2776 6080 2808 6112
rect 2848 6080 2880 6112
rect 2920 6080 2952 6112
rect 2992 6080 3024 6112
rect 3064 6080 3096 6112
rect 3136 6080 3168 6112
rect 3208 6080 3240 6112
rect 3280 6080 3312 6112
rect 3352 6080 3384 6112
rect 3424 6080 3456 6112
rect 3496 6080 3528 6112
rect 3568 6080 3600 6112
rect 3640 6080 3672 6112
rect 3712 6080 3744 6112
rect 3784 6080 3816 6112
rect 3856 6080 3888 6112
rect 3928 6080 3960 6112
rect 40 6008 72 6040
rect 112 6008 144 6040
rect 184 6008 216 6040
rect 256 6008 288 6040
rect 328 6008 360 6040
rect 400 6008 432 6040
rect 472 6008 504 6040
rect 544 6008 576 6040
rect 616 6008 648 6040
rect 688 6008 720 6040
rect 760 6008 792 6040
rect 832 6008 864 6040
rect 904 6008 936 6040
rect 976 6008 1008 6040
rect 1048 6008 1080 6040
rect 1120 6008 1152 6040
rect 1192 6008 1224 6040
rect 1264 6008 1296 6040
rect 1336 6008 1368 6040
rect 1408 6008 1440 6040
rect 1480 6008 1512 6040
rect 1552 6008 1584 6040
rect 1624 6008 1656 6040
rect 1696 6008 1728 6040
rect 1768 6008 1800 6040
rect 1840 6008 1872 6040
rect 1912 6008 1944 6040
rect 1984 6008 2016 6040
rect 2056 6008 2088 6040
rect 2128 6008 2160 6040
rect 2200 6008 2232 6040
rect 2272 6008 2304 6040
rect 2344 6008 2376 6040
rect 2416 6008 2448 6040
rect 2488 6008 2520 6040
rect 2560 6008 2592 6040
rect 2632 6008 2664 6040
rect 2704 6008 2736 6040
rect 2776 6008 2808 6040
rect 2848 6008 2880 6040
rect 2920 6008 2952 6040
rect 2992 6008 3024 6040
rect 3064 6008 3096 6040
rect 3136 6008 3168 6040
rect 3208 6008 3240 6040
rect 3280 6008 3312 6040
rect 3352 6008 3384 6040
rect 3424 6008 3456 6040
rect 3496 6008 3528 6040
rect 3568 6008 3600 6040
rect 3640 6008 3672 6040
rect 3712 6008 3744 6040
rect 3784 6008 3816 6040
rect 3856 6008 3888 6040
rect 3928 6008 3960 6040
rect 40 5936 72 5968
rect 112 5936 144 5968
rect 184 5936 216 5968
rect 256 5936 288 5968
rect 328 5936 360 5968
rect 400 5936 432 5968
rect 472 5936 504 5968
rect 544 5936 576 5968
rect 616 5936 648 5968
rect 688 5936 720 5968
rect 760 5936 792 5968
rect 832 5936 864 5968
rect 904 5936 936 5968
rect 976 5936 1008 5968
rect 1048 5936 1080 5968
rect 1120 5936 1152 5968
rect 1192 5936 1224 5968
rect 1264 5936 1296 5968
rect 1336 5936 1368 5968
rect 1408 5936 1440 5968
rect 1480 5936 1512 5968
rect 1552 5936 1584 5968
rect 1624 5936 1656 5968
rect 1696 5936 1728 5968
rect 1768 5936 1800 5968
rect 1840 5936 1872 5968
rect 1912 5936 1944 5968
rect 1984 5936 2016 5968
rect 2056 5936 2088 5968
rect 2128 5936 2160 5968
rect 2200 5936 2232 5968
rect 2272 5936 2304 5968
rect 2344 5936 2376 5968
rect 2416 5936 2448 5968
rect 2488 5936 2520 5968
rect 2560 5936 2592 5968
rect 2632 5936 2664 5968
rect 2704 5936 2736 5968
rect 2776 5936 2808 5968
rect 2848 5936 2880 5968
rect 2920 5936 2952 5968
rect 2992 5936 3024 5968
rect 3064 5936 3096 5968
rect 3136 5936 3168 5968
rect 3208 5936 3240 5968
rect 3280 5936 3312 5968
rect 3352 5936 3384 5968
rect 3424 5936 3456 5968
rect 3496 5936 3528 5968
rect 3568 5936 3600 5968
rect 3640 5936 3672 5968
rect 3712 5936 3744 5968
rect 3784 5936 3816 5968
rect 3856 5936 3888 5968
rect 3928 5936 3960 5968
rect 40 5864 72 5896
rect 112 5864 144 5896
rect 184 5864 216 5896
rect 256 5864 288 5896
rect 328 5864 360 5896
rect 400 5864 432 5896
rect 472 5864 504 5896
rect 544 5864 576 5896
rect 616 5864 648 5896
rect 688 5864 720 5896
rect 760 5864 792 5896
rect 832 5864 864 5896
rect 904 5864 936 5896
rect 976 5864 1008 5896
rect 1048 5864 1080 5896
rect 1120 5864 1152 5896
rect 1192 5864 1224 5896
rect 1264 5864 1296 5896
rect 1336 5864 1368 5896
rect 1408 5864 1440 5896
rect 1480 5864 1512 5896
rect 1552 5864 1584 5896
rect 1624 5864 1656 5896
rect 1696 5864 1728 5896
rect 1768 5864 1800 5896
rect 1840 5864 1872 5896
rect 1912 5864 1944 5896
rect 1984 5864 2016 5896
rect 2056 5864 2088 5896
rect 2128 5864 2160 5896
rect 2200 5864 2232 5896
rect 2272 5864 2304 5896
rect 2344 5864 2376 5896
rect 2416 5864 2448 5896
rect 2488 5864 2520 5896
rect 2560 5864 2592 5896
rect 2632 5864 2664 5896
rect 2704 5864 2736 5896
rect 2776 5864 2808 5896
rect 2848 5864 2880 5896
rect 2920 5864 2952 5896
rect 2992 5864 3024 5896
rect 3064 5864 3096 5896
rect 3136 5864 3168 5896
rect 3208 5864 3240 5896
rect 3280 5864 3312 5896
rect 3352 5864 3384 5896
rect 3424 5864 3456 5896
rect 3496 5864 3528 5896
rect 3568 5864 3600 5896
rect 3640 5864 3672 5896
rect 3712 5864 3744 5896
rect 3784 5864 3816 5896
rect 3856 5864 3888 5896
rect 3928 5864 3960 5896
rect 40 5792 72 5824
rect 112 5792 144 5824
rect 184 5792 216 5824
rect 256 5792 288 5824
rect 328 5792 360 5824
rect 400 5792 432 5824
rect 472 5792 504 5824
rect 544 5792 576 5824
rect 616 5792 648 5824
rect 688 5792 720 5824
rect 760 5792 792 5824
rect 832 5792 864 5824
rect 904 5792 936 5824
rect 976 5792 1008 5824
rect 1048 5792 1080 5824
rect 1120 5792 1152 5824
rect 1192 5792 1224 5824
rect 1264 5792 1296 5824
rect 1336 5792 1368 5824
rect 1408 5792 1440 5824
rect 1480 5792 1512 5824
rect 1552 5792 1584 5824
rect 1624 5792 1656 5824
rect 1696 5792 1728 5824
rect 1768 5792 1800 5824
rect 1840 5792 1872 5824
rect 1912 5792 1944 5824
rect 1984 5792 2016 5824
rect 2056 5792 2088 5824
rect 2128 5792 2160 5824
rect 2200 5792 2232 5824
rect 2272 5792 2304 5824
rect 2344 5792 2376 5824
rect 2416 5792 2448 5824
rect 2488 5792 2520 5824
rect 2560 5792 2592 5824
rect 2632 5792 2664 5824
rect 2704 5792 2736 5824
rect 2776 5792 2808 5824
rect 2848 5792 2880 5824
rect 2920 5792 2952 5824
rect 2992 5792 3024 5824
rect 3064 5792 3096 5824
rect 3136 5792 3168 5824
rect 3208 5792 3240 5824
rect 3280 5792 3312 5824
rect 3352 5792 3384 5824
rect 3424 5792 3456 5824
rect 3496 5792 3528 5824
rect 3568 5792 3600 5824
rect 3640 5792 3672 5824
rect 3712 5792 3744 5824
rect 3784 5792 3816 5824
rect 3856 5792 3888 5824
rect 3928 5792 3960 5824
rect 40 5720 72 5752
rect 112 5720 144 5752
rect 184 5720 216 5752
rect 256 5720 288 5752
rect 328 5720 360 5752
rect 400 5720 432 5752
rect 472 5720 504 5752
rect 544 5720 576 5752
rect 616 5720 648 5752
rect 688 5720 720 5752
rect 760 5720 792 5752
rect 832 5720 864 5752
rect 904 5720 936 5752
rect 976 5720 1008 5752
rect 1048 5720 1080 5752
rect 1120 5720 1152 5752
rect 1192 5720 1224 5752
rect 1264 5720 1296 5752
rect 1336 5720 1368 5752
rect 1408 5720 1440 5752
rect 1480 5720 1512 5752
rect 1552 5720 1584 5752
rect 1624 5720 1656 5752
rect 1696 5720 1728 5752
rect 1768 5720 1800 5752
rect 1840 5720 1872 5752
rect 1912 5720 1944 5752
rect 1984 5720 2016 5752
rect 2056 5720 2088 5752
rect 2128 5720 2160 5752
rect 2200 5720 2232 5752
rect 2272 5720 2304 5752
rect 2344 5720 2376 5752
rect 2416 5720 2448 5752
rect 2488 5720 2520 5752
rect 2560 5720 2592 5752
rect 2632 5720 2664 5752
rect 2704 5720 2736 5752
rect 2776 5720 2808 5752
rect 2848 5720 2880 5752
rect 2920 5720 2952 5752
rect 2992 5720 3024 5752
rect 3064 5720 3096 5752
rect 3136 5720 3168 5752
rect 3208 5720 3240 5752
rect 3280 5720 3312 5752
rect 3352 5720 3384 5752
rect 3424 5720 3456 5752
rect 3496 5720 3528 5752
rect 3568 5720 3600 5752
rect 3640 5720 3672 5752
rect 3712 5720 3744 5752
rect 3784 5720 3816 5752
rect 3856 5720 3888 5752
rect 3928 5720 3960 5752
rect 40 5648 72 5680
rect 112 5648 144 5680
rect 184 5648 216 5680
rect 256 5648 288 5680
rect 328 5648 360 5680
rect 400 5648 432 5680
rect 472 5648 504 5680
rect 544 5648 576 5680
rect 616 5648 648 5680
rect 688 5648 720 5680
rect 760 5648 792 5680
rect 832 5648 864 5680
rect 904 5648 936 5680
rect 976 5648 1008 5680
rect 1048 5648 1080 5680
rect 1120 5648 1152 5680
rect 1192 5648 1224 5680
rect 1264 5648 1296 5680
rect 1336 5648 1368 5680
rect 1408 5648 1440 5680
rect 1480 5648 1512 5680
rect 1552 5648 1584 5680
rect 1624 5648 1656 5680
rect 1696 5648 1728 5680
rect 1768 5648 1800 5680
rect 1840 5648 1872 5680
rect 1912 5648 1944 5680
rect 1984 5648 2016 5680
rect 2056 5648 2088 5680
rect 2128 5648 2160 5680
rect 2200 5648 2232 5680
rect 2272 5648 2304 5680
rect 2344 5648 2376 5680
rect 2416 5648 2448 5680
rect 2488 5648 2520 5680
rect 2560 5648 2592 5680
rect 2632 5648 2664 5680
rect 2704 5648 2736 5680
rect 2776 5648 2808 5680
rect 2848 5648 2880 5680
rect 2920 5648 2952 5680
rect 2992 5648 3024 5680
rect 3064 5648 3096 5680
rect 3136 5648 3168 5680
rect 3208 5648 3240 5680
rect 3280 5648 3312 5680
rect 3352 5648 3384 5680
rect 3424 5648 3456 5680
rect 3496 5648 3528 5680
rect 3568 5648 3600 5680
rect 3640 5648 3672 5680
rect 3712 5648 3744 5680
rect 3784 5648 3816 5680
rect 3856 5648 3888 5680
rect 3928 5648 3960 5680
rect 40 5576 72 5608
rect 112 5576 144 5608
rect 184 5576 216 5608
rect 256 5576 288 5608
rect 328 5576 360 5608
rect 400 5576 432 5608
rect 472 5576 504 5608
rect 544 5576 576 5608
rect 616 5576 648 5608
rect 688 5576 720 5608
rect 760 5576 792 5608
rect 832 5576 864 5608
rect 904 5576 936 5608
rect 976 5576 1008 5608
rect 1048 5576 1080 5608
rect 1120 5576 1152 5608
rect 1192 5576 1224 5608
rect 1264 5576 1296 5608
rect 1336 5576 1368 5608
rect 1408 5576 1440 5608
rect 1480 5576 1512 5608
rect 1552 5576 1584 5608
rect 1624 5576 1656 5608
rect 1696 5576 1728 5608
rect 1768 5576 1800 5608
rect 1840 5576 1872 5608
rect 1912 5576 1944 5608
rect 1984 5576 2016 5608
rect 2056 5576 2088 5608
rect 2128 5576 2160 5608
rect 2200 5576 2232 5608
rect 2272 5576 2304 5608
rect 2344 5576 2376 5608
rect 2416 5576 2448 5608
rect 2488 5576 2520 5608
rect 2560 5576 2592 5608
rect 2632 5576 2664 5608
rect 2704 5576 2736 5608
rect 2776 5576 2808 5608
rect 2848 5576 2880 5608
rect 2920 5576 2952 5608
rect 2992 5576 3024 5608
rect 3064 5576 3096 5608
rect 3136 5576 3168 5608
rect 3208 5576 3240 5608
rect 3280 5576 3312 5608
rect 3352 5576 3384 5608
rect 3424 5576 3456 5608
rect 3496 5576 3528 5608
rect 3568 5576 3600 5608
rect 3640 5576 3672 5608
rect 3712 5576 3744 5608
rect 3784 5576 3816 5608
rect 3856 5576 3888 5608
rect 3928 5576 3960 5608
rect 40 5504 72 5536
rect 112 5504 144 5536
rect 184 5504 216 5536
rect 256 5504 288 5536
rect 328 5504 360 5536
rect 400 5504 432 5536
rect 472 5504 504 5536
rect 544 5504 576 5536
rect 616 5504 648 5536
rect 688 5504 720 5536
rect 760 5504 792 5536
rect 832 5504 864 5536
rect 904 5504 936 5536
rect 976 5504 1008 5536
rect 1048 5504 1080 5536
rect 1120 5504 1152 5536
rect 1192 5504 1224 5536
rect 1264 5504 1296 5536
rect 1336 5504 1368 5536
rect 1408 5504 1440 5536
rect 1480 5504 1512 5536
rect 1552 5504 1584 5536
rect 1624 5504 1656 5536
rect 1696 5504 1728 5536
rect 1768 5504 1800 5536
rect 1840 5504 1872 5536
rect 1912 5504 1944 5536
rect 1984 5504 2016 5536
rect 2056 5504 2088 5536
rect 2128 5504 2160 5536
rect 2200 5504 2232 5536
rect 2272 5504 2304 5536
rect 2344 5504 2376 5536
rect 2416 5504 2448 5536
rect 2488 5504 2520 5536
rect 2560 5504 2592 5536
rect 2632 5504 2664 5536
rect 2704 5504 2736 5536
rect 2776 5504 2808 5536
rect 2848 5504 2880 5536
rect 2920 5504 2952 5536
rect 2992 5504 3024 5536
rect 3064 5504 3096 5536
rect 3136 5504 3168 5536
rect 3208 5504 3240 5536
rect 3280 5504 3312 5536
rect 3352 5504 3384 5536
rect 3424 5504 3456 5536
rect 3496 5504 3528 5536
rect 3568 5504 3600 5536
rect 3640 5504 3672 5536
rect 3712 5504 3744 5536
rect 3784 5504 3816 5536
rect 3856 5504 3888 5536
rect 3928 5504 3960 5536
rect 40 5432 72 5464
rect 112 5432 144 5464
rect 184 5432 216 5464
rect 256 5432 288 5464
rect 328 5432 360 5464
rect 400 5432 432 5464
rect 472 5432 504 5464
rect 544 5432 576 5464
rect 616 5432 648 5464
rect 688 5432 720 5464
rect 760 5432 792 5464
rect 832 5432 864 5464
rect 904 5432 936 5464
rect 976 5432 1008 5464
rect 1048 5432 1080 5464
rect 1120 5432 1152 5464
rect 1192 5432 1224 5464
rect 1264 5432 1296 5464
rect 1336 5432 1368 5464
rect 1408 5432 1440 5464
rect 1480 5432 1512 5464
rect 1552 5432 1584 5464
rect 1624 5432 1656 5464
rect 1696 5432 1728 5464
rect 1768 5432 1800 5464
rect 1840 5432 1872 5464
rect 1912 5432 1944 5464
rect 1984 5432 2016 5464
rect 2056 5432 2088 5464
rect 2128 5432 2160 5464
rect 2200 5432 2232 5464
rect 2272 5432 2304 5464
rect 2344 5432 2376 5464
rect 2416 5432 2448 5464
rect 2488 5432 2520 5464
rect 2560 5432 2592 5464
rect 2632 5432 2664 5464
rect 2704 5432 2736 5464
rect 2776 5432 2808 5464
rect 2848 5432 2880 5464
rect 2920 5432 2952 5464
rect 2992 5432 3024 5464
rect 3064 5432 3096 5464
rect 3136 5432 3168 5464
rect 3208 5432 3240 5464
rect 3280 5432 3312 5464
rect 3352 5432 3384 5464
rect 3424 5432 3456 5464
rect 3496 5432 3528 5464
rect 3568 5432 3600 5464
rect 3640 5432 3672 5464
rect 3712 5432 3744 5464
rect 3784 5432 3816 5464
rect 3856 5432 3888 5464
rect 3928 5432 3960 5464
rect 40 5360 72 5392
rect 112 5360 144 5392
rect 184 5360 216 5392
rect 256 5360 288 5392
rect 328 5360 360 5392
rect 400 5360 432 5392
rect 472 5360 504 5392
rect 544 5360 576 5392
rect 616 5360 648 5392
rect 688 5360 720 5392
rect 760 5360 792 5392
rect 832 5360 864 5392
rect 904 5360 936 5392
rect 976 5360 1008 5392
rect 1048 5360 1080 5392
rect 1120 5360 1152 5392
rect 1192 5360 1224 5392
rect 1264 5360 1296 5392
rect 1336 5360 1368 5392
rect 1408 5360 1440 5392
rect 1480 5360 1512 5392
rect 1552 5360 1584 5392
rect 1624 5360 1656 5392
rect 1696 5360 1728 5392
rect 1768 5360 1800 5392
rect 1840 5360 1872 5392
rect 1912 5360 1944 5392
rect 1984 5360 2016 5392
rect 2056 5360 2088 5392
rect 2128 5360 2160 5392
rect 2200 5360 2232 5392
rect 2272 5360 2304 5392
rect 2344 5360 2376 5392
rect 2416 5360 2448 5392
rect 2488 5360 2520 5392
rect 2560 5360 2592 5392
rect 2632 5360 2664 5392
rect 2704 5360 2736 5392
rect 2776 5360 2808 5392
rect 2848 5360 2880 5392
rect 2920 5360 2952 5392
rect 2992 5360 3024 5392
rect 3064 5360 3096 5392
rect 3136 5360 3168 5392
rect 3208 5360 3240 5392
rect 3280 5360 3312 5392
rect 3352 5360 3384 5392
rect 3424 5360 3456 5392
rect 3496 5360 3528 5392
rect 3568 5360 3600 5392
rect 3640 5360 3672 5392
rect 3712 5360 3744 5392
rect 3784 5360 3816 5392
rect 3856 5360 3888 5392
rect 3928 5360 3960 5392
rect 40 5288 72 5320
rect 112 5288 144 5320
rect 184 5288 216 5320
rect 256 5288 288 5320
rect 328 5288 360 5320
rect 400 5288 432 5320
rect 472 5288 504 5320
rect 544 5288 576 5320
rect 616 5288 648 5320
rect 688 5288 720 5320
rect 760 5288 792 5320
rect 832 5288 864 5320
rect 904 5288 936 5320
rect 976 5288 1008 5320
rect 1048 5288 1080 5320
rect 1120 5288 1152 5320
rect 1192 5288 1224 5320
rect 1264 5288 1296 5320
rect 1336 5288 1368 5320
rect 1408 5288 1440 5320
rect 1480 5288 1512 5320
rect 1552 5288 1584 5320
rect 1624 5288 1656 5320
rect 1696 5288 1728 5320
rect 1768 5288 1800 5320
rect 1840 5288 1872 5320
rect 1912 5288 1944 5320
rect 1984 5288 2016 5320
rect 2056 5288 2088 5320
rect 2128 5288 2160 5320
rect 2200 5288 2232 5320
rect 2272 5288 2304 5320
rect 2344 5288 2376 5320
rect 2416 5288 2448 5320
rect 2488 5288 2520 5320
rect 2560 5288 2592 5320
rect 2632 5288 2664 5320
rect 2704 5288 2736 5320
rect 2776 5288 2808 5320
rect 2848 5288 2880 5320
rect 2920 5288 2952 5320
rect 2992 5288 3024 5320
rect 3064 5288 3096 5320
rect 3136 5288 3168 5320
rect 3208 5288 3240 5320
rect 3280 5288 3312 5320
rect 3352 5288 3384 5320
rect 3424 5288 3456 5320
rect 3496 5288 3528 5320
rect 3568 5288 3600 5320
rect 3640 5288 3672 5320
rect 3712 5288 3744 5320
rect 3784 5288 3816 5320
rect 3856 5288 3888 5320
rect 3928 5288 3960 5320
rect 40 5216 72 5248
rect 112 5216 144 5248
rect 184 5216 216 5248
rect 256 5216 288 5248
rect 328 5216 360 5248
rect 400 5216 432 5248
rect 472 5216 504 5248
rect 544 5216 576 5248
rect 616 5216 648 5248
rect 688 5216 720 5248
rect 760 5216 792 5248
rect 832 5216 864 5248
rect 904 5216 936 5248
rect 976 5216 1008 5248
rect 1048 5216 1080 5248
rect 1120 5216 1152 5248
rect 1192 5216 1224 5248
rect 1264 5216 1296 5248
rect 1336 5216 1368 5248
rect 1408 5216 1440 5248
rect 1480 5216 1512 5248
rect 1552 5216 1584 5248
rect 1624 5216 1656 5248
rect 1696 5216 1728 5248
rect 1768 5216 1800 5248
rect 1840 5216 1872 5248
rect 1912 5216 1944 5248
rect 1984 5216 2016 5248
rect 2056 5216 2088 5248
rect 2128 5216 2160 5248
rect 2200 5216 2232 5248
rect 2272 5216 2304 5248
rect 2344 5216 2376 5248
rect 2416 5216 2448 5248
rect 2488 5216 2520 5248
rect 2560 5216 2592 5248
rect 2632 5216 2664 5248
rect 2704 5216 2736 5248
rect 2776 5216 2808 5248
rect 2848 5216 2880 5248
rect 2920 5216 2952 5248
rect 2992 5216 3024 5248
rect 3064 5216 3096 5248
rect 3136 5216 3168 5248
rect 3208 5216 3240 5248
rect 3280 5216 3312 5248
rect 3352 5216 3384 5248
rect 3424 5216 3456 5248
rect 3496 5216 3528 5248
rect 3568 5216 3600 5248
rect 3640 5216 3672 5248
rect 3712 5216 3744 5248
rect 3784 5216 3816 5248
rect 3856 5216 3888 5248
rect 3928 5216 3960 5248
rect 40 5144 72 5176
rect 112 5144 144 5176
rect 184 5144 216 5176
rect 256 5144 288 5176
rect 328 5144 360 5176
rect 400 5144 432 5176
rect 472 5144 504 5176
rect 544 5144 576 5176
rect 616 5144 648 5176
rect 688 5144 720 5176
rect 760 5144 792 5176
rect 832 5144 864 5176
rect 904 5144 936 5176
rect 976 5144 1008 5176
rect 1048 5144 1080 5176
rect 1120 5144 1152 5176
rect 1192 5144 1224 5176
rect 1264 5144 1296 5176
rect 1336 5144 1368 5176
rect 1408 5144 1440 5176
rect 1480 5144 1512 5176
rect 1552 5144 1584 5176
rect 1624 5144 1656 5176
rect 1696 5144 1728 5176
rect 1768 5144 1800 5176
rect 1840 5144 1872 5176
rect 1912 5144 1944 5176
rect 1984 5144 2016 5176
rect 2056 5144 2088 5176
rect 2128 5144 2160 5176
rect 2200 5144 2232 5176
rect 2272 5144 2304 5176
rect 2344 5144 2376 5176
rect 2416 5144 2448 5176
rect 2488 5144 2520 5176
rect 2560 5144 2592 5176
rect 2632 5144 2664 5176
rect 2704 5144 2736 5176
rect 2776 5144 2808 5176
rect 2848 5144 2880 5176
rect 2920 5144 2952 5176
rect 2992 5144 3024 5176
rect 3064 5144 3096 5176
rect 3136 5144 3168 5176
rect 3208 5144 3240 5176
rect 3280 5144 3312 5176
rect 3352 5144 3384 5176
rect 3424 5144 3456 5176
rect 3496 5144 3528 5176
rect 3568 5144 3600 5176
rect 3640 5144 3672 5176
rect 3712 5144 3744 5176
rect 3784 5144 3816 5176
rect 3856 5144 3888 5176
rect 3928 5144 3960 5176
rect 40 5072 72 5104
rect 112 5072 144 5104
rect 184 5072 216 5104
rect 256 5072 288 5104
rect 328 5072 360 5104
rect 400 5072 432 5104
rect 472 5072 504 5104
rect 544 5072 576 5104
rect 616 5072 648 5104
rect 688 5072 720 5104
rect 760 5072 792 5104
rect 832 5072 864 5104
rect 904 5072 936 5104
rect 976 5072 1008 5104
rect 1048 5072 1080 5104
rect 1120 5072 1152 5104
rect 1192 5072 1224 5104
rect 1264 5072 1296 5104
rect 1336 5072 1368 5104
rect 1408 5072 1440 5104
rect 1480 5072 1512 5104
rect 1552 5072 1584 5104
rect 1624 5072 1656 5104
rect 1696 5072 1728 5104
rect 1768 5072 1800 5104
rect 1840 5072 1872 5104
rect 1912 5072 1944 5104
rect 1984 5072 2016 5104
rect 2056 5072 2088 5104
rect 2128 5072 2160 5104
rect 2200 5072 2232 5104
rect 2272 5072 2304 5104
rect 2344 5072 2376 5104
rect 2416 5072 2448 5104
rect 2488 5072 2520 5104
rect 2560 5072 2592 5104
rect 2632 5072 2664 5104
rect 2704 5072 2736 5104
rect 2776 5072 2808 5104
rect 2848 5072 2880 5104
rect 2920 5072 2952 5104
rect 2992 5072 3024 5104
rect 3064 5072 3096 5104
rect 3136 5072 3168 5104
rect 3208 5072 3240 5104
rect 3280 5072 3312 5104
rect 3352 5072 3384 5104
rect 3424 5072 3456 5104
rect 3496 5072 3528 5104
rect 3568 5072 3600 5104
rect 3640 5072 3672 5104
rect 3712 5072 3744 5104
rect 3784 5072 3816 5104
rect 3856 5072 3888 5104
rect 3928 5072 3960 5104
rect 40 5000 72 5032
rect 112 5000 144 5032
rect 184 5000 216 5032
rect 256 5000 288 5032
rect 328 5000 360 5032
rect 400 5000 432 5032
rect 472 5000 504 5032
rect 544 5000 576 5032
rect 616 5000 648 5032
rect 688 5000 720 5032
rect 760 5000 792 5032
rect 832 5000 864 5032
rect 904 5000 936 5032
rect 976 5000 1008 5032
rect 1048 5000 1080 5032
rect 1120 5000 1152 5032
rect 1192 5000 1224 5032
rect 1264 5000 1296 5032
rect 1336 5000 1368 5032
rect 1408 5000 1440 5032
rect 1480 5000 1512 5032
rect 1552 5000 1584 5032
rect 1624 5000 1656 5032
rect 1696 5000 1728 5032
rect 1768 5000 1800 5032
rect 1840 5000 1872 5032
rect 1912 5000 1944 5032
rect 1984 5000 2016 5032
rect 2056 5000 2088 5032
rect 2128 5000 2160 5032
rect 2200 5000 2232 5032
rect 2272 5000 2304 5032
rect 2344 5000 2376 5032
rect 2416 5000 2448 5032
rect 2488 5000 2520 5032
rect 2560 5000 2592 5032
rect 2632 5000 2664 5032
rect 2704 5000 2736 5032
rect 2776 5000 2808 5032
rect 2848 5000 2880 5032
rect 2920 5000 2952 5032
rect 2992 5000 3024 5032
rect 3064 5000 3096 5032
rect 3136 5000 3168 5032
rect 3208 5000 3240 5032
rect 3280 5000 3312 5032
rect 3352 5000 3384 5032
rect 3424 5000 3456 5032
rect 3496 5000 3528 5032
rect 3568 5000 3600 5032
rect 3640 5000 3672 5032
rect 3712 5000 3744 5032
rect 3784 5000 3816 5032
rect 3856 5000 3888 5032
rect 3928 5000 3960 5032
rect 40 4928 72 4960
rect 112 4928 144 4960
rect 184 4928 216 4960
rect 256 4928 288 4960
rect 328 4928 360 4960
rect 400 4928 432 4960
rect 472 4928 504 4960
rect 544 4928 576 4960
rect 616 4928 648 4960
rect 688 4928 720 4960
rect 760 4928 792 4960
rect 832 4928 864 4960
rect 904 4928 936 4960
rect 976 4928 1008 4960
rect 1048 4928 1080 4960
rect 1120 4928 1152 4960
rect 1192 4928 1224 4960
rect 1264 4928 1296 4960
rect 1336 4928 1368 4960
rect 1408 4928 1440 4960
rect 1480 4928 1512 4960
rect 1552 4928 1584 4960
rect 1624 4928 1656 4960
rect 1696 4928 1728 4960
rect 1768 4928 1800 4960
rect 1840 4928 1872 4960
rect 1912 4928 1944 4960
rect 1984 4928 2016 4960
rect 2056 4928 2088 4960
rect 2128 4928 2160 4960
rect 2200 4928 2232 4960
rect 2272 4928 2304 4960
rect 2344 4928 2376 4960
rect 2416 4928 2448 4960
rect 2488 4928 2520 4960
rect 2560 4928 2592 4960
rect 2632 4928 2664 4960
rect 2704 4928 2736 4960
rect 2776 4928 2808 4960
rect 2848 4928 2880 4960
rect 2920 4928 2952 4960
rect 2992 4928 3024 4960
rect 3064 4928 3096 4960
rect 3136 4928 3168 4960
rect 3208 4928 3240 4960
rect 3280 4928 3312 4960
rect 3352 4928 3384 4960
rect 3424 4928 3456 4960
rect 3496 4928 3528 4960
rect 3568 4928 3600 4960
rect 3640 4928 3672 4960
rect 3712 4928 3744 4960
rect 3784 4928 3816 4960
rect 3856 4928 3888 4960
rect 3928 4928 3960 4960
rect 40 4856 72 4888
rect 112 4856 144 4888
rect 184 4856 216 4888
rect 256 4856 288 4888
rect 328 4856 360 4888
rect 400 4856 432 4888
rect 472 4856 504 4888
rect 544 4856 576 4888
rect 616 4856 648 4888
rect 688 4856 720 4888
rect 760 4856 792 4888
rect 832 4856 864 4888
rect 904 4856 936 4888
rect 976 4856 1008 4888
rect 1048 4856 1080 4888
rect 1120 4856 1152 4888
rect 1192 4856 1224 4888
rect 1264 4856 1296 4888
rect 1336 4856 1368 4888
rect 1408 4856 1440 4888
rect 1480 4856 1512 4888
rect 1552 4856 1584 4888
rect 1624 4856 1656 4888
rect 1696 4856 1728 4888
rect 1768 4856 1800 4888
rect 1840 4856 1872 4888
rect 1912 4856 1944 4888
rect 1984 4856 2016 4888
rect 2056 4856 2088 4888
rect 2128 4856 2160 4888
rect 2200 4856 2232 4888
rect 2272 4856 2304 4888
rect 2344 4856 2376 4888
rect 2416 4856 2448 4888
rect 2488 4856 2520 4888
rect 2560 4856 2592 4888
rect 2632 4856 2664 4888
rect 2704 4856 2736 4888
rect 2776 4856 2808 4888
rect 2848 4856 2880 4888
rect 2920 4856 2952 4888
rect 2992 4856 3024 4888
rect 3064 4856 3096 4888
rect 3136 4856 3168 4888
rect 3208 4856 3240 4888
rect 3280 4856 3312 4888
rect 3352 4856 3384 4888
rect 3424 4856 3456 4888
rect 3496 4856 3528 4888
rect 3568 4856 3600 4888
rect 3640 4856 3672 4888
rect 3712 4856 3744 4888
rect 3784 4856 3816 4888
rect 3856 4856 3888 4888
rect 3928 4856 3960 4888
rect 40 4784 72 4816
rect 112 4784 144 4816
rect 184 4784 216 4816
rect 256 4784 288 4816
rect 328 4784 360 4816
rect 400 4784 432 4816
rect 472 4784 504 4816
rect 544 4784 576 4816
rect 616 4784 648 4816
rect 688 4784 720 4816
rect 760 4784 792 4816
rect 832 4784 864 4816
rect 904 4784 936 4816
rect 976 4784 1008 4816
rect 1048 4784 1080 4816
rect 1120 4784 1152 4816
rect 1192 4784 1224 4816
rect 1264 4784 1296 4816
rect 1336 4784 1368 4816
rect 1408 4784 1440 4816
rect 1480 4784 1512 4816
rect 1552 4784 1584 4816
rect 1624 4784 1656 4816
rect 1696 4784 1728 4816
rect 1768 4784 1800 4816
rect 1840 4784 1872 4816
rect 1912 4784 1944 4816
rect 1984 4784 2016 4816
rect 2056 4784 2088 4816
rect 2128 4784 2160 4816
rect 2200 4784 2232 4816
rect 2272 4784 2304 4816
rect 2344 4784 2376 4816
rect 2416 4784 2448 4816
rect 2488 4784 2520 4816
rect 2560 4784 2592 4816
rect 2632 4784 2664 4816
rect 2704 4784 2736 4816
rect 2776 4784 2808 4816
rect 2848 4784 2880 4816
rect 2920 4784 2952 4816
rect 2992 4784 3024 4816
rect 3064 4784 3096 4816
rect 3136 4784 3168 4816
rect 3208 4784 3240 4816
rect 3280 4784 3312 4816
rect 3352 4784 3384 4816
rect 3424 4784 3456 4816
rect 3496 4784 3528 4816
rect 3568 4784 3600 4816
rect 3640 4784 3672 4816
rect 3712 4784 3744 4816
rect 3784 4784 3816 4816
rect 3856 4784 3888 4816
rect 3928 4784 3960 4816
rect 40 4712 72 4744
rect 112 4712 144 4744
rect 184 4712 216 4744
rect 256 4712 288 4744
rect 328 4712 360 4744
rect 400 4712 432 4744
rect 472 4712 504 4744
rect 544 4712 576 4744
rect 616 4712 648 4744
rect 688 4712 720 4744
rect 760 4712 792 4744
rect 832 4712 864 4744
rect 904 4712 936 4744
rect 976 4712 1008 4744
rect 1048 4712 1080 4744
rect 1120 4712 1152 4744
rect 1192 4712 1224 4744
rect 1264 4712 1296 4744
rect 1336 4712 1368 4744
rect 1408 4712 1440 4744
rect 1480 4712 1512 4744
rect 1552 4712 1584 4744
rect 1624 4712 1656 4744
rect 1696 4712 1728 4744
rect 1768 4712 1800 4744
rect 1840 4712 1872 4744
rect 1912 4712 1944 4744
rect 1984 4712 2016 4744
rect 2056 4712 2088 4744
rect 2128 4712 2160 4744
rect 2200 4712 2232 4744
rect 2272 4712 2304 4744
rect 2344 4712 2376 4744
rect 2416 4712 2448 4744
rect 2488 4712 2520 4744
rect 2560 4712 2592 4744
rect 2632 4712 2664 4744
rect 2704 4712 2736 4744
rect 2776 4712 2808 4744
rect 2848 4712 2880 4744
rect 2920 4712 2952 4744
rect 2992 4712 3024 4744
rect 3064 4712 3096 4744
rect 3136 4712 3168 4744
rect 3208 4712 3240 4744
rect 3280 4712 3312 4744
rect 3352 4712 3384 4744
rect 3424 4712 3456 4744
rect 3496 4712 3528 4744
rect 3568 4712 3600 4744
rect 3640 4712 3672 4744
rect 3712 4712 3744 4744
rect 3784 4712 3816 4744
rect 3856 4712 3888 4744
rect 3928 4712 3960 4744
rect 40 4640 72 4672
rect 112 4640 144 4672
rect 184 4640 216 4672
rect 256 4640 288 4672
rect 328 4640 360 4672
rect 400 4640 432 4672
rect 472 4640 504 4672
rect 544 4640 576 4672
rect 616 4640 648 4672
rect 688 4640 720 4672
rect 760 4640 792 4672
rect 832 4640 864 4672
rect 904 4640 936 4672
rect 976 4640 1008 4672
rect 1048 4640 1080 4672
rect 1120 4640 1152 4672
rect 1192 4640 1224 4672
rect 1264 4640 1296 4672
rect 1336 4640 1368 4672
rect 1408 4640 1440 4672
rect 1480 4640 1512 4672
rect 1552 4640 1584 4672
rect 1624 4640 1656 4672
rect 1696 4640 1728 4672
rect 1768 4640 1800 4672
rect 1840 4640 1872 4672
rect 1912 4640 1944 4672
rect 1984 4640 2016 4672
rect 2056 4640 2088 4672
rect 2128 4640 2160 4672
rect 2200 4640 2232 4672
rect 2272 4640 2304 4672
rect 2344 4640 2376 4672
rect 2416 4640 2448 4672
rect 2488 4640 2520 4672
rect 2560 4640 2592 4672
rect 2632 4640 2664 4672
rect 2704 4640 2736 4672
rect 2776 4640 2808 4672
rect 2848 4640 2880 4672
rect 2920 4640 2952 4672
rect 2992 4640 3024 4672
rect 3064 4640 3096 4672
rect 3136 4640 3168 4672
rect 3208 4640 3240 4672
rect 3280 4640 3312 4672
rect 3352 4640 3384 4672
rect 3424 4640 3456 4672
rect 3496 4640 3528 4672
rect 3568 4640 3600 4672
rect 3640 4640 3672 4672
rect 3712 4640 3744 4672
rect 3784 4640 3816 4672
rect 3856 4640 3888 4672
rect 3928 4640 3960 4672
rect 40 4568 72 4600
rect 112 4568 144 4600
rect 184 4568 216 4600
rect 256 4568 288 4600
rect 328 4568 360 4600
rect 400 4568 432 4600
rect 472 4568 504 4600
rect 544 4568 576 4600
rect 616 4568 648 4600
rect 688 4568 720 4600
rect 760 4568 792 4600
rect 832 4568 864 4600
rect 904 4568 936 4600
rect 976 4568 1008 4600
rect 1048 4568 1080 4600
rect 1120 4568 1152 4600
rect 1192 4568 1224 4600
rect 1264 4568 1296 4600
rect 1336 4568 1368 4600
rect 1408 4568 1440 4600
rect 1480 4568 1512 4600
rect 1552 4568 1584 4600
rect 1624 4568 1656 4600
rect 1696 4568 1728 4600
rect 1768 4568 1800 4600
rect 1840 4568 1872 4600
rect 1912 4568 1944 4600
rect 1984 4568 2016 4600
rect 2056 4568 2088 4600
rect 2128 4568 2160 4600
rect 2200 4568 2232 4600
rect 2272 4568 2304 4600
rect 2344 4568 2376 4600
rect 2416 4568 2448 4600
rect 2488 4568 2520 4600
rect 2560 4568 2592 4600
rect 2632 4568 2664 4600
rect 2704 4568 2736 4600
rect 2776 4568 2808 4600
rect 2848 4568 2880 4600
rect 2920 4568 2952 4600
rect 2992 4568 3024 4600
rect 3064 4568 3096 4600
rect 3136 4568 3168 4600
rect 3208 4568 3240 4600
rect 3280 4568 3312 4600
rect 3352 4568 3384 4600
rect 3424 4568 3456 4600
rect 3496 4568 3528 4600
rect 3568 4568 3600 4600
rect 3640 4568 3672 4600
rect 3712 4568 3744 4600
rect 3784 4568 3816 4600
rect 3856 4568 3888 4600
rect 3928 4568 3960 4600
rect 40 4496 72 4528
rect 112 4496 144 4528
rect 184 4496 216 4528
rect 256 4496 288 4528
rect 328 4496 360 4528
rect 400 4496 432 4528
rect 472 4496 504 4528
rect 544 4496 576 4528
rect 616 4496 648 4528
rect 688 4496 720 4528
rect 760 4496 792 4528
rect 832 4496 864 4528
rect 904 4496 936 4528
rect 976 4496 1008 4528
rect 1048 4496 1080 4528
rect 1120 4496 1152 4528
rect 1192 4496 1224 4528
rect 1264 4496 1296 4528
rect 1336 4496 1368 4528
rect 1408 4496 1440 4528
rect 1480 4496 1512 4528
rect 1552 4496 1584 4528
rect 1624 4496 1656 4528
rect 1696 4496 1728 4528
rect 1768 4496 1800 4528
rect 1840 4496 1872 4528
rect 1912 4496 1944 4528
rect 1984 4496 2016 4528
rect 2056 4496 2088 4528
rect 2128 4496 2160 4528
rect 2200 4496 2232 4528
rect 2272 4496 2304 4528
rect 2344 4496 2376 4528
rect 2416 4496 2448 4528
rect 2488 4496 2520 4528
rect 2560 4496 2592 4528
rect 2632 4496 2664 4528
rect 2704 4496 2736 4528
rect 2776 4496 2808 4528
rect 2848 4496 2880 4528
rect 2920 4496 2952 4528
rect 2992 4496 3024 4528
rect 3064 4496 3096 4528
rect 3136 4496 3168 4528
rect 3208 4496 3240 4528
rect 3280 4496 3312 4528
rect 3352 4496 3384 4528
rect 3424 4496 3456 4528
rect 3496 4496 3528 4528
rect 3568 4496 3600 4528
rect 3640 4496 3672 4528
rect 3712 4496 3744 4528
rect 3784 4496 3816 4528
rect 3856 4496 3888 4528
rect 3928 4496 3960 4528
rect 40 4424 72 4456
rect 112 4424 144 4456
rect 184 4424 216 4456
rect 256 4424 288 4456
rect 328 4424 360 4456
rect 400 4424 432 4456
rect 472 4424 504 4456
rect 544 4424 576 4456
rect 616 4424 648 4456
rect 688 4424 720 4456
rect 760 4424 792 4456
rect 832 4424 864 4456
rect 904 4424 936 4456
rect 976 4424 1008 4456
rect 1048 4424 1080 4456
rect 1120 4424 1152 4456
rect 1192 4424 1224 4456
rect 1264 4424 1296 4456
rect 1336 4424 1368 4456
rect 1408 4424 1440 4456
rect 1480 4424 1512 4456
rect 1552 4424 1584 4456
rect 1624 4424 1656 4456
rect 1696 4424 1728 4456
rect 1768 4424 1800 4456
rect 1840 4424 1872 4456
rect 1912 4424 1944 4456
rect 1984 4424 2016 4456
rect 2056 4424 2088 4456
rect 2128 4424 2160 4456
rect 2200 4424 2232 4456
rect 2272 4424 2304 4456
rect 2344 4424 2376 4456
rect 2416 4424 2448 4456
rect 2488 4424 2520 4456
rect 2560 4424 2592 4456
rect 2632 4424 2664 4456
rect 2704 4424 2736 4456
rect 2776 4424 2808 4456
rect 2848 4424 2880 4456
rect 2920 4424 2952 4456
rect 2992 4424 3024 4456
rect 3064 4424 3096 4456
rect 3136 4424 3168 4456
rect 3208 4424 3240 4456
rect 3280 4424 3312 4456
rect 3352 4424 3384 4456
rect 3424 4424 3456 4456
rect 3496 4424 3528 4456
rect 3568 4424 3600 4456
rect 3640 4424 3672 4456
rect 3712 4424 3744 4456
rect 3784 4424 3816 4456
rect 3856 4424 3888 4456
rect 3928 4424 3960 4456
rect 40 4352 72 4384
rect 112 4352 144 4384
rect 184 4352 216 4384
rect 256 4352 288 4384
rect 328 4352 360 4384
rect 400 4352 432 4384
rect 472 4352 504 4384
rect 544 4352 576 4384
rect 616 4352 648 4384
rect 688 4352 720 4384
rect 760 4352 792 4384
rect 832 4352 864 4384
rect 904 4352 936 4384
rect 976 4352 1008 4384
rect 1048 4352 1080 4384
rect 1120 4352 1152 4384
rect 1192 4352 1224 4384
rect 1264 4352 1296 4384
rect 1336 4352 1368 4384
rect 1408 4352 1440 4384
rect 1480 4352 1512 4384
rect 1552 4352 1584 4384
rect 1624 4352 1656 4384
rect 1696 4352 1728 4384
rect 1768 4352 1800 4384
rect 1840 4352 1872 4384
rect 1912 4352 1944 4384
rect 1984 4352 2016 4384
rect 2056 4352 2088 4384
rect 2128 4352 2160 4384
rect 2200 4352 2232 4384
rect 2272 4352 2304 4384
rect 2344 4352 2376 4384
rect 2416 4352 2448 4384
rect 2488 4352 2520 4384
rect 2560 4352 2592 4384
rect 2632 4352 2664 4384
rect 2704 4352 2736 4384
rect 2776 4352 2808 4384
rect 2848 4352 2880 4384
rect 2920 4352 2952 4384
rect 2992 4352 3024 4384
rect 3064 4352 3096 4384
rect 3136 4352 3168 4384
rect 3208 4352 3240 4384
rect 3280 4352 3312 4384
rect 3352 4352 3384 4384
rect 3424 4352 3456 4384
rect 3496 4352 3528 4384
rect 3568 4352 3600 4384
rect 3640 4352 3672 4384
rect 3712 4352 3744 4384
rect 3784 4352 3816 4384
rect 3856 4352 3888 4384
rect 3928 4352 3960 4384
rect 40 4280 72 4312
rect 112 4280 144 4312
rect 184 4280 216 4312
rect 256 4280 288 4312
rect 328 4280 360 4312
rect 400 4280 432 4312
rect 472 4280 504 4312
rect 544 4280 576 4312
rect 616 4280 648 4312
rect 688 4280 720 4312
rect 760 4280 792 4312
rect 832 4280 864 4312
rect 904 4280 936 4312
rect 976 4280 1008 4312
rect 1048 4280 1080 4312
rect 1120 4280 1152 4312
rect 1192 4280 1224 4312
rect 1264 4280 1296 4312
rect 1336 4280 1368 4312
rect 1408 4280 1440 4312
rect 1480 4280 1512 4312
rect 1552 4280 1584 4312
rect 1624 4280 1656 4312
rect 1696 4280 1728 4312
rect 1768 4280 1800 4312
rect 1840 4280 1872 4312
rect 1912 4280 1944 4312
rect 1984 4280 2016 4312
rect 2056 4280 2088 4312
rect 2128 4280 2160 4312
rect 2200 4280 2232 4312
rect 2272 4280 2304 4312
rect 2344 4280 2376 4312
rect 2416 4280 2448 4312
rect 2488 4280 2520 4312
rect 2560 4280 2592 4312
rect 2632 4280 2664 4312
rect 2704 4280 2736 4312
rect 2776 4280 2808 4312
rect 2848 4280 2880 4312
rect 2920 4280 2952 4312
rect 2992 4280 3024 4312
rect 3064 4280 3096 4312
rect 3136 4280 3168 4312
rect 3208 4280 3240 4312
rect 3280 4280 3312 4312
rect 3352 4280 3384 4312
rect 3424 4280 3456 4312
rect 3496 4280 3528 4312
rect 3568 4280 3600 4312
rect 3640 4280 3672 4312
rect 3712 4280 3744 4312
rect 3784 4280 3816 4312
rect 3856 4280 3888 4312
rect 3928 4280 3960 4312
rect 40 4208 72 4240
rect 112 4208 144 4240
rect 184 4208 216 4240
rect 256 4208 288 4240
rect 328 4208 360 4240
rect 400 4208 432 4240
rect 472 4208 504 4240
rect 544 4208 576 4240
rect 616 4208 648 4240
rect 688 4208 720 4240
rect 760 4208 792 4240
rect 832 4208 864 4240
rect 904 4208 936 4240
rect 976 4208 1008 4240
rect 1048 4208 1080 4240
rect 1120 4208 1152 4240
rect 1192 4208 1224 4240
rect 1264 4208 1296 4240
rect 1336 4208 1368 4240
rect 1408 4208 1440 4240
rect 1480 4208 1512 4240
rect 1552 4208 1584 4240
rect 1624 4208 1656 4240
rect 1696 4208 1728 4240
rect 1768 4208 1800 4240
rect 1840 4208 1872 4240
rect 1912 4208 1944 4240
rect 1984 4208 2016 4240
rect 2056 4208 2088 4240
rect 2128 4208 2160 4240
rect 2200 4208 2232 4240
rect 2272 4208 2304 4240
rect 2344 4208 2376 4240
rect 2416 4208 2448 4240
rect 2488 4208 2520 4240
rect 2560 4208 2592 4240
rect 2632 4208 2664 4240
rect 2704 4208 2736 4240
rect 2776 4208 2808 4240
rect 2848 4208 2880 4240
rect 2920 4208 2952 4240
rect 2992 4208 3024 4240
rect 3064 4208 3096 4240
rect 3136 4208 3168 4240
rect 3208 4208 3240 4240
rect 3280 4208 3312 4240
rect 3352 4208 3384 4240
rect 3424 4208 3456 4240
rect 3496 4208 3528 4240
rect 3568 4208 3600 4240
rect 3640 4208 3672 4240
rect 3712 4208 3744 4240
rect 3784 4208 3816 4240
rect 3856 4208 3888 4240
rect 3928 4208 3960 4240
rect 40 4136 72 4168
rect 112 4136 144 4168
rect 184 4136 216 4168
rect 256 4136 288 4168
rect 328 4136 360 4168
rect 400 4136 432 4168
rect 472 4136 504 4168
rect 544 4136 576 4168
rect 616 4136 648 4168
rect 688 4136 720 4168
rect 760 4136 792 4168
rect 832 4136 864 4168
rect 904 4136 936 4168
rect 976 4136 1008 4168
rect 1048 4136 1080 4168
rect 1120 4136 1152 4168
rect 1192 4136 1224 4168
rect 1264 4136 1296 4168
rect 1336 4136 1368 4168
rect 1408 4136 1440 4168
rect 1480 4136 1512 4168
rect 1552 4136 1584 4168
rect 1624 4136 1656 4168
rect 1696 4136 1728 4168
rect 1768 4136 1800 4168
rect 1840 4136 1872 4168
rect 1912 4136 1944 4168
rect 1984 4136 2016 4168
rect 2056 4136 2088 4168
rect 2128 4136 2160 4168
rect 2200 4136 2232 4168
rect 2272 4136 2304 4168
rect 2344 4136 2376 4168
rect 2416 4136 2448 4168
rect 2488 4136 2520 4168
rect 2560 4136 2592 4168
rect 2632 4136 2664 4168
rect 2704 4136 2736 4168
rect 2776 4136 2808 4168
rect 2848 4136 2880 4168
rect 2920 4136 2952 4168
rect 2992 4136 3024 4168
rect 3064 4136 3096 4168
rect 3136 4136 3168 4168
rect 3208 4136 3240 4168
rect 3280 4136 3312 4168
rect 3352 4136 3384 4168
rect 3424 4136 3456 4168
rect 3496 4136 3528 4168
rect 3568 4136 3600 4168
rect 3640 4136 3672 4168
rect 3712 4136 3744 4168
rect 3784 4136 3816 4168
rect 3856 4136 3888 4168
rect 3928 4136 3960 4168
rect 40 4064 72 4096
rect 112 4064 144 4096
rect 184 4064 216 4096
rect 256 4064 288 4096
rect 328 4064 360 4096
rect 400 4064 432 4096
rect 472 4064 504 4096
rect 544 4064 576 4096
rect 616 4064 648 4096
rect 688 4064 720 4096
rect 760 4064 792 4096
rect 832 4064 864 4096
rect 904 4064 936 4096
rect 976 4064 1008 4096
rect 1048 4064 1080 4096
rect 1120 4064 1152 4096
rect 1192 4064 1224 4096
rect 1264 4064 1296 4096
rect 1336 4064 1368 4096
rect 1408 4064 1440 4096
rect 1480 4064 1512 4096
rect 1552 4064 1584 4096
rect 1624 4064 1656 4096
rect 1696 4064 1728 4096
rect 1768 4064 1800 4096
rect 1840 4064 1872 4096
rect 1912 4064 1944 4096
rect 1984 4064 2016 4096
rect 2056 4064 2088 4096
rect 2128 4064 2160 4096
rect 2200 4064 2232 4096
rect 2272 4064 2304 4096
rect 2344 4064 2376 4096
rect 2416 4064 2448 4096
rect 2488 4064 2520 4096
rect 2560 4064 2592 4096
rect 2632 4064 2664 4096
rect 2704 4064 2736 4096
rect 2776 4064 2808 4096
rect 2848 4064 2880 4096
rect 2920 4064 2952 4096
rect 2992 4064 3024 4096
rect 3064 4064 3096 4096
rect 3136 4064 3168 4096
rect 3208 4064 3240 4096
rect 3280 4064 3312 4096
rect 3352 4064 3384 4096
rect 3424 4064 3456 4096
rect 3496 4064 3528 4096
rect 3568 4064 3600 4096
rect 3640 4064 3672 4096
rect 3712 4064 3744 4096
rect 3784 4064 3816 4096
rect 3856 4064 3888 4096
rect 3928 4064 3960 4096
rect 40 3992 72 4024
rect 112 3992 144 4024
rect 184 3992 216 4024
rect 256 3992 288 4024
rect 328 3992 360 4024
rect 400 3992 432 4024
rect 472 3992 504 4024
rect 544 3992 576 4024
rect 616 3992 648 4024
rect 688 3992 720 4024
rect 760 3992 792 4024
rect 832 3992 864 4024
rect 904 3992 936 4024
rect 976 3992 1008 4024
rect 1048 3992 1080 4024
rect 1120 3992 1152 4024
rect 1192 3992 1224 4024
rect 1264 3992 1296 4024
rect 1336 3992 1368 4024
rect 1408 3992 1440 4024
rect 1480 3992 1512 4024
rect 1552 3992 1584 4024
rect 1624 3992 1656 4024
rect 1696 3992 1728 4024
rect 1768 3992 1800 4024
rect 1840 3992 1872 4024
rect 1912 3992 1944 4024
rect 1984 3992 2016 4024
rect 2056 3992 2088 4024
rect 2128 3992 2160 4024
rect 2200 3992 2232 4024
rect 2272 3992 2304 4024
rect 2344 3992 2376 4024
rect 2416 3992 2448 4024
rect 2488 3992 2520 4024
rect 2560 3992 2592 4024
rect 2632 3992 2664 4024
rect 2704 3992 2736 4024
rect 2776 3992 2808 4024
rect 2848 3992 2880 4024
rect 2920 3992 2952 4024
rect 2992 3992 3024 4024
rect 3064 3992 3096 4024
rect 3136 3992 3168 4024
rect 3208 3992 3240 4024
rect 3280 3992 3312 4024
rect 3352 3992 3384 4024
rect 3424 3992 3456 4024
rect 3496 3992 3528 4024
rect 3568 3992 3600 4024
rect 3640 3992 3672 4024
rect 3712 3992 3744 4024
rect 3784 3992 3816 4024
rect 3856 3992 3888 4024
rect 3928 3992 3960 4024
rect 40 3920 72 3952
rect 112 3920 144 3952
rect 184 3920 216 3952
rect 256 3920 288 3952
rect 328 3920 360 3952
rect 400 3920 432 3952
rect 472 3920 504 3952
rect 544 3920 576 3952
rect 616 3920 648 3952
rect 688 3920 720 3952
rect 760 3920 792 3952
rect 832 3920 864 3952
rect 904 3920 936 3952
rect 976 3920 1008 3952
rect 1048 3920 1080 3952
rect 1120 3920 1152 3952
rect 1192 3920 1224 3952
rect 1264 3920 1296 3952
rect 1336 3920 1368 3952
rect 1408 3920 1440 3952
rect 1480 3920 1512 3952
rect 1552 3920 1584 3952
rect 1624 3920 1656 3952
rect 1696 3920 1728 3952
rect 1768 3920 1800 3952
rect 1840 3920 1872 3952
rect 1912 3920 1944 3952
rect 1984 3920 2016 3952
rect 2056 3920 2088 3952
rect 2128 3920 2160 3952
rect 2200 3920 2232 3952
rect 2272 3920 2304 3952
rect 2344 3920 2376 3952
rect 2416 3920 2448 3952
rect 2488 3920 2520 3952
rect 2560 3920 2592 3952
rect 2632 3920 2664 3952
rect 2704 3920 2736 3952
rect 2776 3920 2808 3952
rect 2848 3920 2880 3952
rect 2920 3920 2952 3952
rect 2992 3920 3024 3952
rect 3064 3920 3096 3952
rect 3136 3920 3168 3952
rect 3208 3920 3240 3952
rect 3280 3920 3312 3952
rect 3352 3920 3384 3952
rect 3424 3920 3456 3952
rect 3496 3920 3528 3952
rect 3568 3920 3600 3952
rect 3640 3920 3672 3952
rect 3712 3920 3744 3952
rect 3784 3920 3816 3952
rect 3856 3920 3888 3952
rect 3928 3920 3960 3952
rect 40 3848 72 3880
rect 112 3848 144 3880
rect 184 3848 216 3880
rect 256 3848 288 3880
rect 328 3848 360 3880
rect 400 3848 432 3880
rect 472 3848 504 3880
rect 544 3848 576 3880
rect 616 3848 648 3880
rect 688 3848 720 3880
rect 760 3848 792 3880
rect 832 3848 864 3880
rect 904 3848 936 3880
rect 976 3848 1008 3880
rect 1048 3848 1080 3880
rect 1120 3848 1152 3880
rect 1192 3848 1224 3880
rect 1264 3848 1296 3880
rect 1336 3848 1368 3880
rect 1408 3848 1440 3880
rect 1480 3848 1512 3880
rect 1552 3848 1584 3880
rect 1624 3848 1656 3880
rect 1696 3848 1728 3880
rect 1768 3848 1800 3880
rect 1840 3848 1872 3880
rect 1912 3848 1944 3880
rect 1984 3848 2016 3880
rect 2056 3848 2088 3880
rect 2128 3848 2160 3880
rect 2200 3848 2232 3880
rect 2272 3848 2304 3880
rect 2344 3848 2376 3880
rect 2416 3848 2448 3880
rect 2488 3848 2520 3880
rect 2560 3848 2592 3880
rect 2632 3848 2664 3880
rect 2704 3848 2736 3880
rect 2776 3848 2808 3880
rect 2848 3848 2880 3880
rect 2920 3848 2952 3880
rect 2992 3848 3024 3880
rect 3064 3848 3096 3880
rect 3136 3848 3168 3880
rect 3208 3848 3240 3880
rect 3280 3848 3312 3880
rect 3352 3848 3384 3880
rect 3424 3848 3456 3880
rect 3496 3848 3528 3880
rect 3568 3848 3600 3880
rect 3640 3848 3672 3880
rect 3712 3848 3744 3880
rect 3784 3848 3816 3880
rect 3856 3848 3888 3880
rect 3928 3848 3960 3880
rect 40 3776 72 3808
rect 112 3776 144 3808
rect 184 3776 216 3808
rect 256 3776 288 3808
rect 328 3776 360 3808
rect 400 3776 432 3808
rect 472 3776 504 3808
rect 544 3776 576 3808
rect 616 3776 648 3808
rect 688 3776 720 3808
rect 760 3776 792 3808
rect 832 3776 864 3808
rect 904 3776 936 3808
rect 976 3776 1008 3808
rect 1048 3776 1080 3808
rect 1120 3776 1152 3808
rect 1192 3776 1224 3808
rect 1264 3776 1296 3808
rect 1336 3776 1368 3808
rect 1408 3776 1440 3808
rect 1480 3776 1512 3808
rect 1552 3776 1584 3808
rect 1624 3776 1656 3808
rect 1696 3776 1728 3808
rect 1768 3776 1800 3808
rect 1840 3776 1872 3808
rect 1912 3776 1944 3808
rect 1984 3776 2016 3808
rect 2056 3776 2088 3808
rect 2128 3776 2160 3808
rect 2200 3776 2232 3808
rect 2272 3776 2304 3808
rect 2344 3776 2376 3808
rect 2416 3776 2448 3808
rect 2488 3776 2520 3808
rect 2560 3776 2592 3808
rect 2632 3776 2664 3808
rect 2704 3776 2736 3808
rect 2776 3776 2808 3808
rect 2848 3776 2880 3808
rect 2920 3776 2952 3808
rect 2992 3776 3024 3808
rect 3064 3776 3096 3808
rect 3136 3776 3168 3808
rect 3208 3776 3240 3808
rect 3280 3776 3312 3808
rect 3352 3776 3384 3808
rect 3424 3776 3456 3808
rect 3496 3776 3528 3808
rect 3568 3776 3600 3808
rect 3640 3776 3672 3808
rect 3712 3776 3744 3808
rect 3784 3776 3816 3808
rect 3856 3776 3888 3808
rect 3928 3776 3960 3808
rect 40 3704 72 3736
rect 112 3704 144 3736
rect 184 3704 216 3736
rect 256 3704 288 3736
rect 328 3704 360 3736
rect 400 3704 432 3736
rect 472 3704 504 3736
rect 544 3704 576 3736
rect 616 3704 648 3736
rect 688 3704 720 3736
rect 760 3704 792 3736
rect 832 3704 864 3736
rect 904 3704 936 3736
rect 976 3704 1008 3736
rect 1048 3704 1080 3736
rect 1120 3704 1152 3736
rect 1192 3704 1224 3736
rect 1264 3704 1296 3736
rect 1336 3704 1368 3736
rect 1408 3704 1440 3736
rect 1480 3704 1512 3736
rect 1552 3704 1584 3736
rect 1624 3704 1656 3736
rect 1696 3704 1728 3736
rect 1768 3704 1800 3736
rect 1840 3704 1872 3736
rect 1912 3704 1944 3736
rect 1984 3704 2016 3736
rect 2056 3704 2088 3736
rect 2128 3704 2160 3736
rect 2200 3704 2232 3736
rect 2272 3704 2304 3736
rect 2344 3704 2376 3736
rect 2416 3704 2448 3736
rect 2488 3704 2520 3736
rect 2560 3704 2592 3736
rect 2632 3704 2664 3736
rect 2704 3704 2736 3736
rect 2776 3704 2808 3736
rect 2848 3704 2880 3736
rect 2920 3704 2952 3736
rect 2992 3704 3024 3736
rect 3064 3704 3096 3736
rect 3136 3704 3168 3736
rect 3208 3704 3240 3736
rect 3280 3704 3312 3736
rect 3352 3704 3384 3736
rect 3424 3704 3456 3736
rect 3496 3704 3528 3736
rect 3568 3704 3600 3736
rect 3640 3704 3672 3736
rect 3712 3704 3744 3736
rect 3784 3704 3816 3736
rect 3856 3704 3888 3736
rect 3928 3704 3960 3736
rect 40 3632 72 3664
rect 112 3632 144 3664
rect 184 3632 216 3664
rect 256 3632 288 3664
rect 328 3632 360 3664
rect 400 3632 432 3664
rect 472 3632 504 3664
rect 544 3632 576 3664
rect 616 3632 648 3664
rect 688 3632 720 3664
rect 760 3632 792 3664
rect 832 3632 864 3664
rect 904 3632 936 3664
rect 976 3632 1008 3664
rect 1048 3632 1080 3664
rect 1120 3632 1152 3664
rect 1192 3632 1224 3664
rect 1264 3632 1296 3664
rect 1336 3632 1368 3664
rect 1408 3632 1440 3664
rect 1480 3632 1512 3664
rect 1552 3632 1584 3664
rect 1624 3632 1656 3664
rect 1696 3632 1728 3664
rect 1768 3632 1800 3664
rect 1840 3632 1872 3664
rect 1912 3632 1944 3664
rect 1984 3632 2016 3664
rect 2056 3632 2088 3664
rect 2128 3632 2160 3664
rect 2200 3632 2232 3664
rect 2272 3632 2304 3664
rect 2344 3632 2376 3664
rect 2416 3632 2448 3664
rect 2488 3632 2520 3664
rect 2560 3632 2592 3664
rect 2632 3632 2664 3664
rect 2704 3632 2736 3664
rect 2776 3632 2808 3664
rect 2848 3632 2880 3664
rect 2920 3632 2952 3664
rect 2992 3632 3024 3664
rect 3064 3632 3096 3664
rect 3136 3632 3168 3664
rect 3208 3632 3240 3664
rect 3280 3632 3312 3664
rect 3352 3632 3384 3664
rect 3424 3632 3456 3664
rect 3496 3632 3528 3664
rect 3568 3632 3600 3664
rect 3640 3632 3672 3664
rect 3712 3632 3744 3664
rect 3784 3632 3816 3664
rect 3856 3632 3888 3664
rect 3928 3632 3960 3664
rect 40 3560 72 3592
rect 112 3560 144 3592
rect 184 3560 216 3592
rect 256 3560 288 3592
rect 328 3560 360 3592
rect 400 3560 432 3592
rect 472 3560 504 3592
rect 544 3560 576 3592
rect 616 3560 648 3592
rect 688 3560 720 3592
rect 760 3560 792 3592
rect 832 3560 864 3592
rect 904 3560 936 3592
rect 976 3560 1008 3592
rect 1048 3560 1080 3592
rect 1120 3560 1152 3592
rect 1192 3560 1224 3592
rect 1264 3560 1296 3592
rect 1336 3560 1368 3592
rect 1408 3560 1440 3592
rect 1480 3560 1512 3592
rect 1552 3560 1584 3592
rect 1624 3560 1656 3592
rect 1696 3560 1728 3592
rect 1768 3560 1800 3592
rect 1840 3560 1872 3592
rect 1912 3560 1944 3592
rect 1984 3560 2016 3592
rect 2056 3560 2088 3592
rect 2128 3560 2160 3592
rect 2200 3560 2232 3592
rect 2272 3560 2304 3592
rect 2344 3560 2376 3592
rect 2416 3560 2448 3592
rect 2488 3560 2520 3592
rect 2560 3560 2592 3592
rect 2632 3560 2664 3592
rect 2704 3560 2736 3592
rect 2776 3560 2808 3592
rect 2848 3560 2880 3592
rect 2920 3560 2952 3592
rect 2992 3560 3024 3592
rect 3064 3560 3096 3592
rect 3136 3560 3168 3592
rect 3208 3560 3240 3592
rect 3280 3560 3312 3592
rect 3352 3560 3384 3592
rect 3424 3560 3456 3592
rect 3496 3560 3528 3592
rect 3568 3560 3600 3592
rect 3640 3560 3672 3592
rect 3712 3560 3744 3592
rect 3784 3560 3816 3592
rect 3856 3560 3888 3592
rect 3928 3560 3960 3592
rect 40 3488 72 3520
rect 112 3488 144 3520
rect 184 3488 216 3520
rect 256 3488 288 3520
rect 328 3488 360 3520
rect 400 3488 432 3520
rect 472 3488 504 3520
rect 544 3488 576 3520
rect 616 3488 648 3520
rect 688 3488 720 3520
rect 760 3488 792 3520
rect 832 3488 864 3520
rect 904 3488 936 3520
rect 976 3488 1008 3520
rect 1048 3488 1080 3520
rect 1120 3488 1152 3520
rect 1192 3488 1224 3520
rect 1264 3488 1296 3520
rect 1336 3488 1368 3520
rect 1408 3488 1440 3520
rect 1480 3488 1512 3520
rect 1552 3488 1584 3520
rect 1624 3488 1656 3520
rect 1696 3488 1728 3520
rect 1768 3488 1800 3520
rect 1840 3488 1872 3520
rect 1912 3488 1944 3520
rect 1984 3488 2016 3520
rect 2056 3488 2088 3520
rect 2128 3488 2160 3520
rect 2200 3488 2232 3520
rect 2272 3488 2304 3520
rect 2344 3488 2376 3520
rect 2416 3488 2448 3520
rect 2488 3488 2520 3520
rect 2560 3488 2592 3520
rect 2632 3488 2664 3520
rect 2704 3488 2736 3520
rect 2776 3488 2808 3520
rect 2848 3488 2880 3520
rect 2920 3488 2952 3520
rect 2992 3488 3024 3520
rect 3064 3488 3096 3520
rect 3136 3488 3168 3520
rect 3208 3488 3240 3520
rect 3280 3488 3312 3520
rect 3352 3488 3384 3520
rect 3424 3488 3456 3520
rect 3496 3488 3528 3520
rect 3568 3488 3600 3520
rect 3640 3488 3672 3520
rect 3712 3488 3744 3520
rect 3784 3488 3816 3520
rect 3856 3488 3888 3520
rect 3928 3488 3960 3520
rect 40 3416 72 3448
rect 112 3416 144 3448
rect 184 3416 216 3448
rect 256 3416 288 3448
rect 328 3416 360 3448
rect 400 3416 432 3448
rect 472 3416 504 3448
rect 544 3416 576 3448
rect 616 3416 648 3448
rect 688 3416 720 3448
rect 760 3416 792 3448
rect 832 3416 864 3448
rect 904 3416 936 3448
rect 976 3416 1008 3448
rect 1048 3416 1080 3448
rect 1120 3416 1152 3448
rect 1192 3416 1224 3448
rect 1264 3416 1296 3448
rect 1336 3416 1368 3448
rect 1408 3416 1440 3448
rect 1480 3416 1512 3448
rect 1552 3416 1584 3448
rect 1624 3416 1656 3448
rect 1696 3416 1728 3448
rect 1768 3416 1800 3448
rect 1840 3416 1872 3448
rect 1912 3416 1944 3448
rect 1984 3416 2016 3448
rect 2056 3416 2088 3448
rect 2128 3416 2160 3448
rect 2200 3416 2232 3448
rect 2272 3416 2304 3448
rect 2344 3416 2376 3448
rect 2416 3416 2448 3448
rect 2488 3416 2520 3448
rect 2560 3416 2592 3448
rect 2632 3416 2664 3448
rect 2704 3416 2736 3448
rect 2776 3416 2808 3448
rect 2848 3416 2880 3448
rect 2920 3416 2952 3448
rect 2992 3416 3024 3448
rect 3064 3416 3096 3448
rect 3136 3416 3168 3448
rect 3208 3416 3240 3448
rect 3280 3416 3312 3448
rect 3352 3416 3384 3448
rect 3424 3416 3456 3448
rect 3496 3416 3528 3448
rect 3568 3416 3600 3448
rect 3640 3416 3672 3448
rect 3712 3416 3744 3448
rect 3784 3416 3816 3448
rect 3856 3416 3888 3448
rect 3928 3416 3960 3448
rect 40 3344 72 3376
rect 112 3344 144 3376
rect 184 3344 216 3376
rect 256 3344 288 3376
rect 328 3344 360 3376
rect 400 3344 432 3376
rect 472 3344 504 3376
rect 544 3344 576 3376
rect 616 3344 648 3376
rect 688 3344 720 3376
rect 760 3344 792 3376
rect 832 3344 864 3376
rect 904 3344 936 3376
rect 976 3344 1008 3376
rect 1048 3344 1080 3376
rect 1120 3344 1152 3376
rect 1192 3344 1224 3376
rect 1264 3344 1296 3376
rect 1336 3344 1368 3376
rect 1408 3344 1440 3376
rect 1480 3344 1512 3376
rect 1552 3344 1584 3376
rect 1624 3344 1656 3376
rect 1696 3344 1728 3376
rect 1768 3344 1800 3376
rect 1840 3344 1872 3376
rect 1912 3344 1944 3376
rect 1984 3344 2016 3376
rect 2056 3344 2088 3376
rect 2128 3344 2160 3376
rect 2200 3344 2232 3376
rect 2272 3344 2304 3376
rect 2344 3344 2376 3376
rect 2416 3344 2448 3376
rect 2488 3344 2520 3376
rect 2560 3344 2592 3376
rect 2632 3344 2664 3376
rect 2704 3344 2736 3376
rect 2776 3344 2808 3376
rect 2848 3344 2880 3376
rect 2920 3344 2952 3376
rect 2992 3344 3024 3376
rect 3064 3344 3096 3376
rect 3136 3344 3168 3376
rect 3208 3344 3240 3376
rect 3280 3344 3312 3376
rect 3352 3344 3384 3376
rect 3424 3344 3456 3376
rect 3496 3344 3528 3376
rect 3568 3344 3600 3376
rect 3640 3344 3672 3376
rect 3712 3344 3744 3376
rect 3784 3344 3816 3376
rect 3856 3344 3888 3376
rect 3928 3344 3960 3376
rect 40 3272 72 3304
rect 112 3272 144 3304
rect 184 3272 216 3304
rect 256 3272 288 3304
rect 328 3272 360 3304
rect 400 3272 432 3304
rect 472 3272 504 3304
rect 544 3272 576 3304
rect 616 3272 648 3304
rect 688 3272 720 3304
rect 760 3272 792 3304
rect 832 3272 864 3304
rect 904 3272 936 3304
rect 976 3272 1008 3304
rect 1048 3272 1080 3304
rect 1120 3272 1152 3304
rect 1192 3272 1224 3304
rect 1264 3272 1296 3304
rect 1336 3272 1368 3304
rect 1408 3272 1440 3304
rect 1480 3272 1512 3304
rect 1552 3272 1584 3304
rect 1624 3272 1656 3304
rect 1696 3272 1728 3304
rect 1768 3272 1800 3304
rect 1840 3272 1872 3304
rect 1912 3272 1944 3304
rect 1984 3272 2016 3304
rect 2056 3272 2088 3304
rect 2128 3272 2160 3304
rect 2200 3272 2232 3304
rect 2272 3272 2304 3304
rect 2344 3272 2376 3304
rect 2416 3272 2448 3304
rect 2488 3272 2520 3304
rect 2560 3272 2592 3304
rect 2632 3272 2664 3304
rect 2704 3272 2736 3304
rect 2776 3272 2808 3304
rect 2848 3272 2880 3304
rect 2920 3272 2952 3304
rect 2992 3272 3024 3304
rect 3064 3272 3096 3304
rect 3136 3272 3168 3304
rect 3208 3272 3240 3304
rect 3280 3272 3312 3304
rect 3352 3272 3384 3304
rect 3424 3272 3456 3304
rect 3496 3272 3528 3304
rect 3568 3272 3600 3304
rect 3640 3272 3672 3304
rect 3712 3272 3744 3304
rect 3784 3272 3816 3304
rect 3856 3272 3888 3304
rect 3928 3272 3960 3304
rect 40 3200 72 3232
rect 112 3200 144 3232
rect 184 3200 216 3232
rect 256 3200 288 3232
rect 328 3200 360 3232
rect 400 3200 432 3232
rect 472 3200 504 3232
rect 544 3200 576 3232
rect 616 3200 648 3232
rect 688 3200 720 3232
rect 760 3200 792 3232
rect 832 3200 864 3232
rect 904 3200 936 3232
rect 976 3200 1008 3232
rect 1048 3200 1080 3232
rect 1120 3200 1152 3232
rect 1192 3200 1224 3232
rect 1264 3200 1296 3232
rect 1336 3200 1368 3232
rect 1408 3200 1440 3232
rect 1480 3200 1512 3232
rect 1552 3200 1584 3232
rect 1624 3200 1656 3232
rect 1696 3200 1728 3232
rect 1768 3200 1800 3232
rect 1840 3200 1872 3232
rect 1912 3200 1944 3232
rect 1984 3200 2016 3232
rect 2056 3200 2088 3232
rect 2128 3200 2160 3232
rect 2200 3200 2232 3232
rect 2272 3200 2304 3232
rect 2344 3200 2376 3232
rect 2416 3200 2448 3232
rect 2488 3200 2520 3232
rect 2560 3200 2592 3232
rect 2632 3200 2664 3232
rect 2704 3200 2736 3232
rect 2776 3200 2808 3232
rect 2848 3200 2880 3232
rect 2920 3200 2952 3232
rect 2992 3200 3024 3232
rect 3064 3200 3096 3232
rect 3136 3200 3168 3232
rect 3208 3200 3240 3232
rect 3280 3200 3312 3232
rect 3352 3200 3384 3232
rect 3424 3200 3456 3232
rect 3496 3200 3528 3232
rect 3568 3200 3600 3232
rect 3640 3200 3672 3232
rect 3712 3200 3744 3232
rect 3784 3200 3816 3232
rect 3856 3200 3888 3232
rect 3928 3200 3960 3232
rect 40 3128 72 3160
rect 112 3128 144 3160
rect 184 3128 216 3160
rect 256 3128 288 3160
rect 328 3128 360 3160
rect 400 3128 432 3160
rect 472 3128 504 3160
rect 544 3128 576 3160
rect 616 3128 648 3160
rect 688 3128 720 3160
rect 760 3128 792 3160
rect 832 3128 864 3160
rect 904 3128 936 3160
rect 976 3128 1008 3160
rect 1048 3128 1080 3160
rect 1120 3128 1152 3160
rect 1192 3128 1224 3160
rect 1264 3128 1296 3160
rect 1336 3128 1368 3160
rect 1408 3128 1440 3160
rect 1480 3128 1512 3160
rect 1552 3128 1584 3160
rect 1624 3128 1656 3160
rect 1696 3128 1728 3160
rect 1768 3128 1800 3160
rect 1840 3128 1872 3160
rect 1912 3128 1944 3160
rect 1984 3128 2016 3160
rect 2056 3128 2088 3160
rect 2128 3128 2160 3160
rect 2200 3128 2232 3160
rect 2272 3128 2304 3160
rect 2344 3128 2376 3160
rect 2416 3128 2448 3160
rect 2488 3128 2520 3160
rect 2560 3128 2592 3160
rect 2632 3128 2664 3160
rect 2704 3128 2736 3160
rect 2776 3128 2808 3160
rect 2848 3128 2880 3160
rect 2920 3128 2952 3160
rect 2992 3128 3024 3160
rect 3064 3128 3096 3160
rect 3136 3128 3168 3160
rect 3208 3128 3240 3160
rect 3280 3128 3312 3160
rect 3352 3128 3384 3160
rect 3424 3128 3456 3160
rect 3496 3128 3528 3160
rect 3568 3128 3600 3160
rect 3640 3128 3672 3160
rect 3712 3128 3744 3160
rect 3784 3128 3816 3160
rect 3856 3128 3888 3160
rect 3928 3128 3960 3160
rect 40 3056 72 3088
rect 112 3056 144 3088
rect 184 3056 216 3088
rect 256 3056 288 3088
rect 328 3056 360 3088
rect 400 3056 432 3088
rect 472 3056 504 3088
rect 544 3056 576 3088
rect 616 3056 648 3088
rect 688 3056 720 3088
rect 760 3056 792 3088
rect 832 3056 864 3088
rect 904 3056 936 3088
rect 976 3056 1008 3088
rect 1048 3056 1080 3088
rect 1120 3056 1152 3088
rect 1192 3056 1224 3088
rect 1264 3056 1296 3088
rect 1336 3056 1368 3088
rect 1408 3056 1440 3088
rect 1480 3056 1512 3088
rect 1552 3056 1584 3088
rect 1624 3056 1656 3088
rect 1696 3056 1728 3088
rect 1768 3056 1800 3088
rect 1840 3056 1872 3088
rect 1912 3056 1944 3088
rect 1984 3056 2016 3088
rect 2056 3056 2088 3088
rect 2128 3056 2160 3088
rect 2200 3056 2232 3088
rect 2272 3056 2304 3088
rect 2344 3056 2376 3088
rect 2416 3056 2448 3088
rect 2488 3056 2520 3088
rect 2560 3056 2592 3088
rect 2632 3056 2664 3088
rect 2704 3056 2736 3088
rect 2776 3056 2808 3088
rect 2848 3056 2880 3088
rect 2920 3056 2952 3088
rect 2992 3056 3024 3088
rect 3064 3056 3096 3088
rect 3136 3056 3168 3088
rect 3208 3056 3240 3088
rect 3280 3056 3312 3088
rect 3352 3056 3384 3088
rect 3424 3056 3456 3088
rect 3496 3056 3528 3088
rect 3568 3056 3600 3088
rect 3640 3056 3672 3088
rect 3712 3056 3744 3088
rect 3784 3056 3816 3088
rect 3856 3056 3888 3088
rect 3928 3056 3960 3088
rect 40 2984 72 3016
rect 112 2984 144 3016
rect 184 2984 216 3016
rect 256 2984 288 3016
rect 328 2984 360 3016
rect 400 2984 432 3016
rect 472 2984 504 3016
rect 544 2984 576 3016
rect 616 2984 648 3016
rect 688 2984 720 3016
rect 760 2984 792 3016
rect 832 2984 864 3016
rect 904 2984 936 3016
rect 976 2984 1008 3016
rect 1048 2984 1080 3016
rect 1120 2984 1152 3016
rect 1192 2984 1224 3016
rect 1264 2984 1296 3016
rect 1336 2984 1368 3016
rect 1408 2984 1440 3016
rect 1480 2984 1512 3016
rect 1552 2984 1584 3016
rect 1624 2984 1656 3016
rect 1696 2984 1728 3016
rect 1768 2984 1800 3016
rect 1840 2984 1872 3016
rect 1912 2984 1944 3016
rect 1984 2984 2016 3016
rect 2056 2984 2088 3016
rect 2128 2984 2160 3016
rect 2200 2984 2232 3016
rect 2272 2984 2304 3016
rect 2344 2984 2376 3016
rect 2416 2984 2448 3016
rect 2488 2984 2520 3016
rect 2560 2984 2592 3016
rect 2632 2984 2664 3016
rect 2704 2984 2736 3016
rect 2776 2984 2808 3016
rect 2848 2984 2880 3016
rect 2920 2984 2952 3016
rect 2992 2984 3024 3016
rect 3064 2984 3096 3016
rect 3136 2984 3168 3016
rect 3208 2984 3240 3016
rect 3280 2984 3312 3016
rect 3352 2984 3384 3016
rect 3424 2984 3456 3016
rect 3496 2984 3528 3016
rect 3568 2984 3600 3016
rect 3640 2984 3672 3016
rect 3712 2984 3744 3016
rect 3784 2984 3816 3016
rect 3856 2984 3888 3016
rect 3928 2984 3960 3016
rect 40 2912 72 2944
rect 112 2912 144 2944
rect 184 2912 216 2944
rect 256 2912 288 2944
rect 328 2912 360 2944
rect 400 2912 432 2944
rect 472 2912 504 2944
rect 544 2912 576 2944
rect 616 2912 648 2944
rect 688 2912 720 2944
rect 760 2912 792 2944
rect 832 2912 864 2944
rect 904 2912 936 2944
rect 976 2912 1008 2944
rect 1048 2912 1080 2944
rect 1120 2912 1152 2944
rect 1192 2912 1224 2944
rect 1264 2912 1296 2944
rect 1336 2912 1368 2944
rect 1408 2912 1440 2944
rect 1480 2912 1512 2944
rect 1552 2912 1584 2944
rect 1624 2912 1656 2944
rect 1696 2912 1728 2944
rect 1768 2912 1800 2944
rect 1840 2912 1872 2944
rect 1912 2912 1944 2944
rect 1984 2912 2016 2944
rect 2056 2912 2088 2944
rect 2128 2912 2160 2944
rect 2200 2912 2232 2944
rect 2272 2912 2304 2944
rect 2344 2912 2376 2944
rect 2416 2912 2448 2944
rect 2488 2912 2520 2944
rect 2560 2912 2592 2944
rect 2632 2912 2664 2944
rect 2704 2912 2736 2944
rect 2776 2912 2808 2944
rect 2848 2912 2880 2944
rect 2920 2912 2952 2944
rect 2992 2912 3024 2944
rect 3064 2912 3096 2944
rect 3136 2912 3168 2944
rect 3208 2912 3240 2944
rect 3280 2912 3312 2944
rect 3352 2912 3384 2944
rect 3424 2912 3456 2944
rect 3496 2912 3528 2944
rect 3568 2912 3600 2944
rect 3640 2912 3672 2944
rect 3712 2912 3744 2944
rect 3784 2912 3816 2944
rect 3856 2912 3888 2944
rect 3928 2912 3960 2944
rect 40 2840 72 2872
rect 112 2840 144 2872
rect 184 2840 216 2872
rect 256 2840 288 2872
rect 328 2840 360 2872
rect 400 2840 432 2872
rect 472 2840 504 2872
rect 544 2840 576 2872
rect 616 2840 648 2872
rect 688 2840 720 2872
rect 760 2840 792 2872
rect 832 2840 864 2872
rect 904 2840 936 2872
rect 976 2840 1008 2872
rect 1048 2840 1080 2872
rect 1120 2840 1152 2872
rect 1192 2840 1224 2872
rect 1264 2840 1296 2872
rect 1336 2840 1368 2872
rect 1408 2840 1440 2872
rect 1480 2840 1512 2872
rect 1552 2840 1584 2872
rect 1624 2840 1656 2872
rect 1696 2840 1728 2872
rect 1768 2840 1800 2872
rect 1840 2840 1872 2872
rect 1912 2840 1944 2872
rect 1984 2840 2016 2872
rect 2056 2840 2088 2872
rect 2128 2840 2160 2872
rect 2200 2840 2232 2872
rect 2272 2840 2304 2872
rect 2344 2840 2376 2872
rect 2416 2840 2448 2872
rect 2488 2840 2520 2872
rect 2560 2840 2592 2872
rect 2632 2840 2664 2872
rect 2704 2840 2736 2872
rect 2776 2840 2808 2872
rect 2848 2840 2880 2872
rect 2920 2840 2952 2872
rect 2992 2840 3024 2872
rect 3064 2840 3096 2872
rect 3136 2840 3168 2872
rect 3208 2840 3240 2872
rect 3280 2840 3312 2872
rect 3352 2840 3384 2872
rect 3424 2840 3456 2872
rect 3496 2840 3528 2872
rect 3568 2840 3600 2872
rect 3640 2840 3672 2872
rect 3712 2840 3744 2872
rect 3784 2840 3816 2872
rect 3856 2840 3888 2872
rect 3928 2840 3960 2872
rect 40 2768 72 2800
rect 112 2768 144 2800
rect 184 2768 216 2800
rect 256 2768 288 2800
rect 328 2768 360 2800
rect 400 2768 432 2800
rect 472 2768 504 2800
rect 544 2768 576 2800
rect 616 2768 648 2800
rect 688 2768 720 2800
rect 760 2768 792 2800
rect 832 2768 864 2800
rect 904 2768 936 2800
rect 976 2768 1008 2800
rect 1048 2768 1080 2800
rect 1120 2768 1152 2800
rect 1192 2768 1224 2800
rect 1264 2768 1296 2800
rect 1336 2768 1368 2800
rect 1408 2768 1440 2800
rect 1480 2768 1512 2800
rect 1552 2768 1584 2800
rect 1624 2768 1656 2800
rect 1696 2768 1728 2800
rect 1768 2768 1800 2800
rect 1840 2768 1872 2800
rect 1912 2768 1944 2800
rect 1984 2768 2016 2800
rect 2056 2768 2088 2800
rect 2128 2768 2160 2800
rect 2200 2768 2232 2800
rect 2272 2768 2304 2800
rect 2344 2768 2376 2800
rect 2416 2768 2448 2800
rect 2488 2768 2520 2800
rect 2560 2768 2592 2800
rect 2632 2768 2664 2800
rect 2704 2768 2736 2800
rect 2776 2768 2808 2800
rect 2848 2768 2880 2800
rect 2920 2768 2952 2800
rect 2992 2768 3024 2800
rect 3064 2768 3096 2800
rect 3136 2768 3168 2800
rect 3208 2768 3240 2800
rect 3280 2768 3312 2800
rect 3352 2768 3384 2800
rect 3424 2768 3456 2800
rect 3496 2768 3528 2800
rect 3568 2768 3600 2800
rect 3640 2768 3672 2800
rect 3712 2768 3744 2800
rect 3784 2768 3816 2800
rect 3856 2768 3888 2800
rect 3928 2768 3960 2800
rect 40 2696 72 2728
rect 112 2696 144 2728
rect 184 2696 216 2728
rect 256 2696 288 2728
rect 328 2696 360 2728
rect 400 2696 432 2728
rect 472 2696 504 2728
rect 544 2696 576 2728
rect 616 2696 648 2728
rect 688 2696 720 2728
rect 760 2696 792 2728
rect 832 2696 864 2728
rect 904 2696 936 2728
rect 976 2696 1008 2728
rect 1048 2696 1080 2728
rect 1120 2696 1152 2728
rect 1192 2696 1224 2728
rect 1264 2696 1296 2728
rect 1336 2696 1368 2728
rect 1408 2696 1440 2728
rect 1480 2696 1512 2728
rect 1552 2696 1584 2728
rect 1624 2696 1656 2728
rect 1696 2696 1728 2728
rect 1768 2696 1800 2728
rect 1840 2696 1872 2728
rect 1912 2696 1944 2728
rect 1984 2696 2016 2728
rect 2056 2696 2088 2728
rect 2128 2696 2160 2728
rect 2200 2696 2232 2728
rect 2272 2696 2304 2728
rect 2344 2696 2376 2728
rect 2416 2696 2448 2728
rect 2488 2696 2520 2728
rect 2560 2696 2592 2728
rect 2632 2696 2664 2728
rect 2704 2696 2736 2728
rect 2776 2696 2808 2728
rect 2848 2696 2880 2728
rect 2920 2696 2952 2728
rect 2992 2696 3024 2728
rect 3064 2696 3096 2728
rect 3136 2696 3168 2728
rect 3208 2696 3240 2728
rect 3280 2696 3312 2728
rect 3352 2696 3384 2728
rect 3424 2696 3456 2728
rect 3496 2696 3528 2728
rect 3568 2696 3600 2728
rect 3640 2696 3672 2728
rect 3712 2696 3744 2728
rect 3784 2696 3816 2728
rect 3856 2696 3888 2728
rect 3928 2696 3960 2728
rect 40 2624 72 2656
rect 112 2624 144 2656
rect 184 2624 216 2656
rect 256 2624 288 2656
rect 328 2624 360 2656
rect 400 2624 432 2656
rect 472 2624 504 2656
rect 544 2624 576 2656
rect 616 2624 648 2656
rect 688 2624 720 2656
rect 760 2624 792 2656
rect 832 2624 864 2656
rect 904 2624 936 2656
rect 976 2624 1008 2656
rect 1048 2624 1080 2656
rect 1120 2624 1152 2656
rect 1192 2624 1224 2656
rect 1264 2624 1296 2656
rect 1336 2624 1368 2656
rect 1408 2624 1440 2656
rect 1480 2624 1512 2656
rect 1552 2624 1584 2656
rect 1624 2624 1656 2656
rect 1696 2624 1728 2656
rect 1768 2624 1800 2656
rect 1840 2624 1872 2656
rect 1912 2624 1944 2656
rect 1984 2624 2016 2656
rect 2056 2624 2088 2656
rect 2128 2624 2160 2656
rect 2200 2624 2232 2656
rect 2272 2624 2304 2656
rect 2344 2624 2376 2656
rect 2416 2624 2448 2656
rect 2488 2624 2520 2656
rect 2560 2624 2592 2656
rect 2632 2624 2664 2656
rect 2704 2624 2736 2656
rect 2776 2624 2808 2656
rect 2848 2624 2880 2656
rect 2920 2624 2952 2656
rect 2992 2624 3024 2656
rect 3064 2624 3096 2656
rect 3136 2624 3168 2656
rect 3208 2624 3240 2656
rect 3280 2624 3312 2656
rect 3352 2624 3384 2656
rect 3424 2624 3456 2656
rect 3496 2624 3528 2656
rect 3568 2624 3600 2656
rect 3640 2624 3672 2656
rect 3712 2624 3744 2656
rect 3784 2624 3816 2656
rect 3856 2624 3888 2656
rect 3928 2624 3960 2656
rect 40 2552 72 2584
rect 112 2552 144 2584
rect 184 2552 216 2584
rect 256 2552 288 2584
rect 328 2552 360 2584
rect 400 2552 432 2584
rect 472 2552 504 2584
rect 544 2552 576 2584
rect 616 2552 648 2584
rect 688 2552 720 2584
rect 760 2552 792 2584
rect 832 2552 864 2584
rect 904 2552 936 2584
rect 976 2552 1008 2584
rect 1048 2552 1080 2584
rect 1120 2552 1152 2584
rect 1192 2552 1224 2584
rect 1264 2552 1296 2584
rect 1336 2552 1368 2584
rect 1408 2552 1440 2584
rect 1480 2552 1512 2584
rect 1552 2552 1584 2584
rect 1624 2552 1656 2584
rect 1696 2552 1728 2584
rect 1768 2552 1800 2584
rect 1840 2552 1872 2584
rect 1912 2552 1944 2584
rect 1984 2552 2016 2584
rect 2056 2552 2088 2584
rect 2128 2552 2160 2584
rect 2200 2552 2232 2584
rect 2272 2552 2304 2584
rect 2344 2552 2376 2584
rect 2416 2552 2448 2584
rect 2488 2552 2520 2584
rect 2560 2552 2592 2584
rect 2632 2552 2664 2584
rect 2704 2552 2736 2584
rect 2776 2552 2808 2584
rect 2848 2552 2880 2584
rect 2920 2552 2952 2584
rect 2992 2552 3024 2584
rect 3064 2552 3096 2584
rect 3136 2552 3168 2584
rect 3208 2552 3240 2584
rect 3280 2552 3312 2584
rect 3352 2552 3384 2584
rect 3424 2552 3456 2584
rect 3496 2552 3528 2584
rect 3568 2552 3600 2584
rect 3640 2552 3672 2584
rect 3712 2552 3744 2584
rect 3784 2552 3816 2584
rect 3856 2552 3888 2584
rect 3928 2552 3960 2584
rect 40 2480 72 2512
rect 112 2480 144 2512
rect 184 2480 216 2512
rect 256 2480 288 2512
rect 328 2480 360 2512
rect 400 2480 432 2512
rect 472 2480 504 2512
rect 544 2480 576 2512
rect 616 2480 648 2512
rect 688 2480 720 2512
rect 760 2480 792 2512
rect 832 2480 864 2512
rect 904 2480 936 2512
rect 976 2480 1008 2512
rect 1048 2480 1080 2512
rect 1120 2480 1152 2512
rect 1192 2480 1224 2512
rect 1264 2480 1296 2512
rect 1336 2480 1368 2512
rect 1408 2480 1440 2512
rect 1480 2480 1512 2512
rect 1552 2480 1584 2512
rect 1624 2480 1656 2512
rect 1696 2480 1728 2512
rect 1768 2480 1800 2512
rect 1840 2480 1872 2512
rect 1912 2480 1944 2512
rect 1984 2480 2016 2512
rect 2056 2480 2088 2512
rect 2128 2480 2160 2512
rect 2200 2480 2232 2512
rect 2272 2480 2304 2512
rect 2344 2480 2376 2512
rect 2416 2480 2448 2512
rect 2488 2480 2520 2512
rect 2560 2480 2592 2512
rect 2632 2480 2664 2512
rect 2704 2480 2736 2512
rect 2776 2480 2808 2512
rect 2848 2480 2880 2512
rect 2920 2480 2952 2512
rect 2992 2480 3024 2512
rect 3064 2480 3096 2512
rect 3136 2480 3168 2512
rect 3208 2480 3240 2512
rect 3280 2480 3312 2512
rect 3352 2480 3384 2512
rect 3424 2480 3456 2512
rect 3496 2480 3528 2512
rect 3568 2480 3600 2512
rect 3640 2480 3672 2512
rect 3712 2480 3744 2512
rect 3784 2480 3816 2512
rect 3856 2480 3888 2512
rect 3928 2480 3960 2512
rect 40 2408 72 2440
rect 112 2408 144 2440
rect 184 2408 216 2440
rect 256 2408 288 2440
rect 328 2408 360 2440
rect 400 2408 432 2440
rect 472 2408 504 2440
rect 544 2408 576 2440
rect 616 2408 648 2440
rect 688 2408 720 2440
rect 760 2408 792 2440
rect 832 2408 864 2440
rect 904 2408 936 2440
rect 976 2408 1008 2440
rect 1048 2408 1080 2440
rect 1120 2408 1152 2440
rect 1192 2408 1224 2440
rect 1264 2408 1296 2440
rect 1336 2408 1368 2440
rect 1408 2408 1440 2440
rect 1480 2408 1512 2440
rect 1552 2408 1584 2440
rect 1624 2408 1656 2440
rect 1696 2408 1728 2440
rect 1768 2408 1800 2440
rect 1840 2408 1872 2440
rect 1912 2408 1944 2440
rect 1984 2408 2016 2440
rect 2056 2408 2088 2440
rect 2128 2408 2160 2440
rect 2200 2408 2232 2440
rect 2272 2408 2304 2440
rect 2344 2408 2376 2440
rect 2416 2408 2448 2440
rect 2488 2408 2520 2440
rect 2560 2408 2592 2440
rect 2632 2408 2664 2440
rect 2704 2408 2736 2440
rect 2776 2408 2808 2440
rect 2848 2408 2880 2440
rect 2920 2408 2952 2440
rect 2992 2408 3024 2440
rect 3064 2408 3096 2440
rect 3136 2408 3168 2440
rect 3208 2408 3240 2440
rect 3280 2408 3312 2440
rect 3352 2408 3384 2440
rect 3424 2408 3456 2440
rect 3496 2408 3528 2440
rect 3568 2408 3600 2440
rect 3640 2408 3672 2440
rect 3712 2408 3744 2440
rect 3784 2408 3816 2440
rect 3856 2408 3888 2440
rect 3928 2408 3960 2440
rect 40 2336 72 2368
rect 112 2336 144 2368
rect 184 2336 216 2368
rect 256 2336 288 2368
rect 328 2336 360 2368
rect 400 2336 432 2368
rect 472 2336 504 2368
rect 544 2336 576 2368
rect 616 2336 648 2368
rect 688 2336 720 2368
rect 760 2336 792 2368
rect 832 2336 864 2368
rect 904 2336 936 2368
rect 976 2336 1008 2368
rect 1048 2336 1080 2368
rect 1120 2336 1152 2368
rect 1192 2336 1224 2368
rect 1264 2336 1296 2368
rect 1336 2336 1368 2368
rect 1408 2336 1440 2368
rect 1480 2336 1512 2368
rect 1552 2336 1584 2368
rect 1624 2336 1656 2368
rect 1696 2336 1728 2368
rect 1768 2336 1800 2368
rect 1840 2336 1872 2368
rect 1912 2336 1944 2368
rect 1984 2336 2016 2368
rect 2056 2336 2088 2368
rect 2128 2336 2160 2368
rect 2200 2336 2232 2368
rect 2272 2336 2304 2368
rect 2344 2336 2376 2368
rect 2416 2336 2448 2368
rect 2488 2336 2520 2368
rect 2560 2336 2592 2368
rect 2632 2336 2664 2368
rect 2704 2336 2736 2368
rect 2776 2336 2808 2368
rect 2848 2336 2880 2368
rect 2920 2336 2952 2368
rect 2992 2336 3024 2368
rect 3064 2336 3096 2368
rect 3136 2336 3168 2368
rect 3208 2336 3240 2368
rect 3280 2336 3312 2368
rect 3352 2336 3384 2368
rect 3424 2336 3456 2368
rect 3496 2336 3528 2368
rect 3568 2336 3600 2368
rect 3640 2336 3672 2368
rect 3712 2336 3744 2368
rect 3784 2336 3816 2368
rect 3856 2336 3888 2368
rect 3928 2336 3960 2368
rect 40 2264 72 2296
rect 112 2264 144 2296
rect 184 2264 216 2296
rect 256 2264 288 2296
rect 328 2264 360 2296
rect 400 2264 432 2296
rect 472 2264 504 2296
rect 544 2264 576 2296
rect 616 2264 648 2296
rect 688 2264 720 2296
rect 760 2264 792 2296
rect 832 2264 864 2296
rect 904 2264 936 2296
rect 976 2264 1008 2296
rect 1048 2264 1080 2296
rect 1120 2264 1152 2296
rect 1192 2264 1224 2296
rect 1264 2264 1296 2296
rect 1336 2264 1368 2296
rect 1408 2264 1440 2296
rect 1480 2264 1512 2296
rect 1552 2264 1584 2296
rect 1624 2264 1656 2296
rect 1696 2264 1728 2296
rect 1768 2264 1800 2296
rect 1840 2264 1872 2296
rect 1912 2264 1944 2296
rect 1984 2264 2016 2296
rect 2056 2264 2088 2296
rect 2128 2264 2160 2296
rect 2200 2264 2232 2296
rect 2272 2264 2304 2296
rect 2344 2264 2376 2296
rect 2416 2264 2448 2296
rect 2488 2264 2520 2296
rect 2560 2264 2592 2296
rect 2632 2264 2664 2296
rect 2704 2264 2736 2296
rect 2776 2264 2808 2296
rect 2848 2264 2880 2296
rect 2920 2264 2952 2296
rect 2992 2264 3024 2296
rect 3064 2264 3096 2296
rect 3136 2264 3168 2296
rect 3208 2264 3240 2296
rect 3280 2264 3312 2296
rect 3352 2264 3384 2296
rect 3424 2264 3456 2296
rect 3496 2264 3528 2296
rect 3568 2264 3600 2296
rect 3640 2264 3672 2296
rect 3712 2264 3744 2296
rect 3784 2264 3816 2296
rect 3856 2264 3888 2296
rect 3928 2264 3960 2296
rect 40 2192 72 2224
rect 112 2192 144 2224
rect 184 2192 216 2224
rect 256 2192 288 2224
rect 328 2192 360 2224
rect 400 2192 432 2224
rect 472 2192 504 2224
rect 544 2192 576 2224
rect 616 2192 648 2224
rect 688 2192 720 2224
rect 760 2192 792 2224
rect 832 2192 864 2224
rect 904 2192 936 2224
rect 976 2192 1008 2224
rect 1048 2192 1080 2224
rect 1120 2192 1152 2224
rect 1192 2192 1224 2224
rect 1264 2192 1296 2224
rect 1336 2192 1368 2224
rect 1408 2192 1440 2224
rect 1480 2192 1512 2224
rect 1552 2192 1584 2224
rect 1624 2192 1656 2224
rect 1696 2192 1728 2224
rect 1768 2192 1800 2224
rect 1840 2192 1872 2224
rect 1912 2192 1944 2224
rect 1984 2192 2016 2224
rect 2056 2192 2088 2224
rect 2128 2192 2160 2224
rect 2200 2192 2232 2224
rect 2272 2192 2304 2224
rect 2344 2192 2376 2224
rect 2416 2192 2448 2224
rect 2488 2192 2520 2224
rect 2560 2192 2592 2224
rect 2632 2192 2664 2224
rect 2704 2192 2736 2224
rect 2776 2192 2808 2224
rect 2848 2192 2880 2224
rect 2920 2192 2952 2224
rect 2992 2192 3024 2224
rect 3064 2192 3096 2224
rect 3136 2192 3168 2224
rect 3208 2192 3240 2224
rect 3280 2192 3312 2224
rect 3352 2192 3384 2224
rect 3424 2192 3456 2224
rect 3496 2192 3528 2224
rect 3568 2192 3600 2224
rect 3640 2192 3672 2224
rect 3712 2192 3744 2224
rect 3784 2192 3816 2224
rect 3856 2192 3888 2224
rect 3928 2192 3960 2224
rect 40 2120 72 2152
rect 112 2120 144 2152
rect 184 2120 216 2152
rect 256 2120 288 2152
rect 328 2120 360 2152
rect 400 2120 432 2152
rect 472 2120 504 2152
rect 544 2120 576 2152
rect 616 2120 648 2152
rect 688 2120 720 2152
rect 760 2120 792 2152
rect 832 2120 864 2152
rect 904 2120 936 2152
rect 976 2120 1008 2152
rect 1048 2120 1080 2152
rect 1120 2120 1152 2152
rect 1192 2120 1224 2152
rect 1264 2120 1296 2152
rect 1336 2120 1368 2152
rect 1408 2120 1440 2152
rect 1480 2120 1512 2152
rect 1552 2120 1584 2152
rect 1624 2120 1656 2152
rect 1696 2120 1728 2152
rect 1768 2120 1800 2152
rect 1840 2120 1872 2152
rect 1912 2120 1944 2152
rect 1984 2120 2016 2152
rect 2056 2120 2088 2152
rect 2128 2120 2160 2152
rect 2200 2120 2232 2152
rect 2272 2120 2304 2152
rect 2344 2120 2376 2152
rect 2416 2120 2448 2152
rect 2488 2120 2520 2152
rect 2560 2120 2592 2152
rect 2632 2120 2664 2152
rect 2704 2120 2736 2152
rect 2776 2120 2808 2152
rect 2848 2120 2880 2152
rect 2920 2120 2952 2152
rect 2992 2120 3024 2152
rect 3064 2120 3096 2152
rect 3136 2120 3168 2152
rect 3208 2120 3240 2152
rect 3280 2120 3312 2152
rect 3352 2120 3384 2152
rect 3424 2120 3456 2152
rect 3496 2120 3528 2152
rect 3568 2120 3600 2152
rect 3640 2120 3672 2152
rect 3712 2120 3744 2152
rect 3784 2120 3816 2152
rect 3856 2120 3888 2152
rect 3928 2120 3960 2152
rect 40 2048 72 2080
rect 112 2048 144 2080
rect 184 2048 216 2080
rect 256 2048 288 2080
rect 328 2048 360 2080
rect 400 2048 432 2080
rect 472 2048 504 2080
rect 544 2048 576 2080
rect 616 2048 648 2080
rect 688 2048 720 2080
rect 760 2048 792 2080
rect 832 2048 864 2080
rect 904 2048 936 2080
rect 976 2048 1008 2080
rect 1048 2048 1080 2080
rect 1120 2048 1152 2080
rect 1192 2048 1224 2080
rect 1264 2048 1296 2080
rect 1336 2048 1368 2080
rect 1408 2048 1440 2080
rect 1480 2048 1512 2080
rect 1552 2048 1584 2080
rect 1624 2048 1656 2080
rect 1696 2048 1728 2080
rect 1768 2048 1800 2080
rect 1840 2048 1872 2080
rect 1912 2048 1944 2080
rect 1984 2048 2016 2080
rect 2056 2048 2088 2080
rect 2128 2048 2160 2080
rect 2200 2048 2232 2080
rect 2272 2048 2304 2080
rect 2344 2048 2376 2080
rect 2416 2048 2448 2080
rect 2488 2048 2520 2080
rect 2560 2048 2592 2080
rect 2632 2048 2664 2080
rect 2704 2048 2736 2080
rect 2776 2048 2808 2080
rect 2848 2048 2880 2080
rect 2920 2048 2952 2080
rect 2992 2048 3024 2080
rect 3064 2048 3096 2080
rect 3136 2048 3168 2080
rect 3208 2048 3240 2080
rect 3280 2048 3312 2080
rect 3352 2048 3384 2080
rect 3424 2048 3456 2080
rect 3496 2048 3528 2080
rect 3568 2048 3600 2080
rect 3640 2048 3672 2080
rect 3712 2048 3744 2080
rect 3784 2048 3816 2080
rect 3856 2048 3888 2080
rect 3928 2048 3960 2080
rect 40 1976 72 2008
rect 112 1976 144 2008
rect 184 1976 216 2008
rect 256 1976 288 2008
rect 328 1976 360 2008
rect 400 1976 432 2008
rect 472 1976 504 2008
rect 544 1976 576 2008
rect 616 1976 648 2008
rect 688 1976 720 2008
rect 760 1976 792 2008
rect 832 1976 864 2008
rect 904 1976 936 2008
rect 976 1976 1008 2008
rect 1048 1976 1080 2008
rect 1120 1976 1152 2008
rect 1192 1976 1224 2008
rect 1264 1976 1296 2008
rect 1336 1976 1368 2008
rect 1408 1976 1440 2008
rect 1480 1976 1512 2008
rect 1552 1976 1584 2008
rect 1624 1976 1656 2008
rect 1696 1976 1728 2008
rect 1768 1976 1800 2008
rect 1840 1976 1872 2008
rect 1912 1976 1944 2008
rect 1984 1976 2016 2008
rect 2056 1976 2088 2008
rect 2128 1976 2160 2008
rect 2200 1976 2232 2008
rect 2272 1976 2304 2008
rect 2344 1976 2376 2008
rect 2416 1976 2448 2008
rect 2488 1976 2520 2008
rect 2560 1976 2592 2008
rect 2632 1976 2664 2008
rect 2704 1976 2736 2008
rect 2776 1976 2808 2008
rect 2848 1976 2880 2008
rect 2920 1976 2952 2008
rect 2992 1976 3024 2008
rect 3064 1976 3096 2008
rect 3136 1976 3168 2008
rect 3208 1976 3240 2008
rect 3280 1976 3312 2008
rect 3352 1976 3384 2008
rect 3424 1976 3456 2008
rect 3496 1976 3528 2008
rect 3568 1976 3600 2008
rect 3640 1976 3672 2008
rect 3712 1976 3744 2008
rect 3784 1976 3816 2008
rect 3856 1976 3888 2008
rect 3928 1976 3960 2008
rect 40 1904 72 1936
rect 112 1904 144 1936
rect 184 1904 216 1936
rect 256 1904 288 1936
rect 328 1904 360 1936
rect 400 1904 432 1936
rect 472 1904 504 1936
rect 544 1904 576 1936
rect 616 1904 648 1936
rect 688 1904 720 1936
rect 760 1904 792 1936
rect 832 1904 864 1936
rect 904 1904 936 1936
rect 976 1904 1008 1936
rect 1048 1904 1080 1936
rect 1120 1904 1152 1936
rect 1192 1904 1224 1936
rect 1264 1904 1296 1936
rect 1336 1904 1368 1936
rect 1408 1904 1440 1936
rect 1480 1904 1512 1936
rect 1552 1904 1584 1936
rect 1624 1904 1656 1936
rect 1696 1904 1728 1936
rect 1768 1904 1800 1936
rect 1840 1904 1872 1936
rect 1912 1904 1944 1936
rect 1984 1904 2016 1936
rect 2056 1904 2088 1936
rect 2128 1904 2160 1936
rect 2200 1904 2232 1936
rect 2272 1904 2304 1936
rect 2344 1904 2376 1936
rect 2416 1904 2448 1936
rect 2488 1904 2520 1936
rect 2560 1904 2592 1936
rect 2632 1904 2664 1936
rect 2704 1904 2736 1936
rect 2776 1904 2808 1936
rect 2848 1904 2880 1936
rect 2920 1904 2952 1936
rect 2992 1904 3024 1936
rect 3064 1904 3096 1936
rect 3136 1904 3168 1936
rect 3208 1904 3240 1936
rect 3280 1904 3312 1936
rect 3352 1904 3384 1936
rect 3424 1904 3456 1936
rect 3496 1904 3528 1936
rect 3568 1904 3600 1936
rect 3640 1904 3672 1936
rect 3712 1904 3744 1936
rect 3784 1904 3816 1936
rect 3856 1904 3888 1936
rect 3928 1904 3960 1936
rect 40 1832 72 1864
rect 112 1832 144 1864
rect 184 1832 216 1864
rect 256 1832 288 1864
rect 328 1832 360 1864
rect 400 1832 432 1864
rect 472 1832 504 1864
rect 544 1832 576 1864
rect 616 1832 648 1864
rect 688 1832 720 1864
rect 760 1832 792 1864
rect 832 1832 864 1864
rect 904 1832 936 1864
rect 976 1832 1008 1864
rect 1048 1832 1080 1864
rect 1120 1832 1152 1864
rect 1192 1832 1224 1864
rect 1264 1832 1296 1864
rect 1336 1832 1368 1864
rect 1408 1832 1440 1864
rect 1480 1832 1512 1864
rect 1552 1832 1584 1864
rect 1624 1832 1656 1864
rect 1696 1832 1728 1864
rect 1768 1832 1800 1864
rect 1840 1832 1872 1864
rect 1912 1832 1944 1864
rect 1984 1832 2016 1864
rect 2056 1832 2088 1864
rect 2128 1832 2160 1864
rect 2200 1832 2232 1864
rect 2272 1832 2304 1864
rect 2344 1832 2376 1864
rect 2416 1832 2448 1864
rect 2488 1832 2520 1864
rect 2560 1832 2592 1864
rect 2632 1832 2664 1864
rect 2704 1832 2736 1864
rect 2776 1832 2808 1864
rect 2848 1832 2880 1864
rect 2920 1832 2952 1864
rect 2992 1832 3024 1864
rect 3064 1832 3096 1864
rect 3136 1832 3168 1864
rect 3208 1832 3240 1864
rect 3280 1832 3312 1864
rect 3352 1832 3384 1864
rect 3424 1832 3456 1864
rect 3496 1832 3528 1864
rect 3568 1832 3600 1864
rect 3640 1832 3672 1864
rect 3712 1832 3744 1864
rect 3784 1832 3816 1864
rect 3856 1832 3888 1864
rect 3928 1832 3960 1864
rect 40 1760 72 1792
rect 112 1760 144 1792
rect 184 1760 216 1792
rect 256 1760 288 1792
rect 328 1760 360 1792
rect 400 1760 432 1792
rect 472 1760 504 1792
rect 544 1760 576 1792
rect 616 1760 648 1792
rect 688 1760 720 1792
rect 760 1760 792 1792
rect 832 1760 864 1792
rect 904 1760 936 1792
rect 976 1760 1008 1792
rect 1048 1760 1080 1792
rect 1120 1760 1152 1792
rect 1192 1760 1224 1792
rect 1264 1760 1296 1792
rect 1336 1760 1368 1792
rect 1408 1760 1440 1792
rect 1480 1760 1512 1792
rect 1552 1760 1584 1792
rect 1624 1760 1656 1792
rect 1696 1760 1728 1792
rect 1768 1760 1800 1792
rect 1840 1760 1872 1792
rect 1912 1760 1944 1792
rect 1984 1760 2016 1792
rect 2056 1760 2088 1792
rect 2128 1760 2160 1792
rect 2200 1760 2232 1792
rect 2272 1760 2304 1792
rect 2344 1760 2376 1792
rect 2416 1760 2448 1792
rect 2488 1760 2520 1792
rect 2560 1760 2592 1792
rect 2632 1760 2664 1792
rect 2704 1760 2736 1792
rect 2776 1760 2808 1792
rect 2848 1760 2880 1792
rect 2920 1760 2952 1792
rect 2992 1760 3024 1792
rect 3064 1760 3096 1792
rect 3136 1760 3168 1792
rect 3208 1760 3240 1792
rect 3280 1760 3312 1792
rect 3352 1760 3384 1792
rect 3424 1760 3456 1792
rect 3496 1760 3528 1792
rect 3568 1760 3600 1792
rect 3640 1760 3672 1792
rect 3712 1760 3744 1792
rect 3784 1760 3816 1792
rect 3856 1760 3888 1792
rect 3928 1760 3960 1792
rect 40 1688 72 1720
rect 112 1688 144 1720
rect 184 1688 216 1720
rect 256 1688 288 1720
rect 328 1688 360 1720
rect 400 1688 432 1720
rect 472 1688 504 1720
rect 544 1688 576 1720
rect 616 1688 648 1720
rect 688 1688 720 1720
rect 760 1688 792 1720
rect 832 1688 864 1720
rect 904 1688 936 1720
rect 976 1688 1008 1720
rect 1048 1688 1080 1720
rect 1120 1688 1152 1720
rect 1192 1688 1224 1720
rect 1264 1688 1296 1720
rect 1336 1688 1368 1720
rect 1408 1688 1440 1720
rect 1480 1688 1512 1720
rect 1552 1688 1584 1720
rect 1624 1688 1656 1720
rect 1696 1688 1728 1720
rect 1768 1688 1800 1720
rect 1840 1688 1872 1720
rect 1912 1688 1944 1720
rect 1984 1688 2016 1720
rect 2056 1688 2088 1720
rect 2128 1688 2160 1720
rect 2200 1688 2232 1720
rect 2272 1688 2304 1720
rect 2344 1688 2376 1720
rect 2416 1688 2448 1720
rect 2488 1688 2520 1720
rect 2560 1688 2592 1720
rect 2632 1688 2664 1720
rect 2704 1688 2736 1720
rect 2776 1688 2808 1720
rect 2848 1688 2880 1720
rect 2920 1688 2952 1720
rect 2992 1688 3024 1720
rect 3064 1688 3096 1720
rect 3136 1688 3168 1720
rect 3208 1688 3240 1720
rect 3280 1688 3312 1720
rect 3352 1688 3384 1720
rect 3424 1688 3456 1720
rect 3496 1688 3528 1720
rect 3568 1688 3600 1720
rect 3640 1688 3672 1720
rect 3712 1688 3744 1720
rect 3784 1688 3816 1720
rect 3856 1688 3888 1720
rect 3928 1688 3960 1720
rect 40 1616 72 1648
rect 112 1616 144 1648
rect 184 1616 216 1648
rect 256 1616 288 1648
rect 328 1616 360 1648
rect 400 1616 432 1648
rect 472 1616 504 1648
rect 544 1616 576 1648
rect 616 1616 648 1648
rect 688 1616 720 1648
rect 760 1616 792 1648
rect 832 1616 864 1648
rect 904 1616 936 1648
rect 976 1616 1008 1648
rect 1048 1616 1080 1648
rect 1120 1616 1152 1648
rect 1192 1616 1224 1648
rect 1264 1616 1296 1648
rect 1336 1616 1368 1648
rect 1408 1616 1440 1648
rect 1480 1616 1512 1648
rect 1552 1616 1584 1648
rect 1624 1616 1656 1648
rect 1696 1616 1728 1648
rect 1768 1616 1800 1648
rect 1840 1616 1872 1648
rect 1912 1616 1944 1648
rect 1984 1616 2016 1648
rect 2056 1616 2088 1648
rect 2128 1616 2160 1648
rect 2200 1616 2232 1648
rect 2272 1616 2304 1648
rect 2344 1616 2376 1648
rect 2416 1616 2448 1648
rect 2488 1616 2520 1648
rect 2560 1616 2592 1648
rect 2632 1616 2664 1648
rect 2704 1616 2736 1648
rect 2776 1616 2808 1648
rect 2848 1616 2880 1648
rect 2920 1616 2952 1648
rect 2992 1616 3024 1648
rect 3064 1616 3096 1648
rect 3136 1616 3168 1648
rect 3208 1616 3240 1648
rect 3280 1616 3312 1648
rect 3352 1616 3384 1648
rect 3424 1616 3456 1648
rect 3496 1616 3528 1648
rect 3568 1616 3600 1648
rect 3640 1616 3672 1648
rect 3712 1616 3744 1648
rect 3784 1616 3816 1648
rect 3856 1616 3888 1648
rect 3928 1616 3960 1648
rect 40 1544 72 1576
rect 112 1544 144 1576
rect 184 1544 216 1576
rect 256 1544 288 1576
rect 328 1544 360 1576
rect 400 1544 432 1576
rect 472 1544 504 1576
rect 544 1544 576 1576
rect 616 1544 648 1576
rect 688 1544 720 1576
rect 760 1544 792 1576
rect 832 1544 864 1576
rect 904 1544 936 1576
rect 976 1544 1008 1576
rect 1048 1544 1080 1576
rect 1120 1544 1152 1576
rect 1192 1544 1224 1576
rect 1264 1544 1296 1576
rect 1336 1544 1368 1576
rect 1408 1544 1440 1576
rect 1480 1544 1512 1576
rect 1552 1544 1584 1576
rect 1624 1544 1656 1576
rect 1696 1544 1728 1576
rect 1768 1544 1800 1576
rect 1840 1544 1872 1576
rect 1912 1544 1944 1576
rect 1984 1544 2016 1576
rect 2056 1544 2088 1576
rect 2128 1544 2160 1576
rect 2200 1544 2232 1576
rect 2272 1544 2304 1576
rect 2344 1544 2376 1576
rect 2416 1544 2448 1576
rect 2488 1544 2520 1576
rect 2560 1544 2592 1576
rect 2632 1544 2664 1576
rect 2704 1544 2736 1576
rect 2776 1544 2808 1576
rect 2848 1544 2880 1576
rect 2920 1544 2952 1576
rect 2992 1544 3024 1576
rect 3064 1544 3096 1576
rect 3136 1544 3168 1576
rect 3208 1544 3240 1576
rect 3280 1544 3312 1576
rect 3352 1544 3384 1576
rect 3424 1544 3456 1576
rect 3496 1544 3528 1576
rect 3568 1544 3600 1576
rect 3640 1544 3672 1576
rect 3712 1544 3744 1576
rect 3784 1544 3816 1576
rect 3856 1544 3888 1576
rect 3928 1544 3960 1576
rect 40 1472 72 1504
rect 112 1472 144 1504
rect 184 1472 216 1504
rect 256 1472 288 1504
rect 328 1472 360 1504
rect 400 1472 432 1504
rect 472 1472 504 1504
rect 544 1472 576 1504
rect 616 1472 648 1504
rect 688 1472 720 1504
rect 760 1472 792 1504
rect 832 1472 864 1504
rect 904 1472 936 1504
rect 976 1472 1008 1504
rect 1048 1472 1080 1504
rect 1120 1472 1152 1504
rect 1192 1472 1224 1504
rect 1264 1472 1296 1504
rect 1336 1472 1368 1504
rect 1408 1472 1440 1504
rect 1480 1472 1512 1504
rect 1552 1472 1584 1504
rect 1624 1472 1656 1504
rect 1696 1472 1728 1504
rect 1768 1472 1800 1504
rect 1840 1472 1872 1504
rect 1912 1472 1944 1504
rect 1984 1472 2016 1504
rect 2056 1472 2088 1504
rect 2128 1472 2160 1504
rect 2200 1472 2232 1504
rect 2272 1472 2304 1504
rect 2344 1472 2376 1504
rect 2416 1472 2448 1504
rect 2488 1472 2520 1504
rect 2560 1472 2592 1504
rect 2632 1472 2664 1504
rect 2704 1472 2736 1504
rect 2776 1472 2808 1504
rect 2848 1472 2880 1504
rect 2920 1472 2952 1504
rect 2992 1472 3024 1504
rect 3064 1472 3096 1504
rect 3136 1472 3168 1504
rect 3208 1472 3240 1504
rect 3280 1472 3312 1504
rect 3352 1472 3384 1504
rect 3424 1472 3456 1504
rect 3496 1472 3528 1504
rect 3568 1472 3600 1504
rect 3640 1472 3672 1504
rect 3712 1472 3744 1504
rect 3784 1472 3816 1504
rect 3856 1472 3888 1504
rect 3928 1472 3960 1504
rect 40 1400 72 1432
rect 112 1400 144 1432
rect 184 1400 216 1432
rect 256 1400 288 1432
rect 328 1400 360 1432
rect 400 1400 432 1432
rect 472 1400 504 1432
rect 544 1400 576 1432
rect 616 1400 648 1432
rect 688 1400 720 1432
rect 760 1400 792 1432
rect 832 1400 864 1432
rect 904 1400 936 1432
rect 976 1400 1008 1432
rect 1048 1400 1080 1432
rect 1120 1400 1152 1432
rect 1192 1400 1224 1432
rect 1264 1400 1296 1432
rect 1336 1400 1368 1432
rect 1408 1400 1440 1432
rect 1480 1400 1512 1432
rect 1552 1400 1584 1432
rect 1624 1400 1656 1432
rect 1696 1400 1728 1432
rect 1768 1400 1800 1432
rect 1840 1400 1872 1432
rect 1912 1400 1944 1432
rect 1984 1400 2016 1432
rect 2056 1400 2088 1432
rect 2128 1400 2160 1432
rect 2200 1400 2232 1432
rect 2272 1400 2304 1432
rect 2344 1400 2376 1432
rect 2416 1400 2448 1432
rect 2488 1400 2520 1432
rect 2560 1400 2592 1432
rect 2632 1400 2664 1432
rect 2704 1400 2736 1432
rect 2776 1400 2808 1432
rect 2848 1400 2880 1432
rect 2920 1400 2952 1432
rect 2992 1400 3024 1432
rect 3064 1400 3096 1432
rect 3136 1400 3168 1432
rect 3208 1400 3240 1432
rect 3280 1400 3312 1432
rect 3352 1400 3384 1432
rect 3424 1400 3456 1432
rect 3496 1400 3528 1432
rect 3568 1400 3600 1432
rect 3640 1400 3672 1432
rect 3712 1400 3744 1432
rect 3784 1400 3816 1432
rect 3856 1400 3888 1432
rect 3928 1400 3960 1432
rect 40 1328 72 1360
rect 112 1328 144 1360
rect 184 1328 216 1360
rect 256 1328 288 1360
rect 328 1328 360 1360
rect 400 1328 432 1360
rect 472 1328 504 1360
rect 544 1328 576 1360
rect 616 1328 648 1360
rect 688 1328 720 1360
rect 760 1328 792 1360
rect 832 1328 864 1360
rect 904 1328 936 1360
rect 976 1328 1008 1360
rect 1048 1328 1080 1360
rect 1120 1328 1152 1360
rect 1192 1328 1224 1360
rect 1264 1328 1296 1360
rect 1336 1328 1368 1360
rect 1408 1328 1440 1360
rect 1480 1328 1512 1360
rect 1552 1328 1584 1360
rect 1624 1328 1656 1360
rect 1696 1328 1728 1360
rect 1768 1328 1800 1360
rect 1840 1328 1872 1360
rect 1912 1328 1944 1360
rect 1984 1328 2016 1360
rect 2056 1328 2088 1360
rect 2128 1328 2160 1360
rect 2200 1328 2232 1360
rect 2272 1328 2304 1360
rect 2344 1328 2376 1360
rect 2416 1328 2448 1360
rect 2488 1328 2520 1360
rect 2560 1328 2592 1360
rect 2632 1328 2664 1360
rect 2704 1328 2736 1360
rect 2776 1328 2808 1360
rect 2848 1328 2880 1360
rect 2920 1328 2952 1360
rect 2992 1328 3024 1360
rect 3064 1328 3096 1360
rect 3136 1328 3168 1360
rect 3208 1328 3240 1360
rect 3280 1328 3312 1360
rect 3352 1328 3384 1360
rect 3424 1328 3456 1360
rect 3496 1328 3528 1360
rect 3568 1328 3600 1360
rect 3640 1328 3672 1360
rect 3712 1328 3744 1360
rect 3784 1328 3816 1360
rect 3856 1328 3888 1360
rect 3928 1328 3960 1360
rect 40 1256 72 1288
rect 112 1256 144 1288
rect 184 1256 216 1288
rect 256 1256 288 1288
rect 328 1256 360 1288
rect 400 1256 432 1288
rect 472 1256 504 1288
rect 544 1256 576 1288
rect 616 1256 648 1288
rect 688 1256 720 1288
rect 760 1256 792 1288
rect 832 1256 864 1288
rect 904 1256 936 1288
rect 976 1256 1008 1288
rect 1048 1256 1080 1288
rect 1120 1256 1152 1288
rect 1192 1256 1224 1288
rect 1264 1256 1296 1288
rect 1336 1256 1368 1288
rect 1408 1256 1440 1288
rect 1480 1256 1512 1288
rect 1552 1256 1584 1288
rect 1624 1256 1656 1288
rect 1696 1256 1728 1288
rect 1768 1256 1800 1288
rect 1840 1256 1872 1288
rect 1912 1256 1944 1288
rect 1984 1256 2016 1288
rect 2056 1256 2088 1288
rect 2128 1256 2160 1288
rect 2200 1256 2232 1288
rect 2272 1256 2304 1288
rect 2344 1256 2376 1288
rect 2416 1256 2448 1288
rect 2488 1256 2520 1288
rect 2560 1256 2592 1288
rect 2632 1256 2664 1288
rect 2704 1256 2736 1288
rect 2776 1256 2808 1288
rect 2848 1256 2880 1288
rect 2920 1256 2952 1288
rect 2992 1256 3024 1288
rect 3064 1256 3096 1288
rect 3136 1256 3168 1288
rect 3208 1256 3240 1288
rect 3280 1256 3312 1288
rect 3352 1256 3384 1288
rect 3424 1256 3456 1288
rect 3496 1256 3528 1288
rect 3568 1256 3600 1288
rect 3640 1256 3672 1288
rect 3712 1256 3744 1288
rect 3784 1256 3816 1288
rect 3856 1256 3888 1288
rect 3928 1256 3960 1288
rect 0 33416 4000 33430
rect 0 33384 112 33416
rect 144 33384 184 33416
rect 216 33384 256 33416
rect 288 33384 328 33416
rect 360 33384 400 33416
rect 432 33384 472 33416
rect 504 33384 544 33416
rect 576 33384 616 33416
rect 648 33384 688 33416
rect 720 33384 760 33416
rect 792 33384 832 33416
rect 864 33384 904 33416
rect 936 33384 976 33416
rect 1008 33384 1048 33416
rect 1080 33384 1120 33416
rect 1152 33384 1192 33416
rect 1224 33384 1264 33416
rect 1296 33384 1336 33416
rect 1368 33384 1408 33416
rect 1440 33384 1480 33416
rect 1512 33384 1552 33416
rect 1584 33384 1624 33416
rect 1656 33384 1696 33416
rect 1728 33384 1768 33416
rect 1800 33384 1840 33416
rect 1872 33384 1912 33416
rect 1944 33384 1984 33416
rect 2016 33384 2056 33416
rect 2088 33384 2128 33416
rect 2160 33384 2200 33416
rect 2232 33384 2272 33416
rect 2304 33384 2344 33416
rect 2376 33384 2416 33416
rect 2448 33384 2488 33416
rect 2520 33384 2560 33416
rect 2592 33384 2632 33416
rect 2664 33384 2704 33416
rect 2736 33384 2776 33416
rect 2808 33384 2848 33416
rect 2880 33384 2920 33416
rect 2952 33384 2992 33416
rect 3024 33384 3064 33416
rect 3096 33384 3136 33416
rect 3168 33384 3208 33416
rect 3240 33384 3280 33416
rect 3312 33384 3352 33416
rect 3384 33384 3424 33416
rect 3456 33384 3496 33416
rect 3528 33384 3568 33416
rect 3600 33384 3640 33416
rect 3672 33384 3712 33416
rect 3744 33384 3784 33416
rect 3816 33384 3856 33416
rect 3888 33384 4000 33416
rect 0 33370 4000 33384
rect 0 29716 4000 29730
rect 0 29684 112 29716
rect 144 29684 184 29716
rect 216 29684 256 29716
rect 288 29684 328 29716
rect 360 29684 400 29716
rect 432 29684 472 29716
rect 504 29684 544 29716
rect 576 29684 616 29716
rect 648 29684 688 29716
rect 720 29684 760 29716
rect 792 29684 832 29716
rect 864 29684 904 29716
rect 936 29684 976 29716
rect 1008 29684 1048 29716
rect 1080 29684 1120 29716
rect 1152 29684 1192 29716
rect 1224 29684 1264 29716
rect 1296 29684 1336 29716
rect 1368 29684 1408 29716
rect 1440 29684 1480 29716
rect 1512 29684 1552 29716
rect 1584 29684 1624 29716
rect 1656 29684 1696 29716
rect 1728 29684 1768 29716
rect 1800 29684 1840 29716
rect 1872 29684 1912 29716
rect 1944 29684 1984 29716
rect 2016 29684 2056 29716
rect 2088 29684 2128 29716
rect 2160 29684 2200 29716
rect 2232 29684 2272 29716
rect 2304 29684 2344 29716
rect 2376 29684 2416 29716
rect 2448 29684 2488 29716
rect 2520 29684 2560 29716
rect 2592 29684 2632 29716
rect 2664 29684 2704 29716
rect 2736 29684 2776 29716
rect 2808 29684 2848 29716
rect 2880 29684 2920 29716
rect 2952 29684 2992 29716
rect 3024 29684 3064 29716
rect 3096 29684 3136 29716
rect 3168 29684 3208 29716
rect 3240 29684 3280 29716
rect 3312 29684 3352 29716
rect 3384 29684 3424 29716
rect 3456 29684 3496 29716
rect 3528 29684 3568 29716
rect 3600 29684 3640 29716
rect 3672 29684 3712 29716
rect 3744 29684 3784 29716
rect 3816 29684 3856 29716
rect 3888 29684 4000 29716
rect 0 29670 4000 29684
rect 0 12144 4000 12200
rect 0 12112 40 12144
rect 72 12112 112 12144
rect 144 12112 184 12144
rect 216 12112 256 12144
rect 288 12112 328 12144
rect 360 12112 400 12144
rect 432 12112 472 12144
rect 504 12112 544 12144
rect 576 12112 616 12144
rect 648 12112 688 12144
rect 720 12112 760 12144
rect 792 12112 832 12144
rect 864 12112 904 12144
rect 936 12112 976 12144
rect 1008 12112 1048 12144
rect 1080 12112 1120 12144
rect 1152 12112 1192 12144
rect 1224 12112 1264 12144
rect 1296 12112 1336 12144
rect 1368 12112 1408 12144
rect 1440 12112 1480 12144
rect 1512 12112 1552 12144
rect 1584 12112 1624 12144
rect 1656 12112 1696 12144
rect 1728 12112 1768 12144
rect 1800 12112 1840 12144
rect 1872 12112 1912 12144
rect 1944 12112 1984 12144
rect 2016 12112 2056 12144
rect 2088 12112 2128 12144
rect 2160 12112 2200 12144
rect 2232 12112 2272 12144
rect 2304 12112 2344 12144
rect 2376 12112 2416 12144
rect 2448 12112 2488 12144
rect 2520 12112 2560 12144
rect 2592 12112 2632 12144
rect 2664 12112 2704 12144
rect 2736 12112 2776 12144
rect 2808 12112 2848 12144
rect 2880 12112 2920 12144
rect 2952 12112 2992 12144
rect 3024 12112 3064 12144
rect 3096 12112 3136 12144
rect 3168 12112 3208 12144
rect 3240 12112 3280 12144
rect 3312 12112 3352 12144
rect 3384 12112 3424 12144
rect 3456 12112 3496 12144
rect 3528 12112 3568 12144
rect 3600 12112 3640 12144
rect 3672 12112 3712 12144
rect 3744 12112 3784 12144
rect 3816 12112 3856 12144
rect 3888 12112 3928 12144
rect 3960 12112 4000 12144
rect 0 12072 4000 12112
rect 0 12040 40 12072
rect 72 12040 112 12072
rect 144 12040 184 12072
rect 216 12040 256 12072
rect 288 12040 328 12072
rect 360 12040 400 12072
rect 432 12040 472 12072
rect 504 12040 544 12072
rect 576 12040 616 12072
rect 648 12040 688 12072
rect 720 12040 760 12072
rect 792 12040 832 12072
rect 864 12040 904 12072
rect 936 12040 976 12072
rect 1008 12040 1048 12072
rect 1080 12040 1120 12072
rect 1152 12040 1192 12072
rect 1224 12040 1264 12072
rect 1296 12040 1336 12072
rect 1368 12040 1408 12072
rect 1440 12040 1480 12072
rect 1512 12040 1552 12072
rect 1584 12040 1624 12072
rect 1656 12040 1696 12072
rect 1728 12040 1768 12072
rect 1800 12040 1840 12072
rect 1872 12040 1912 12072
rect 1944 12040 1984 12072
rect 2016 12040 2056 12072
rect 2088 12040 2128 12072
rect 2160 12040 2200 12072
rect 2232 12040 2272 12072
rect 2304 12040 2344 12072
rect 2376 12040 2416 12072
rect 2448 12040 2488 12072
rect 2520 12040 2560 12072
rect 2592 12040 2632 12072
rect 2664 12040 2704 12072
rect 2736 12040 2776 12072
rect 2808 12040 2848 12072
rect 2880 12040 2920 12072
rect 2952 12040 2992 12072
rect 3024 12040 3064 12072
rect 3096 12040 3136 12072
rect 3168 12040 3208 12072
rect 3240 12040 3280 12072
rect 3312 12040 3352 12072
rect 3384 12040 3424 12072
rect 3456 12040 3496 12072
rect 3528 12040 3568 12072
rect 3600 12040 3640 12072
rect 3672 12040 3712 12072
rect 3744 12040 3784 12072
rect 3816 12040 3856 12072
rect 3888 12040 3928 12072
rect 3960 12040 4000 12072
rect 0 12000 4000 12040
rect 0 11968 40 12000
rect 72 11968 112 12000
rect 144 11968 184 12000
rect 216 11968 256 12000
rect 288 11968 328 12000
rect 360 11968 400 12000
rect 432 11968 472 12000
rect 504 11968 544 12000
rect 576 11968 616 12000
rect 648 11968 688 12000
rect 720 11968 760 12000
rect 792 11968 832 12000
rect 864 11968 904 12000
rect 936 11968 976 12000
rect 1008 11968 1048 12000
rect 1080 11968 1120 12000
rect 1152 11968 1192 12000
rect 1224 11968 1264 12000
rect 1296 11968 1336 12000
rect 1368 11968 1408 12000
rect 1440 11968 1480 12000
rect 1512 11968 1552 12000
rect 1584 11968 1624 12000
rect 1656 11968 1696 12000
rect 1728 11968 1768 12000
rect 1800 11968 1840 12000
rect 1872 11968 1912 12000
rect 1944 11968 1984 12000
rect 2016 11968 2056 12000
rect 2088 11968 2128 12000
rect 2160 11968 2200 12000
rect 2232 11968 2272 12000
rect 2304 11968 2344 12000
rect 2376 11968 2416 12000
rect 2448 11968 2488 12000
rect 2520 11968 2560 12000
rect 2592 11968 2632 12000
rect 2664 11968 2704 12000
rect 2736 11968 2776 12000
rect 2808 11968 2848 12000
rect 2880 11968 2920 12000
rect 2952 11968 2992 12000
rect 3024 11968 3064 12000
rect 3096 11968 3136 12000
rect 3168 11968 3208 12000
rect 3240 11968 3280 12000
rect 3312 11968 3352 12000
rect 3384 11968 3424 12000
rect 3456 11968 3496 12000
rect 3528 11968 3568 12000
rect 3600 11968 3640 12000
rect 3672 11968 3712 12000
rect 3744 11968 3784 12000
rect 3816 11968 3856 12000
rect 3888 11968 3928 12000
rect 3960 11968 4000 12000
rect 0 11928 4000 11968
rect 0 11896 40 11928
rect 72 11896 112 11928
rect 144 11896 184 11928
rect 216 11896 256 11928
rect 288 11896 328 11928
rect 360 11896 400 11928
rect 432 11896 472 11928
rect 504 11896 544 11928
rect 576 11896 616 11928
rect 648 11896 688 11928
rect 720 11896 760 11928
rect 792 11896 832 11928
rect 864 11896 904 11928
rect 936 11896 976 11928
rect 1008 11896 1048 11928
rect 1080 11896 1120 11928
rect 1152 11896 1192 11928
rect 1224 11896 1264 11928
rect 1296 11896 1336 11928
rect 1368 11896 1408 11928
rect 1440 11896 1480 11928
rect 1512 11896 1552 11928
rect 1584 11896 1624 11928
rect 1656 11896 1696 11928
rect 1728 11896 1768 11928
rect 1800 11896 1840 11928
rect 1872 11896 1912 11928
rect 1944 11896 1984 11928
rect 2016 11896 2056 11928
rect 2088 11896 2128 11928
rect 2160 11896 2200 11928
rect 2232 11896 2272 11928
rect 2304 11896 2344 11928
rect 2376 11896 2416 11928
rect 2448 11896 2488 11928
rect 2520 11896 2560 11928
rect 2592 11896 2632 11928
rect 2664 11896 2704 11928
rect 2736 11896 2776 11928
rect 2808 11896 2848 11928
rect 2880 11896 2920 11928
rect 2952 11896 2992 11928
rect 3024 11896 3064 11928
rect 3096 11896 3136 11928
rect 3168 11896 3208 11928
rect 3240 11896 3280 11928
rect 3312 11896 3352 11928
rect 3384 11896 3424 11928
rect 3456 11896 3496 11928
rect 3528 11896 3568 11928
rect 3600 11896 3640 11928
rect 3672 11896 3712 11928
rect 3744 11896 3784 11928
rect 3816 11896 3856 11928
rect 3888 11896 3928 11928
rect 3960 11896 4000 11928
rect 0 11856 4000 11896
rect 0 11824 40 11856
rect 72 11824 112 11856
rect 144 11824 184 11856
rect 216 11824 256 11856
rect 288 11824 328 11856
rect 360 11824 400 11856
rect 432 11824 472 11856
rect 504 11824 544 11856
rect 576 11824 616 11856
rect 648 11824 688 11856
rect 720 11824 760 11856
rect 792 11824 832 11856
rect 864 11824 904 11856
rect 936 11824 976 11856
rect 1008 11824 1048 11856
rect 1080 11824 1120 11856
rect 1152 11824 1192 11856
rect 1224 11824 1264 11856
rect 1296 11824 1336 11856
rect 1368 11824 1408 11856
rect 1440 11824 1480 11856
rect 1512 11824 1552 11856
rect 1584 11824 1624 11856
rect 1656 11824 1696 11856
rect 1728 11824 1768 11856
rect 1800 11824 1840 11856
rect 1872 11824 1912 11856
rect 1944 11824 1984 11856
rect 2016 11824 2056 11856
rect 2088 11824 2128 11856
rect 2160 11824 2200 11856
rect 2232 11824 2272 11856
rect 2304 11824 2344 11856
rect 2376 11824 2416 11856
rect 2448 11824 2488 11856
rect 2520 11824 2560 11856
rect 2592 11824 2632 11856
rect 2664 11824 2704 11856
rect 2736 11824 2776 11856
rect 2808 11824 2848 11856
rect 2880 11824 2920 11856
rect 2952 11824 2992 11856
rect 3024 11824 3064 11856
rect 3096 11824 3136 11856
rect 3168 11824 3208 11856
rect 3240 11824 3280 11856
rect 3312 11824 3352 11856
rect 3384 11824 3424 11856
rect 3456 11824 3496 11856
rect 3528 11824 3568 11856
rect 3600 11824 3640 11856
rect 3672 11824 3712 11856
rect 3744 11824 3784 11856
rect 3816 11824 3856 11856
rect 3888 11824 3928 11856
rect 3960 11824 4000 11856
rect 0 11784 4000 11824
rect 0 11752 40 11784
rect 72 11752 112 11784
rect 144 11752 184 11784
rect 216 11752 256 11784
rect 288 11752 328 11784
rect 360 11752 400 11784
rect 432 11752 472 11784
rect 504 11752 544 11784
rect 576 11752 616 11784
rect 648 11752 688 11784
rect 720 11752 760 11784
rect 792 11752 832 11784
rect 864 11752 904 11784
rect 936 11752 976 11784
rect 1008 11752 1048 11784
rect 1080 11752 1120 11784
rect 1152 11752 1192 11784
rect 1224 11752 1264 11784
rect 1296 11752 1336 11784
rect 1368 11752 1408 11784
rect 1440 11752 1480 11784
rect 1512 11752 1552 11784
rect 1584 11752 1624 11784
rect 1656 11752 1696 11784
rect 1728 11752 1768 11784
rect 1800 11752 1840 11784
rect 1872 11752 1912 11784
rect 1944 11752 1984 11784
rect 2016 11752 2056 11784
rect 2088 11752 2128 11784
rect 2160 11752 2200 11784
rect 2232 11752 2272 11784
rect 2304 11752 2344 11784
rect 2376 11752 2416 11784
rect 2448 11752 2488 11784
rect 2520 11752 2560 11784
rect 2592 11752 2632 11784
rect 2664 11752 2704 11784
rect 2736 11752 2776 11784
rect 2808 11752 2848 11784
rect 2880 11752 2920 11784
rect 2952 11752 2992 11784
rect 3024 11752 3064 11784
rect 3096 11752 3136 11784
rect 3168 11752 3208 11784
rect 3240 11752 3280 11784
rect 3312 11752 3352 11784
rect 3384 11752 3424 11784
rect 3456 11752 3496 11784
rect 3528 11752 3568 11784
rect 3600 11752 3640 11784
rect 3672 11752 3712 11784
rect 3744 11752 3784 11784
rect 3816 11752 3856 11784
rect 3888 11752 3928 11784
rect 3960 11752 4000 11784
rect 0 11712 4000 11752
rect 0 11680 40 11712
rect 72 11680 112 11712
rect 144 11680 184 11712
rect 216 11680 256 11712
rect 288 11680 328 11712
rect 360 11680 400 11712
rect 432 11680 472 11712
rect 504 11680 544 11712
rect 576 11680 616 11712
rect 648 11680 688 11712
rect 720 11680 760 11712
rect 792 11680 832 11712
rect 864 11680 904 11712
rect 936 11680 976 11712
rect 1008 11680 1048 11712
rect 1080 11680 1120 11712
rect 1152 11680 1192 11712
rect 1224 11680 1264 11712
rect 1296 11680 1336 11712
rect 1368 11680 1408 11712
rect 1440 11680 1480 11712
rect 1512 11680 1552 11712
rect 1584 11680 1624 11712
rect 1656 11680 1696 11712
rect 1728 11680 1768 11712
rect 1800 11680 1840 11712
rect 1872 11680 1912 11712
rect 1944 11680 1984 11712
rect 2016 11680 2056 11712
rect 2088 11680 2128 11712
rect 2160 11680 2200 11712
rect 2232 11680 2272 11712
rect 2304 11680 2344 11712
rect 2376 11680 2416 11712
rect 2448 11680 2488 11712
rect 2520 11680 2560 11712
rect 2592 11680 2632 11712
rect 2664 11680 2704 11712
rect 2736 11680 2776 11712
rect 2808 11680 2848 11712
rect 2880 11680 2920 11712
rect 2952 11680 2992 11712
rect 3024 11680 3064 11712
rect 3096 11680 3136 11712
rect 3168 11680 3208 11712
rect 3240 11680 3280 11712
rect 3312 11680 3352 11712
rect 3384 11680 3424 11712
rect 3456 11680 3496 11712
rect 3528 11680 3568 11712
rect 3600 11680 3640 11712
rect 3672 11680 3712 11712
rect 3744 11680 3784 11712
rect 3816 11680 3856 11712
rect 3888 11680 3928 11712
rect 3960 11680 4000 11712
rect 0 11640 4000 11680
rect 0 11608 40 11640
rect 72 11608 112 11640
rect 144 11608 184 11640
rect 216 11608 256 11640
rect 288 11608 328 11640
rect 360 11608 400 11640
rect 432 11608 472 11640
rect 504 11608 544 11640
rect 576 11608 616 11640
rect 648 11608 688 11640
rect 720 11608 760 11640
rect 792 11608 832 11640
rect 864 11608 904 11640
rect 936 11608 976 11640
rect 1008 11608 1048 11640
rect 1080 11608 1120 11640
rect 1152 11608 1192 11640
rect 1224 11608 1264 11640
rect 1296 11608 1336 11640
rect 1368 11608 1408 11640
rect 1440 11608 1480 11640
rect 1512 11608 1552 11640
rect 1584 11608 1624 11640
rect 1656 11608 1696 11640
rect 1728 11608 1768 11640
rect 1800 11608 1840 11640
rect 1872 11608 1912 11640
rect 1944 11608 1984 11640
rect 2016 11608 2056 11640
rect 2088 11608 2128 11640
rect 2160 11608 2200 11640
rect 2232 11608 2272 11640
rect 2304 11608 2344 11640
rect 2376 11608 2416 11640
rect 2448 11608 2488 11640
rect 2520 11608 2560 11640
rect 2592 11608 2632 11640
rect 2664 11608 2704 11640
rect 2736 11608 2776 11640
rect 2808 11608 2848 11640
rect 2880 11608 2920 11640
rect 2952 11608 2992 11640
rect 3024 11608 3064 11640
rect 3096 11608 3136 11640
rect 3168 11608 3208 11640
rect 3240 11608 3280 11640
rect 3312 11608 3352 11640
rect 3384 11608 3424 11640
rect 3456 11608 3496 11640
rect 3528 11608 3568 11640
rect 3600 11608 3640 11640
rect 3672 11608 3712 11640
rect 3744 11608 3784 11640
rect 3816 11608 3856 11640
rect 3888 11608 3928 11640
rect 3960 11608 4000 11640
rect 0 11568 4000 11608
rect 0 11536 40 11568
rect 72 11536 112 11568
rect 144 11536 184 11568
rect 216 11536 256 11568
rect 288 11536 328 11568
rect 360 11536 400 11568
rect 432 11536 472 11568
rect 504 11536 544 11568
rect 576 11536 616 11568
rect 648 11536 688 11568
rect 720 11536 760 11568
rect 792 11536 832 11568
rect 864 11536 904 11568
rect 936 11536 976 11568
rect 1008 11536 1048 11568
rect 1080 11536 1120 11568
rect 1152 11536 1192 11568
rect 1224 11536 1264 11568
rect 1296 11536 1336 11568
rect 1368 11536 1408 11568
rect 1440 11536 1480 11568
rect 1512 11536 1552 11568
rect 1584 11536 1624 11568
rect 1656 11536 1696 11568
rect 1728 11536 1768 11568
rect 1800 11536 1840 11568
rect 1872 11536 1912 11568
rect 1944 11536 1984 11568
rect 2016 11536 2056 11568
rect 2088 11536 2128 11568
rect 2160 11536 2200 11568
rect 2232 11536 2272 11568
rect 2304 11536 2344 11568
rect 2376 11536 2416 11568
rect 2448 11536 2488 11568
rect 2520 11536 2560 11568
rect 2592 11536 2632 11568
rect 2664 11536 2704 11568
rect 2736 11536 2776 11568
rect 2808 11536 2848 11568
rect 2880 11536 2920 11568
rect 2952 11536 2992 11568
rect 3024 11536 3064 11568
rect 3096 11536 3136 11568
rect 3168 11536 3208 11568
rect 3240 11536 3280 11568
rect 3312 11536 3352 11568
rect 3384 11536 3424 11568
rect 3456 11536 3496 11568
rect 3528 11536 3568 11568
rect 3600 11536 3640 11568
rect 3672 11536 3712 11568
rect 3744 11536 3784 11568
rect 3816 11536 3856 11568
rect 3888 11536 3928 11568
rect 3960 11536 4000 11568
rect 0 11496 4000 11536
rect 0 11464 40 11496
rect 72 11464 112 11496
rect 144 11464 184 11496
rect 216 11464 256 11496
rect 288 11464 328 11496
rect 360 11464 400 11496
rect 432 11464 472 11496
rect 504 11464 544 11496
rect 576 11464 616 11496
rect 648 11464 688 11496
rect 720 11464 760 11496
rect 792 11464 832 11496
rect 864 11464 904 11496
rect 936 11464 976 11496
rect 1008 11464 1048 11496
rect 1080 11464 1120 11496
rect 1152 11464 1192 11496
rect 1224 11464 1264 11496
rect 1296 11464 1336 11496
rect 1368 11464 1408 11496
rect 1440 11464 1480 11496
rect 1512 11464 1552 11496
rect 1584 11464 1624 11496
rect 1656 11464 1696 11496
rect 1728 11464 1768 11496
rect 1800 11464 1840 11496
rect 1872 11464 1912 11496
rect 1944 11464 1984 11496
rect 2016 11464 2056 11496
rect 2088 11464 2128 11496
rect 2160 11464 2200 11496
rect 2232 11464 2272 11496
rect 2304 11464 2344 11496
rect 2376 11464 2416 11496
rect 2448 11464 2488 11496
rect 2520 11464 2560 11496
rect 2592 11464 2632 11496
rect 2664 11464 2704 11496
rect 2736 11464 2776 11496
rect 2808 11464 2848 11496
rect 2880 11464 2920 11496
rect 2952 11464 2992 11496
rect 3024 11464 3064 11496
rect 3096 11464 3136 11496
rect 3168 11464 3208 11496
rect 3240 11464 3280 11496
rect 3312 11464 3352 11496
rect 3384 11464 3424 11496
rect 3456 11464 3496 11496
rect 3528 11464 3568 11496
rect 3600 11464 3640 11496
rect 3672 11464 3712 11496
rect 3744 11464 3784 11496
rect 3816 11464 3856 11496
rect 3888 11464 3928 11496
rect 3960 11464 4000 11496
rect 0 11424 4000 11464
rect 0 11392 40 11424
rect 72 11392 112 11424
rect 144 11392 184 11424
rect 216 11392 256 11424
rect 288 11392 328 11424
rect 360 11392 400 11424
rect 432 11392 472 11424
rect 504 11392 544 11424
rect 576 11392 616 11424
rect 648 11392 688 11424
rect 720 11392 760 11424
rect 792 11392 832 11424
rect 864 11392 904 11424
rect 936 11392 976 11424
rect 1008 11392 1048 11424
rect 1080 11392 1120 11424
rect 1152 11392 1192 11424
rect 1224 11392 1264 11424
rect 1296 11392 1336 11424
rect 1368 11392 1408 11424
rect 1440 11392 1480 11424
rect 1512 11392 1552 11424
rect 1584 11392 1624 11424
rect 1656 11392 1696 11424
rect 1728 11392 1768 11424
rect 1800 11392 1840 11424
rect 1872 11392 1912 11424
rect 1944 11392 1984 11424
rect 2016 11392 2056 11424
rect 2088 11392 2128 11424
rect 2160 11392 2200 11424
rect 2232 11392 2272 11424
rect 2304 11392 2344 11424
rect 2376 11392 2416 11424
rect 2448 11392 2488 11424
rect 2520 11392 2560 11424
rect 2592 11392 2632 11424
rect 2664 11392 2704 11424
rect 2736 11392 2776 11424
rect 2808 11392 2848 11424
rect 2880 11392 2920 11424
rect 2952 11392 2992 11424
rect 3024 11392 3064 11424
rect 3096 11392 3136 11424
rect 3168 11392 3208 11424
rect 3240 11392 3280 11424
rect 3312 11392 3352 11424
rect 3384 11392 3424 11424
rect 3456 11392 3496 11424
rect 3528 11392 3568 11424
rect 3600 11392 3640 11424
rect 3672 11392 3712 11424
rect 3744 11392 3784 11424
rect 3816 11392 3856 11424
rect 3888 11392 3928 11424
rect 3960 11392 4000 11424
rect 0 11352 4000 11392
rect 0 11320 40 11352
rect 72 11320 112 11352
rect 144 11320 184 11352
rect 216 11320 256 11352
rect 288 11320 328 11352
rect 360 11320 400 11352
rect 432 11320 472 11352
rect 504 11320 544 11352
rect 576 11320 616 11352
rect 648 11320 688 11352
rect 720 11320 760 11352
rect 792 11320 832 11352
rect 864 11320 904 11352
rect 936 11320 976 11352
rect 1008 11320 1048 11352
rect 1080 11320 1120 11352
rect 1152 11320 1192 11352
rect 1224 11320 1264 11352
rect 1296 11320 1336 11352
rect 1368 11320 1408 11352
rect 1440 11320 1480 11352
rect 1512 11320 1552 11352
rect 1584 11320 1624 11352
rect 1656 11320 1696 11352
rect 1728 11320 1768 11352
rect 1800 11320 1840 11352
rect 1872 11320 1912 11352
rect 1944 11320 1984 11352
rect 2016 11320 2056 11352
rect 2088 11320 2128 11352
rect 2160 11320 2200 11352
rect 2232 11320 2272 11352
rect 2304 11320 2344 11352
rect 2376 11320 2416 11352
rect 2448 11320 2488 11352
rect 2520 11320 2560 11352
rect 2592 11320 2632 11352
rect 2664 11320 2704 11352
rect 2736 11320 2776 11352
rect 2808 11320 2848 11352
rect 2880 11320 2920 11352
rect 2952 11320 2992 11352
rect 3024 11320 3064 11352
rect 3096 11320 3136 11352
rect 3168 11320 3208 11352
rect 3240 11320 3280 11352
rect 3312 11320 3352 11352
rect 3384 11320 3424 11352
rect 3456 11320 3496 11352
rect 3528 11320 3568 11352
rect 3600 11320 3640 11352
rect 3672 11320 3712 11352
rect 3744 11320 3784 11352
rect 3816 11320 3856 11352
rect 3888 11320 3928 11352
rect 3960 11320 4000 11352
rect 0 11280 4000 11320
rect 0 11248 40 11280
rect 72 11248 112 11280
rect 144 11248 184 11280
rect 216 11248 256 11280
rect 288 11248 328 11280
rect 360 11248 400 11280
rect 432 11248 472 11280
rect 504 11248 544 11280
rect 576 11248 616 11280
rect 648 11248 688 11280
rect 720 11248 760 11280
rect 792 11248 832 11280
rect 864 11248 904 11280
rect 936 11248 976 11280
rect 1008 11248 1048 11280
rect 1080 11248 1120 11280
rect 1152 11248 1192 11280
rect 1224 11248 1264 11280
rect 1296 11248 1336 11280
rect 1368 11248 1408 11280
rect 1440 11248 1480 11280
rect 1512 11248 1552 11280
rect 1584 11248 1624 11280
rect 1656 11248 1696 11280
rect 1728 11248 1768 11280
rect 1800 11248 1840 11280
rect 1872 11248 1912 11280
rect 1944 11248 1984 11280
rect 2016 11248 2056 11280
rect 2088 11248 2128 11280
rect 2160 11248 2200 11280
rect 2232 11248 2272 11280
rect 2304 11248 2344 11280
rect 2376 11248 2416 11280
rect 2448 11248 2488 11280
rect 2520 11248 2560 11280
rect 2592 11248 2632 11280
rect 2664 11248 2704 11280
rect 2736 11248 2776 11280
rect 2808 11248 2848 11280
rect 2880 11248 2920 11280
rect 2952 11248 2992 11280
rect 3024 11248 3064 11280
rect 3096 11248 3136 11280
rect 3168 11248 3208 11280
rect 3240 11248 3280 11280
rect 3312 11248 3352 11280
rect 3384 11248 3424 11280
rect 3456 11248 3496 11280
rect 3528 11248 3568 11280
rect 3600 11248 3640 11280
rect 3672 11248 3712 11280
rect 3744 11248 3784 11280
rect 3816 11248 3856 11280
rect 3888 11248 3928 11280
rect 3960 11248 4000 11280
rect 0 11208 4000 11248
rect 0 11176 40 11208
rect 72 11176 112 11208
rect 144 11176 184 11208
rect 216 11176 256 11208
rect 288 11176 328 11208
rect 360 11176 400 11208
rect 432 11176 472 11208
rect 504 11176 544 11208
rect 576 11176 616 11208
rect 648 11176 688 11208
rect 720 11176 760 11208
rect 792 11176 832 11208
rect 864 11176 904 11208
rect 936 11176 976 11208
rect 1008 11176 1048 11208
rect 1080 11176 1120 11208
rect 1152 11176 1192 11208
rect 1224 11176 1264 11208
rect 1296 11176 1336 11208
rect 1368 11176 1408 11208
rect 1440 11176 1480 11208
rect 1512 11176 1552 11208
rect 1584 11176 1624 11208
rect 1656 11176 1696 11208
rect 1728 11176 1768 11208
rect 1800 11176 1840 11208
rect 1872 11176 1912 11208
rect 1944 11176 1984 11208
rect 2016 11176 2056 11208
rect 2088 11176 2128 11208
rect 2160 11176 2200 11208
rect 2232 11176 2272 11208
rect 2304 11176 2344 11208
rect 2376 11176 2416 11208
rect 2448 11176 2488 11208
rect 2520 11176 2560 11208
rect 2592 11176 2632 11208
rect 2664 11176 2704 11208
rect 2736 11176 2776 11208
rect 2808 11176 2848 11208
rect 2880 11176 2920 11208
rect 2952 11176 2992 11208
rect 3024 11176 3064 11208
rect 3096 11176 3136 11208
rect 3168 11176 3208 11208
rect 3240 11176 3280 11208
rect 3312 11176 3352 11208
rect 3384 11176 3424 11208
rect 3456 11176 3496 11208
rect 3528 11176 3568 11208
rect 3600 11176 3640 11208
rect 3672 11176 3712 11208
rect 3744 11176 3784 11208
rect 3816 11176 3856 11208
rect 3888 11176 3928 11208
rect 3960 11176 4000 11208
rect 0 11136 4000 11176
rect 0 11104 40 11136
rect 72 11104 112 11136
rect 144 11104 184 11136
rect 216 11104 256 11136
rect 288 11104 328 11136
rect 360 11104 400 11136
rect 432 11104 472 11136
rect 504 11104 544 11136
rect 576 11104 616 11136
rect 648 11104 688 11136
rect 720 11104 760 11136
rect 792 11104 832 11136
rect 864 11104 904 11136
rect 936 11104 976 11136
rect 1008 11104 1048 11136
rect 1080 11104 1120 11136
rect 1152 11104 1192 11136
rect 1224 11104 1264 11136
rect 1296 11104 1336 11136
rect 1368 11104 1408 11136
rect 1440 11104 1480 11136
rect 1512 11104 1552 11136
rect 1584 11104 1624 11136
rect 1656 11104 1696 11136
rect 1728 11104 1768 11136
rect 1800 11104 1840 11136
rect 1872 11104 1912 11136
rect 1944 11104 1984 11136
rect 2016 11104 2056 11136
rect 2088 11104 2128 11136
rect 2160 11104 2200 11136
rect 2232 11104 2272 11136
rect 2304 11104 2344 11136
rect 2376 11104 2416 11136
rect 2448 11104 2488 11136
rect 2520 11104 2560 11136
rect 2592 11104 2632 11136
rect 2664 11104 2704 11136
rect 2736 11104 2776 11136
rect 2808 11104 2848 11136
rect 2880 11104 2920 11136
rect 2952 11104 2992 11136
rect 3024 11104 3064 11136
rect 3096 11104 3136 11136
rect 3168 11104 3208 11136
rect 3240 11104 3280 11136
rect 3312 11104 3352 11136
rect 3384 11104 3424 11136
rect 3456 11104 3496 11136
rect 3528 11104 3568 11136
rect 3600 11104 3640 11136
rect 3672 11104 3712 11136
rect 3744 11104 3784 11136
rect 3816 11104 3856 11136
rect 3888 11104 3928 11136
rect 3960 11104 4000 11136
rect 0 11064 4000 11104
rect 0 11032 40 11064
rect 72 11032 112 11064
rect 144 11032 184 11064
rect 216 11032 256 11064
rect 288 11032 328 11064
rect 360 11032 400 11064
rect 432 11032 472 11064
rect 504 11032 544 11064
rect 576 11032 616 11064
rect 648 11032 688 11064
rect 720 11032 760 11064
rect 792 11032 832 11064
rect 864 11032 904 11064
rect 936 11032 976 11064
rect 1008 11032 1048 11064
rect 1080 11032 1120 11064
rect 1152 11032 1192 11064
rect 1224 11032 1264 11064
rect 1296 11032 1336 11064
rect 1368 11032 1408 11064
rect 1440 11032 1480 11064
rect 1512 11032 1552 11064
rect 1584 11032 1624 11064
rect 1656 11032 1696 11064
rect 1728 11032 1768 11064
rect 1800 11032 1840 11064
rect 1872 11032 1912 11064
rect 1944 11032 1984 11064
rect 2016 11032 2056 11064
rect 2088 11032 2128 11064
rect 2160 11032 2200 11064
rect 2232 11032 2272 11064
rect 2304 11032 2344 11064
rect 2376 11032 2416 11064
rect 2448 11032 2488 11064
rect 2520 11032 2560 11064
rect 2592 11032 2632 11064
rect 2664 11032 2704 11064
rect 2736 11032 2776 11064
rect 2808 11032 2848 11064
rect 2880 11032 2920 11064
rect 2952 11032 2992 11064
rect 3024 11032 3064 11064
rect 3096 11032 3136 11064
rect 3168 11032 3208 11064
rect 3240 11032 3280 11064
rect 3312 11032 3352 11064
rect 3384 11032 3424 11064
rect 3456 11032 3496 11064
rect 3528 11032 3568 11064
rect 3600 11032 3640 11064
rect 3672 11032 3712 11064
rect 3744 11032 3784 11064
rect 3816 11032 3856 11064
rect 3888 11032 3928 11064
rect 3960 11032 4000 11064
rect 0 10992 4000 11032
rect 0 10960 40 10992
rect 72 10960 112 10992
rect 144 10960 184 10992
rect 216 10960 256 10992
rect 288 10960 328 10992
rect 360 10960 400 10992
rect 432 10960 472 10992
rect 504 10960 544 10992
rect 576 10960 616 10992
rect 648 10960 688 10992
rect 720 10960 760 10992
rect 792 10960 832 10992
rect 864 10960 904 10992
rect 936 10960 976 10992
rect 1008 10960 1048 10992
rect 1080 10960 1120 10992
rect 1152 10960 1192 10992
rect 1224 10960 1264 10992
rect 1296 10960 1336 10992
rect 1368 10960 1408 10992
rect 1440 10960 1480 10992
rect 1512 10960 1552 10992
rect 1584 10960 1624 10992
rect 1656 10960 1696 10992
rect 1728 10960 1768 10992
rect 1800 10960 1840 10992
rect 1872 10960 1912 10992
rect 1944 10960 1984 10992
rect 2016 10960 2056 10992
rect 2088 10960 2128 10992
rect 2160 10960 2200 10992
rect 2232 10960 2272 10992
rect 2304 10960 2344 10992
rect 2376 10960 2416 10992
rect 2448 10960 2488 10992
rect 2520 10960 2560 10992
rect 2592 10960 2632 10992
rect 2664 10960 2704 10992
rect 2736 10960 2776 10992
rect 2808 10960 2848 10992
rect 2880 10960 2920 10992
rect 2952 10960 2992 10992
rect 3024 10960 3064 10992
rect 3096 10960 3136 10992
rect 3168 10960 3208 10992
rect 3240 10960 3280 10992
rect 3312 10960 3352 10992
rect 3384 10960 3424 10992
rect 3456 10960 3496 10992
rect 3528 10960 3568 10992
rect 3600 10960 3640 10992
rect 3672 10960 3712 10992
rect 3744 10960 3784 10992
rect 3816 10960 3856 10992
rect 3888 10960 3928 10992
rect 3960 10960 4000 10992
rect 0 10920 4000 10960
rect 0 10888 40 10920
rect 72 10888 112 10920
rect 144 10888 184 10920
rect 216 10888 256 10920
rect 288 10888 328 10920
rect 360 10888 400 10920
rect 432 10888 472 10920
rect 504 10888 544 10920
rect 576 10888 616 10920
rect 648 10888 688 10920
rect 720 10888 760 10920
rect 792 10888 832 10920
rect 864 10888 904 10920
rect 936 10888 976 10920
rect 1008 10888 1048 10920
rect 1080 10888 1120 10920
rect 1152 10888 1192 10920
rect 1224 10888 1264 10920
rect 1296 10888 1336 10920
rect 1368 10888 1408 10920
rect 1440 10888 1480 10920
rect 1512 10888 1552 10920
rect 1584 10888 1624 10920
rect 1656 10888 1696 10920
rect 1728 10888 1768 10920
rect 1800 10888 1840 10920
rect 1872 10888 1912 10920
rect 1944 10888 1984 10920
rect 2016 10888 2056 10920
rect 2088 10888 2128 10920
rect 2160 10888 2200 10920
rect 2232 10888 2272 10920
rect 2304 10888 2344 10920
rect 2376 10888 2416 10920
rect 2448 10888 2488 10920
rect 2520 10888 2560 10920
rect 2592 10888 2632 10920
rect 2664 10888 2704 10920
rect 2736 10888 2776 10920
rect 2808 10888 2848 10920
rect 2880 10888 2920 10920
rect 2952 10888 2992 10920
rect 3024 10888 3064 10920
rect 3096 10888 3136 10920
rect 3168 10888 3208 10920
rect 3240 10888 3280 10920
rect 3312 10888 3352 10920
rect 3384 10888 3424 10920
rect 3456 10888 3496 10920
rect 3528 10888 3568 10920
rect 3600 10888 3640 10920
rect 3672 10888 3712 10920
rect 3744 10888 3784 10920
rect 3816 10888 3856 10920
rect 3888 10888 3928 10920
rect 3960 10888 4000 10920
rect 0 10848 4000 10888
rect 0 10816 40 10848
rect 72 10816 112 10848
rect 144 10816 184 10848
rect 216 10816 256 10848
rect 288 10816 328 10848
rect 360 10816 400 10848
rect 432 10816 472 10848
rect 504 10816 544 10848
rect 576 10816 616 10848
rect 648 10816 688 10848
rect 720 10816 760 10848
rect 792 10816 832 10848
rect 864 10816 904 10848
rect 936 10816 976 10848
rect 1008 10816 1048 10848
rect 1080 10816 1120 10848
rect 1152 10816 1192 10848
rect 1224 10816 1264 10848
rect 1296 10816 1336 10848
rect 1368 10816 1408 10848
rect 1440 10816 1480 10848
rect 1512 10816 1552 10848
rect 1584 10816 1624 10848
rect 1656 10816 1696 10848
rect 1728 10816 1768 10848
rect 1800 10816 1840 10848
rect 1872 10816 1912 10848
rect 1944 10816 1984 10848
rect 2016 10816 2056 10848
rect 2088 10816 2128 10848
rect 2160 10816 2200 10848
rect 2232 10816 2272 10848
rect 2304 10816 2344 10848
rect 2376 10816 2416 10848
rect 2448 10816 2488 10848
rect 2520 10816 2560 10848
rect 2592 10816 2632 10848
rect 2664 10816 2704 10848
rect 2736 10816 2776 10848
rect 2808 10816 2848 10848
rect 2880 10816 2920 10848
rect 2952 10816 2992 10848
rect 3024 10816 3064 10848
rect 3096 10816 3136 10848
rect 3168 10816 3208 10848
rect 3240 10816 3280 10848
rect 3312 10816 3352 10848
rect 3384 10816 3424 10848
rect 3456 10816 3496 10848
rect 3528 10816 3568 10848
rect 3600 10816 3640 10848
rect 3672 10816 3712 10848
rect 3744 10816 3784 10848
rect 3816 10816 3856 10848
rect 3888 10816 3928 10848
rect 3960 10816 4000 10848
rect 0 10776 4000 10816
rect 0 10744 40 10776
rect 72 10744 112 10776
rect 144 10744 184 10776
rect 216 10744 256 10776
rect 288 10744 328 10776
rect 360 10744 400 10776
rect 432 10744 472 10776
rect 504 10744 544 10776
rect 576 10744 616 10776
rect 648 10744 688 10776
rect 720 10744 760 10776
rect 792 10744 832 10776
rect 864 10744 904 10776
rect 936 10744 976 10776
rect 1008 10744 1048 10776
rect 1080 10744 1120 10776
rect 1152 10744 1192 10776
rect 1224 10744 1264 10776
rect 1296 10744 1336 10776
rect 1368 10744 1408 10776
rect 1440 10744 1480 10776
rect 1512 10744 1552 10776
rect 1584 10744 1624 10776
rect 1656 10744 1696 10776
rect 1728 10744 1768 10776
rect 1800 10744 1840 10776
rect 1872 10744 1912 10776
rect 1944 10744 1984 10776
rect 2016 10744 2056 10776
rect 2088 10744 2128 10776
rect 2160 10744 2200 10776
rect 2232 10744 2272 10776
rect 2304 10744 2344 10776
rect 2376 10744 2416 10776
rect 2448 10744 2488 10776
rect 2520 10744 2560 10776
rect 2592 10744 2632 10776
rect 2664 10744 2704 10776
rect 2736 10744 2776 10776
rect 2808 10744 2848 10776
rect 2880 10744 2920 10776
rect 2952 10744 2992 10776
rect 3024 10744 3064 10776
rect 3096 10744 3136 10776
rect 3168 10744 3208 10776
rect 3240 10744 3280 10776
rect 3312 10744 3352 10776
rect 3384 10744 3424 10776
rect 3456 10744 3496 10776
rect 3528 10744 3568 10776
rect 3600 10744 3640 10776
rect 3672 10744 3712 10776
rect 3744 10744 3784 10776
rect 3816 10744 3856 10776
rect 3888 10744 3928 10776
rect 3960 10744 4000 10776
rect 0 10704 4000 10744
rect 0 10672 40 10704
rect 72 10672 112 10704
rect 144 10672 184 10704
rect 216 10672 256 10704
rect 288 10672 328 10704
rect 360 10672 400 10704
rect 432 10672 472 10704
rect 504 10672 544 10704
rect 576 10672 616 10704
rect 648 10672 688 10704
rect 720 10672 760 10704
rect 792 10672 832 10704
rect 864 10672 904 10704
rect 936 10672 976 10704
rect 1008 10672 1048 10704
rect 1080 10672 1120 10704
rect 1152 10672 1192 10704
rect 1224 10672 1264 10704
rect 1296 10672 1336 10704
rect 1368 10672 1408 10704
rect 1440 10672 1480 10704
rect 1512 10672 1552 10704
rect 1584 10672 1624 10704
rect 1656 10672 1696 10704
rect 1728 10672 1768 10704
rect 1800 10672 1840 10704
rect 1872 10672 1912 10704
rect 1944 10672 1984 10704
rect 2016 10672 2056 10704
rect 2088 10672 2128 10704
rect 2160 10672 2200 10704
rect 2232 10672 2272 10704
rect 2304 10672 2344 10704
rect 2376 10672 2416 10704
rect 2448 10672 2488 10704
rect 2520 10672 2560 10704
rect 2592 10672 2632 10704
rect 2664 10672 2704 10704
rect 2736 10672 2776 10704
rect 2808 10672 2848 10704
rect 2880 10672 2920 10704
rect 2952 10672 2992 10704
rect 3024 10672 3064 10704
rect 3096 10672 3136 10704
rect 3168 10672 3208 10704
rect 3240 10672 3280 10704
rect 3312 10672 3352 10704
rect 3384 10672 3424 10704
rect 3456 10672 3496 10704
rect 3528 10672 3568 10704
rect 3600 10672 3640 10704
rect 3672 10672 3712 10704
rect 3744 10672 3784 10704
rect 3816 10672 3856 10704
rect 3888 10672 3928 10704
rect 3960 10672 4000 10704
rect 0 10632 4000 10672
rect 0 10600 40 10632
rect 72 10600 112 10632
rect 144 10600 184 10632
rect 216 10600 256 10632
rect 288 10600 328 10632
rect 360 10600 400 10632
rect 432 10600 472 10632
rect 504 10600 544 10632
rect 576 10600 616 10632
rect 648 10600 688 10632
rect 720 10600 760 10632
rect 792 10600 832 10632
rect 864 10600 904 10632
rect 936 10600 976 10632
rect 1008 10600 1048 10632
rect 1080 10600 1120 10632
rect 1152 10600 1192 10632
rect 1224 10600 1264 10632
rect 1296 10600 1336 10632
rect 1368 10600 1408 10632
rect 1440 10600 1480 10632
rect 1512 10600 1552 10632
rect 1584 10600 1624 10632
rect 1656 10600 1696 10632
rect 1728 10600 1768 10632
rect 1800 10600 1840 10632
rect 1872 10600 1912 10632
rect 1944 10600 1984 10632
rect 2016 10600 2056 10632
rect 2088 10600 2128 10632
rect 2160 10600 2200 10632
rect 2232 10600 2272 10632
rect 2304 10600 2344 10632
rect 2376 10600 2416 10632
rect 2448 10600 2488 10632
rect 2520 10600 2560 10632
rect 2592 10600 2632 10632
rect 2664 10600 2704 10632
rect 2736 10600 2776 10632
rect 2808 10600 2848 10632
rect 2880 10600 2920 10632
rect 2952 10600 2992 10632
rect 3024 10600 3064 10632
rect 3096 10600 3136 10632
rect 3168 10600 3208 10632
rect 3240 10600 3280 10632
rect 3312 10600 3352 10632
rect 3384 10600 3424 10632
rect 3456 10600 3496 10632
rect 3528 10600 3568 10632
rect 3600 10600 3640 10632
rect 3672 10600 3712 10632
rect 3744 10600 3784 10632
rect 3816 10600 3856 10632
rect 3888 10600 3928 10632
rect 3960 10600 4000 10632
rect 0 10560 4000 10600
rect 0 10528 40 10560
rect 72 10528 112 10560
rect 144 10528 184 10560
rect 216 10528 256 10560
rect 288 10528 328 10560
rect 360 10528 400 10560
rect 432 10528 472 10560
rect 504 10528 544 10560
rect 576 10528 616 10560
rect 648 10528 688 10560
rect 720 10528 760 10560
rect 792 10528 832 10560
rect 864 10528 904 10560
rect 936 10528 976 10560
rect 1008 10528 1048 10560
rect 1080 10528 1120 10560
rect 1152 10528 1192 10560
rect 1224 10528 1264 10560
rect 1296 10528 1336 10560
rect 1368 10528 1408 10560
rect 1440 10528 1480 10560
rect 1512 10528 1552 10560
rect 1584 10528 1624 10560
rect 1656 10528 1696 10560
rect 1728 10528 1768 10560
rect 1800 10528 1840 10560
rect 1872 10528 1912 10560
rect 1944 10528 1984 10560
rect 2016 10528 2056 10560
rect 2088 10528 2128 10560
rect 2160 10528 2200 10560
rect 2232 10528 2272 10560
rect 2304 10528 2344 10560
rect 2376 10528 2416 10560
rect 2448 10528 2488 10560
rect 2520 10528 2560 10560
rect 2592 10528 2632 10560
rect 2664 10528 2704 10560
rect 2736 10528 2776 10560
rect 2808 10528 2848 10560
rect 2880 10528 2920 10560
rect 2952 10528 2992 10560
rect 3024 10528 3064 10560
rect 3096 10528 3136 10560
rect 3168 10528 3208 10560
rect 3240 10528 3280 10560
rect 3312 10528 3352 10560
rect 3384 10528 3424 10560
rect 3456 10528 3496 10560
rect 3528 10528 3568 10560
rect 3600 10528 3640 10560
rect 3672 10528 3712 10560
rect 3744 10528 3784 10560
rect 3816 10528 3856 10560
rect 3888 10528 3928 10560
rect 3960 10528 4000 10560
rect 0 10488 4000 10528
rect 0 10456 40 10488
rect 72 10456 112 10488
rect 144 10456 184 10488
rect 216 10456 256 10488
rect 288 10456 328 10488
rect 360 10456 400 10488
rect 432 10456 472 10488
rect 504 10456 544 10488
rect 576 10456 616 10488
rect 648 10456 688 10488
rect 720 10456 760 10488
rect 792 10456 832 10488
rect 864 10456 904 10488
rect 936 10456 976 10488
rect 1008 10456 1048 10488
rect 1080 10456 1120 10488
rect 1152 10456 1192 10488
rect 1224 10456 1264 10488
rect 1296 10456 1336 10488
rect 1368 10456 1408 10488
rect 1440 10456 1480 10488
rect 1512 10456 1552 10488
rect 1584 10456 1624 10488
rect 1656 10456 1696 10488
rect 1728 10456 1768 10488
rect 1800 10456 1840 10488
rect 1872 10456 1912 10488
rect 1944 10456 1984 10488
rect 2016 10456 2056 10488
rect 2088 10456 2128 10488
rect 2160 10456 2200 10488
rect 2232 10456 2272 10488
rect 2304 10456 2344 10488
rect 2376 10456 2416 10488
rect 2448 10456 2488 10488
rect 2520 10456 2560 10488
rect 2592 10456 2632 10488
rect 2664 10456 2704 10488
rect 2736 10456 2776 10488
rect 2808 10456 2848 10488
rect 2880 10456 2920 10488
rect 2952 10456 2992 10488
rect 3024 10456 3064 10488
rect 3096 10456 3136 10488
rect 3168 10456 3208 10488
rect 3240 10456 3280 10488
rect 3312 10456 3352 10488
rect 3384 10456 3424 10488
rect 3456 10456 3496 10488
rect 3528 10456 3568 10488
rect 3600 10456 3640 10488
rect 3672 10456 3712 10488
rect 3744 10456 3784 10488
rect 3816 10456 3856 10488
rect 3888 10456 3928 10488
rect 3960 10456 4000 10488
rect 0 10416 4000 10456
rect 0 10384 40 10416
rect 72 10384 112 10416
rect 144 10384 184 10416
rect 216 10384 256 10416
rect 288 10384 328 10416
rect 360 10384 400 10416
rect 432 10384 472 10416
rect 504 10384 544 10416
rect 576 10384 616 10416
rect 648 10384 688 10416
rect 720 10384 760 10416
rect 792 10384 832 10416
rect 864 10384 904 10416
rect 936 10384 976 10416
rect 1008 10384 1048 10416
rect 1080 10384 1120 10416
rect 1152 10384 1192 10416
rect 1224 10384 1264 10416
rect 1296 10384 1336 10416
rect 1368 10384 1408 10416
rect 1440 10384 1480 10416
rect 1512 10384 1552 10416
rect 1584 10384 1624 10416
rect 1656 10384 1696 10416
rect 1728 10384 1768 10416
rect 1800 10384 1840 10416
rect 1872 10384 1912 10416
rect 1944 10384 1984 10416
rect 2016 10384 2056 10416
rect 2088 10384 2128 10416
rect 2160 10384 2200 10416
rect 2232 10384 2272 10416
rect 2304 10384 2344 10416
rect 2376 10384 2416 10416
rect 2448 10384 2488 10416
rect 2520 10384 2560 10416
rect 2592 10384 2632 10416
rect 2664 10384 2704 10416
rect 2736 10384 2776 10416
rect 2808 10384 2848 10416
rect 2880 10384 2920 10416
rect 2952 10384 2992 10416
rect 3024 10384 3064 10416
rect 3096 10384 3136 10416
rect 3168 10384 3208 10416
rect 3240 10384 3280 10416
rect 3312 10384 3352 10416
rect 3384 10384 3424 10416
rect 3456 10384 3496 10416
rect 3528 10384 3568 10416
rect 3600 10384 3640 10416
rect 3672 10384 3712 10416
rect 3744 10384 3784 10416
rect 3816 10384 3856 10416
rect 3888 10384 3928 10416
rect 3960 10384 4000 10416
rect 0 10344 4000 10384
rect 0 10312 40 10344
rect 72 10312 112 10344
rect 144 10312 184 10344
rect 216 10312 256 10344
rect 288 10312 328 10344
rect 360 10312 400 10344
rect 432 10312 472 10344
rect 504 10312 544 10344
rect 576 10312 616 10344
rect 648 10312 688 10344
rect 720 10312 760 10344
rect 792 10312 832 10344
rect 864 10312 904 10344
rect 936 10312 976 10344
rect 1008 10312 1048 10344
rect 1080 10312 1120 10344
rect 1152 10312 1192 10344
rect 1224 10312 1264 10344
rect 1296 10312 1336 10344
rect 1368 10312 1408 10344
rect 1440 10312 1480 10344
rect 1512 10312 1552 10344
rect 1584 10312 1624 10344
rect 1656 10312 1696 10344
rect 1728 10312 1768 10344
rect 1800 10312 1840 10344
rect 1872 10312 1912 10344
rect 1944 10312 1984 10344
rect 2016 10312 2056 10344
rect 2088 10312 2128 10344
rect 2160 10312 2200 10344
rect 2232 10312 2272 10344
rect 2304 10312 2344 10344
rect 2376 10312 2416 10344
rect 2448 10312 2488 10344
rect 2520 10312 2560 10344
rect 2592 10312 2632 10344
rect 2664 10312 2704 10344
rect 2736 10312 2776 10344
rect 2808 10312 2848 10344
rect 2880 10312 2920 10344
rect 2952 10312 2992 10344
rect 3024 10312 3064 10344
rect 3096 10312 3136 10344
rect 3168 10312 3208 10344
rect 3240 10312 3280 10344
rect 3312 10312 3352 10344
rect 3384 10312 3424 10344
rect 3456 10312 3496 10344
rect 3528 10312 3568 10344
rect 3600 10312 3640 10344
rect 3672 10312 3712 10344
rect 3744 10312 3784 10344
rect 3816 10312 3856 10344
rect 3888 10312 3928 10344
rect 3960 10312 4000 10344
rect 0 10272 4000 10312
rect 0 10240 40 10272
rect 72 10240 112 10272
rect 144 10240 184 10272
rect 216 10240 256 10272
rect 288 10240 328 10272
rect 360 10240 400 10272
rect 432 10240 472 10272
rect 504 10240 544 10272
rect 576 10240 616 10272
rect 648 10240 688 10272
rect 720 10240 760 10272
rect 792 10240 832 10272
rect 864 10240 904 10272
rect 936 10240 976 10272
rect 1008 10240 1048 10272
rect 1080 10240 1120 10272
rect 1152 10240 1192 10272
rect 1224 10240 1264 10272
rect 1296 10240 1336 10272
rect 1368 10240 1408 10272
rect 1440 10240 1480 10272
rect 1512 10240 1552 10272
rect 1584 10240 1624 10272
rect 1656 10240 1696 10272
rect 1728 10240 1768 10272
rect 1800 10240 1840 10272
rect 1872 10240 1912 10272
rect 1944 10240 1984 10272
rect 2016 10240 2056 10272
rect 2088 10240 2128 10272
rect 2160 10240 2200 10272
rect 2232 10240 2272 10272
rect 2304 10240 2344 10272
rect 2376 10240 2416 10272
rect 2448 10240 2488 10272
rect 2520 10240 2560 10272
rect 2592 10240 2632 10272
rect 2664 10240 2704 10272
rect 2736 10240 2776 10272
rect 2808 10240 2848 10272
rect 2880 10240 2920 10272
rect 2952 10240 2992 10272
rect 3024 10240 3064 10272
rect 3096 10240 3136 10272
rect 3168 10240 3208 10272
rect 3240 10240 3280 10272
rect 3312 10240 3352 10272
rect 3384 10240 3424 10272
rect 3456 10240 3496 10272
rect 3528 10240 3568 10272
rect 3600 10240 3640 10272
rect 3672 10240 3712 10272
rect 3744 10240 3784 10272
rect 3816 10240 3856 10272
rect 3888 10240 3928 10272
rect 3960 10240 4000 10272
rect 0 10200 4000 10240
rect 0 10168 40 10200
rect 72 10168 112 10200
rect 144 10168 184 10200
rect 216 10168 256 10200
rect 288 10168 328 10200
rect 360 10168 400 10200
rect 432 10168 472 10200
rect 504 10168 544 10200
rect 576 10168 616 10200
rect 648 10168 688 10200
rect 720 10168 760 10200
rect 792 10168 832 10200
rect 864 10168 904 10200
rect 936 10168 976 10200
rect 1008 10168 1048 10200
rect 1080 10168 1120 10200
rect 1152 10168 1192 10200
rect 1224 10168 1264 10200
rect 1296 10168 1336 10200
rect 1368 10168 1408 10200
rect 1440 10168 1480 10200
rect 1512 10168 1552 10200
rect 1584 10168 1624 10200
rect 1656 10168 1696 10200
rect 1728 10168 1768 10200
rect 1800 10168 1840 10200
rect 1872 10168 1912 10200
rect 1944 10168 1984 10200
rect 2016 10168 2056 10200
rect 2088 10168 2128 10200
rect 2160 10168 2200 10200
rect 2232 10168 2272 10200
rect 2304 10168 2344 10200
rect 2376 10168 2416 10200
rect 2448 10168 2488 10200
rect 2520 10168 2560 10200
rect 2592 10168 2632 10200
rect 2664 10168 2704 10200
rect 2736 10168 2776 10200
rect 2808 10168 2848 10200
rect 2880 10168 2920 10200
rect 2952 10168 2992 10200
rect 3024 10168 3064 10200
rect 3096 10168 3136 10200
rect 3168 10168 3208 10200
rect 3240 10168 3280 10200
rect 3312 10168 3352 10200
rect 3384 10168 3424 10200
rect 3456 10168 3496 10200
rect 3528 10168 3568 10200
rect 3600 10168 3640 10200
rect 3672 10168 3712 10200
rect 3744 10168 3784 10200
rect 3816 10168 3856 10200
rect 3888 10168 3928 10200
rect 3960 10168 4000 10200
rect 0 10128 4000 10168
rect 0 10096 40 10128
rect 72 10096 112 10128
rect 144 10096 184 10128
rect 216 10096 256 10128
rect 288 10096 328 10128
rect 360 10096 400 10128
rect 432 10096 472 10128
rect 504 10096 544 10128
rect 576 10096 616 10128
rect 648 10096 688 10128
rect 720 10096 760 10128
rect 792 10096 832 10128
rect 864 10096 904 10128
rect 936 10096 976 10128
rect 1008 10096 1048 10128
rect 1080 10096 1120 10128
rect 1152 10096 1192 10128
rect 1224 10096 1264 10128
rect 1296 10096 1336 10128
rect 1368 10096 1408 10128
rect 1440 10096 1480 10128
rect 1512 10096 1552 10128
rect 1584 10096 1624 10128
rect 1656 10096 1696 10128
rect 1728 10096 1768 10128
rect 1800 10096 1840 10128
rect 1872 10096 1912 10128
rect 1944 10096 1984 10128
rect 2016 10096 2056 10128
rect 2088 10096 2128 10128
rect 2160 10096 2200 10128
rect 2232 10096 2272 10128
rect 2304 10096 2344 10128
rect 2376 10096 2416 10128
rect 2448 10096 2488 10128
rect 2520 10096 2560 10128
rect 2592 10096 2632 10128
rect 2664 10096 2704 10128
rect 2736 10096 2776 10128
rect 2808 10096 2848 10128
rect 2880 10096 2920 10128
rect 2952 10096 2992 10128
rect 3024 10096 3064 10128
rect 3096 10096 3136 10128
rect 3168 10096 3208 10128
rect 3240 10096 3280 10128
rect 3312 10096 3352 10128
rect 3384 10096 3424 10128
rect 3456 10096 3496 10128
rect 3528 10096 3568 10128
rect 3600 10096 3640 10128
rect 3672 10096 3712 10128
rect 3744 10096 3784 10128
rect 3816 10096 3856 10128
rect 3888 10096 3928 10128
rect 3960 10096 4000 10128
rect 0 10056 4000 10096
rect 0 10024 40 10056
rect 72 10024 112 10056
rect 144 10024 184 10056
rect 216 10024 256 10056
rect 288 10024 328 10056
rect 360 10024 400 10056
rect 432 10024 472 10056
rect 504 10024 544 10056
rect 576 10024 616 10056
rect 648 10024 688 10056
rect 720 10024 760 10056
rect 792 10024 832 10056
rect 864 10024 904 10056
rect 936 10024 976 10056
rect 1008 10024 1048 10056
rect 1080 10024 1120 10056
rect 1152 10024 1192 10056
rect 1224 10024 1264 10056
rect 1296 10024 1336 10056
rect 1368 10024 1408 10056
rect 1440 10024 1480 10056
rect 1512 10024 1552 10056
rect 1584 10024 1624 10056
rect 1656 10024 1696 10056
rect 1728 10024 1768 10056
rect 1800 10024 1840 10056
rect 1872 10024 1912 10056
rect 1944 10024 1984 10056
rect 2016 10024 2056 10056
rect 2088 10024 2128 10056
rect 2160 10024 2200 10056
rect 2232 10024 2272 10056
rect 2304 10024 2344 10056
rect 2376 10024 2416 10056
rect 2448 10024 2488 10056
rect 2520 10024 2560 10056
rect 2592 10024 2632 10056
rect 2664 10024 2704 10056
rect 2736 10024 2776 10056
rect 2808 10024 2848 10056
rect 2880 10024 2920 10056
rect 2952 10024 2992 10056
rect 3024 10024 3064 10056
rect 3096 10024 3136 10056
rect 3168 10024 3208 10056
rect 3240 10024 3280 10056
rect 3312 10024 3352 10056
rect 3384 10024 3424 10056
rect 3456 10024 3496 10056
rect 3528 10024 3568 10056
rect 3600 10024 3640 10056
rect 3672 10024 3712 10056
rect 3744 10024 3784 10056
rect 3816 10024 3856 10056
rect 3888 10024 3928 10056
rect 3960 10024 4000 10056
rect 0 9984 4000 10024
rect 0 9952 40 9984
rect 72 9952 112 9984
rect 144 9952 184 9984
rect 216 9952 256 9984
rect 288 9952 328 9984
rect 360 9952 400 9984
rect 432 9952 472 9984
rect 504 9952 544 9984
rect 576 9952 616 9984
rect 648 9952 688 9984
rect 720 9952 760 9984
rect 792 9952 832 9984
rect 864 9952 904 9984
rect 936 9952 976 9984
rect 1008 9952 1048 9984
rect 1080 9952 1120 9984
rect 1152 9952 1192 9984
rect 1224 9952 1264 9984
rect 1296 9952 1336 9984
rect 1368 9952 1408 9984
rect 1440 9952 1480 9984
rect 1512 9952 1552 9984
rect 1584 9952 1624 9984
rect 1656 9952 1696 9984
rect 1728 9952 1768 9984
rect 1800 9952 1840 9984
rect 1872 9952 1912 9984
rect 1944 9952 1984 9984
rect 2016 9952 2056 9984
rect 2088 9952 2128 9984
rect 2160 9952 2200 9984
rect 2232 9952 2272 9984
rect 2304 9952 2344 9984
rect 2376 9952 2416 9984
rect 2448 9952 2488 9984
rect 2520 9952 2560 9984
rect 2592 9952 2632 9984
rect 2664 9952 2704 9984
rect 2736 9952 2776 9984
rect 2808 9952 2848 9984
rect 2880 9952 2920 9984
rect 2952 9952 2992 9984
rect 3024 9952 3064 9984
rect 3096 9952 3136 9984
rect 3168 9952 3208 9984
rect 3240 9952 3280 9984
rect 3312 9952 3352 9984
rect 3384 9952 3424 9984
rect 3456 9952 3496 9984
rect 3528 9952 3568 9984
rect 3600 9952 3640 9984
rect 3672 9952 3712 9984
rect 3744 9952 3784 9984
rect 3816 9952 3856 9984
rect 3888 9952 3928 9984
rect 3960 9952 4000 9984
rect 0 9912 4000 9952
rect 0 9880 40 9912
rect 72 9880 112 9912
rect 144 9880 184 9912
rect 216 9880 256 9912
rect 288 9880 328 9912
rect 360 9880 400 9912
rect 432 9880 472 9912
rect 504 9880 544 9912
rect 576 9880 616 9912
rect 648 9880 688 9912
rect 720 9880 760 9912
rect 792 9880 832 9912
rect 864 9880 904 9912
rect 936 9880 976 9912
rect 1008 9880 1048 9912
rect 1080 9880 1120 9912
rect 1152 9880 1192 9912
rect 1224 9880 1264 9912
rect 1296 9880 1336 9912
rect 1368 9880 1408 9912
rect 1440 9880 1480 9912
rect 1512 9880 1552 9912
rect 1584 9880 1624 9912
rect 1656 9880 1696 9912
rect 1728 9880 1768 9912
rect 1800 9880 1840 9912
rect 1872 9880 1912 9912
rect 1944 9880 1984 9912
rect 2016 9880 2056 9912
rect 2088 9880 2128 9912
rect 2160 9880 2200 9912
rect 2232 9880 2272 9912
rect 2304 9880 2344 9912
rect 2376 9880 2416 9912
rect 2448 9880 2488 9912
rect 2520 9880 2560 9912
rect 2592 9880 2632 9912
rect 2664 9880 2704 9912
rect 2736 9880 2776 9912
rect 2808 9880 2848 9912
rect 2880 9880 2920 9912
rect 2952 9880 2992 9912
rect 3024 9880 3064 9912
rect 3096 9880 3136 9912
rect 3168 9880 3208 9912
rect 3240 9880 3280 9912
rect 3312 9880 3352 9912
rect 3384 9880 3424 9912
rect 3456 9880 3496 9912
rect 3528 9880 3568 9912
rect 3600 9880 3640 9912
rect 3672 9880 3712 9912
rect 3744 9880 3784 9912
rect 3816 9880 3856 9912
rect 3888 9880 3928 9912
rect 3960 9880 4000 9912
rect 0 9840 4000 9880
rect 0 9808 40 9840
rect 72 9808 112 9840
rect 144 9808 184 9840
rect 216 9808 256 9840
rect 288 9808 328 9840
rect 360 9808 400 9840
rect 432 9808 472 9840
rect 504 9808 544 9840
rect 576 9808 616 9840
rect 648 9808 688 9840
rect 720 9808 760 9840
rect 792 9808 832 9840
rect 864 9808 904 9840
rect 936 9808 976 9840
rect 1008 9808 1048 9840
rect 1080 9808 1120 9840
rect 1152 9808 1192 9840
rect 1224 9808 1264 9840
rect 1296 9808 1336 9840
rect 1368 9808 1408 9840
rect 1440 9808 1480 9840
rect 1512 9808 1552 9840
rect 1584 9808 1624 9840
rect 1656 9808 1696 9840
rect 1728 9808 1768 9840
rect 1800 9808 1840 9840
rect 1872 9808 1912 9840
rect 1944 9808 1984 9840
rect 2016 9808 2056 9840
rect 2088 9808 2128 9840
rect 2160 9808 2200 9840
rect 2232 9808 2272 9840
rect 2304 9808 2344 9840
rect 2376 9808 2416 9840
rect 2448 9808 2488 9840
rect 2520 9808 2560 9840
rect 2592 9808 2632 9840
rect 2664 9808 2704 9840
rect 2736 9808 2776 9840
rect 2808 9808 2848 9840
rect 2880 9808 2920 9840
rect 2952 9808 2992 9840
rect 3024 9808 3064 9840
rect 3096 9808 3136 9840
rect 3168 9808 3208 9840
rect 3240 9808 3280 9840
rect 3312 9808 3352 9840
rect 3384 9808 3424 9840
rect 3456 9808 3496 9840
rect 3528 9808 3568 9840
rect 3600 9808 3640 9840
rect 3672 9808 3712 9840
rect 3744 9808 3784 9840
rect 3816 9808 3856 9840
rect 3888 9808 3928 9840
rect 3960 9808 4000 9840
rect 0 9768 4000 9808
rect 0 9736 40 9768
rect 72 9736 112 9768
rect 144 9736 184 9768
rect 216 9736 256 9768
rect 288 9736 328 9768
rect 360 9736 400 9768
rect 432 9736 472 9768
rect 504 9736 544 9768
rect 576 9736 616 9768
rect 648 9736 688 9768
rect 720 9736 760 9768
rect 792 9736 832 9768
rect 864 9736 904 9768
rect 936 9736 976 9768
rect 1008 9736 1048 9768
rect 1080 9736 1120 9768
rect 1152 9736 1192 9768
rect 1224 9736 1264 9768
rect 1296 9736 1336 9768
rect 1368 9736 1408 9768
rect 1440 9736 1480 9768
rect 1512 9736 1552 9768
rect 1584 9736 1624 9768
rect 1656 9736 1696 9768
rect 1728 9736 1768 9768
rect 1800 9736 1840 9768
rect 1872 9736 1912 9768
rect 1944 9736 1984 9768
rect 2016 9736 2056 9768
rect 2088 9736 2128 9768
rect 2160 9736 2200 9768
rect 2232 9736 2272 9768
rect 2304 9736 2344 9768
rect 2376 9736 2416 9768
rect 2448 9736 2488 9768
rect 2520 9736 2560 9768
rect 2592 9736 2632 9768
rect 2664 9736 2704 9768
rect 2736 9736 2776 9768
rect 2808 9736 2848 9768
rect 2880 9736 2920 9768
rect 2952 9736 2992 9768
rect 3024 9736 3064 9768
rect 3096 9736 3136 9768
rect 3168 9736 3208 9768
rect 3240 9736 3280 9768
rect 3312 9736 3352 9768
rect 3384 9736 3424 9768
rect 3456 9736 3496 9768
rect 3528 9736 3568 9768
rect 3600 9736 3640 9768
rect 3672 9736 3712 9768
rect 3744 9736 3784 9768
rect 3816 9736 3856 9768
rect 3888 9736 3928 9768
rect 3960 9736 4000 9768
rect 0 9696 4000 9736
rect 0 9664 40 9696
rect 72 9664 112 9696
rect 144 9664 184 9696
rect 216 9664 256 9696
rect 288 9664 328 9696
rect 360 9664 400 9696
rect 432 9664 472 9696
rect 504 9664 544 9696
rect 576 9664 616 9696
rect 648 9664 688 9696
rect 720 9664 760 9696
rect 792 9664 832 9696
rect 864 9664 904 9696
rect 936 9664 976 9696
rect 1008 9664 1048 9696
rect 1080 9664 1120 9696
rect 1152 9664 1192 9696
rect 1224 9664 1264 9696
rect 1296 9664 1336 9696
rect 1368 9664 1408 9696
rect 1440 9664 1480 9696
rect 1512 9664 1552 9696
rect 1584 9664 1624 9696
rect 1656 9664 1696 9696
rect 1728 9664 1768 9696
rect 1800 9664 1840 9696
rect 1872 9664 1912 9696
rect 1944 9664 1984 9696
rect 2016 9664 2056 9696
rect 2088 9664 2128 9696
rect 2160 9664 2200 9696
rect 2232 9664 2272 9696
rect 2304 9664 2344 9696
rect 2376 9664 2416 9696
rect 2448 9664 2488 9696
rect 2520 9664 2560 9696
rect 2592 9664 2632 9696
rect 2664 9664 2704 9696
rect 2736 9664 2776 9696
rect 2808 9664 2848 9696
rect 2880 9664 2920 9696
rect 2952 9664 2992 9696
rect 3024 9664 3064 9696
rect 3096 9664 3136 9696
rect 3168 9664 3208 9696
rect 3240 9664 3280 9696
rect 3312 9664 3352 9696
rect 3384 9664 3424 9696
rect 3456 9664 3496 9696
rect 3528 9664 3568 9696
rect 3600 9664 3640 9696
rect 3672 9664 3712 9696
rect 3744 9664 3784 9696
rect 3816 9664 3856 9696
rect 3888 9664 3928 9696
rect 3960 9664 4000 9696
rect 0 9624 4000 9664
rect 0 9592 40 9624
rect 72 9592 112 9624
rect 144 9592 184 9624
rect 216 9592 256 9624
rect 288 9592 328 9624
rect 360 9592 400 9624
rect 432 9592 472 9624
rect 504 9592 544 9624
rect 576 9592 616 9624
rect 648 9592 688 9624
rect 720 9592 760 9624
rect 792 9592 832 9624
rect 864 9592 904 9624
rect 936 9592 976 9624
rect 1008 9592 1048 9624
rect 1080 9592 1120 9624
rect 1152 9592 1192 9624
rect 1224 9592 1264 9624
rect 1296 9592 1336 9624
rect 1368 9592 1408 9624
rect 1440 9592 1480 9624
rect 1512 9592 1552 9624
rect 1584 9592 1624 9624
rect 1656 9592 1696 9624
rect 1728 9592 1768 9624
rect 1800 9592 1840 9624
rect 1872 9592 1912 9624
rect 1944 9592 1984 9624
rect 2016 9592 2056 9624
rect 2088 9592 2128 9624
rect 2160 9592 2200 9624
rect 2232 9592 2272 9624
rect 2304 9592 2344 9624
rect 2376 9592 2416 9624
rect 2448 9592 2488 9624
rect 2520 9592 2560 9624
rect 2592 9592 2632 9624
rect 2664 9592 2704 9624
rect 2736 9592 2776 9624
rect 2808 9592 2848 9624
rect 2880 9592 2920 9624
rect 2952 9592 2992 9624
rect 3024 9592 3064 9624
rect 3096 9592 3136 9624
rect 3168 9592 3208 9624
rect 3240 9592 3280 9624
rect 3312 9592 3352 9624
rect 3384 9592 3424 9624
rect 3456 9592 3496 9624
rect 3528 9592 3568 9624
rect 3600 9592 3640 9624
rect 3672 9592 3712 9624
rect 3744 9592 3784 9624
rect 3816 9592 3856 9624
rect 3888 9592 3928 9624
rect 3960 9592 4000 9624
rect 0 9552 4000 9592
rect 0 9520 40 9552
rect 72 9520 112 9552
rect 144 9520 184 9552
rect 216 9520 256 9552
rect 288 9520 328 9552
rect 360 9520 400 9552
rect 432 9520 472 9552
rect 504 9520 544 9552
rect 576 9520 616 9552
rect 648 9520 688 9552
rect 720 9520 760 9552
rect 792 9520 832 9552
rect 864 9520 904 9552
rect 936 9520 976 9552
rect 1008 9520 1048 9552
rect 1080 9520 1120 9552
rect 1152 9520 1192 9552
rect 1224 9520 1264 9552
rect 1296 9520 1336 9552
rect 1368 9520 1408 9552
rect 1440 9520 1480 9552
rect 1512 9520 1552 9552
rect 1584 9520 1624 9552
rect 1656 9520 1696 9552
rect 1728 9520 1768 9552
rect 1800 9520 1840 9552
rect 1872 9520 1912 9552
rect 1944 9520 1984 9552
rect 2016 9520 2056 9552
rect 2088 9520 2128 9552
rect 2160 9520 2200 9552
rect 2232 9520 2272 9552
rect 2304 9520 2344 9552
rect 2376 9520 2416 9552
rect 2448 9520 2488 9552
rect 2520 9520 2560 9552
rect 2592 9520 2632 9552
rect 2664 9520 2704 9552
rect 2736 9520 2776 9552
rect 2808 9520 2848 9552
rect 2880 9520 2920 9552
rect 2952 9520 2992 9552
rect 3024 9520 3064 9552
rect 3096 9520 3136 9552
rect 3168 9520 3208 9552
rect 3240 9520 3280 9552
rect 3312 9520 3352 9552
rect 3384 9520 3424 9552
rect 3456 9520 3496 9552
rect 3528 9520 3568 9552
rect 3600 9520 3640 9552
rect 3672 9520 3712 9552
rect 3744 9520 3784 9552
rect 3816 9520 3856 9552
rect 3888 9520 3928 9552
rect 3960 9520 4000 9552
rect 0 9480 4000 9520
rect 0 9448 40 9480
rect 72 9448 112 9480
rect 144 9448 184 9480
rect 216 9448 256 9480
rect 288 9448 328 9480
rect 360 9448 400 9480
rect 432 9448 472 9480
rect 504 9448 544 9480
rect 576 9448 616 9480
rect 648 9448 688 9480
rect 720 9448 760 9480
rect 792 9448 832 9480
rect 864 9448 904 9480
rect 936 9448 976 9480
rect 1008 9448 1048 9480
rect 1080 9448 1120 9480
rect 1152 9448 1192 9480
rect 1224 9448 1264 9480
rect 1296 9448 1336 9480
rect 1368 9448 1408 9480
rect 1440 9448 1480 9480
rect 1512 9448 1552 9480
rect 1584 9448 1624 9480
rect 1656 9448 1696 9480
rect 1728 9448 1768 9480
rect 1800 9448 1840 9480
rect 1872 9448 1912 9480
rect 1944 9448 1984 9480
rect 2016 9448 2056 9480
rect 2088 9448 2128 9480
rect 2160 9448 2200 9480
rect 2232 9448 2272 9480
rect 2304 9448 2344 9480
rect 2376 9448 2416 9480
rect 2448 9448 2488 9480
rect 2520 9448 2560 9480
rect 2592 9448 2632 9480
rect 2664 9448 2704 9480
rect 2736 9448 2776 9480
rect 2808 9448 2848 9480
rect 2880 9448 2920 9480
rect 2952 9448 2992 9480
rect 3024 9448 3064 9480
rect 3096 9448 3136 9480
rect 3168 9448 3208 9480
rect 3240 9448 3280 9480
rect 3312 9448 3352 9480
rect 3384 9448 3424 9480
rect 3456 9448 3496 9480
rect 3528 9448 3568 9480
rect 3600 9448 3640 9480
rect 3672 9448 3712 9480
rect 3744 9448 3784 9480
rect 3816 9448 3856 9480
rect 3888 9448 3928 9480
rect 3960 9448 4000 9480
rect 0 9408 4000 9448
rect 0 9376 40 9408
rect 72 9376 112 9408
rect 144 9376 184 9408
rect 216 9376 256 9408
rect 288 9376 328 9408
rect 360 9376 400 9408
rect 432 9376 472 9408
rect 504 9376 544 9408
rect 576 9376 616 9408
rect 648 9376 688 9408
rect 720 9376 760 9408
rect 792 9376 832 9408
rect 864 9376 904 9408
rect 936 9376 976 9408
rect 1008 9376 1048 9408
rect 1080 9376 1120 9408
rect 1152 9376 1192 9408
rect 1224 9376 1264 9408
rect 1296 9376 1336 9408
rect 1368 9376 1408 9408
rect 1440 9376 1480 9408
rect 1512 9376 1552 9408
rect 1584 9376 1624 9408
rect 1656 9376 1696 9408
rect 1728 9376 1768 9408
rect 1800 9376 1840 9408
rect 1872 9376 1912 9408
rect 1944 9376 1984 9408
rect 2016 9376 2056 9408
rect 2088 9376 2128 9408
rect 2160 9376 2200 9408
rect 2232 9376 2272 9408
rect 2304 9376 2344 9408
rect 2376 9376 2416 9408
rect 2448 9376 2488 9408
rect 2520 9376 2560 9408
rect 2592 9376 2632 9408
rect 2664 9376 2704 9408
rect 2736 9376 2776 9408
rect 2808 9376 2848 9408
rect 2880 9376 2920 9408
rect 2952 9376 2992 9408
rect 3024 9376 3064 9408
rect 3096 9376 3136 9408
rect 3168 9376 3208 9408
rect 3240 9376 3280 9408
rect 3312 9376 3352 9408
rect 3384 9376 3424 9408
rect 3456 9376 3496 9408
rect 3528 9376 3568 9408
rect 3600 9376 3640 9408
rect 3672 9376 3712 9408
rect 3744 9376 3784 9408
rect 3816 9376 3856 9408
rect 3888 9376 3928 9408
rect 3960 9376 4000 9408
rect 0 9336 4000 9376
rect 0 9304 40 9336
rect 72 9304 112 9336
rect 144 9304 184 9336
rect 216 9304 256 9336
rect 288 9304 328 9336
rect 360 9304 400 9336
rect 432 9304 472 9336
rect 504 9304 544 9336
rect 576 9304 616 9336
rect 648 9304 688 9336
rect 720 9304 760 9336
rect 792 9304 832 9336
rect 864 9304 904 9336
rect 936 9304 976 9336
rect 1008 9304 1048 9336
rect 1080 9304 1120 9336
rect 1152 9304 1192 9336
rect 1224 9304 1264 9336
rect 1296 9304 1336 9336
rect 1368 9304 1408 9336
rect 1440 9304 1480 9336
rect 1512 9304 1552 9336
rect 1584 9304 1624 9336
rect 1656 9304 1696 9336
rect 1728 9304 1768 9336
rect 1800 9304 1840 9336
rect 1872 9304 1912 9336
rect 1944 9304 1984 9336
rect 2016 9304 2056 9336
rect 2088 9304 2128 9336
rect 2160 9304 2200 9336
rect 2232 9304 2272 9336
rect 2304 9304 2344 9336
rect 2376 9304 2416 9336
rect 2448 9304 2488 9336
rect 2520 9304 2560 9336
rect 2592 9304 2632 9336
rect 2664 9304 2704 9336
rect 2736 9304 2776 9336
rect 2808 9304 2848 9336
rect 2880 9304 2920 9336
rect 2952 9304 2992 9336
rect 3024 9304 3064 9336
rect 3096 9304 3136 9336
rect 3168 9304 3208 9336
rect 3240 9304 3280 9336
rect 3312 9304 3352 9336
rect 3384 9304 3424 9336
rect 3456 9304 3496 9336
rect 3528 9304 3568 9336
rect 3600 9304 3640 9336
rect 3672 9304 3712 9336
rect 3744 9304 3784 9336
rect 3816 9304 3856 9336
rect 3888 9304 3928 9336
rect 3960 9304 4000 9336
rect 0 9264 4000 9304
rect 0 9232 40 9264
rect 72 9232 112 9264
rect 144 9232 184 9264
rect 216 9232 256 9264
rect 288 9232 328 9264
rect 360 9232 400 9264
rect 432 9232 472 9264
rect 504 9232 544 9264
rect 576 9232 616 9264
rect 648 9232 688 9264
rect 720 9232 760 9264
rect 792 9232 832 9264
rect 864 9232 904 9264
rect 936 9232 976 9264
rect 1008 9232 1048 9264
rect 1080 9232 1120 9264
rect 1152 9232 1192 9264
rect 1224 9232 1264 9264
rect 1296 9232 1336 9264
rect 1368 9232 1408 9264
rect 1440 9232 1480 9264
rect 1512 9232 1552 9264
rect 1584 9232 1624 9264
rect 1656 9232 1696 9264
rect 1728 9232 1768 9264
rect 1800 9232 1840 9264
rect 1872 9232 1912 9264
rect 1944 9232 1984 9264
rect 2016 9232 2056 9264
rect 2088 9232 2128 9264
rect 2160 9232 2200 9264
rect 2232 9232 2272 9264
rect 2304 9232 2344 9264
rect 2376 9232 2416 9264
rect 2448 9232 2488 9264
rect 2520 9232 2560 9264
rect 2592 9232 2632 9264
rect 2664 9232 2704 9264
rect 2736 9232 2776 9264
rect 2808 9232 2848 9264
rect 2880 9232 2920 9264
rect 2952 9232 2992 9264
rect 3024 9232 3064 9264
rect 3096 9232 3136 9264
rect 3168 9232 3208 9264
rect 3240 9232 3280 9264
rect 3312 9232 3352 9264
rect 3384 9232 3424 9264
rect 3456 9232 3496 9264
rect 3528 9232 3568 9264
rect 3600 9232 3640 9264
rect 3672 9232 3712 9264
rect 3744 9232 3784 9264
rect 3816 9232 3856 9264
rect 3888 9232 3928 9264
rect 3960 9232 4000 9264
rect 0 9192 4000 9232
rect 0 9160 40 9192
rect 72 9160 112 9192
rect 144 9160 184 9192
rect 216 9160 256 9192
rect 288 9160 328 9192
rect 360 9160 400 9192
rect 432 9160 472 9192
rect 504 9160 544 9192
rect 576 9160 616 9192
rect 648 9160 688 9192
rect 720 9160 760 9192
rect 792 9160 832 9192
rect 864 9160 904 9192
rect 936 9160 976 9192
rect 1008 9160 1048 9192
rect 1080 9160 1120 9192
rect 1152 9160 1192 9192
rect 1224 9160 1264 9192
rect 1296 9160 1336 9192
rect 1368 9160 1408 9192
rect 1440 9160 1480 9192
rect 1512 9160 1552 9192
rect 1584 9160 1624 9192
rect 1656 9160 1696 9192
rect 1728 9160 1768 9192
rect 1800 9160 1840 9192
rect 1872 9160 1912 9192
rect 1944 9160 1984 9192
rect 2016 9160 2056 9192
rect 2088 9160 2128 9192
rect 2160 9160 2200 9192
rect 2232 9160 2272 9192
rect 2304 9160 2344 9192
rect 2376 9160 2416 9192
rect 2448 9160 2488 9192
rect 2520 9160 2560 9192
rect 2592 9160 2632 9192
rect 2664 9160 2704 9192
rect 2736 9160 2776 9192
rect 2808 9160 2848 9192
rect 2880 9160 2920 9192
rect 2952 9160 2992 9192
rect 3024 9160 3064 9192
rect 3096 9160 3136 9192
rect 3168 9160 3208 9192
rect 3240 9160 3280 9192
rect 3312 9160 3352 9192
rect 3384 9160 3424 9192
rect 3456 9160 3496 9192
rect 3528 9160 3568 9192
rect 3600 9160 3640 9192
rect 3672 9160 3712 9192
rect 3744 9160 3784 9192
rect 3816 9160 3856 9192
rect 3888 9160 3928 9192
rect 3960 9160 4000 9192
rect 0 9120 4000 9160
rect 0 9088 40 9120
rect 72 9088 112 9120
rect 144 9088 184 9120
rect 216 9088 256 9120
rect 288 9088 328 9120
rect 360 9088 400 9120
rect 432 9088 472 9120
rect 504 9088 544 9120
rect 576 9088 616 9120
rect 648 9088 688 9120
rect 720 9088 760 9120
rect 792 9088 832 9120
rect 864 9088 904 9120
rect 936 9088 976 9120
rect 1008 9088 1048 9120
rect 1080 9088 1120 9120
rect 1152 9088 1192 9120
rect 1224 9088 1264 9120
rect 1296 9088 1336 9120
rect 1368 9088 1408 9120
rect 1440 9088 1480 9120
rect 1512 9088 1552 9120
rect 1584 9088 1624 9120
rect 1656 9088 1696 9120
rect 1728 9088 1768 9120
rect 1800 9088 1840 9120
rect 1872 9088 1912 9120
rect 1944 9088 1984 9120
rect 2016 9088 2056 9120
rect 2088 9088 2128 9120
rect 2160 9088 2200 9120
rect 2232 9088 2272 9120
rect 2304 9088 2344 9120
rect 2376 9088 2416 9120
rect 2448 9088 2488 9120
rect 2520 9088 2560 9120
rect 2592 9088 2632 9120
rect 2664 9088 2704 9120
rect 2736 9088 2776 9120
rect 2808 9088 2848 9120
rect 2880 9088 2920 9120
rect 2952 9088 2992 9120
rect 3024 9088 3064 9120
rect 3096 9088 3136 9120
rect 3168 9088 3208 9120
rect 3240 9088 3280 9120
rect 3312 9088 3352 9120
rect 3384 9088 3424 9120
rect 3456 9088 3496 9120
rect 3528 9088 3568 9120
rect 3600 9088 3640 9120
rect 3672 9088 3712 9120
rect 3744 9088 3784 9120
rect 3816 9088 3856 9120
rect 3888 9088 3928 9120
rect 3960 9088 4000 9120
rect 0 9048 4000 9088
rect 0 9016 40 9048
rect 72 9016 112 9048
rect 144 9016 184 9048
rect 216 9016 256 9048
rect 288 9016 328 9048
rect 360 9016 400 9048
rect 432 9016 472 9048
rect 504 9016 544 9048
rect 576 9016 616 9048
rect 648 9016 688 9048
rect 720 9016 760 9048
rect 792 9016 832 9048
rect 864 9016 904 9048
rect 936 9016 976 9048
rect 1008 9016 1048 9048
rect 1080 9016 1120 9048
rect 1152 9016 1192 9048
rect 1224 9016 1264 9048
rect 1296 9016 1336 9048
rect 1368 9016 1408 9048
rect 1440 9016 1480 9048
rect 1512 9016 1552 9048
rect 1584 9016 1624 9048
rect 1656 9016 1696 9048
rect 1728 9016 1768 9048
rect 1800 9016 1840 9048
rect 1872 9016 1912 9048
rect 1944 9016 1984 9048
rect 2016 9016 2056 9048
rect 2088 9016 2128 9048
rect 2160 9016 2200 9048
rect 2232 9016 2272 9048
rect 2304 9016 2344 9048
rect 2376 9016 2416 9048
rect 2448 9016 2488 9048
rect 2520 9016 2560 9048
rect 2592 9016 2632 9048
rect 2664 9016 2704 9048
rect 2736 9016 2776 9048
rect 2808 9016 2848 9048
rect 2880 9016 2920 9048
rect 2952 9016 2992 9048
rect 3024 9016 3064 9048
rect 3096 9016 3136 9048
rect 3168 9016 3208 9048
rect 3240 9016 3280 9048
rect 3312 9016 3352 9048
rect 3384 9016 3424 9048
rect 3456 9016 3496 9048
rect 3528 9016 3568 9048
rect 3600 9016 3640 9048
rect 3672 9016 3712 9048
rect 3744 9016 3784 9048
rect 3816 9016 3856 9048
rect 3888 9016 3928 9048
rect 3960 9016 4000 9048
rect 0 8976 4000 9016
rect 0 8944 40 8976
rect 72 8944 112 8976
rect 144 8944 184 8976
rect 216 8944 256 8976
rect 288 8944 328 8976
rect 360 8944 400 8976
rect 432 8944 472 8976
rect 504 8944 544 8976
rect 576 8944 616 8976
rect 648 8944 688 8976
rect 720 8944 760 8976
rect 792 8944 832 8976
rect 864 8944 904 8976
rect 936 8944 976 8976
rect 1008 8944 1048 8976
rect 1080 8944 1120 8976
rect 1152 8944 1192 8976
rect 1224 8944 1264 8976
rect 1296 8944 1336 8976
rect 1368 8944 1408 8976
rect 1440 8944 1480 8976
rect 1512 8944 1552 8976
rect 1584 8944 1624 8976
rect 1656 8944 1696 8976
rect 1728 8944 1768 8976
rect 1800 8944 1840 8976
rect 1872 8944 1912 8976
rect 1944 8944 1984 8976
rect 2016 8944 2056 8976
rect 2088 8944 2128 8976
rect 2160 8944 2200 8976
rect 2232 8944 2272 8976
rect 2304 8944 2344 8976
rect 2376 8944 2416 8976
rect 2448 8944 2488 8976
rect 2520 8944 2560 8976
rect 2592 8944 2632 8976
rect 2664 8944 2704 8976
rect 2736 8944 2776 8976
rect 2808 8944 2848 8976
rect 2880 8944 2920 8976
rect 2952 8944 2992 8976
rect 3024 8944 3064 8976
rect 3096 8944 3136 8976
rect 3168 8944 3208 8976
rect 3240 8944 3280 8976
rect 3312 8944 3352 8976
rect 3384 8944 3424 8976
rect 3456 8944 3496 8976
rect 3528 8944 3568 8976
rect 3600 8944 3640 8976
rect 3672 8944 3712 8976
rect 3744 8944 3784 8976
rect 3816 8944 3856 8976
rect 3888 8944 3928 8976
rect 3960 8944 4000 8976
rect 0 8904 4000 8944
rect 0 8872 40 8904
rect 72 8872 112 8904
rect 144 8872 184 8904
rect 216 8872 256 8904
rect 288 8872 328 8904
rect 360 8872 400 8904
rect 432 8872 472 8904
rect 504 8872 544 8904
rect 576 8872 616 8904
rect 648 8872 688 8904
rect 720 8872 760 8904
rect 792 8872 832 8904
rect 864 8872 904 8904
rect 936 8872 976 8904
rect 1008 8872 1048 8904
rect 1080 8872 1120 8904
rect 1152 8872 1192 8904
rect 1224 8872 1264 8904
rect 1296 8872 1336 8904
rect 1368 8872 1408 8904
rect 1440 8872 1480 8904
rect 1512 8872 1552 8904
rect 1584 8872 1624 8904
rect 1656 8872 1696 8904
rect 1728 8872 1768 8904
rect 1800 8872 1840 8904
rect 1872 8872 1912 8904
rect 1944 8872 1984 8904
rect 2016 8872 2056 8904
rect 2088 8872 2128 8904
rect 2160 8872 2200 8904
rect 2232 8872 2272 8904
rect 2304 8872 2344 8904
rect 2376 8872 2416 8904
rect 2448 8872 2488 8904
rect 2520 8872 2560 8904
rect 2592 8872 2632 8904
rect 2664 8872 2704 8904
rect 2736 8872 2776 8904
rect 2808 8872 2848 8904
rect 2880 8872 2920 8904
rect 2952 8872 2992 8904
rect 3024 8872 3064 8904
rect 3096 8872 3136 8904
rect 3168 8872 3208 8904
rect 3240 8872 3280 8904
rect 3312 8872 3352 8904
rect 3384 8872 3424 8904
rect 3456 8872 3496 8904
rect 3528 8872 3568 8904
rect 3600 8872 3640 8904
rect 3672 8872 3712 8904
rect 3744 8872 3784 8904
rect 3816 8872 3856 8904
rect 3888 8872 3928 8904
rect 3960 8872 4000 8904
rect 0 8832 4000 8872
rect 0 8800 40 8832
rect 72 8800 112 8832
rect 144 8800 184 8832
rect 216 8800 256 8832
rect 288 8800 328 8832
rect 360 8800 400 8832
rect 432 8800 472 8832
rect 504 8800 544 8832
rect 576 8800 616 8832
rect 648 8800 688 8832
rect 720 8800 760 8832
rect 792 8800 832 8832
rect 864 8800 904 8832
rect 936 8800 976 8832
rect 1008 8800 1048 8832
rect 1080 8800 1120 8832
rect 1152 8800 1192 8832
rect 1224 8800 1264 8832
rect 1296 8800 1336 8832
rect 1368 8800 1408 8832
rect 1440 8800 1480 8832
rect 1512 8800 1552 8832
rect 1584 8800 1624 8832
rect 1656 8800 1696 8832
rect 1728 8800 1768 8832
rect 1800 8800 1840 8832
rect 1872 8800 1912 8832
rect 1944 8800 1984 8832
rect 2016 8800 2056 8832
rect 2088 8800 2128 8832
rect 2160 8800 2200 8832
rect 2232 8800 2272 8832
rect 2304 8800 2344 8832
rect 2376 8800 2416 8832
rect 2448 8800 2488 8832
rect 2520 8800 2560 8832
rect 2592 8800 2632 8832
rect 2664 8800 2704 8832
rect 2736 8800 2776 8832
rect 2808 8800 2848 8832
rect 2880 8800 2920 8832
rect 2952 8800 2992 8832
rect 3024 8800 3064 8832
rect 3096 8800 3136 8832
rect 3168 8800 3208 8832
rect 3240 8800 3280 8832
rect 3312 8800 3352 8832
rect 3384 8800 3424 8832
rect 3456 8800 3496 8832
rect 3528 8800 3568 8832
rect 3600 8800 3640 8832
rect 3672 8800 3712 8832
rect 3744 8800 3784 8832
rect 3816 8800 3856 8832
rect 3888 8800 3928 8832
rect 3960 8800 4000 8832
rect 0 8760 4000 8800
rect 0 8728 40 8760
rect 72 8728 112 8760
rect 144 8728 184 8760
rect 216 8728 256 8760
rect 288 8728 328 8760
rect 360 8728 400 8760
rect 432 8728 472 8760
rect 504 8728 544 8760
rect 576 8728 616 8760
rect 648 8728 688 8760
rect 720 8728 760 8760
rect 792 8728 832 8760
rect 864 8728 904 8760
rect 936 8728 976 8760
rect 1008 8728 1048 8760
rect 1080 8728 1120 8760
rect 1152 8728 1192 8760
rect 1224 8728 1264 8760
rect 1296 8728 1336 8760
rect 1368 8728 1408 8760
rect 1440 8728 1480 8760
rect 1512 8728 1552 8760
rect 1584 8728 1624 8760
rect 1656 8728 1696 8760
rect 1728 8728 1768 8760
rect 1800 8728 1840 8760
rect 1872 8728 1912 8760
rect 1944 8728 1984 8760
rect 2016 8728 2056 8760
rect 2088 8728 2128 8760
rect 2160 8728 2200 8760
rect 2232 8728 2272 8760
rect 2304 8728 2344 8760
rect 2376 8728 2416 8760
rect 2448 8728 2488 8760
rect 2520 8728 2560 8760
rect 2592 8728 2632 8760
rect 2664 8728 2704 8760
rect 2736 8728 2776 8760
rect 2808 8728 2848 8760
rect 2880 8728 2920 8760
rect 2952 8728 2992 8760
rect 3024 8728 3064 8760
rect 3096 8728 3136 8760
rect 3168 8728 3208 8760
rect 3240 8728 3280 8760
rect 3312 8728 3352 8760
rect 3384 8728 3424 8760
rect 3456 8728 3496 8760
rect 3528 8728 3568 8760
rect 3600 8728 3640 8760
rect 3672 8728 3712 8760
rect 3744 8728 3784 8760
rect 3816 8728 3856 8760
rect 3888 8728 3928 8760
rect 3960 8728 4000 8760
rect 0 8688 4000 8728
rect 0 8656 40 8688
rect 72 8656 112 8688
rect 144 8656 184 8688
rect 216 8656 256 8688
rect 288 8656 328 8688
rect 360 8656 400 8688
rect 432 8656 472 8688
rect 504 8656 544 8688
rect 576 8656 616 8688
rect 648 8656 688 8688
rect 720 8656 760 8688
rect 792 8656 832 8688
rect 864 8656 904 8688
rect 936 8656 976 8688
rect 1008 8656 1048 8688
rect 1080 8656 1120 8688
rect 1152 8656 1192 8688
rect 1224 8656 1264 8688
rect 1296 8656 1336 8688
rect 1368 8656 1408 8688
rect 1440 8656 1480 8688
rect 1512 8656 1552 8688
rect 1584 8656 1624 8688
rect 1656 8656 1696 8688
rect 1728 8656 1768 8688
rect 1800 8656 1840 8688
rect 1872 8656 1912 8688
rect 1944 8656 1984 8688
rect 2016 8656 2056 8688
rect 2088 8656 2128 8688
rect 2160 8656 2200 8688
rect 2232 8656 2272 8688
rect 2304 8656 2344 8688
rect 2376 8656 2416 8688
rect 2448 8656 2488 8688
rect 2520 8656 2560 8688
rect 2592 8656 2632 8688
rect 2664 8656 2704 8688
rect 2736 8656 2776 8688
rect 2808 8656 2848 8688
rect 2880 8656 2920 8688
rect 2952 8656 2992 8688
rect 3024 8656 3064 8688
rect 3096 8656 3136 8688
rect 3168 8656 3208 8688
rect 3240 8656 3280 8688
rect 3312 8656 3352 8688
rect 3384 8656 3424 8688
rect 3456 8656 3496 8688
rect 3528 8656 3568 8688
rect 3600 8656 3640 8688
rect 3672 8656 3712 8688
rect 3744 8656 3784 8688
rect 3816 8656 3856 8688
rect 3888 8656 3928 8688
rect 3960 8656 4000 8688
rect 0 8616 4000 8656
rect 0 8584 40 8616
rect 72 8584 112 8616
rect 144 8584 184 8616
rect 216 8584 256 8616
rect 288 8584 328 8616
rect 360 8584 400 8616
rect 432 8584 472 8616
rect 504 8584 544 8616
rect 576 8584 616 8616
rect 648 8584 688 8616
rect 720 8584 760 8616
rect 792 8584 832 8616
rect 864 8584 904 8616
rect 936 8584 976 8616
rect 1008 8584 1048 8616
rect 1080 8584 1120 8616
rect 1152 8584 1192 8616
rect 1224 8584 1264 8616
rect 1296 8584 1336 8616
rect 1368 8584 1408 8616
rect 1440 8584 1480 8616
rect 1512 8584 1552 8616
rect 1584 8584 1624 8616
rect 1656 8584 1696 8616
rect 1728 8584 1768 8616
rect 1800 8584 1840 8616
rect 1872 8584 1912 8616
rect 1944 8584 1984 8616
rect 2016 8584 2056 8616
rect 2088 8584 2128 8616
rect 2160 8584 2200 8616
rect 2232 8584 2272 8616
rect 2304 8584 2344 8616
rect 2376 8584 2416 8616
rect 2448 8584 2488 8616
rect 2520 8584 2560 8616
rect 2592 8584 2632 8616
rect 2664 8584 2704 8616
rect 2736 8584 2776 8616
rect 2808 8584 2848 8616
rect 2880 8584 2920 8616
rect 2952 8584 2992 8616
rect 3024 8584 3064 8616
rect 3096 8584 3136 8616
rect 3168 8584 3208 8616
rect 3240 8584 3280 8616
rect 3312 8584 3352 8616
rect 3384 8584 3424 8616
rect 3456 8584 3496 8616
rect 3528 8584 3568 8616
rect 3600 8584 3640 8616
rect 3672 8584 3712 8616
rect 3744 8584 3784 8616
rect 3816 8584 3856 8616
rect 3888 8584 3928 8616
rect 3960 8584 4000 8616
rect 0 8544 4000 8584
rect 0 8512 40 8544
rect 72 8512 112 8544
rect 144 8512 184 8544
rect 216 8512 256 8544
rect 288 8512 328 8544
rect 360 8512 400 8544
rect 432 8512 472 8544
rect 504 8512 544 8544
rect 576 8512 616 8544
rect 648 8512 688 8544
rect 720 8512 760 8544
rect 792 8512 832 8544
rect 864 8512 904 8544
rect 936 8512 976 8544
rect 1008 8512 1048 8544
rect 1080 8512 1120 8544
rect 1152 8512 1192 8544
rect 1224 8512 1264 8544
rect 1296 8512 1336 8544
rect 1368 8512 1408 8544
rect 1440 8512 1480 8544
rect 1512 8512 1552 8544
rect 1584 8512 1624 8544
rect 1656 8512 1696 8544
rect 1728 8512 1768 8544
rect 1800 8512 1840 8544
rect 1872 8512 1912 8544
rect 1944 8512 1984 8544
rect 2016 8512 2056 8544
rect 2088 8512 2128 8544
rect 2160 8512 2200 8544
rect 2232 8512 2272 8544
rect 2304 8512 2344 8544
rect 2376 8512 2416 8544
rect 2448 8512 2488 8544
rect 2520 8512 2560 8544
rect 2592 8512 2632 8544
rect 2664 8512 2704 8544
rect 2736 8512 2776 8544
rect 2808 8512 2848 8544
rect 2880 8512 2920 8544
rect 2952 8512 2992 8544
rect 3024 8512 3064 8544
rect 3096 8512 3136 8544
rect 3168 8512 3208 8544
rect 3240 8512 3280 8544
rect 3312 8512 3352 8544
rect 3384 8512 3424 8544
rect 3456 8512 3496 8544
rect 3528 8512 3568 8544
rect 3600 8512 3640 8544
rect 3672 8512 3712 8544
rect 3744 8512 3784 8544
rect 3816 8512 3856 8544
rect 3888 8512 3928 8544
rect 3960 8512 4000 8544
rect 0 8472 4000 8512
rect 0 8440 40 8472
rect 72 8440 112 8472
rect 144 8440 184 8472
rect 216 8440 256 8472
rect 288 8440 328 8472
rect 360 8440 400 8472
rect 432 8440 472 8472
rect 504 8440 544 8472
rect 576 8440 616 8472
rect 648 8440 688 8472
rect 720 8440 760 8472
rect 792 8440 832 8472
rect 864 8440 904 8472
rect 936 8440 976 8472
rect 1008 8440 1048 8472
rect 1080 8440 1120 8472
rect 1152 8440 1192 8472
rect 1224 8440 1264 8472
rect 1296 8440 1336 8472
rect 1368 8440 1408 8472
rect 1440 8440 1480 8472
rect 1512 8440 1552 8472
rect 1584 8440 1624 8472
rect 1656 8440 1696 8472
rect 1728 8440 1768 8472
rect 1800 8440 1840 8472
rect 1872 8440 1912 8472
rect 1944 8440 1984 8472
rect 2016 8440 2056 8472
rect 2088 8440 2128 8472
rect 2160 8440 2200 8472
rect 2232 8440 2272 8472
rect 2304 8440 2344 8472
rect 2376 8440 2416 8472
rect 2448 8440 2488 8472
rect 2520 8440 2560 8472
rect 2592 8440 2632 8472
rect 2664 8440 2704 8472
rect 2736 8440 2776 8472
rect 2808 8440 2848 8472
rect 2880 8440 2920 8472
rect 2952 8440 2992 8472
rect 3024 8440 3064 8472
rect 3096 8440 3136 8472
rect 3168 8440 3208 8472
rect 3240 8440 3280 8472
rect 3312 8440 3352 8472
rect 3384 8440 3424 8472
rect 3456 8440 3496 8472
rect 3528 8440 3568 8472
rect 3600 8440 3640 8472
rect 3672 8440 3712 8472
rect 3744 8440 3784 8472
rect 3816 8440 3856 8472
rect 3888 8440 3928 8472
rect 3960 8440 4000 8472
rect 0 8400 4000 8440
rect 0 8368 40 8400
rect 72 8368 112 8400
rect 144 8368 184 8400
rect 216 8368 256 8400
rect 288 8368 328 8400
rect 360 8368 400 8400
rect 432 8368 472 8400
rect 504 8368 544 8400
rect 576 8368 616 8400
rect 648 8368 688 8400
rect 720 8368 760 8400
rect 792 8368 832 8400
rect 864 8368 904 8400
rect 936 8368 976 8400
rect 1008 8368 1048 8400
rect 1080 8368 1120 8400
rect 1152 8368 1192 8400
rect 1224 8368 1264 8400
rect 1296 8368 1336 8400
rect 1368 8368 1408 8400
rect 1440 8368 1480 8400
rect 1512 8368 1552 8400
rect 1584 8368 1624 8400
rect 1656 8368 1696 8400
rect 1728 8368 1768 8400
rect 1800 8368 1840 8400
rect 1872 8368 1912 8400
rect 1944 8368 1984 8400
rect 2016 8368 2056 8400
rect 2088 8368 2128 8400
rect 2160 8368 2200 8400
rect 2232 8368 2272 8400
rect 2304 8368 2344 8400
rect 2376 8368 2416 8400
rect 2448 8368 2488 8400
rect 2520 8368 2560 8400
rect 2592 8368 2632 8400
rect 2664 8368 2704 8400
rect 2736 8368 2776 8400
rect 2808 8368 2848 8400
rect 2880 8368 2920 8400
rect 2952 8368 2992 8400
rect 3024 8368 3064 8400
rect 3096 8368 3136 8400
rect 3168 8368 3208 8400
rect 3240 8368 3280 8400
rect 3312 8368 3352 8400
rect 3384 8368 3424 8400
rect 3456 8368 3496 8400
rect 3528 8368 3568 8400
rect 3600 8368 3640 8400
rect 3672 8368 3712 8400
rect 3744 8368 3784 8400
rect 3816 8368 3856 8400
rect 3888 8368 3928 8400
rect 3960 8368 4000 8400
rect 0 8328 4000 8368
rect 0 8296 40 8328
rect 72 8296 112 8328
rect 144 8296 184 8328
rect 216 8296 256 8328
rect 288 8296 328 8328
rect 360 8296 400 8328
rect 432 8296 472 8328
rect 504 8296 544 8328
rect 576 8296 616 8328
rect 648 8296 688 8328
rect 720 8296 760 8328
rect 792 8296 832 8328
rect 864 8296 904 8328
rect 936 8296 976 8328
rect 1008 8296 1048 8328
rect 1080 8296 1120 8328
rect 1152 8296 1192 8328
rect 1224 8296 1264 8328
rect 1296 8296 1336 8328
rect 1368 8296 1408 8328
rect 1440 8296 1480 8328
rect 1512 8296 1552 8328
rect 1584 8296 1624 8328
rect 1656 8296 1696 8328
rect 1728 8296 1768 8328
rect 1800 8296 1840 8328
rect 1872 8296 1912 8328
rect 1944 8296 1984 8328
rect 2016 8296 2056 8328
rect 2088 8296 2128 8328
rect 2160 8296 2200 8328
rect 2232 8296 2272 8328
rect 2304 8296 2344 8328
rect 2376 8296 2416 8328
rect 2448 8296 2488 8328
rect 2520 8296 2560 8328
rect 2592 8296 2632 8328
rect 2664 8296 2704 8328
rect 2736 8296 2776 8328
rect 2808 8296 2848 8328
rect 2880 8296 2920 8328
rect 2952 8296 2992 8328
rect 3024 8296 3064 8328
rect 3096 8296 3136 8328
rect 3168 8296 3208 8328
rect 3240 8296 3280 8328
rect 3312 8296 3352 8328
rect 3384 8296 3424 8328
rect 3456 8296 3496 8328
rect 3528 8296 3568 8328
rect 3600 8296 3640 8328
rect 3672 8296 3712 8328
rect 3744 8296 3784 8328
rect 3816 8296 3856 8328
rect 3888 8296 3928 8328
rect 3960 8296 4000 8328
rect 0 8256 4000 8296
rect 0 8224 40 8256
rect 72 8224 112 8256
rect 144 8224 184 8256
rect 216 8224 256 8256
rect 288 8224 328 8256
rect 360 8224 400 8256
rect 432 8224 472 8256
rect 504 8224 544 8256
rect 576 8224 616 8256
rect 648 8224 688 8256
rect 720 8224 760 8256
rect 792 8224 832 8256
rect 864 8224 904 8256
rect 936 8224 976 8256
rect 1008 8224 1048 8256
rect 1080 8224 1120 8256
rect 1152 8224 1192 8256
rect 1224 8224 1264 8256
rect 1296 8224 1336 8256
rect 1368 8224 1408 8256
rect 1440 8224 1480 8256
rect 1512 8224 1552 8256
rect 1584 8224 1624 8256
rect 1656 8224 1696 8256
rect 1728 8224 1768 8256
rect 1800 8224 1840 8256
rect 1872 8224 1912 8256
rect 1944 8224 1984 8256
rect 2016 8224 2056 8256
rect 2088 8224 2128 8256
rect 2160 8224 2200 8256
rect 2232 8224 2272 8256
rect 2304 8224 2344 8256
rect 2376 8224 2416 8256
rect 2448 8224 2488 8256
rect 2520 8224 2560 8256
rect 2592 8224 2632 8256
rect 2664 8224 2704 8256
rect 2736 8224 2776 8256
rect 2808 8224 2848 8256
rect 2880 8224 2920 8256
rect 2952 8224 2992 8256
rect 3024 8224 3064 8256
rect 3096 8224 3136 8256
rect 3168 8224 3208 8256
rect 3240 8224 3280 8256
rect 3312 8224 3352 8256
rect 3384 8224 3424 8256
rect 3456 8224 3496 8256
rect 3528 8224 3568 8256
rect 3600 8224 3640 8256
rect 3672 8224 3712 8256
rect 3744 8224 3784 8256
rect 3816 8224 3856 8256
rect 3888 8224 3928 8256
rect 3960 8224 4000 8256
rect 0 8184 4000 8224
rect 0 8152 40 8184
rect 72 8152 112 8184
rect 144 8152 184 8184
rect 216 8152 256 8184
rect 288 8152 328 8184
rect 360 8152 400 8184
rect 432 8152 472 8184
rect 504 8152 544 8184
rect 576 8152 616 8184
rect 648 8152 688 8184
rect 720 8152 760 8184
rect 792 8152 832 8184
rect 864 8152 904 8184
rect 936 8152 976 8184
rect 1008 8152 1048 8184
rect 1080 8152 1120 8184
rect 1152 8152 1192 8184
rect 1224 8152 1264 8184
rect 1296 8152 1336 8184
rect 1368 8152 1408 8184
rect 1440 8152 1480 8184
rect 1512 8152 1552 8184
rect 1584 8152 1624 8184
rect 1656 8152 1696 8184
rect 1728 8152 1768 8184
rect 1800 8152 1840 8184
rect 1872 8152 1912 8184
rect 1944 8152 1984 8184
rect 2016 8152 2056 8184
rect 2088 8152 2128 8184
rect 2160 8152 2200 8184
rect 2232 8152 2272 8184
rect 2304 8152 2344 8184
rect 2376 8152 2416 8184
rect 2448 8152 2488 8184
rect 2520 8152 2560 8184
rect 2592 8152 2632 8184
rect 2664 8152 2704 8184
rect 2736 8152 2776 8184
rect 2808 8152 2848 8184
rect 2880 8152 2920 8184
rect 2952 8152 2992 8184
rect 3024 8152 3064 8184
rect 3096 8152 3136 8184
rect 3168 8152 3208 8184
rect 3240 8152 3280 8184
rect 3312 8152 3352 8184
rect 3384 8152 3424 8184
rect 3456 8152 3496 8184
rect 3528 8152 3568 8184
rect 3600 8152 3640 8184
rect 3672 8152 3712 8184
rect 3744 8152 3784 8184
rect 3816 8152 3856 8184
rect 3888 8152 3928 8184
rect 3960 8152 4000 8184
rect 0 8112 4000 8152
rect 0 8080 40 8112
rect 72 8080 112 8112
rect 144 8080 184 8112
rect 216 8080 256 8112
rect 288 8080 328 8112
rect 360 8080 400 8112
rect 432 8080 472 8112
rect 504 8080 544 8112
rect 576 8080 616 8112
rect 648 8080 688 8112
rect 720 8080 760 8112
rect 792 8080 832 8112
rect 864 8080 904 8112
rect 936 8080 976 8112
rect 1008 8080 1048 8112
rect 1080 8080 1120 8112
rect 1152 8080 1192 8112
rect 1224 8080 1264 8112
rect 1296 8080 1336 8112
rect 1368 8080 1408 8112
rect 1440 8080 1480 8112
rect 1512 8080 1552 8112
rect 1584 8080 1624 8112
rect 1656 8080 1696 8112
rect 1728 8080 1768 8112
rect 1800 8080 1840 8112
rect 1872 8080 1912 8112
rect 1944 8080 1984 8112
rect 2016 8080 2056 8112
rect 2088 8080 2128 8112
rect 2160 8080 2200 8112
rect 2232 8080 2272 8112
rect 2304 8080 2344 8112
rect 2376 8080 2416 8112
rect 2448 8080 2488 8112
rect 2520 8080 2560 8112
rect 2592 8080 2632 8112
rect 2664 8080 2704 8112
rect 2736 8080 2776 8112
rect 2808 8080 2848 8112
rect 2880 8080 2920 8112
rect 2952 8080 2992 8112
rect 3024 8080 3064 8112
rect 3096 8080 3136 8112
rect 3168 8080 3208 8112
rect 3240 8080 3280 8112
rect 3312 8080 3352 8112
rect 3384 8080 3424 8112
rect 3456 8080 3496 8112
rect 3528 8080 3568 8112
rect 3600 8080 3640 8112
rect 3672 8080 3712 8112
rect 3744 8080 3784 8112
rect 3816 8080 3856 8112
rect 3888 8080 3928 8112
rect 3960 8080 4000 8112
rect 0 8040 4000 8080
rect 0 8008 40 8040
rect 72 8008 112 8040
rect 144 8008 184 8040
rect 216 8008 256 8040
rect 288 8008 328 8040
rect 360 8008 400 8040
rect 432 8008 472 8040
rect 504 8008 544 8040
rect 576 8008 616 8040
rect 648 8008 688 8040
rect 720 8008 760 8040
rect 792 8008 832 8040
rect 864 8008 904 8040
rect 936 8008 976 8040
rect 1008 8008 1048 8040
rect 1080 8008 1120 8040
rect 1152 8008 1192 8040
rect 1224 8008 1264 8040
rect 1296 8008 1336 8040
rect 1368 8008 1408 8040
rect 1440 8008 1480 8040
rect 1512 8008 1552 8040
rect 1584 8008 1624 8040
rect 1656 8008 1696 8040
rect 1728 8008 1768 8040
rect 1800 8008 1840 8040
rect 1872 8008 1912 8040
rect 1944 8008 1984 8040
rect 2016 8008 2056 8040
rect 2088 8008 2128 8040
rect 2160 8008 2200 8040
rect 2232 8008 2272 8040
rect 2304 8008 2344 8040
rect 2376 8008 2416 8040
rect 2448 8008 2488 8040
rect 2520 8008 2560 8040
rect 2592 8008 2632 8040
rect 2664 8008 2704 8040
rect 2736 8008 2776 8040
rect 2808 8008 2848 8040
rect 2880 8008 2920 8040
rect 2952 8008 2992 8040
rect 3024 8008 3064 8040
rect 3096 8008 3136 8040
rect 3168 8008 3208 8040
rect 3240 8008 3280 8040
rect 3312 8008 3352 8040
rect 3384 8008 3424 8040
rect 3456 8008 3496 8040
rect 3528 8008 3568 8040
rect 3600 8008 3640 8040
rect 3672 8008 3712 8040
rect 3744 8008 3784 8040
rect 3816 8008 3856 8040
rect 3888 8008 3928 8040
rect 3960 8008 4000 8040
rect 0 7968 4000 8008
rect 0 7936 40 7968
rect 72 7936 112 7968
rect 144 7936 184 7968
rect 216 7936 256 7968
rect 288 7936 328 7968
rect 360 7936 400 7968
rect 432 7936 472 7968
rect 504 7936 544 7968
rect 576 7936 616 7968
rect 648 7936 688 7968
rect 720 7936 760 7968
rect 792 7936 832 7968
rect 864 7936 904 7968
rect 936 7936 976 7968
rect 1008 7936 1048 7968
rect 1080 7936 1120 7968
rect 1152 7936 1192 7968
rect 1224 7936 1264 7968
rect 1296 7936 1336 7968
rect 1368 7936 1408 7968
rect 1440 7936 1480 7968
rect 1512 7936 1552 7968
rect 1584 7936 1624 7968
rect 1656 7936 1696 7968
rect 1728 7936 1768 7968
rect 1800 7936 1840 7968
rect 1872 7936 1912 7968
rect 1944 7936 1984 7968
rect 2016 7936 2056 7968
rect 2088 7936 2128 7968
rect 2160 7936 2200 7968
rect 2232 7936 2272 7968
rect 2304 7936 2344 7968
rect 2376 7936 2416 7968
rect 2448 7936 2488 7968
rect 2520 7936 2560 7968
rect 2592 7936 2632 7968
rect 2664 7936 2704 7968
rect 2736 7936 2776 7968
rect 2808 7936 2848 7968
rect 2880 7936 2920 7968
rect 2952 7936 2992 7968
rect 3024 7936 3064 7968
rect 3096 7936 3136 7968
rect 3168 7936 3208 7968
rect 3240 7936 3280 7968
rect 3312 7936 3352 7968
rect 3384 7936 3424 7968
rect 3456 7936 3496 7968
rect 3528 7936 3568 7968
rect 3600 7936 3640 7968
rect 3672 7936 3712 7968
rect 3744 7936 3784 7968
rect 3816 7936 3856 7968
rect 3888 7936 3928 7968
rect 3960 7936 4000 7968
rect 0 7896 4000 7936
rect 0 7864 40 7896
rect 72 7864 112 7896
rect 144 7864 184 7896
rect 216 7864 256 7896
rect 288 7864 328 7896
rect 360 7864 400 7896
rect 432 7864 472 7896
rect 504 7864 544 7896
rect 576 7864 616 7896
rect 648 7864 688 7896
rect 720 7864 760 7896
rect 792 7864 832 7896
rect 864 7864 904 7896
rect 936 7864 976 7896
rect 1008 7864 1048 7896
rect 1080 7864 1120 7896
rect 1152 7864 1192 7896
rect 1224 7864 1264 7896
rect 1296 7864 1336 7896
rect 1368 7864 1408 7896
rect 1440 7864 1480 7896
rect 1512 7864 1552 7896
rect 1584 7864 1624 7896
rect 1656 7864 1696 7896
rect 1728 7864 1768 7896
rect 1800 7864 1840 7896
rect 1872 7864 1912 7896
rect 1944 7864 1984 7896
rect 2016 7864 2056 7896
rect 2088 7864 2128 7896
rect 2160 7864 2200 7896
rect 2232 7864 2272 7896
rect 2304 7864 2344 7896
rect 2376 7864 2416 7896
rect 2448 7864 2488 7896
rect 2520 7864 2560 7896
rect 2592 7864 2632 7896
rect 2664 7864 2704 7896
rect 2736 7864 2776 7896
rect 2808 7864 2848 7896
rect 2880 7864 2920 7896
rect 2952 7864 2992 7896
rect 3024 7864 3064 7896
rect 3096 7864 3136 7896
rect 3168 7864 3208 7896
rect 3240 7864 3280 7896
rect 3312 7864 3352 7896
rect 3384 7864 3424 7896
rect 3456 7864 3496 7896
rect 3528 7864 3568 7896
rect 3600 7864 3640 7896
rect 3672 7864 3712 7896
rect 3744 7864 3784 7896
rect 3816 7864 3856 7896
rect 3888 7864 3928 7896
rect 3960 7864 4000 7896
rect 0 7824 4000 7864
rect 0 7792 40 7824
rect 72 7792 112 7824
rect 144 7792 184 7824
rect 216 7792 256 7824
rect 288 7792 328 7824
rect 360 7792 400 7824
rect 432 7792 472 7824
rect 504 7792 544 7824
rect 576 7792 616 7824
rect 648 7792 688 7824
rect 720 7792 760 7824
rect 792 7792 832 7824
rect 864 7792 904 7824
rect 936 7792 976 7824
rect 1008 7792 1048 7824
rect 1080 7792 1120 7824
rect 1152 7792 1192 7824
rect 1224 7792 1264 7824
rect 1296 7792 1336 7824
rect 1368 7792 1408 7824
rect 1440 7792 1480 7824
rect 1512 7792 1552 7824
rect 1584 7792 1624 7824
rect 1656 7792 1696 7824
rect 1728 7792 1768 7824
rect 1800 7792 1840 7824
rect 1872 7792 1912 7824
rect 1944 7792 1984 7824
rect 2016 7792 2056 7824
rect 2088 7792 2128 7824
rect 2160 7792 2200 7824
rect 2232 7792 2272 7824
rect 2304 7792 2344 7824
rect 2376 7792 2416 7824
rect 2448 7792 2488 7824
rect 2520 7792 2560 7824
rect 2592 7792 2632 7824
rect 2664 7792 2704 7824
rect 2736 7792 2776 7824
rect 2808 7792 2848 7824
rect 2880 7792 2920 7824
rect 2952 7792 2992 7824
rect 3024 7792 3064 7824
rect 3096 7792 3136 7824
rect 3168 7792 3208 7824
rect 3240 7792 3280 7824
rect 3312 7792 3352 7824
rect 3384 7792 3424 7824
rect 3456 7792 3496 7824
rect 3528 7792 3568 7824
rect 3600 7792 3640 7824
rect 3672 7792 3712 7824
rect 3744 7792 3784 7824
rect 3816 7792 3856 7824
rect 3888 7792 3928 7824
rect 3960 7792 4000 7824
rect 0 7752 4000 7792
rect 0 7720 40 7752
rect 72 7720 112 7752
rect 144 7720 184 7752
rect 216 7720 256 7752
rect 288 7720 328 7752
rect 360 7720 400 7752
rect 432 7720 472 7752
rect 504 7720 544 7752
rect 576 7720 616 7752
rect 648 7720 688 7752
rect 720 7720 760 7752
rect 792 7720 832 7752
rect 864 7720 904 7752
rect 936 7720 976 7752
rect 1008 7720 1048 7752
rect 1080 7720 1120 7752
rect 1152 7720 1192 7752
rect 1224 7720 1264 7752
rect 1296 7720 1336 7752
rect 1368 7720 1408 7752
rect 1440 7720 1480 7752
rect 1512 7720 1552 7752
rect 1584 7720 1624 7752
rect 1656 7720 1696 7752
rect 1728 7720 1768 7752
rect 1800 7720 1840 7752
rect 1872 7720 1912 7752
rect 1944 7720 1984 7752
rect 2016 7720 2056 7752
rect 2088 7720 2128 7752
rect 2160 7720 2200 7752
rect 2232 7720 2272 7752
rect 2304 7720 2344 7752
rect 2376 7720 2416 7752
rect 2448 7720 2488 7752
rect 2520 7720 2560 7752
rect 2592 7720 2632 7752
rect 2664 7720 2704 7752
rect 2736 7720 2776 7752
rect 2808 7720 2848 7752
rect 2880 7720 2920 7752
rect 2952 7720 2992 7752
rect 3024 7720 3064 7752
rect 3096 7720 3136 7752
rect 3168 7720 3208 7752
rect 3240 7720 3280 7752
rect 3312 7720 3352 7752
rect 3384 7720 3424 7752
rect 3456 7720 3496 7752
rect 3528 7720 3568 7752
rect 3600 7720 3640 7752
rect 3672 7720 3712 7752
rect 3744 7720 3784 7752
rect 3816 7720 3856 7752
rect 3888 7720 3928 7752
rect 3960 7720 4000 7752
rect 0 7680 4000 7720
rect 0 7648 40 7680
rect 72 7648 112 7680
rect 144 7648 184 7680
rect 216 7648 256 7680
rect 288 7648 328 7680
rect 360 7648 400 7680
rect 432 7648 472 7680
rect 504 7648 544 7680
rect 576 7648 616 7680
rect 648 7648 688 7680
rect 720 7648 760 7680
rect 792 7648 832 7680
rect 864 7648 904 7680
rect 936 7648 976 7680
rect 1008 7648 1048 7680
rect 1080 7648 1120 7680
rect 1152 7648 1192 7680
rect 1224 7648 1264 7680
rect 1296 7648 1336 7680
rect 1368 7648 1408 7680
rect 1440 7648 1480 7680
rect 1512 7648 1552 7680
rect 1584 7648 1624 7680
rect 1656 7648 1696 7680
rect 1728 7648 1768 7680
rect 1800 7648 1840 7680
rect 1872 7648 1912 7680
rect 1944 7648 1984 7680
rect 2016 7648 2056 7680
rect 2088 7648 2128 7680
rect 2160 7648 2200 7680
rect 2232 7648 2272 7680
rect 2304 7648 2344 7680
rect 2376 7648 2416 7680
rect 2448 7648 2488 7680
rect 2520 7648 2560 7680
rect 2592 7648 2632 7680
rect 2664 7648 2704 7680
rect 2736 7648 2776 7680
rect 2808 7648 2848 7680
rect 2880 7648 2920 7680
rect 2952 7648 2992 7680
rect 3024 7648 3064 7680
rect 3096 7648 3136 7680
rect 3168 7648 3208 7680
rect 3240 7648 3280 7680
rect 3312 7648 3352 7680
rect 3384 7648 3424 7680
rect 3456 7648 3496 7680
rect 3528 7648 3568 7680
rect 3600 7648 3640 7680
rect 3672 7648 3712 7680
rect 3744 7648 3784 7680
rect 3816 7648 3856 7680
rect 3888 7648 3928 7680
rect 3960 7648 4000 7680
rect 0 7608 4000 7648
rect 0 7576 40 7608
rect 72 7576 112 7608
rect 144 7576 184 7608
rect 216 7576 256 7608
rect 288 7576 328 7608
rect 360 7576 400 7608
rect 432 7576 472 7608
rect 504 7576 544 7608
rect 576 7576 616 7608
rect 648 7576 688 7608
rect 720 7576 760 7608
rect 792 7576 832 7608
rect 864 7576 904 7608
rect 936 7576 976 7608
rect 1008 7576 1048 7608
rect 1080 7576 1120 7608
rect 1152 7576 1192 7608
rect 1224 7576 1264 7608
rect 1296 7576 1336 7608
rect 1368 7576 1408 7608
rect 1440 7576 1480 7608
rect 1512 7576 1552 7608
rect 1584 7576 1624 7608
rect 1656 7576 1696 7608
rect 1728 7576 1768 7608
rect 1800 7576 1840 7608
rect 1872 7576 1912 7608
rect 1944 7576 1984 7608
rect 2016 7576 2056 7608
rect 2088 7576 2128 7608
rect 2160 7576 2200 7608
rect 2232 7576 2272 7608
rect 2304 7576 2344 7608
rect 2376 7576 2416 7608
rect 2448 7576 2488 7608
rect 2520 7576 2560 7608
rect 2592 7576 2632 7608
rect 2664 7576 2704 7608
rect 2736 7576 2776 7608
rect 2808 7576 2848 7608
rect 2880 7576 2920 7608
rect 2952 7576 2992 7608
rect 3024 7576 3064 7608
rect 3096 7576 3136 7608
rect 3168 7576 3208 7608
rect 3240 7576 3280 7608
rect 3312 7576 3352 7608
rect 3384 7576 3424 7608
rect 3456 7576 3496 7608
rect 3528 7576 3568 7608
rect 3600 7576 3640 7608
rect 3672 7576 3712 7608
rect 3744 7576 3784 7608
rect 3816 7576 3856 7608
rect 3888 7576 3928 7608
rect 3960 7576 4000 7608
rect 0 7536 4000 7576
rect 0 7504 40 7536
rect 72 7504 112 7536
rect 144 7504 184 7536
rect 216 7504 256 7536
rect 288 7504 328 7536
rect 360 7504 400 7536
rect 432 7504 472 7536
rect 504 7504 544 7536
rect 576 7504 616 7536
rect 648 7504 688 7536
rect 720 7504 760 7536
rect 792 7504 832 7536
rect 864 7504 904 7536
rect 936 7504 976 7536
rect 1008 7504 1048 7536
rect 1080 7504 1120 7536
rect 1152 7504 1192 7536
rect 1224 7504 1264 7536
rect 1296 7504 1336 7536
rect 1368 7504 1408 7536
rect 1440 7504 1480 7536
rect 1512 7504 1552 7536
rect 1584 7504 1624 7536
rect 1656 7504 1696 7536
rect 1728 7504 1768 7536
rect 1800 7504 1840 7536
rect 1872 7504 1912 7536
rect 1944 7504 1984 7536
rect 2016 7504 2056 7536
rect 2088 7504 2128 7536
rect 2160 7504 2200 7536
rect 2232 7504 2272 7536
rect 2304 7504 2344 7536
rect 2376 7504 2416 7536
rect 2448 7504 2488 7536
rect 2520 7504 2560 7536
rect 2592 7504 2632 7536
rect 2664 7504 2704 7536
rect 2736 7504 2776 7536
rect 2808 7504 2848 7536
rect 2880 7504 2920 7536
rect 2952 7504 2992 7536
rect 3024 7504 3064 7536
rect 3096 7504 3136 7536
rect 3168 7504 3208 7536
rect 3240 7504 3280 7536
rect 3312 7504 3352 7536
rect 3384 7504 3424 7536
rect 3456 7504 3496 7536
rect 3528 7504 3568 7536
rect 3600 7504 3640 7536
rect 3672 7504 3712 7536
rect 3744 7504 3784 7536
rect 3816 7504 3856 7536
rect 3888 7504 3928 7536
rect 3960 7504 4000 7536
rect 0 7464 4000 7504
rect 0 7432 40 7464
rect 72 7432 112 7464
rect 144 7432 184 7464
rect 216 7432 256 7464
rect 288 7432 328 7464
rect 360 7432 400 7464
rect 432 7432 472 7464
rect 504 7432 544 7464
rect 576 7432 616 7464
rect 648 7432 688 7464
rect 720 7432 760 7464
rect 792 7432 832 7464
rect 864 7432 904 7464
rect 936 7432 976 7464
rect 1008 7432 1048 7464
rect 1080 7432 1120 7464
rect 1152 7432 1192 7464
rect 1224 7432 1264 7464
rect 1296 7432 1336 7464
rect 1368 7432 1408 7464
rect 1440 7432 1480 7464
rect 1512 7432 1552 7464
rect 1584 7432 1624 7464
rect 1656 7432 1696 7464
rect 1728 7432 1768 7464
rect 1800 7432 1840 7464
rect 1872 7432 1912 7464
rect 1944 7432 1984 7464
rect 2016 7432 2056 7464
rect 2088 7432 2128 7464
rect 2160 7432 2200 7464
rect 2232 7432 2272 7464
rect 2304 7432 2344 7464
rect 2376 7432 2416 7464
rect 2448 7432 2488 7464
rect 2520 7432 2560 7464
rect 2592 7432 2632 7464
rect 2664 7432 2704 7464
rect 2736 7432 2776 7464
rect 2808 7432 2848 7464
rect 2880 7432 2920 7464
rect 2952 7432 2992 7464
rect 3024 7432 3064 7464
rect 3096 7432 3136 7464
rect 3168 7432 3208 7464
rect 3240 7432 3280 7464
rect 3312 7432 3352 7464
rect 3384 7432 3424 7464
rect 3456 7432 3496 7464
rect 3528 7432 3568 7464
rect 3600 7432 3640 7464
rect 3672 7432 3712 7464
rect 3744 7432 3784 7464
rect 3816 7432 3856 7464
rect 3888 7432 3928 7464
rect 3960 7432 4000 7464
rect 0 7392 4000 7432
rect 0 7360 40 7392
rect 72 7360 112 7392
rect 144 7360 184 7392
rect 216 7360 256 7392
rect 288 7360 328 7392
rect 360 7360 400 7392
rect 432 7360 472 7392
rect 504 7360 544 7392
rect 576 7360 616 7392
rect 648 7360 688 7392
rect 720 7360 760 7392
rect 792 7360 832 7392
rect 864 7360 904 7392
rect 936 7360 976 7392
rect 1008 7360 1048 7392
rect 1080 7360 1120 7392
rect 1152 7360 1192 7392
rect 1224 7360 1264 7392
rect 1296 7360 1336 7392
rect 1368 7360 1408 7392
rect 1440 7360 1480 7392
rect 1512 7360 1552 7392
rect 1584 7360 1624 7392
rect 1656 7360 1696 7392
rect 1728 7360 1768 7392
rect 1800 7360 1840 7392
rect 1872 7360 1912 7392
rect 1944 7360 1984 7392
rect 2016 7360 2056 7392
rect 2088 7360 2128 7392
rect 2160 7360 2200 7392
rect 2232 7360 2272 7392
rect 2304 7360 2344 7392
rect 2376 7360 2416 7392
rect 2448 7360 2488 7392
rect 2520 7360 2560 7392
rect 2592 7360 2632 7392
rect 2664 7360 2704 7392
rect 2736 7360 2776 7392
rect 2808 7360 2848 7392
rect 2880 7360 2920 7392
rect 2952 7360 2992 7392
rect 3024 7360 3064 7392
rect 3096 7360 3136 7392
rect 3168 7360 3208 7392
rect 3240 7360 3280 7392
rect 3312 7360 3352 7392
rect 3384 7360 3424 7392
rect 3456 7360 3496 7392
rect 3528 7360 3568 7392
rect 3600 7360 3640 7392
rect 3672 7360 3712 7392
rect 3744 7360 3784 7392
rect 3816 7360 3856 7392
rect 3888 7360 3928 7392
rect 3960 7360 4000 7392
rect 0 7320 4000 7360
rect 0 7288 40 7320
rect 72 7288 112 7320
rect 144 7288 184 7320
rect 216 7288 256 7320
rect 288 7288 328 7320
rect 360 7288 400 7320
rect 432 7288 472 7320
rect 504 7288 544 7320
rect 576 7288 616 7320
rect 648 7288 688 7320
rect 720 7288 760 7320
rect 792 7288 832 7320
rect 864 7288 904 7320
rect 936 7288 976 7320
rect 1008 7288 1048 7320
rect 1080 7288 1120 7320
rect 1152 7288 1192 7320
rect 1224 7288 1264 7320
rect 1296 7288 1336 7320
rect 1368 7288 1408 7320
rect 1440 7288 1480 7320
rect 1512 7288 1552 7320
rect 1584 7288 1624 7320
rect 1656 7288 1696 7320
rect 1728 7288 1768 7320
rect 1800 7288 1840 7320
rect 1872 7288 1912 7320
rect 1944 7288 1984 7320
rect 2016 7288 2056 7320
rect 2088 7288 2128 7320
rect 2160 7288 2200 7320
rect 2232 7288 2272 7320
rect 2304 7288 2344 7320
rect 2376 7288 2416 7320
rect 2448 7288 2488 7320
rect 2520 7288 2560 7320
rect 2592 7288 2632 7320
rect 2664 7288 2704 7320
rect 2736 7288 2776 7320
rect 2808 7288 2848 7320
rect 2880 7288 2920 7320
rect 2952 7288 2992 7320
rect 3024 7288 3064 7320
rect 3096 7288 3136 7320
rect 3168 7288 3208 7320
rect 3240 7288 3280 7320
rect 3312 7288 3352 7320
rect 3384 7288 3424 7320
rect 3456 7288 3496 7320
rect 3528 7288 3568 7320
rect 3600 7288 3640 7320
rect 3672 7288 3712 7320
rect 3744 7288 3784 7320
rect 3816 7288 3856 7320
rect 3888 7288 3928 7320
rect 3960 7288 4000 7320
rect 0 7248 4000 7288
rect 0 7216 40 7248
rect 72 7216 112 7248
rect 144 7216 184 7248
rect 216 7216 256 7248
rect 288 7216 328 7248
rect 360 7216 400 7248
rect 432 7216 472 7248
rect 504 7216 544 7248
rect 576 7216 616 7248
rect 648 7216 688 7248
rect 720 7216 760 7248
rect 792 7216 832 7248
rect 864 7216 904 7248
rect 936 7216 976 7248
rect 1008 7216 1048 7248
rect 1080 7216 1120 7248
rect 1152 7216 1192 7248
rect 1224 7216 1264 7248
rect 1296 7216 1336 7248
rect 1368 7216 1408 7248
rect 1440 7216 1480 7248
rect 1512 7216 1552 7248
rect 1584 7216 1624 7248
rect 1656 7216 1696 7248
rect 1728 7216 1768 7248
rect 1800 7216 1840 7248
rect 1872 7216 1912 7248
rect 1944 7216 1984 7248
rect 2016 7216 2056 7248
rect 2088 7216 2128 7248
rect 2160 7216 2200 7248
rect 2232 7216 2272 7248
rect 2304 7216 2344 7248
rect 2376 7216 2416 7248
rect 2448 7216 2488 7248
rect 2520 7216 2560 7248
rect 2592 7216 2632 7248
rect 2664 7216 2704 7248
rect 2736 7216 2776 7248
rect 2808 7216 2848 7248
rect 2880 7216 2920 7248
rect 2952 7216 2992 7248
rect 3024 7216 3064 7248
rect 3096 7216 3136 7248
rect 3168 7216 3208 7248
rect 3240 7216 3280 7248
rect 3312 7216 3352 7248
rect 3384 7216 3424 7248
rect 3456 7216 3496 7248
rect 3528 7216 3568 7248
rect 3600 7216 3640 7248
rect 3672 7216 3712 7248
rect 3744 7216 3784 7248
rect 3816 7216 3856 7248
rect 3888 7216 3928 7248
rect 3960 7216 4000 7248
rect 0 7176 4000 7216
rect 0 7144 40 7176
rect 72 7144 112 7176
rect 144 7144 184 7176
rect 216 7144 256 7176
rect 288 7144 328 7176
rect 360 7144 400 7176
rect 432 7144 472 7176
rect 504 7144 544 7176
rect 576 7144 616 7176
rect 648 7144 688 7176
rect 720 7144 760 7176
rect 792 7144 832 7176
rect 864 7144 904 7176
rect 936 7144 976 7176
rect 1008 7144 1048 7176
rect 1080 7144 1120 7176
rect 1152 7144 1192 7176
rect 1224 7144 1264 7176
rect 1296 7144 1336 7176
rect 1368 7144 1408 7176
rect 1440 7144 1480 7176
rect 1512 7144 1552 7176
rect 1584 7144 1624 7176
rect 1656 7144 1696 7176
rect 1728 7144 1768 7176
rect 1800 7144 1840 7176
rect 1872 7144 1912 7176
rect 1944 7144 1984 7176
rect 2016 7144 2056 7176
rect 2088 7144 2128 7176
rect 2160 7144 2200 7176
rect 2232 7144 2272 7176
rect 2304 7144 2344 7176
rect 2376 7144 2416 7176
rect 2448 7144 2488 7176
rect 2520 7144 2560 7176
rect 2592 7144 2632 7176
rect 2664 7144 2704 7176
rect 2736 7144 2776 7176
rect 2808 7144 2848 7176
rect 2880 7144 2920 7176
rect 2952 7144 2992 7176
rect 3024 7144 3064 7176
rect 3096 7144 3136 7176
rect 3168 7144 3208 7176
rect 3240 7144 3280 7176
rect 3312 7144 3352 7176
rect 3384 7144 3424 7176
rect 3456 7144 3496 7176
rect 3528 7144 3568 7176
rect 3600 7144 3640 7176
rect 3672 7144 3712 7176
rect 3744 7144 3784 7176
rect 3816 7144 3856 7176
rect 3888 7144 3928 7176
rect 3960 7144 4000 7176
rect 0 7104 4000 7144
rect 0 7072 40 7104
rect 72 7072 112 7104
rect 144 7072 184 7104
rect 216 7072 256 7104
rect 288 7072 328 7104
rect 360 7072 400 7104
rect 432 7072 472 7104
rect 504 7072 544 7104
rect 576 7072 616 7104
rect 648 7072 688 7104
rect 720 7072 760 7104
rect 792 7072 832 7104
rect 864 7072 904 7104
rect 936 7072 976 7104
rect 1008 7072 1048 7104
rect 1080 7072 1120 7104
rect 1152 7072 1192 7104
rect 1224 7072 1264 7104
rect 1296 7072 1336 7104
rect 1368 7072 1408 7104
rect 1440 7072 1480 7104
rect 1512 7072 1552 7104
rect 1584 7072 1624 7104
rect 1656 7072 1696 7104
rect 1728 7072 1768 7104
rect 1800 7072 1840 7104
rect 1872 7072 1912 7104
rect 1944 7072 1984 7104
rect 2016 7072 2056 7104
rect 2088 7072 2128 7104
rect 2160 7072 2200 7104
rect 2232 7072 2272 7104
rect 2304 7072 2344 7104
rect 2376 7072 2416 7104
rect 2448 7072 2488 7104
rect 2520 7072 2560 7104
rect 2592 7072 2632 7104
rect 2664 7072 2704 7104
rect 2736 7072 2776 7104
rect 2808 7072 2848 7104
rect 2880 7072 2920 7104
rect 2952 7072 2992 7104
rect 3024 7072 3064 7104
rect 3096 7072 3136 7104
rect 3168 7072 3208 7104
rect 3240 7072 3280 7104
rect 3312 7072 3352 7104
rect 3384 7072 3424 7104
rect 3456 7072 3496 7104
rect 3528 7072 3568 7104
rect 3600 7072 3640 7104
rect 3672 7072 3712 7104
rect 3744 7072 3784 7104
rect 3816 7072 3856 7104
rect 3888 7072 3928 7104
rect 3960 7072 4000 7104
rect 0 7032 4000 7072
rect 0 7000 40 7032
rect 72 7000 112 7032
rect 144 7000 184 7032
rect 216 7000 256 7032
rect 288 7000 328 7032
rect 360 7000 400 7032
rect 432 7000 472 7032
rect 504 7000 544 7032
rect 576 7000 616 7032
rect 648 7000 688 7032
rect 720 7000 760 7032
rect 792 7000 832 7032
rect 864 7000 904 7032
rect 936 7000 976 7032
rect 1008 7000 1048 7032
rect 1080 7000 1120 7032
rect 1152 7000 1192 7032
rect 1224 7000 1264 7032
rect 1296 7000 1336 7032
rect 1368 7000 1408 7032
rect 1440 7000 1480 7032
rect 1512 7000 1552 7032
rect 1584 7000 1624 7032
rect 1656 7000 1696 7032
rect 1728 7000 1768 7032
rect 1800 7000 1840 7032
rect 1872 7000 1912 7032
rect 1944 7000 1984 7032
rect 2016 7000 2056 7032
rect 2088 7000 2128 7032
rect 2160 7000 2200 7032
rect 2232 7000 2272 7032
rect 2304 7000 2344 7032
rect 2376 7000 2416 7032
rect 2448 7000 2488 7032
rect 2520 7000 2560 7032
rect 2592 7000 2632 7032
rect 2664 7000 2704 7032
rect 2736 7000 2776 7032
rect 2808 7000 2848 7032
rect 2880 7000 2920 7032
rect 2952 7000 2992 7032
rect 3024 7000 3064 7032
rect 3096 7000 3136 7032
rect 3168 7000 3208 7032
rect 3240 7000 3280 7032
rect 3312 7000 3352 7032
rect 3384 7000 3424 7032
rect 3456 7000 3496 7032
rect 3528 7000 3568 7032
rect 3600 7000 3640 7032
rect 3672 7000 3712 7032
rect 3744 7000 3784 7032
rect 3816 7000 3856 7032
rect 3888 7000 3928 7032
rect 3960 7000 4000 7032
rect 0 6960 4000 7000
rect 0 6928 40 6960
rect 72 6928 112 6960
rect 144 6928 184 6960
rect 216 6928 256 6960
rect 288 6928 328 6960
rect 360 6928 400 6960
rect 432 6928 472 6960
rect 504 6928 544 6960
rect 576 6928 616 6960
rect 648 6928 688 6960
rect 720 6928 760 6960
rect 792 6928 832 6960
rect 864 6928 904 6960
rect 936 6928 976 6960
rect 1008 6928 1048 6960
rect 1080 6928 1120 6960
rect 1152 6928 1192 6960
rect 1224 6928 1264 6960
rect 1296 6928 1336 6960
rect 1368 6928 1408 6960
rect 1440 6928 1480 6960
rect 1512 6928 1552 6960
rect 1584 6928 1624 6960
rect 1656 6928 1696 6960
rect 1728 6928 1768 6960
rect 1800 6928 1840 6960
rect 1872 6928 1912 6960
rect 1944 6928 1984 6960
rect 2016 6928 2056 6960
rect 2088 6928 2128 6960
rect 2160 6928 2200 6960
rect 2232 6928 2272 6960
rect 2304 6928 2344 6960
rect 2376 6928 2416 6960
rect 2448 6928 2488 6960
rect 2520 6928 2560 6960
rect 2592 6928 2632 6960
rect 2664 6928 2704 6960
rect 2736 6928 2776 6960
rect 2808 6928 2848 6960
rect 2880 6928 2920 6960
rect 2952 6928 2992 6960
rect 3024 6928 3064 6960
rect 3096 6928 3136 6960
rect 3168 6928 3208 6960
rect 3240 6928 3280 6960
rect 3312 6928 3352 6960
rect 3384 6928 3424 6960
rect 3456 6928 3496 6960
rect 3528 6928 3568 6960
rect 3600 6928 3640 6960
rect 3672 6928 3712 6960
rect 3744 6928 3784 6960
rect 3816 6928 3856 6960
rect 3888 6928 3928 6960
rect 3960 6928 4000 6960
rect 0 6888 4000 6928
rect 0 6856 40 6888
rect 72 6856 112 6888
rect 144 6856 184 6888
rect 216 6856 256 6888
rect 288 6856 328 6888
rect 360 6856 400 6888
rect 432 6856 472 6888
rect 504 6856 544 6888
rect 576 6856 616 6888
rect 648 6856 688 6888
rect 720 6856 760 6888
rect 792 6856 832 6888
rect 864 6856 904 6888
rect 936 6856 976 6888
rect 1008 6856 1048 6888
rect 1080 6856 1120 6888
rect 1152 6856 1192 6888
rect 1224 6856 1264 6888
rect 1296 6856 1336 6888
rect 1368 6856 1408 6888
rect 1440 6856 1480 6888
rect 1512 6856 1552 6888
rect 1584 6856 1624 6888
rect 1656 6856 1696 6888
rect 1728 6856 1768 6888
rect 1800 6856 1840 6888
rect 1872 6856 1912 6888
rect 1944 6856 1984 6888
rect 2016 6856 2056 6888
rect 2088 6856 2128 6888
rect 2160 6856 2200 6888
rect 2232 6856 2272 6888
rect 2304 6856 2344 6888
rect 2376 6856 2416 6888
rect 2448 6856 2488 6888
rect 2520 6856 2560 6888
rect 2592 6856 2632 6888
rect 2664 6856 2704 6888
rect 2736 6856 2776 6888
rect 2808 6856 2848 6888
rect 2880 6856 2920 6888
rect 2952 6856 2992 6888
rect 3024 6856 3064 6888
rect 3096 6856 3136 6888
rect 3168 6856 3208 6888
rect 3240 6856 3280 6888
rect 3312 6856 3352 6888
rect 3384 6856 3424 6888
rect 3456 6856 3496 6888
rect 3528 6856 3568 6888
rect 3600 6856 3640 6888
rect 3672 6856 3712 6888
rect 3744 6856 3784 6888
rect 3816 6856 3856 6888
rect 3888 6856 3928 6888
rect 3960 6856 4000 6888
rect 0 6800 4000 6856
rect 0 6544 4000 6600
rect 0 6512 40 6544
rect 72 6512 112 6544
rect 144 6512 184 6544
rect 216 6512 256 6544
rect 288 6512 328 6544
rect 360 6512 400 6544
rect 432 6512 472 6544
rect 504 6512 544 6544
rect 576 6512 616 6544
rect 648 6512 688 6544
rect 720 6512 760 6544
rect 792 6512 832 6544
rect 864 6512 904 6544
rect 936 6512 976 6544
rect 1008 6512 1048 6544
rect 1080 6512 1120 6544
rect 1152 6512 1192 6544
rect 1224 6512 1264 6544
rect 1296 6512 1336 6544
rect 1368 6512 1408 6544
rect 1440 6512 1480 6544
rect 1512 6512 1552 6544
rect 1584 6512 1624 6544
rect 1656 6512 1696 6544
rect 1728 6512 1768 6544
rect 1800 6512 1840 6544
rect 1872 6512 1912 6544
rect 1944 6512 1984 6544
rect 2016 6512 2056 6544
rect 2088 6512 2128 6544
rect 2160 6512 2200 6544
rect 2232 6512 2272 6544
rect 2304 6512 2344 6544
rect 2376 6512 2416 6544
rect 2448 6512 2488 6544
rect 2520 6512 2560 6544
rect 2592 6512 2632 6544
rect 2664 6512 2704 6544
rect 2736 6512 2776 6544
rect 2808 6512 2848 6544
rect 2880 6512 2920 6544
rect 2952 6512 2992 6544
rect 3024 6512 3064 6544
rect 3096 6512 3136 6544
rect 3168 6512 3208 6544
rect 3240 6512 3280 6544
rect 3312 6512 3352 6544
rect 3384 6512 3424 6544
rect 3456 6512 3496 6544
rect 3528 6512 3568 6544
rect 3600 6512 3640 6544
rect 3672 6512 3712 6544
rect 3744 6512 3784 6544
rect 3816 6512 3856 6544
rect 3888 6512 3928 6544
rect 3960 6512 4000 6544
rect 0 6472 4000 6512
rect 0 6440 40 6472
rect 72 6440 112 6472
rect 144 6440 184 6472
rect 216 6440 256 6472
rect 288 6440 328 6472
rect 360 6440 400 6472
rect 432 6440 472 6472
rect 504 6440 544 6472
rect 576 6440 616 6472
rect 648 6440 688 6472
rect 720 6440 760 6472
rect 792 6440 832 6472
rect 864 6440 904 6472
rect 936 6440 976 6472
rect 1008 6440 1048 6472
rect 1080 6440 1120 6472
rect 1152 6440 1192 6472
rect 1224 6440 1264 6472
rect 1296 6440 1336 6472
rect 1368 6440 1408 6472
rect 1440 6440 1480 6472
rect 1512 6440 1552 6472
rect 1584 6440 1624 6472
rect 1656 6440 1696 6472
rect 1728 6440 1768 6472
rect 1800 6440 1840 6472
rect 1872 6440 1912 6472
rect 1944 6440 1984 6472
rect 2016 6440 2056 6472
rect 2088 6440 2128 6472
rect 2160 6440 2200 6472
rect 2232 6440 2272 6472
rect 2304 6440 2344 6472
rect 2376 6440 2416 6472
rect 2448 6440 2488 6472
rect 2520 6440 2560 6472
rect 2592 6440 2632 6472
rect 2664 6440 2704 6472
rect 2736 6440 2776 6472
rect 2808 6440 2848 6472
rect 2880 6440 2920 6472
rect 2952 6440 2992 6472
rect 3024 6440 3064 6472
rect 3096 6440 3136 6472
rect 3168 6440 3208 6472
rect 3240 6440 3280 6472
rect 3312 6440 3352 6472
rect 3384 6440 3424 6472
rect 3456 6440 3496 6472
rect 3528 6440 3568 6472
rect 3600 6440 3640 6472
rect 3672 6440 3712 6472
rect 3744 6440 3784 6472
rect 3816 6440 3856 6472
rect 3888 6440 3928 6472
rect 3960 6440 4000 6472
rect 0 6400 4000 6440
rect 0 6368 40 6400
rect 72 6368 112 6400
rect 144 6368 184 6400
rect 216 6368 256 6400
rect 288 6368 328 6400
rect 360 6368 400 6400
rect 432 6368 472 6400
rect 504 6368 544 6400
rect 576 6368 616 6400
rect 648 6368 688 6400
rect 720 6368 760 6400
rect 792 6368 832 6400
rect 864 6368 904 6400
rect 936 6368 976 6400
rect 1008 6368 1048 6400
rect 1080 6368 1120 6400
rect 1152 6368 1192 6400
rect 1224 6368 1264 6400
rect 1296 6368 1336 6400
rect 1368 6368 1408 6400
rect 1440 6368 1480 6400
rect 1512 6368 1552 6400
rect 1584 6368 1624 6400
rect 1656 6368 1696 6400
rect 1728 6368 1768 6400
rect 1800 6368 1840 6400
rect 1872 6368 1912 6400
rect 1944 6368 1984 6400
rect 2016 6368 2056 6400
rect 2088 6368 2128 6400
rect 2160 6368 2200 6400
rect 2232 6368 2272 6400
rect 2304 6368 2344 6400
rect 2376 6368 2416 6400
rect 2448 6368 2488 6400
rect 2520 6368 2560 6400
rect 2592 6368 2632 6400
rect 2664 6368 2704 6400
rect 2736 6368 2776 6400
rect 2808 6368 2848 6400
rect 2880 6368 2920 6400
rect 2952 6368 2992 6400
rect 3024 6368 3064 6400
rect 3096 6368 3136 6400
rect 3168 6368 3208 6400
rect 3240 6368 3280 6400
rect 3312 6368 3352 6400
rect 3384 6368 3424 6400
rect 3456 6368 3496 6400
rect 3528 6368 3568 6400
rect 3600 6368 3640 6400
rect 3672 6368 3712 6400
rect 3744 6368 3784 6400
rect 3816 6368 3856 6400
rect 3888 6368 3928 6400
rect 3960 6368 4000 6400
rect 0 6328 4000 6368
rect 0 6296 40 6328
rect 72 6296 112 6328
rect 144 6296 184 6328
rect 216 6296 256 6328
rect 288 6296 328 6328
rect 360 6296 400 6328
rect 432 6296 472 6328
rect 504 6296 544 6328
rect 576 6296 616 6328
rect 648 6296 688 6328
rect 720 6296 760 6328
rect 792 6296 832 6328
rect 864 6296 904 6328
rect 936 6296 976 6328
rect 1008 6296 1048 6328
rect 1080 6296 1120 6328
rect 1152 6296 1192 6328
rect 1224 6296 1264 6328
rect 1296 6296 1336 6328
rect 1368 6296 1408 6328
rect 1440 6296 1480 6328
rect 1512 6296 1552 6328
rect 1584 6296 1624 6328
rect 1656 6296 1696 6328
rect 1728 6296 1768 6328
rect 1800 6296 1840 6328
rect 1872 6296 1912 6328
rect 1944 6296 1984 6328
rect 2016 6296 2056 6328
rect 2088 6296 2128 6328
rect 2160 6296 2200 6328
rect 2232 6296 2272 6328
rect 2304 6296 2344 6328
rect 2376 6296 2416 6328
rect 2448 6296 2488 6328
rect 2520 6296 2560 6328
rect 2592 6296 2632 6328
rect 2664 6296 2704 6328
rect 2736 6296 2776 6328
rect 2808 6296 2848 6328
rect 2880 6296 2920 6328
rect 2952 6296 2992 6328
rect 3024 6296 3064 6328
rect 3096 6296 3136 6328
rect 3168 6296 3208 6328
rect 3240 6296 3280 6328
rect 3312 6296 3352 6328
rect 3384 6296 3424 6328
rect 3456 6296 3496 6328
rect 3528 6296 3568 6328
rect 3600 6296 3640 6328
rect 3672 6296 3712 6328
rect 3744 6296 3784 6328
rect 3816 6296 3856 6328
rect 3888 6296 3928 6328
rect 3960 6296 4000 6328
rect 0 6256 4000 6296
rect 0 6224 40 6256
rect 72 6224 112 6256
rect 144 6224 184 6256
rect 216 6224 256 6256
rect 288 6224 328 6256
rect 360 6224 400 6256
rect 432 6224 472 6256
rect 504 6224 544 6256
rect 576 6224 616 6256
rect 648 6224 688 6256
rect 720 6224 760 6256
rect 792 6224 832 6256
rect 864 6224 904 6256
rect 936 6224 976 6256
rect 1008 6224 1048 6256
rect 1080 6224 1120 6256
rect 1152 6224 1192 6256
rect 1224 6224 1264 6256
rect 1296 6224 1336 6256
rect 1368 6224 1408 6256
rect 1440 6224 1480 6256
rect 1512 6224 1552 6256
rect 1584 6224 1624 6256
rect 1656 6224 1696 6256
rect 1728 6224 1768 6256
rect 1800 6224 1840 6256
rect 1872 6224 1912 6256
rect 1944 6224 1984 6256
rect 2016 6224 2056 6256
rect 2088 6224 2128 6256
rect 2160 6224 2200 6256
rect 2232 6224 2272 6256
rect 2304 6224 2344 6256
rect 2376 6224 2416 6256
rect 2448 6224 2488 6256
rect 2520 6224 2560 6256
rect 2592 6224 2632 6256
rect 2664 6224 2704 6256
rect 2736 6224 2776 6256
rect 2808 6224 2848 6256
rect 2880 6224 2920 6256
rect 2952 6224 2992 6256
rect 3024 6224 3064 6256
rect 3096 6224 3136 6256
rect 3168 6224 3208 6256
rect 3240 6224 3280 6256
rect 3312 6224 3352 6256
rect 3384 6224 3424 6256
rect 3456 6224 3496 6256
rect 3528 6224 3568 6256
rect 3600 6224 3640 6256
rect 3672 6224 3712 6256
rect 3744 6224 3784 6256
rect 3816 6224 3856 6256
rect 3888 6224 3928 6256
rect 3960 6224 4000 6256
rect 0 6184 4000 6224
rect 0 6152 40 6184
rect 72 6152 112 6184
rect 144 6152 184 6184
rect 216 6152 256 6184
rect 288 6152 328 6184
rect 360 6152 400 6184
rect 432 6152 472 6184
rect 504 6152 544 6184
rect 576 6152 616 6184
rect 648 6152 688 6184
rect 720 6152 760 6184
rect 792 6152 832 6184
rect 864 6152 904 6184
rect 936 6152 976 6184
rect 1008 6152 1048 6184
rect 1080 6152 1120 6184
rect 1152 6152 1192 6184
rect 1224 6152 1264 6184
rect 1296 6152 1336 6184
rect 1368 6152 1408 6184
rect 1440 6152 1480 6184
rect 1512 6152 1552 6184
rect 1584 6152 1624 6184
rect 1656 6152 1696 6184
rect 1728 6152 1768 6184
rect 1800 6152 1840 6184
rect 1872 6152 1912 6184
rect 1944 6152 1984 6184
rect 2016 6152 2056 6184
rect 2088 6152 2128 6184
rect 2160 6152 2200 6184
rect 2232 6152 2272 6184
rect 2304 6152 2344 6184
rect 2376 6152 2416 6184
rect 2448 6152 2488 6184
rect 2520 6152 2560 6184
rect 2592 6152 2632 6184
rect 2664 6152 2704 6184
rect 2736 6152 2776 6184
rect 2808 6152 2848 6184
rect 2880 6152 2920 6184
rect 2952 6152 2992 6184
rect 3024 6152 3064 6184
rect 3096 6152 3136 6184
rect 3168 6152 3208 6184
rect 3240 6152 3280 6184
rect 3312 6152 3352 6184
rect 3384 6152 3424 6184
rect 3456 6152 3496 6184
rect 3528 6152 3568 6184
rect 3600 6152 3640 6184
rect 3672 6152 3712 6184
rect 3744 6152 3784 6184
rect 3816 6152 3856 6184
rect 3888 6152 3928 6184
rect 3960 6152 4000 6184
rect 0 6112 4000 6152
rect 0 6080 40 6112
rect 72 6080 112 6112
rect 144 6080 184 6112
rect 216 6080 256 6112
rect 288 6080 328 6112
rect 360 6080 400 6112
rect 432 6080 472 6112
rect 504 6080 544 6112
rect 576 6080 616 6112
rect 648 6080 688 6112
rect 720 6080 760 6112
rect 792 6080 832 6112
rect 864 6080 904 6112
rect 936 6080 976 6112
rect 1008 6080 1048 6112
rect 1080 6080 1120 6112
rect 1152 6080 1192 6112
rect 1224 6080 1264 6112
rect 1296 6080 1336 6112
rect 1368 6080 1408 6112
rect 1440 6080 1480 6112
rect 1512 6080 1552 6112
rect 1584 6080 1624 6112
rect 1656 6080 1696 6112
rect 1728 6080 1768 6112
rect 1800 6080 1840 6112
rect 1872 6080 1912 6112
rect 1944 6080 1984 6112
rect 2016 6080 2056 6112
rect 2088 6080 2128 6112
rect 2160 6080 2200 6112
rect 2232 6080 2272 6112
rect 2304 6080 2344 6112
rect 2376 6080 2416 6112
rect 2448 6080 2488 6112
rect 2520 6080 2560 6112
rect 2592 6080 2632 6112
rect 2664 6080 2704 6112
rect 2736 6080 2776 6112
rect 2808 6080 2848 6112
rect 2880 6080 2920 6112
rect 2952 6080 2992 6112
rect 3024 6080 3064 6112
rect 3096 6080 3136 6112
rect 3168 6080 3208 6112
rect 3240 6080 3280 6112
rect 3312 6080 3352 6112
rect 3384 6080 3424 6112
rect 3456 6080 3496 6112
rect 3528 6080 3568 6112
rect 3600 6080 3640 6112
rect 3672 6080 3712 6112
rect 3744 6080 3784 6112
rect 3816 6080 3856 6112
rect 3888 6080 3928 6112
rect 3960 6080 4000 6112
rect 0 6040 4000 6080
rect 0 6008 40 6040
rect 72 6008 112 6040
rect 144 6008 184 6040
rect 216 6008 256 6040
rect 288 6008 328 6040
rect 360 6008 400 6040
rect 432 6008 472 6040
rect 504 6008 544 6040
rect 576 6008 616 6040
rect 648 6008 688 6040
rect 720 6008 760 6040
rect 792 6008 832 6040
rect 864 6008 904 6040
rect 936 6008 976 6040
rect 1008 6008 1048 6040
rect 1080 6008 1120 6040
rect 1152 6008 1192 6040
rect 1224 6008 1264 6040
rect 1296 6008 1336 6040
rect 1368 6008 1408 6040
rect 1440 6008 1480 6040
rect 1512 6008 1552 6040
rect 1584 6008 1624 6040
rect 1656 6008 1696 6040
rect 1728 6008 1768 6040
rect 1800 6008 1840 6040
rect 1872 6008 1912 6040
rect 1944 6008 1984 6040
rect 2016 6008 2056 6040
rect 2088 6008 2128 6040
rect 2160 6008 2200 6040
rect 2232 6008 2272 6040
rect 2304 6008 2344 6040
rect 2376 6008 2416 6040
rect 2448 6008 2488 6040
rect 2520 6008 2560 6040
rect 2592 6008 2632 6040
rect 2664 6008 2704 6040
rect 2736 6008 2776 6040
rect 2808 6008 2848 6040
rect 2880 6008 2920 6040
rect 2952 6008 2992 6040
rect 3024 6008 3064 6040
rect 3096 6008 3136 6040
rect 3168 6008 3208 6040
rect 3240 6008 3280 6040
rect 3312 6008 3352 6040
rect 3384 6008 3424 6040
rect 3456 6008 3496 6040
rect 3528 6008 3568 6040
rect 3600 6008 3640 6040
rect 3672 6008 3712 6040
rect 3744 6008 3784 6040
rect 3816 6008 3856 6040
rect 3888 6008 3928 6040
rect 3960 6008 4000 6040
rect 0 5968 4000 6008
rect 0 5936 40 5968
rect 72 5936 112 5968
rect 144 5936 184 5968
rect 216 5936 256 5968
rect 288 5936 328 5968
rect 360 5936 400 5968
rect 432 5936 472 5968
rect 504 5936 544 5968
rect 576 5936 616 5968
rect 648 5936 688 5968
rect 720 5936 760 5968
rect 792 5936 832 5968
rect 864 5936 904 5968
rect 936 5936 976 5968
rect 1008 5936 1048 5968
rect 1080 5936 1120 5968
rect 1152 5936 1192 5968
rect 1224 5936 1264 5968
rect 1296 5936 1336 5968
rect 1368 5936 1408 5968
rect 1440 5936 1480 5968
rect 1512 5936 1552 5968
rect 1584 5936 1624 5968
rect 1656 5936 1696 5968
rect 1728 5936 1768 5968
rect 1800 5936 1840 5968
rect 1872 5936 1912 5968
rect 1944 5936 1984 5968
rect 2016 5936 2056 5968
rect 2088 5936 2128 5968
rect 2160 5936 2200 5968
rect 2232 5936 2272 5968
rect 2304 5936 2344 5968
rect 2376 5936 2416 5968
rect 2448 5936 2488 5968
rect 2520 5936 2560 5968
rect 2592 5936 2632 5968
rect 2664 5936 2704 5968
rect 2736 5936 2776 5968
rect 2808 5936 2848 5968
rect 2880 5936 2920 5968
rect 2952 5936 2992 5968
rect 3024 5936 3064 5968
rect 3096 5936 3136 5968
rect 3168 5936 3208 5968
rect 3240 5936 3280 5968
rect 3312 5936 3352 5968
rect 3384 5936 3424 5968
rect 3456 5936 3496 5968
rect 3528 5936 3568 5968
rect 3600 5936 3640 5968
rect 3672 5936 3712 5968
rect 3744 5936 3784 5968
rect 3816 5936 3856 5968
rect 3888 5936 3928 5968
rect 3960 5936 4000 5968
rect 0 5896 4000 5936
rect 0 5864 40 5896
rect 72 5864 112 5896
rect 144 5864 184 5896
rect 216 5864 256 5896
rect 288 5864 328 5896
rect 360 5864 400 5896
rect 432 5864 472 5896
rect 504 5864 544 5896
rect 576 5864 616 5896
rect 648 5864 688 5896
rect 720 5864 760 5896
rect 792 5864 832 5896
rect 864 5864 904 5896
rect 936 5864 976 5896
rect 1008 5864 1048 5896
rect 1080 5864 1120 5896
rect 1152 5864 1192 5896
rect 1224 5864 1264 5896
rect 1296 5864 1336 5896
rect 1368 5864 1408 5896
rect 1440 5864 1480 5896
rect 1512 5864 1552 5896
rect 1584 5864 1624 5896
rect 1656 5864 1696 5896
rect 1728 5864 1768 5896
rect 1800 5864 1840 5896
rect 1872 5864 1912 5896
rect 1944 5864 1984 5896
rect 2016 5864 2056 5896
rect 2088 5864 2128 5896
rect 2160 5864 2200 5896
rect 2232 5864 2272 5896
rect 2304 5864 2344 5896
rect 2376 5864 2416 5896
rect 2448 5864 2488 5896
rect 2520 5864 2560 5896
rect 2592 5864 2632 5896
rect 2664 5864 2704 5896
rect 2736 5864 2776 5896
rect 2808 5864 2848 5896
rect 2880 5864 2920 5896
rect 2952 5864 2992 5896
rect 3024 5864 3064 5896
rect 3096 5864 3136 5896
rect 3168 5864 3208 5896
rect 3240 5864 3280 5896
rect 3312 5864 3352 5896
rect 3384 5864 3424 5896
rect 3456 5864 3496 5896
rect 3528 5864 3568 5896
rect 3600 5864 3640 5896
rect 3672 5864 3712 5896
rect 3744 5864 3784 5896
rect 3816 5864 3856 5896
rect 3888 5864 3928 5896
rect 3960 5864 4000 5896
rect 0 5824 4000 5864
rect 0 5792 40 5824
rect 72 5792 112 5824
rect 144 5792 184 5824
rect 216 5792 256 5824
rect 288 5792 328 5824
rect 360 5792 400 5824
rect 432 5792 472 5824
rect 504 5792 544 5824
rect 576 5792 616 5824
rect 648 5792 688 5824
rect 720 5792 760 5824
rect 792 5792 832 5824
rect 864 5792 904 5824
rect 936 5792 976 5824
rect 1008 5792 1048 5824
rect 1080 5792 1120 5824
rect 1152 5792 1192 5824
rect 1224 5792 1264 5824
rect 1296 5792 1336 5824
rect 1368 5792 1408 5824
rect 1440 5792 1480 5824
rect 1512 5792 1552 5824
rect 1584 5792 1624 5824
rect 1656 5792 1696 5824
rect 1728 5792 1768 5824
rect 1800 5792 1840 5824
rect 1872 5792 1912 5824
rect 1944 5792 1984 5824
rect 2016 5792 2056 5824
rect 2088 5792 2128 5824
rect 2160 5792 2200 5824
rect 2232 5792 2272 5824
rect 2304 5792 2344 5824
rect 2376 5792 2416 5824
rect 2448 5792 2488 5824
rect 2520 5792 2560 5824
rect 2592 5792 2632 5824
rect 2664 5792 2704 5824
rect 2736 5792 2776 5824
rect 2808 5792 2848 5824
rect 2880 5792 2920 5824
rect 2952 5792 2992 5824
rect 3024 5792 3064 5824
rect 3096 5792 3136 5824
rect 3168 5792 3208 5824
rect 3240 5792 3280 5824
rect 3312 5792 3352 5824
rect 3384 5792 3424 5824
rect 3456 5792 3496 5824
rect 3528 5792 3568 5824
rect 3600 5792 3640 5824
rect 3672 5792 3712 5824
rect 3744 5792 3784 5824
rect 3816 5792 3856 5824
rect 3888 5792 3928 5824
rect 3960 5792 4000 5824
rect 0 5752 4000 5792
rect 0 5720 40 5752
rect 72 5720 112 5752
rect 144 5720 184 5752
rect 216 5720 256 5752
rect 288 5720 328 5752
rect 360 5720 400 5752
rect 432 5720 472 5752
rect 504 5720 544 5752
rect 576 5720 616 5752
rect 648 5720 688 5752
rect 720 5720 760 5752
rect 792 5720 832 5752
rect 864 5720 904 5752
rect 936 5720 976 5752
rect 1008 5720 1048 5752
rect 1080 5720 1120 5752
rect 1152 5720 1192 5752
rect 1224 5720 1264 5752
rect 1296 5720 1336 5752
rect 1368 5720 1408 5752
rect 1440 5720 1480 5752
rect 1512 5720 1552 5752
rect 1584 5720 1624 5752
rect 1656 5720 1696 5752
rect 1728 5720 1768 5752
rect 1800 5720 1840 5752
rect 1872 5720 1912 5752
rect 1944 5720 1984 5752
rect 2016 5720 2056 5752
rect 2088 5720 2128 5752
rect 2160 5720 2200 5752
rect 2232 5720 2272 5752
rect 2304 5720 2344 5752
rect 2376 5720 2416 5752
rect 2448 5720 2488 5752
rect 2520 5720 2560 5752
rect 2592 5720 2632 5752
rect 2664 5720 2704 5752
rect 2736 5720 2776 5752
rect 2808 5720 2848 5752
rect 2880 5720 2920 5752
rect 2952 5720 2992 5752
rect 3024 5720 3064 5752
rect 3096 5720 3136 5752
rect 3168 5720 3208 5752
rect 3240 5720 3280 5752
rect 3312 5720 3352 5752
rect 3384 5720 3424 5752
rect 3456 5720 3496 5752
rect 3528 5720 3568 5752
rect 3600 5720 3640 5752
rect 3672 5720 3712 5752
rect 3744 5720 3784 5752
rect 3816 5720 3856 5752
rect 3888 5720 3928 5752
rect 3960 5720 4000 5752
rect 0 5680 4000 5720
rect 0 5648 40 5680
rect 72 5648 112 5680
rect 144 5648 184 5680
rect 216 5648 256 5680
rect 288 5648 328 5680
rect 360 5648 400 5680
rect 432 5648 472 5680
rect 504 5648 544 5680
rect 576 5648 616 5680
rect 648 5648 688 5680
rect 720 5648 760 5680
rect 792 5648 832 5680
rect 864 5648 904 5680
rect 936 5648 976 5680
rect 1008 5648 1048 5680
rect 1080 5648 1120 5680
rect 1152 5648 1192 5680
rect 1224 5648 1264 5680
rect 1296 5648 1336 5680
rect 1368 5648 1408 5680
rect 1440 5648 1480 5680
rect 1512 5648 1552 5680
rect 1584 5648 1624 5680
rect 1656 5648 1696 5680
rect 1728 5648 1768 5680
rect 1800 5648 1840 5680
rect 1872 5648 1912 5680
rect 1944 5648 1984 5680
rect 2016 5648 2056 5680
rect 2088 5648 2128 5680
rect 2160 5648 2200 5680
rect 2232 5648 2272 5680
rect 2304 5648 2344 5680
rect 2376 5648 2416 5680
rect 2448 5648 2488 5680
rect 2520 5648 2560 5680
rect 2592 5648 2632 5680
rect 2664 5648 2704 5680
rect 2736 5648 2776 5680
rect 2808 5648 2848 5680
rect 2880 5648 2920 5680
rect 2952 5648 2992 5680
rect 3024 5648 3064 5680
rect 3096 5648 3136 5680
rect 3168 5648 3208 5680
rect 3240 5648 3280 5680
rect 3312 5648 3352 5680
rect 3384 5648 3424 5680
rect 3456 5648 3496 5680
rect 3528 5648 3568 5680
rect 3600 5648 3640 5680
rect 3672 5648 3712 5680
rect 3744 5648 3784 5680
rect 3816 5648 3856 5680
rect 3888 5648 3928 5680
rect 3960 5648 4000 5680
rect 0 5608 4000 5648
rect 0 5576 40 5608
rect 72 5576 112 5608
rect 144 5576 184 5608
rect 216 5576 256 5608
rect 288 5576 328 5608
rect 360 5576 400 5608
rect 432 5576 472 5608
rect 504 5576 544 5608
rect 576 5576 616 5608
rect 648 5576 688 5608
rect 720 5576 760 5608
rect 792 5576 832 5608
rect 864 5576 904 5608
rect 936 5576 976 5608
rect 1008 5576 1048 5608
rect 1080 5576 1120 5608
rect 1152 5576 1192 5608
rect 1224 5576 1264 5608
rect 1296 5576 1336 5608
rect 1368 5576 1408 5608
rect 1440 5576 1480 5608
rect 1512 5576 1552 5608
rect 1584 5576 1624 5608
rect 1656 5576 1696 5608
rect 1728 5576 1768 5608
rect 1800 5576 1840 5608
rect 1872 5576 1912 5608
rect 1944 5576 1984 5608
rect 2016 5576 2056 5608
rect 2088 5576 2128 5608
rect 2160 5576 2200 5608
rect 2232 5576 2272 5608
rect 2304 5576 2344 5608
rect 2376 5576 2416 5608
rect 2448 5576 2488 5608
rect 2520 5576 2560 5608
rect 2592 5576 2632 5608
rect 2664 5576 2704 5608
rect 2736 5576 2776 5608
rect 2808 5576 2848 5608
rect 2880 5576 2920 5608
rect 2952 5576 2992 5608
rect 3024 5576 3064 5608
rect 3096 5576 3136 5608
rect 3168 5576 3208 5608
rect 3240 5576 3280 5608
rect 3312 5576 3352 5608
rect 3384 5576 3424 5608
rect 3456 5576 3496 5608
rect 3528 5576 3568 5608
rect 3600 5576 3640 5608
rect 3672 5576 3712 5608
rect 3744 5576 3784 5608
rect 3816 5576 3856 5608
rect 3888 5576 3928 5608
rect 3960 5576 4000 5608
rect 0 5536 4000 5576
rect 0 5504 40 5536
rect 72 5504 112 5536
rect 144 5504 184 5536
rect 216 5504 256 5536
rect 288 5504 328 5536
rect 360 5504 400 5536
rect 432 5504 472 5536
rect 504 5504 544 5536
rect 576 5504 616 5536
rect 648 5504 688 5536
rect 720 5504 760 5536
rect 792 5504 832 5536
rect 864 5504 904 5536
rect 936 5504 976 5536
rect 1008 5504 1048 5536
rect 1080 5504 1120 5536
rect 1152 5504 1192 5536
rect 1224 5504 1264 5536
rect 1296 5504 1336 5536
rect 1368 5504 1408 5536
rect 1440 5504 1480 5536
rect 1512 5504 1552 5536
rect 1584 5504 1624 5536
rect 1656 5504 1696 5536
rect 1728 5504 1768 5536
rect 1800 5504 1840 5536
rect 1872 5504 1912 5536
rect 1944 5504 1984 5536
rect 2016 5504 2056 5536
rect 2088 5504 2128 5536
rect 2160 5504 2200 5536
rect 2232 5504 2272 5536
rect 2304 5504 2344 5536
rect 2376 5504 2416 5536
rect 2448 5504 2488 5536
rect 2520 5504 2560 5536
rect 2592 5504 2632 5536
rect 2664 5504 2704 5536
rect 2736 5504 2776 5536
rect 2808 5504 2848 5536
rect 2880 5504 2920 5536
rect 2952 5504 2992 5536
rect 3024 5504 3064 5536
rect 3096 5504 3136 5536
rect 3168 5504 3208 5536
rect 3240 5504 3280 5536
rect 3312 5504 3352 5536
rect 3384 5504 3424 5536
rect 3456 5504 3496 5536
rect 3528 5504 3568 5536
rect 3600 5504 3640 5536
rect 3672 5504 3712 5536
rect 3744 5504 3784 5536
rect 3816 5504 3856 5536
rect 3888 5504 3928 5536
rect 3960 5504 4000 5536
rect 0 5464 4000 5504
rect 0 5432 40 5464
rect 72 5432 112 5464
rect 144 5432 184 5464
rect 216 5432 256 5464
rect 288 5432 328 5464
rect 360 5432 400 5464
rect 432 5432 472 5464
rect 504 5432 544 5464
rect 576 5432 616 5464
rect 648 5432 688 5464
rect 720 5432 760 5464
rect 792 5432 832 5464
rect 864 5432 904 5464
rect 936 5432 976 5464
rect 1008 5432 1048 5464
rect 1080 5432 1120 5464
rect 1152 5432 1192 5464
rect 1224 5432 1264 5464
rect 1296 5432 1336 5464
rect 1368 5432 1408 5464
rect 1440 5432 1480 5464
rect 1512 5432 1552 5464
rect 1584 5432 1624 5464
rect 1656 5432 1696 5464
rect 1728 5432 1768 5464
rect 1800 5432 1840 5464
rect 1872 5432 1912 5464
rect 1944 5432 1984 5464
rect 2016 5432 2056 5464
rect 2088 5432 2128 5464
rect 2160 5432 2200 5464
rect 2232 5432 2272 5464
rect 2304 5432 2344 5464
rect 2376 5432 2416 5464
rect 2448 5432 2488 5464
rect 2520 5432 2560 5464
rect 2592 5432 2632 5464
rect 2664 5432 2704 5464
rect 2736 5432 2776 5464
rect 2808 5432 2848 5464
rect 2880 5432 2920 5464
rect 2952 5432 2992 5464
rect 3024 5432 3064 5464
rect 3096 5432 3136 5464
rect 3168 5432 3208 5464
rect 3240 5432 3280 5464
rect 3312 5432 3352 5464
rect 3384 5432 3424 5464
rect 3456 5432 3496 5464
rect 3528 5432 3568 5464
rect 3600 5432 3640 5464
rect 3672 5432 3712 5464
rect 3744 5432 3784 5464
rect 3816 5432 3856 5464
rect 3888 5432 3928 5464
rect 3960 5432 4000 5464
rect 0 5392 4000 5432
rect 0 5360 40 5392
rect 72 5360 112 5392
rect 144 5360 184 5392
rect 216 5360 256 5392
rect 288 5360 328 5392
rect 360 5360 400 5392
rect 432 5360 472 5392
rect 504 5360 544 5392
rect 576 5360 616 5392
rect 648 5360 688 5392
rect 720 5360 760 5392
rect 792 5360 832 5392
rect 864 5360 904 5392
rect 936 5360 976 5392
rect 1008 5360 1048 5392
rect 1080 5360 1120 5392
rect 1152 5360 1192 5392
rect 1224 5360 1264 5392
rect 1296 5360 1336 5392
rect 1368 5360 1408 5392
rect 1440 5360 1480 5392
rect 1512 5360 1552 5392
rect 1584 5360 1624 5392
rect 1656 5360 1696 5392
rect 1728 5360 1768 5392
rect 1800 5360 1840 5392
rect 1872 5360 1912 5392
rect 1944 5360 1984 5392
rect 2016 5360 2056 5392
rect 2088 5360 2128 5392
rect 2160 5360 2200 5392
rect 2232 5360 2272 5392
rect 2304 5360 2344 5392
rect 2376 5360 2416 5392
rect 2448 5360 2488 5392
rect 2520 5360 2560 5392
rect 2592 5360 2632 5392
rect 2664 5360 2704 5392
rect 2736 5360 2776 5392
rect 2808 5360 2848 5392
rect 2880 5360 2920 5392
rect 2952 5360 2992 5392
rect 3024 5360 3064 5392
rect 3096 5360 3136 5392
rect 3168 5360 3208 5392
rect 3240 5360 3280 5392
rect 3312 5360 3352 5392
rect 3384 5360 3424 5392
rect 3456 5360 3496 5392
rect 3528 5360 3568 5392
rect 3600 5360 3640 5392
rect 3672 5360 3712 5392
rect 3744 5360 3784 5392
rect 3816 5360 3856 5392
rect 3888 5360 3928 5392
rect 3960 5360 4000 5392
rect 0 5320 4000 5360
rect 0 5288 40 5320
rect 72 5288 112 5320
rect 144 5288 184 5320
rect 216 5288 256 5320
rect 288 5288 328 5320
rect 360 5288 400 5320
rect 432 5288 472 5320
rect 504 5288 544 5320
rect 576 5288 616 5320
rect 648 5288 688 5320
rect 720 5288 760 5320
rect 792 5288 832 5320
rect 864 5288 904 5320
rect 936 5288 976 5320
rect 1008 5288 1048 5320
rect 1080 5288 1120 5320
rect 1152 5288 1192 5320
rect 1224 5288 1264 5320
rect 1296 5288 1336 5320
rect 1368 5288 1408 5320
rect 1440 5288 1480 5320
rect 1512 5288 1552 5320
rect 1584 5288 1624 5320
rect 1656 5288 1696 5320
rect 1728 5288 1768 5320
rect 1800 5288 1840 5320
rect 1872 5288 1912 5320
rect 1944 5288 1984 5320
rect 2016 5288 2056 5320
rect 2088 5288 2128 5320
rect 2160 5288 2200 5320
rect 2232 5288 2272 5320
rect 2304 5288 2344 5320
rect 2376 5288 2416 5320
rect 2448 5288 2488 5320
rect 2520 5288 2560 5320
rect 2592 5288 2632 5320
rect 2664 5288 2704 5320
rect 2736 5288 2776 5320
rect 2808 5288 2848 5320
rect 2880 5288 2920 5320
rect 2952 5288 2992 5320
rect 3024 5288 3064 5320
rect 3096 5288 3136 5320
rect 3168 5288 3208 5320
rect 3240 5288 3280 5320
rect 3312 5288 3352 5320
rect 3384 5288 3424 5320
rect 3456 5288 3496 5320
rect 3528 5288 3568 5320
rect 3600 5288 3640 5320
rect 3672 5288 3712 5320
rect 3744 5288 3784 5320
rect 3816 5288 3856 5320
rect 3888 5288 3928 5320
rect 3960 5288 4000 5320
rect 0 5248 4000 5288
rect 0 5216 40 5248
rect 72 5216 112 5248
rect 144 5216 184 5248
rect 216 5216 256 5248
rect 288 5216 328 5248
rect 360 5216 400 5248
rect 432 5216 472 5248
rect 504 5216 544 5248
rect 576 5216 616 5248
rect 648 5216 688 5248
rect 720 5216 760 5248
rect 792 5216 832 5248
rect 864 5216 904 5248
rect 936 5216 976 5248
rect 1008 5216 1048 5248
rect 1080 5216 1120 5248
rect 1152 5216 1192 5248
rect 1224 5216 1264 5248
rect 1296 5216 1336 5248
rect 1368 5216 1408 5248
rect 1440 5216 1480 5248
rect 1512 5216 1552 5248
rect 1584 5216 1624 5248
rect 1656 5216 1696 5248
rect 1728 5216 1768 5248
rect 1800 5216 1840 5248
rect 1872 5216 1912 5248
rect 1944 5216 1984 5248
rect 2016 5216 2056 5248
rect 2088 5216 2128 5248
rect 2160 5216 2200 5248
rect 2232 5216 2272 5248
rect 2304 5216 2344 5248
rect 2376 5216 2416 5248
rect 2448 5216 2488 5248
rect 2520 5216 2560 5248
rect 2592 5216 2632 5248
rect 2664 5216 2704 5248
rect 2736 5216 2776 5248
rect 2808 5216 2848 5248
rect 2880 5216 2920 5248
rect 2952 5216 2992 5248
rect 3024 5216 3064 5248
rect 3096 5216 3136 5248
rect 3168 5216 3208 5248
rect 3240 5216 3280 5248
rect 3312 5216 3352 5248
rect 3384 5216 3424 5248
rect 3456 5216 3496 5248
rect 3528 5216 3568 5248
rect 3600 5216 3640 5248
rect 3672 5216 3712 5248
rect 3744 5216 3784 5248
rect 3816 5216 3856 5248
rect 3888 5216 3928 5248
rect 3960 5216 4000 5248
rect 0 5176 4000 5216
rect 0 5144 40 5176
rect 72 5144 112 5176
rect 144 5144 184 5176
rect 216 5144 256 5176
rect 288 5144 328 5176
rect 360 5144 400 5176
rect 432 5144 472 5176
rect 504 5144 544 5176
rect 576 5144 616 5176
rect 648 5144 688 5176
rect 720 5144 760 5176
rect 792 5144 832 5176
rect 864 5144 904 5176
rect 936 5144 976 5176
rect 1008 5144 1048 5176
rect 1080 5144 1120 5176
rect 1152 5144 1192 5176
rect 1224 5144 1264 5176
rect 1296 5144 1336 5176
rect 1368 5144 1408 5176
rect 1440 5144 1480 5176
rect 1512 5144 1552 5176
rect 1584 5144 1624 5176
rect 1656 5144 1696 5176
rect 1728 5144 1768 5176
rect 1800 5144 1840 5176
rect 1872 5144 1912 5176
rect 1944 5144 1984 5176
rect 2016 5144 2056 5176
rect 2088 5144 2128 5176
rect 2160 5144 2200 5176
rect 2232 5144 2272 5176
rect 2304 5144 2344 5176
rect 2376 5144 2416 5176
rect 2448 5144 2488 5176
rect 2520 5144 2560 5176
rect 2592 5144 2632 5176
rect 2664 5144 2704 5176
rect 2736 5144 2776 5176
rect 2808 5144 2848 5176
rect 2880 5144 2920 5176
rect 2952 5144 2992 5176
rect 3024 5144 3064 5176
rect 3096 5144 3136 5176
rect 3168 5144 3208 5176
rect 3240 5144 3280 5176
rect 3312 5144 3352 5176
rect 3384 5144 3424 5176
rect 3456 5144 3496 5176
rect 3528 5144 3568 5176
rect 3600 5144 3640 5176
rect 3672 5144 3712 5176
rect 3744 5144 3784 5176
rect 3816 5144 3856 5176
rect 3888 5144 3928 5176
rect 3960 5144 4000 5176
rect 0 5104 4000 5144
rect 0 5072 40 5104
rect 72 5072 112 5104
rect 144 5072 184 5104
rect 216 5072 256 5104
rect 288 5072 328 5104
rect 360 5072 400 5104
rect 432 5072 472 5104
rect 504 5072 544 5104
rect 576 5072 616 5104
rect 648 5072 688 5104
rect 720 5072 760 5104
rect 792 5072 832 5104
rect 864 5072 904 5104
rect 936 5072 976 5104
rect 1008 5072 1048 5104
rect 1080 5072 1120 5104
rect 1152 5072 1192 5104
rect 1224 5072 1264 5104
rect 1296 5072 1336 5104
rect 1368 5072 1408 5104
rect 1440 5072 1480 5104
rect 1512 5072 1552 5104
rect 1584 5072 1624 5104
rect 1656 5072 1696 5104
rect 1728 5072 1768 5104
rect 1800 5072 1840 5104
rect 1872 5072 1912 5104
rect 1944 5072 1984 5104
rect 2016 5072 2056 5104
rect 2088 5072 2128 5104
rect 2160 5072 2200 5104
rect 2232 5072 2272 5104
rect 2304 5072 2344 5104
rect 2376 5072 2416 5104
rect 2448 5072 2488 5104
rect 2520 5072 2560 5104
rect 2592 5072 2632 5104
rect 2664 5072 2704 5104
rect 2736 5072 2776 5104
rect 2808 5072 2848 5104
rect 2880 5072 2920 5104
rect 2952 5072 2992 5104
rect 3024 5072 3064 5104
rect 3096 5072 3136 5104
rect 3168 5072 3208 5104
rect 3240 5072 3280 5104
rect 3312 5072 3352 5104
rect 3384 5072 3424 5104
rect 3456 5072 3496 5104
rect 3528 5072 3568 5104
rect 3600 5072 3640 5104
rect 3672 5072 3712 5104
rect 3744 5072 3784 5104
rect 3816 5072 3856 5104
rect 3888 5072 3928 5104
rect 3960 5072 4000 5104
rect 0 5032 4000 5072
rect 0 5000 40 5032
rect 72 5000 112 5032
rect 144 5000 184 5032
rect 216 5000 256 5032
rect 288 5000 328 5032
rect 360 5000 400 5032
rect 432 5000 472 5032
rect 504 5000 544 5032
rect 576 5000 616 5032
rect 648 5000 688 5032
rect 720 5000 760 5032
rect 792 5000 832 5032
rect 864 5000 904 5032
rect 936 5000 976 5032
rect 1008 5000 1048 5032
rect 1080 5000 1120 5032
rect 1152 5000 1192 5032
rect 1224 5000 1264 5032
rect 1296 5000 1336 5032
rect 1368 5000 1408 5032
rect 1440 5000 1480 5032
rect 1512 5000 1552 5032
rect 1584 5000 1624 5032
rect 1656 5000 1696 5032
rect 1728 5000 1768 5032
rect 1800 5000 1840 5032
rect 1872 5000 1912 5032
rect 1944 5000 1984 5032
rect 2016 5000 2056 5032
rect 2088 5000 2128 5032
rect 2160 5000 2200 5032
rect 2232 5000 2272 5032
rect 2304 5000 2344 5032
rect 2376 5000 2416 5032
rect 2448 5000 2488 5032
rect 2520 5000 2560 5032
rect 2592 5000 2632 5032
rect 2664 5000 2704 5032
rect 2736 5000 2776 5032
rect 2808 5000 2848 5032
rect 2880 5000 2920 5032
rect 2952 5000 2992 5032
rect 3024 5000 3064 5032
rect 3096 5000 3136 5032
rect 3168 5000 3208 5032
rect 3240 5000 3280 5032
rect 3312 5000 3352 5032
rect 3384 5000 3424 5032
rect 3456 5000 3496 5032
rect 3528 5000 3568 5032
rect 3600 5000 3640 5032
rect 3672 5000 3712 5032
rect 3744 5000 3784 5032
rect 3816 5000 3856 5032
rect 3888 5000 3928 5032
rect 3960 5000 4000 5032
rect 0 4960 4000 5000
rect 0 4928 40 4960
rect 72 4928 112 4960
rect 144 4928 184 4960
rect 216 4928 256 4960
rect 288 4928 328 4960
rect 360 4928 400 4960
rect 432 4928 472 4960
rect 504 4928 544 4960
rect 576 4928 616 4960
rect 648 4928 688 4960
rect 720 4928 760 4960
rect 792 4928 832 4960
rect 864 4928 904 4960
rect 936 4928 976 4960
rect 1008 4928 1048 4960
rect 1080 4928 1120 4960
rect 1152 4928 1192 4960
rect 1224 4928 1264 4960
rect 1296 4928 1336 4960
rect 1368 4928 1408 4960
rect 1440 4928 1480 4960
rect 1512 4928 1552 4960
rect 1584 4928 1624 4960
rect 1656 4928 1696 4960
rect 1728 4928 1768 4960
rect 1800 4928 1840 4960
rect 1872 4928 1912 4960
rect 1944 4928 1984 4960
rect 2016 4928 2056 4960
rect 2088 4928 2128 4960
rect 2160 4928 2200 4960
rect 2232 4928 2272 4960
rect 2304 4928 2344 4960
rect 2376 4928 2416 4960
rect 2448 4928 2488 4960
rect 2520 4928 2560 4960
rect 2592 4928 2632 4960
rect 2664 4928 2704 4960
rect 2736 4928 2776 4960
rect 2808 4928 2848 4960
rect 2880 4928 2920 4960
rect 2952 4928 2992 4960
rect 3024 4928 3064 4960
rect 3096 4928 3136 4960
rect 3168 4928 3208 4960
rect 3240 4928 3280 4960
rect 3312 4928 3352 4960
rect 3384 4928 3424 4960
rect 3456 4928 3496 4960
rect 3528 4928 3568 4960
rect 3600 4928 3640 4960
rect 3672 4928 3712 4960
rect 3744 4928 3784 4960
rect 3816 4928 3856 4960
rect 3888 4928 3928 4960
rect 3960 4928 4000 4960
rect 0 4888 4000 4928
rect 0 4856 40 4888
rect 72 4856 112 4888
rect 144 4856 184 4888
rect 216 4856 256 4888
rect 288 4856 328 4888
rect 360 4856 400 4888
rect 432 4856 472 4888
rect 504 4856 544 4888
rect 576 4856 616 4888
rect 648 4856 688 4888
rect 720 4856 760 4888
rect 792 4856 832 4888
rect 864 4856 904 4888
rect 936 4856 976 4888
rect 1008 4856 1048 4888
rect 1080 4856 1120 4888
rect 1152 4856 1192 4888
rect 1224 4856 1264 4888
rect 1296 4856 1336 4888
rect 1368 4856 1408 4888
rect 1440 4856 1480 4888
rect 1512 4856 1552 4888
rect 1584 4856 1624 4888
rect 1656 4856 1696 4888
rect 1728 4856 1768 4888
rect 1800 4856 1840 4888
rect 1872 4856 1912 4888
rect 1944 4856 1984 4888
rect 2016 4856 2056 4888
rect 2088 4856 2128 4888
rect 2160 4856 2200 4888
rect 2232 4856 2272 4888
rect 2304 4856 2344 4888
rect 2376 4856 2416 4888
rect 2448 4856 2488 4888
rect 2520 4856 2560 4888
rect 2592 4856 2632 4888
rect 2664 4856 2704 4888
rect 2736 4856 2776 4888
rect 2808 4856 2848 4888
rect 2880 4856 2920 4888
rect 2952 4856 2992 4888
rect 3024 4856 3064 4888
rect 3096 4856 3136 4888
rect 3168 4856 3208 4888
rect 3240 4856 3280 4888
rect 3312 4856 3352 4888
rect 3384 4856 3424 4888
rect 3456 4856 3496 4888
rect 3528 4856 3568 4888
rect 3600 4856 3640 4888
rect 3672 4856 3712 4888
rect 3744 4856 3784 4888
rect 3816 4856 3856 4888
rect 3888 4856 3928 4888
rect 3960 4856 4000 4888
rect 0 4816 4000 4856
rect 0 4784 40 4816
rect 72 4784 112 4816
rect 144 4784 184 4816
rect 216 4784 256 4816
rect 288 4784 328 4816
rect 360 4784 400 4816
rect 432 4784 472 4816
rect 504 4784 544 4816
rect 576 4784 616 4816
rect 648 4784 688 4816
rect 720 4784 760 4816
rect 792 4784 832 4816
rect 864 4784 904 4816
rect 936 4784 976 4816
rect 1008 4784 1048 4816
rect 1080 4784 1120 4816
rect 1152 4784 1192 4816
rect 1224 4784 1264 4816
rect 1296 4784 1336 4816
rect 1368 4784 1408 4816
rect 1440 4784 1480 4816
rect 1512 4784 1552 4816
rect 1584 4784 1624 4816
rect 1656 4784 1696 4816
rect 1728 4784 1768 4816
rect 1800 4784 1840 4816
rect 1872 4784 1912 4816
rect 1944 4784 1984 4816
rect 2016 4784 2056 4816
rect 2088 4784 2128 4816
rect 2160 4784 2200 4816
rect 2232 4784 2272 4816
rect 2304 4784 2344 4816
rect 2376 4784 2416 4816
rect 2448 4784 2488 4816
rect 2520 4784 2560 4816
rect 2592 4784 2632 4816
rect 2664 4784 2704 4816
rect 2736 4784 2776 4816
rect 2808 4784 2848 4816
rect 2880 4784 2920 4816
rect 2952 4784 2992 4816
rect 3024 4784 3064 4816
rect 3096 4784 3136 4816
rect 3168 4784 3208 4816
rect 3240 4784 3280 4816
rect 3312 4784 3352 4816
rect 3384 4784 3424 4816
rect 3456 4784 3496 4816
rect 3528 4784 3568 4816
rect 3600 4784 3640 4816
rect 3672 4784 3712 4816
rect 3744 4784 3784 4816
rect 3816 4784 3856 4816
rect 3888 4784 3928 4816
rect 3960 4784 4000 4816
rect 0 4744 4000 4784
rect 0 4712 40 4744
rect 72 4712 112 4744
rect 144 4712 184 4744
rect 216 4712 256 4744
rect 288 4712 328 4744
rect 360 4712 400 4744
rect 432 4712 472 4744
rect 504 4712 544 4744
rect 576 4712 616 4744
rect 648 4712 688 4744
rect 720 4712 760 4744
rect 792 4712 832 4744
rect 864 4712 904 4744
rect 936 4712 976 4744
rect 1008 4712 1048 4744
rect 1080 4712 1120 4744
rect 1152 4712 1192 4744
rect 1224 4712 1264 4744
rect 1296 4712 1336 4744
rect 1368 4712 1408 4744
rect 1440 4712 1480 4744
rect 1512 4712 1552 4744
rect 1584 4712 1624 4744
rect 1656 4712 1696 4744
rect 1728 4712 1768 4744
rect 1800 4712 1840 4744
rect 1872 4712 1912 4744
rect 1944 4712 1984 4744
rect 2016 4712 2056 4744
rect 2088 4712 2128 4744
rect 2160 4712 2200 4744
rect 2232 4712 2272 4744
rect 2304 4712 2344 4744
rect 2376 4712 2416 4744
rect 2448 4712 2488 4744
rect 2520 4712 2560 4744
rect 2592 4712 2632 4744
rect 2664 4712 2704 4744
rect 2736 4712 2776 4744
rect 2808 4712 2848 4744
rect 2880 4712 2920 4744
rect 2952 4712 2992 4744
rect 3024 4712 3064 4744
rect 3096 4712 3136 4744
rect 3168 4712 3208 4744
rect 3240 4712 3280 4744
rect 3312 4712 3352 4744
rect 3384 4712 3424 4744
rect 3456 4712 3496 4744
rect 3528 4712 3568 4744
rect 3600 4712 3640 4744
rect 3672 4712 3712 4744
rect 3744 4712 3784 4744
rect 3816 4712 3856 4744
rect 3888 4712 3928 4744
rect 3960 4712 4000 4744
rect 0 4672 4000 4712
rect 0 4640 40 4672
rect 72 4640 112 4672
rect 144 4640 184 4672
rect 216 4640 256 4672
rect 288 4640 328 4672
rect 360 4640 400 4672
rect 432 4640 472 4672
rect 504 4640 544 4672
rect 576 4640 616 4672
rect 648 4640 688 4672
rect 720 4640 760 4672
rect 792 4640 832 4672
rect 864 4640 904 4672
rect 936 4640 976 4672
rect 1008 4640 1048 4672
rect 1080 4640 1120 4672
rect 1152 4640 1192 4672
rect 1224 4640 1264 4672
rect 1296 4640 1336 4672
rect 1368 4640 1408 4672
rect 1440 4640 1480 4672
rect 1512 4640 1552 4672
rect 1584 4640 1624 4672
rect 1656 4640 1696 4672
rect 1728 4640 1768 4672
rect 1800 4640 1840 4672
rect 1872 4640 1912 4672
rect 1944 4640 1984 4672
rect 2016 4640 2056 4672
rect 2088 4640 2128 4672
rect 2160 4640 2200 4672
rect 2232 4640 2272 4672
rect 2304 4640 2344 4672
rect 2376 4640 2416 4672
rect 2448 4640 2488 4672
rect 2520 4640 2560 4672
rect 2592 4640 2632 4672
rect 2664 4640 2704 4672
rect 2736 4640 2776 4672
rect 2808 4640 2848 4672
rect 2880 4640 2920 4672
rect 2952 4640 2992 4672
rect 3024 4640 3064 4672
rect 3096 4640 3136 4672
rect 3168 4640 3208 4672
rect 3240 4640 3280 4672
rect 3312 4640 3352 4672
rect 3384 4640 3424 4672
rect 3456 4640 3496 4672
rect 3528 4640 3568 4672
rect 3600 4640 3640 4672
rect 3672 4640 3712 4672
rect 3744 4640 3784 4672
rect 3816 4640 3856 4672
rect 3888 4640 3928 4672
rect 3960 4640 4000 4672
rect 0 4600 4000 4640
rect 0 4568 40 4600
rect 72 4568 112 4600
rect 144 4568 184 4600
rect 216 4568 256 4600
rect 288 4568 328 4600
rect 360 4568 400 4600
rect 432 4568 472 4600
rect 504 4568 544 4600
rect 576 4568 616 4600
rect 648 4568 688 4600
rect 720 4568 760 4600
rect 792 4568 832 4600
rect 864 4568 904 4600
rect 936 4568 976 4600
rect 1008 4568 1048 4600
rect 1080 4568 1120 4600
rect 1152 4568 1192 4600
rect 1224 4568 1264 4600
rect 1296 4568 1336 4600
rect 1368 4568 1408 4600
rect 1440 4568 1480 4600
rect 1512 4568 1552 4600
rect 1584 4568 1624 4600
rect 1656 4568 1696 4600
rect 1728 4568 1768 4600
rect 1800 4568 1840 4600
rect 1872 4568 1912 4600
rect 1944 4568 1984 4600
rect 2016 4568 2056 4600
rect 2088 4568 2128 4600
rect 2160 4568 2200 4600
rect 2232 4568 2272 4600
rect 2304 4568 2344 4600
rect 2376 4568 2416 4600
rect 2448 4568 2488 4600
rect 2520 4568 2560 4600
rect 2592 4568 2632 4600
rect 2664 4568 2704 4600
rect 2736 4568 2776 4600
rect 2808 4568 2848 4600
rect 2880 4568 2920 4600
rect 2952 4568 2992 4600
rect 3024 4568 3064 4600
rect 3096 4568 3136 4600
rect 3168 4568 3208 4600
rect 3240 4568 3280 4600
rect 3312 4568 3352 4600
rect 3384 4568 3424 4600
rect 3456 4568 3496 4600
rect 3528 4568 3568 4600
rect 3600 4568 3640 4600
rect 3672 4568 3712 4600
rect 3744 4568 3784 4600
rect 3816 4568 3856 4600
rect 3888 4568 3928 4600
rect 3960 4568 4000 4600
rect 0 4528 4000 4568
rect 0 4496 40 4528
rect 72 4496 112 4528
rect 144 4496 184 4528
rect 216 4496 256 4528
rect 288 4496 328 4528
rect 360 4496 400 4528
rect 432 4496 472 4528
rect 504 4496 544 4528
rect 576 4496 616 4528
rect 648 4496 688 4528
rect 720 4496 760 4528
rect 792 4496 832 4528
rect 864 4496 904 4528
rect 936 4496 976 4528
rect 1008 4496 1048 4528
rect 1080 4496 1120 4528
rect 1152 4496 1192 4528
rect 1224 4496 1264 4528
rect 1296 4496 1336 4528
rect 1368 4496 1408 4528
rect 1440 4496 1480 4528
rect 1512 4496 1552 4528
rect 1584 4496 1624 4528
rect 1656 4496 1696 4528
rect 1728 4496 1768 4528
rect 1800 4496 1840 4528
rect 1872 4496 1912 4528
rect 1944 4496 1984 4528
rect 2016 4496 2056 4528
rect 2088 4496 2128 4528
rect 2160 4496 2200 4528
rect 2232 4496 2272 4528
rect 2304 4496 2344 4528
rect 2376 4496 2416 4528
rect 2448 4496 2488 4528
rect 2520 4496 2560 4528
rect 2592 4496 2632 4528
rect 2664 4496 2704 4528
rect 2736 4496 2776 4528
rect 2808 4496 2848 4528
rect 2880 4496 2920 4528
rect 2952 4496 2992 4528
rect 3024 4496 3064 4528
rect 3096 4496 3136 4528
rect 3168 4496 3208 4528
rect 3240 4496 3280 4528
rect 3312 4496 3352 4528
rect 3384 4496 3424 4528
rect 3456 4496 3496 4528
rect 3528 4496 3568 4528
rect 3600 4496 3640 4528
rect 3672 4496 3712 4528
rect 3744 4496 3784 4528
rect 3816 4496 3856 4528
rect 3888 4496 3928 4528
rect 3960 4496 4000 4528
rect 0 4456 4000 4496
rect 0 4424 40 4456
rect 72 4424 112 4456
rect 144 4424 184 4456
rect 216 4424 256 4456
rect 288 4424 328 4456
rect 360 4424 400 4456
rect 432 4424 472 4456
rect 504 4424 544 4456
rect 576 4424 616 4456
rect 648 4424 688 4456
rect 720 4424 760 4456
rect 792 4424 832 4456
rect 864 4424 904 4456
rect 936 4424 976 4456
rect 1008 4424 1048 4456
rect 1080 4424 1120 4456
rect 1152 4424 1192 4456
rect 1224 4424 1264 4456
rect 1296 4424 1336 4456
rect 1368 4424 1408 4456
rect 1440 4424 1480 4456
rect 1512 4424 1552 4456
rect 1584 4424 1624 4456
rect 1656 4424 1696 4456
rect 1728 4424 1768 4456
rect 1800 4424 1840 4456
rect 1872 4424 1912 4456
rect 1944 4424 1984 4456
rect 2016 4424 2056 4456
rect 2088 4424 2128 4456
rect 2160 4424 2200 4456
rect 2232 4424 2272 4456
rect 2304 4424 2344 4456
rect 2376 4424 2416 4456
rect 2448 4424 2488 4456
rect 2520 4424 2560 4456
rect 2592 4424 2632 4456
rect 2664 4424 2704 4456
rect 2736 4424 2776 4456
rect 2808 4424 2848 4456
rect 2880 4424 2920 4456
rect 2952 4424 2992 4456
rect 3024 4424 3064 4456
rect 3096 4424 3136 4456
rect 3168 4424 3208 4456
rect 3240 4424 3280 4456
rect 3312 4424 3352 4456
rect 3384 4424 3424 4456
rect 3456 4424 3496 4456
rect 3528 4424 3568 4456
rect 3600 4424 3640 4456
rect 3672 4424 3712 4456
rect 3744 4424 3784 4456
rect 3816 4424 3856 4456
rect 3888 4424 3928 4456
rect 3960 4424 4000 4456
rect 0 4384 4000 4424
rect 0 4352 40 4384
rect 72 4352 112 4384
rect 144 4352 184 4384
rect 216 4352 256 4384
rect 288 4352 328 4384
rect 360 4352 400 4384
rect 432 4352 472 4384
rect 504 4352 544 4384
rect 576 4352 616 4384
rect 648 4352 688 4384
rect 720 4352 760 4384
rect 792 4352 832 4384
rect 864 4352 904 4384
rect 936 4352 976 4384
rect 1008 4352 1048 4384
rect 1080 4352 1120 4384
rect 1152 4352 1192 4384
rect 1224 4352 1264 4384
rect 1296 4352 1336 4384
rect 1368 4352 1408 4384
rect 1440 4352 1480 4384
rect 1512 4352 1552 4384
rect 1584 4352 1624 4384
rect 1656 4352 1696 4384
rect 1728 4352 1768 4384
rect 1800 4352 1840 4384
rect 1872 4352 1912 4384
rect 1944 4352 1984 4384
rect 2016 4352 2056 4384
rect 2088 4352 2128 4384
rect 2160 4352 2200 4384
rect 2232 4352 2272 4384
rect 2304 4352 2344 4384
rect 2376 4352 2416 4384
rect 2448 4352 2488 4384
rect 2520 4352 2560 4384
rect 2592 4352 2632 4384
rect 2664 4352 2704 4384
rect 2736 4352 2776 4384
rect 2808 4352 2848 4384
rect 2880 4352 2920 4384
rect 2952 4352 2992 4384
rect 3024 4352 3064 4384
rect 3096 4352 3136 4384
rect 3168 4352 3208 4384
rect 3240 4352 3280 4384
rect 3312 4352 3352 4384
rect 3384 4352 3424 4384
rect 3456 4352 3496 4384
rect 3528 4352 3568 4384
rect 3600 4352 3640 4384
rect 3672 4352 3712 4384
rect 3744 4352 3784 4384
rect 3816 4352 3856 4384
rect 3888 4352 3928 4384
rect 3960 4352 4000 4384
rect 0 4312 4000 4352
rect 0 4280 40 4312
rect 72 4280 112 4312
rect 144 4280 184 4312
rect 216 4280 256 4312
rect 288 4280 328 4312
rect 360 4280 400 4312
rect 432 4280 472 4312
rect 504 4280 544 4312
rect 576 4280 616 4312
rect 648 4280 688 4312
rect 720 4280 760 4312
rect 792 4280 832 4312
rect 864 4280 904 4312
rect 936 4280 976 4312
rect 1008 4280 1048 4312
rect 1080 4280 1120 4312
rect 1152 4280 1192 4312
rect 1224 4280 1264 4312
rect 1296 4280 1336 4312
rect 1368 4280 1408 4312
rect 1440 4280 1480 4312
rect 1512 4280 1552 4312
rect 1584 4280 1624 4312
rect 1656 4280 1696 4312
rect 1728 4280 1768 4312
rect 1800 4280 1840 4312
rect 1872 4280 1912 4312
rect 1944 4280 1984 4312
rect 2016 4280 2056 4312
rect 2088 4280 2128 4312
rect 2160 4280 2200 4312
rect 2232 4280 2272 4312
rect 2304 4280 2344 4312
rect 2376 4280 2416 4312
rect 2448 4280 2488 4312
rect 2520 4280 2560 4312
rect 2592 4280 2632 4312
rect 2664 4280 2704 4312
rect 2736 4280 2776 4312
rect 2808 4280 2848 4312
rect 2880 4280 2920 4312
rect 2952 4280 2992 4312
rect 3024 4280 3064 4312
rect 3096 4280 3136 4312
rect 3168 4280 3208 4312
rect 3240 4280 3280 4312
rect 3312 4280 3352 4312
rect 3384 4280 3424 4312
rect 3456 4280 3496 4312
rect 3528 4280 3568 4312
rect 3600 4280 3640 4312
rect 3672 4280 3712 4312
rect 3744 4280 3784 4312
rect 3816 4280 3856 4312
rect 3888 4280 3928 4312
rect 3960 4280 4000 4312
rect 0 4240 4000 4280
rect 0 4208 40 4240
rect 72 4208 112 4240
rect 144 4208 184 4240
rect 216 4208 256 4240
rect 288 4208 328 4240
rect 360 4208 400 4240
rect 432 4208 472 4240
rect 504 4208 544 4240
rect 576 4208 616 4240
rect 648 4208 688 4240
rect 720 4208 760 4240
rect 792 4208 832 4240
rect 864 4208 904 4240
rect 936 4208 976 4240
rect 1008 4208 1048 4240
rect 1080 4208 1120 4240
rect 1152 4208 1192 4240
rect 1224 4208 1264 4240
rect 1296 4208 1336 4240
rect 1368 4208 1408 4240
rect 1440 4208 1480 4240
rect 1512 4208 1552 4240
rect 1584 4208 1624 4240
rect 1656 4208 1696 4240
rect 1728 4208 1768 4240
rect 1800 4208 1840 4240
rect 1872 4208 1912 4240
rect 1944 4208 1984 4240
rect 2016 4208 2056 4240
rect 2088 4208 2128 4240
rect 2160 4208 2200 4240
rect 2232 4208 2272 4240
rect 2304 4208 2344 4240
rect 2376 4208 2416 4240
rect 2448 4208 2488 4240
rect 2520 4208 2560 4240
rect 2592 4208 2632 4240
rect 2664 4208 2704 4240
rect 2736 4208 2776 4240
rect 2808 4208 2848 4240
rect 2880 4208 2920 4240
rect 2952 4208 2992 4240
rect 3024 4208 3064 4240
rect 3096 4208 3136 4240
rect 3168 4208 3208 4240
rect 3240 4208 3280 4240
rect 3312 4208 3352 4240
rect 3384 4208 3424 4240
rect 3456 4208 3496 4240
rect 3528 4208 3568 4240
rect 3600 4208 3640 4240
rect 3672 4208 3712 4240
rect 3744 4208 3784 4240
rect 3816 4208 3856 4240
rect 3888 4208 3928 4240
rect 3960 4208 4000 4240
rect 0 4168 4000 4208
rect 0 4136 40 4168
rect 72 4136 112 4168
rect 144 4136 184 4168
rect 216 4136 256 4168
rect 288 4136 328 4168
rect 360 4136 400 4168
rect 432 4136 472 4168
rect 504 4136 544 4168
rect 576 4136 616 4168
rect 648 4136 688 4168
rect 720 4136 760 4168
rect 792 4136 832 4168
rect 864 4136 904 4168
rect 936 4136 976 4168
rect 1008 4136 1048 4168
rect 1080 4136 1120 4168
rect 1152 4136 1192 4168
rect 1224 4136 1264 4168
rect 1296 4136 1336 4168
rect 1368 4136 1408 4168
rect 1440 4136 1480 4168
rect 1512 4136 1552 4168
rect 1584 4136 1624 4168
rect 1656 4136 1696 4168
rect 1728 4136 1768 4168
rect 1800 4136 1840 4168
rect 1872 4136 1912 4168
rect 1944 4136 1984 4168
rect 2016 4136 2056 4168
rect 2088 4136 2128 4168
rect 2160 4136 2200 4168
rect 2232 4136 2272 4168
rect 2304 4136 2344 4168
rect 2376 4136 2416 4168
rect 2448 4136 2488 4168
rect 2520 4136 2560 4168
rect 2592 4136 2632 4168
rect 2664 4136 2704 4168
rect 2736 4136 2776 4168
rect 2808 4136 2848 4168
rect 2880 4136 2920 4168
rect 2952 4136 2992 4168
rect 3024 4136 3064 4168
rect 3096 4136 3136 4168
rect 3168 4136 3208 4168
rect 3240 4136 3280 4168
rect 3312 4136 3352 4168
rect 3384 4136 3424 4168
rect 3456 4136 3496 4168
rect 3528 4136 3568 4168
rect 3600 4136 3640 4168
rect 3672 4136 3712 4168
rect 3744 4136 3784 4168
rect 3816 4136 3856 4168
rect 3888 4136 3928 4168
rect 3960 4136 4000 4168
rect 0 4096 4000 4136
rect 0 4064 40 4096
rect 72 4064 112 4096
rect 144 4064 184 4096
rect 216 4064 256 4096
rect 288 4064 328 4096
rect 360 4064 400 4096
rect 432 4064 472 4096
rect 504 4064 544 4096
rect 576 4064 616 4096
rect 648 4064 688 4096
rect 720 4064 760 4096
rect 792 4064 832 4096
rect 864 4064 904 4096
rect 936 4064 976 4096
rect 1008 4064 1048 4096
rect 1080 4064 1120 4096
rect 1152 4064 1192 4096
rect 1224 4064 1264 4096
rect 1296 4064 1336 4096
rect 1368 4064 1408 4096
rect 1440 4064 1480 4096
rect 1512 4064 1552 4096
rect 1584 4064 1624 4096
rect 1656 4064 1696 4096
rect 1728 4064 1768 4096
rect 1800 4064 1840 4096
rect 1872 4064 1912 4096
rect 1944 4064 1984 4096
rect 2016 4064 2056 4096
rect 2088 4064 2128 4096
rect 2160 4064 2200 4096
rect 2232 4064 2272 4096
rect 2304 4064 2344 4096
rect 2376 4064 2416 4096
rect 2448 4064 2488 4096
rect 2520 4064 2560 4096
rect 2592 4064 2632 4096
rect 2664 4064 2704 4096
rect 2736 4064 2776 4096
rect 2808 4064 2848 4096
rect 2880 4064 2920 4096
rect 2952 4064 2992 4096
rect 3024 4064 3064 4096
rect 3096 4064 3136 4096
rect 3168 4064 3208 4096
rect 3240 4064 3280 4096
rect 3312 4064 3352 4096
rect 3384 4064 3424 4096
rect 3456 4064 3496 4096
rect 3528 4064 3568 4096
rect 3600 4064 3640 4096
rect 3672 4064 3712 4096
rect 3744 4064 3784 4096
rect 3816 4064 3856 4096
rect 3888 4064 3928 4096
rect 3960 4064 4000 4096
rect 0 4024 4000 4064
rect 0 3992 40 4024
rect 72 3992 112 4024
rect 144 3992 184 4024
rect 216 3992 256 4024
rect 288 3992 328 4024
rect 360 3992 400 4024
rect 432 3992 472 4024
rect 504 3992 544 4024
rect 576 3992 616 4024
rect 648 3992 688 4024
rect 720 3992 760 4024
rect 792 3992 832 4024
rect 864 3992 904 4024
rect 936 3992 976 4024
rect 1008 3992 1048 4024
rect 1080 3992 1120 4024
rect 1152 3992 1192 4024
rect 1224 3992 1264 4024
rect 1296 3992 1336 4024
rect 1368 3992 1408 4024
rect 1440 3992 1480 4024
rect 1512 3992 1552 4024
rect 1584 3992 1624 4024
rect 1656 3992 1696 4024
rect 1728 3992 1768 4024
rect 1800 3992 1840 4024
rect 1872 3992 1912 4024
rect 1944 3992 1984 4024
rect 2016 3992 2056 4024
rect 2088 3992 2128 4024
rect 2160 3992 2200 4024
rect 2232 3992 2272 4024
rect 2304 3992 2344 4024
rect 2376 3992 2416 4024
rect 2448 3992 2488 4024
rect 2520 3992 2560 4024
rect 2592 3992 2632 4024
rect 2664 3992 2704 4024
rect 2736 3992 2776 4024
rect 2808 3992 2848 4024
rect 2880 3992 2920 4024
rect 2952 3992 2992 4024
rect 3024 3992 3064 4024
rect 3096 3992 3136 4024
rect 3168 3992 3208 4024
rect 3240 3992 3280 4024
rect 3312 3992 3352 4024
rect 3384 3992 3424 4024
rect 3456 3992 3496 4024
rect 3528 3992 3568 4024
rect 3600 3992 3640 4024
rect 3672 3992 3712 4024
rect 3744 3992 3784 4024
rect 3816 3992 3856 4024
rect 3888 3992 3928 4024
rect 3960 3992 4000 4024
rect 0 3952 4000 3992
rect 0 3920 40 3952
rect 72 3920 112 3952
rect 144 3920 184 3952
rect 216 3920 256 3952
rect 288 3920 328 3952
rect 360 3920 400 3952
rect 432 3920 472 3952
rect 504 3920 544 3952
rect 576 3920 616 3952
rect 648 3920 688 3952
rect 720 3920 760 3952
rect 792 3920 832 3952
rect 864 3920 904 3952
rect 936 3920 976 3952
rect 1008 3920 1048 3952
rect 1080 3920 1120 3952
rect 1152 3920 1192 3952
rect 1224 3920 1264 3952
rect 1296 3920 1336 3952
rect 1368 3920 1408 3952
rect 1440 3920 1480 3952
rect 1512 3920 1552 3952
rect 1584 3920 1624 3952
rect 1656 3920 1696 3952
rect 1728 3920 1768 3952
rect 1800 3920 1840 3952
rect 1872 3920 1912 3952
rect 1944 3920 1984 3952
rect 2016 3920 2056 3952
rect 2088 3920 2128 3952
rect 2160 3920 2200 3952
rect 2232 3920 2272 3952
rect 2304 3920 2344 3952
rect 2376 3920 2416 3952
rect 2448 3920 2488 3952
rect 2520 3920 2560 3952
rect 2592 3920 2632 3952
rect 2664 3920 2704 3952
rect 2736 3920 2776 3952
rect 2808 3920 2848 3952
rect 2880 3920 2920 3952
rect 2952 3920 2992 3952
rect 3024 3920 3064 3952
rect 3096 3920 3136 3952
rect 3168 3920 3208 3952
rect 3240 3920 3280 3952
rect 3312 3920 3352 3952
rect 3384 3920 3424 3952
rect 3456 3920 3496 3952
rect 3528 3920 3568 3952
rect 3600 3920 3640 3952
rect 3672 3920 3712 3952
rect 3744 3920 3784 3952
rect 3816 3920 3856 3952
rect 3888 3920 3928 3952
rect 3960 3920 4000 3952
rect 0 3880 4000 3920
rect 0 3848 40 3880
rect 72 3848 112 3880
rect 144 3848 184 3880
rect 216 3848 256 3880
rect 288 3848 328 3880
rect 360 3848 400 3880
rect 432 3848 472 3880
rect 504 3848 544 3880
rect 576 3848 616 3880
rect 648 3848 688 3880
rect 720 3848 760 3880
rect 792 3848 832 3880
rect 864 3848 904 3880
rect 936 3848 976 3880
rect 1008 3848 1048 3880
rect 1080 3848 1120 3880
rect 1152 3848 1192 3880
rect 1224 3848 1264 3880
rect 1296 3848 1336 3880
rect 1368 3848 1408 3880
rect 1440 3848 1480 3880
rect 1512 3848 1552 3880
rect 1584 3848 1624 3880
rect 1656 3848 1696 3880
rect 1728 3848 1768 3880
rect 1800 3848 1840 3880
rect 1872 3848 1912 3880
rect 1944 3848 1984 3880
rect 2016 3848 2056 3880
rect 2088 3848 2128 3880
rect 2160 3848 2200 3880
rect 2232 3848 2272 3880
rect 2304 3848 2344 3880
rect 2376 3848 2416 3880
rect 2448 3848 2488 3880
rect 2520 3848 2560 3880
rect 2592 3848 2632 3880
rect 2664 3848 2704 3880
rect 2736 3848 2776 3880
rect 2808 3848 2848 3880
rect 2880 3848 2920 3880
rect 2952 3848 2992 3880
rect 3024 3848 3064 3880
rect 3096 3848 3136 3880
rect 3168 3848 3208 3880
rect 3240 3848 3280 3880
rect 3312 3848 3352 3880
rect 3384 3848 3424 3880
rect 3456 3848 3496 3880
rect 3528 3848 3568 3880
rect 3600 3848 3640 3880
rect 3672 3848 3712 3880
rect 3744 3848 3784 3880
rect 3816 3848 3856 3880
rect 3888 3848 3928 3880
rect 3960 3848 4000 3880
rect 0 3808 4000 3848
rect 0 3776 40 3808
rect 72 3776 112 3808
rect 144 3776 184 3808
rect 216 3776 256 3808
rect 288 3776 328 3808
rect 360 3776 400 3808
rect 432 3776 472 3808
rect 504 3776 544 3808
rect 576 3776 616 3808
rect 648 3776 688 3808
rect 720 3776 760 3808
rect 792 3776 832 3808
rect 864 3776 904 3808
rect 936 3776 976 3808
rect 1008 3776 1048 3808
rect 1080 3776 1120 3808
rect 1152 3776 1192 3808
rect 1224 3776 1264 3808
rect 1296 3776 1336 3808
rect 1368 3776 1408 3808
rect 1440 3776 1480 3808
rect 1512 3776 1552 3808
rect 1584 3776 1624 3808
rect 1656 3776 1696 3808
rect 1728 3776 1768 3808
rect 1800 3776 1840 3808
rect 1872 3776 1912 3808
rect 1944 3776 1984 3808
rect 2016 3776 2056 3808
rect 2088 3776 2128 3808
rect 2160 3776 2200 3808
rect 2232 3776 2272 3808
rect 2304 3776 2344 3808
rect 2376 3776 2416 3808
rect 2448 3776 2488 3808
rect 2520 3776 2560 3808
rect 2592 3776 2632 3808
rect 2664 3776 2704 3808
rect 2736 3776 2776 3808
rect 2808 3776 2848 3808
rect 2880 3776 2920 3808
rect 2952 3776 2992 3808
rect 3024 3776 3064 3808
rect 3096 3776 3136 3808
rect 3168 3776 3208 3808
rect 3240 3776 3280 3808
rect 3312 3776 3352 3808
rect 3384 3776 3424 3808
rect 3456 3776 3496 3808
rect 3528 3776 3568 3808
rect 3600 3776 3640 3808
rect 3672 3776 3712 3808
rect 3744 3776 3784 3808
rect 3816 3776 3856 3808
rect 3888 3776 3928 3808
rect 3960 3776 4000 3808
rect 0 3736 4000 3776
rect 0 3704 40 3736
rect 72 3704 112 3736
rect 144 3704 184 3736
rect 216 3704 256 3736
rect 288 3704 328 3736
rect 360 3704 400 3736
rect 432 3704 472 3736
rect 504 3704 544 3736
rect 576 3704 616 3736
rect 648 3704 688 3736
rect 720 3704 760 3736
rect 792 3704 832 3736
rect 864 3704 904 3736
rect 936 3704 976 3736
rect 1008 3704 1048 3736
rect 1080 3704 1120 3736
rect 1152 3704 1192 3736
rect 1224 3704 1264 3736
rect 1296 3704 1336 3736
rect 1368 3704 1408 3736
rect 1440 3704 1480 3736
rect 1512 3704 1552 3736
rect 1584 3704 1624 3736
rect 1656 3704 1696 3736
rect 1728 3704 1768 3736
rect 1800 3704 1840 3736
rect 1872 3704 1912 3736
rect 1944 3704 1984 3736
rect 2016 3704 2056 3736
rect 2088 3704 2128 3736
rect 2160 3704 2200 3736
rect 2232 3704 2272 3736
rect 2304 3704 2344 3736
rect 2376 3704 2416 3736
rect 2448 3704 2488 3736
rect 2520 3704 2560 3736
rect 2592 3704 2632 3736
rect 2664 3704 2704 3736
rect 2736 3704 2776 3736
rect 2808 3704 2848 3736
rect 2880 3704 2920 3736
rect 2952 3704 2992 3736
rect 3024 3704 3064 3736
rect 3096 3704 3136 3736
rect 3168 3704 3208 3736
rect 3240 3704 3280 3736
rect 3312 3704 3352 3736
rect 3384 3704 3424 3736
rect 3456 3704 3496 3736
rect 3528 3704 3568 3736
rect 3600 3704 3640 3736
rect 3672 3704 3712 3736
rect 3744 3704 3784 3736
rect 3816 3704 3856 3736
rect 3888 3704 3928 3736
rect 3960 3704 4000 3736
rect 0 3664 4000 3704
rect 0 3632 40 3664
rect 72 3632 112 3664
rect 144 3632 184 3664
rect 216 3632 256 3664
rect 288 3632 328 3664
rect 360 3632 400 3664
rect 432 3632 472 3664
rect 504 3632 544 3664
rect 576 3632 616 3664
rect 648 3632 688 3664
rect 720 3632 760 3664
rect 792 3632 832 3664
rect 864 3632 904 3664
rect 936 3632 976 3664
rect 1008 3632 1048 3664
rect 1080 3632 1120 3664
rect 1152 3632 1192 3664
rect 1224 3632 1264 3664
rect 1296 3632 1336 3664
rect 1368 3632 1408 3664
rect 1440 3632 1480 3664
rect 1512 3632 1552 3664
rect 1584 3632 1624 3664
rect 1656 3632 1696 3664
rect 1728 3632 1768 3664
rect 1800 3632 1840 3664
rect 1872 3632 1912 3664
rect 1944 3632 1984 3664
rect 2016 3632 2056 3664
rect 2088 3632 2128 3664
rect 2160 3632 2200 3664
rect 2232 3632 2272 3664
rect 2304 3632 2344 3664
rect 2376 3632 2416 3664
rect 2448 3632 2488 3664
rect 2520 3632 2560 3664
rect 2592 3632 2632 3664
rect 2664 3632 2704 3664
rect 2736 3632 2776 3664
rect 2808 3632 2848 3664
rect 2880 3632 2920 3664
rect 2952 3632 2992 3664
rect 3024 3632 3064 3664
rect 3096 3632 3136 3664
rect 3168 3632 3208 3664
rect 3240 3632 3280 3664
rect 3312 3632 3352 3664
rect 3384 3632 3424 3664
rect 3456 3632 3496 3664
rect 3528 3632 3568 3664
rect 3600 3632 3640 3664
rect 3672 3632 3712 3664
rect 3744 3632 3784 3664
rect 3816 3632 3856 3664
rect 3888 3632 3928 3664
rect 3960 3632 4000 3664
rect 0 3592 4000 3632
rect 0 3560 40 3592
rect 72 3560 112 3592
rect 144 3560 184 3592
rect 216 3560 256 3592
rect 288 3560 328 3592
rect 360 3560 400 3592
rect 432 3560 472 3592
rect 504 3560 544 3592
rect 576 3560 616 3592
rect 648 3560 688 3592
rect 720 3560 760 3592
rect 792 3560 832 3592
rect 864 3560 904 3592
rect 936 3560 976 3592
rect 1008 3560 1048 3592
rect 1080 3560 1120 3592
rect 1152 3560 1192 3592
rect 1224 3560 1264 3592
rect 1296 3560 1336 3592
rect 1368 3560 1408 3592
rect 1440 3560 1480 3592
rect 1512 3560 1552 3592
rect 1584 3560 1624 3592
rect 1656 3560 1696 3592
rect 1728 3560 1768 3592
rect 1800 3560 1840 3592
rect 1872 3560 1912 3592
rect 1944 3560 1984 3592
rect 2016 3560 2056 3592
rect 2088 3560 2128 3592
rect 2160 3560 2200 3592
rect 2232 3560 2272 3592
rect 2304 3560 2344 3592
rect 2376 3560 2416 3592
rect 2448 3560 2488 3592
rect 2520 3560 2560 3592
rect 2592 3560 2632 3592
rect 2664 3560 2704 3592
rect 2736 3560 2776 3592
rect 2808 3560 2848 3592
rect 2880 3560 2920 3592
rect 2952 3560 2992 3592
rect 3024 3560 3064 3592
rect 3096 3560 3136 3592
rect 3168 3560 3208 3592
rect 3240 3560 3280 3592
rect 3312 3560 3352 3592
rect 3384 3560 3424 3592
rect 3456 3560 3496 3592
rect 3528 3560 3568 3592
rect 3600 3560 3640 3592
rect 3672 3560 3712 3592
rect 3744 3560 3784 3592
rect 3816 3560 3856 3592
rect 3888 3560 3928 3592
rect 3960 3560 4000 3592
rect 0 3520 4000 3560
rect 0 3488 40 3520
rect 72 3488 112 3520
rect 144 3488 184 3520
rect 216 3488 256 3520
rect 288 3488 328 3520
rect 360 3488 400 3520
rect 432 3488 472 3520
rect 504 3488 544 3520
rect 576 3488 616 3520
rect 648 3488 688 3520
rect 720 3488 760 3520
rect 792 3488 832 3520
rect 864 3488 904 3520
rect 936 3488 976 3520
rect 1008 3488 1048 3520
rect 1080 3488 1120 3520
rect 1152 3488 1192 3520
rect 1224 3488 1264 3520
rect 1296 3488 1336 3520
rect 1368 3488 1408 3520
rect 1440 3488 1480 3520
rect 1512 3488 1552 3520
rect 1584 3488 1624 3520
rect 1656 3488 1696 3520
rect 1728 3488 1768 3520
rect 1800 3488 1840 3520
rect 1872 3488 1912 3520
rect 1944 3488 1984 3520
rect 2016 3488 2056 3520
rect 2088 3488 2128 3520
rect 2160 3488 2200 3520
rect 2232 3488 2272 3520
rect 2304 3488 2344 3520
rect 2376 3488 2416 3520
rect 2448 3488 2488 3520
rect 2520 3488 2560 3520
rect 2592 3488 2632 3520
rect 2664 3488 2704 3520
rect 2736 3488 2776 3520
rect 2808 3488 2848 3520
rect 2880 3488 2920 3520
rect 2952 3488 2992 3520
rect 3024 3488 3064 3520
rect 3096 3488 3136 3520
rect 3168 3488 3208 3520
rect 3240 3488 3280 3520
rect 3312 3488 3352 3520
rect 3384 3488 3424 3520
rect 3456 3488 3496 3520
rect 3528 3488 3568 3520
rect 3600 3488 3640 3520
rect 3672 3488 3712 3520
rect 3744 3488 3784 3520
rect 3816 3488 3856 3520
rect 3888 3488 3928 3520
rect 3960 3488 4000 3520
rect 0 3448 4000 3488
rect 0 3416 40 3448
rect 72 3416 112 3448
rect 144 3416 184 3448
rect 216 3416 256 3448
rect 288 3416 328 3448
rect 360 3416 400 3448
rect 432 3416 472 3448
rect 504 3416 544 3448
rect 576 3416 616 3448
rect 648 3416 688 3448
rect 720 3416 760 3448
rect 792 3416 832 3448
rect 864 3416 904 3448
rect 936 3416 976 3448
rect 1008 3416 1048 3448
rect 1080 3416 1120 3448
rect 1152 3416 1192 3448
rect 1224 3416 1264 3448
rect 1296 3416 1336 3448
rect 1368 3416 1408 3448
rect 1440 3416 1480 3448
rect 1512 3416 1552 3448
rect 1584 3416 1624 3448
rect 1656 3416 1696 3448
rect 1728 3416 1768 3448
rect 1800 3416 1840 3448
rect 1872 3416 1912 3448
rect 1944 3416 1984 3448
rect 2016 3416 2056 3448
rect 2088 3416 2128 3448
rect 2160 3416 2200 3448
rect 2232 3416 2272 3448
rect 2304 3416 2344 3448
rect 2376 3416 2416 3448
rect 2448 3416 2488 3448
rect 2520 3416 2560 3448
rect 2592 3416 2632 3448
rect 2664 3416 2704 3448
rect 2736 3416 2776 3448
rect 2808 3416 2848 3448
rect 2880 3416 2920 3448
rect 2952 3416 2992 3448
rect 3024 3416 3064 3448
rect 3096 3416 3136 3448
rect 3168 3416 3208 3448
rect 3240 3416 3280 3448
rect 3312 3416 3352 3448
rect 3384 3416 3424 3448
rect 3456 3416 3496 3448
rect 3528 3416 3568 3448
rect 3600 3416 3640 3448
rect 3672 3416 3712 3448
rect 3744 3416 3784 3448
rect 3816 3416 3856 3448
rect 3888 3416 3928 3448
rect 3960 3416 4000 3448
rect 0 3376 4000 3416
rect 0 3344 40 3376
rect 72 3344 112 3376
rect 144 3344 184 3376
rect 216 3344 256 3376
rect 288 3344 328 3376
rect 360 3344 400 3376
rect 432 3344 472 3376
rect 504 3344 544 3376
rect 576 3344 616 3376
rect 648 3344 688 3376
rect 720 3344 760 3376
rect 792 3344 832 3376
rect 864 3344 904 3376
rect 936 3344 976 3376
rect 1008 3344 1048 3376
rect 1080 3344 1120 3376
rect 1152 3344 1192 3376
rect 1224 3344 1264 3376
rect 1296 3344 1336 3376
rect 1368 3344 1408 3376
rect 1440 3344 1480 3376
rect 1512 3344 1552 3376
rect 1584 3344 1624 3376
rect 1656 3344 1696 3376
rect 1728 3344 1768 3376
rect 1800 3344 1840 3376
rect 1872 3344 1912 3376
rect 1944 3344 1984 3376
rect 2016 3344 2056 3376
rect 2088 3344 2128 3376
rect 2160 3344 2200 3376
rect 2232 3344 2272 3376
rect 2304 3344 2344 3376
rect 2376 3344 2416 3376
rect 2448 3344 2488 3376
rect 2520 3344 2560 3376
rect 2592 3344 2632 3376
rect 2664 3344 2704 3376
rect 2736 3344 2776 3376
rect 2808 3344 2848 3376
rect 2880 3344 2920 3376
rect 2952 3344 2992 3376
rect 3024 3344 3064 3376
rect 3096 3344 3136 3376
rect 3168 3344 3208 3376
rect 3240 3344 3280 3376
rect 3312 3344 3352 3376
rect 3384 3344 3424 3376
rect 3456 3344 3496 3376
rect 3528 3344 3568 3376
rect 3600 3344 3640 3376
rect 3672 3344 3712 3376
rect 3744 3344 3784 3376
rect 3816 3344 3856 3376
rect 3888 3344 3928 3376
rect 3960 3344 4000 3376
rect 0 3304 4000 3344
rect 0 3272 40 3304
rect 72 3272 112 3304
rect 144 3272 184 3304
rect 216 3272 256 3304
rect 288 3272 328 3304
rect 360 3272 400 3304
rect 432 3272 472 3304
rect 504 3272 544 3304
rect 576 3272 616 3304
rect 648 3272 688 3304
rect 720 3272 760 3304
rect 792 3272 832 3304
rect 864 3272 904 3304
rect 936 3272 976 3304
rect 1008 3272 1048 3304
rect 1080 3272 1120 3304
rect 1152 3272 1192 3304
rect 1224 3272 1264 3304
rect 1296 3272 1336 3304
rect 1368 3272 1408 3304
rect 1440 3272 1480 3304
rect 1512 3272 1552 3304
rect 1584 3272 1624 3304
rect 1656 3272 1696 3304
rect 1728 3272 1768 3304
rect 1800 3272 1840 3304
rect 1872 3272 1912 3304
rect 1944 3272 1984 3304
rect 2016 3272 2056 3304
rect 2088 3272 2128 3304
rect 2160 3272 2200 3304
rect 2232 3272 2272 3304
rect 2304 3272 2344 3304
rect 2376 3272 2416 3304
rect 2448 3272 2488 3304
rect 2520 3272 2560 3304
rect 2592 3272 2632 3304
rect 2664 3272 2704 3304
rect 2736 3272 2776 3304
rect 2808 3272 2848 3304
rect 2880 3272 2920 3304
rect 2952 3272 2992 3304
rect 3024 3272 3064 3304
rect 3096 3272 3136 3304
rect 3168 3272 3208 3304
rect 3240 3272 3280 3304
rect 3312 3272 3352 3304
rect 3384 3272 3424 3304
rect 3456 3272 3496 3304
rect 3528 3272 3568 3304
rect 3600 3272 3640 3304
rect 3672 3272 3712 3304
rect 3744 3272 3784 3304
rect 3816 3272 3856 3304
rect 3888 3272 3928 3304
rect 3960 3272 4000 3304
rect 0 3232 4000 3272
rect 0 3200 40 3232
rect 72 3200 112 3232
rect 144 3200 184 3232
rect 216 3200 256 3232
rect 288 3200 328 3232
rect 360 3200 400 3232
rect 432 3200 472 3232
rect 504 3200 544 3232
rect 576 3200 616 3232
rect 648 3200 688 3232
rect 720 3200 760 3232
rect 792 3200 832 3232
rect 864 3200 904 3232
rect 936 3200 976 3232
rect 1008 3200 1048 3232
rect 1080 3200 1120 3232
rect 1152 3200 1192 3232
rect 1224 3200 1264 3232
rect 1296 3200 1336 3232
rect 1368 3200 1408 3232
rect 1440 3200 1480 3232
rect 1512 3200 1552 3232
rect 1584 3200 1624 3232
rect 1656 3200 1696 3232
rect 1728 3200 1768 3232
rect 1800 3200 1840 3232
rect 1872 3200 1912 3232
rect 1944 3200 1984 3232
rect 2016 3200 2056 3232
rect 2088 3200 2128 3232
rect 2160 3200 2200 3232
rect 2232 3200 2272 3232
rect 2304 3200 2344 3232
rect 2376 3200 2416 3232
rect 2448 3200 2488 3232
rect 2520 3200 2560 3232
rect 2592 3200 2632 3232
rect 2664 3200 2704 3232
rect 2736 3200 2776 3232
rect 2808 3200 2848 3232
rect 2880 3200 2920 3232
rect 2952 3200 2992 3232
rect 3024 3200 3064 3232
rect 3096 3200 3136 3232
rect 3168 3200 3208 3232
rect 3240 3200 3280 3232
rect 3312 3200 3352 3232
rect 3384 3200 3424 3232
rect 3456 3200 3496 3232
rect 3528 3200 3568 3232
rect 3600 3200 3640 3232
rect 3672 3200 3712 3232
rect 3744 3200 3784 3232
rect 3816 3200 3856 3232
rect 3888 3200 3928 3232
rect 3960 3200 4000 3232
rect 0 3160 4000 3200
rect 0 3128 40 3160
rect 72 3128 112 3160
rect 144 3128 184 3160
rect 216 3128 256 3160
rect 288 3128 328 3160
rect 360 3128 400 3160
rect 432 3128 472 3160
rect 504 3128 544 3160
rect 576 3128 616 3160
rect 648 3128 688 3160
rect 720 3128 760 3160
rect 792 3128 832 3160
rect 864 3128 904 3160
rect 936 3128 976 3160
rect 1008 3128 1048 3160
rect 1080 3128 1120 3160
rect 1152 3128 1192 3160
rect 1224 3128 1264 3160
rect 1296 3128 1336 3160
rect 1368 3128 1408 3160
rect 1440 3128 1480 3160
rect 1512 3128 1552 3160
rect 1584 3128 1624 3160
rect 1656 3128 1696 3160
rect 1728 3128 1768 3160
rect 1800 3128 1840 3160
rect 1872 3128 1912 3160
rect 1944 3128 1984 3160
rect 2016 3128 2056 3160
rect 2088 3128 2128 3160
rect 2160 3128 2200 3160
rect 2232 3128 2272 3160
rect 2304 3128 2344 3160
rect 2376 3128 2416 3160
rect 2448 3128 2488 3160
rect 2520 3128 2560 3160
rect 2592 3128 2632 3160
rect 2664 3128 2704 3160
rect 2736 3128 2776 3160
rect 2808 3128 2848 3160
rect 2880 3128 2920 3160
rect 2952 3128 2992 3160
rect 3024 3128 3064 3160
rect 3096 3128 3136 3160
rect 3168 3128 3208 3160
rect 3240 3128 3280 3160
rect 3312 3128 3352 3160
rect 3384 3128 3424 3160
rect 3456 3128 3496 3160
rect 3528 3128 3568 3160
rect 3600 3128 3640 3160
rect 3672 3128 3712 3160
rect 3744 3128 3784 3160
rect 3816 3128 3856 3160
rect 3888 3128 3928 3160
rect 3960 3128 4000 3160
rect 0 3088 4000 3128
rect 0 3056 40 3088
rect 72 3056 112 3088
rect 144 3056 184 3088
rect 216 3056 256 3088
rect 288 3056 328 3088
rect 360 3056 400 3088
rect 432 3056 472 3088
rect 504 3056 544 3088
rect 576 3056 616 3088
rect 648 3056 688 3088
rect 720 3056 760 3088
rect 792 3056 832 3088
rect 864 3056 904 3088
rect 936 3056 976 3088
rect 1008 3056 1048 3088
rect 1080 3056 1120 3088
rect 1152 3056 1192 3088
rect 1224 3056 1264 3088
rect 1296 3056 1336 3088
rect 1368 3056 1408 3088
rect 1440 3056 1480 3088
rect 1512 3056 1552 3088
rect 1584 3056 1624 3088
rect 1656 3056 1696 3088
rect 1728 3056 1768 3088
rect 1800 3056 1840 3088
rect 1872 3056 1912 3088
rect 1944 3056 1984 3088
rect 2016 3056 2056 3088
rect 2088 3056 2128 3088
rect 2160 3056 2200 3088
rect 2232 3056 2272 3088
rect 2304 3056 2344 3088
rect 2376 3056 2416 3088
rect 2448 3056 2488 3088
rect 2520 3056 2560 3088
rect 2592 3056 2632 3088
rect 2664 3056 2704 3088
rect 2736 3056 2776 3088
rect 2808 3056 2848 3088
rect 2880 3056 2920 3088
rect 2952 3056 2992 3088
rect 3024 3056 3064 3088
rect 3096 3056 3136 3088
rect 3168 3056 3208 3088
rect 3240 3056 3280 3088
rect 3312 3056 3352 3088
rect 3384 3056 3424 3088
rect 3456 3056 3496 3088
rect 3528 3056 3568 3088
rect 3600 3056 3640 3088
rect 3672 3056 3712 3088
rect 3744 3056 3784 3088
rect 3816 3056 3856 3088
rect 3888 3056 3928 3088
rect 3960 3056 4000 3088
rect 0 3016 4000 3056
rect 0 2984 40 3016
rect 72 2984 112 3016
rect 144 2984 184 3016
rect 216 2984 256 3016
rect 288 2984 328 3016
rect 360 2984 400 3016
rect 432 2984 472 3016
rect 504 2984 544 3016
rect 576 2984 616 3016
rect 648 2984 688 3016
rect 720 2984 760 3016
rect 792 2984 832 3016
rect 864 2984 904 3016
rect 936 2984 976 3016
rect 1008 2984 1048 3016
rect 1080 2984 1120 3016
rect 1152 2984 1192 3016
rect 1224 2984 1264 3016
rect 1296 2984 1336 3016
rect 1368 2984 1408 3016
rect 1440 2984 1480 3016
rect 1512 2984 1552 3016
rect 1584 2984 1624 3016
rect 1656 2984 1696 3016
rect 1728 2984 1768 3016
rect 1800 2984 1840 3016
rect 1872 2984 1912 3016
rect 1944 2984 1984 3016
rect 2016 2984 2056 3016
rect 2088 2984 2128 3016
rect 2160 2984 2200 3016
rect 2232 2984 2272 3016
rect 2304 2984 2344 3016
rect 2376 2984 2416 3016
rect 2448 2984 2488 3016
rect 2520 2984 2560 3016
rect 2592 2984 2632 3016
rect 2664 2984 2704 3016
rect 2736 2984 2776 3016
rect 2808 2984 2848 3016
rect 2880 2984 2920 3016
rect 2952 2984 2992 3016
rect 3024 2984 3064 3016
rect 3096 2984 3136 3016
rect 3168 2984 3208 3016
rect 3240 2984 3280 3016
rect 3312 2984 3352 3016
rect 3384 2984 3424 3016
rect 3456 2984 3496 3016
rect 3528 2984 3568 3016
rect 3600 2984 3640 3016
rect 3672 2984 3712 3016
rect 3744 2984 3784 3016
rect 3816 2984 3856 3016
rect 3888 2984 3928 3016
rect 3960 2984 4000 3016
rect 0 2944 4000 2984
rect 0 2912 40 2944
rect 72 2912 112 2944
rect 144 2912 184 2944
rect 216 2912 256 2944
rect 288 2912 328 2944
rect 360 2912 400 2944
rect 432 2912 472 2944
rect 504 2912 544 2944
rect 576 2912 616 2944
rect 648 2912 688 2944
rect 720 2912 760 2944
rect 792 2912 832 2944
rect 864 2912 904 2944
rect 936 2912 976 2944
rect 1008 2912 1048 2944
rect 1080 2912 1120 2944
rect 1152 2912 1192 2944
rect 1224 2912 1264 2944
rect 1296 2912 1336 2944
rect 1368 2912 1408 2944
rect 1440 2912 1480 2944
rect 1512 2912 1552 2944
rect 1584 2912 1624 2944
rect 1656 2912 1696 2944
rect 1728 2912 1768 2944
rect 1800 2912 1840 2944
rect 1872 2912 1912 2944
rect 1944 2912 1984 2944
rect 2016 2912 2056 2944
rect 2088 2912 2128 2944
rect 2160 2912 2200 2944
rect 2232 2912 2272 2944
rect 2304 2912 2344 2944
rect 2376 2912 2416 2944
rect 2448 2912 2488 2944
rect 2520 2912 2560 2944
rect 2592 2912 2632 2944
rect 2664 2912 2704 2944
rect 2736 2912 2776 2944
rect 2808 2912 2848 2944
rect 2880 2912 2920 2944
rect 2952 2912 2992 2944
rect 3024 2912 3064 2944
rect 3096 2912 3136 2944
rect 3168 2912 3208 2944
rect 3240 2912 3280 2944
rect 3312 2912 3352 2944
rect 3384 2912 3424 2944
rect 3456 2912 3496 2944
rect 3528 2912 3568 2944
rect 3600 2912 3640 2944
rect 3672 2912 3712 2944
rect 3744 2912 3784 2944
rect 3816 2912 3856 2944
rect 3888 2912 3928 2944
rect 3960 2912 4000 2944
rect 0 2872 4000 2912
rect 0 2840 40 2872
rect 72 2840 112 2872
rect 144 2840 184 2872
rect 216 2840 256 2872
rect 288 2840 328 2872
rect 360 2840 400 2872
rect 432 2840 472 2872
rect 504 2840 544 2872
rect 576 2840 616 2872
rect 648 2840 688 2872
rect 720 2840 760 2872
rect 792 2840 832 2872
rect 864 2840 904 2872
rect 936 2840 976 2872
rect 1008 2840 1048 2872
rect 1080 2840 1120 2872
rect 1152 2840 1192 2872
rect 1224 2840 1264 2872
rect 1296 2840 1336 2872
rect 1368 2840 1408 2872
rect 1440 2840 1480 2872
rect 1512 2840 1552 2872
rect 1584 2840 1624 2872
rect 1656 2840 1696 2872
rect 1728 2840 1768 2872
rect 1800 2840 1840 2872
rect 1872 2840 1912 2872
rect 1944 2840 1984 2872
rect 2016 2840 2056 2872
rect 2088 2840 2128 2872
rect 2160 2840 2200 2872
rect 2232 2840 2272 2872
rect 2304 2840 2344 2872
rect 2376 2840 2416 2872
rect 2448 2840 2488 2872
rect 2520 2840 2560 2872
rect 2592 2840 2632 2872
rect 2664 2840 2704 2872
rect 2736 2840 2776 2872
rect 2808 2840 2848 2872
rect 2880 2840 2920 2872
rect 2952 2840 2992 2872
rect 3024 2840 3064 2872
rect 3096 2840 3136 2872
rect 3168 2840 3208 2872
rect 3240 2840 3280 2872
rect 3312 2840 3352 2872
rect 3384 2840 3424 2872
rect 3456 2840 3496 2872
rect 3528 2840 3568 2872
rect 3600 2840 3640 2872
rect 3672 2840 3712 2872
rect 3744 2840 3784 2872
rect 3816 2840 3856 2872
rect 3888 2840 3928 2872
rect 3960 2840 4000 2872
rect 0 2800 4000 2840
rect 0 2768 40 2800
rect 72 2768 112 2800
rect 144 2768 184 2800
rect 216 2768 256 2800
rect 288 2768 328 2800
rect 360 2768 400 2800
rect 432 2768 472 2800
rect 504 2768 544 2800
rect 576 2768 616 2800
rect 648 2768 688 2800
rect 720 2768 760 2800
rect 792 2768 832 2800
rect 864 2768 904 2800
rect 936 2768 976 2800
rect 1008 2768 1048 2800
rect 1080 2768 1120 2800
rect 1152 2768 1192 2800
rect 1224 2768 1264 2800
rect 1296 2768 1336 2800
rect 1368 2768 1408 2800
rect 1440 2768 1480 2800
rect 1512 2768 1552 2800
rect 1584 2768 1624 2800
rect 1656 2768 1696 2800
rect 1728 2768 1768 2800
rect 1800 2768 1840 2800
rect 1872 2768 1912 2800
rect 1944 2768 1984 2800
rect 2016 2768 2056 2800
rect 2088 2768 2128 2800
rect 2160 2768 2200 2800
rect 2232 2768 2272 2800
rect 2304 2768 2344 2800
rect 2376 2768 2416 2800
rect 2448 2768 2488 2800
rect 2520 2768 2560 2800
rect 2592 2768 2632 2800
rect 2664 2768 2704 2800
rect 2736 2768 2776 2800
rect 2808 2768 2848 2800
rect 2880 2768 2920 2800
rect 2952 2768 2992 2800
rect 3024 2768 3064 2800
rect 3096 2768 3136 2800
rect 3168 2768 3208 2800
rect 3240 2768 3280 2800
rect 3312 2768 3352 2800
rect 3384 2768 3424 2800
rect 3456 2768 3496 2800
rect 3528 2768 3568 2800
rect 3600 2768 3640 2800
rect 3672 2768 3712 2800
rect 3744 2768 3784 2800
rect 3816 2768 3856 2800
rect 3888 2768 3928 2800
rect 3960 2768 4000 2800
rect 0 2728 4000 2768
rect 0 2696 40 2728
rect 72 2696 112 2728
rect 144 2696 184 2728
rect 216 2696 256 2728
rect 288 2696 328 2728
rect 360 2696 400 2728
rect 432 2696 472 2728
rect 504 2696 544 2728
rect 576 2696 616 2728
rect 648 2696 688 2728
rect 720 2696 760 2728
rect 792 2696 832 2728
rect 864 2696 904 2728
rect 936 2696 976 2728
rect 1008 2696 1048 2728
rect 1080 2696 1120 2728
rect 1152 2696 1192 2728
rect 1224 2696 1264 2728
rect 1296 2696 1336 2728
rect 1368 2696 1408 2728
rect 1440 2696 1480 2728
rect 1512 2696 1552 2728
rect 1584 2696 1624 2728
rect 1656 2696 1696 2728
rect 1728 2696 1768 2728
rect 1800 2696 1840 2728
rect 1872 2696 1912 2728
rect 1944 2696 1984 2728
rect 2016 2696 2056 2728
rect 2088 2696 2128 2728
rect 2160 2696 2200 2728
rect 2232 2696 2272 2728
rect 2304 2696 2344 2728
rect 2376 2696 2416 2728
rect 2448 2696 2488 2728
rect 2520 2696 2560 2728
rect 2592 2696 2632 2728
rect 2664 2696 2704 2728
rect 2736 2696 2776 2728
rect 2808 2696 2848 2728
rect 2880 2696 2920 2728
rect 2952 2696 2992 2728
rect 3024 2696 3064 2728
rect 3096 2696 3136 2728
rect 3168 2696 3208 2728
rect 3240 2696 3280 2728
rect 3312 2696 3352 2728
rect 3384 2696 3424 2728
rect 3456 2696 3496 2728
rect 3528 2696 3568 2728
rect 3600 2696 3640 2728
rect 3672 2696 3712 2728
rect 3744 2696 3784 2728
rect 3816 2696 3856 2728
rect 3888 2696 3928 2728
rect 3960 2696 4000 2728
rect 0 2656 4000 2696
rect 0 2624 40 2656
rect 72 2624 112 2656
rect 144 2624 184 2656
rect 216 2624 256 2656
rect 288 2624 328 2656
rect 360 2624 400 2656
rect 432 2624 472 2656
rect 504 2624 544 2656
rect 576 2624 616 2656
rect 648 2624 688 2656
rect 720 2624 760 2656
rect 792 2624 832 2656
rect 864 2624 904 2656
rect 936 2624 976 2656
rect 1008 2624 1048 2656
rect 1080 2624 1120 2656
rect 1152 2624 1192 2656
rect 1224 2624 1264 2656
rect 1296 2624 1336 2656
rect 1368 2624 1408 2656
rect 1440 2624 1480 2656
rect 1512 2624 1552 2656
rect 1584 2624 1624 2656
rect 1656 2624 1696 2656
rect 1728 2624 1768 2656
rect 1800 2624 1840 2656
rect 1872 2624 1912 2656
rect 1944 2624 1984 2656
rect 2016 2624 2056 2656
rect 2088 2624 2128 2656
rect 2160 2624 2200 2656
rect 2232 2624 2272 2656
rect 2304 2624 2344 2656
rect 2376 2624 2416 2656
rect 2448 2624 2488 2656
rect 2520 2624 2560 2656
rect 2592 2624 2632 2656
rect 2664 2624 2704 2656
rect 2736 2624 2776 2656
rect 2808 2624 2848 2656
rect 2880 2624 2920 2656
rect 2952 2624 2992 2656
rect 3024 2624 3064 2656
rect 3096 2624 3136 2656
rect 3168 2624 3208 2656
rect 3240 2624 3280 2656
rect 3312 2624 3352 2656
rect 3384 2624 3424 2656
rect 3456 2624 3496 2656
rect 3528 2624 3568 2656
rect 3600 2624 3640 2656
rect 3672 2624 3712 2656
rect 3744 2624 3784 2656
rect 3816 2624 3856 2656
rect 3888 2624 3928 2656
rect 3960 2624 4000 2656
rect 0 2584 4000 2624
rect 0 2552 40 2584
rect 72 2552 112 2584
rect 144 2552 184 2584
rect 216 2552 256 2584
rect 288 2552 328 2584
rect 360 2552 400 2584
rect 432 2552 472 2584
rect 504 2552 544 2584
rect 576 2552 616 2584
rect 648 2552 688 2584
rect 720 2552 760 2584
rect 792 2552 832 2584
rect 864 2552 904 2584
rect 936 2552 976 2584
rect 1008 2552 1048 2584
rect 1080 2552 1120 2584
rect 1152 2552 1192 2584
rect 1224 2552 1264 2584
rect 1296 2552 1336 2584
rect 1368 2552 1408 2584
rect 1440 2552 1480 2584
rect 1512 2552 1552 2584
rect 1584 2552 1624 2584
rect 1656 2552 1696 2584
rect 1728 2552 1768 2584
rect 1800 2552 1840 2584
rect 1872 2552 1912 2584
rect 1944 2552 1984 2584
rect 2016 2552 2056 2584
rect 2088 2552 2128 2584
rect 2160 2552 2200 2584
rect 2232 2552 2272 2584
rect 2304 2552 2344 2584
rect 2376 2552 2416 2584
rect 2448 2552 2488 2584
rect 2520 2552 2560 2584
rect 2592 2552 2632 2584
rect 2664 2552 2704 2584
rect 2736 2552 2776 2584
rect 2808 2552 2848 2584
rect 2880 2552 2920 2584
rect 2952 2552 2992 2584
rect 3024 2552 3064 2584
rect 3096 2552 3136 2584
rect 3168 2552 3208 2584
rect 3240 2552 3280 2584
rect 3312 2552 3352 2584
rect 3384 2552 3424 2584
rect 3456 2552 3496 2584
rect 3528 2552 3568 2584
rect 3600 2552 3640 2584
rect 3672 2552 3712 2584
rect 3744 2552 3784 2584
rect 3816 2552 3856 2584
rect 3888 2552 3928 2584
rect 3960 2552 4000 2584
rect 0 2512 4000 2552
rect 0 2480 40 2512
rect 72 2480 112 2512
rect 144 2480 184 2512
rect 216 2480 256 2512
rect 288 2480 328 2512
rect 360 2480 400 2512
rect 432 2480 472 2512
rect 504 2480 544 2512
rect 576 2480 616 2512
rect 648 2480 688 2512
rect 720 2480 760 2512
rect 792 2480 832 2512
rect 864 2480 904 2512
rect 936 2480 976 2512
rect 1008 2480 1048 2512
rect 1080 2480 1120 2512
rect 1152 2480 1192 2512
rect 1224 2480 1264 2512
rect 1296 2480 1336 2512
rect 1368 2480 1408 2512
rect 1440 2480 1480 2512
rect 1512 2480 1552 2512
rect 1584 2480 1624 2512
rect 1656 2480 1696 2512
rect 1728 2480 1768 2512
rect 1800 2480 1840 2512
rect 1872 2480 1912 2512
rect 1944 2480 1984 2512
rect 2016 2480 2056 2512
rect 2088 2480 2128 2512
rect 2160 2480 2200 2512
rect 2232 2480 2272 2512
rect 2304 2480 2344 2512
rect 2376 2480 2416 2512
rect 2448 2480 2488 2512
rect 2520 2480 2560 2512
rect 2592 2480 2632 2512
rect 2664 2480 2704 2512
rect 2736 2480 2776 2512
rect 2808 2480 2848 2512
rect 2880 2480 2920 2512
rect 2952 2480 2992 2512
rect 3024 2480 3064 2512
rect 3096 2480 3136 2512
rect 3168 2480 3208 2512
rect 3240 2480 3280 2512
rect 3312 2480 3352 2512
rect 3384 2480 3424 2512
rect 3456 2480 3496 2512
rect 3528 2480 3568 2512
rect 3600 2480 3640 2512
rect 3672 2480 3712 2512
rect 3744 2480 3784 2512
rect 3816 2480 3856 2512
rect 3888 2480 3928 2512
rect 3960 2480 4000 2512
rect 0 2440 4000 2480
rect 0 2408 40 2440
rect 72 2408 112 2440
rect 144 2408 184 2440
rect 216 2408 256 2440
rect 288 2408 328 2440
rect 360 2408 400 2440
rect 432 2408 472 2440
rect 504 2408 544 2440
rect 576 2408 616 2440
rect 648 2408 688 2440
rect 720 2408 760 2440
rect 792 2408 832 2440
rect 864 2408 904 2440
rect 936 2408 976 2440
rect 1008 2408 1048 2440
rect 1080 2408 1120 2440
rect 1152 2408 1192 2440
rect 1224 2408 1264 2440
rect 1296 2408 1336 2440
rect 1368 2408 1408 2440
rect 1440 2408 1480 2440
rect 1512 2408 1552 2440
rect 1584 2408 1624 2440
rect 1656 2408 1696 2440
rect 1728 2408 1768 2440
rect 1800 2408 1840 2440
rect 1872 2408 1912 2440
rect 1944 2408 1984 2440
rect 2016 2408 2056 2440
rect 2088 2408 2128 2440
rect 2160 2408 2200 2440
rect 2232 2408 2272 2440
rect 2304 2408 2344 2440
rect 2376 2408 2416 2440
rect 2448 2408 2488 2440
rect 2520 2408 2560 2440
rect 2592 2408 2632 2440
rect 2664 2408 2704 2440
rect 2736 2408 2776 2440
rect 2808 2408 2848 2440
rect 2880 2408 2920 2440
rect 2952 2408 2992 2440
rect 3024 2408 3064 2440
rect 3096 2408 3136 2440
rect 3168 2408 3208 2440
rect 3240 2408 3280 2440
rect 3312 2408 3352 2440
rect 3384 2408 3424 2440
rect 3456 2408 3496 2440
rect 3528 2408 3568 2440
rect 3600 2408 3640 2440
rect 3672 2408 3712 2440
rect 3744 2408 3784 2440
rect 3816 2408 3856 2440
rect 3888 2408 3928 2440
rect 3960 2408 4000 2440
rect 0 2368 4000 2408
rect 0 2336 40 2368
rect 72 2336 112 2368
rect 144 2336 184 2368
rect 216 2336 256 2368
rect 288 2336 328 2368
rect 360 2336 400 2368
rect 432 2336 472 2368
rect 504 2336 544 2368
rect 576 2336 616 2368
rect 648 2336 688 2368
rect 720 2336 760 2368
rect 792 2336 832 2368
rect 864 2336 904 2368
rect 936 2336 976 2368
rect 1008 2336 1048 2368
rect 1080 2336 1120 2368
rect 1152 2336 1192 2368
rect 1224 2336 1264 2368
rect 1296 2336 1336 2368
rect 1368 2336 1408 2368
rect 1440 2336 1480 2368
rect 1512 2336 1552 2368
rect 1584 2336 1624 2368
rect 1656 2336 1696 2368
rect 1728 2336 1768 2368
rect 1800 2336 1840 2368
rect 1872 2336 1912 2368
rect 1944 2336 1984 2368
rect 2016 2336 2056 2368
rect 2088 2336 2128 2368
rect 2160 2336 2200 2368
rect 2232 2336 2272 2368
rect 2304 2336 2344 2368
rect 2376 2336 2416 2368
rect 2448 2336 2488 2368
rect 2520 2336 2560 2368
rect 2592 2336 2632 2368
rect 2664 2336 2704 2368
rect 2736 2336 2776 2368
rect 2808 2336 2848 2368
rect 2880 2336 2920 2368
rect 2952 2336 2992 2368
rect 3024 2336 3064 2368
rect 3096 2336 3136 2368
rect 3168 2336 3208 2368
rect 3240 2336 3280 2368
rect 3312 2336 3352 2368
rect 3384 2336 3424 2368
rect 3456 2336 3496 2368
rect 3528 2336 3568 2368
rect 3600 2336 3640 2368
rect 3672 2336 3712 2368
rect 3744 2336 3784 2368
rect 3816 2336 3856 2368
rect 3888 2336 3928 2368
rect 3960 2336 4000 2368
rect 0 2296 4000 2336
rect 0 2264 40 2296
rect 72 2264 112 2296
rect 144 2264 184 2296
rect 216 2264 256 2296
rect 288 2264 328 2296
rect 360 2264 400 2296
rect 432 2264 472 2296
rect 504 2264 544 2296
rect 576 2264 616 2296
rect 648 2264 688 2296
rect 720 2264 760 2296
rect 792 2264 832 2296
rect 864 2264 904 2296
rect 936 2264 976 2296
rect 1008 2264 1048 2296
rect 1080 2264 1120 2296
rect 1152 2264 1192 2296
rect 1224 2264 1264 2296
rect 1296 2264 1336 2296
rect 1368 2264 1408 2296
rect 1440 2264 1480 2296
rect 1512 2264 1552 2296
rect 1584 2264 1624 2296
rect 1656 2264 1696 2296
rect 1728 2264 1768 2296
rect 1800 2264 1840 2296
rect 1872 2264 1912 2296
rect 1944 2264 1984 2296
rect 2016 2264 2056 2296
rect 2088 2264 2128 2296
rect 2160 2264 2200 2296
rect 2232 2264 2272 2296
rect 2304 2264 2344 2296
rect 2376 2264 2416 2296
rect 2448 2264 2488 2296
rect 2520 2264 2560 2296
rect 2592 2264 2632 2296
rect 2664 2264 2704 2296
rect 2736 2264 2776 2296
rect 2808 2264 2848 2296
rect 2880 2264 2920 2296
rect 2952 2264 2992 2296
rect 3024 2264 3064 2296
rect 3096 2264 3136 2296
rect 3168 2264 3208 2296
rect 3240 2264 3280 2296
rect 3312 2264 3352 2296
rect 3384 2264 3424 2296
rect 3456 2264 3496 2296
rect 3528 2264 3568 2296
rect 3600 2264 3640 2296
rect 3672 2264 3712 2296
rect 3744 2264 3784 2296
rect 3816 2264 3856 2296
rect 3888 2264 3928 2296
rect 3960 2264 4000 2296
rect 0 2224 4000 2264
rect 0 2192 40 2224
rect 72 2192 112 2224
rect 144 2192 184 2224
rect 216 2192 256 2224
rect 288 2192 328 2224
rect 360 2192 400 2224
rect 432 2192 472 2224
rect 504 2192 544 2224
rect 576 2192 616 2224
rect 648 2192 688 2224
rect 720 2192 760 2224
rect 792 2192 832 2224
rect 864 2192 904 2224
rect 936 2192 976 2224
rect 1008 2192 1048 2224
rect 1080 2192 1120 2224
rect 1152 2192 1192 2224
rect 1224 2192 1264 2224
rect 1296 2192 1336 2224
rect 1368 2192 1408 2224
rect 1440 2192 1480 2224
rect 1512 2192 1552 2224
rect 1584 2192 1624 2224
rect 1656 2192 1696 2224
rect 1728 2192 1768 2224
rect 1800 2192 1840 2224
rect 1872 2192 1912 2224
rect 1944 2192 1984 2224
rect 2016 2192 2056 2224
rect 2088 2192 2128 2224
rect 2160 2192 2200 2224
rect 2232 2192 2272 2224
rect 2304 2192 2344 2224
rect 2376 2192 2416 2224
rect 2448 2192 2488 2224
rect 2520 2192 2560 2224
rect 2592 2192 2632 2224
rect 2664 2192 2704 2224
rect 2736 2192 2776 2224
rect 2808 2192 2848 2224
rect 2880 2192 2920 2224
rect 2952 2192 2992 2224
rect 3024 2192 3064 2224
rect 3096 2192 3136 2224
rect 3168 2192 3208 2224
rect 3240 2192 3280 2224
rect 3312 2192 3352 2224
rect 3384 2192 3424 2224
rect 3456 2192 3496 2224
rect 3528 2192 3568 2224
rect 3600 2192 3640 2224
rect 3672 2192 3712 2224
rect 3744 2192 3784 2224
rect 3816 2192 3856 2224
rect 3888 2192 3928 2224
rect 3960 2192 4000 2224
rect 0 2152 4000 2192
rect 0 2120 40 2152
rect 72 2120 112 2152
rect 144 2120 184 2152
rect 216 2120 256 2152
rect 288 2120 328 2152
rect 360 2120 400 2152
rect 432 2120 472 2152
rect 504 2120 544 2152
rect 576 2120 616 2152
rect 648 2120 688 2152
rect 720 2120 760 2152
rect 792 2120 832 2152
rect 864 2120 904 2152
rect 936 2120 976 2152
rect 1008 2120 1048 2152
rect 1080 2120 1120 2152
rect 1152 2120 1192 2152
rect 1224 2120 1264 2152
rect 1296 2120 1336 2152
rect 1368 2120 1408 2152
rect 1440 2120 1480 2152
rect 1512 2120 1552 2152
rect 1584 2120 1624 2152
rect 1656 2120 1696 2152
rect 1728 2120 1768 2152
rect 1800 2120 1840 2152
rect 1872 2120 1912 2152
rect 1944 2120 1984 2152
rect 2016 2120 2056 2152
rect 2088 2120 2128 2152
rect 2160 2120 2200 2152
rect 2232 2120 2272 2152
rect 2304 2120 2344 2152
rect 2376 2120 2416 2152
rect 2448 2120 2488 2152
rect 2520 2120 2560 2152
rect 2592 2120 2632 2152
rect 2664 2120 2704 2152
rect 2736 2120 2776 2152
rect 2808 2120 2848 2152
rect 2880 2120 2920 2152
rect 2952 2120 2992 2152
rect 3024 2120 3064 2152
rect 3096 2120 3136 2152
rect 3168 2120 3208 2152
rect 3240 2120 3280 2152
rect 3312 2120 3352 2152
rect 3384 2120 3424 2152
rect 3456 2120 3496 2152
rect 3528 2120 3568 2152
rect 3600 2120 3640 2152
rect 3672 2120 3712 2152
rect 3744 2120 3784 2152
rect 3816 2120 3856 2152
rect 3888 2120 3928 2152
rect 3960 2120 4000 2152
rect 0 2080 4000 2120
rect 0 2048 40 2080
rect 72 2048 112 2080
rect 144 2048 184 2080
rect 216 2048 256 2080
rect 288 2048 328 2080
rect 360 2048 400 2080
rect 432 2048 472 2080
rect 504 2048 544 2080
rect 576 2048 616 2080
rect 648 2048 688 2080
rect 720 2048 760 2080
rect 792 2048 832 2080
rect 864 2048 904 2080
rect 936 2048 976 2080
rect 1008 2048 1048 2080
rect 1080 2048 1120 2080
rect 1152 2048 1192 2080
rect 1224 2048 1264 2080
rect 1296 2048 1336 2080
rect 1368 2048 1408 2080
rect 1440 2048 1480 2080
rect 1512 2048 1552 2080
rect 1584 2048 1624 2080
rect 1656 2048 1696 2080
rect 1728 2048 1768 2080
rect 1800 2048 1840 2080
rect 1872 2048 1912 2080
rect 1944 2048 1984 2080
rect 2016 2048 2056 2080
rect 2088 2048 2128 2080
rect 2160 2048 2200 2080
rect 2232 2048 2272 2080
rect 2304 2048 2344 2080
rect 2376 2048 2416 2080
rect 2448 2048 2488 2080
rect 2520 2048 2560 2080
rect 2592 2048 2632 2080
rect 2664 2048 2704 2080
rect 2736 2048 2776 2080
rect 2808 2048 2848 2080
rect 2880 2048 2920 2080
rect 2952 2048 2992 2080
rect 3024 2048 3064 2080
rect 3096 2048 3136 2080
rect 3168 2048 3208 2080
rect 3240 2048 3280 2080
rect 3312 2048 3352 2080
rect 3384 2048 3424 2080
rect 3456 2048 3496 2080
rect 3528 2048 3568 2080
rect 3600 2048 3640 2080
rect 3672 2048 3712 2080
rect 3744 2048 3784 2080
rect 3816 2048 3856 2080
rect 3888 2048 3928 2080
rect 3960 2048 4000 2080
rect 0 2008 4000 2048
rect 0 1976 40 2008
rect 72 1976 112 2008
rect 144 1976 184 2008
rect 216 1976 256 2008
rect 288 1976 328 2008
rect 360 1976 400 2008
rect 432 1976 472 2008
rect 504 1976 544 2008
rect 576 1976 616 2008
rect 648 1976 688 2008
rect 720 1976 760 2008
rect 792 1976 832 2008
rect 864 1976 904 2008
rect 936 1976 976 2008
rect 1008 1976 1048 2008
rect 1080 1976 1120 2008
rect 1152 1976 1192 2008
rect 1224 1976 1264 2008
rect 1296 1976 1336 2008
rect 1368 1976 1408 2008
rect 1440 1976 1480 2008
rect 1512 1976 1552 2008
rect 1584 1976 1624 2008
rect 1656 1976 1696 2008
rect 1728 1976 1768 2008
rect 1800 1976 1840 2008
rect 1872 1976 1912 2008
rect 1944 1976 1984 2008
rect 2016 1976 2056 2008
rect 2088 1976 2128 2008
rect 2160 1976 2200 2008
rect 2232 1976 2272 2008
rect 2304 1976 2344 2008
rect 2376 1976 2416 2008
rect 2448 1976 2488 2008
rect 2520 1976 2560 2008
rect 2592 1976 2632 2008
rect 2664 1976 2704 2008
rect 2736 1976 2776 2008
rect 2808 1976 2848 2008
rect 2880 1976 2920 2008
rect 2952 1976 2992 2008
rect 3024 1976 3064 2008
rect 3096 1976 3136 2008
rect 3168 1976 3208 2008
rect 3240 1976 3280 2008
rect 3312 1976 3352 2008
rect 3384 1976 3424 2008
rect 3456 1976 3496 2008
rect 3528 1976 3568 2008
rect 3600 1976 3640 2008
rect 3672 1976 3712 2008
rect 3744 1976 3784 2008
rect 3816 1976 3856 2008
rect 3888 1976 3928 2008
rect 3960 1976 4000 2008
rect 0 1936 4000 1976
rect 0 1904 40 1936
rect 72 1904 112 1936
rect 144 1904 184 1936
rect 216 1904 256 1936
rect 288 1904 328 1936
rect 360 1904 400 1936
rect 432 1904 472 1936
rect 504 1904 544 1936
rect 576 1904 616 1936
rect 648 1904 688 1936
rect 720 1904 760 1936
rect 792 1904 832 1936
rect 864 1904 904 1936
rect 936 1904 976 1936
rect 1008 1904 1048 1936
rect 1080 1904 1120 1936
rect 1152 1904 1192 1936
rect 1224 1904 1264 1936
rect 1296 1904 1336 1936
rect 1368 1904 1408 1936
rect 1440 1904 1480 1936
rect 1512 1904 1552 1936
rect 1584 1904 1624 1936
rect 1656 1904 1696 1936
rect 1728 1904 1768 1936
rect 1800 1904 1840 1936
rect 1872 1904 1912 1936
rect 1944 1904 1984 1936
rect 2016 1904 2056 1936
rect 2088 1904 2128 1936
rect 2160 1904 2200 1936
rect 2232 1904 2272 1936
rect 2304 1904 2344 1936
rect 2376 1904 2416 1936
rect 2448 1904 2488 1936
rect 2520 1904 2560 1936
rect 2592 1904 2632 1936
rect 2664 1904 2704 1936
rect 2736 1904 2776 1936
rect 2808 1904 2848 1936
rect 2880 1904 2920 1936
rect 2952 1904 2992 1936
rect 3024 1904 3064 1936
rect 3096 1904 3136 1936
rect 3168 1904 3208 1936
rect 3240 1904 3280 1936
rect 3312 1904 3352 1936
rect 3384 1904 3424 1936
rect 3456 1904 3496 1936
rect 3528 1904 3568 1936
rect 3600 1904 3640 1936
rect 3672 1904 3712 1936
rect 3744 1904 3784 1936
rect 3816 1904 3856 1936
rect 3888 1904 3928 1936
rect 3960 1904 4000 1936
rect 0 1864 4000 1904
rect 0 1832 40 1864
rect 72 1832 112 1864
rect 144 1832 184 1864
rect 216 1832 256 1864
rect 288 1832 328 1864
rect 360 1832 400 1864
rect 432 1832 472 1864
rect 504 1832 544 1864
rect 576 1832 616 1864
rect 648 1832 688 1864
rect 720 1832 760 1864
rect 792 1832 832 1864
rect 864 1832 904 1864
rect 936 1832 976 1864
rect 1008 1832 1048 1864
rect 1080 1832 1120 1864
rect 1152 1832 1192 1864
rect 1224 1832 1264 1864
rect 1296 1832 1336 1864
rect 1368 1832 1408 1864
rect 1440 1832 1480 1864
rect 1512 1832 1552 1864
rect 1584 1832 1624 1864
rect 1656 1832 1696 1864
rect 1728 1832 1768 1864
rect 1800 1832 1840 1864
rect 1872 1832 1912 1864
rect 1944 1832 1984 1864
rect 2016 1832 2056 1864
rect 2088 1832 2128 1864
rect 2160 1832 2200 1864
rect 2232 1832 2272 1864
rect 2304 1832 2344 1864
rect 2376 1832 2416 1864
rect 2448 1832 2488 1864
rect 2520 1832 2560 1864
rect 2592 1832 2632 1864
rect 2664 1832 2704 1864
rect 2736 1832 2776 1864
rect 2808 1832 2848 1864
rect 2880 1832 2920 1864
rect 2952 1832 2992 1864
rect 3024 1832 3064 1864
rect 3096 1832 3136 1864
rect 3168 1832 3208 1864
rect 3240 1832 3280 1864
rect 3312 1832 3352 1864
rect 3384 1832 3424 1864
rect 3456 1832 3496 1864
rect 3528 1832 3568 1864
rect 3600 1832 3640 1864
rect 3672 1832 3712 1864
rect 3744 1832 3784 1864
rect 3816 1832 3856 1864
rect 3888 1832 3928 1864
rect 3960 1832 4000 1864
rect 0 1792 4000 1832
rect 0 1760 40 1792
rect 72 1760 112 1792
rect 144 1760 184 1792
rect 216 1760 256 1792
rect 288 1760 328 1792
rect 360 1760 400 1792
rect 432 1760 472 1792
rect 504 1760 544 1792
rect 576 1760 616 1792
rect 648 1760 688 1792
rect 720 1760 760 1792
rect 792 1760 832 1792
rect 864 1760 904 1792
rect 936 1760 976 1792
rect 1008 1760 1048 1792
rect 1080 1760 1120 1792
rect 1152 1760 1192 1792
rect 1224 1760 1264 1792
rect 1296 1760 1336 1792
rect 1368 1760 1408 1792
rect 1440 1760 1480 1792
rect 1512 1760 1552 1792
rect 1584 1760 1624 1792
rect 1656 1760 1696 1792
rect 1728 1760 1768 1792
rect 1800 1760 1840 1792
rect 1872 1760 1912 1792
rect 1944 1760 1984 1792
rect 2016 1760 2056 1792
rect 2088 1760 2128 1792
rect 2160 1760 2200 1792
rect 2232 1760 2272 1792
rect 2304 1760 2344 1792
rect 2376 1760 2416 1792
rect 2448 1760 2488 1792
rect 2520 1760 2560 1792
rect 2592 1760 2632 1792
rect 2664 1760 2704 1792
rect 2736 1760 2776 1792
rect 2808 1760 2848 1792
rect 2880 1760 2920 1792
rect 2952 1760 2992 1792
rect 3024 1760 3064 1792
rect 3096 1760 3136 1792
rect 3168 1760 3208 1792
rect 3240 1760 3280 1792
rect 3312 1760 3352 1792
rect 3384 1760 3424 1792
rect 3456 1760 3496 1792
rect 3528 1760 3568 1792
rect 3600 1760 3640 1792
rect 3672 1760 3712 1792
rect 3744 1760 3784 1792
rect 3816 1760 3856 1792
rect 3888 1760 3928 1792
rect 3960 1760 4000 1792
rect 0 1720 4000 1760
rect 0 1688 40 1720
rect 72 1688 112 1720
rect 144 1688 184 1720
rect 216 1688 256 1720
rect 288 1688 328 1720
rect 360 1688 400 1720
rect 432 1688 472 1720
rect 504 1688 544 1720
rect 576 1688 616 1720
rect 648 1688 688 1720
rect 720 1688 760 1720
rect 792 1688 832 1720
rect 864 1688 904 1720
rect 936 1688 976 1720
rect 1008 1688 1048 1720
rect 1080 1688 1120 1720
rect 1152 1688 1192 1720
rect 1224 1688 1264 1720
rect 1296 1688 1336 1720
rect 1368 1688 1408 1720
rect 1440 1688 1480 1720
rect 1512 1688 1552 1720
rect 1584 1688 1624 1720
rect 1656 1688 1696 1720
rect 1728 1688 1768 1720
rect 1800 1688 1840 1720
rect 1872 1688 1912 1720
rect 1944 1688 1984 1720
rect 2016 1688 2056 1720
rect 2088 1688 2128 1720
rect 2160 1688 2200 1720
rect 2232 1688 2272 1720
rect 2304 1688 2344 1720
rect 2376 1688 2416 1720
rect 2448 1688 2488 1720
rect 2520 1688 2560 1720
rect 2592 1688 2632 1720
rect 2664 1688 2704 1720
rect 2736 1688 2776 1720
rect 2808 1688 2848 1720
rect 2880 1688 2920 1720
rect 2952 1688 2992 1720
rect 3024 1688 3064 1720
rect 3096 1688 3136 1720
rect 3168 1688 3208 1720
rect 3240 1688 3280 1720
rect 3312 1688 3352 1720
rect 3384 1688 3424 1720
rect 3456 1688 3496 1720
rect 3528 1688 3568 1720
rect 3600 1688 3640 1720
rect 3672 1688 3712 1720
rect 3744 1688 3784 1720
rect 3816 1688 3856 1720
rect 3888 1688 3928 1720
rect 3960 1688 4000 1720
rect 0 1648 4000 1688
rect 0 1616 40 1648
rect 72 1616 112 1648
rect 144 1616 184 1648
rect 216 1616 256 1648
rect 288 1616 328 1648
rect 360 1616 400 1648
rect 432 1616 472 1648
rect 504 1616 544 1648
rect 576 1616 616 1648
rect 648 1616 688 1648
rect 720 1616 760 1648
rect 792 1616 832 1648
rect 864 1616 904 1648
rect 936 1616 976 1648
rect 1008 1616 1048 1648
rect 1080 1616 1120 1648
rect 1152 1616 1192 1648
rect 1224 1616 1264 1648
rect 1296 1616 1336 1648
rect 1368 1616 1408 1648
rect 1440 1616 1480 1648
rect 1512 1616 1552 1648
rect 1584 1616 1624 1648
rect 1656 1616 1696 1648
rect 1728 1616 1768 1648
rect 1800 1616 1840 1648
rect 1872 1616 1912 1648
rect 1944 1616 1984 1648
rect 2016 1616 2056 1648
rect 2088 1616 2128 1648
rect 2160 1616 2200 1648
rect 2232 1616 2272 1648
rect 2304 1616 2344 1648
rect 2376 1616 2416 1648
rect 2448 1616 2488 1648
rect 2520 1616 2560 1648
rect 2592 1616 2632 1648
rect 2664 1616 2704 1648
rect 2736 1616 2776 1648
rect 2808 1616 2848 1648
rect 2880 1616 2920 1648
rect 2952 1616 2992 1648
rect 3024 1616 3064 1648
rect 3096 1616 3136 1648
rect 3168 1616 3208 1648
rect 3240 1616 3280 1648
rect 3312 1616 3352 1648
rect 3384 1616 3424 1648
rect 3456 1616 3496 1648
rect 3528 1616 3568 1648
rect 3600 1616 3640 1648
rect 3672 1616 3712 1648
rect 3744 1616 3784 1648
rect 3816 1616 3856 1648
rect 3888 1616 3928 1648
rect 3960 1616 4000 1648
rect 0 1576 4000 1616
rect 0 1544 40 1576
rect 72 1544 112 1576
rect 144 1544 184 1576
rect 216 1544 256 1576
rect 288 1544 328 1576
rect 360 1544 400 1576
rect 432 1544 472 1576
rect 504 1544 544 1576
rect 576 1544 616 1576
rect 648 1544 688 1576
rect 720 1544 760 1576
rect 792 1544 832 1576
rect 864 1544 904 1576
rect 936 1544 976 1576
rect 1008 1544 1048 1576
rect 1080 1544 1120 1576
rect 1152 1544 1192 1576
rect 1224 1544 1264 1576
rect 1296 1544 1336 1576
rect 1368 1544 1408 1576
rect 1440 1544 1480 1576
rect 1512 1544 1552 1576
rect 1584 1544 1624 1576
rect 1656 1544 1696 1576
rect 1728 1544 1768 1576
rect 1800 1544 1840 1576
rect 1872 1544 1912 1576
rect 1944 1544 1984 1576
rect 2016 1544 2056 1576
rect 2088 1544 2128 1576
rect 2160 1544 2200 1576
rect 2232 1544 2272 1576
rect 2304 1544 2344 1576
rect 2376 1544 2416 1576
rect 2448 1544 2488 1576
rect 2520 1544 2560 1576
rect 2592 1544 2632 1576
rect 2664 1544 2704 1576
rect 2736 1544 2776 1576
rect 2808 1544 2848 1576
rect 2880 1544 2920 1576
rect 2952 1544 2992 1576
rect 3024 1544 3064 1576
rect 3096 1544 3136 1576
rect 3168 1544 3208 1576
rect 3240 1544 3280 1576
rect 3312 1544 3352 1576
rect 3384 1544 3424 1576
rect 3456 1544 3496 1576
rect 3528 1544 3568 1576
rect 3600 1544 3640 1576
rect 3672 1544 3712 1576
rect 3744 1544 3784 1576
rect 3816 1544 3856 1576
rect 3888 1544 3928 1576
rect 3960 1544 4000 1576
rect 0 1504 4000 1544
rect 0 1472 40 1504
rect 72 1472 112 1504
rect 144 1472 184 1504
rect 216 1472 256 1504
rect 288 1472 328 1504
rect 360 1472 400 1504
rect 432 1472 472 1504
rect 504 1472 544 1504
rect 576 1472 616 1504
rect 648 1472 688 1504
rect 720 1472 760 1504
rect 792 1472 832 1504
rect 864 1472 904 1504
rect 936 1472 976 1504
rect 1008 1472 1048 1504
rect 1080 1472 1120 1504
rect 1152 1472 1192 1504
rect 1224 1472 1264 1504
rect 1296 1472 1336 1504
rect 1368 1472 1408 1504
rect 1440 1472 1480 1504
rect 1512 1472 1552 1504
rect 1584 1472 1624 1504
rect 1656 1472 1696 1504
rect 1728 1472 1768 1504
rect 1800 1472 1840 1504
rect 1872 1472 1912 1504
rect 1944 1472 1984 1504
rect 2016 1472 2056 1504
rect 2088 1472 2128 1504
rect 2160 1472 2200 1504
rect 2232 1472 2272 1504
rect 2304 1472 2344 1504
rect 2376 1472 2416 1504
rect 2448 1472 2488 1504
rect 2520 1472 2560 1504
rect 2592 1472 2632 1504
rect 2664 1472 2704 1504
rect 2736 1472 2776 1504
rect 2808 1472 2848 1504
rect 2880 1472 2920 1504
rect 2952 1472 2992 1504
rect 3024 1472 3064 1504
rect 3096 1472 3136 1504
rect 3168 1472 3208 1504
rect 3240 1472 3280 1504
rect 3312 1472 3352 1504
rect 3384 1472 3424 1504
rect 3456 1472 3496 1504
rect 3528 1472 3568 1504
rect 3600 1472 3640 1504
rect 3672 1472 3712 1504
rect 3744 1472 3784 1504
rect 3816 1472 3856 1504
rect 3888 1472 3928 1504
rect 3960 1472 4000 1504
rect 0 1432 4000 1472
rect 0 1400 40 1432
rect 72 1400 112 1432
rect 144 1400 184 1432
rect 216 1400 256 1432
rect 288 1400 328 1432
rect 360 1400 400 1432
rect 432 1400 472 1432
rect 504 1400 544 1432
rect 576 1400 616 1432
rect 648 1400 688 1432
rect 720 1400 760 1432
rect 792 1400 832 1432
rect 864 1400 904 1432
rect 936 1400 976 1432
rect 1008 1400 1048 1432
rect 1080 1400 1120 1432
rect 1152 1400 1192 1432
rect 1224 1400 1264 1432
rect 1296 1400 1336 1432
rect 1368 1400 1408 1432
rect 1440 1400 1480 1432
rect 1512 1400 1552 1432
rect 1584 1400 1624 1432
rect 1656 1400 1696 1432
rect 1728 1400 1768 1432
rect 1800 1400 1840 1432
rect 1872 1400 1912 1432
rect 1944 1400 1984 1432
rect 2016 1400 2056 1432
rect 2088 1400 2128 1432
rect 2160 1400 2200 1432
rect 2232 1400 2272 1432
rect 2304 1400 2344 1432
rect 2376 1400 2416 1432
rect 2448 1400 2488 1432
rect 2520 1400 2560 1432
rect 2592 1400 2632 1432
rect 2664 1400 2704 1432
rect 2736 1400 2776 1432
rect 2808 1400 2848 1432
rect 2880 1400 2920 1432
rect 2952 1400 2992 1432
rect 3024 1400 3064 1432
rect 3096 1400 3136 1432
rect 3168 1400 3208 1432
rect 3240 1400 3280 1432
rect 3312 1400 3352 1432
rect 3384 1400 3424 1432
rect 3456 1400 3496 1432
rect 3528 1400 3568 1432
rect 3600 1400 3640 1432
rect 3672 1400 3712 1432
rect 3744 1400 3784 1432
rect 3816 1400 3856 1432
rect 3888 1400 3928 1432
rect 3960 1400 4000 1432
rect 0 1360 4000 1400
rect 0 1328 40 1360
rect 72 1328 112 1360
rect 144 1328 184 1360
rect 216 1328 256 1360
rect 288 1328 328 1360
rect 360 1328 400 1360
rect 432 1328 472 1360
rect 504 1328 544 1360
rect 576 1328 616 1360
rect 648 1328 688 1360
rect 720 1328 760 1360
rect 792 1328 832 1360
rect 864 1328 904 1360
rect 936 1328 976 1360
rect 1008 1328 1048 1360
rect 1080 1328 1120 1360
rect 1152 1328 1192 1360
rect 1224 1328 1264 1360
rect 1296 1328 1336 1360
rect 1368 1328 1408 1360
rect 1440 1328 1480 1360
rect 1512 1328 1552 1360
rect 1584 1328 1624 1360
rect 1656 1328 1696 1360
rect 1728 1328 1768 1360
rect 1800 1328 1840 1360
rect 1872 1328 1912 1360
rect 1944 1328 1984 1360
rect 2016 1328 2056 1360
rect 2088 1328 2128 1360
rect 2160 1328 2200 1360
rect 2232 1328 2272 1360
rect 2304 1328 2344 1360
rect 2376 1328 2416 1360
rect 2448 1328 2488 1360
rect 2520 1328 2560 1360
rect 2592 1328 2632 1360
rect 2664 1328 2704 1360
rect 2736 1328 2776 1360
rect 2808 1328 2848 1360
rect 2880 1328 2920 1360
rect 2952 1328 2992 1360
rect 3024 1328 3064 1360
rect 3096 1328 3136 1360
rect 3168 1328 3208 1360
rect 3240 1328 3280 1360
rect 3312 1328 3352 1360
rect 3384 1328 3424 1360
rect 3456 1328 3496 1360
rect 3528 1328 3568 1360
rect 3600 1328 3640 1360
rect 3672 1328 3712 1360
rect 3744 1328 3784 1360
rect 3816 1328 3856 1360
rect 3888 1328 3928 1360
rect 3960 1328 4000 1360
rect 0 1288 4000 1328
rect 0 1256 40 1288
rect 72 1256 112 1288
rect 144 1256 184 1288
rect 216 1256 256 1288
rect 288 1256 328 1288
rect 360 1256 400 1288
rect 432 1256 472 1288
rect 504 1256 544 1288
rect 576 1256 616 1288
rect 648 1256 688 1288
rect 720 1256 760 1288
rect 792 1256 832 1288
rect 864 1256 904 1288
rect 936 1256 976 1288
rect 1008 1256 1048 1288
rect 1080 1256 1120 1288
rect 1152 1256 1192 1288
rect 1224 1256 1264 1288
rect 1296 1256 1336 1288
rect 1368 1256 1408 1288
rect 1440 1256 1480 1288
rect 1512 1256 1552 1288
rect 1584 1256 1624 1288
rect 1656 1256 1696 1288
rect 1728 1256 1768 1288
rect 1800 1256 1840 1288
rect 1872 1256 1912 1288
rect 1944 1256 1984 1288
rect 2016 1256 2056 1288
rect 2088 1256 2128 1288
rect 2160 1256 2200 1288
rect 2232 1256 2272 1288
rect 2304 1256 2344 1288
rect 2376 1256 2416 1288
rect 2448 1256 2488 1288
rect 2520 1256 2560 1288
rect 2592 1256 2632 1288
rect 2664 1256 2704 1288
rect 2736 1256 2776 1288
rect 2808 1256 2848 1288
rect 2880 1256 2920 1288
rect 2952 1256 2992 1288
rect 3024 1256 3064 1288
rect 3096 1256 3136 1288
rect 3168 1256 3208 1288
rect 3240 1256 3280 1288
rect 3312 1256 3352 1288
rect 3384 1256 3424 1288
rect 3456 1256 3496 1288
rect 3528 1256 3568 1288
rect 3600 1256 3640 1288
rect 3672 1256 3712 1288
rect 3744 1256 3784 1288
rect 3816 1256 3856 1288
rect 3888 1256 3928 1288
rect 3960 1256 4000 1288
rect 0 1200 4000 1256
<< psubdiffcont >>
rect 112 31384 144 31416
rect 112 27939 144 27971
rect 112 22842 144 22874
rect 112 17816 144 17848
<< nsubdiffcont >>
rect 112 33384 144 33416
rect 112 29684 144 29716
rect 40 12112 72 12144
rect 40 6512 72 6544
<< metal1 >>
rect 184 33384 216 33416
rect 256 33384 288 33416
rect 328 33384 360 33416
rect 400 33384 432 33416
rect 472 33384 504 33416
rect 544 33384 576 33416
rect 616 33384 648 33416
rect 688 33384 720 33416
rect 760 33384 792 33416
rect 832 33384 864 33416
rect 904 33384 936 33416
rect 976 33384 1008 33416
rect 1048 33384 1080 33416
rect 1120 33384 1152 33416
rect 1192 33384 1224 33416
rect 1264 33384 1296 33416
rect 1336 33384 1368 33416
rect 1408 33384 1440 33416
rect 1480 33384 1512 33416
rect 1552 33384 1584 33416
rect 1624 33384 1656 33416
rect 1696 33384 1728 33416
rect 1768 33384 1800 33416
rect 1840 33384 1872 33416
rect 1912 33384 1944 33416
rect 1984 33384 2016 33416
rect 2056 33384 2088 33416
rect 2128 33384 2160 33416
rect 2200 33384 2232 33416
rect 2272 33384 2304 33416
rect 2344 33384 2376 33416
rect 2416 33384 2448 33416
rect 2488 33384 2520 33416
rect 2560 33384 2592 33416
rect 2632 33384 2664 33416
rect 2704 33384 2736 33416
rect 2776 33384 2808 33416
rect 2848 33384 2880 33416
rect 2920 33384 2952 33416
rect 2992 33384 3024 33416
rect 3064 33384 3096 33416
rect 3136 33384 3168 33416
rect 3208 33384 3240 33416
rect 3280 33384 3312 33416
rect 3352 33384 3384 33416
rect 3424 33384 3456 33416
rect 3496 33384 3528 33416
rect 3568 33384 3600 33416
rect 3640 33384 3672 33416
rect 3712 33384 3744 33416
rect 3784 33384 3816 33416
rect 3856 33384 3888 33416
rect 184 29684 216 29716
rect 256 29684 288 29716
rect 328 29684 360 29716
rect 400 29684 432 29716
rect 472 29684 504 29716
rect 544 29684 576 29716
rect 616 29684 648 29716
rect 688 29684 720 29716
rect 760 29684 792 29716
rect 832 29684 864 29716
rect 904 29684 936 29716
rect 976 29684 1008 29716
rect 1048 29684 1080 29716
rect 1120 29684 1152 29716
rect 1192 29684 1224 29716
rect 1264 29684 1296 29716
rect 1336 29684 1368 29716
rect 1408 29684 1440 29716
rect 1480 29684 1512 29716
rect 1552 29684 1584 29716
rect 1624 29684 1656 29716
rect 1696 29684 1728 29716
rect 1768 29684 1800 29716
rect 1840 29684 1872 29716
rect 1912 29684 1944 29716
rect 1984 29684 2016 29716
rect 2056 29684 2088 29716
rect 2128 29684 2160 29716
rect 2200 29684 2232 29716
rect 2272 29684 2304 29716
rect 2344 29684 2376 29716
rect 2416 29684 2448 29716
rect 2488 29684 2520 29716
rect 2560 29684 2592 29716
rect 2632 29684 2664 29716
rect 2704 29684 2736 29716
rect 2776 29684 2808 29716
rect 2848 29684 2880 29716
rect 2920 29684 2952 29716
rect 2992 29684 3024 29716
rect 3064 29684 3096 29716
rect 3136 29684 3168 29716
rect 3208 29684 3240 29716
rect 3280 29684 3312 29716
rect 3352 29684 3384 29716
rect 3424 29684 3456 29716
rect 3496 29684 3528 29716
rect 3568 29684 3600 29716
rect 3640 29684 3672 29716
rect 3712 29684 3744 29716
rect 3784 29684 3816 29716
rect 3856 29684 3888 29716
rect 112 12112 144 12144
rect 184 12112 216 12144
rect 256 12112 288 12144
rect 328 12112 360 12144
rect 400 12112 432 12144
rect 472 12112 504 12144
rect 544 12112 576 12144
rect 616 12112 648 12144
rect 688 12112 720 12144
rect 760 12112 792 12144
rect 832 12112 864 12144
rect 904 12112 936 12144
rect 976 12112 1008 12144
rect 1048 12112 1080 12144
rect 1120 12112 1152 12144
rect 1192 12112 1224 12144
rect 1264 12112 1296 12144
rect 1336 12112 1368 12144
rect 1408 12112 1440 12144
rect 1480 12112 1512 12144
rect 1552 12112 1584 12144
rect 1624 12112 1656 12144
rect 1696 12112 1728 12144
rect 1768 12112 1800 12144
rect 1840 12112 1872 12144
rect 1912 12112 1944 12144
rect 1984 12112 2016 12144
rect 2056 12112 2088 12144
rect 2128 12112 2160 12144
rect 2200 12112 2232 12144
rect 2272 12112 2304 12144
rect 2344 12112 2376 12144
rect 2416 12112 2448 12144
rect 2488 12112 2520 12144
rect 2560 12112 2592 12144
rect 2632 12112 2664 12144
rect 2704 12112 2736 12144
rect 2776 12112 2808 12144
rect 2848 12112 2880 12144
rect 2920 12112 2952 12144
rect 2992 12112 3024 12144
rect 3064 12112 3096 12144
rect 3136 12112 3168 12144
rect 3208 12112 3240 12144
rect 3280 12112 3312 12144
rect 3352 12112 3384 12144
rect 3424 12112 3456 12144
rect 3496 12112 3528 12144
rect 3568 12112 3600 12144
rect 3640 12112 3672 12144
rect 3712 12112 3744 12144
rect 3784 12112 3816 12144
rect 3856 12112 3888 12144
rect 3928 12112 3960 12144
rect 40 12040 72 12072
rect 112 12040 144 12072
rect 184 12040 216 12072
rect 256 12040 288 12072
rect 328 12040 360 12072
rect 400 12040 432 12072
rect 472 12040 504 12072
rect 544 12040 576 12072
rect 616 12040 648 12072
rect 688 12040 720 12072
rect 760 12040 792 12072
rect 832 12040 864 12072
rect 904 12040 936 12072
rect 976 12040 1008 12072
rect 1048 12040 1080 12072
rect 1120 12040 1152 12072
rect 1192 12040 1224 12072
rect 1264 12040 1296 12072
rect 1336 12040 1368 12072
rect 1408 12040 1440 12072
rect 1480 12040 1512 12072
rect 1552 12040 1584 12072
rect 1624 12040 1656 12072
rect 1696 12040 1728 12072
rect 1768 12040 1800 12072
rect 1840 12040 1872 12072
rect 1912 12040 1944 12072
rect 1984 12040 2016 12072
rect 2056 12040 2088 12072
rect 2128 12040 2160 12072
rect 2200 12040 2232 12072
rect 2272 12040 2304 12072
rect 2344 12040 2376 12072
rect 2416 12040 2448 12072
rect 2488 12040 2520 12072
rect 2560 12040 2592 12072
rect 2632 12040 2664 12072
rect 2704 12040 2736 12072
rect 2776 12040 2808 12072
rect 2848 12040 2880 12072
rect 2920 12040 2952 12072
rect 2992 12040 3024 12072
rect 3064 12040 3096 12072
rect 3136 12040 3168 12072
rect 3208 12040 3240 12072
rect 3280 12040 3312 12072
rect 3352 12040 3384 12072
rect 3424 12040 3456 12072
rect 3496 12040 3528 12072
rect 3568 12040 3600 12072
rect 3640 12040 3672 12072
rect 3712 12040 3744 12072
rect 3784 12040 3816 12072
rect 3856 12040 3888 12072
rect 3928 12040 3960 12072
rect 40 11968 72 12000
rect 112 11968 144 12000
rect 184 11968 216 12000
rect 256 11968 288 12000
rect 328 11968 360 12000
rect 400 11968 432 12000
rect 472 11968 504 12000
rect 544 11968 576 12000
rect 616 11968 648 12000
rect 688 11968 720 12000
rect 760 11968 792 12000
rect 832 11968 864 12000
rect 904 11968 936 12000
rect 976 11968 1008 12000
rect 1048 11968 1080 12000
rect 1120 11968 1152 12000
rect 1192 11968 1224 12000
rect 1264 11968 1296 12000
rect 1336 11968 1368 12000
rect 1408 11968 1440 12000
rect 1480 11968 1512 12000
rect 1552 11968 1584 12000
rect 1624 11968 1656 12000
rect 1696 11968 1728 12000
rect 1768 11968 1800 12000
rect 1840 11968 1872 12000
rect 1912 11968 1944 12000
rect 1984 11968 2016 12000
rect 2056 11968 2088 12000
rect 2128 11968 2160 12000
rect 2200 11968 2232 12000
rect 2272 11968 2304 12000
rect 2344 11968 2376 12000
rect 2416 11968 2448 12000
rect 2488 11968 2520 12000
rect 2560 11968 2592 12000
rect 2632 11968 2664 12000
rect 2704 11968 2736 12000
rect 2776 11968 2808 12000
rect 2848 11968 2880 12000
rect 2920 11968 2952 12000
rect 2992 11968 3024 12000
rect 3064 11968 3096 12000
rect 3136 11968 3168 12000
rect 3208 11968 3240 12000
rect 3280 11968 3312 12000
rect 3352 11968 3384 12000
rect 3424 11968 3456 12000
rect 3496 11968 3528 12000
rect 3568 11968 3600 12000
rect 3640 11968 3672 12000
rect 3712 11968 3744 12000
rect 3784 11968 3816 12000
rect 3856 11968 3888 12000
rect 3928 11968 3960 12000
rect 40 11896 72 11928
rect 112 11896 144 11928
rect 184 11896 216 11928
rect 256 11896 288 11928
rect 328 11896 360 11928
rect 400 11896 432 11928
rect 472 11896 504 11928
rect 544 11896 576 11928
rect 616 11896 648 11928
rect 688 11896 720 11928
rect 760 11896 792 11928
rect 832 11896 864 11928
rect 904 11896 936 11928
rect 976 11896 1008 11928
rect 1048 11896 1080 11928
rect 1120 11896 1152 11928
rect 1192 11896 1224 11928
rect 1264 11896 1296 11928
rect 1336 11896 1368 11928
rect 1408 11896 1440 11928
rect 1480 11896 1512 11928
rect 1552 11896 1584 11928
rect 1624 11896 1656 11928
rect 1696 11896 1728 11928
rect 1768 11896 1800 11928
rect 1840 11896 1872 11928
rect 1912 11896 1944 11928
rect 1984 11896 2016 11928
rect 2056 11896 2088 11928
rect 2128 11896 2160 11928
rect 2200 11896 2232 11928
rect 2272 11896 2304 11928
rect 2344 11896 2376 11928
rect 2416 11896 2448 11928
rect 2488 11896 2520 11928
rect 2560 11896 2592 11928
rect 2632 11896 2664 11928
rect 2704 11896 2736 11928
rect 2776 11896 2808 11928
rect 2848 11896 2880 11928
rect 2920 11896 2952 11928
rect 2992 11896 3024 11928
rect 3064 11896 3096 11928
rect 3136 11896 3168 11928
rect 3208 11896 3240 11928
rect 3280 11896 3312 11928
rect 3352 11896 3384 11928
rect 3424 11896 3456 11928
rect 3496 11896 3528 11928
rect 3568 11896 3600 11928
rect 3640 11896 3672 11928
rect 3712 11896 3744 11928
rect 3784 11896 3816 11928
rect 3856 11896 3888 11928
rect 3928 11896 3960 11928
rect 40 11824 72 11856
rect 112 11824 144 11856
rect 184 11824 216 11856
rect 256 11824 288 11856
rect 328 11824 360 11856
rect 400 11824 432 11856
rect 472 11824 504 11856
rect 544 11824 576 11856
rect 616 11824 648 11856
rect 688 11824 720 11856
rect 760 11824 792 11856
rect 832 11824 864 11856
rect 904 11824 936 11856
rect 976 11824 1008 11856
rect 1048 11824 1080 11856
rect 1120 11824 1152 11856
rect 1192 11824 1224 11856
rect 1264 11824 1296 11856
rect 1336 11824 1368 11856
rect 1408 11824 1440 11856
rect 1480 11824 1512 11856
rect 1552 11824 1584 11856
rect 1624 11824 1656 11856
rect 1696 11824 1728 11856
rect 1768 11824 1800 11856
rect 1840 11824 1872 11856
rect 1912 11824 1944 11856
rect 1984 11824 2016 11856
rect 2056 11824 2088 11856
rect 2128 11824 2160 11856
rect 2200 11824 2232 11856
rect 2272 11824 2304 11856
rect 2344 11824 2376 11856
rect 2416 11824 2448 11856
rect 2488 11824 2520 11856
rect 2560 11824 2592 11856
rect 2632 11824 2664 11856
rect 2704 11824 2736 11856
rect 2776 11824 2808 11856
rect 2848 11824 2880 11856
rect 2920 11824 2952 11856
rect 2992 11824 3024 11856
rect 3064 11824 3096 11856
rect 3136 11824 3168 11856
rect 3208 11824 3240 11856
rect 3280 11824 3312 11856
rect 3352 11824 3384 11856
rect 3424 11824 3456 11856
rect 3496 11824 3528 11856
rect 3568 11824 3600 11856
rect 3640 11824 3672 11856
rect 3712 11824 3744 11856
rect 3784 11824 3816 11856
rect 3856 11824 3888 11856
rect 3928 11824 3960 11856
rect 40 11752 72 11784
rect 112 11752 144 11784
rect 184 11752 216 11784
rect 256 11752 288 11784
rect 328 11752 360 11784
rect 400 11752 432 11784
rect 472 11752 504 11784
rect 544 11752 576 11784
rect 616 11752 648 11784
rect 688 11752 720 11784
rect 760 11752 792 11784
rect 832 11752 864 11784
rect 904 11752 936 11784
rect 976 11752 1008 11784
rect 1048 11752 1080 11784
rect 1120 11752 1152 11784
rect 1192 11752 1224 11784
rect 1264 11752 1296 11784
rect 1336 11752 1368 11784
rect 1408 11752 1440 11784
rect 1480 11752 1512 11784
rect 1552 11752 1584 11784
rect 1624 11752 1656 11784
rect 1696 11752 1728 11784
rect 1768 11752 1800 11784
rect 1840 11752 1872 11784
rect 1912 11752 1944 11784
rect 1984 11752 2016 11784
rect 2056 11752 2088 11784
rect 2128 11752 2160 11784
rect 2200 11752 2232 11784
rect 2272 11752 2304 11784
rect 2344 11752 2376 11784
rect 2416 11752 2448 11784
rect 2488 11752 2520 11784
rect 2560 11752 2592 11784
rect 2632 11752 2664 11784
rect 2704 11752 2736 11784
rect 2776 11752 2808 11784
rect 2848 11752 2880 11784
rect 2920 11752 2952 11784
rect 2992 11752 3024 11784
rect 3064 11752 3096 11784
rect 3136 11752 3168 11784
rect 3208 11752 3240 11784
rect 3280 11752 3312 11784
rect 3352 11752 3384 11784
rect 3424 11752 3456 11784
rect 3496 11752 3528 11784
rect 3568 11752 3600 11784
rect 3640 11752 3672 11784
rect 3712 11752 3744 11784
rect 3784 11752 3816 11784
rect 3856 11752 3888 11784
rect 3928 11752 3960 11784
rect 40 11680 72 11712
rect 112 11680 144 11712
rect 184 11680 216 11712
rect 256 11680 288 11712
rect 328 11680 360 11712
rect 400 11680 432 11712
rect 472 11680 504 11712
rect 544 11680 576 11712
rect 616 11680 648 11712
rect 688 11680 720 11712
rect 760 11680 792 11712
rect 832 11680 864 11712
rect 904 11680 936 11712
rect 976 11680 1008 11712
rect 1048 11680 1080 11712
rect 1120 11680 1152 11712
rect 1192 11680 1224 11712
rect 1264 11680 1296 11712
rect 1336 11680 1368 11712
rect 1408 11680 1440 11712
rect 1480 11680 1512 11712
rect 1552 11680 1584 11712
rect 1624 11680 1656 11712
rect 1696 11680 1728 11712
rect 1768 11680 1800 11712
rect 1840 11680 1872 11712
rect 1912 11680 1944 11712
rect 1984 11680 2016 11712
rect 2056 11680 2088 11712
rect 2128 11680 2160 11712
rect 2200 11680 2232 11712
rect 2272 11680 2304 11712
rect 2344 11680 2376 11712
rect 2416 11680 2448 11712
rect 2488 11680 2520 11712
rect 2560 11680 2592 11712
rect 2632 11680 2664 11712
rect 2704 11680 2736 11712
rect 2776 11680 2808 11712
rect 2848 11680 2880 11712
rect 2920 11680 2952 11712
rect 2992 11680 3024 11712
rect 3064 11680 3096 11712
rect 3136 11680 3168 11712
rect 3208 11680 3240 11712
rect 3280 11680 3312 11712
rect 3352 11680 3384 11712
rect 3424 11680 3456 11712
rect 3496 11680 3528 11712
rect 3568 11680 3600 11712
rect 3640 11680 3672 11712
rect 3712 11680 3744 11712
rect 3784 11680 3816 11712
rect 3856 11680 3888 11712
rect 3928 11680 3960 11712
rect 40 11608 72 11640
rect 112 11608 144 11640
rect 184 11608 216 11640
rect 256 11608 288 11640
rect 328 11608 360 11640
rect 400 11608 432 11640
rect 472 11608 504 11640
rect 544 11608 576 11640
rect 616 11608 648 11640
rect 688 11608 720 11640
rect 760 11608 792 11640
rect 832 11608 864 11640
rect 904 11608 936 11640
rect 976 11608 1008 11640
rect 1048 11608 1080 11640
rect 1120 11608 1152 11640
rect 1192 11608 1224 11640
rect 1264 11608 1296 11640
rect 1336 11608 1368 11640
rect 1408 11608 1440 11640
rect 1480 11608 1512 11640
rect 1552 11608 1584 11640
rect 1624 11608 1656 11640
rect 1696 11608 1728 11640
rect 1768 11608 1800 11640
rect 1840 11608 1872 11640
rect 1912 11608 1944 11640
rect 1984 11608 2016 11640
rect 2056 11608 2088 11640
rect 2128 11608 2160 11640
rect 2200 11608 2232 11640
rect 2272 11608 2304 11640
rect 2344 11608 2376 11640
rect 2416 11608 2448 11640
rect 2488 11608 2520 11640
rect 2560 11608 2592 11640
rect 2632 11608 2664 11640
rect 2704 11608 2736 11640
rect 2776 11608 2808 11640
rect 2848 11608 2880 11640
rect 2920 11608 2952 11640
rect 2992 11608 3024 11640
rect 3064 11608 3096 11640
rect 3136 11608 3168 11640
rect 3208 11608 3240 11640
rect 3280 11608 3312 11640
rect 3352 11608 3384 11640
rect 3424 11608 3456 11640
rect 3496 11608 3528 11640
rect 3568 11608 3600 11640
rect 3640 11608 3672 11640
rect 3712 11608 3744 11640
rect 3784 11608 3816 11640
rect 3856 11608 3888 11640
rect 3928 11608 3960 11640
rect 40 11536 72 11568
rect 112 11536 144 11568
rect 184 11536 216 11568
rect 256 11536 288 11568
rect 328 11536 360 11568
rect 400 11536 432 11568
rect 472 11536 504 11568
rect 544 11536 576 11568
rect 616 11536 648 11568
rect 688 11536 720 11568
rect 760 11536 792 11568
rect 832 11536 864 11568
rect 904 11536 936 11568
rect 976 11536 1008 11568
rect 1048 11536 1080 11568
rect 1120 11536 1152 11568
rect 1192 11536 1224 11568
rect 1264 11536 1296 11568
rect 1336 11536 1368 11568
rect 1408 11536 1440 11568
rect 1480 11536 1512 11568
rect 1552 11536 1584 11568
rect 1624 11536 1656 11568
rect 1696 11536 1728 11568
rect 1768 11536 1800 11568
rect 1840 11536 1872 11568
rect 1912 11536 1944 11568
rect 1984 11536 2016 11568
rect 2056 11536 2088 11568
rect 2128 11536 2160 11568
rect 2200 11536 2232 11568
rect 2272 11536 2304 11568
rect 2344 11536 2376 11568
rect 2416 11536 2448 11568
rect 2488 11536 2520 11568
rect 2560 11536 2592 11568
rect 2632 11536 2664 11568
rect 2704 11536 2736 11568
rect 2776 11536 2808 11568
rect 2848 11536 2880 11568
rect 2920 11536 2952 11568
rect 2992 11536 3024 11568
rect 3064 11536 3096 11568
rect 3136 11536 3168 11568
rect 3208 11536 3240 11568
rect 3280 11536 3312 11568
rect 3352 11536 3384 11568
rect 3424 11536 3456 11568
rect 3496 11536 3528 11568
rect 3568 11536 3600 11568
rect 3640 11536 3672 11568
rect 3712 11536 3744 11568
rect 3784 11536 3816 11568
rect 3856 11536 3888 11568
rect 3928 11536 3960 11568
rect 40 11464 72 11496
rect 112 11464 144 11496
rect 184 11464 216 11496
rect 256 11464 288 11496
rect 328 11464 360 11496
rect 400 11464 432 11496
rect 472 11464 504 11496
rect 544 11464 576 11496
rect 616 11464 648 11496
rect 688 11464 720 11496
rect 760 11464 792 11496
rect 832 11464 864 11496
rect 904 11464 936 11496
rect 976 11464 1008 11496
rect 1048 11464 1080 11496
rect 1120 11464 1152 11496
rect 1192 11464 1224 11496
rect 1264 11464 1296 11496
rect 1336 11464 1368 11496
rect 1408 11464 1440 11496
rect 1480 11464 1512 11496
rect 1552 11464 1584 11496
rect 1624 11464 1656 11496
rect 1696 11464 1728 11496
rect 1768 11464 1800 11496
rect 1840 11464 1872 11496
rect 1912 11464 1944 11496
rect 1984 11464 2016 11496
rect 2056 11464 2088 11496
rect 2128 11464 2160 11496
rect 2200 11464 2232 11496
rect 2272 11464 2304 11496
rect 2344 11464 2376 11496
rect 2416 11464 2448 11496
rect 2488 11464 2520 11496
rect 2560 11464 2592 11496
rect 2632 11464 2664 11496
rect 2704 11464 2736 11496
rect 2776 11464 2808 11496
rect 2848 11464 2880 11496
rect 2920 11464 2952 11496
rect 2992 11464 3024 11496
rect 3064 11464 3096 11496
rect 3136 11464 3168 11496
rect 3208 11464 3240 11496
rect 3280 11464 3312 11496
rect 3352 11464 3384 11496
rect 3424 11464 3456 11496
rect 3496 11464 3528 11496
rect 3568 11464 3600 11496
rect 3640 11464 3672 11496
rect 3712 11464 3744 11496
rect 3784 11464 3816 11496
rect 3856 11464 3888 11496
rect 3928 11464 3960 11496
rect 40 11392 72 11424
rect 112 11392 144 11424
rect 184 11392 216 11424
rect 256 11392 288 11424
rect 328 11392 360 11424
rect 400 11392 432 11424
rect 472 11392 504 11424
rect 544 11392 576 11424
rect 616 11392 648 11424
rect 688 11392 720 11424
rect 760 11392 792 11424
rect 832 11392 864 11424
rect 904 11392 936 11424
rect 976 11392 1008 11424
rect 1048 11392 1080 11424
rect 1120 11392 1152 11424
rect 1192 11392 1224 11424
rect 1264 11392 1296 11424
rect 1336 11392 1368 11424
rect 1408 11392 1440 11424
rect 1480 11392 1512 11424
rect 1552 11392 1584 11424
rect 1624 11392 1656 11424
rect 1696 11392 1728 11424
rect 1768 11392 1800 11424
rect 1840 11392 1872 11424
rect 1912 11392 1944 11424
rect 1984 11392 2016 11424
rect 2056 11392 2088 11424
rect 2128 11392 2160 11424
rect 2200 11392 2232 11424
rect 2272 11392 2304 11424
rect 2344 11392 2376 11424
rect 2416 11392 2448 11424
rect 2488 11392 2520 11424
rect 2560 11392 2592 11424
rect 2632 11392 2664 11424
rect 2704 11392 2736 11424
rect 2776 11392 2808 11424
rect 2848 11392 2880 11424
rect 2920 11392 2952 11424
rect 2992 11392 3024 11424
rect 3064 11392 3096 11424
rect 3136 11392 3168 11424
rect 3208 11392 3240 11424
rect 3280 11392 3312 11424
rect 3352 11392 3384 11424
rect 3424 11392 3456 11424
rect 3496 11392 3528 11424
rect 3568 11392 3600 11424
rect 3640 11392 3672 11424
rect 3712 11392 3744 11424
rect 3784 11392 3816 11424
rect 3856 11392 3888 11424
rect 3928 11392 3960 11424
rect 40 11320 72 11352
rect 112 11320 144 11352
rect 184 11320 216 11352
rect 256 11320 288 11352
rect 328 11320 360 11352
rect 400 11320 432 11352
rect 472 11320 504 11352
rect 544 11320 576 11352
rect 616 11320 648 11352
rect 688 11320 720 11352
rect 760 11320 792 11352
rect 832 11320 864 11352
rect 904 11320 936 11352
rect 976 11320 1008 11352
rect 1048 11320 1080 11352
rect 1120 11320 1152 11352
rect 1192 11320 1224 11352
rect 1264 11320 1296 11352
rect 1336 11320 1368 11352
rect 1408 11320 1440 11352
rect 1480 11320 1512 11352
rect 1552 11320 1584 11352
rect 1624 11320 1656 11352
rect 1696 11320 1728 11352
rect 1768 11320 1800 11352
rect 1840 11320 1872 11352
rect 1912 11320 1944 11352
rect 1984 11320 2016 11352
rect 2056 11320 2088 11352
rect 2128 11320 2160 11352
rect 2200 11320 2232 11352
rect 2272 11320 2304 11352
rect 2344 11320 2376 11352
rect 2416 11320 2448 11352
rect 2488 11320 2520 11352
rect 2560 11320 2592 11352
rect 2632 11320 2664 11352
rect 2704 11320 2736 11352
rect 2776 11320 2808 11352
rect 2848 11320 2880 11352
rect 2920 11320 2952 11352
rect 2992 11320 3024 11352
rect 3064 11320 3096 11352
rect 3136 11320 3168 11352
rect 3208 11320 3240 11352
rect 3280 11320 3312 11352
rect 3352 11320 3384 11352
rect 3424 11320 3456 11352
rect 3496 11320 3528 11352
rect 3568 11320 3600 11352
rect 3640 11320 3672 11352
rect 3712 11320 3744 11352
rect 3784 11320 3816 11352
rect 3856 11320 3888 11352
rect 3928 11320 3960 11352
rect 40 11248 72 11280
rect 112 11248 144 11280
rect 184 11248 216 11280
rect 256 11248 288 11280
rect 328 11248 360 11280
rect 400 11248 432 11280
rect 472 11248 504 11280
rect 544 11248 576 11280
rect 616 11248 648 11280
rect 688 11248 720 11280
rect 760 11248 792 11280
rect 832 11248 864 11280
rect 904 11248 936 11280
rect 976 11248 1008 11280
rect 1048 11248 1080 11280
rect 1120 11248 1152 11280
rect 1192 11248 1224 11280
rect 1264 11248 1296 11280
rect 1336 11248 1368 11280
rect 1408 11248 1440 11280
rect 1480 11248 1512 11280
rect 1552 11248 1584 11280
rect 1624 11248 1656 11280
rect 1696 11248 1728 11280
rect 1768 11248 1800 11280
rect 1840 11248 1872 11280
rect 1912 11248 1944 11280
rect 1984 11248 2016 11280
rect 2056 11248 2088 11280
rect 2128 11248 2160 11280
rect 2200 11248 2232 11280
rect 2272 11248 2304 11280
rect 2344 11248 2376 11280
rect 2416 11248 2448 11280
rect 2488 11248 2520 11280
rect 2560 11248 2592 11280
rect 2632 11248 2664 11280
rect 2704 11248 2736 11280
rect 2776 11248 2808 11280
rect 2848 11248 2880 11280
rect 2920 11248 2952 11280
rect 2992 11248 3024 11280
rect 3064 11248 3096 11280
rect 3136 11248 3168 11280
rect 3208 11248 3240 11280
rect 3280 11248 3312 11280
rect 3352 11248 3384 11280
rect 3424 11248 3456 11280
rect 3496 11248 3528 11280
rect 3568 11248 3600 11280
rect 3640 11248 3672 11280
rect 3712 11248 3744 11280
rect 3784 11248 3816 11280
rect 3856 11248 3888 11280
rect 3928 11248 3960 11280
rect 40 11176 72 11208
rect 112 11176 144 11208
rect 184 11176 216 11208
rect 256 11176 288 11208
rect 328 11176 360 11208
rect 400 11176 432 11208
rect 472 11176 504 11208
rect 544 11176 576 11208
rect 616 11176 648 11208
rect 688 11176 720 11208
rect 760 11176 792 11208
rect 832 11176 864 11208
rect 904 11176 936 11208
rect 976 11176 1008 11208
rect 1048 11176 1080 11208
rect 1120 11176 1152 11208
rect 1192 11176 1224 11208
rect 1264 11176 1296 11208
rect 1336 11176 1368 11208
rect 1408 11176 1440 11208
rect 1480 11176 1512 11208
rect 1552 11176 1584 11208
rect 1624 11176 1656 11208
rect 1696 11176 1728 11208
rect 1768 11176 1800 11208
rect 1840 11176 1872 11208
rect 1912 11176 1944 11208
rect 1984 11176 2016 11208
rect 2056 11176 2088 11208
rect 2128 11176 2160 11208
rect 2200 11176 2232 11208
rect 2272 11176 2304 11208
rect 2344 11176 2376 11208
rect 2416 11176 2448 11208
rect 2488 11176 2520 11208
rect 2560 11176 2592 11208
rect 2632 11176 2664 11208
rect 2704 11176 2736 11208
rect 2776 11176 2808 11208
rect 2848 11176 2880 11208
rect 2920 11176 2952 11208
rect 2992 11176 3024 11208
rect 3064 11176 3096 11208
rect 3136 11176 3168 11208
rect 3208 11176 3240 11208
rect 3280 11176 3312 11208
rect 3352 11176 3384 11208
rect 3424 11176 3456 11208
rect 3496 11176 3528 11208
rect 3568 11176 3600 11208
rect 3640 11176 3672 11208
rect 3712 11176 3744 11208
rect 3784 11176 3816 11208
rect 3856 11176 3888 11208
rect 3928 11176 3960 11208
rect 40 11104 72 11136
rect 112 11104 144 11136
rect 184 11104 216 11136
rect 256 11104 288 11136
rect 328 11104 360 11136
rect 400 11104 432 11136
rect 472 11104 504 11136
rect 544 11104 576 11136
rect 616 11104 648 11136
rect 688 11104 720 11136
rect 760 11104 792 11136
rect 832 11104 864 11136
rect 904 11104 936 11136
rect 976 11104 1008 11136
rect 1048 11104 1080 11136
rect 1120 11104 1152 11136
rect 1192 11104 1224 11136
rect 1264 11104 1296 11136
rect 1336 11104 1368 11136
rect 1408 11104 1440 11136
rect 1480 11104 1512 11136
rect 1552 11104 1584 11136
rect 1624 11104 1656 11136
rect 1696 11104 1728 11136
rect 1768 11104 1800 11136
rect 1840 11104 1872 11136
rect 1912 11104 1944 11136
rect 1984 11104 2016 11136
rect 2056 11104 2088 11136
rect 2128 11104 2160 11136
rect 2200 11104 2232 11136
rect 2272 11104 2304 11136
rect 2344 11104 2376 11136
rect 2416 11104 2448 11136
rect 2488 11104 2520 11136
rect 2560 11104 2592 11136
rect 2632 11104 2664 11136
rect 2704 11104 2736 11136
rect 2776 11104 2808 11136
rect 2848 11104 2880 11136
rect 2920 11104 2952 11136
rect 2992 11104 3024 11136
rect 3064 11104 3096 11136
rect 3136 11104 3168 11136
rect 3208 11104 3240 11136
rect 3280 11104 3312 11136
rect 3352 11104 3384 11136
rect 3424 11104 3456 11136
rect 3496 11104 3528 11136
rect 3568 11104 3600 11136
rect 3640 11104 3672 11136
rect 3712 11104 3744 11136
rect 3784 11104 3816 11136
rect 3856 11104 3888 11136
rect 3928 11104 3960 11136
rect 40 11032 72 11064
rect 112 11032 144 11064
rect 184 11032 216 11064
rect 256 11032 288 11064
rect 328 11032 360 11064
rect 400 11032 432 11064
rect 472 11032 504 11064
rect 544 11032 576 11064
rect 616 11032 648 11064
rect 688 11032 720 11064
rect 760 11032 792 11064
rect 832 11032 864 11064
rect 904 11032 936 11064
rect 976 11032 1008 11064
rect 1048 11032 1080 11064
rect 1120 11032 1152 11064
rect 1192 11032 1224 11064
rect 1264 11032 1296 11064
rect 1336 11032 1368 11064
rect 1408 11032 1440 11064
rect 1480 11032 1512 11064
rect 1552 11032 1584 11064
rect 1624 11032 1656 11064
rect 1696 11032 1728 11064
rect 1768 11032 1800 11064
rect 1840 11032 1872 11064
rect 1912 11032 1944 11064
rect 1984 11032 2016 11064
rect 2056 11032 2088 11064
rect 2128 11032 2160 11064
rect 2200 11032 2232 11064
rect 2272 11032 2304 11064
rect 2344 11032 2376 11064
rect 2416 11032 2448 11064
rect 2488 11032 2520 11064
rect 2560 11032 2592 11064
rect 2632 11032 2664 11064
rect 2704 11032 2736 11064
rect 2776 11032 2808 11064
rect 2848 11032 2880 11064
rect 2920 11032 2952 11064
rect 2992 11032 3024 11064
rect 3064 11032 3096 11064
rect 3136 11032 3168 11064
rect 3208 11032 3240 11064
rect 3280 11032 3312 11064
rect 3352 11032 3384 11064
rect 3424 11032 3456 11064
rect 3496 11032 3528 11064
rect 3568 11032 3600 11064
rect 3640 11032 3672 11064
rect 3712 11032 3744 11064
rect 3784 11032 3816 11064
rect 3856 11032 3888 11064
rect 3928 11032 3960 11064
rect 40 10960 72 10992
rect 112 10960 144 10992
rect 184 10960 216 10992
rect 256 10960 288 10992
rect 328 10960 360 10992
rect 400 10960 432 10992
rect 472 10960 504 10992
rect 544 10960 576 10992
rect 616 10960 648 10992
rect 688 10960 720 10992
rect 760 10960 792 10992
rect 832 10960 864 10992
rect 904 10960 936 10992
rect 976 10960 1008 10992
rect 1048 10960 1080 10992
rect 1120 10960 1152 10992
rect 1192 10960 1224 10992
rect 1264 10960 1296 10992
rect 1336 10960 1368 10992
rect 1408 10960 1440 10992
rect 1480 10960 1512 10992
rect 1552 10960 1584 10992
rect 1624 10960 1656 10992
rect 1696 10960 1728 10992
rect 1768 10960 1800 10992
rect 1840 10960 1872 10992
rect 1912 10960 1944 10992
rect 1984 10960 2016 10992
rect 2056 10960 2088 10992
rect 2128 10960 2160 10992
rect 2200 10960 2232 10992
rect 2272 10960 2304 10992
rect 2344 10960 2376 10992
rect 2416 10960 2448 10992
rect 2488 10960 2520 10992
rect 2560 10960 2592 10992
rect 2632 10960 2664 10992
rect 2704 10960 2736 10992
rect 2776 10960 2808 10992
rect 2848 10960 2880 10992
rect 2920 10960 2952 10992
rect 2992 10960 3024 10992
rect 3064 10960 3096 10992
rect 3136 10960 3168 10992
rect 3208 10960 3240 10992
rect 3280 10960 3312 10992
rect 3352 10960 3384 10992
rect 3424 10960 3456 10992
rect 3496 10960 3528 10992
rect 3568 10960 3600 10992
rect 3640 10960 3672 10992
rect 3712 10960 3744 10992
rect 3784 10960 3816 10992
rect 3856 10960 3888 10992
rect 3928 10960 3960 10992
rect 40 10888 72 10920
rect 112 10888 144 10920
rect 184 10888 216 10920
rect 256 10888 288 10920
rect 328 10888 360 10920
rect 400 10888 432 10920
rect 472 10888 504 10920
rect 544 10888 576 10920
rect 616 10888 648 10920
rect 688 10888 720 10920
rect 760 10888 792 10920
rect 832 10888 864 10920
rect 904 10888 936 10920
rect 976 10888 1008 10920
rect 1048 10888 1080 10920
rect 1120 10888 1152 10920
rect 1192 10888 1224 10920
rect 1264 10888 1296 10920
rect 1336 10888 1368 10920
rect 1408 10888 1440 10920
rect 1480 10888 1512 10920
rect 1552 10888 1584 10920
rect 1624 10888 1656 10920
rect 1696 10888 1728 10920
rect 1768 10888 1800 10920
rect 1840 10888 1872 10920
rect 1912 10888 1944 10920
rect 1984 10888 2016 10920
rect 2056 10888 2088 10920
rect 2128 10888 2160 10920
rect 2200 10888 2232 10920
rect 2272 10888 2304 10920
rect 2344 10888 2376 10920
rect 2416 10888 2448 10920
rect 2488 10888 2520 10920
rect 2560 10888 2592 10920
rect 2632 10888 2664 10920
rect 2704 10888 2736 10920
rect 2776 10888 2808 10920
rect 2848 10888 2880 10920
rect 2920 10888 2952 10920
rect 2992 10888 3024 10920
rect 3064 10888 3096 10920
rect 3136 10888 3168 10920
rect 3208 10888 3240 10920
rect 3280 10888 3312 10920
rect 3352 10888 3384 10920
rect 3424 10888 3456 10920
rect 3496 10888 3528 10920
rect 3568 10888 3600 10920
rect 3640 10888 3672 10920
rect 3712 10888 3744 10920
rect 3784 10888 3816 10920
rect 3856 10888 3888 10920
rect 3928 10888 3960 10920
rect 40 10816 72 10848
rect 112 10816 144 10848
rect 184 10816 216 10848
rect 256 10816 288 10848
rect 328 10816 360 10848
rect 400 10816 432 10848
rect 472 10816 504 10848
rect 544 10816 576 10848
rect 616 10816 648 10848
rect 688 10816 720 10848
rect 760 10816 792 10848
rect 832 10816 864 10848
rect 904 10816 936 10848
rect 976 10816 1008 10848
rect 1048 10816 1080 10848
rect 1120 10816 1152 10848
rect 1192 10816 1224 10848
rect 1264 10816 1296 10848
rect 1336 10816 1368 10848
rect 1408 10816 1440 10848
rect 1480 10816 1512 10848
rect 1552 10816 1584 10848
rect 1624 10816 1656 10848
rect 1696 10816 1728 10848
rect 1768 10816 1800 10848
rect 1840 10816 1872 10848
rect 1912 10816 1944 10848
rect 1984 10816 2016 10848
rect 2056 10816 2088 10848
rect 2128 10816 2160 10848
rect 2200 10816 2232 10848
rect 2272 10816 2304 10848
rect 2344 10816 2376 10848
rect 2416 10816 2448 10848
rect 2488 10816 2520 10848
rect 2560 10816 2592 10848
rect 2632 10816 2664 10848
rect 2704 10816 2736 10848
rect 2776 10816 2808 10848
rect 2848 10816 2880 10848
rect 2920 10816 2952 10848
rect 2992 10816 3024 10848
rect 3064 10816 3096 10848
rect 3136 10816 3168 10848
rect 3208 10816 3240 10848
rect 3280 10816 3312 10848
rect 3352 10816 3384 10848
rect 3424 10816 3456 10848
rect 3496 10816 3528 10848
rect 3568 10816 3600 10848
rect 3640 10816 3672 10848
rect 3712 10816 3744 10848
rect 3784 10816 3816 10848
rect 3856 10816 3888 10848
rect 3928 10816 3960 10848
rect 40 10744 72 10776
rect 112 10744 144 10776
rect 184 10744 216 10776
rect 256 10744 288 10776
rect 328 10744 360 10776
rect 400 10744 432 10776
rect 472 10744 504 10776
rect 544 10744 576 10776
rect 616 10744 648 10776
rect 688 10744 720 10776
rect 760 10744 792 10776
rect 832 10744 864 10776
rect 904 10744 936 10776
rect 976 10744 1008 10776
rect 1048 10744 1080 10776
rect 1120 10744 1152 10776
rect 1192 10744 1224 10776
rect 1264 10744 1296 10776
rect 1336 10744 1368 10776
rect 1408 10744 1440 10776
rect 1480 10744 1512 10776
rect 1552 10744 1584 10776
rect 1624 10744 1656 10776
rect 1696 10744 1728 10776
rect 1768 10744 1800 10776
rect 1840 10744 1872 10776
rect 1912 10744 1944 10776
rect 1984 10744 2016 10776
rect 2056 10744 2088 10776
rect 2128 10744 2160 10776
rect 2200 10744 2232 10776
rect 2272 10744 2304 10776
rect 2344 10744 2376 10776
rect 2416 10744 2448 10776
rect 2488 10744 2520 10776
rect 2560 10744 2592 10776
rect 2632 10744 2664 10776
rect 2704 10744 2736 10776
rect 2776 10744 2808 10776
rect 2848 10744 2880 10776
rect 2920 10744 2952 10776
rect 2992 10744 3024 10776
rect 3064 10744 3096 10776
rect 3136 10744 3168 10776
rect 3208 10744 3240 10776
rect 3280 10744 3312 10776
rect 3352 10744 3384 10776
rect 3424 10744 3456 10776
rect 3496 10744 3528 10776
rect 3568 10744 3600 10776
rect 3640 10744 3672 10776
rect 3712 10744 3744 10776
rect 3784 10744 3816 10776
rect 3856 10744 3888 10776
rect 3928 10744 3960 10776
rect 40 10672 72 10704
rect 112 10672 144 10704
rect 184 10672 216 10704
rect 256 10672 288 10704
rect 328 10672 360 10704
rect 400 10672 432 10704
rect 472 10672 504 10704
rect 544 10672 576 10704
rect 616 10672 648 10704
rect 688 10672 720 10704
rect 760 10672 792 10704
rect 832 10672 864 10704
rect 904 10672 936 10704
rect 976 10672 1008 10704
rect 1048 10672 1080 10704
rect 1120 10672 1152 10704
rect 1192 10672 1224 10704
rect 1264 10672 1296 10704
rect 1336 10672 1368 10704
rect 1408 10672 1440 10704
rect 1480 10672 1512 10704
rect 1552 10672 1584 10704
rect 1624 10672 1656 10704
rect 1696 10672 1728 10704
rect 1768 10672 1800 10704
rect 1840 10672 1872 10704
rect 1912 10672 1944 10704
rect 1984 10672 2016 10704
rect 2056 10672 2088 10704
rect 2128 10672 2160 10704
rect 2200 10672 2232 10704
rect 2272 10672 2304 10704
rect 2344 10672 2376 10704
rect 2416 10672 2448 10704
rect 2488 10672 2520 10704
rect 2560 10672 2592 10704
rect 2632 10672 2664 10704
rect 2704 10672 2736 10704
rect 2776 10672 2808 10704
rect 2848 10672 2880 10704
rect 2920 10672 2952 10704
rect 2992 10672 3024 10704
rect 3064 10672 3096 10704
rect 3136 10672 3168 10704
rect 3208 10672 3240 10704
rect 3280 10672 3312 10704
rect 3352 10672 3384 10704
rect 3424 10672 3456 10704
rect 3496 10672 3528 10704
rect 3568 10672 3600 10704
rect 3640 10672 3672 10704
rect 3712 10672 3744 10704
rect 3784 10672 3816 10704
rect 3856 10672 3888 10704
rect 3928 10672 3960 10704
rect 40 10600 72 10632
rect 112 10600 144 10632
rect 184 10600 216 10632
rect 256 10600 288 10632
rect 328 10600 360 10632
rect 400 10600 432 10632
rect 472 10600 504 10632
rect 544 10600 576 10632
rect 616 10600 648 10632
rect 688 10600 720 10632
rect 760 10600 792 10632
rect 832 10600 864 10632
rect 904 10600 936 10632
rect 976 10600 1008 10632
rect 1048 10600 1080 10632
rect 1120 10600 1152 10632
rect 1192 10600 1224 10632
rect 1264 10600 1296 10632
rect 1336 10600 1368 10632
rect 1408 10600 1440 10632
rect 1480 10600 1512 10632
rect 1552 10600 1584 10632
rect 1624 10600 1656 10632
rect 1696 10600 1728 10632
rect 1768 10600 1800 10632
rect 1840 10600 1872 10632
rect 1912 10600 1944 10632
rect 1984 10600 2016 10632
rect 2056 10600 2088 10632
rect 2128 10600 2160 10632
rect 2200 10600 2232 10632
rect 2272 10600 2304 10632
rect 2344 10600 2376 10632
rect 2416 10600 2448 10632
rect 2488 10600 2520 10632
rect 2560 10600 2592 10632
rect 2632 10600 2664 10632
rect 2704 10600 2736 10632
rect 2776 10600 2808 10632
rect 2848 10600 2880 10632
rect 2920 10600 2952 10632
rect 2992 10600 3024 10632
rect 3064 10600 3096 10632
rect 3136 10600 3168 10632
rect 3208 10600 3240 10632
rect 3280 10600 3312 10632
rect 3352 10600 3384 10632
rect 3424 10600 3456 10632
rect 3496 10600 3528 10632
rect 3568 10600 3600 10632
rect 3640 10600 3672 10632
rect 3712 10600 3744 10632
rect 3784 10600 3816 10632
rect 3856 10600 3888 10632
rect 3928 10600 3960 10632
rect 40 10528 72 10560
rect 112 10528 144 10560
rect 184 10528 216 10560
rect 256 10528 288 10560
rect 328 10528 360 10560
rect 400 10528 432 10560
rect 472 10528 504 10560
rect 544 10528 576 10560
rect 616 10528 648 10560
rect 688 10528 720 10560
rect 760 10528 792 10560
rect 832 10528 864 10560
rect 904 10528 936 10560
rect 976 10528 1008 10560
rect 1048 10528 1080 10560
rect 1120 10528 1152 10560
rect 1192 10528 1224 10560
rect 1264 10528 1296 10560
rect 1336 10528 1368 10560
rect 1408 10528 1440 10560
rect 1480 10528 1512 10560
rect 1552 10528 1584 10560
rect 1624 10528 1656 10560
rect 1696 10528 1728 10560
rect 1768 10528 1800 10560
rect 1840 10528 1872 10560
rect 1912 10528 1944 10560
rect 1984 10528 2016 10560
rect 2056 10528 2088 10560
rect 2128 10528 2160 10560
rect 2200 10528 2232 10560
rect 2272 10528 2304 10560
rect 2344 10528 2376 10560
rect 2416 10528 2448 10560
rect 2488 10528 2520 10560
rect 2560 10528 2592 10560
rect 2632 10528 2664 10560
rect 2704 10528 2736 10560
rect 2776 10528 2808 10560
rect 2848 10528 2880 10560
rect 2920 10528 2952 10560
rect 2992 10528 3024 10560
rect 3064 10528 3096 10560
rect 3136 10528 3168 10560
rect 3208 10528 3240 10560
rect 3280 10528 3312 10560
rect 3352 10528 3384 10560
rect 3424 10528 3456 10560
rect 3496 10528 3528 10560
rect 3568 10528 3600 10560
rect 3640 10528 3672 10560
rect 3712 10528 3744 10560
rect 3784 10528 3816 10560
rect 3856 10528 3888 10560
rect 3928 10528 3960 10560
rect 40 10456 72 10488
rect 112 10456 144 10488
rect 184 10456 216 10488
rect 256 10456 288 10488
rect 328 10456 360 10488
rect 400 10456 432 10488
rect 472 10456 504 10488
rect 544 10456 576 10488
rect 616 10456 648 10488
rect 688 10456 720 10488
rect 760 10456 792 10488
rect 832 10456 864 10488
rect 904 10456 936 10488
rect 976 10456 1008 10488
rect 1048 10456 1080 10488
rect 1120 10456 1152 10488
rect 1192 10456 1224 10488
rect 1264 10456 1296 10488
rect 1336 10456 1368 10488
rect 1408 10456 1440 10488
rect 1480 10456 1512 10488
rect 1552 10456 1584 10488
rect 1624 10456 1656 10488
rect 1696 10456 1728 10488
rect 1768 10456 1800 10488
rect 1840 10456 1872 10488
rect 1912 10456 1944 10488
rect 1984 10456 2016 10488
rect 2056 10456 2088 10488
rect 2128 10456 2160 10488
rect 2200 10456 2232 10488
rect 2272 10456 2304 10488
rect 2344 10456 2376 10488
rect 2416 10456 2448 10488
rect 2488 10456 2520 10488
rect 2560 10456 2592 10488
rect 2632 10456 2664 10488
rect 2704 10456 2736 10488
rect 2776 10456 2808 10488
rect 2848 10456 2880 10488
rect 2920 10456 2952 10488
rect 2992 10456 3024 10488
rect 3064 10456 3096 10488
rect 3136 10456 3168 10488
rect 3208 10456 3240 10488
rect 3280 10456 3312 10488
rect 3352 10456 3384 10488
rect 3424 10456 3456 10488
rect 3496 10456 3528 10488
rect 3568 10456 3600 10488
rect 3640 10456 3672 10488
rect 3712 10456 3744 10488
rect 3784 10456 3816 10488
rect 3856 10456 3888 10488
rect 3928 10456 3960 10488
rect 40 10384 72 10416
rect 112 10384 144 10416
rect 184 10384 216 10416
rect 256 10384 288 10416
rect 328 10384 360 10416
rect 400 10384 432 10416
rect 472 10384 504 10416
rect 544 10384 576 10416
rect 616 10384 648 10416
rect 688 10384 720 10416
rect 760 10384 792 10416
rect 832 10384 864 10416
rect 904 10384 936 10416
rect 976 10384 1008 10416
rect 1048 10384 1080 10416
rect 1120 10384 1152 10416
rect 1192 10384 1224 10416
rect 1264 10384 1296 10416
rect 1336 10384 1368 10416
rect 1408 10384 1440 10416
rect 1480 10384 1512 10416
rect 1552 10384 1584 10416
rect 1624 10384 1656 10416
rect 1696 10384 1728 10416
rect 1768 10384 1800 10416
rect 1840 10384 1872 10416
rect 1912 10384 1944 10416
rect 1984 10384 2016 10416
rect 2056 10384 2088 10416
rect 2128 10384 2160 10416
rect 2200 10384 2232 10416
rect 2272 10384 2304 10416
rect 2344 10384 2376 10416
rect 2416 10384 2448 10416
rect 2488 10384 2520 10416
rect 2560 10384 2592 10416
rect 2632 10384 2664 10416
rect 2704 10384 2736 10416
rect 2776 10384 2808 10416
rect 2848 10384 2880 10416
rect 2920 10384 2952 10416
rect 2992 10384 3024 10416
rect 3064 10384 3096 10416
rect 3136 10384 3168 10416
rect 3208 10384 3240 10416
rect 3280 10384 3312 10416
rect 3352 10384 3384 10416
rect 3424 10384 3456 10416
rect 3496 10384 3528 10416
rect 3568 10384 3600 10416
rect 3640 10384 3672 10416
rect 3712 10384 3744 10416
rect 3784 10384 3816 10416
rect 3856 10384 3888 10416
rect 3928 10384 3960 10416
rect 40 10312 72 10344
rect 112 10312 144 10344
rect 184 10312 216 10344
rect 256 10312 288 10344
rect 328 10312 360 10344
rect 400 10312 432 10344
rect 472 10312 504 10344
rect 544 10312 576 10344
rect 616 10312 648 10344
rect 688 10312 720 10344
rect 760 10312 792 10344
rect 832 10312 864 10344
rect 904 10312 936 10344
rect 976 10312 1008 10344
rect 1048 10312 1080 10344
rect 1120 10312 1152 10344
rect 1192 10312 1224 10344
rect 1264 10312 1296 10344
rect 1336 10312 1368 10344
rect 1408 10312 1440 10344
rect 1480 10312 1512 10344
rect 1552 10312 1584 10344
rect 1624 10312 1656 10344
rect 1696 10312 1728 10344
rect 1768 10312 1800 10344
rect 1840 10312 1872 10344
rect 1912 10312 1944 10344
rect 1984 10312 2016 10344
rect 2056 10312 2088 10344
rect 2128 10312 2160 10344
rect 2200 10312 2232 10344
rect 2272 10312 2304 10344
rect 2344 10312 2376 10344
rect 2416 10312 2448 10344
rect 2488 10312 2520 10344
rect 2560 10312 2592 10344
rect 2632 10312 2664 10344
rect 2704 10312 2736 10344
rect 2776 10312 2808 10344
rect 2848 10312 2880 10344
rect 2920 10312 2952 10344
rect 2992 10312 3024 10344
rect 3064 10312 3096 10344
rect 3136 10312 3168 10344
rect 3208 10312 3240 10344
rect 3280 10312 3312 10344
rect 3352 10312 3384 10344
rect 3424 10312 3456 10344
rect 3496 10312 3528 10344
rect 3568 10312 3600 10344
rect 3640 10312 3672 10344
rect 3712 10312 3744 10344
rect 3784 10312 3816 10344
rect 3856 10312 3888 10344
rect 3928 10312 3960 10344
rect 40 10240 72 10272
rect 112 10240 144 10272
rect 184 10240 216 10272
rect 256 10240 288 10272
rect 328 10240 360 10272
rect 400 10240 432 10272
rect 472 10240 504 10272
rect 544 10240 576 10272
rect 616 10240 648 10272
rect 688 10240 720 10272
rect 760 10240 792 10272
rect 832 10240 864 10272
rect 904 10240 936 10272
rect 976 10240 1008 10272
rect 1048 10240 1080 10272
rect 1120 10240 1152 10272
rect 1192 10240 1224 10272
rect 1264 10240 1296 10272
rect 1336 10240 1368 10272
rect 1408 10240 1440 10272
rect 1480 10240 1512 10272
rect 1552 10240 1584 10272
rect 1624 10240 1656 10272
rect 1696 10240 1728 10272
rect 1768 10240 1800 10272
rect 1840 10240 1872 10272
rect 1912 10240 1944 10272
rect 1984 10240 2016 10272
rect 2056 10240 2088 10272
rect 2128 10240 2160 10272
rect 2200 10240 2232 10272
rect 2272 10240 2304 10272
rect 2344 10240 2376 10272
rect 2416 10240 2448 10272
rect 2488 10240 2520 10272
rect 2560 10240 2592 10272
rect 2632 10240 2664 10272
rect 2704 10240 2736 10272
rect 2776 10240 2808 10272
rect 2848 10240 2880 10272
rect 2920 10240 2952 10272
rect 2992 10240 3024 10272
rect 3064 10240 3096 10272
rect 3136 10240 3168 10272
rect 3208 10240 3240 10272
rect 3280 10240 3312 10272
rect 3352 10240 3384 10272
rect 3424 10240 3456 10272
rect 3496 10240 3528 10272
rect 3568 10240 3600 10272
rect 3640 10240 3672 10272
rect 3712 10240 3744 10272
rect 3784 10240 3816 10272
rect 3856 10240 3888 10272
rect 3928 10240 3960 10272
rect 40 10168 72 10200
rect 112 10168 144 10200
rect 184 10168 216 10200
rect 256 10168 288 10200
rect 328 10168 360 10200
rect 400 10168 432 10200
rect 472 10168 504 10200
rect 544 10168 576 10200
rect 616 10168 648 10200
rect 688 10168 720 10200
rect 760 10168 792 10200
rect 832 10168 864 10200
rect 904 10168 936 10200
rect 976 10168 1008 10200
rect 1048 10168 1080 10200
rect 1120 10168 1152 10200
rect 1192 10168 1224 10200
rect 1264 10168 1296 10200
rect 1336 10168 1368 10200
rect 1408 10168 1440 10200
rect 1480 10168 1512 10200
rect 1552 10168 1584 10200
rect 1624 10168 1656 10200
rect 1696 10168 1728 10200
rect 1768 10168 1800 10200
rect 1840 10168 1872 10200
rect 1912 10168 1944 10200
rect 1984 10168 2016 10200
rect 2056 10168 2088 10200
rect 2128 10168 2160 10200
rect 2200 10168 2232 10200
rect 2272 10168 2304 10200
rect 2344 10168 2376 10200
rect 2416 10168 2448 10200
rect 2488 10168 2520 10200
rect 2560 10168 2592 10200
rect 2632 10168 2664 10200
rect 2704 10168 2736 10200
rect 2776 10168 2808 10200
rect 2848 10168 2880 10200
rect 2920 10168 2952 10200
rect 2992 10168 3024 10200
rect 3064 10168 3096 10200
rect 3136 10168 3168 10200
rect 3208 10168 3240 10200
rect 3280 10168 3312 10200
rect 3352 10168 3384 10200
rect 3424 10168 3456 10200
rect 3496 10168 3528 10200
rect 3568 10168 3600 10200
rect 3640 10168 3672 10200
rect 3712 10168 3744 10200
rect 3784 10168 3816 10200
rect 3856 10168 3888 10200
rect 3928 10168 3960 10200
rect 40 10096 72 10128
rect 112 10096 144 10128
rect 184 10096 216 10128
rect 256 10096 288 10128
rect 328 10096 360 10128
rect 400 10096 432 10128
rect 472 10096 504 10128
rect 544 10096 576 10128
rect 616 10096 648 10128
rect 688 10096 720 10128
rect 760 10096 792 10128
rect 832 10096 864 10128
rect 904 10096 936 10128
rect 976 10096 1008 10128
rect 1048 10096 1080 10128
rect 1120 10096 1152 10128
rect 1192 10096 1224 10128
rect 1264 10096 1296 10128
rect 1336 10096 1368 10128
rect 1408 10096 1440 10128
rect 1480 10096 1512 10128
rect 1552 10096 1584 10128
rect 1624 10096 1656 10128
rect 1696 10096 1728 10128
rect 1768 10096 1800 10128
rect 1840 10096 1872 10128
rect 1912 10096 1944 10128
rect 1984 10096 2016 10128
rect 2056 10096 2088 10128
rect 2128 10096 2160 10128
rect 2200 10096 2232 10128
rect 2272 10096 2304 10128
rect 2344 10096 2376 10128
rect 2416 10096 2448 10128
rect 2488 10096 2520 10128
rect 2560 10096 2592 10128
rect 2632 10096 2664 10128
rect 2704 10096 2736 10128
rect 2776 10096 2808 10128
rect 2848 10096 2880 10128
rect 2920 10096 2952 10128
rect 2992 10096 3024 10128
rect 3064 10096 3096 10128
rect 3136 10096 3168 10128
rect 3208 10096 3240 10128
rect 3280 10096 3312 10128
rect 3352 10096 3384 10128
rect 3424 10096 3456 10128
rect 3496 10096 3528 10128
rect 3568 10096 3600 10128
rect 3640 10096 3672 10128
rect 3712 10096 3744 10128
rect 3784 10096 3816 10128
rect 3856 10096 3888 10128
rect 3928 10096 3960 10128
rect 40 10024 72 10056
rect 112 10024 144 10056
rect 184 10024 216 10056
rect 256 10024 288 10056
rect 328 10024 360 10056
rect 400 10024 432 10056
rect 472 10024 504 10056
rect 544 10024 576 10056
rect 616 10024 648 10056
rect 688 10024 720 10056
rect 760 10024 792 10056
rect 832 10024 864 10056
rect 904 10024 936 10056
rect 976 10024 1008 10056
rect 1048 10024 1080 10056
rect 1120 10024 1152 10056
rect 1192 10024 1224 10056
rect 1264 10024 1296 10056
rect 1336 10024 1368 10056
rect 1408 10024 1440 10056
rect 1480 10024 1512 10056
rect 1552 10024 1584 10056
rect 1624 10024 1656 10056
rect 1696 10024 1728 10056
rect 1768 10024 1800 10056
rect 1840 10024 1872 10056
rect 1912 10024 1944 10056
rect 1984 10024 2016 10056
rect 2056 10024 2088 10056
rect 2128 10024 2160 10056
rect 2200 10024 2232 10056
rect 2272 10024 2304 10056
rect 2344 10024 2376 10056
rect 2416 10024 2448 10056
rect 2488 10024 2520 10056
rect 2560 10024 2592 10056
rect 2632 10024 2664 10056
rect 2704 10024 2736 10056
rect 2776 10024 2808 10056
rect 2848 10024 2880 10056
rect 2920 10024 2952 10056
rect 2992 10024 3024 10056
rect 3064 10024 3096 10056
rect 3136 10024 3168 10056
rect 3208 10024 3240 10056
rect 3280 10024 3312 10056
rect 3352 10024 3384 10056
rect 3424 10024 3456 10056
rect 3496 10024 3528 10056
rect 3568 10024 3600 10056
rect 3640 10024 3672 10056
rect 3712 10024 3744 10056
rect 3784 10024 3816 10056
rect 3856 10024 3888 10056
rect 3928 10024 3960 10056
rect 40 9952 72 9984
rect 112 9952 144 9984
rect 184 9952 216 9984
rect 256 9952 288 9984
rect 328 9952 360 9984
rect 400 9952 432 9984
rect 472 9952 504 9984
rect 544 9952 576 9984
rect 616 9952 648 9984
rect 688 9952 720 9984
rect 760 9952 792 9984
rect 832 9952 864 9984
rect 904 9952 936 9984
rect 976 9952 1008 9984
rect 1048 9952 1080 9984
rect 1120 9952 1152 9984
rect 1192 9952 1224 9984
rect 1264 9952 1296 9984
rect 1336 9952 1368 9984
rect 1408 9952 1440 9984
rect 1480 9952 1512 9984
rect 1552 9952 1584 9984
rect 1624 9952 1656 9984
rect 1696 9952 1728 9984
rect 1768 9952 1800 9984
rect 1840 9952 1872 9984
rect 1912 9952 1944 9984
rect 1984 9952 2016 9984
rect 2056 9952 2088 9984
rect 2128 9952 2160 9984
rect 2200 9952 2232 9984
rect 2272 9952 2304 9984
rect 2344 9952 2376 9984
rect 2416 9952 2448 9984
rect 2488 9952 2520 9984
rect 2560 9952 2592 9984
rect 2632 9952 2664 9984
rect 2704 9952 2736 9984
rect 2776 9952 2808 9984
rect 2848 9952 2880 9984
rect 2920 9952 2952 9984
rect 2992 9952 3024 9984
rect 3064 9952 3096 9984
rect 3136 9952 3168 9984
rect 3208 9952 3240 9984
rect 3280 9952 3312 9984
rect 3352 9952 3384 9984
rect 3424 9952 3456 9984
rect 3496 9952 3528 9984
rect 3568 9952 3600 9984
rect 3640 9952 3672 9984
rect 3712 9952 3744 9984
rect 3784 9952 3816 9984
rect 3856 9952 3888 9984
rect 3928 9952 3960 9984
rect 40 9880 72 9912
rect 112 9880 144 9912
rect 184 9880 216 9912
rect 256 9880 288 9912
rect 328 9880 360 9912
rect 400 9880 432 9912
rect 472 9880 504 9912
rect 544 9880 576 9912
rect 616 9880 648 9912
rect 688 9880 720 9912
rect 760 9880 792 9912
rect 832 9880 864 9912
rect 904 9880 936 9912
rect 976 9880 1008 9912
rect 1048 9880 1080 9912
rect 1120 9880 1152 9912
rect 1192 9880 1224 9912
rect 1264 9880 1296 9912
rect 1336 9880 1368 9912
rect 1408 9880 1440 9912
rect 1480 9880 1512 9912
rect 1552 9880 1584 9912
rect 1624 9880 1656 9912
rect 1696 9880 1728 9912
rect 1768 9880 1800 9912
rect 1840 9880 1872 9912
rect 1912 9880 1944 9912
rect 1984 9880 2016 9912
rect 2056 9880 2088 9912
rect 2128 9880 2160 9912
rect 2200 9880 2232 9912
rect 2272 9880 2304 9912
rect 2344 9880 2376 9912
rect 2416 9880 2448 9912
rect 2488 9880 2520 9912
rect 2560 9880 2592 9912
rect 2632 9880 2664 9912
rect 2704 9880 2736 9912
rect 2776 9880 2808 9912
rect 2848 9880 2880 9912
rect 2920 9880 2952 9912
rect 2992 9880 3024 9912
rect 3064 9880 3096 9912
rect 3136 9880 3168 9912
rect 3208 9880 3240 9912
rect 3280 9880 3312 9912
rect 3352 9880 3384 9912
rect 3424 9880 3456 9912
rect 3496 9880 3528 9912
rect 3568 9880 3600 9912
rect 3640 9880 3672 9912
rect 3712 9880 3744 9912
rect 3784 9880 3816 9912
rect 3856 9880 3888 9912
rect 3928 9880 3960 9912
rect 40 9808 72 9840
rect 112 9808 144 9840
rect 184 9808 216 9840
rect 256 9808 288 9840
rect 328 9808 360 9840
rect 400 9808 432 9840
rect 472 9808 504 9840
rect 544 9808 576 9840
rect 616 9808 648 9840
rect 688 9808 720 9840
rect 760 9808 792 9840
rect 832 9808 864 9840
rect 904 9808 936 9840
rect 976 9808 1008 9840
rect 1048 9808 1080 9840
rect 1120 9808 1152 9840
rect 1192 9808 1224 9840
rect 1264 9808 1296 9840
rect 1336 9808 1368 9840
rect 1408 9808 1440 9840
rect 1480 9808 1512 9840
rect 1552 9808 1584 9840
rect 1624 9808 1656 9840
rect 1696 9808 1728 9840
rect 1768 9808 1800 9840
rect 1840 9808 1872 9840
rect 1912 9808 1944 9840
rect 1984 9808 2016 9840
rect 2056 9808 2088 9840
rect 2128 9808 2160 9840
rect 2200 9808 2232 9840
rect 2272 9808 2304 9840
rect 2344 9808 2376 9840
rect 2416 9808 2448 9840
rect 2488 9808 2520 9840
rect 2560 9808 2592 9840
rect 2632 9808 2664 9840
rect 2704 9808 2736 9840
rect 2776 9808 2808 9840
rect 2848 9808 2880 9840
rect 2920 9808 2952 9840
rect 2992 9808 3024 9840
rect 3064 9808 3096 9840
rect 3136 9808 3168 9840
rect 3208 9808 3240 9840
rect 3280 9808 3312 9840
rect 3352 9808 3384 9840
rect 3424 9808 3456 9840
rect 3496 9808 3528 9840
rect 3568 9808 3600 9840
rect 3640 9808 3672 9840
rect 3712 9808 3744 9840
rect 3784 9808 3816 9840
rect 3856 9808 3888 9840
rect 3928 9808 3960 9840
rect 40 9736 72 9768
rect 112 9736 144 9768
rect 184 9736 216 9768
rect 256 9736 288 9768
rect 328 9736 360 9768
rect 400 9736 432 9768
rect 472 9736 504 9768
rect 544 9736 576 9768
rect 616 9736 648 9768
rect 688 9736 720 9768
rect 760 9736 792 9768
rect 832 9736 864 9768
rect 904 9736 936 9768
rect 976 9736 1008 9768
rect 1048 9736 1080 9768
rect 1120 9736 1152 9768
rect 1192 9736 1224 9768
rect 1264 9736 1296 9768
rect 1336 9736 1368 9768
rect 1408 9736 1440 9768
rect 1480 9736 1512 9768
rect 1552 9736 1584 9768
rect 1624 9736 1656 9768
rect 1696 9736 1728 9768
rect 1768 9736 1800 9768
rect 1840 9736 1872 9768
rect 1912 9736 1944 9768
rect 1984 9736 2016 9768
rect 2056 9736 2088 9768
rect 2128 9736 2160 9768
rect 2200 9736 2232 9768
rect 2272 9736 2304 9768
rect 2344 9736 2376 9768
rect 2416 9736 2448 9768
rect 2488 9736 2520 9768
rect 2560 9736 2592 9768
rect 2632 9736 2664 9768
rect 2704 9736 2736 9768
rect 2776 9736 2808 9768
rect 2848 9736 2880 9768
rect 2920 9736 2952 9768
rect 2992 9736 3024 9768
rect 3064 9736 3096 9768
rect 3136 9736 3168 9768
rect 3208 9736 3240 9768
rect 3280 9736 3312 9768
rect 3352 9736 3384 9768
rect 3424 9736 3456 9768
rect 3496 9736 3528 9768
rect 3568 9736 3600 9768
rect 3640 9736 3672 9768
rect 3712 9736 3744 9768
rect 3784 9736 3816 9768
rect 3856 9736 3888 9768
rect 3928 9736 3960 9768
rect 40 9664 72 9696
rect 112 9664 144 9696
rect 184 9664 216 9696
rect 256 9664 288 9696
rect 328 9664 360 9696
rect 400 9664 432 9696
rect 472 9664 504 9696
rect 544 9664 576 9696
rect 616 9664 648 9696
rect 688 9664 720 9696
rect 760 9664 792 9696
rect 832 9664 864 9696
rect 904 9664 936 9696
rect 976 9664 1008 9696
rect 1048 9664 1080 9696
rect 1120 9664 1152 9696
rect 1192 9664 1224 9696
rect 1264 9664 1296 9696
rect 1336 9664 1368 9696
rect 1408 9664 1440 9696
rect 1480 9664 1512 9696
rect 1552 9664 1584 9696
rect 1624 9664 1656 9696
rect 1696 9664 1728 9696
rect 1768 9664 1800 9696
rect 1840 9664 1872 9696
rect 1912 9664 1944 9696
rect 1984 9664 2016 9696
rect 2056 9664 2088 9696
rect 2128 9664 2160 9696
rect 2200 9664 2232 9696
rect 2272 9664 2304 9696
rect 2344 9664 2376 9696
rect 2416 9664 2448 9696
rect 2488 9664 2520 9696
rect 2560 9664 2592 9696
rect 2632 9664 2664 9696
rect 2704 9664 2736 9696
rect 2776 9664 2808 9696
rect 2848 9664 2880 9696
rect 2920 9664 2952 9696
rect 2992 9664 3024 9696
rect 3064 9664 3096 9696
rect 3136 9664 3168 9696
rect 3208 9664 3240 9696
rect 3280 9664 3312 9696
rect 3352 9664 3384 9696
rect 3424 9664 3456 9696
rect 3496 9664 3528 9696
rect 3568 9664 3600 9696
rect 3640 9664 3672 9696
rect 3712 9664 3744 9696
rect 3784 9664 3816 9696
rect 3856 9664 3888 9696
rect 3928 9664 3960 9696
rect 40 9592 72 9624
rect 112 9592 144 9624
rect 184 9592 216 9624
rect 256 9592 288 9624
rect 328 9592 360 9624
rect 400 9592 432 9624
rect 472 9592 504 9624
rect 544 9592 576 9624
rect 616 9592 648 9624
rect 688 9592 720 9624
rect 760 9592 792 9624
rect 832 9592 864 9624
rect 904 9592 936 9624
rect 976 9592 1008 9624
rect 1048 9592 1080 9624
rect 1120 9592 1152 9624
rect 1192 9592 1224 9624
rect 1264 9592 1296 9624
rect 1336 9592 1368 9624
rect 1408 9592 1440 9624
rect 1480 9592 1512 9624
rect 1552 9592 1584 9624
rect 1624 9592 1656 9624
rect 1696 9592 1728 9624
rect 1768 9592 1800 9624
rect 1840 9592 1872 9624
rect 1912 9592 1944 9624
rect 1984 9592 2016 9624
rect 2056 9592 2088 9624
rect 2128 9592 2160 9624
rect 2200 9592 2232 9624
rect 2272 9592 2304 9624
rect 2344 9592 2376 9624
rect 2416 9592 2448 9624
rect 2488 9592 2520 9624
rect 2560 9592 2592 9624
rect 2632 9592 2664 9624
rect 2704 9592 2736 9624
rect 2776 9592 2808 9624
rect 2848 9592 2880 9624
rect 2920 9592 2952 9624
rect 2992 9592 3024 9624
rect 3064 9592 3096 9624
rect 3136 9592 3168 9624
rect 3208 9592 3240 9624
rect 3280 9592 3312 9624
rect 3352 9592 3384 9624
rect 3424 9592 3456 9624
rect 3496 9592 3528 9624
rect 3568 9592 3600 9624
rect 3640 9592 3672 9624
rect 3712 9592 3744 9624
rect 3784 9592 3816 9624
rect 3856 9592 3888 9624
rect 3928 9592 3960 9624
rect 40 9520 72 9552
rect 112 9520 144 9552
rect 184 9520 216 9552
rect 256 9520 288 9552
rect 328 9520 360 9552
rect 400 9520 432 9552
rect 472 9520 504 9552
rect 544 9520 576 9552
rect 616 9520 648 9552
rect 688 9520 720 9552
rect 760 9520 792 9552
rect 832 9520 864 9552
rect 904 9520 936 9552
rect 976 9520 1008 9552
rect 1048 9520 1080 9552
rect 1120 9520 1152 9552
rect 1192 9520 1224 9552
rect 1264 9520 1296 9552
rect 1336 9520 1368 9552
rect 1408 9520 1440 9552
rect 1480 9520 1512 9552
rect 1552 9520 1584 9552
rect 1624 9520 1656 9552
rect 1696 9520 1728 9552
rect 1768 9520 1800 9552
rect 1840 9520 1872 9552
rect 1912 9520 1944 9552
rect 1984 9520 2016 9552
rect 2056 9520 2088 9552
rect 2128 9520 2160 9552
rect 2200 9520 2232 9552
rect 2272 9520 2304 9552
rect 2344 9520 2376 9552
rect 2416 9520 2448 9552
rect 2488 9520 2520 9552
rect 2560 9520 2592 9552
rect 2632 9520 2664 9552
rect 2704 9520 2736 9552
rect 2776 9520 2808 9552
rect 2848 9520 2880 9552
rect 2920 9520 2952 9552
rect 2992 9520 3024 9552
rect 3064 9520 3096 9552
rect 3136 9520 3168 9552
rect 3208 9520 3240 9552
rect 3280 9520 3312 9552
rect 3352 9520 3384 9552
rect 3424 9520 3456 9552
rect 3496 9520 3528 9552
rect 3568 9520 3600 9552
rect 3640 9520 3672 9552
rect 3712 9520 3744 9552
rect 3784 9520 3816 9552
rect 3856 9520 3888 9552
rect 3928 9520 3960 9552
rect 40 9448 72 9480
rect 112 9448 144 9480
rect 184 9448 216 9480
rect 256 9448 288 9480
rect 328 9448 360 9480
rect 400 9448 432 9480
rect 472 9448 504 9480
rect 544 9448 576 9480
rect 616 9448 648 9480
rect 688 9448 720 9480
rect 760 9448 792 9480
rect 832 9448 864 9480
rect 904 9448 936 9480
rect 976 9448 1008 9480
rect 1048 9448 1080 9480
rect 1120 9448 1152 9480
rect 1192 9448 1224 9480
rect 1264 9448 1296 9480
rect 1336 9448 1368 9480
rect 1408 9448 1440 9480
rect 1480 9448 1512 9480
rect 1552 9448 1584 9480
rect 1624 9448 1656 9480
rect 1696 9448 1728 9480
rect 1768 9448 1800 9480
rect 1840 9448 1872 9480
rect 1912 9448 1944 9480
rect 1984 9448 2016 9480
rect 2056 9448 2088 9480
rect 2128 9448 2160 9480
rect 2200 9448 2232 9480
rect 2272 9448 2304 9480
rect 2344 9448 2376 9480
rect 2416 9448 2448 9480
rect 2488 9448 2520 9480
rect 2560 9448 2592 9480
rect 2632 9448 2664 9480
rect 2704 9448 2736 9480
rect 2776 9448 2808 9480
rect 2848 9448 2880 9480
rect 2920 9448 2952 9480
rect 2992 9448 3024 9480
rect 3064 9448 3096 9480
rect 3136 9448 3168 9480
rect 3208 9448 3240 9480
rect 3280 9448 3312 9480
rect 3352 9448 3384 9480
rect 3424 9448 3456 9480
rect 3496 9448 3528 9480
rect 3568 9448 3600 9480
rect 3640 9448 3672 9480
rect 3712 9448 3744 9480
rect 3784 9448 3816 9480
rect 3856 9448 3888 9480
rect 3928 9448 3960 9480
rect 40 9376 72 9408
rect 112 9376 144 9408
rect 184 9376 216 9408
rect 256 9376 288 9408
rect 328 9376 360 9408
rect 400 9376 432 9408
rect 472 9376 504 9408
rect 544 9376 576 9408
rect 616 9376 648 9408
rect 688 9376 720 9408
rect 760 9376 792 9408
rect 832 9376 864 9408
rect 904 9376 936 9408
rect 976 9376 1008 9408
rect 1048 9376 1080 9408
rect 1120 9376 1152 9408
rect 1192 9376 1224 9408
rect 1264 9376 1296 9408
rect 1336 9376 1368 9408
rect 1408 9376 1440 9408
rect 1480 9376 1512 9408
rect 1552 9376 1584 9408
rect 1624 9376 1656 9408
rect 1696 9376 1728 9408
rect 1768 9376 1800 9408
rect 1840 9376 1872 9408
rect 1912 9376 1944 9408
rect 1984 9376 2016 9408
rect 2056 9376 2088 9408
rect 2128 9376 2160 9408
rect 2200 9376 2232 9408
rect 2272 9376 2304 9408
rect 2344 9376 2376 9408
rect 2416 9376 2448 9408
rect 2488 9376 2520 9408
rect 2560 9376 2592 9408
rect 2632 9376 2664 9408
rect 2704 9376 2736 9408
rect 2776 9376 2808 9408
rect 2848 9376 2880 9408
rect 2920 9376 2952 9408
rect 2992 9376 3024 9408
rect 3064 9376 3096 9408
rect 3136 9376 3168 9408
rect 3208 9376 3240 9408
rect 3280 9376 3312 9408
rect 3352 9376 3384 9408
rect 3424 9376 3456 9408
rect 3496 9376 3528 9408
rect 3568 9376 3600 9408
rect 3640 9376 3672 9408
rect 3712 9376 3744 9408
rect 3784 9376 3816 9408
rect 3856 9376 3888 9408
rect 3928 9376 3960 9408
rect 40 9304 72 9336
rect 112 9304 144 9336
rect 184 9304 216 9336
rect 256 9304 288 9336
rect 328 9304 360 9336
rect 400 9304 432 9336
rect 472 9304 504 9336
rect 544 9304 576 9336
rect 616 9304 648 9336
rect 688 9304 720 9336
rect 760 9304 792 9336
rect 832 9304 864 9336
rect 904 9304 936 9336
rect 976 9304 1008 9336
rect 1048 9304 1080 9336
rect 1120 9304 1152 9336
rect 1192 9304 1224 9336
rect 1264 9304 1296 9336
rect 1336 9304 1368 9336
rect 1408 9304 1440 9336
rect 1480 9304 1512 9336
rect 1552 9304 1584 9336
rect 1624 9304 1656 9336
rect 1696 9304 1728 9336
rect 1768 9304 1800 9336
rect 1840 9304 1872 9336
rect 1912 9304 1944 9336
rect 1984 9304 2016 9336
rect 2056 9304 2088 9336
rect 2128 9304 2160 9336
rect 2200 9304 2232 9336
rect 2272 9304 2304 9336
rect 2344 9304 2376 9336
rect 2416 9304 2448 9336
rect 2488 9304 2520 9336
rect 2560 9304 2592 9336
rect 2632 9304 2664 9336
rect 2704 9304 2736 9336
rect 2776 9304 2808 9336
rect 2848 9304 2880 9336
rect 2920 9304 2952 9336
rect 2992 9304 3024 9336
rect 3064 9304 3096 9336
rect 3136 9304 3168 9336
rect 3208 9304 3240 9336
rect 3280 9304 3312 9336
rect 3352 9304 3384 9336
rect 3424 9304 3456 9336
rect 3496 9304 3528 9336
rect 3568 9304 3600 9336
rect 3640 9304 3672 9336
rect 3712 9304 3744 9336
rect 3784 9304 3816 9336
rect 3856 9304 3888 9336
rect 3928 9304 3960 9336
rect 40 9232 72 9264
rect 112 9232 144 9264
rect 184 9232 216 9264
rect 256 9232 288 9264
rect 328 9232 360 9264
rect 400 9232 432 9264
rect 472 9232 504 9264
rect 544 9232 576 9264
rect 616 9232 648 9264
rect 688 9232 720 9264
rect 760 9232 792 9264
rect 832 9232 864 9264
rect 904 9232 936 9264
rect 976 9232 1008 9264
rect 1048 9232 1080 9264
rect 1120 9232 1152 9264
rect 1192 9232 1224 9264
rect 1264 9232 1296 9264
rect 1336 9232 1368 9264
rect 1408 9232 1440 9264
rect 1480 9232 1512 9264
rect 1552 9232 1584 9264
rect 1624 9232 1656 9264
rect 1696 9232 1728 9264
rect 1768 9232 1800 9264
rect 1840 9232 1872 9264
rect 1912 9232 1944 9264
rect 1984 9232 2016 9264
rect 2056 9232 2088 9264
rect 2128 9232 2160 9264
rect 2200 9232 2232 9264
rect 2272 9232 2304 9264
rect 2344 9232 2376 9264
rect 2416 9232 2448 9264
rect 2488 9232 2520 9264
rect 2560 9232 2592 9264
rect 2632 9232 2664 9264
rect 2704 9232 2736 9264
rect 2776 9232 2808 9264
rect 2848 9232 2880 9264
rect 2920 9232 2952 9264
rect 2992 9232 3024 9264
rect 3064 9232 3096 9264
rect 3136 9232 3168 9264
rect 3208 9232 3240 9264
rect 3280 9232 3312 9264
rect 3352 9232 3384 9264
rect 3424 9232 3456 9264
rect 3496 9232 3528 9264
rect 3568 9232 3600 9264
rect 3640 9232 3672 9264
rect 3712 9232 3744 9264
rect 3784 9232 3816 9264
rect 3856 9232 3888 9264
rect 3928 9232 3960 9264
rect 40 9160 72 9192
rect 112 9160 144 9192
rect 184 9160 216 9192
rect 256 9160 288 9192
rect 328 9160 360 9192
rect 400 9160 432 9192
rect 472 9160 504 9192
rect 544 9160 576 9192
rect 616 9160 648 9192
rect 688 9160 720 9192
rect 760 9160 792 9192
rect 832 9160 864 9192
rect 904 9160 936 9192
rect 976 9160 1008 9192
rect 1048 9160 1080 9192
rect 1120 9160 1152 9192
rect 1192 9160 1224 9192
rect 1264 9160 1296 9192
rect 1336 9160 1368 9192
rect 1408 9160 1440 9192
rect 1480 9160 1512 9192
rect 1552 9160 1584 9192
rect 1624 9160 1656 9192
rect 1696 9160 1728 9192
rect 1768 9160 1800 9192
rect 1840 9160 1872 9192
rect 1912 9160 1944 9192
rect 1984 9160 2016 9192
rect 2056 9160 2088 9192
rect 2128 9160 2160 9192
rect 2200 9160 2232 9192
rect 2272 9160 2304 9192
rect 2344 9160 2376 9192
rect 2416 9160 2448 9192
rect 2488 9160 2520 9192
rect 2560 9160 2592 9192
rect 2632 9160 2664 9192
rect 2704 9160 2736 9192
rect 2776 9160 2808 9192
rect 2848 9160 2880 9192
rect 2920 9160 2952 9192
rect 2992 9160 3024 9192
rect 3064 9160 3096 9192
rect 3136 9160 3168 9192
rect 3208 9160 3240 9192
rect 3280 9160 3312 9192
rect 3352 9160 3384 9192
rect 3424 9160 3456 9192
rect 3496 9160 3528 9192
rect 3568 9160 3600 9192
rect 3640 9160 3672 9192
rect 3712 9160 3744 9192
rect 3784 9160 3816 9192
rect 3856 9160 3888 9192
rect 3928 9160 3960 9192
rect 40 9088 72 9120
rect 112 9088 144 9120
rect 184 9088 216 9120
rect 256 9088 288 9120
rect 328 9088 360 9120
rect 400 9088 432 9120
rect 472 9088 504 9120
rect 544 9088 576 9120
rect 616 9088 648 9120
rect 688 9088 720 9120
rect 760 9088 792 9120
rect 832 9088 864 9120
rect 904 9088 936 9120
rect 976 9088 1008 9120
rect 1048 9088 1080 9120
rect 1120 9088 1152 9120
rect 1192 9088 1224 9120
rect 1264 9088 1296 9120
rect 1336 9088 1368 9120
rect 1408 9088 1440 9120
rect 1480 9088 1512 9120
rect 1552 9088 1584 9120
rect 1624 9088 1656 9120
rect 1696 9088 1728 9120
rect 1768 9088 1800 9120
rect 1840 9088 1872 9120
rect 1912 9088 1944 9120
rect 1984 9088 2016 9120
rect 2056 9088 2088 9120
rect 2128 9088 2160 9120
rect 2200 9088 2232 9120
rect 2272 9088 2304 9120
rect 2344 9088 2376 9120
rect 2416 9088 2448 9120
rect 2488 9088 2520 9120
rect 2560 9088 2592 9120
rect 2632 9088 2664 9120
rect 2704 9088 2736 9120
rect 2776 9088 2808 9120
rect 2848 9088 2880 9120
rect 2920 9088 2952 9120
rect 2992 9088 3024 9120
rect 3064 9088 3096 9120
rect 3136 9088 3168 9120
rect 3208 9088 3240 9120
rect 3280 9088 3312 9120
rect 3352 9088 3384 9120
rect 3424 9088 3456 9120
rect 3496 9088 3528 9120
rect 3568 9088 3600 9120
rect 3640 9088 3672 9120
rect 3712 9088 3744 9120
rect 3784 9088 3816 9120
rect 3856 9088 3888 9120
rect 3928 9088 3960 9120
rect 40 9016 72 9048
rect 112 9016 144 9048
rect 184 9016 216 9048
rect 256 9016 288 9048
rect 328 9016 360 9048
rect 400 9016 432 9048
rect 472 9016 504 9048
rect 544 9016 576 9048
rect 616 9016 648 9048
rect 688 9016 720 9048
rect 760 9016 792 9048
rect 832 9016 864 9048
rect 904 9016 936 9048
rect 976 9016 1008 9048
rect 1048 9016 1080 9048
rect 1120 9016 1152 9048
rect 1192 9016 1224 9048
rect 1264 9016 1296 9048
rect 1336 9016 1368 9048
rect 1408 9016 1440 9048
rect 1480 9016 1512 9048
rect 1552 9016 1584 9048
rect 1624 9016 1656 9048
rect 1696 9016 1728 9048
rect 1768 9016 1800 9048
rect 1840 9016 1872 9048
rect 1912 9016 1944 9048
rect 1984 9016 2016 9048
rect 2056 9016 2088 9048
rect 2128 9016 2160 9048
rect 2200 9016 2232 9048
rect 2272 9016 2304 9048
rect 2344 9016 2376 9048
rect 2416 9016 2448 9048
rect 2488 9016 2520 9048
rect 2560 9016 2592 9048
rect 2632 9016 2664 9048
rect 2704 9016 2736 9048
rect 2776 9016 2808 9048
rect 2848 9016 2880 9048
rect 2920 9016 2952 9048
rect 2992 9016 3024 9048
rect 3064 9016 3096 9048
rect 3136 9016 3168 9048
rect 3208 9016 3240 9048
rect 3280 9016 3312 9048
rect 3352 9016 3384 9048
rect 3424 9016 3456 9048
rect 3496 9016 3528 9048
rect 3568 9016 3600 9048
rect 3640 9016 3672 9048
rect 3712 9016 3744 9048
rect 3784 9016 3816 9048
rect 3856 9016 3888 9048
rect 3928 9016 3960 9048
rect 40 8944 72 8976
rect 112 8944 144 8976
rect 184 8944 216 8976
rect 256 8944 288 8976
rect 328 8944 360 8976
rect 400 8944 432 8976
rect 472 8944 504 8976
rect 544 8944 576 8976
rect 616 8944 648 8976
rect 688 8944 720 8976
rect 760 8944 792 8976
rect 832 8944 864 8976
rect 904 8944 936 8976
rect 976 8944 1008 8976
rect 1048 8944 1080 8976
rect 1120 8944 1152 8976
rect 1192 8944 1224 8976
rect 1264 8944 1296 8976
rect 1336 8944 1368 8976
rect 1408 8944 1440 8976
rect 1480 8944 1512 8976
rect 1552 8944 1584 8976
rect 1624 8944 1656 8976
rect 1696 8944 1728 8976
rect 1768 8944 1800 8976
rect 1840 8944 1872 8976
rect 1912 8944 1944 8976
rect 1984 8944 2016 8976
rect 2056 8944 2088 8976
rect 2128 8944 2160 8976
rect 2200 8944 2232 8976
rect 2272 8944 2304 8976
rect 2344 8944 2376 8976
rect 2416 8944 2448 8976
rect 2488 8944 2520 8976
rect 2560 8944 2592 8976
rect 2632 8944 2664 8976
rect 2704 8944 2736 8976
rect 2776 8944 2808 8976
rect 2848 8944 2880 8976
rect 2920 8944 2952 8976
rect 2992 8944 3024 8976
rect 3064 8944 3096 8976
rect 3136 8944 3168 8976
rect 3208 8944 3240 8976
rect 3280 8944 3312 8976
rect 3352 8944 3384 8976
rect 3424 8944 3456 8976
rect 3496 8944 3528 8976
rect 3568 8944 3600 8976
rect 3640 8944 3672 8976
rect 3712 8944 3744 8976
rect 3784 8944 3816 8976
rect 3856 8944 3888 8976
rect 3928 8944 3960 8976
rect 40 8872 72 8904
rect 112 8872 144 8904
rect 184 8872 216 8904
rect 256 8872 288 8904
rect 328 8872 360 8904
rect 400 8872 432 8904
rect 472 8872 504 8904
rect 544 8872 576 8904
rect 616 8872 648 8904
rect 688 8872 720 8904
rect 760 8872 792 8904
rect 832 8872 864 8904
rect 904 8872 936 8904
rect 976 8872 1008 8904
rect 1048 8872 1080 8904
rect 1120 8872 1152 8904
rect 1192 8872 1224 8904
rect 1264 8872 1296 8904
rect 1336 8872 1368 8904
rect 1408 8872 1440 8904
rect 1480 8872 1512 8904
rect 1552 8872 1584 8904
rect 1624 8872 1656 8904
rect 1696 8872 1728 8904
rect 1768 8872 1800 8904
rect 1840 8872 1872 8904
rect 1912 8872 1944 8904
rect 1984 8872 2016 8904
rect 2056 8872 2088 8904
rect 2128 8872 2160 8904
rect 2200 8872 2232 8904
rect 2272 8872 2304 8904
rect 2344 8872 2376 8904
rect 2416 8872 2448 8904
rect 2488 8872 2520 8904
rect 2560 8872 2592 8904
rect 2632 8872 2664 8904
rect 2704 8872 2736 8904
rect 2776 8872 2808 8904
rect 2848 8872 2880 8904
rect 2920 8872 2952 8904
rect 2992 8872 3024 8904
rect 3064 8872 3096 8904
rect 3136 8872 3168 8904
rect 3208 8872 3240 8904
rect 3280 8872 3312 8904
rect 3352 8872 3384 8904
rect 3424 8872 3456 8904
rect 3496 8872 3528 8904
rect 3568 8872 3600 8904
rect 3640 8872 3672 8904
rect 3712 8872 3744 8904
rect 3784 8872 3816 8904
rect 3856 8872 3888 8904
rect 3928 8872 3960 8904
rect 40 8800 72 8832
rect 112 8800 144 8832
rect 184 8800 216 8832
rect 256 8800 288 8832
rect 328 8800 360 8832
rect 400 8800 432 8832
rect 472 8800 504 8832
rect 544 8800 576 8832
rect 616 8800 648 8832
rect 688 8800 720 8832
rect 760 8800 792 8832
rect 832 8800 864 8832
rect 904 8800 936 8832
rect 976 8800 1008 8832
rect 1048 8800 1080 8832
rect 1120 8800 1152 8832
rect 1192 8800 1224 8832
rect 1264 8800 1296 8832
rect 1336 8800 1368 8832
rect 1408 8800 1440 8832
rect 1480 8800 1512 8832
rect 1552 8800 1584 8832
rect 1624 8800 1656 8832
rect 1696 8800 1728 8832
rect 1768 8800 1800 8832
rect 1840 8800 1872 8832
rect 1912 8800 1944 8832
rect 1984 8800 2016 8832
rect 2056 8800 2088 8832
rect 2128 8800 2160 8832
rect 2200 8800 2232 8832
rect 2272 8800 2304 8832
rect 2344 8800 2376 8832
rect 2416 8800 2448 8832
rect 2488 8800 2520 8832
rect 2560 8800 2592 8832
rect 2632 8800 2664 8832
rect 2704 8800 2736 8832
rect 2776 8800 2808 8832
rect 2848 8800 2880 8832
rect 2920 8800 2952 8832
rect 2992 8800 3024 8832
rect 3064 8800 3096 8832
rect 3136 8800 3168 8832
rect 3208 8800 3240 8832
rect 3280 8800 3312 8832
rect 3352 8800 3384 8832
rect 3424 8800 3456 8832
rect 3496 8800 3528 8832
rect 3568 8800 3600 8832
rect 3640 8800 3672 8832
rect 3712 8800 3744 8832
rect 3784 8800 3816 8832
rect 3856 8800 3888 8832
rect 3928 8800 3960 8832
rect 40 8728 72 8760
rect 112 8728 144 8760
rect 184 8728 216 8760
rect 256 8728 288 8760
rect 328 8728 360 8760
rect 400 8728 432 8760
rect 472 8728 504 8760
rect 544 8728 576 8760
rect 616 8728 648 8760
rect 688 8728 720 8760
rect 760 8728 792 8760
rect 832 8728 864 8760
rect 904 8728 936 8760
rect 976 8728 1008 8760
rect 1048 8728 1080 8760
rect 1120 8728 1152 8760
rect 1192 8728 1224 8760
rect 1264 8728 1296 8760
rect 1336 8728 1368 8760
rect 1408 8728 1440 8760
rect 1480 8728 1512 8760
rect 1552 8728 1584 8760
rect 1624 8728 1656 8760
rect 1696 8728 1728 8760
rect 1768 8728 1800 8760
rect 1840 8728 1872 8760
rect 1912 8728 1944 8760
rect 1984 8728 2016 8760
rect 2056 8728 2088 8760
rect 2128 8728 2160 8760
rect 2200 8728 2232 8760
rect 2272 8728 2304 8760
rect 2344 8728 2376 8760
rect 2416 8728 2448 8760
rect 2488 8728 2520 8760
rect 2560 8728 2592 8760
rect 2632 8728 2664 8760
rect 2704 8728 2736 8760
rect 2776 8728 2808 8760
rect 2848 8728 2880 8760
rect 2920 8728 2952 8760
rect 2992 8728 3024 8760
rect 3064 8728 3096 8760
rect 3136 8728 3168 8760
rect 3208 8728 3240 8760
rect 3280 8728 3312 8760
rect 3352 8728 3384 8760
rect 3424 8728 3456 8760
rect 3496 8728 3528 8760
rect 3568 8728 3600 8760
rect 3640 8728 3672 8760
rect 3712 8728 3744 8760
rect 3784 8728 3816 8760
rect 3856 8728 3888 8760
rect 3928 8728 3960 8760
rect 40 8656 72 8688
rect 112 8656 144 8688
rect 184 8656 216 8688
rect 256 8656 288 8688
rect 328 8656 360 8688
rect 400 8656 432 8688
rect 472 8656 504 8688
rect 544 8656 576 8688
rect 616 8656 648 8688
rect 688 8656 720 8688
rect 760 8656 792 8688
rect 832 8656 864 8688
rect 904 8656 936 8688
rect 976 8656 1008 8688
rect 1048 8656 1080 8688
rect 1120 8656 1152 8688
rect 1192 8656 1224 8688
rect 1264 8656 1296 8688
rect 1336 8656 1368 8688
rect 1408 8656 1440 8688
rect 1480 8656 1512 8688
rect 1552 8656 1584 8688
rect 1624 8656 1656 8688
rect 1696 8656 1728 8688
rect 1768 8656 1800 8688
rect 1840 8656 1872 8688
rect 1912 8656 1944 8688
rect 1984 8656 2016 8688
rect 2056 8656 2088 8688
rect 2128 8656 2160 8688
rect 2200 8656 2232 8688
rect 2272 8656 2304 8688
rect 2344 8656 2376 8688
rect 2416 8656 2448 8688
rect 2488 8656 2520 8688
rect 2560 8656 2592 8688
rect 2632 8656 2664 8688
rect 2704 8656 2736 8688
rect 2776 8656 2808 8688
rect 2848 8656 2880 8688
rect 2920 8656 2952 8688
rect 2992 8656 3024 8688
rect 3064 8656 3096 8688
rect 3136 8656 3168 8688
rect 3208 8656 3240 8688
rect 3280 8656 3312 8688
rect 3352 8656 3384 8688
rect 3424 8656 3456 8688
rect 3496 8656 3528 8688
rect 3568 8656 3600 8688
rect 3640 8656 3672 8688
rect 3712 8656 3744 8688
rect 3784 8656 3816 8688
rect 3856 8656 3888 8688
rect 3928 8656 3960 8688
rect 40 8584 72 8616
rect 112 8584 144 8616
rect 184 8584 216 8616
rect 256 8584 288 8616
rect 328 8584 360 8616
rect 400 8584 432 8616
rect 472 8584 504 8616
rect 544 8584 576 8616
rect 616 8584 648 8616
rect 688 8584 720 8616
rect 760 8584 792 8616
rect 832 8584 864 8616
rect 904 8584 936 8616
rect 976 8584 1008 8616
rect 1048 8584 1080 8616
rect 1120 8584 1152 8616
rect 1192 8584 1224 8616
rect 1264 8584 1296 8616
rect 1336 8584 1368 8616
rect 1408 8584 1440 8616
rect 1480 8584 1512 8616
rect 1552 8584 1584 8616
rect 1624 8584 1656 8616
rect 1696 8584 1728 8616
rect 1768 8584 1800 8616
rect 1840 8584 1872 8616
rect 1912 8584 1944 8616
rect 1984 8584 2016 8616
rect 2056 8584 2088 8616
rect 2128 8584 2160 8616
rect 2200 8584 2232 8616
rect 2272 8584 2304 8616
rect 2344 8584 2376 8616
rect 2416 8584 2448 8616
rect 2488 8584 2520 8616
rect 2560 8584 2592 8616
rect 2632 8584 2664 8616
rect 2704 8584 2736 8616
rect 2776 8584 2808 8616
rect 2848 8584 2880 8616
rect 2920 8584 2952 8616
rect 2992 8584 3024 8616
rect 3064 8584 3096 8616
rect 3136 8584 3168 8616
rect 3208 8584 3240 8616
rect 3280 8584 3312 8616
rect 3352 8584 3384 8616
rect 3424 8584 3456 8616
rect 3496 8584 3528 8616
rect 3568 8584 3600 8616
rect 3640 8584 3672 8616
rect 3712 8584 3744 8616
rect 3784 8584 3816 8616
rect 3856 8584 3888 8616
rect 3928 8584 3960 8616
rect 40 8512 72 8544
rect 112 8512 144 8544
rect 184 8512 216 8544
rect 256 8512 288 8544
rect 328 8512 360 8544
rect 400 8512 432 8544
rect 472 8512 504 8544
rect 544 8512 576 8544
rect 616 8512 648 8544
rect 688 8512 720 8544
rect 760 8512 792 8544
rect 832 8512 864 8544
rect 904 8512 936 8544
rect 976 8512 1008 8544
rect 1048 8512 1080 8544
rect 1120 8512 1152 8544
rect 1192 8512 1224 8544
rect 1264 8512 1296 8544
rect 1336 8512 1368 8544
rect 1408 8512 1440 8544
rect 1480 8512 1512 8544
rect 1552 8512 1584 8544
rect 1624 8512 1656 8544
rect 1696 8512 1728 8544
rect 1768 8512 1800 8544
rect 1840 8512 1872 8544
rect 1912 8512 1944 8544
rect 1984 8512 2016 8544
rect 2056 8512 2088 8544
rect 2128 8512 2160 8544
rect 2200 8512 2232 8544
rect 2272 8512 2304 8544
rect 2344 8512 2376 8544
rect 2416 8512 2448 8544
rect 2488 8512 2520 8544
rect 2560 8512 2592 8544
rect 2632 8512 2664 8544
rect 2704 8512 2736 8544
rect 2776 8512 2808 8544
rect 2848 8512 2880 8544
rect 2920 8512 2952 8544
rect 2992 8512 3024 8544
rect 3064 8512 3096 8544
rect 3136 8512 3168 8544
rect 3208 8512 3240 8544
rect 3280 8512 3312 8544
rect 3352 8512 3384 8544
rect 3424 8512 3456 8544
rect 3496 8512 3528 8544
rect 3568 8512 3600 8544
rect 3640 8512 3672 8544
rect 3712 8512 3744 8544
rect 3784 8512 3816 8544
rect 3856 8512 3888 8544
rect 3928 8512 3960 8544
rect 40 8440 72 8472
rect 112 8440 144 8472
rect 184 8440 216 8472
rect 256 8440 288 8472
rect 328 8440 360 8472
rect 400 8440 432 8472
rect 472 8440 504 8472
rect 544 8440 576 8472
rect 616 8440 648 8472
rect 688 8440 720 8472
rect 760 8440 792 8472
rect 832 8440 864 8472
rect 904 8440 936 8472
rect 976 8440 1008 8472
rect 1048 8440 1080 8472
rect 1120 8440 1152 8472
rect 1192 8440 1224 8472
rect 1264 8440 1296 8472
rect 1336 8440 1368 8472
rect 1408 8440 1440 8472
rect 1480 8440 1512 8472
rect 1552 8440 1584 8472
rect 1624 8440 1656 8472
rect 1696 8440 1728 8472
rect 1768 8440 1800 8472
rect 1840 8440 1872 8472
rect 1912 8440 1944 8472
rect 1984 8440 2016 8472
rect 2056 8440 2088 8472
rect 2128 8440 2160 8472
rect 2200 8440 2232 8472
rect 2272 8440 2304 8472
rect 2344 8440 2376 8472
rect 2416 8440 2448 8472
rect 2488 8440 2520 8472
rect 2560 8440 2592 8472
rect 2632 8440 2664 8472
rect 2704 8440 2736 8472
rect 2776 8440 2808 8472
rect 2848 8440 2880 8472
rect 2920 8440 2952 8472
rect 2992 8440 3024 8472
rect 3064 8440 3096 8472
rect 3136 8440 3168 8472
rect 3208 8440 3240 8472
rect 3280 8440 3312 8472
rect 3352 8440 3384 8472
rect 3424 8440 3456 8472
rect 3496 8440 3528 8472
rect 3568 8440 3600 8472
rect 3640 8440 3672 8472
rect 3712 8440 3744 8472
rect 3784 8440 3816 8472
rect 3856 8440 3888 8472
rect 3928 8440 3960 8472
rect 40 8368 72 8400
rect 112 8368 144 8400
rect 184 8368 216 8400
rect 256 8368 288 8400
rect 328 8368 360 8400
rect 400 8368 432 8400
rect 472 8368 504 8400
rect 544 8368 576 8400
rect 616 8368 648 8400
rect 688 8368 720 8400
rect 760 8368 792 8400
rect 832 8368 864 8400
rect 904 8368 936 8400
rect 976 8368 1008 8400
rect 1048 8368 1080 8400
rect 1120 8368 1152 8400
rect 1192 8368 1224 8400
rect 1264 8368 1296 8400
rect 1336 8368 1368 8400
rect 1408 8368 1440 8400
rect 1480 8368 1512 8400
rect 1552 8368 1584 8400
rect 1624 8368 1656 8400
rect 1696 8368 1728 8400
rect 1768 8368 1800 8400
rect 1840 8368 1872 8400
rect 1912 8368 1944 8400
rect 1984 8368 2016 8400
rect 2056 8368 2088 8400
rect 2128 8368 2160 8400
rect 2200 8368 2232 8400
rect 2272 8368 2304 8400
rect 2344 8368 2376 8400
rect 2416 8368 2448 8400
rect 2488 8368 2520 8400
rect 2560 8368 2592 8400
rect 2632 8368 2664 8400
rect 2704 8368 2736 8400
rect 2776 8368 2808 8400
rect 2848 8368 2880 8400
rect 2920 8368 2952 8400
rect 2992 8368 3024 8400
rect 3064 8368 3096 8400
rect 3136 8368 3168 8400
rect 3208 8368 3240 8400
rect 3280 8368 3312 8400
rect 3352 8368 3384 8400
rect 3424 8368 3456 8400
rect 3496 8368 3528 8400
rect 3568 8368 3600 8400
rect 3640 8368 3672 8400
rect 3712 8368 3744 8400
rect 3784 8368 3816 8400
rect 3856 8368 3888 8400
rect 3928 8368 3960 8400
rect 40 8296 72 8328
rect 112 8296 144 8328
rect 184 8296 216 8328
rect 256 8296 288 8328
rect 328 8296 360 8328
rect 400 8296 432 8328
rect 472 8296 504 8328
rect 544 8296 576 8328
rect 616 8296 648 8328
rect 688 8296 720 8328
rect 760 8296 792 8328
rect 832 8296 864 8328
rect 904 8296 936 8328
rect 976 8296 1008 8328
rect 1048 8296 1080 8328
rect 1120 8296 1152 8328
rect 1192 8296 1224 8328
rect 1264 8296 1296 8328
rect 1336 8296 1368 8328
rect 1408 8296 1440 8328
rect 1480 8296 1512 8328
rect 1552 8296 1584 8328
rect 1624 8296 1656 8328
rect 1696 8296 1728 8328
rect 1768 8296 1800 8328
rect 1840 8296 1872 8328
rect 1912 8296 1944 8328
rect 1984 8296 2016 8328
rect 2056 8296 2088 8328
rect 2128 8296 2160 8328
rect 2200 8296 2232 8328
rect 2272 8296 2304 8328
rect 2344 8296 2376 8328
rect 2416 8296 2448 8328
rect 2488 8296 2520 8328
rect 2560 8296 2592 8328
rect 2632 8296 2664 8328
rect 2704 8296 2736 8328
rect 2776 8296 2808 8328
rect 2848 8296 2880 8328
rect 2920 8296 2952 8328
rect 2992 8296 3024 8328
rect 3064 8296 3096 8328
rect 3136 8296 3168 8328
rect 3208 8296 3240 8328
rect 3280 8296 3312 8328
rect 3352 8296 3384 8328
rect 3424 8296 3456 8328
rect 3496 8296 3528 8328
rect 3568 8296 3600 8328
rect 3640 8296 3672 8328
rect 3712 8296 3744 8328
rect 3784 8296 3816 8328
rect 3856 8296 3888 8328
rect 3928 8296 3960 8328
rect 40 8224 72 8256
rect 112 8224 144 8256
rect 184 8224 216 8256
rect 256 8224 288 8256
rect 328 8224 360 8256
rect 400 8224 432 8256
rect 472 8224 504 8256
rect 544 8224 576 8256
rect 616 8224 648 8256
rect 688 8224 720 8256
rect 760 8224 792 8256
rect 832 8224 864 8256
rect 904 8224 936 8256
rect 976 8224 1008 8256
rect 1048 8224 1080 8256
rect 1120 8224 1152 8256
rect 1192 8224 1224 8256
rect 1264 8224 1296 8256
rect 1336 8224 1368 8256
rect 1408 8224 1440 8256
rect 1480 8224 1512 8256
rect 1552 8224 1584 8256
rect 1624 8224 1656 8256
rect 1696 8224 1728 8256
rect 1768 8224 1800 8256
rect 1840 8224 1872 8256
rect 1912 8224 1944 8256
rect 1984 8224 2016 8256
rect 2056 8224 2088 8256
rect 2128 8224 2160 8256
rect 2200 8224 2232 8256
rect 2272 8224 2304 8256
rect 2344 8224 2376 8256
rect 2416 8224 2448 8256
rect 2488 8224 2520 8256
rect 2560 8224 2592 8256
rect 2632 8224 2664 8256
rect 2704 8224 2736 8256
rect 2776 8224 2808 8256
rect 2848 8224 2880 8256
rect 2920 8224 2952 8256
rect 2992 8224 3024 8256
rect 3064 8224 3096 8256
rect 3136 8224 3168 8256
rect 3208 8224 3240 8256
rect 3280 8224 3312 8256
rect 3352 8224 3384 8256
rect 3424 8224 3456 8256
rect 3496 8224 3528 8256
rect 3568 8224 3600 8256
rect 3640 8224 3672 8256
rect 3712 8224 3744 8256
rect 3784 8224 3816 8256
rect 3856 8224 3888 8256
rect 3928 8224 3960 8256
rect 40 8152 72 8184
rect 112 8152 144 8184
rect 184 8152 216 8184
rect 256 8152 288 8184
rect 328 8152 360 8184
rect 400 8152 432 8184
rect 472 8152 504 8184
rect 544 8152 576 8184
rect 616 8152 648 8184
rect 688 8152 720 8184
rect 760 8152 792 8184
rect 832 8152 864 8184
rect 904 8152 936 8184
rect 976 8152 1008 8184
rect 1048 8152 1080 8184
rect 1120 8152 1152 8184
rect 1192 8152 1224 8184
rect 1264 8152 1296 8184
rect 1336 8152 1368 8184
rect 1408 8152 1440 8184
rect 1480 8152 1512 8184
rect 1552 8152 1584 8184
rect 1624 8152 1656 8184
rect 1696 8152 1728 8184
rect 1768 8152 1800 8184
rect 1840 8152 1872 8184
rect 1912 8152 1944 8184
rect 1984 8152 2016 8184
rect 2056 8152 2088 8184
rect 2128 8152 2160 8184
rect 2200 8152 2232 8184
rect 2272 8152 2304 8184
rect 2344 8152 2376 8184
rect 2416 8152 2448 8184
rect 2488 8152 2520 8184
rect 2560 8152 2592 8184
rect 2632 8152 2664 8184
rect 2704 8152 2736 8184
rect 2776 8152 2808 8184
rect 2848 8152 2880 8184
rect 2920 8152 2952 8184
rect 2992 8152 3024 8184
rect 3064 8152 3096 8184
rect 3136 8152 3168 8184
rect 3208 8152 3240 8184
rect 3280 8152 3312 8184
rect 3352 8152 3384 8184
rect 3424 8152 3456 8184
rect 3496 8152 3528 8184
rect 3568 8152 3600 8184
rect 3640 8152 3672 8184
rect 3712 8152 3744 8184
rect 3784 8152 3816 8184
rect 3856 8152 3888 8184
rect 3928 8152 3960 8184
rect 40 8080 72 8112
rect 112 8080 144 8112
rect 184 8080 216 8112
rect 256 8080 288 8112
rect 328 8080 360 8112
rect 400 8080 432 8112
rect 472 8080 504 8112
rect 544 8080 576 8112
rect 616 8080 648 8112
rect 688 8080 720 8112
rect 760 8080 792 8112
rect 832 8080 864 8112
rect 904 8080 936 8112
rect 976 8080 1008 8112
rect 1048 8080 1080 8112
rect 1120 8080 1152 8112
rect 1192 8080 1224 8112
rect 1264 8080 1296 8112
rect 1336 8080 1368 8112
rect 1408 8080 1440 8112
rect 1480 8080 1512 8112
rect 1552 8080 1584 8112
rect 1624 8080 1656 8112
rect 1696 8080 1728 8112
rect 1768 8080 1800 8112
rect 1840 8080 1872 8112
rect 1912 8080 1944 8112
rect 1984 8080 2016 8112
rect 2056 8080 2088 8112
rect 2128 8080 2160 8112
rect 2200 8080 2232 8112
rect 2272 8080 2304 8112
rect 2344 8080 2376 8112
rect 2416 8080 2448 8112
rect 2488 8080 2520 8112
rect 2560 8080 2592 8112
rect 2632 8080 2664 8112
rect 2704 8080 2736 8112
rect 2776 8080 2808 8112
rect 2848 8080 2880 8112
rect 2920 8080 2952 8112
rect 2992 8080 3024 8112
rect 3064 8080 3096 8112
rect 3136 8080 3168 8112
rect 3208 8080 3240 8112
rect 3280 8080 3312 8112
rect 3352 8080 3384 8112
rect 3424 8080 3456 8112
rect 3496 8080 3528 8112
rect 3568 8080 3600 8112
rect 3640 8080 3672 8112
rect 3712 8080 3744 8112
rect 3784 8080 3816 8112
rect 3856 8080 3888 8112
rect 3928 8080 3960 8112
rect 40 8008 72 8040
rect 112 8008 144 8040
rect 184 8008 216 8040
rect 256 8008 288 8040
rect 328 8008 360 8040
rect 400 8008 432 8040
rect 472 8008 504 8040
rect 544 8008 576 8040
rect 616 8008 648 8040
rect 688 8008 720 8040
rect 760 8008 792 8040
rect 832 8008 864 8040
rect 904 8008 936 8040
rect 976 8008 1008 8040
rect 1048 8008 1080 8040
rect 1120 8008 1152 8040
rect 1192 8008 1224 8040
rect 1264 8008 1296 8040
rect 1336 8008 1368 8040
rect 1408 8008 1440 8040
rect 1480 8008 1512 8040
rect 1552 8008 1584 8040
rect 1624 8008 1656 8040
rect 1696 8008 1728 8040
rect 1768 8008 1800 8040
rect 1840 8008 1872 8040
rect 1912 8008 1944 8040
rect 1984 8008 2016 8040
rect 2056 8008 2088 8040
rect 2128 8008 2160 8040
rect 2200 8008 2232 8040
rect 2272 8008 2304 8040
rect 2344 8008 2376 8040
rect 2416 8008 2448 8040
rect 2488 8008 2520 8040
rect 2560 8008 2592 8040
rect 2632 8008 2664 8040
rect 2704 8008 2736 8040
rect 2776 8008 2808 8040
rect 2848 8008 2880 8040
rect 2920 8008 2952 8040
rect 2992 8008 3024 8040
rect 3064 8008 3096 8040
rect 3136 8008 3168 8040
rect 3208 8008 3240 8040
rect 3280 8008 3312 8040
rect 3352 8008 3384 8040
rect 3424 8008 3456 8040
rect 3496 8008 3528 8040
rect 3568 8008 3600 8040
rect 3640 8008 3672 8040
rect 3712 8008 3744 8040
rect 3784 8008 3816 8040
rect 3856 8008 3888 8040
rect 3928 8008 3960 8040
rect 40 7936 72 7968
rect 112 7936 144 7968
rect 184 7936 216 7968
rect 256 7936 288 7968
rect 328 7936 360 7968
rect 400 7936 432 7968
rect 472 7936 504 7968
rect 544 7936 576 7968
rect 616 7936 648 7968
rect 688 7936 720 7968
rect 760 7936 792 7968
rect 832 7936 864 7968
rect 904 7936 936 7968
rect 976 7936 1008 7968
rect 1048 7936 1080 7968
rect 1120 7936 1152 7968
rect 1192 7936 1224 7968
rect 1264 7936 1296 7968
rect 1336 7936 1368 7968
rect 1408 7936 1440 7968
rect 1480 7936 1512 7968
rect 1552 7936 1584 7968
rect 1624 7936 1656 7968
rect 1696 7936 1728 7968
rect 1768 7936 1800 7968
rect 1840 7936 1872 7968
rect 1912 7936 1944 7968
rect 1984 7936 2016 7968
rect 2056 7936 2088 7968
rect 2128 7936 2160 7968
rect 2200 7936 2232 7968
rect 2272 7936 2304 7968
rect 2344 7936 2376 7968
rect 2416 7936 2448 7968
rect 2488 7936 2520 7968
rect 2560 7936 2592 7968
rect 2632 7936 2664 7968
rect 2704 7936 2736 7968
rect 2776 7936 2808 7968
rect 2848 7936 2880 7968
rect 2920 7936 2952 7968
rect 2992 7936 3024 7968
rect 3064 7936 3096 7968
rect 3136 7936 3168 7968
rect 3208 7936 3240 7968
rect 3280 7936 3312 7968
rect 3352 7936 3384 7968
rect 3424 7936 3456 7968
rect 3496 7936 3528 7968
rect 3568 7936 3600 7968
rect 3640 7936 3672 7968
rect 3712 7936 3744 7968
rect 3784 7936 3816 7968
rect 3856 7936 3888 7968
rect 3928 7936 3960 7968
rect 40 7864 72 7896
rect 112 7864 144 7896
rect 184 7864 216 7896
rect 256 7864 288 7896
rect 328 7864 360 7896
rect 400 7864 432 7896
rect 472 7864 504 7896
rect 544 7864 576 7896
rect 616 7864 648 7896
rect 688 7864 720 7896
rect 760 7864 792 7896
rect 832 7864 864 7896
rect 904 7864 936 7896
rect 976 7864 1008 7896
rect 1048 7864 1080 7896
rect 1120 7864 1152 7896
rect 1192 7864 1224 7896
rect 1264 7864 1296 7896
rect 1336 7864 1368 7896
rect 1408 7864 1440 7896
rect 1480 7864 1512 7896
rect 1552 7864 1584 7896
rect 1624 7864 1656 7896
rect 1696 7864 1728 7896
rect 1768 7864 1800 7896
rect 1840 7864 1872 7896
rect 1912 7864 1944 7896
rect 1984 7864 2016 7896
rect 2056 7864 2088 7896
rect 2128 7864 2160 7896
rect 2200 7864 2232 7896
rect 2272 7864 2304 7896
rect 2344 7864 2376 7896
rect 2416 7864 2448 7896
rect 2488 7864 2520 7896
rect 2560 7864 2592 7896
rect 2632 7864 2664 7896
rect 2704 7864 2736 7896
rect 2776 7864 2808 7896
rect 2848 7864 2880 7896
rect 2920 7864 2952 7896
rect 2992 7864 3024 7896
rect 3064 7864 3096 7896
rect 3136 7864 3168 7896
rect 3208 7864 3240 7896
rect 3280 7864 3312 7896
rect 3352 7864 3384 7896
rect 3424 7864 3456 7896
rect 3496 7864 3528 7896
rect 3568 7864 3600 7896
rect 3640 7864 3672 7896
rect 3712 7864 3744 7896
rect 3784 7864 3816 7896
rect 3856 7864 3888 7896
rect 3928 7864 3960 7896
rect 40 7792 72 7824
rect 112 7792 144 7824
rect 184 7792 216 7824
rect 256 7792 288 7824
rect 328 7792 360 7824
rect 400 7792 432 7824
rect 472 7792 504 7824
rect 544 7792 576 7824
rect 616 7792 648 7824
rect 688 7792 720 7824
rect 760 7792 792 7824
rect 832 7792 864 7824
rect 904 7792 936 7824
rect 976 7792 1008 7824
rect 1048 7792 1080 7824
rect 1120 7792 1152 7824
rect 1192 7792 1224 7824
rect 1264 7792 1296 7824
rect 1336 7792 1368 7824
rect 1408 7792 1440 7824
rect 1480 7792 1512 7824
rect 1552 7792 1584 7824
rect 1624 7792 1656 7824
rect 1696 7792 1728 7824
rect 1768 7792 1800 7824
rect 1840 7792 1872 7824
rect 1912 7792 1944 7824
rect 1984 7792 2016 7824
rect 2056 7792 2088 7824
rect 2128 7792 2160 7824
rect 2200 7792 2232 7824
rect 2272 7792 2304 7824
rect 2344 7792 2376 7824
rect 2416 7792 2448 7824
rect 2488 7792 2520 7824
rect 2560 7792 2592 7824
rect 2632 7792 2664 7824
rect 2704 7792 2736 7824
rect 2776 7792 2808 7824
rect 2848 7792 2880 7824
rect 2920 7792 2952 7824
rect 2992 7792 3024 7824
rect 3064 7792 3096 7824
rect 3136 7792 3168 7824
rect 3208 7792 3240 7824
rect 3280 7792 3312 7824
rect 3352 7792 3384 7824
rect 3424 7792 3456 7824
rect 3496 7792 3528 7824
rect 3568 7792 3600 7824
rect 3640 7792 3672 7824
rect 3712 7792 3744 7824
rect 3784 7792 3816 7824
rect 3856 7792 3888 7824
rect 3928 7792 3960 7824
rect 40 7720 72 7752
rect 112 7720 144 7752
rect 184 7720 216 7752
rect 256 7720 288 7752
rect 328 7720 360 7752
rect 400 7720 432 7752
rect 472 7720 504 7752
rect 544 7720 576 7752
rect 616 7720 648 7752
rect 688 7720 720 7752
rect 760 7720 792 7752
rect 832 7720 864 7752
rect 904 7720 936 7752
rect 976 7720 1008 7752
rect 1048 7720 1080 7752
rect 1120 7720 1152 7752
rect 1192 7720 1224 7752
rect 1264 7720 1296 7752
rect 1336 7720 1368 7752
rect 1408 7720 1440 7752
rect 1480 7720 1512 7752
rect 1552 7720 1584 7752
rect 1624 7720 1656 7752
rect 1696 7720 1728 7752
rect 1768 7720 1800 7752
rect 1840 7720 1872 7752
rect 1912 7720 1944 7752
rect 1984 7720 2016 7752
rect 2056 7720 2088 7752
rect 2128 7720 2160 7752
rect 2200 7720 2232 7752
rect 2272 7720 2304 7752
rect 2344 7720 2376 7752
rect 2416 7720 2448 7752
rect 2488 7720 2520 7752
rect 2560 7720 2592 7752
rect 2632 7720 2664 7752
rect 2704 7720 2736 7752
rect 2776 7720 2808 7752
rect 2848 7720 2880 7752
rect 2920 7720 2952 7752
rect 2992 7720 3024 7752
rect 3064 7720 3096 7752
rect 3136 7720 3168 7752
rect 3208 7720 3240 7752
rect 3280 7720 3312 7752
rect 3352 7720 3384 7752
rect 3424 7720 3456 7752
rect 3496 7720 3528 7752
rect 3568 7720 3600 7752
rect 3640 7720 3672 7752
rect 3712 7720 3744 7752
rect 3784 7720 3816 7752
rect 3856 7720 3888 7752
rect 3928 7720 3960 7752
rect 40 7648 72 7680
rect 112 7648 144 7680
rect 184 7648 216 7680
rect 256 7648 288 7680
rect 328 7648 360 7680
rect 400 7648 432 7680
rect 472 7648 504 7680
rect 544 7648 576 7680
rect 616 7648 648 7680
rect 688 7648 720 7680
rect 760 7648 792 7680
rect 832 7648 864 7680
rect 904 7648 936 7680
rect 976 7648 1008 7680
rect 1048 7648 1080 7680
rect 1120 7648 1152 7680
rect 1192 7648 1224 7680
rect 1264 7648 1296 7680
rect 1336 7648 1368 7680
rect 1408 7648 1440 7680
rect 1480 7648 1512 7680
rect 1552 7648 1584 7680
rect 1624 7648 1656 7680
rect 1696 7648 1728 7680
rect 1768 7648 1800 7680
rect 1840 7648 1872 7680
rect 1912 7648 1944 7680
rect 1984 7648 2016 7680
rect 2056 7648 2088 7680
rect 2128 7648 2160 7680
rect 2200 7648 2232 7680
rect 2272 7648 2304 7680
rect 2344 7648 2376 7680
rect 2416 7648 2448 7680
rect 2488 7648 2520 7680
rect 2560 7648 2592 7680
rect 2632 7648 2664 7680
rect 2704 7648 2736 7680
rect 2776 7648 2808 7680
rect 2848 7648 2880 7680
rect 2920 7648 2952 7680
rect 2992 7648 3024 7680
rect 3064 7648 3096 7680
rect 3136 7648 3168 7680
rect 3208 7648 3240 7680
rect 3280 7648 3312 7680
rect 3352 7648 3384 7680
rect 3424 7648 3456 7680
rect 3496 7648 3528 7680
rect 3568 7648 3600 7680
rect 3640 7648 3672 7680
rect 3712 7648 3744 7680
rect 3784 7648 3816 7680
rect 3856 7648 3888 7680
rect 3928 7648 3960 7680
rect 40 7576 72 7608
rect 112 7576 144 7608
rect 184 7576 216 7608
rect 256 7576 288 7608
rect 328 7576 360 7608
rect 400 7576 432 7608
rect 472 7576 504 7608
rect 544 7576 576 7608
rect 616 7576 648 7608
rect 688 7576 720 7608
rect 760 7576 792 7608
rect 832 7576 864 7608
rect 904 7576 936 7608
rect 976 7576 1008 7608
rect 1048 7576 1080 7608
rect 1120 7576 1152 7608
rect 1192 7576 1224 7608
rect 1264 7576 1296 7608
rect 1336 7576 1368 7608
rect 1408 7576 1440 7608
rect 1480 7576 1512 7608
rect 1552 7576 1584 7608
rect 1624 7576 1656 7608
rect 1696 7576 1728 7608
rect 1768 7576 1800 7608
rect 1840 7576 1872 7608
rect 1912 7576 1944 7608
rect 1984 7576 2016 7608
rect 2056 7576 2088 7608
rect 2128 7576 2160 7608
rect 2200 7576 2232 7608
rect 2272 7576 2304 7608
rect 2344 7576 2376 7608
rect 2416 7576 2448 7608
rect 2488 7576 2520 7608
rect 2560 7576 2592 7608
rect 2632 7576 2664 7608
rect 2704 7576 2736 7608
rect 2776 7576 2808 7608
rect 2848 7576 2880 7608
rect 2920 7576 2952 7608
rect 2992 7576 3024 7608
rect 3064 7576 3096 7608
rect 3136 7576 3168 7608
rect 3208 7576 3240 7608
rect 3280 7576 3312 7608
rect 3352 7576 3384 7608
rect 3424 7576 3456 7608
rect 3496 7576 3528 7608
rect 3568 7576 3600 7608
rect 3640 7576 3672 7608
rect 3712 7576 3744 7608
rect 3784 7576 3816 7608
rect 3856 7576 3888 7608
rect 3928 7576 3960 7608
rect 40 7504 72 7536
rect 112 7504 144 7536
rect 184 7504 216 7536
rect 256 7504 288 7536
rect 328 7504 360 7536
rect 400 7504 432 7536
rect 472 7504 504 7536
rect 544 7504 576 7536
rect 616 7504 648 7536
rect 688 7504 720 7536
rect 760 7504 792 7536
rect 832 7504 864 7536
rect 904 7504 936 7536
rect 976 7504 1008 7536
rect 1048 7504 1080 7536
rect 1120 7504 1152 7536
rect 1192 7504 1224 7536
rect 1264 7504 1296 7536
rect 1336 7504 1368 7536
rect 1408 7504 1440 7536
rect 1480 7504 1512 7536
rect 1552 7504 1584 7536
rect 1624 7504 1656 7536
rect 1696 7504 1728 7536
rect 1768 7504 1800 7536
rect 1840 7504 1872 7536
rect 1912 7504 1944 7536
rect 1984 7504 2016 7536
rect 2056 7504 2088 7536
rect 2128 7504 2160 7536
rect 2200 7504 2232 7536
rect 2272 7504 2304 7536
rect 2344 7504 2376 7536
rect 2416 7504 2448 7536
rect 2488 7504 2520 7536
rect 2560 7504 2592 7536
rect 2632 7504 2664 7536
rect 2704 7504 2736 7536
rect 2776 7504 2808 7536
rect 2848 7504 2880 7536
rect 2920 7504 2952 7536
rect 2992 7504 3024 7536
rect 3064 7504 3096 7536
rect 3136 7504 3168 7536
rect 3208 7504 3240 7536
rect 3280 7504 3312 7536
rect 3352 7504 3384 7536
rect 3424 7504 3456 7536
rect 3496 7504 3528 7536
rect 3568 7504 3600 7536
rect 3640 7504 3672 7536
rect 3712 7504 3744 7536
rect 3784 7504 3816 7536
rect 3856 7504 3888 7536
rect 3928 7504 3960 7536
rect 40 7432 72 7464
rect 112 7432 144 7464
rect 184 7432 216 7464
rect 256 7432 288 7464
rect 328 7432 360 7464
rect 400 7432 432 7464
rect 472 7432 504 7464
rect 544 7432 576 7464
rect 616 7432 648 7464
rect 688 7432 720 7464
rect 760 7432 792 7464
rect 832 7432 864 7464
rect 904 7432 936 7464
rect 976 7432 1008 7464
rect 1048 7432 1080 7464
rect 1120 7432 1152 7464
rect 1192 7432 1224 7464
rect 1264 7432 1296 7464
rect 1336 7432 1368 7464
rect 1408 7432 1440 7464
rect 1480 7432 1512 7464
rect 1552 7432 1584 7464
rect 1624 7432 1656 7464
rect 1696 7432 1728 7464
rect 1768 7432 1800 7464
rect 1840 7432 1872 7464
rect 1912 7432 1944 7464
rect 1984 7432 2016 7464
rect 2056 7432 2088 7464
rect 2128 7432 2160 7464
rect 2200 7432 2232 7464
rect 2272 7432 2304 7464
rect 2344 7432 2376 7464
rect 2416 7432 2448 7464
rect 2488 7432 2520 7464
rect 2560 7432 2592 7464
rect 2632 7432 2664 7464
rect 2704 7432 2736 7464
rect 2776 7432 2808 7464
rect 2848 7432 2880 7464
rect 2920 7432 2952 7464
rect 2992 7432 3024 7464
rect 3064 7432 3096 7464
rect 3136 7432 3168 7464
rect 3208 7432 3240 7464
rect 3280 7432 3312 7464
rect 3352 7432 3384 7464
rect 3424 7432 3456 7464
rect 3496 7432 3528 7464
rect 3568 7432 3600 7464
rect 3640 7432 3672 7464
rect 3712 7432 3744 7464
rect 3784 7432 3816 7464
rect 3856 7432 3888 7464
rect 3928 7432 3960 7464
rect 40 7360 72 7392
rect 112 7360 144 7392
rect 184 7360 216 7392
rect 256 7360 288 7392
rect 328 7360 360 7392
rect 400 7360 432 7392
rect 472 7360 504 7392
rect 544 7360 576 7392
rect 616 7360 648 7392
rect 688 7360 720 7392
rect 760 7360 792 7392
rect 832 7360 864 7392
rect 904 7360 936 7392
rect 976 7360 1008 7392
rect 1048 7360 1080 7392
rect 1120 7360 1152 7392
rect 1192 7360 1224 7392
rect 1264 7360 1296 7392
rect 1336 7360 1368 7392
rect 1408 7360 1440 7392
rect 1480 7360 1512 7392
rect 1552 7360 1584 7392
rect 1624 7360 1656 7392
rect 1696 7360 1728 7392
rect 1768 7360 1800 7392
rect 1840 7360 1872 7392
rect 1912 7360 1944 7392
rect 1984 7360 2016 7392
rect 2056 7360 2088 7392
rect 2128 7360 2160 7392
rect 2200 7360 2232 7392
rect 2272 7360 2304 7392
rect 2344 7360 2376 7392
rect 2416 7360 2448 7392
rect 2488 7360 2520 7392
rect 2560 7360 2592 7392
rect 2632 7360 2664 7392
rect 2704 7360 2736 7392
rect 2776 7360 2808 7392
rect 2848 7360 2880 7392
rect 2920 7360 2952 7392
rect 2992 7360 3024 7392
rect 3064 7360 3096 7392
rect 3136 7360 3168 7392
rect 3208 7360 3240 7392
rect 3280 7360 3312 7392
rect 3352 7360 3384 7392
rect 3424 7360 3456 7392
rect 3496 7360 3528 7392
rect 3568 7360 3600 7392
rect 3640 7360 3672 7392
rect 3712 7360 3744 7392
rect 3784 7360 3816 7392
rect 3856 7360 3888 7392
rect 3928 7360 3960 7392
rect 40 7288 72 7320
rect 112 7288 144 7320
rect 184 7288 216 7320
rect 256 7288 288 7320
rect 328 7288 360 7320
rect 400 7288 432 7320
rect 472 7288 504 7320
rect 544 7288 576 7320
rect 616 7288 648 7320
rect 688 7288 720 7320
rect 760 7288 792 7320
rect 832 7288 864 7320
rect 904 7288 936 7320
rect 976 7288 1008 7320
rect 1048 7288 1080 7320
rect 1120 7288 1152 7320
rect 1192 7288 1224 7320
rect 1264 7288 1296 7320
rect 1336 7288 1368 7320
rect 1408 7288 1440 7320
rect 1480 7288 1512 7320
rect 1552 7288 1584 7320
rect 1624 7288 1656 7320
rect 1696 7288 1728 7320
rect 1768 7288 1800 7320
rect 1840 7288 1872 7320
rect 1912 7288 1944 7320
rect 1984 7288 2016 7320
rect 2056 7288 2088 7320
rect 2128 7288 2160 7320
rect 2200 7288 2232 7320
rect 2272 7288 2304 7320
rect 2344 7288 2376 7320
rect 2416 7288 2448 7320
rect 2488 7288 2520 7320
rect 2560 7288 2592 7320
rect 2632 7288 2664 7320
rect 2704 7288 2736 7320
rect 2776 7288 2808 7320
rect 2848 7288 2880 7320
rect 2920 7288 2952 7320
rect 2992 7288 3024 7320
rect 3064 7288 3096 7320
rect 3136 7288 3168 7320
rect 3208 7288 3240 7320
rect 3280 7288 3312 7320
rect 3352 7288 3384 7320
rect 3424 7288 3456 7320
rect 3496 7288 3528 7320
rect 3568 7288 3600 7320
rect 3640 7288 3672 7320
rect 3712 7288 3744 7320
rect 3784 7288 3816 7320
rect 3856 7288 3888 7320
rect 3928 7288 3960 7320
rect 40 7216 72 7248
rect 112 7216 144 7248
rect 184 7216 216 7248
rect 256 7216 288 7248
rect 328 7216 360 7248
rect 400 7216 432 7248
rect 472 7216 504 7248
rect 544 7216 576 7248
rect 616 7216 648 7248
rect 688 7216 720 7248
rect 760 7216 792 7248
rect 832 7216 864 7248
rect 904 7216 936 7248
rect 976 7216 1008 7248
rect 1048 7216 1080 7248
rect 1120 7216 1152 7248
rect 1192 7216 1224 7248
rect 1264 7216 1296 7248
rect 1336 7216 1368 7248
rect 1408 7216 1440 7248
rect 1480 7216 1512 7248
rect 1552 7216 1584 7248
rect 1624 7216 1656 7248
rect 1696 7216 1728 7248
rect 1768 7216 1800 7248
rect 1840 7216 1872 7248
rect 1912 7216 1944 7248
rect 1984 7216 2016 7248
rect 2056 7216 2088 7248
rect 2128 7216 2160 7248
rect 2200 7216 2232 7248
rect 2272 7216 2304 7248
rect 2344 7216 2376 7248
rect 2416 7216 2448 7248
rect 2488 7216 2520 7248
rect 2560 7216 2592 7248
rect 2632 7216 2664 7248
rect 2704 7216 2736 7248
rect 2776 7216 2808 7248
rect 2848 7216 2880 7248
rect 2920 7216 2952 7248
rect 2992 7216 3024 7248
rect 3064 7216 3096 7248
rect 3136 7216 3168 7248
rect 3208 7216 3240 7248
rect 3280 7216 3312 7248
rect 3352 7216 3384 7248
rect 3424 7216 3456 7248
rect 3496 7216 3528 7248
rect 3568 7216 3600 7248
rect 3640 7216 3672 7248
rect 3712 7216 3744 7248
rect 3784 7216 3816 7248
rect 3856 7216 3888 7248
rect 3928 7216 3960 7248
rect 40 7144 72 7176
rect 112 7144 144 7176
rect 184 7144 216 7176
rect 256 7144 288 7176
rect 328 7144 360 7176
rect 400 7144 432 7176
rect 472 7144 504 7176
rect 544 7144 576 7176
rect 616 7144 648 7176
rect 688 7144 720 7176
rect 760 7144 792 7176
rect 832 7144 864 7176
rect 904 7144 936 7176
rect 976 7144 1008 7176
rect 1048 7144 1080 7176
rect 1120 7144 1152 7176
rect 1192 7144 1224 7176
rect 1264 7144 1296 7176
rect 1336 7144 1368 7176
rect 1408 7144 1440 7176
rect 1480 7144 1512 7176
rect 1552 7144 1584 7176
rect 1624 7144 1656 7176
rect 1696 7144 1728 7176
rect 1768 7144 1800 7176
rect 1840 7144 1872 7176
rect 1912 7144 1944 7176
rect 1984 7144 2016 7176
rect 2056 7144 2088 7176
rect 2128 7144 2160 7176
rect 2200 7144 2232 7176
rect 2272 7144 2304 7176
rect 2344 7144 2376 7176
rect 2416 7144 2448 7176
rect 2488 7144 2520 7176
rect 2560 7144 2592 7176
rect 2632 7144 2664 7176
rect 2704 7144 2736 7176
rect 2776 7144 2808 7176
rect 2848 7144 2880 7176
rect 2920 7144 2952 7176
rect 2992 7144 3024 7176
rect 3064 7144 3096 7176
rect 3136 7144 3168 7176
rect 3208 7144 3240 7176
rect 3280 7144 3312 7176
rect 3352 7144 3384 7176
rect 3424 7144 3456 7176
rect 3496 7144 3528 7176
rect 3568 7144 3600 7176
rect 3640 7144 3672 7176
rect 3712 7144 3744 7176
rect 3784 7144 3816 7176
rect 3856 7144 3888 7176
rect 3928 7144 3960 7176
rect 40 7072 72 7104
rect 112 7072 144 7104
rect 184 7072 216 7104
rect 256 7072 288 7104
rect 328 7072 360 7104
rect 400 7072 432 7104
rect 472 7072 504 7104
rect 544 7072 576 7104
rect 616 7072 648 7104
rect 688 7072 720 7104
rect 760 7072 792 7104
rect 832 7072 864 7104
rect 904 7072 936 7104
rect 976 7072 1008 7104
rect 1048 7072 1080 7104
rect 1120 7072 1152 7104
rect 1192 7072 1224 7104
rect 1264 7072 1296 7104
rect 1336 7072 1368 7104
rect 1408 7072 1440 7104
rect 1480 7072 1512 7104
rect 1552 7072 1584 7104
rect 1624 7072 1656 7104
rect 1696 7072 1728 7104
rect 1768 7072 1800 7104
rect 1840 7072 1872 7104
rect 1912 7072 1944 7104
rect 1984 7072 2016 7104
rect 2056 7072 2088 7104
rect 2128 7072 2160 7104
rect 2200 7072 2232 7104
rect 2272 7072 2304 7104
rect 2344 7072 2376 7104
rect 2416 7072 2448 7104
rect 2488 7072 2520 7104
rect 2560 7072 2592 7104
rect 2632 7072 2664 7104
rect 2704 7072 2736 7104
rect 2776 7072 2808 7104
rect 2848 7072 2880 7104
rect 2920 7072 2952 7104
rect 2992 7072 3024 7104
rect 3064 7072 3096 7104
rect 3136 7072 3168 7104
rect 3208 7072 3240 7104
rect 3280 7072 3312 7104
rect 3352 7072 3384 7104
rect 3424 7072 3456 7104
rect 3496 7072 3528 7104
rect 3568 7072 3600 7104
rect 3640 7072 3672 7104
rect 3712 7072 3744 7104
rect 3784 7072 3816 7104
rect 3856 7072 3888 7104
rect 3928 7072 3960 7104
rect 40 7000 72 7032
rect 112 7000 144 7032
rect 184 7000 216 7032
rect 256 7000 288 7032
rect 328 7000 360 7032
rect 400 7000 432 7032
rect 472 7000 504 7032
rect 544 7000 576 7032
rect 616 7000 648 7032
rect 688 7000 720 7032
rect 760 7000 792 7032
rect 832 7000 864 7032
rect 904 7000 936 7032
rect 976 7000 1008 7032
rect 1048 7000 1080 7032
rect 1120 7000 1152 7032
rect 1192 7000 1224 7032
rect 1264 7000 1296 7032
rect 1336 7000 1368 7032
rect 1408 7000 1440 7032
rect 1480 7000 1512 7032
rect 1552 7000 1584 7032
rect 1624 7000 1656 7032
rect 1696 7000 1728 7032
rect 1768 7000 1800 7032
rect 1840 7000 1872 7032
rect 1912 7000 1944 7032
rect 1984 7000 2016 7032
rect 2056 7000 2088 7032
rect 2128 7000 2160 7032
rect 2200 7000 2232 7032
rect 2272 7000 2304 7032
rect 2344 7000 2376 7032
rect 2416 7000 2448 7032
rect 2488 7000 2520 7032
rect 2560 7000 2592 7032
rect 2632 7000 2664 7032
rect 2704 7000 2736 7032
rect 2776 7000 2808 7032
rect 2848 7000 2880 7032
rect 2920 7000 2952 7032
rect 2992 7000 3024 7032
rect 3064 7000 3096 7032
rect 3136 7000 3168 7032
rect 3208 7000 3240 7032
rect 3280 7000 3312 7032
rect 3352 7000 3384 7032
rect 3424 7000 3456 7032
rect 3496 7000 3528 7032
rect 3568 7000 3600 7032
rect 3640 7000 3672 7032
rect 3712 7000 3744 7032
rect 3784 7000 3816 7032
rect 3856 7000 3888 7032
rect 3928 7000 3960 7032
rect 40 6928 72 6960
rect 112 6928 144 6960
rect 184 6928 216 6960
rect 256 6928 288 6960
rect 328 6928 360 6960
rect 400 6928 432 6960
rect 472 6928 504 6960
rect 544 6928 576 6960
rect 616 6928 648 6960
rect 688 6928 720 6960
rect 760 6928 792 6960
rect 832 6928 864 6960
rect 904 6928 936 6960
rect 976 6928 1008 6960
rect 1048 6928 1080 6960
rect 1120 6928 1152 6960
rect 1192 6928 1224 6960
rect 1264 6928 1296 6960
rect 1336 6928 1368 6960
rect 1408 6928 1440 6960
rect 1480 6928 1512 6960
rect 1552 6928 1584 6960
rect 1624 6928 1656 6960
rect 1696 6928 1728 6960
rect 1768 6928 1800 6960
rect 1840 6928 1872 6960
rect 1912 6928 1944 6960
rect 1984 6928 2016 6960
rect 2056 6928 2088 6960
rect 2128 6928 2160 6960
rect 2200 6928 2232 6960
rect 2272 6928 2304 6960
rect 2344 6928 2376 6960
rect 2416 6928 2448 6960
rect 2488 6928 2520 6960
rect 2560 6928 2592 6960
rect 2632 6928 2664 6960
rect 2704 6928 2736 6960
rect 2776 6928 2808 6960
rect 2848 6928 2880 6960
rect 2920 6928 2952 6960
rect 2992 6928 3024 6960
rect 3064 6928 3096 6960
rect 3136 6928 3168 6960
rect 3208 6928 3240 6960
rect 3280 6928 3312 6960
rect 3352 6928 3384 6960
rect 3424 6928 3456 6960
rect 3496 6928 3528 6960
rect 3568 6928 3600 6960
rect 3640 6928 3672 6960
rect 3712 6928 3744 6960
rect 3784 6928 3816 6960
rect 3856 6928 3888 6960
rect 3928 6928 3960 6960
rect 40 6856 72 6888
rect 112 6856 144 6888
rect 184 6856 216 6888
rect 256 6856 288 6888
rect 328 6856 360 6888
rect 400 6856 432 6888
rect 472 6856 504 6888
rect 544 6856 576 6888
rect 616 6856 648 6888
rect 688 6856 720 6888
rect 760 6856 792 6888
rect 832 6856 864 6888
rect 904 6856 936 6888
rect 976 6856 1008 6888
rect 1048 6856 1080 6888
rect 1120 6856 1152 6888
rect 1192 6856 1224 6888
rect 1264 6856 1296 6888
rect 1336 6856 1368 6888
rect 1408 6856 1440 6888
rect 1480 6856 1512 6888
rect 1552 6856 1584 6888
rect 1624 6856 1656 6888
rect 1696 6856 1728 6888
rect 1768 6856 1800 6888
rect 1840 6856 1872 6888
rect 1912 6856 1944 6888
rect 1984 6856 2016 6888
rect 2056 6856 2088 6888
rect 2128 6856 2160 6888
rect 2200 6856 2232 6888
rect 2272 6856 2304 6888
rect 2344 6856 2376 6888
rect 2416 6856 2448 6888
rect 2488 6856 2520 6888
rect 2560 6856 2592 6888
rect 2632 6856 2664 6888
rect 2704 6856 2736 6888
rect 2776 6856 2808 6888
rect 2848 6856 2880 6888
rect 2920 6856 2952 6888
rect 2992 6856 3024 6888
rect 3064 6856 3096 6888
rect 3136 6856 3168 6888
rect 3208 6856 3240 6888
rect 3280 6856 3312 6888
rect 3352 6856 3384 6888
rect 3424 6856 3456 6888
rect 3496 6856 3528 6888
rect 3568 6856 3600 6888
rect 3640 6856 3672 6888
rect 3712 6856 3744 6888
rect 3784 6856 3816 6888
rect 3856 6856 3888 6888
rect 3928 6856 3960 6888
rect 112 6512 144 6544
rect 184 6512 216 6544
rect 256 6512 288 6544
rect 328 6512 360 6544
rect 400 6512 432 6544
rect 472 6512 504 6544
rect 544 6512 576 6544
rect 616 6512 648 6544
rect 688 6512 720 6544
rect 760 6512 792 6544
rect 832 6512 864 6544
rect 904 6512 936 6544
rect 976 6512 1008 6544
rect 1048 6512 1080 6544
rect 1120 6512 1152 6544
rect 1192 6512 1224 6544
rect 1264 6512 1296 6544
rect 1336 6512 1368 6544
rect 1408 6512 1440 6544
rect 1480 6512 1512 6544
rect 1552 6512 1584 6544
rect 1624 6512 1656 6544
rect 1696 6512 1728 6544
rect 1768 6512 1800 6544
rect 1840 6512 1872 6544
rect 1912 6512 1944 6544
rect 1984 6512 2016 6544
rect 2056 6512 2088 6544
rect 2128 6512 2160 6544
rect 2200 6512 2232 6544
rect 2272 6512 2304 6544
rect 2344 6512 2376 6544
rect 2416 6512 2448 6544
rect 2488 6512 2520 6544
rect 2560 6512 2592 6544
rect 2632 6512 2664 6544
rect 2704 6512 2736 6544
rect 2776 6512 2808 6544
rect 2848 6512 2880 6544
rect 2920 6512 2952 6544
rect 2992 6512 3024 6544
rect 3064 6512 3096 6544
rect 3136 6512 3168 6544
rect 3208 6512 3240 6544
rect 3280 6512 3312 6544
rect 3352 6512 3384 6544
rect 3424 6512 3456 6544
rect 3496 6512 3528 6544
rect 3568 6512 3600 6544
rect 3640 6512 3672 6544
rect 3712 6512 3744 6544
rect 3784 6512 3816 6544
rect 3856 6512 3888 6544
rect 3928 6512 3960 6544
rect 40 6440 72 6472
rect 112 6440 144 6472
rect 184 6440 216 6472
rect 256 6440 288 6472
rect 328 6440 360 6472
rect 400 6440 432 6472
rect 472 6440 504 6472
rect 544 6440 576 6472
rect 616 6440 648 6472
rect 688 6440 720 6472
rect 760 6440 792 6472
rect 832 6440 864 6472
rect 904 6440 936 6472
rect 976 6440 1008 6472
rect 1048 6440 1080 6472
rect 1120 6440 1152 6472
rect 1192 6440 1224 6472
rect 1264 6440 1296 6472
rect 1336 6440 1368 6472
rect 1408 6440 1440 6472
rect 1480 6440 1512 6472
rect 1552 6440 1584 6472
rect 1624 6440 1656 6472
rect 1696 6440 1728 6472
rect 1768 6440 1800 6472
rect 1840 6440 1872 6472
rect 1912 6440 1944 6472
rect 1984 6440 2016 6472
rect 2056 6440 2088 6472
rect 2128 6440 2160 6472
rect 2200 6440 2232 6472
rect 2272 6440 2304 6472
rect 2344 6440 2376 6472
rect 2416 6440 2448 6472
rect 2488 6440 2520 6472
rect 2560 6440 2592 6472
rect 2632 6440 2664 6472
rect 2704 6440 2736 6472
rect 2776 6440 2808 6472
rect 2848 6440 2880 6472
rect 2920 6440 2952 6472
rect 2992 6440 3024 6472
rect 3064 6440 3096 6472
rect 3136 6440 3168 6472
rect 3208 6440 3240 6472
rect 3280 6440 3312 6472
rect 3352 6440 3384 6472
rect 3424 6440 3456 6472
rect 3496 6440 3528 6472
rect 3568 6440 3600 6472
rect 3640 6440 3672 6472
rect 3712 6440 3744 6472
rect 3784 6440 3816 6472
rect 3856 6440 3888 6472
rect 3928 6440 3960 6472
rect 40 6368 72 6400
rect 112 6368 144 6400
rect 184 6368 216 6400
rect 256 6368 288 6400
rect 328 6368 360 6400
rect 400 6368 432 6400
rect 472 6368 504 6400
rect 544 6368 576 6400
rect 616 6368 648 6400
rect 688 6368 720 6400
rect 760 6368 792 6400
rect 832 6368 864 6400
rect 904 6368 936 6400
rect 976 6368 1008 6400
rect 1048 6368 1080 6400
rect 1120 6368 1152 6400
rect 1192 6368 1224 6400
rect 1264 6368 1296 6400
rect 1336 6368 1368 6400
rect 1408 6368 1440 6400
rect 1480 6368 1512 6400
rect 1552 6368 1584 6400
rect 1624 6368 1656 6400
rect 1696 6368 1728 6400
rect 1768 6368 1800 6400
rect 1840 6368 1872 6400
rect 1912 6368 1944 6400
rect 1984 6368 2016 6400
rect 2056 6368 2088 6400
rect 2128 6368 2160 6400
rect 2200 6368 2232 6400
rect 2272 6368 2304 6400
rect 2344 6368 2376 6400
rect 2416 6368 2448 6400
rect 2488 6368 2520 6400
rect 2560 6368 2592 6400
rect 2632 6368 2664 6400
rect 2704 6368 2736 6400
rect 2776 6368 2808 6400
rect 2848 6368 2880 6400
rect 2920 6368 2952 6400
rect 2992 6368 3024 6400
rect 3064 6368 3096 6400
rect 3136 6368 3168 6400
rect 3208 6368 3240 6400
rect 3280 6368 3312 6400
rect 3352 6368 3384 6400
rect 3424 6368 3456 6400
rect 3496 6368 3528 6400
rect 3568 6368 3600 6400
rect 3640 6368 3672 6400
rect 3712 6368 3744 6400
rect 3784 6368 3816 6400
rect 3856 6368 3888 6400
rect 3928 6368 3960 6400
rect 40 6296 72 6328
rect 112 6296 144 6328
rect 184 6296 216 6328
rect 256 6296 288 6328
rect 328 6296 360 6328
rect 400 6296 432 6328
rect 472 6296 504 6328
rect 544 6296 576 6328
rect 616 6296 648 6328
rect 688 6296 720 6328
rect 760 6296 792 6328
rect 832 6296 864 6328
rect 904 6296 936 6328
rect 976 6296 1008 6328
rect 1048 6296 1080 6328
rect 1120 6296 1152 6328
rect 1192 6296 1224 6328
rect 1264 6296 1296 6328
rect 1336 6296 1368 6328
rect 1408 6296 1440 6328
rect 1480 6296 1512 6328
rect 1552 6296 1584 6328
rect 1624 6296 1656 6328
rect 1696 6296 1728 6328
rect 1768 6296 1800 6328
rect 1840 6296 1872 6328
rect 1912 6296 1944 6328
rect 1984 6296 2016 6328
rect 2056 6296 2088 6328
rect 2128 6296 2160 6328
rect 2200 6296 2232 6328
rect 2272 6296 2304 6328
rect 2344 6296 2376 6328
rect 2416 6296 2448 6328
rect 2488 6296 2520 6328
rect 2560 6296 2592 6328
rect 2632 6296 2664 6328
rect 2704 6296 2736 6328
rect 2776 6296 2808 6328
rect 2848 6296 2880 6328
rect 2920 6296 2952 6328
rect 2992 6296 3024 6328
rect 3064 6296 3096 6328
rect 3136 6296 3168 6328
rect 3208 6296 3240 6328
rect 3280 6296 3312 6328
rect 3352 6296 3384 6328
rect 3424 6296 3456 6328
rect 3496 6296 3528 6328
rect 3568 6296 3600 6328
rect 3640 6296 3672 6328
rect 3712 6296 3744 6328
rect 3784 6296 3816 6328
rect 3856 6296 3888 6328
rect 3928 6296 3960 6328
rect 40 6224 72 6256
rect 112 6224 144 6256
rect 184 6224 216 6256
rect 256 6224 288 6256
rect 328 6224 360 6256
rect 400 6224 432 6256
rect 472 6224 504 6256
rect 544 6224 576 6256
rect 616 6224 648 6256
rect 688 6224 720 6256
rect 760 6224 792 6256
rect 832 6224 864 6256
rect 904 6224 936 6256
rect 976 6224 1008 6256
rect 1048 6224 1080 6256
rect 1120 6224 1152 6256
rect 1192 6224 1224 6256
rect 1264 6224 1296 6256
rect 1336 6224 1368 6256
rect 1408 6224 1440 6256
rect 1480 6224 1512 6256
rect 1552 6224 1584 6256
rect 1624 6224 1656 6256
rect 1696 6224 1728 6256
rect 1768 6224 1800 6256
rect 1840 6224 1872 6256
rect 1912 6224 1944 6256
rect 1984 6224 2016 6256
rect 2056 6224 2088 6256
rect 2128 6224 2160 6256
rect 2200 6224 2232 6256
rect 2272 6224 2304 6256
rect 2344 6224 2376 6256
rect 2416 6224 2448 6256
rect 2488 6224 2520 6256
rect 2560 6224 2592 6256
rect 2632 6224 2664 6256
rect 2704 6224 2736 6256
rect 2776 6224 2808 6256
rect 2848 6224 2880 6256
rect 2920 6224 2952 6256
rect 2992 6224 3024 6256
rect 3064 6224 3096 6256
rect 3136 6224 3168 6256
rect 3208 6224 3240 6256
rect 3280 6224 3312 6256
rect 3352 6224 3384 6256
rect 3424 6224 3456 6256
rect 3496 6224 3528 6256
rect 3568 6224 3600 6256
rect 3640 6224 3672 6256
rect 3712 6224 3744 6256
rect 3784 6224 3816 6256
rect 3856 6224 3888 6256
rect 3928 6224 3960 6256
rect 40 6152 72 6184
rect 112 6152 144 6184
rect 184 6152 216 6184
rect 256 6152 288 6184
rect 328 6152 360 6184
rect 400 6152 432 6184
rect 472 6152 504 6184
rect 544 6152 576 6184
rect 616 6152 648 6184
rect 688 6152 720 6184
rect 760 6152 792 6184
rect 832 6152 864 6184
rect 904 6152 936 6184
rect 976 6152 1008 6184
rect 1048 6152 1080 6184
rect 1120 6152 1152 6184
rect 1192 6152 1224 6184
rect 1264 6152 1296 6184
rect 1336 6152 1368 6184
rect 1408 6152 1440 6184
rect 1480 6152 1512 6184
rect 1552 6152 1584 6184
rect 1624 6152 1656 6184
rect 1696 6152 1728 6184
rect 1768 6152 1800 6184
rect 1840 6152 1872 6184
rect 1912 6152 1944 6184
rect 1984 6152 2016 6184
rect 2056 6152 2088 6184
rect 2128 6152 2160 6184
rect 2200 6152 2232 6184
rect 2272 6152 2304 6184
rect 2344 6152 2376 6184
rect 2416 6152 2448 6184
rect 2488 6152 2520 6184
rect 2560 6152 2592 6184
rect 2632 6152 2664 6184
rect 2704 6152 2736 6184
rect 2776 6152 2808 6184
rect 2848 6152 2880 6184
rect 2920 6152 2952 6184
rect 2992 6152 3024 6184
rect 3064 6152 3096 6184
rect 3136 6152 3168 6184
rect 3208 6152 3240 6184
rect 3280 6152 3312 6184
rect 3352 6152 3384 6184
rect 3424 6152 3456 6184
rect 3496 6152 3528 6184
rect 3568 6152 3600 6184
rect 3640 6152 3672 6184
rect 3712 6152 3744 6184
rect 3784 6152 3816 6184
rect 3856 6152 3888 6184
rect 3928 6152 3960 6184
rect 40 6080 72 6112
rect 112 6080 144 6112
rect 184 6080 216 6112
rect 256 6080 288 6112
rect 328 6080 360 6112
rect 400 6080 432 6112
rect 472 6080 504 6112
rect 544 6080 576 6112
rect 616 6080 648 6112
rect 688 6080 720 6112
rect 760 6080 792 6112
rect 832 6080 864 6112
rect 904 6080 936 6112
rect 976 6080 1008 6112
rect 1048 6080 1080 6112
rect 1120 6080 1152 6112
rect 1192 6080 1224 6112
rect 1264 6080 1296 6112
rect 1336 6080 1368 6112
rect 1408 6080 1440 6112
rect 1480 6080 1512 6112
rect 1552 6080 1584 6112
rect 1624 6080 1656 6112
rect 1696 6080 1728 6112
rect 1768 6080 1800 6112
rect 1840 6080 1872 6112
rect 1912 6080 1944 6112
rect 1984 6080 2016 6112
rect 2056 6080 2088 6112
rect 2128 6080 2160 6112
rect 2200 6080 2232 6112
rect 2272 6080 2304 6112
rect 2344 6080 2376 6112
rect 2416 6080 2448 6112
rect 2488 6080 2520 6112
rect 2560 6080 2592 6112
rect 2632 6080 2664 6112
rect 2704 6080 2736 6112
rect 2776 6080 2808 6112
rect 2848 6080 2880 6112
rect 2920 6080 2952 6112
rect 2992 6080 3024 6112
rect 3064 6080 3096 6112
rect 3136 6080 3168 6112
rect 3208 6080 3240 6112
rect 3280 6080 3312 6112
rect 3352 6080 3384 6112
rect 3424 6080 3456 6112
rect 3496 6080 3528 6112
rect 3568 6080 3600 6112
rect 3640 6080 3672 6112
rect 3712 6080 3744 6112
rect 3784 6080 3816 6112
rect 3856 6080 3888 6112
rect 3928 6080 3960 6112
rect 40 6008 72 6040
rect 112 6008 144 6040
rect 184 6008 216 6040
rect 256 6008 288 6040
rect 328 6008 360 6040
rect 400 6008 432 6040
rect 472 6008 504 6040
rect 544 6008 576 6040
rect 616 6008 648 6040
rect 688 6008 720 6040
rect 760 6008 792 6040
rect 832 6008 864 6040
rect 904 6008 936 6040
rect 976 6008 1008 6040
rect 1048 6008 1080 6040
rect 1120 6008 1152 6040
rect 1192 6008 1224 6040
rect 1264 6008 1296 6040
rect 1336 6008 1368 6040
rect 1408 6008 1440 6040
rect 1480 6008 1512 6040
rect 1552 6008 1584 6040
rect 1624 6008 1656 6040
rect 1696 6008 1728 6040
rect 1768 6008 1800 6040
rect 1840 6008 1872 6040
rect 1912 6008 1944 6040
rect 1984 6008 2016 6040
rect 2056 6008 2088 6040
rect 2128 6008 2160 6040
rect 2200 6008 2232 6040
rect 2272 6008 2304 6040
rect 2344 6008 2376 6040
rect 2416 6008 2448 6040
rect 2488 6008 2520 6040
rect 2560 6008 2592 6040
rect 2632 6008 2664 6040
rect 2704 6008 2736 6040
rect 2776 6008 2808 6040
rect 2848 6008 2880 6040
rect 2920 6008 2952 6040
rect 2992 6008 3024 6040
rect 3064 6008 3096 6040
rect 3136 6008 3168 6040
rect 3208 6008 3240 6040
rect 3280 6008 3312 6040
rect 3352 6008 3384 6040
rect 3424 6008 3456 6040
rect 3496 6008 3528 6040
rect 3568 6008 3600 6040
rect 3640 6008 3672 6040
rect 3712 6008 3744 6040
rect 3784 6008 3816 6040
rect 3856 6008 3888 6040
rect 3928 6008 3960 6040
rect 40 5936 72 5968
rect 112 5936 144 5968
rect 184 5936 216 5968
rect 256 5936 288 5968
rect 328 5936 360 5968
rect 400 5936 432 5968
rect 472 5936 504 5968
rect 544 5936 576 5968
rect 616 5936 648 5968
rect 688 5936 720 5968
rect 760 5936 792 5968
rect 832 5936 864 5968
rect 904 5936 936 5968
rect 976 5936 1008 5968
rect 1048 5936 1080 5968
rect 1120 5936 1152 5968
rect 1192 5936 1224 5968
rect 1264 5936 1296 5968
rect 1336 5936 1368 5968
rect 1408 5936 1440 5968
rect 1480 5936 1512 5968
rect 1552 5936 1584 5968
rect 1624 5936 1656 5968
rect 1696 5936 1728 5968
rect 1768 5936 1800 5968
rect 1840 5936 1872 5968
rect 1912 5936 1944 5968
rect 1984 5936 2016 5968
rect 2056 5936 2088 5968
rect 2128 5936 2160 5968
rect 2200 5936 2232 5968
rect 2272 5936 2304 5968
rect 2344 5936 2376 5968
rect 2416 5936 2448 5968
rect 2488 5936 2520 5968
rect 2560 5936 2592 5968
rect 2632 5936 2664 5968
rect 2704 5936 2736 5968
rect 2776 5936 2808 5968
rect 2848 5936 2880 5968
rect 2920 5936 2952 5968
rect 2992 5936 3024 5968
rect 3064 5936 3096 5968
rect 3136 5936 3168 5968
rect 3208 5936 3240 5968
rect 3280 5936 3312 5968
rect 3352 5936 3384 5968
rect 3424 5936 3456 5968
rect 3496 5936 3528 5968
rect 3568 5936 3600 5968
rect 3640 5936 3672 5968
rect 3712 5936 3744 5968
rect 3784 5936 3816 5968
rect 3856 5936 3888 5968
rect 3928 5936 3960 5968
rect 40 5864 72 5896
rect 112 5864 144 5896
rect 184 5864 216 5896
rect 256 5864 288 5896
rect 328 5864 360 5896
rect 400 5864 432 5896
rect 472 5864 504 5896
rect 544 5864 576 5896
rect 616 5864 648 5896
rect 688 5864 720 5896
rect 760 5864 792 5896
rect 832 5864 864 5896
rect 904 5864 936 5896
rect 976 5864 1008 5896
rect 1048 5864 1080 5896
rect 1120 5864 1152 5896
rect 1192 5864 1224 5896
rect 1264 5864 1296 5896
rect 1336 5864 1368 5896
rect 1408 5864 1440 5896
rect 1480 5864 1512 5896
rect 1552 5864 1584 5896
rect 1624 5864 1656 5896
rect 1696 5864 1728 5896
rect 1768 5864 1800 5896
rect 1840 5864 1872 5896
rect 1912 5864 1944 5896
rect 1984 5864 2016 5896
rect 2056 5864 2088 5896
rect 2128 5864 2160 5896
rect 2200 5864 2232 5896
rect 2272 5864 2304 5896
rect 2344 5864 2376 5896
rect 2416 5864 2448 5896
rect 2488 5864 2520 5896
rect 2560 5864 2592 5896
rect 2632 5864 2664 5896
rect 2704 5864 2736 5896
rect 2776 5864 2808 5896
rect 2848 5864 2880 5896
rect 2920 5864 2952 5896
rect 2992 5864 3024 5896
rect 3064 5864 3096 5896
rect 3136 5864 3168 5896
rect 3208 5864 3240 5896
rect 3280 5864 3312 5896
rect 3352 5864 3384 5896
rect 3424 5864 3456 5896
rect 3496 5864 3528 5896
rect 3568 5864 3600 5896
rect 3640 5864 3672 5896
rect 3712 5864 3744 5896
rect 3784 5864 3816 5896
rect 3856 5864 3888 5896
rect 3928 5864 3960 5896
rect 40 5792 72 5824
rect 112 5792 144 5824
rect 184 5792 216 5824
rect 256 5792 288 5824
rect 328 5792 360 5824
rect 400 5792 432 5824
rect 472 5792 504 5824
rect 544 5792 576 5824
rect 616 5792 648 5824
rect 688 5792 720 5824
rect 760 5792 792 5824
rect 832 5792 864 5824
rect 904 5792 936 5824
rect 976 5792 1008 5824
rect 1048 5792 1080 5824
rect 1120 5792 1152 5824
rect 1192 5792 1224 5824
rect 1264 5792 1296 5824
rect 1336 5792 1368 5824
rect 1408 5792 1440 5824
rect 1480 5792 1512 5824
rect 1552 5792 1584 5824
rect 1624 5792 1656 5824
rect 1696 5792 1728 5824
rect 1768 5792 1800 5824
rect 1840 5792 1872 5824
rect 1912 5792 1944 5824
rect 1984 5792 2016 5824
rect 2056 5792 2088 5824
rect 2128 5792 2160 5824
rect 2200 5792 2232 5824
rect 2272 5792 2304 5824
rect 2344 5792 2376 5824
rect 2416 5792 2448 5824
rect 2488 5792 2520 5824
rect 2560 5792 2592 5824
rect 2632 5792 2664 5824
rect 2704 5792 2736 5824
rect 2776 5792 2808 5824
rect 2848 5792 2880 5824
rect 2920 5792 2952 5824
rect 2992 5792 3024 5824
rect 3064 5792 3096 5824
rect 3136 5792 3168 5824
rect 3208 5792 3240 5824
rect 3280 5792 3312 5824
rect 3352 5792 3384 5824
rect 3424 5792 3456 5824
rect 3496 5792 3528 5824
rect 3568 5792 3600 5824
rect 3640 5792 3672 5824
rect 3712 5792 3744 5824
rect 3784 5792 3816 5824
rect 3856 5792 3888 5824
rect 3928 5792 3960 5824
rect 40 5720 72 5752
rect 112 5720 144 5752
rect 184 5720 216 5752
rect 256 5720 288 5752
rect 328 5720 360 5752
rect 400 5720 432 5752
rect 472 5720 504 5752
rect 544 5720 576 5752
rect 616 5720 648 5752
rect 688 5720 720 5752
rect 760 5720 792 5752
rect 832 5720 864 5752
rect 904 5720 936 5752
rect 976 5720 1008 5752
rect 1048 5720 1080 5752
rect 1120 5720 1152 5752
rect 1192 5720 1224 5752
rect 1264 5720 1296 5752
rect 1336 5720 1368 5752
rect 1408 5720 1440 5752
rect 1480 5720 1512 5752
rect 1552 5720 1584 5752
rect 1624 5720 1656 5752
rect 1696 5720 1728 5752
rect 1768 5720 1800 5752
rect 1840 5720 1872 5752
rect 1912 5720 1944 5752
rect 1984 5720 2016 5752
rect 2056 5720 2088 5752
rect 2128 5720 2160 5752
rect 2200 5720 2232 5752
rect 2272 5720 2304 5752
rect 2344 5720 2376 5752
rect 2416 5720 2448 5752
rect 2488 5720 2520 5752
rect 2560 5720 2592 5752
rect 2632 5720 2664 5752
rect 2704 5720 2736 5752
rect 2776 5720 2808 5752
rect 2848 5720 2880 5752
rect 2920 5720 2952 5752
rect 2992 5720 3024 5752
rect 3064 5720 3096 5752
rect 3136 5720 3168 5752
rect 3208 5720 3240 5752
rect 3280 5720 3312 5752
rect 3352 5720 3384 5752
rect 3424 5720 3456 5752
rect 3496 5720 3528 5752
rect 3568 5720 3600 5752
rect 3640 5720 3672 5752
rect 3712 5720 3744 5752
rect 3784 5720 3816 5752
rect 3856 5720 3888 5752
rect 3928 5720 3960 5752
rect 40 5648 72 5680
rect 112 5648 144 5680
rect 184 5648 216 5680
rect 256 5648 288 5680
rect 328 5648 360 5680
rect 400 5648 432 5680
rect 472 5648 504 5680
rect 544 5648 576 5680
rect 616 5648 648 5680
rect 688 5648 720 5680
rect 760 5648 792 5680
rect 832 5648 864 5680
rect 904 5648 936 5680
rect 976 5648 1008 5680
rect 1048 5648 1080 5680
rect 1120 5648 1152 5680
rect 1192 5648 1224 5680
rect 1264 5648 1296 5680
rect 1336 5648 1368 5680
rect 1408 5648 1440 5680
rect 1480 5648 1512 5680
rect 1552 5648 1584 5680
rect 1624 5648 1656 5680
rect 1696 5648 1728 5680
rect 1768 5648 1800 5680
rect 1840 5648 1872 5680
rect 1912 5648 1944 5680
rect 1984 5648 2016 5680
rect 2056 5648 2088 5680
rect 2128 5648 2160 5680
rect 2200 5648 2232 5680
rect 2272 5648 2304 5680
rect 2344 5648 2376 5680
rect 2416 5648 2448 5680
rect 2488 5648 2520 5680
rect 2560 5648 2592 5680
rect 2632 5648 2664 5680
rect 2704 5648 2736 5680
rect 2776 5648 2808 5680
rect 2848 5648 2880 5680
rect 2920 5648 2952 5680
rect 2992 5648 3024 5680
rect 3064 5648 3096 5680
rect 3136 5648 3168 5680
rect 3208 5648 3240 5680
rect 3280 5648 3312 5680
rect 3352 5648 3384 5680
rect 3424 5648 3456 5680
rect 3496 5648 3528 5680
rect 3568 5648 3600 5680
rect 3640 5648 3672 5680
rect 3712 5648 3744 5680
rect 3784 5648 3816 5680
rect 3856 5648 3888 5680
rect 3928 5648 3960 5680
rect 40 5576 72 5608
rect 112 5576 144 5608
rect 184 5576 216 5608
rect 256 5576 288 5608
rect 328 5576 360 5608
rect 400 5576 432 5608
rect 472 5576 504 5608
rect 544 5576 576 5608
rect 616 5576 648 5608
rect 688 5576 720 5608
rect 760 5576 792 5608
rect 832 5576 864 5608
rect 904 5576 936 5608
rect 976 5576 1008 5608
rect 1048 5576 1080 5608
rect 1120 5576 1152 5608
rect 1192 5576 1224 5608
rect 1264 5576 1296 5608
rect 1336 5576 1368 5608
rect 1408 5576 1440 5608
rect 1480 5576 1512 5608
rect 1552 5576 1584 5608
rect 1624 5576 1656 5608
rect 1696 5576 1728 5608
rect 1768 5576 1800 5608
rect 1840 5576 1872 5608
rect 1912 5576 1944 5608
rect 1984 5576 2016 5608
rect 2056 5576 2088 5608
rect 2128 5576 2160 5608
rect 2200 5576 2232 5608
rect 2272 5576 2304 5608
rect 2344 5576 2376 5608
rect 2416 5576 2448 5608
rect 2488 5576 2520 5608
rect 2560 5576 2592 5608
rect 2632 5576 2664 5608
rect 2704 5576 2736 5608
rect 2776 5576 2808 5608
rect 2848 5576 2880 5608
rect 2920 5576 2952 5608
rect 2992 5576 3024 5608
rect 3064 5576 3096 5608
rect 3136 5576 3168 5608
rect 3208 5576 3240 5608
rect 3280 5576 3312 5608
rect 3352 5576 3384 5608
rect 3424 5576 3456 5608
rect 3496 5576 3528 5608
rect 3568 5576 3600 5608
rect 3640 5576 3672 5608
rect 3712 5576 3744 5608
rect 3784 5576 3816 5608
rect 3856 5576 3888 5608
rect 3928 5576 3960 5608
rect 40 5504 72 5536
rect 112 5504 144 5536
rect 184 5504 216 5536
rect 256 5504 288 5536
rect 328 5504 360 5536
rect 400 5504 432 5536
rect 472 5504 504 5536
rect 544 5504 576 5536
rect 616 5504 648 5536
rect 688 5504 720 5536
rect 760 5504 792 5536
rect 832 5504 864 5536
rect 904 5504 936 5536
rect 976 5504 1008 5536
rect 1048 5504 1080 5536
rect 1120 5504 1152 5536
rect 1192 5504 1224 5536
rect 1264 5504 1296 5536
rect 1336 5504 1368 5536
rect 1408 5504 1440 5536
rect 1480 5504 1512 5536
rect 1552 5504 1584 5536
rect 1624 5504 1656 5536
rect 1696 5504 1728 5536
rect 1768 5504 1800 5536
rect 1840 5504 1872 5536
rect 1912 5504 1944 5536
rect 1984 5504 2016 5536
rect 2056 5504 2088 5536
rect 2128 5504 2160 5536
rect 2200 5504 2232 5536
rect 2272 5504 2304 5536
rect 2344 5504 2376 5536
rect 2416 5504 2448 5536
rect 2488 5504 2520 5536
rect 2560 5504 2592 5536
rect 2632 5504 2664 5536
rect 2704 5504 2736 5536
rect 2776 5504 2808 5536
rect 2848 5504 2880 5536
rect 2920 5504 2952 5536
rect 2992 5504 3024 5536
rect 3064 5504 3096 5536
rect 3136 5504 3168 5536
rect 3208 5504 3240 5536
rect 3280 5504 3312 5536
rect 3352 5504 3384 5536
rect 3424 5504 3456 5536
rect 3496 5504 3528 5536
rect 3568 5504 3600 5536
rect 3640 5504 3672 5536
rect 3712 5504 3744 5536
rect 3784 5504 3816 5536
rect 3856 5504 3888 5536
rect 3928 5504 3960 5536
rect 40 5432 72 5464
rect 112 5432 144 5464
rect 184 5432 216 5464
rect 256 5432 288 5464
rect 328 5432 360 5464
rect 400 5432 432 5464
rect 472 5432 504 5464
rect 544 5432 576 5464
rect 616 5432 648 5464
rect 688 5432 720 5464
rect 760 5432 792 5464
rect 832 5432 864 5464
rect 904 5432 936 5464
rect 976 5432 1008 5464
rect 1048 5432 1080 5464
rect 1120 5432 1152 5464
rect 1192 5432 1224 5464
rect 1264 5432 1296 5464
rect 1336 5432 1368 5464
rect 1408 5432 1440 5464
rect 1480 5432 1512 5464
rect 1552 5432 1584 5464
rect 1624 5432 1656 5464
rect 1696 5432 1728 5464
rect 1768 5432 1800 5464
rect 1840 5432 1872 5464
rect 1912 5432 1944 5464
rect 1984 5432 2016 5464
rect 2056 5432 2088 5464
rect 2128 5432 2160 5464
rect 2200 5432 2232 5464
rect 2272 5432 2304 5464
rect 2344 5432 2376 5464
rect 2416 5432 2448 5464
rect 2488 5432 2520 5464
rect 2560 5432 2592 5464
rect 2632 5432 2664 5464
rect 2704 5432 2736 5464
rect 2776 5432 2808 5464
rect 2848 5432 2880 5464
rect 2920 5432 2952 5464
rect 2992 5432 3024 5464
rect 3064 5432 3096 5464
rect 3136 5432 3168 5464
rect 3208 5432 3240 5464
rect 3280 5432 3312 5464
rect 3352 5432 3384 5464
rect 3424 5432 3456 5464
rect 3496 5432 3528 5464
rect 3568 5432 3600 5464
rect 3640 5432 3672 5464
rect 3712 5432 3744 5464
rect 3784 5432 3816 5464
rect 3856 5432 3888 5464
rect 3928 5432 3960 5464
rect 40 5360 72 5392
rect 112 5360 144 5392
rect 184 5360 216 5392
rect 256 5360 288 5392
rect 328 5360 360 5392
rect 400 5360 432 5392
rect 472 5360 504 5392
rect 544 5360 576 5392
rect 616 5360 648 5392
rect 688 5360 720 5392
rect 760 5360 792 5392
rect 832 5360 864 5392
rect 904 5360 936 5392
rect 976 5360 1008 5392
rect 1048 5360 1080 5392
rect 1120 5360 1152 5392
rect 1192 5360 1224 5392
rect 1264 5360 1296 5392
rect 1336 5360 1368 5392
rect 1408 5360 1440 5392
rect 1480 5360 1512 5392
rect 1552 5360 1584 5392
rect 1624 5360 1656 5392
rect 1696 5360 1728 5392
rect 1768 5360 1800 5392
rect 1840 5360 1872 5392
rect 1912 5360 1944 5392
rect 1984 5360 2016 5392
rect 2056 5360 2088 5392
rect 2128 5360 2160 5392
rect 2200 5360 2232 5392
rect 2272 5360 2304 5392
rect 2344 5360 2376 5392
rect 2416 5360 2448 5392
rect 2488 5360 2520 5392
rect 2560 5360 2592 5392
rect 2632 5360 2664 5392
rect 2704 5360 2736 5392
rect 2776 5360 2808 5392
rect 2848 5360 2880 5392
rect 2920 5360 2952 5392
rect 2992 5360 3024 5392
rect 3064 5360 3096 5392
rect 3136 5360 3168 5392
rect 3208 5360 3240 5392
rect 3280 5360 3312 5392
rect 3352 5360 3384 5392
rect 3424 5360 3456 5392
rect 3496 5360 3528 5392
rect 3568 5360 3600 5392
rect 3640 5360 3672 5392
rect 3712 5360 3744 5392
rect 3784 5360 3816 5392
rect 3856 5360 3888 5392
rect 3928 5360 3960 5392
rect 40 5288 72 5320
rect 112 5288 144 5320
rect 184 5288 216 5320
rect 256 5288 288 5320
rect 328 5288 360 5320
rect 400 5288 432 5320
rect 472 5288 504 5320
rect 544 5288 576 5320
rect 616 5288 648 5320
rect 688 5288 720 5320
rect 760 5288 792 5320
rect 832 5288 864 5320
rect 904 5288 936 5320
rect 976 5288 1008 5320
rect 1048 5288 1080 5320
rect 1120 5288 1152 5320
rect 1192 5288 1224 5320
rect 1264 5288 1296 5320
rect 1336 5288 1368 5320
rect 1408 5288 1440 5320
rect 1480 5288 1512 5320
rect 1552 5288 1584 5320
rect 1624 5288 1656 5320
rect 1696 5288 1728 5320
rect 1768 5288 1800 5320
rect 1840 5288 1872 5320
rect 1912 5288 1944 5320
rect 1984 5288 2016 5320
rect 2056 5288 2088 5320
rect 2128 5288 2160 5320
rect 2200 5288 2232 5320
rect 2272 5288 2304 5320
rect 2344 5288 2376 5320
rect 2416 5288 2448 5320
rect 2488 5288 2520 5320
rect 2560 5288 2592 5320
rect 2632 5288 2664 5320
rect 2704 5288 2736 5320
rect 2776 5288 2808 5320
rect 2848 5288 2880 5320
rect 2920 5288 2952 5320
rect 2992 5288 3024 5320
rect 3064 5288 3096 5320
rect 3136 5288 3168 5320
rect 3208 5288 3240 5320
rect 3280 5288 3312 5320
rect 3352 5288 3384 5320
rect 3424 5288 3456 5320
rect 3496 5288 3528 5320
rect 3568 5288 3600 5320
rect 3640 5288 3672 5320
rect 3712 5288 3744 5320
rect 3784 5288 3816 5320
rect 3856 5288 3888 5320
rect 3928 5288 3960 5320
rect 40 5216 72 5248
rect 112 5216 144 5248
rect 184 5216 216 5248
rect 256 5216 288 5248
rect 328 5216 360 5248
rect 400 5216 432 5248
rect 472 5216 504 5248
rect 544 5216 576 5248
rect 616 5216 648 5248
rect 688 5216 720 5248
rect 760 5216 792 5248
rect 832 5216 864 5248
rect 904 5216 936 5248
rect 976 5216 1008 5248
rect 1048 5216 1080 5248
rect 1120 5216 1152 5248
rect 1192 5216 1224 5248
rect 1264 5216 1296 5248
rect 1336 5216 1368 5248
rect 1408 5216 1440 5248
rect 1480 5216 1512 5248
rect 1552 5216 1584 5248
rect 1624 5216 1656 5248
rect 1696 5216 1728 5248
rect 1768 5216 1800 5248
rect 1840 5216 1872 5248
rect 1912 5216 1944 5248
rect 1984 5216 2016 5248
rect 2056 5216 2088 5248
rect 2128 5216 2160 5248
rect 2200 5216 2232 5248
rect 2272 5216 2304 5248
rect 2344 5216 2376 5248
rect 2416 5216 2448 5248
rect 2488 5216 2520 5248
rect 2560 5216 2592 5248
rect 2632 5216 2664 5248
rect 2704 5216 2736 5248
rect 2776 5216 2808 5248
rect 2848 5216 2880 5248
rect 2920 5216 2952 5248
rect 2992 5216 3024 5248
rect 3064 5216 3096 5248
rect 3136 5216 3168 5248
rect 3208 5216 3240 5248
rect 3280 5216 3312 5248
rect 3352 5216 3384 5248
rect 3424 5216 3456 5248
rect 3496 5216 3528 5248
rect 3568 5216 3600 5248
rect 3640 5216 3672 5248
rect 3712 5216 3744 5248
rect 3784 5216 3816 5248
rect 3856 5216 3888 5248
rect 3928 5216 3960 5248
rect 40 5144 72 5176
rect 112 5144 144 5176
rect 184 5144 216 5176
rect 256 5144 288 5176
rect 328 5144 360 5176
rect 400 5144 432 5176
rect 472 5144 504 5176
rect 544 5144 576 5176
rect 616 5144 648 5176
rect 688 5144 720 5176
rect 760 5144 792 5176
rect 832 5144 864 5176
rect 904 5144 936 5176
rect 976 5144 1008 5176
rect 1048 5144 1080 5176
rect 1120 5144 1152 5176
rect 1192 5144 1224 5176
rect 1264 5144 1296 5176
rect 1336 5144 1368 5176
rect 1408 5144 1440 5176
rect 1480 5144 1512 5176
rect 1552 5144 1584 5176
rect 1624 5144 1656 5176
rect 1696 5144 1728 5176
rect 1768 5144 1800 5176
rect 1840 5144 1872 5176
rect 1912 5144 1944 5176
rect 1984 5144 2016 5176
rect 2056 5144 2088 5176
rect 2128 5144 2160 5176
rect 2200 5144 2232 5176
rect 2272 5144 2304 5176
rect 2344 5144 2376 5176
rect 2416 5144 2448 5176
rect 2488 5144 2520 5176
rect 2560 5144 2592 5176
rect 2632 5144 2664 5176
rect 2704 5144 2736 5176
rect 2776 5144 2808 5176
rect 2848 5144 2880 5176
rect 2920 5144 2952 5176
rect 2992 5144 3024 5176
rect 3064 5144 3096 5176
rect 3136 5144 3168 5176
rect 3208 5144 3240 5176
rect 3280 5144 3312 5176
rect 3352 5144 3384 5176
rect 3424 5144 3456 5176
rect 3496 5144 3528 5176
rect 3568 5144 3600 5176
rect 3640 5144 3672 5176
rect 3712 5144 3744 5176
rect 3784 5144 3816 5176
rect 3856 5144 3888 5176
rect 3928 5144 3960 5176
rect 40 5072 72 5104
rect 112 5072 144 5104
rect 184 5072 216 5104
rect 256 5072 288 5104
rect 328 5072 360 5104
rect 400 5072 432 5104
rect 472 5072 504 5104
rect 544 5072 576 5104
rect 616 5072 648 5104
rect 688 5072 720 5104
rect 760 5072 792 5104
rect 832 5072 864 5104
rect 904 5072 936 5104
rect 976 5072 1008 5104
rect 1048 5072 1080 5104
rect 1120 5072 1152 5104
rect 1192 5072 1224 5104
rect 1264 5072 1296 5104
rect 1336 5072 1368 5104
rect 1408 5072 1440 5104
rect 1480 5072 1512 5104
rect 1552 5072 1584 5104
rect 1624 5072 1656 5104
rect 1696 5072 1728 5104
rect 1768 5072 1800 5104
rect 1840 5072 1872 5104
rect 1912 5072 1944 5104
rect 1984 5072 2016 5104
rect 2056 5072 2088 5104
rect 2128 5072 2160 5104
rect 2200 5072 2232 5104
rect 2272 5072 2304 5104
rect 2344 5072 2376 5104
rect 2416 5072 2448 5104
rect 2488 5072 2520 5104
rect 2560 5072 2592 5104
rect 2632 5072 2664 5104
rect 2704 5072 2736 5104
rect 2776 5072 2808 5104
rect 2848 5072 2880 5104
rect 2920 5072 2952 5104
rect 2992 5072 3024 5104
rect 3064 5072 3096 5104
rect 3136 5072 3168 5104
rect 3208 5072 3240 5104
rect 3280 5072 3312 5104
rect 3352 5072 3384 5104
rect 3424 5072 3456 5104
rect 3496 5072 3528 5104
rect 3568 5072 3600 5104
rect 3640 5072 3672 5104
rect 3712 5072 3744 5104
rect 3784 5072 3816 5104
rect 3856 5072 3888 5104
rect 3928 5072 3960 5104
rect 40 5000 72 5032
rect 112 5000 144 5032
rect 184 5000 216 5032
rect 256 5000 288 5032
rect 328 5000 360 5032
rect 400 5000 432 5032
rect 472 5000 504 5032
rect 544 5000 576 5032
rect 616 5000 648 5032
rect 688 5000 720 5032
rect 760 5000 792 5032
rect 832 5000 864 5032
rect 904 5000 936 5032
rect 976 5000 1008 5032
rect 1048 5000 1080 5032
rect 1120 5000 1152 5032
rect 1192 5000 1224 5032
rect 1264 5000 1296 5032
rect 1336 5000 1368 5032
rect 1408 5000 1440 5032
rect 1480 5000 1512 5032
rect 1552 5000 1584 5032
rect 1624 5000 1656 5032
rect 1696 5000 1728 5032
rect 1768 5000 1800 5032
rect 1840 5000 1872 5032
rect 1912 5000 1944 5032
rect 1984 5000 2016 5032
rect 2056 5000 2088 5032
rect 2128 5000 2160 5032
rect 2200 5000 2232 5032
rect 2272 5000 2304 5032
rect 2344 5000 2376 5032
rect 2416 5000 2448 5032
rect 2488 5000 2520 5032
rect 2560 5000 2592 5032
rect 2632 5000 2664 5032
rect 2704 5000 2736 5032
rect 2776 5000 2808 5032
rect 2848 5000 2880 5032
rect 2920 5000 2952 5032
rect 2992 5000 3024 5032
rect 3064 5000 3096 5032
rect 3136 5000 3168 5032
rect 3208 5000 3240 5032
rect 3280 5000 3312 5032
rect 3352 5000 3384 5032
rect 3424 5000 3456 5032
rect 3496 5000 3528 5032
rect 3568 5000 3600 5032
rect 3640 5000 3672 5032
rect 3712 5000 3744 5032
rect 3784 5000 3816 5032
rect 3856 5000 3888 5032
rect 3928 5000 3960 5032
rect 40 4928 72 4960
rect 112 4928 144 4960
rect 184 4928 216 4960
rect 256 4928 288 4960
rect 328 4928 360 4960
rect 400 4928 432 4960
rect 472 4928 504 4960
rect 544 4928 576 4960
rect 616 4928 648 4960
rect 688 4928 720 4960
rect 760 4928 792 4960
rect 832 4928 864 4960
rect 904 4928 936 4960
rect 976 4928 1008 4960
rect 1048 4928 1080 4960
rect 1120 4928 1152 4960
rect 1192 4928 1224 4960
rect 1264 4928 1296 4960
rect 1336 4928 1368 4960
rect 1408 4928 1440 4960
rect 1480 4928 1512 4960
rect 1552 4928 1584 4960
rect 1624 4928 1656 4960
rect 1696 4928 1728 4960
rect 1768 4928 1800 4960
rect 1840 4928 1872 4960
rect 1912 4928 1944 4960
rect 1984 4928 2016 4960
rect 2056 4928 2088 4960
rect 2128 4928 2160 4960
rect 2200 4928 2232 4960
rect 2272 4928 2304 4960
rect 2344 4928 2376 4960
rect 2416 4928 2448 4960
rect 2488 4928 2520 4960
rect 2560 4928 2592 4960
rect 2632 4928 2664 4960
rect 2704 4928 2736 4960
rect 2776 4928 2808 4960
rect 2848 4928 2880 4960
rect 2920 4928 2952 4960
rect 2992 4928 3024 4960
rect 3064 4928 3096 4960
rect 3136 4928 3168 4960
rect 3208 4928 3240 4960
rect 3280 4928 3312 4960
rect 3352 4928 3384 4960
rect 3424 4928 3456 4960
rect 3496 4928 3528 4960
rect 3568 4928 3600 4960
rect 3640 4928 3672 4960
rect 3712 4928 3744 4960
rect 3784 4928 3816 4960
rect 3856 4928 3888 4960
rect 3928 4928 3960 4960
rect 40 4856 72 4888
rect 112 4856 144 4888
rect 184 4856 216 4888
rect 256 4856 288 4888
rect 328 4856 360 4888
rect 400 4856 432 4888
rect 472 4856 504 4888
rect 544 4856 576 4888
rect 616 4856 648 4888
rect 688 4856 720 4888
rect 760 4856 792 4888
rect 832 4856 864 4888
rect 904 4856 936 4888
rect 976 4856 1008 4888
rect 1048 4856 1080 4888
rect 1120 4856 1152 4888
rect 1192 4856 1224 4888
rect 1264 4856 1296 4888
rect 1336 4856 1368 4888
rect 1408 4856 1440 4888
rect 1480 4856 1512 4888
rect 1552 4856 1584 4888
rect 1624 4856 1656 4888
rect 1696 4856 1728 4888
rect 1768 4856 1800 4888
rect 1840 4856 1872 4888
rect 1912 4856 1944 4888
rect 1984 4856 2016 4888
rect 2056 4856 2088 4888
rect 2128 4856 2160 4888
rect 2200 4856 2232 4888
rect 2272 4856 2304 4888
rect 2344 4856 2376 4888
rect 2416 4856 2448 4888
rect 2488 4856 2520 4888
rect 2560 4856 2592 4888
rect 2632 4856 2664 4888
rect 2704 4856 2736 4888
rect 2776 4856 2808 4888
rect 2848 4856 2880 4888
rect 2920 4856 2952 4888
rect 2992 4856 3024 4888
rect 3064 4856 3096 4888
rect 3136 4856 3168 4888
rect 3208 4856 3240 4888
rect 3280 4856 3312 4888
rect 3352 4856 3384 4888
rect 3424 4856 3456 4888
rect 3496 4856 3528 4888
rect 3568 4856 3600 4888
rect 3640 4856 3672 4888
rect 3712 4856 3744 4888
rect 3784 4856 3816 4888
rect 3856 4856 3888 4888
rect 3928 4856 3960 4888
rect 40 4784 72 4816
rect 112 4784 144 4816
rect 184 4784 216 4816
rect 256 4784 288 4816
rect 328 4784 360 4816
rect 400 4784 432 4816
rect 472 4784 504 4816
rect 544 4784 576 4816
rect 616 4784 648 4816
rect 688 4784 720 4816
rect 760 4784 792 4816
rect 832 4784 864 4816
rect 904 4784 936 4816
rect 976 4784 1008 4816
rect 1048 4784 1080 4816
rect 1120 4784 1152 4816
rect 1192 4784 1224 4816
rect 1264 4784 1296 4816
rect 1336 4784 1368 4816
rect 1408 4784 1440 4816
rect 1480 4784 1512 4816
rect 1552 4784 1584 4816
rect 1624 4784 1656 4816
rect 1696 4784 1728 4816
rect 1768 4784 1800 4816
rect 1840 4784 1872 4816
rect 1912 4784 1944 4816
rect 1984 4784 2016 4816
rect 2056 4784 2088 4816
rect 2128 4784 2160 4816
rect 2200 4784 2232 4816
rect 2272 4784 2304 4816
rect 2344 4784 2376 4816
rect 2416 4784 2448 4816
rect 2488 4784 2520 4816
rect 2560 4784 2592 4816
rect 2632 4784 2664 4816
rect 2704 4784 2736 4816
rect 2776 4784 2808 4816
rect 2848 4784 2880 4816
rect 2920 4784 2952 4816
rect 2992 4784 3024 4816
rect 3064 4784 3096 4816
rect 3136 4784 3168 4816
rect 3208 4784 3240 4816
rect 3280 4784 3312 4816
rect 3352 4784 3384 4816
rect 3424 4784 3456 4816
rect 3496 4784 3528 4816
rect 3568 4784 3600 4816
rect 3640 4784 3672 4816
rect 3712 4784 3744 4816
rect 3784 4784 3816 4816
rect 3856 4784 3888 4816
rect 3928 4784 3960 4816
rect 40 4712 72 4744
rect 112 4712 144 4744
rect 184 4712 216 4744
rect 256 4712 288 4744
rect 328 4712 360 4744
rect 400 4712 432 4744
rect 472 4712 504 4744
rect 544 4712 576 4744
rect 616 4712 648 4744
rect 688 4712 720 4744
rect 760 4712 792 4744
rect 832 4712 864 4744
rect 904 4712 936 4744
rect 976 4712 1008 4744
rect 1048 4712 1080 4744
rect 1120 4712 1152 4744
rect 1192 4712 1224 4744
rect 1264 4712 1296 4744
rect 1336 4712 1368 4744
rect 1408 4712 1440 4744
rect 1480 4712 1512 4744
rect 1552 4712 1584 4744
rect 1624 4712 1656 4744
rect 1696 4712 1728 4744
rect 1768 4712 1800 4744
rect 1840 4712 1872 4744
rect 1912 4712 1944 4744
rect 1984 4712 2016 4744
rect 2056 4712 2088 4744
rect 2128 4712 2160 4744
rect 2200 4712 2232 4744
rect 2272 4712 2304 4744
rect 2344 4712 2376 4744
rect 2416 4712 2448 4744
rect 2488 4712 2520 4744
rect 2560 4712 2592 4744
rect 2632 4712 2664 4744
rect 2704 4712 2736 4744
rect 2776 4712 2808 4744
rect 2848 4712 2880 4744
rect 2920 4712 2952 4744
rect 2992 4712 3024 4744
rect 3064 4712 3096 4744
rect 3136 4712 3168 4744
rect 3208 4712 3240 4744
rect 3280 4712 3312 4744
rect 3352 4712 3384 4744
rect 3424 4712 3456 4744
rect 3496 4712 3528 4744
rect 3568 4712 3600 4744
rect 3640 4712 3672 4744
rect 3712 4712 3744 4744
rect 3784 4712 3816 4744
rect 3856 4712 3888 4744
rect 3928 4712 3960 4744
rect 40 4640 72 4672
rect 112 4640 144 4672
rect 184 4640 216 4672
rect 256 4640 288 4672
rect 328 4640 360 4672
rect 400 4640 432 4672
rect 472 4640 504 4672
rect 544 4640 576 4672
rect 616 4640 648 4672
rect 688 4640 720 4672
rect 760 4640 792 4672
rect 832 4640 864 4672
rect 904 4640 936 4672
rect 976 4640 1008 4672
rect 1048 4640 1080 4672
rect 1120 4640 1152 4672
rect 1192 4640 1224 4672
rect 1264 4640 1296 4672
rect 1336 4640 1368 4672
rect 1408 4640 1440 4672
rect 1480 4640 1512 4672
rect 1552 4640 1584 4672
rect 1624 4640 1656 4672
rect 1696 4640 1728 4672
rect 1768 4640 1800 4672
rect 1840 4640 1872 4672
rect 1912 4640 1944 4672
rect 1984 4640 2016 4672
rect 2056 4640 2088 4672
rect 2128 4640 2160 4672
rect 2200 4640 2232 4672
rect 2272 4640 2304 4672
rect 2344 4640 2376 4672
rect 2416 4640 2448 4672
rect 2488 4640 2520 4672
rect 2560 4640 2592 4672
rect 2632 4640 2664 4672
rect 2704 4640 2736 4672
rect 2776 4640 2808 4672
rect 2848 4640 2880 4672
rect 2920 4640 2952 4672
rect 2992 4640 3024 4672
rect 3064 4640 3096 4672
rect 3136 4640 3168 4672
rect 3208 4640 3240 4672
rect 3280 4640 3312 4672
rect 3352 4640 3384 4672
rect 3424 4640 3456 4672
rect 3496 4640 3528 4672
rect 3568 4640 3600 4672
rect 3640 4640 3672 4672
rect 3712 4640 3744 4672
rect 3784 4640 3816 4672
rect 3856 4640 3888 4672
rect 3928 4640 3960 4672
rect 40 4568 72 4600
rect 112 4568 144 4600
rect 184 4568 216 4600
rect 256 4568 288 4600
rect 328 4568 360 4600
rect 400 4568 432 4600
rect 472 4568 504 4600
rect 544 4568 576 4600
rect 616 4568 648 4600
rect 688 4568 720 4600
rect 760 4568 792 4600
rect 832 4568 864 4600
rect 904 4568 936 4600
rect 976 4568 1008 4600
rect 1048 4568 1080 4600
rect 1120 4568 1152 4600
rect 1192 4568 1224 4600
rect 1264 4568 1296 4600
rect 1336 4568 1368 4600
rect 1408 4568 1440 4600
rect 1480 4568 1512 4600
rect 1552 4568 1584 4600
rect 1624 4568 1656 4600
rect 1696 4568 1728 4600
rect 1768 4568 1800 4600
rect 1840 4568 1872 4600
rect 1912 4568 1944 4600
rect 1984 4568 2016 4600
rect 2056 4568 2088 4600
rect 2128 4568 2160 4600
rect 2200 4568 2232 4600
rect 2272 4568 2304 4600
rect 2344 4568 2376 4600
rect 2416 4568 2448 4600
rect 2488 4568 2520 4600
rect 2560 4568 2592 4600
rect 2632 4568 2664 4600
rect 2704 4568 2736 4600
rect 2776 4568 2808 4600
rect 2848 4568 2880 4600
rect 2920 4568 2952 4600
rect 2992 4568 3024 4600
rect 3064 4568 3096 4600
rect 3136 4568 3168 4600
rect 3208 4568 3240 4600
rect 3280 4568 3312 4600
rect 3352 4568 3384 4600
rect 3424 4568 3456 4600
rect 3496 4568 3528 4600
rect 3568 4568 3600 4600
rect 3640 4568 3672 4600
rect 3712 4568 3744 4600
rect 3784 4568 3816 4600
rect 3856 4568 3888 4600
rect 3928 4568 3960 4600
rect 40 4496 72 4528
rect 112 4496 144 4528
rect 184 4496 216 4528
rect 256 4496 288 4528
rect 328 4496 360 4528
rect 400 4496 432 4528
rect 472 4496 504 4528
rect 544 4496 576 4528
rect 616 4496 648 4528
rect 688 4496 720 4528
rect 760 4496 792 4528
rect 832 4496 864 4528
rect 904 4496 936 4528
rect 976 4496 1008 4528
rect 1048 4496 1080 4528
rect 1120 4496 1152 4528
rect 1192 4496 1224 4528
rect 1264 4496 1296 4528
rect 1336 4496 1368 4528
rect 1408 4496 1440 4528
rect 1480 4496 1512 4528
rect 1552 4496 1584 4528
rect 1624 4496 1656 4528
rect 1696 4496 1728 4528
rect 1768 4496 1800 4528
rect 1840 4496 1872 4528
rect 1912 4496 1944 4528
rect 1984 4496 2016 4528
rect 2056 4496 2088 4528
rect 2128 4496 2160 4528
rect 2200 4496 2232 4528
rect 2272 4496 2304 4528
rect 2344 4496 2376 4528
rect 2416 4496 2448 4528
rect 2488 4496 2520 4528
rect 2560 4496 2592 4528
rect 2632 4496 2664 4528
rect 2704 4496 2736 4528
rect 2776 4496 2808 4528
rect 2848 4496 2880 4528
rect 2920 4496 2952 4528
rect 2992 4496 3024 4528
rect 3064 4496 3096 4528
rect 3136 4496 3168 4528
rect 3208 4496 3240 4528
rect 3280 4496 3312 4528
rect 3352 4496 3384 4528
rect 3424 4496 3456 4528
rect 3496 4496 3528 4528
rect 3568 4496 3600 4528
rect 3640 4496 3672 4528
rect 3712 4496 3744 4528
rect 3784 4496 3816 4528
rect 3856 4496 3888 4528
rect 3928 4496 3960 4528
rect 40 4424 72 4456
rect 112 4424 144 4456
rect 184 4424 216 4456
rect 256 4424 288 4456
rect 328 4424 360 4456
rect 400 4424 432 4456
rect 472 4424 504 4456
rect 544 4424 576 4456
rect 616 4424 648 4456
rect 688 4424 720 4456
rect 760 4424 792 4456
rect 832 4424 864 4456
rect 904 4424 936 4456
rect 976 4424 1008 4456
rect 1048 4424 1080 4456
rect 1120 4424 1152 4456
rect 1192 4424 1224 4456
rect 1264 4424 1296 4456
rect 1336 4424 1368 4456
rect 1408 4424 1440 4456
rect 1480 4424 1512 4456
rect 1552 4424 1584 4456
rect 1624 4424 1656 4456
rect 1696 4424 1728 4456
rect 1768 4424 1800 4456
rect 1840 4424 1872 4456
rect 1912 4424 1944 4456
rect 1984 4424 2016 4456
rect 2056 4424 2088 4456
rect 2128 4424 2160 4456
rect 2200 4424 2232 4456
rect 2272 4424 2304 4456
rect 2344 4424 2376 4456
rect 2416 4424 2448 4456
rect 2488 4424 2520 4456
rect 2560 4424 2592 4456
rect 2632 4424 2664 4456
rect 2704 4424 2736 4456
rect 2776 4424 2808 4456
rect 2848 4424 2880 4456
rect 2920 4424 2952 4456
rect 2992 4424 3024 4456
rect 3064 4424 3096 4456
rect 3136 4424 3168 4456
rect 3208 4424 3240 4456
rect 3280 4424 3312 4456
rect 3352 4424 3384 4456
rect 3424 4424 3456 4456
rect 3496 4424 3528 4456
rect 3568 4424 3600 4456
rect 3640 4424 3672 4456
rect 3712 4424 3744 4456
rect 3784 4424 3816 4456
rect 3856 4424 3888 4456
rect 3928 4424 3960 4456
rect 40 4352 72 4384
rect 112 4352 144 4384
rect 184 4352 216 4384
rect 256 4352 288 4384
rect 328 4352 360 4384
rect 400 4352 432 4384
rect 472 4352 504 4384
rect 544 4352 576 4384
rect 616 4352 648 4384
rect 688 4352 720 4384
rect 760 4352 792 4384
rect 832 4352 864 4384
rect 904 4352 936 4384
rect 976 4352 1008 4384
rect 1048 4352 1080 4384
rect 1120 4352 1152 4384
rect 1192 4352 1224 4384
rect 1264 4352 1296 4384
rect 1336 4352 1368 4384
rect 1408 4352 1440 4384
rect 1480 4352 1512 4384
rect 1552 4352 1584 4384
rect 1624 4352 1656 4384
rect 1696 4352 1728 4384
rect 1768 4352 1800 4384
rect 1840 4352 1872 4384
rect 1912 4352 1944 4384
rect 1984 4352 2016 4384
rect 2056 4352 2088 4384
rect 2128 4352 2160 4384
rect 2200 4352 2232 4384
rect 2272 4352 2304 4384
rect 2344 4352 2376 4384
rect 2416 4352 2448 4384
rect 2488 4352 2520 4384
rect 2560 4352 2592 4384
rect 2632 4352 2664 4384
rect 2704 4352 2736 4384
rect 2776 4352 2808 4384
rect 2848 4352 2880 4384
rect 2920 4352 2952 4384
rect 2992 4352 3024 4384
rect 3064 4352 3096 4384
rect 3136 4352 3168 4384
rect 3208 4352 3240 4384
rect 3280 4352 3312 4384
rect 3352 4352 3384 4384
rect 3424 4352 3456 4384
rect 3496 4352 3528 4384
rect 3568 4352 3600 4384
rect 3640 4352 3672 4384
rect 3712 4352 3744 4384
rect 3784 4352 3816 4384
rect 3856 4352 3888 4384
rect 3928 4352 3960 4384
rect 40 4280 72 4312
rect 112 4280 144 4312
rect 184 4280 216 4312
rect 256 4280 288 4312
rect 328 4280 360 4312
rect 400 4280 432 4312
rect 472 4280 504 4312
rect 544 4280 576 4312
rect 616 4280 648 4312
rect 688 4280 720 4312
rect 760 4280 792 4312
rect 832 4280 864 4312
rect 904 4280 936 4312
rect 976 4280 1008 4312
rect 1048 4280 1080 4312
rect 1120 4280 1152 4312
rect 1192 4280 1224 4312
rect 1264 4280 1296 4312
rect 1336 4280 1368 4312
rect 1408 4280 1440 4312
rect 1480 4280 1512 4312
rect 1552 4280 1584 4312
rect 1624 4280 1656 4312
rect 1696 4280 1728 4312
rect 1768 4280 1800 4312
rect 1840 4280 1872 4312
rect 1912 4280 1944 4312
rect 1984 4280 2016 4312
rect 2056 4280 2088 4312
rect 2128 4280 2160 4312
rect 2200 4280 2232 4312
rect 2272 4280 2304 4312
rect 2344 4280 2376 4312
rect 2416 4280 2448 4312
rect 2488 4280 2520 4312
rect 2560 4280 2592 4312
rect 2632 4280 2664 4312
rect 2704 4280 2736 4312
rect 2776 4280 2808 4312
rect 2848 4280 2880 4312
rect 2920 4280 2952 4312
rect 2992 4280 3024 4312
rect 3064 4280 3096 4312
rect 3136 4280 3168 4312
rect 3208 4280 3240 4312
rect 3280 4280 3312 4312
rect 3352 4280 3384 4312
rect 3424 4280 3456 4312
rect 3496 4280 3528 4312
rect 3568 4280 3600 4312
rect 3640 4280 3672 4312
rect 3712 4280 3744 4312
rect 3784 4280 3816 4312
rect 3856 4280 3888 4312
rect 3928 4280 3960 4312
rect 40 4208 72 4240
rect 112 4208 144 4240
rect 184 4208 216 4240
rect 256 4208 288 4240
rect 328 4208 360 4240
rect 400 4208 432 4240
rect 472 4208 504 4240
rect 544 4208 576 4240
rect 616 4208 648 4240
rect 688 4208 720 4240
rect 760 4208 792 4240
rect 832 4208 864 4240
rect 904 4208 936 4240
rect 976 4208 1008 4240
rect 1048 4208 1080 4240
rect 1120 4208 1152 4240
rect 1192 4208 1224 4240
rect 1264 4208 1296 4240
rect 1336 4208 1368 4240
rect 1408 4208 1440 4240
rect 1480 4208 1512 4240
rect 1552 4208 1584 4240
rect 1624 4208 1656 4240
rect 1696 4208 1728 4240
rect 1768 4208 1800 4240
rect 1840 4208 1872 4240
rect 1912 4208 1944 4240
rect 1984 4208 2016 4240
rect 2056 4208 2088 4240
rect 2128 4208 2160 4240
rect 2200 4208 2232 4240
rect 2272 4208 2304 4240
rect 2344 4208 2376 4240
rect 2416 4208 2448 4240
rect 2488 4208 2520 4240
rect 2560 4208 2592 4240
rect 2632 4208 2664 4240
rect 2704 4208 2736 4240
rect 2776 4208 2808 4240
rect 2848 4208 2880 4240
rect 2920 4208 2952 4240
rect 2992 4208 3024 4240
rect 3064 4208 3096 4240
rect 3136 4208 3168 4240
rect 3208 4208 3240 4240
rect 3280 4208 3312 4240
rect 3352 4208 3384 4240
rect 3424 4208 3456 4240
rect 3496 4208 3528 4240
rect 3568 4208 3600 4240
rect 3640 4208 3672 4240
rect 3712 4208 3744 4240
rect 3784 4208 3816 4240
rect 3856 4208 3888 4240
rect 3928 4208 3960 4240
rect 40 4136 72 4168
rect 112 4136 144 4168
rect 184 4136 216 4168
rect 256 4136 288 4168
rect 328 4136 360 4168
rect 400 4136 432 4168
rect 472 4136 504 4168
rect 544 4136 576 4168
rect 616 4136 648 4168
rect 688 4136 720 4168
rect 760 4136 792 4168
rect 832 4136 864 4168
rect 904 4136 936 4168
rect 976 4136 1008 4168
rect 1048 4136 1080 4168
rect 1120 4136 1152 4168
rect 1192 4136 1224 4168
rect 1264 4136 1296 4168
rect 1336 4136 1368 4168
rect 1408 4136 1440 4168
rect 1480 4136 1512 4168
rect 1552 4136 1584 4168
rect 1624 4136 1656 4168
rect 1696 4136 1728 4168
rect 1768 4136 1800 4168
rect 1840 4136 1872 4168
rect 1912 4136 1944 4168
rect 1984 4136 2016 4168
rect 2056 4136 2088 4168
rect 2128 4136 2160 4168
rect 2200 4136 2232 4168
rect 2272 4136 2304 4168
rect 2344 4136 2376 4168
rect 2416 4136 2448 4168
rect 2488 4136 2520 4168
rect 2560 4136 2592 4168
rect 2632 4136 2664 4168
rect 2704 4136 2736 4168
rect 2776 4136 2808 4168
rect 2848 4136 2880 4168
rect 2920 4136 2952 4168
rect 2992 4136 3024 4168
rect 3064 4136 3096 4168
rect 3136 4136 3168 4168
rect 3208 4136 3240 4168
rect 3280 4136 3312 4168
rect 3352 4136 3384 4168
rect 3424 4136 3456 4168
rect 3496 4136 3528 4168
rect 3568 4136 3600 4168
rect 3640 4136 3672 4168
rect 3712 4136 3744 4168
rect 3784 4136 3816 4168
rect 3856 4136 3888 4168
rect 3928 4136 3960 4168
rect 40 4064 72 4096
rect 112 4064 144 4096
rect 184 4064 216 4096
rect 256 4064 288 4096
rect 328 4064 360 4096
rect 400 4064 432 4096
rect 472 4064 504 4096
rect 544 4064 576 4096
rect 616 4064 648 4096
rect 688 4064 720 4096
rect 760 4064 792 4096
rect 832 4064 864 4096
rect 904 4064 936 4096
rect 976 4064 1008 4096
rect 1048 4064 1080 4096
rect 1120 4064 1152 4096
rect 1192 4064 1224 4096
rect 1264 4064 1296 4096
rect 1336 4064 1368 4096
rect 1408 4064 1440 4096
rect 1480 4064 1512 4096
rect 1552 4064 1584 4096
rect 1624 4064 1656 4096
rect 1696 4064 1728 4096
rect 1768 4064 1800 4096
rect 1840 4064 1872 4096
rect 1912 4064 1944 4096
rect 1984 4064 2016 4096
rect 2056 4064 2088 4096
rect 2128 4064 2160 4096
rect 2200 4064 2232 4096
rect 2272 4064 2304 4096
rect 2344 4064 2376 4096
rect 2416 4064 2448 4096
rect 2488 4064 2520 4096
rect 2560 4064 2592 4096
rect 2632 4064 2664 4096
rect 2704 4064 2736 4096
rect 2776 4064 2808 4096
rect 2848 4064 2880 4096
rect 2920 4064 2952 4096
rect 2992 4064 3024 4096
rect 3064 4064 3096 4096
rect 3136 4064 3168 4096
rect 3208 4064 3240 4096
rect 3280 4064 3312 4096
rect 3352 4064 3384 4096
rect 3424 4064 3456 4096
rect 3496 4064 3528 4096
rect 3568 4064 3600 4096
rect 3640 4064 3672 4096
rect 3712 4064 3744 4096
rect 3784 4064 3816 4096
rect 3856 4064 3888 4096
rect 3928 4064 3960 4096
rect 40 3992 72 4024
rect 112 3992 144 4024
rect 184 3992 216 4024
rect 256 3992 288 4024
rect 328 3992 360 4024
rect 400 3992 432 4024
rect 472 3992 504 4024
rect 544 3992 576 4024
rect 616 3992 648 4024
rect 688 3992 720 4024
rect 760 3992 792 4024
rect 832 3992 864 4024
rect 904 3992 936 4024
rect 976 3992 1008 4024
rect 1048 3992 1080 4024
rect 1120 3992 1152 4024
rect 1192 3992 1224 4024
rect 1264 3992 1296 4024
rect 1336 3992 1368 4024
rect 1408 3992 1440 4024
rect 1480 3992 1512 4024
rect 1552 3992 1584 4024
rect 1624 3992 1656 4024
rect 1696 3992 1728 4024
rect 1768 3992 1800 4024
rect 1840 3992 1872 4024
rect 1912 3992 1944 4024
rect 1984 3992 2016 4024
rect 2056 3992 2088 4024
rect 2128 3992 2160 4024
rect 2200 3992 2232 4024
rect 2272 3992 2304 4024
rect 2344 3992 2376 4024
rect 2416 3992 2448 4024
rect 2488 3992 2520 4024
rect 2560 3992 2592 4024
rect 2632 3992 2664 4024
rect 2704 3992 2736 4024
rect 2776 3992 2808 4024
rect 2848 3992 2880 4024
rect 2920 3992 2952 4024
rect 2992 3992 3024 4024
rect 3064 3992 3096 4024
rect 3136 3992 3168 4024
rect 3208 3992 3240 4024
rect 3280 3992 3312 4024
rect 3352 3992 3384 4024
rect 3424 3992 3456 4024
rect 3496 3992 3528 4024
rect 3568 3992 3600 4024
rect 3640 3992 3672 4024
rect 3712 3992 3744 4024
rect 3784 3992 3816 4024
rect 3856 3992 3888 4024
rect 3928 3992 3960 4024
rect 40 3920 72 3952
rect 112 3920 144 3952
rect 184 3920 216 3952
rect 256 3920 288 3952
rect 328 3920 360 3952
rect 400 3920 432 3952
rect 472 3920 504 3952
rect 544 3920 576 3952
rect 616 3920 648 3952
rect 688 3920 720 3952
rect 760 3920 792 3952
rect 832 3920 864 3952
rect 904 3920 936 3952
rect 976 3920 1008 3952
rect 1048 3920 1080 3952
rect 1120 3920 1152 3952
rect 1192 3920 1224 3952
rect 1264 3920 1296 3952
rect 1336 3920 1368 3952
rect 1408 3920 1440 3952
rect 1480 3920 1512 3952
rect 1552 3920 1584 3952
rect 1624 3920 1656 3952
rect 1696 3920 1728 3952
rect 1768 3920 1800 3952
rect 1840 3920 1872 3952
rect 1912 3920 1944 3952
rect 1984 3920 2016 3952
rect 2056 3920 2088 3952
rect 2128 3920 2160 3952
rect 2200 3920 2232 3952
rect 2272 3920 2304 3952
rect 2344 3920 2376 3952
rect 2416 3920 2448 3952
rect 2488 3920 2520 3952
rect 2560 3920 2592 3952
rect 2632 3920 2664 3952
rect 2704 3920 2736 3952
rect 2776 3920 2808 3952
rect 2848 3920 2880 3952
rect 2920 3920 2952 3952
rect 2992 3920 3024 3952
rect 3064 3920 3096 3952
rect 3136 3920 3168 3952
rect 3208 3920 3240 3952
rect 3280 3920 3312 3952
rect 3352 3920 3384 3952
rect 3424 3920 3456 3952
rect 3496 3920 3528 3952
rect 3568 3920 3600 3952
rect 3640 3920 3672 3952
rect 3712 3920 3744 3952
rect 3784 3920 3816 3952
rect 3856 3920 3888 3952
rect 3928 3920 3960 3952
rect 40 3848 72 3880
rect 112 3848 144 3880
rect 184 3848 216 3880
rect 256 3848 288 3880
rect 328 3848 360 3880
rect 400 3848 432 3880
rect 472 3848 504 3880
rect 544 3848 576 3880
rect 616 3848 648 3880
rect 688 3848 720 3880
rect 760 3848 792 3880
rect 832 3848 864 3880
rect 904 3848 936 3880
rect 976 3848 1008 3880
rect 1048 3848 1080 3880
rect 1120 3848 1152 3880
rect 1192 3848 1224 3880
rect 1264 3848 1296 3880
rect 1336 3848 1368 3880
rect 1408 3848 1440 3880
rect 1480 3848 1512 3880
rect 1552 3848 1584 3880
rect 1624 3848 1656 3880
rect 1696 3848 1728 3880
rect 1768 3848 1800 3880
rect 1840 3848 1872 3880
rect 1912 3848 1944 3880
rect 1984 3848 2016 3880
rect 2056 3848 2088 3880
rect 2128 3848 2160 3880
rect 2200 3848 2232 3880
rect 2272 3848 2304 3880
rect 2344 3848 2376 3880
rect 2416 3848 2448 3880
rect 2488 3848 2520 3880
rect 2560 3848 2592 3880
rect 2632 3848 2664 3880
rect 2704 3848 2736 3880
rect 2776 3848 2808 3880
rect 2848 3848 2880 3880
rect 2920 3848 2952 3880
rect 2992 3848 3024 3880
rect 3064 3848 3096 3880
rect 3136 3848 3168 3880
rect 3208 3848 3240 3880
rect 3280 3848 3312 3880
rect 3352 3848 3384 3880
rect 3424 3848 3456 3880
rect 3496 3848 3528 3880
rect 3568 3848 3600 3880
rect 3640 3848 3672 3880
rect 3712 3848 3744 3880
rect 3784 3848 3816 3880
rect 3856 3848 3888 3880
rect 3928 3848 3960 3880
rect 40 3776 72 3808
rect 112 3776 144 3808
rect 184 3776 216 3808
rect 256 3776 288 3808
rect 328 3776 360 3808
rect 400 3776 432 3808
rect 472 3776 504 3808
rect 544 3776 576 3808
rect 616 3776 648 3808
rect 688 3776 720 3808
rect 760 3776 792 3808
rect 832 3776 864 3808
rect 904 3776 936 3808
rect 976 3776 1008 3808
rect 1048 3776 1080 3808
rect 1120 3776 1152 3808
rect 1192 3776 1224 3808
rect 1264 3776 1296 3808
rect 1336 3776 1368 3808
rect 1408 3776 1440 3808
rect 1480 3776 1512 3808
rect 1552 3776 1584 3808
rect 1624 3776 1656 3808
rect 1696 3776 1728 3808
rect 1768 3776 1800 3808
rect 1840 3776 1872 3808
rect 1912 3776 1944 3808
rect 1984 3776 2016 3808
rect 2056 3776 2088 3808
rect 2128 3776 2160 3808
rect 2200 3776 2232 3808
rect 2272 3776 2304 3808
rect 2344 3776 2376 3808
rect 2416 3776 2448 3808
rect 2488 3776 2520 3808
rect 2560 3776 2592 3808
rect 2632 3776 2664 3808
rect 2704 3776 2736 3808
rect 2776 3776 2808 3808
rect 2848 3776 2880 3808
rect 2920 3776 2952 3808
rect 2992 3776 3024 3808
rect 3064 3776 3096 3808
rect 3136 3776 3168 3808
rect 3208 3776 3240 3808
rect 3280 3776 3312 3808
rect 3352 3776 3384 3808
rect 3424 3776 3456 3808
rect 3496 3776 3528 3808
rect 3568 3776 3600 3808
rect 3640 3776 3672 3808
rect 3712 3776 3744 3808
rect 3784 3776 3816 3808
rect 3856 3776 3888 3808
rect 3928 3776 3960 3808
rect 40 3704 72 3736
rect 112 3704 144 3736
rect 184 3704 216 3736
rect 256 3704 288 3736
rect 328 3704 360 3736
rect 400 3704 432 3736
rect 472 3704 504 3736
rect 544 3704 576 3736
rect 616 3704 648 3736
rect 688 3704 720 3736
rect 760 3704 792 3736
rect 832 3704 864 3736
rect 904 3704 936 3736
rect 976 3704 1008 3736
rect 1048 3704 1080 3736
rect 1120 3704 1152 3736
rect 1192 3704 1224 3736
rect 1264 3704 1296 3736
rect 1336 3704 1368 3736
rect 1408 3704 1440 3736
rect 1480 3704 1512 3736
rect 1552 3704 1584 3736
rect 1624 3704 1656 3736
rect 1696 3704 1728 3736
rect 1768 3704 1800 3736
rect 1840 3704 1872 3736
rect 1912 3704 1944 3736
rect 1984 3704 2016 3736
rect 2056 3704 2088 3736
rect 2128 3704 2160 3736
rect 2200 3704 2232 3736
rect 2272 3704 2304 3736
rect 2344 3704 2376 3736
rect 2416 3704 2448 3736
rect 2488 3704 2520 3736
rect 2560 3704 2592 3736
rect 2632 3704 2664 3736
rect 2704 3704 2736 3736
rect 2776 3704 2808 3736
rect 2848 3704 2880 3736
rect 2920 3704 2952 3736
rect 2992 3704 3024 3736
rect 3064 3704 3096 3736
rect 3136 3704 3168 3736
rect 3208 3704 3240 3736
rect 3280 3704 3312 3736
rect 3352 3704 3384 3736
rect 3424 3704 3456 3736
rect 3496 3704 3528 3736
rect 3568 3704 3600 3736
rect 3640 3704 3672 3736
rect 3712 3704 3744 3736
rect 3784 3704 3816 3736
rect 3856 3704 3888 3736
rect 3928 3704 3960 3736
rect 40 3632 72 3664
rect 112 3632 144 3664
rect 184 3632 216 3664
rect 256 3632 288 3664
rect 328 3632 360 3664
rect 400 3632 432 3664
rect 472 3632 504 3664
rect 544 3632 576 3664
rect 616 3632 648 3664
rect 688 3632 720 3664
rect 760 3632 792 3664
rect 832 3632 864 3664
rect 904 3632 936 3664
rect 976 3632 1008 3664
rect 1048 3632 1080 3664
rect 1120 3632 1152 3664
rect 1192 3632 1224 3664
rect 1264 3632 1296 3664
rect 1336 3632 1368 3664
rect 1408 3632 1440 3664
rect 1480 3632 1512 3664
rect 1552 3632 1584 3664
rect 1624 3632 1656 3664
rect 1696 3632 1728 3664
rect 1768 3632 1800 3664
rect 1840 3632 1872 3664
rect 1912 3632 1944 3664
rect 1984 3632 2016 3664
rect 2056 3632 2088 3664
rect 2128 3632 2160 3664
rect 2200 3632 2232 3664
rect 2272 3632 2304 3664
rect 2344 3632 2376 3664
rect 2416 3632 2448 3664
rect 2488 3632 2520 3664
rect 2560 3632 2592 3664
rect 2632 3632 2664 3664
rect 2704 3632 2736 3664
rect 2776 3632 2808 3664
rect 2848 3632 2880 3664
rect 2920 3632 2952 3664
rect 2992 3632 3024 3664
rect 3064 3632 3096 3664
rect 3136 3632 3168 3664
rect 3208 3632 3240 3664
rect 3280 3632 3312 3664
rect 3352 3632 3384 3664
rect 3424 3632 3456 3664
rect 3496 3632 3528 3664
rect 3568 3632 3600 3664
rect 3640 3632 3672 3664
rect 3712 3632 3744 3664
rect 3784 3632 3816 3664
rect 3856 3632 3888 3664
rect 3928 3632 3960 3664
rect 40 3560 72 3592
rect 112 3560 144 3592
rect 184 3560 216 3592
rect 256 3560 288 3592
rect 328 3560 360 3592
rect 400 3560 432 3592
rect 472 3560 504 3592
rect 544 3560 576 3592
rect 616 3560 648 3592
rect 688 3560 720 3592
rect 760 3560 792 3592
rect 832 3560 864 3592
rect 904 3560 936 3592
rect 976 3560 1008 3592
rect 1048 3560 1080 3592
rect 1120 3560 1152 3592
rect 1192 3560 1224 3592
rect 1264 3560 1296 3592
rect 1336 3560 1368 3592
rect 1408 3560 1440 3592
rect 1480 3560 1512 3592
rect 1552 3560 1584 3592
rect 1624 3560 1656 3592
rect 1696 3560 1728 3592
rect 1768 3560 1800 3592
rect 1840 3560 1872 3592
rect 1912 3560 1944 3592
rect 1984 3560 2016 3592
rect 2056 3560 2088 3592
rect 2128 3560 2160 3592
rect 2200 3560 2232 3592
rect 2272 3560 2304 3592
rect 2344 3560 2376 3592
rect 2416 3560 2448 3592
rect 2488 3560 2520 3592
rect 2560 3560 2592 3592
rect 2632 3560 2664 3592
rect 2704 3560 2736 3592
rect 2776 3560 2808 3592
rect 2848 3560 2880 3592
rect 2920 3560 2952 3592
rect 2992 3560 3024 3592
rect 3064 3560 3096 3592
rect 3136 3560 3168 3592
rect 3208 3560 3240 3592
rect 3280 3560 3312 3592
rect 3352 3560 3384 3592
rect 3424 3560 3456 3592
rect 3496 3560 3528 3592
rect 3568 3560 3600 3592
rect 3640 3560 3672 3592
rect 3712 3560 3744 3592
rect 3784 3560 3816 3592
rect 3856 3560 3888 3592
rect 3928 3560 3960 3592
rect 40 3488 72 3520
rect 112 3488 144 3520
rect 184 3488 216 3520
rect 256 3488 288 3520
rect 328 3488 360 3520
rect 400 3488 432 3520
rect 472 3488 504 3520
rect 544 3488 576 3520
rect 616 3488 648 3520
rect 688 3488 720 3520
rect 760 3488 792 3520
rect 832 3488 864 3520
rect 904 3488 936 3520
rect 976 3488 1008 3520
rect 1048 3488 1080 3520
rect 1120 3488 1152 3520
rect 1192 3488 1224 3520
rect 1264 3488 1296 3520
rect 1336 3488 1368 3520
rect 1408 3488 1440 3520
rect 1480 3488 1512 3520
rect 1552 3488 1584 3520
rect 1624 3488 1656 3520
rect 1696 3488 1728 3520
rect 1768 3488 1800 3520
rect 1840 3488 1872 3520
rect 1912 3488 1944 3520
rect 1984 3488 2016 3520
rect 2056 3488 2088 3520
rect 2128 3488 2160 3520
rect 2200 3488 2232 3520
rect 2272 3488 2304 3520
rect 2344 3488 2376 3520
rect 2416 3488 2448 3520
rect 2488 3488 2520 3520
rect 2560 3488 2592 3520
rect 2632 3488 2664 3520
rect 2704 3488 2736 3520
rect 2776 3488 2808 3520
rect 2848 3488 2880 3520
rect 2920 3488 2952 3520
rect 2992 3488 3024 3520
rect 3064 3488 3096 3520
rect 3136 3488 3168 3520
rect 3208 3488 3240 3520
rect 3280 3488 3312 3520
rect 3352 3488 3384 3520
rect 3424 3488 3456 3520
rect 3496 3488 3528 3520
rect 3568 3488 3600 3520
rect 3640 3488 3672 3520
rect 3712 3488 3744 3520
rect 3784 3488 3816 3520
rect 3856 3488 3888 3520
rect 3928 3488 3960 3520
rect 40 3416 72 3448
rect 112 3416 144 3448
rect 184 3416 216 3448
rect 256 3416 288 3448
rect 328 3416 360 3448
rect 400 3416 432 3448
rect 472 3416 504 3448
rect 544 3416 576 3448
rect 616 3416 648 3448
rect 688 3416 720 3448
rect 760 3416 792 3448
rect 832 3416 864 3448
rect 904 3416 936 3448
rect 976 3416 1008 3448
rect 1048 3416 1080 3448
rect 1120 3416 1152 3448
rect 1192 3416 1224 3448
rect 1264 3416 1296 3448
rect 1336 3416 1368 3448
rect 1408 3416 1440 3448
rect 1480 3416 1512 3448
rect 1552 3416 1584 3448
rect 1624 3416 1656 3448
rect 1696 3416 1728 3448
rect 1768 3416 1800 3448
rect 1840 3416 1872 3448
rect 1912 3416 1944 3448
rect 1984 3416 2016 3448
rect 2056 3416 2088 3448
rect 2128 3416 2160 3448
rect 2200 3416 2232 3448
rect 2272 3416 2304 3448
rect 2344 3416 2376 3448
rect 2416 3416 2448 3448
rect 2488 3416 2520 3448
rect 2560 3416 2592 3448
rect 2632 3416 2664 3448
rect 2704 3416 2736 3448
rect 2776 3416 2808 3448
rect 2848 3416 2880 3448
rect 2920 3416 2952 3448
rect 2992 3416 3024 3448
rect 3064 3416 3096 3448
rect 3136 3416 3168 3448
rect 3208 3416 3240 3448
rect 3280 3416 3312 3448
rect 3352 3416 3384 3448
rect 3424 3416 3456 3448
rect 3496 3416 3528 3448
rect 3568 3416 3600 3448
rect 3640 3416 3672 3448
rect 3712 3416 3744 3448
rect 3784 3416 3816 3448
rect 3856 3416 3888 3448
rect 3928 3416 3960 3448
rect 40 3344 72 3376
rect 112 3344 144 3376
rect 184 3344 216 3376
rect 256 3344 288 3376
rect 328 3344 360 3376
rect 400 3344 432 3376
rect 472 3344 504 3376
rect 544 3344 576 3376
rect 616 3344 648 3376
rect 688 3344 720 3376
rect 760 3344 792 3376
rect 832 3344 864 3376
rect 904 3344 936 3376
rect 976 3344 1008 3376
rect 1048 3344 1080 3376
rect 1120 3344 1152 3376
rect 1192 3344 1224 3376
rect 1264 3344 1296 3376
rect 1336 3344 1368 3376
rect 1408 3344 1440 3376
rect 1480 3344 1512 3376
rect 1552 3344 1584 3376
rect 1624 3344 1656 3376
rect 1696 3344 1728 3376
rect 1768 3344 1800 3376
rect 1840 3344 1872 3376
rect 1912 3344 1944 3376
rect 1984 3344 2016 3376
rect 2056 3344 2088 3376
rect 2128 3344 2160 3376
rect 2200 3344 2232 3376
rect 2272 3344 2304 3376
rect 2344 3344 2376 3376
rect 2416 3344 2448 3376
rect 2488 3344 2520 3376
rect 2560 3344 2592 3376
rect 2632 3344 2664 3376
rect 2704 3344 2736 3376
rect 2776 3344 2808 3376
rect 2848 3344 2880 3376
rect 2920 3344 2952 3376
rect 2992 3344 3024 3376
rect 3064 3344 3096 3376
rect 3136 3344 3168 3376
rect 3208 3344 3240 3376
rect 3280 3344 3312 3376
rect 3352 3344 3384 3376
rect 3424 3344 3456 3376
rect 3496 3344 3528 3376
rect 3568 3344 3600 3376
rect 3640 3344 3672 3376
rect 3712 3344 3744 3376
rect 3784 3344 3816 3376
rect 3856 3344 3888 3376
rect 3928 3344 3960 3376
rect 40 3272 72 3304
rect 112 3272 144 3304
rect 184 3272 216 3304
rect 256 3272 288 3304
rect 328 3272 360 3304
rect 400 3272 432 3304
rect 472 3272 504 3304
rect 544 3272 576 3304
rect 616 3272 648 3304
rect 688 3272 720 3304
rect 760 3272 792 3304
rect 832 3272 864 3304
rect 904 3272 936 3304
rect 976 3272 1008 3304
rect 1048 3272 1080 3304
rect 1120 3272 1152 3304
rect 1192 3272 1224 3304
rect 1264 3272 1296 3304
rect 1336 3272 1368 3304
rect 1408 3272 1440 3304
rect 1480 3272 1512 3304
rect 1552 3272 1584 3304
rect 1624 3272 1656 3304
rect 1696 3272 1728 3304
rect 1768 3272 1800 3304
rect 1840 3272 1872 3304
rect 1912 3272 1944 3304
rect 1984 3272 2016 3304
rect 2056 3272 2088 3304
rect 2128 3272 2160 3304
rect 2200 3272 2232 3304
rect 2272 3272 2304 3304
rect 2344 3272 2376 3304
rect 2416 3272 2448 3304
rect 2488 3272 2520 3304
rect 2560 3272 2592 3304
rect 2632 3272 2664 3304
rect 2704 3272 2736 3304
rect 2776 3272 2808 3304
rect 2848 3272 2880 3304
rect 2920 3272 2952 3304
rect 2992 3272 3024 3304
rect 3064 3272 3096 3304
rect 3136 3272 3168 3304
rect 3208 3272 3240 3304
rect 3280 3272 3312 3304
rect 3352 3272 3384 3304
rect 3424 3272 3456 3304
rect 3496 3272 3528 3304
rect 3568 3272 3600 3304
rect 3640 3272 3672 3304
rect 3712 3272 3744 3304
rect 3784 3272 3816 3304
rect 3856 3272 3888 3304
rect 3928 3272 3960 3304
rect 40 3200 72 3232
rect 112 3200 144 3232
rect 184 3200 216 3232
rect 256 3200 288 3232
rect 328 3200 360 3232
rect 400 3200 432 3232
rect 472 3200 504 3232
rect 544 3200 576 3232
rect 616 3200 648 3232
rect 688 3200 720 3232
rect 760 3200 792 3232
rect 832 3200 864 3232
rect 904 3200 936 3232
rect 976 3200 1008 3232
rect 1048 3200 1080 3232
rect 1120 3200 1152 3232
rect 1192 3200 1224 3232
rect 1264 3200 1296 3232
rect 1336 3200 1368 3232
rect 1408 3200 1440 3232
rect 1480 3200 1512 3232
rect 1552 3200 1584 3232
rect 1624 3200 1656 3232
rect 1696 3200 1728 3232
rect 1768 3200 1800 3232
rect 1840 3200 1872 3232
rect 1912 3200 1944 3232
rect 1984 3200 2016 3232
rect 2056 3200 2088 3232
rect 2128 3200 2160 3232
rect 2200 3200 2232 3232
rect 2272 3200 2304 3232
rect 2344 3200 2376 3232
rect 2416 3200 2448 3232
rect 2488 3200 2520 3232
rect 2560 3200 2592 3232
rect 2632 3200 2664 3232
rect 2704 3200 2736 3232
rect 2776 3200 2808 3232
rect 2848 3200 2880 3232
rect 2920 3200 2952 3232
rect 2992 3200 3024 3232
rect 3064 3200 3096 3232
rect 3136 3200 3168 3232
rect 3208 3200 3240 3232
rect 3280 3200 3312 3232
rect 3352 3200 3384 3232
rect 3424 3200 3456 3232
rect 3496 3200 3528 3232
rect 3568 3200 3600 3232
rect 3640 3200 3672 3232
rect 3712 3200 3744 3232
rect 3784 3200 3816 3232
rect 3856 3200 3888 3232
rect 3928 3200 3960 3232
rect 40 3128 72 3160
rect 112 3128 144 3160
rect 184 3128 216 3160
rect 256 3128 288 3160
rect 328 3128 360 3160
rect 400 3128 432 3160
rect 472 3128 504 3160
rect 544 3128 576 3160
rect 616 3128 648 3160
rect 688 3128 720 3160
rect 760 3128 792 3160
rect 832 3128 864 3160
rect 904 3128 936 3160
rect 976 3128 1008 3160
rect 1048 3128 1080 3160
rect 1120 3128 1152 3160
rect 1192 3128 1224 3160
rect 1264 3128 1296 3160
rect 1336 3128 1368 3160
rect 1408 3128 1440 3160
rect 1480 3128 1512 3160
rect 1552 3128 1584 3160
rect 1624 3128 1656 3160
rect 1696 3128 1728 3160
rect 1768 3128 1800 3160
rect 1840 3128 1872 3160
rect 1912 3128 1944 3160
rect 1984 3128 2016 3160
rect 2056 3128 2088 3160
rect 2128 3128 2160 3160
rect 2200 3128 2232 3160
rect 2272 3128 2304 3160
rect 2344 3128 2376 3160
rect 2416 3128 2448 3160
rect 2488 3128 2520 3160
rect 2560 3128 2592 3160
rect 2632 3128 2664 3160
rect 2704 3128 2736 3160
rect 2776 3128 2808 3160
rect 2848 3128 2880 3160
rect 2920 3128 2952 3160
rect 2992 3128 3024 3160
rect 3064 3128 3096 3160
rect 3136 3128 3168 3160
rect 3208 3128 3240 3160
rect 3280 3128 3312 3160
rect 3352 3128 3384 3160
rect 3424 3128 3456 3160
rect 3496 3128 3528 3160
rect 3568 3128 3600 3160
rect 3640 3128 3672 3160
rect 3712 3128 3744 3160
rect 3784 3128 3816 3160
rect 3856 3128 3888 3160
rect 3928 3128 3960 3160
rect 40 3056 72 3088
rect 112 3056 144 3088
rect 184 3056 216 3088
rect 256 3056 288 3088
rect 328 3056 360 3088
rect 400 3056 432 3088
rect 472 3056 504 3088
rect 544 3056 576 3088
rect 616 3056 648 3088
rect 688 3056 720 3088
rect 760 3056 792 3088
rect 832 3056 864 3088
rect 904 3056 936 3088
rect 976 3056 1008 3088
rect 1048 3056 1080 3088
rect 1120 3056 1152 3088
rect 1192 3056 1224 3088
rect 1264 3056 1296 3088
rect 1336 3056 1368 3088
rect 1408 3056 1440 3088
rect 1480 3056 1512 3088
rect 1552 3056 1584 3088
rect 1624 3056 1656 3088
rect 1696 3056 1728 3088
rect 1768 3056 1800 3088
rect 1840 3056 1872 3088
rect 1912 3056 1944 3088
rect 1984 3056 2016 3088
rect 2056 3056 2088 3088
rect 2128 3056 2160 3088
rect 2200 3056 2232 3088
rect 2272 3056 2304 3088
rect 2344 3056 2376 3088
rect 2416 3056 2448 3088
rect 2488 3056 2520 3088
rect 2560 3056 2592 3088
rect 2632 3056 2664 3088
rect 2704 3056 2736 3088
rect 2776 3056 2808 3088
rect 2848 3056 2880 3088
rect 2920 3056 2952 3088
rect 2992 3056 3024 3088
rect 3064 3056 3096 3088
rect 3136 3056 3168 3088
rect 3208 3056 3240 3088
rect 3280 3056 3312 3088
rect 3352 3056 3384 3088
rect 3424 3056 3456 3088
rect 3496 3056 3528 3088
rect 3568 3056 3600 3088
rect 3640 3056 3672 3088
rect 3712 3056 3744 3088
rect 3784 3056 3816 3088
rect 3856 3056 3888 3088
rect 3928 3056 3960 3088
rect 40 2984 72 3016
rect 112 2984 144 3016
rect 184 2984 216 3016
rect 256 2984 288 3016
rect 328 2984 360 3016
rect 400 2984 432 3016
rect 472 2984 504 3016
rect 544 2984 576 3016
rect 616 2984 648 3016
rect 688 2984 720 3016
rect 760 2984 792 3016
rect 832 2984 864 3016
rect 904 2984 936 3016
rect 976 2984 1008 3016
rect 1048 2984 1080 3016
rect 1120 2984 1152 3016
rect 1192 2984 1224 3016
rect 1264 2984 1296 3016
rect 1336 2984 1368 3016
rect 1408 2984 1440 3016
rect 1480 2984 1512 3016
rect 1552 2984 1584 3016
rect 1624 2984 1656 3016
rect 1696 2984 1728 3016
rect 1768 2984 1800 3016
rect 1840 2984 1872 3016
rect 1912 2984 1944 3016
rect 1984 2984 2016 3016
rect 2056 2984 2088 3016
rect 2128 2984 2160 3016
rect 2200 2984 2232 3016
rect 2272 2984 2304 3016
rect 2344 2984 2376 3016
rect 2416 2984 2448 3016
rect 2488 2984 2520 3016
rect 2560 2984 2592 3016
rect 2632 2984 2664 3016
rect 2704 2984 2736 3016
rect 2776 2984 2808 3016
rect 2848 2984 2880 3016
rect 2920 2984 2952 3016
rect 2992 2984 3024 3016
rect 3064 2984 3096 3016
rect 3136 2984 3168 3016
rect 3208 2984 3240 3016
rect 3280 2984 3312 3016
rect 3352 2984 3384 3016
rect 3424 2984 3456 3016
rect 3496 2984 3528 3016
rect 3568 2984 3600 3016
rect 3640 2984 3672 3016
rect 3712 2984 3744 3016
rect 3784 2984 3816 3016
rect 3856 2984 3888 3016
rect 3928 2984 3960 3016
rect 40 2912 72 2944
rect 112 2912 144 2944
rect 184 2912 216 2944
rect 256 2912 288 2944
rect 328 2912 360 2944
rect 400 2912 432 2944
rect 472 2912 504 2944
rect 544 2912 576 2944
rect 616 2912 648 2944
rect 688 2912 720 2944
rect 760 2912 792 2944
rect 832 2912 864 2944
rect 904 2912 936 2944
rect 976 2912 1008 2944
rect 1048 2912 1080 2944
rect 1120 2912 1152 2944
rect 1192 2912 1224 2944
rect 1264 2912 1296 2944
rect 1336 2912 1368 2944
rect 1408 2912 1440 2944
rect 1480 2912 1512 2944
rect 1552 2912 1584 2944
rect 1624 2912 1656 2944
rect 1696 2912 1728 2944
rect 1768 2912 1800 2944
rect 1840 2912 1872 2944
rect 1912 2912 1944 2944
rect 1984 2912 2016 2944
rect 2056 2912 2088 2944
rect 2128 2912 2160 2944
rect 2200 2912 2232 2944
rect 2272 2912 2304 2944
rect 2344 2912 2376 2944
rect 2416 2912 2448 2944
rect 2488 2912 2520 2944
rect 2560 2912 2592 2944
rect 2632 2912 2664 2944
rect 2704 2912 2736 2944
rect 2776 2912 2808 2944
rect 2848 2912 2880 2944
rect 2920 2912 2952 2944
rect 2992 2912 3024 2944
rect 3064 2912 3096 2944
rect 3136 2912 3168 2944
rect 3208 2912 3240 2944
rect 3280 2912 3312 2944
rect 3352 2912 3384 2944
rect 3424 2912 3456 2944
rect 3496 2912 3528 2944
rect 3568 2912 3600 2944
rect 3640 2912 3672 2944
rect 3712 2912 3744 2944
rect 3784 2912 3816 2944
rect 3856 2912 3888 2944
rect 3928 2912 3960 2944
rect 40 2840 72 2872
rect 112 2840 144 2872
rect 184 2840 216 2872
rect 256 2840 288 2872
rect 328 2840 360 2872
rect 400 2840 432 2872
rect 472 2840 504 2872
rect 544 2840 576 2872
rect 616 2840 648 2872
rect 688 2840 720 2872
rect 760 2840 792 2872
rect 832 2840 864 2872
rect 904 2840 936 2872
rect 976 2840 1008 2872
rect 1048 2840 1080 2872
rect 1120 2840 1152 2872
rect 1192 2840 1224 2872
rect 1264 2840 1296 2872
rect 1336 2840 1368 2872
rect 1408 2840 1440 2872
rect 1480 2840 1512 2872
rect 1552 2840 1584 2872
rect 1624 2840 1656 2872
rect 1696 2840 1728 2872
rect 1768 2840 1800 2872
rect 1840 2840 1872 2872
rect 1912 2840 1944 2872
rect 1984 2840 2016 2872
rect 2056 2840 2088 2872
rect 2128 2840 2160 2872
rect 2200 2840 2232 2872
rect 2272 2840 2304 2872
rect 2344 2840 2376 2872
rect 2416 2840 2448 2872
rect 2488 2840 2520 2872
rect 2560 2840 2592 2872
rect 2632 2840 2664 2872
rect 2704 2840 2736 2872
rect 2776 2840 2808 2872
rect 2848 2840 2880 2872
rect 2920 2840 2952 2872
rect 2992 2840 3024 2872
rect 3064 2840 3096 2872
rect 3136 2840 3168 2872
rect 3208 2840 3240 2872
rect 3280 2840 3312 2872
rect 3352 2840 3384 2872
rect 3424 2840 3456 2872
rect 3496 2840 3528 2872
rect 3568 2840 3600 2872
rect 3640 2840 3672 2872
rect 3712 2840 3744 2872
rect 3784 2840 3816 2872
rect 3856 2840 3888 2872
rect 3928 2840 3960 2872
rect 40 2768 72 2800
rect 112 2768 144 2800
rect 184 2768 216 2800
rect 256 2768 288 2800
rect 328 2768 360 2800
rect 400 2768 432 2800
rect 472 2768 504 2800
rect 544 2768 576 2800
rect 616 2768 648 2800
rect 688 2768 720 2800
rect 760 2768 792 2800
rect 832 2768 864 2800
rect 904 2768 936 2800
rect 976 2768 1008 2800
rect 1048 2768 1080 2800
rect 1120 2768 1152 2800
rect 1192 2768 1224 2800
rect 1264 2768 1296 2800
rect 1336 2768 1368 2800
rect 1408 2768 1440 2800
rect 1480 2768 1512 2800
rect 1552 2768 1584 2800
rect 1624 2768 1656 2800
rect 1696 2768 1728 2800
rect 1768 2768 1800 2800
rect 1840 2768 1872 2800
rect 1912 2768 1944 2800
rect 1984 2768 2016 2800
rect 2056 2768 2088 2800
rect 2128 2768 2160 2800
rect 2200 2768 2232 2800
rect 2272 2768 2304 2800
rect 2344 2768 2376 2800
rect 2416 2768 2448 2800
rect 2488 2768 2520 2800
rect 2560 2768 2592 2800
rect 2632 2768 2664 2800
rect 2704 2768 2736 2800
rect 2776 2768 2808 2800
rect 2848 2768 2880 2800
rect 2920 2768 2952 2800
rect 2992 2768 3024 2800
rect 3064 2768 3096 2800
rect 3136 2768 3168 2800
rect 3208 2768 3240 2800
rect 3280 2768 3312 2800
rect 3352 2768 3384 2800
rect 3424 2768 3456 2800
rect 3496 2768 3528 2800
rect 3568 2768 3600 2800
rect 3640 2768 3672 2800
rect 3712 2768 3744 2800
rect 3784 2768 3816 2800
rect 3856 2768 3888 2800
rect 3928 2768 3960 2800
rect 40 2696 72 2728
rect 112 2696 144 2728
rect 184 2696 216 2728
rect 256 2696 288 2728
rect 328 2696 360 2728
rect 400 2696 432 2728
rect 472 2696 504 2728
rect 544 2696 576 2728
rect 616 2696 648 2728
rect 688 2696 720 2728
rect 760 2696 792 2728
rect 832 2696 864 2728
rect 904 2696 936 2728
rect 976 2696 1008 2728
rect 1048 2696 1080 2728
rect 1120 2696 1152 2728
rect 1192 2696 1224 2728
rect 1264 2696 1296 2728
rect 1336 2696 1368 2728
rect 1408 2696 1440 2728
rect 1480 2696 1512 2728
rect 1552 2696 1584 2728
rect 1624 2696 1656 2728
rect 1696 2696 1728 2728
rect 1768 2696 1800 2728
rect 1840 2696 1872 2728
rect 1912 2696 1944 2728
rect 1984 2696 2016 2728
rect 2056 2696 2088 2728
rect 2128 2696 2160 2728
rect 2200 2696 2232 2728
rect 2272 2696 2304 2728
rect 2344 2696 2376 2728
rect 2416 2696 2448 2728
rect 2488 2696 2520 2728
rect 2560 2696 2592 2728
rect 2632 2696 2664 2728
rect 2704 2696 2736 2728
rect 2776 2696 2808 2728
rect 2848 2696 2880 2728
rect 2920 2696 2952 2728
rect 2992 2696 3024 2728
rect 3064 2696 3096 2728
rect 3136 2696 3168 2728
rect 3208 2696 3240 2728
rect 3280 2696 3312 2728
rect 3352 2696 3384 2728
rect 3424 2696 3456 2728
rect 3496 2696 3528 2728
rect 3568 2696 3600 2728
rect 3640 2696 3672 2728
rect 3712 2696 3744 2728
rect 3784 2696 3816 2728
rect 3856 2696 3888 2728
rect 3928 2696 3960 2728
rect 40 2624 72 2656
rect 112 2624 144 2656
rect 184 2624 216 2656
rect 256 2624 288 2656
rect 328 2624 360 2656
rect 400 2624 432 2656
rect 472 2624 504 2656
rect 544 2624 576 2656
rect 616 2624 648 2656
rect 688 2624 720 2656
rect 760 2624 792 2656
rect 832 2624 864 2656
rect 904 2624 936 2656
rect 976 2624 1008 2656
rect 1048 2624 1080 2656
rect 1120 2624 1152 2656
rect 1192 2624 1224 2656
rect 1264 2624 1296 2656
rect 1336 2624 1368 2656
rect 1408 2624 1440 2656
rect 1480 2624 1512 2656
rect 1552 2624 1584 2656
rect 1624 2624 1656 2656
rect 1696 2624 1728 2656
rect 1768 2624 1800 2656
rect 1840 2624 1872 2656
rect 1912 2624 1944 2656
rect 1984 2624 2016 2656
rect 2056 2624 2088 2656
rect 2128 2624 2160 2656
rect 2200 2624 2232 2656
rect 2272 2624 2304 2656
rect 2344 2624 2376 2656
rect 2416 2624 2448 2656
rect 2488 2624 2520 2656
rect 2560 2624 2592 2656
rect 2632 2624 2664 2656
rect 2704 2624 2736 2656
rect 2776 2624 2808 2656
rect 2848 2624 2880 2656
rect 2920 2624 2952 2656
rect 2992 2624 3024 2656
rect 3064 2624 3096 2656
rect 3136 2624 3168 2656
rect 3208 2624 3240 2656
rect 3280 2624 3312 2656
rect 3352 2624 3384 2656
rect 3424 2624 3456 2656
rect 3496 2624 3528 2656
rect 3568 2624 3600 2656
rect 3640 2624 3672 2656
rect 3712 2624 3744 2656
rect 3784 2624 3816 2656
rect 3856 2624 3888 2656
rect 3928 2624 3960 2656
rect 40 2552 72 2584
rect 112 2552 144 2584
rect 184 2552 216 2584
rect 256 2552 288 2584
rect 328 2552 360 2584
rect 400 2552 432 2584
rect 472 2552 504 2584
rect 544 2552 576 2584
rect 616 2552 648 2584
rect 688 2552 720 2584
rect 760 2552 792 2584
rect 832 2552 864 2584
rect 904 2552 936 2584
rect 976 2552 1008 2584
rect 1048 2552 1080 2584
rect 1120 2552 1152 2584
rect 1192 2552 1224 2584
rect 1264 2552 1296 2584
rect 1336 2552 1368 2584
rect 1408 2552 1440 2584
rect 1480 2552 1512 2584
rect 1552 2552 1584 2584
rect 1624 2552 1656 2584
rect 1696 2552 1728 2584
rect 1768 2552 1800 2584
rect 1840 2552 1872 2584
rect 1912 2552 1944 2584
rect 1984 2552 2016 2584
rect 2056 2552 2088 2584
rect 2128 2552 2160 2584
rect 2200 2552 2232 2584
rect 2272 2552 2304 2584
rect 2344 2552 2376 2584
rect 2416 2552 2448 2584
rect 2488 2552 2520 2584
rect 2560 2552 2592 2584
rect 2632 2552 2664 2584
rect 2704 2552 2736 2584
rect 2776 2552 2808 2584
rect 2848 2552 2880 2584
rect 2920 2552 2952 2584
rect 2992 2552 3024 2584
rect 3064 2552 3096 2584
rect 3136 2552 3168 2584
rect 3208 2552 3240 2584
rect 3280 2552 3312 2584
rect 3352 2552 3384 2584
rect 3424 2552 3456 2584
rect 3496 2552 3528 2584
rect 3568 2552 3600 2584
rect 3640 2552 3672 2584
rect 3712 2552 3744 2584
rect 3784 2552 3816 2584
rect 3856 2552 3888 2584
rect 3928 2552 3960 2584
rect 40 2480 72 2512
rect 112 2480 144 2512
rect 184 2480 216 2512
rect 256 2480 288 2512
rect 328 2480 360 2512
rect 400 2480 432 2512
rect 472 2480 504 2512
rect 544 2480 576 2512
rect 616 2480 648 2512
rect 688 2480 720 2512
rect 760 2480 792 2512
rect 832 2480 864 2512
rect 904 2480 936 2512
rect 976 2480 1008 2512
rect 1048 2480 1080 2512
rect 1120 2480 1152 2512
rect 1192 2480 1224 2512
rect 1264 2480 1296 2512
rect 1336 2480 1368 2512
rect 1408 2480 1440 2512
rect 1480 2480 1512 2512
rect 1552 2480 1584 2512
rect 1624 2480 1656 2512
rect 1696 2480 1728 2512
rect 1768 2480 1800 2512
rect 1840 2480 1872 2512
rect 1912 2480 1944 2512
rect 1984 2480 2016 2512
rect 2056 2480 2088 2512
rect 2128 2480 2160 2512
rect 2200 2480 2232 2512
rect 2272 2480 2304 2512
rect 2344 2480 2376 2512
rect 2416 2480 2448 2512
rect 2488 2480 2520 2512
rect 2560 2480 2592 2512
rect 2632 2480 2664 2512
rect 2704 2480 2736 2512
rect 2776 2480 2808 2512
rect 2848 2480 2880 2512
rect 2920 2480 2952 2512
rect 2992 2480 3024 2512
rect 3064 2480 3096 2512
rect 3136 2480 3168 2512
rect 3208 2480 3240 2512
rect 3280 2480 3312 2512
rect 3352 2480 3384 2512
rect 3424 2480 3456 2512
rect 3496 2480 3528 2512
rect 3568 2480 3600 2512
rect 3640 2480 3672 2512
rect 3712 2480 3744 2512
rect 3784 2480 3816 2512
rect 3856 2480 3888 2512
rect 3928 2480 3960 2512
rect 40 2408 72 2440
rect 112 2408 144 2440
rect 184 2408 216 2440
rect 256 2408 288 2440
rect 328 2408 360 2440
rect 400 2408 432 2440
rect 472 2408 504 2440
rect 544 2408 576 2440
rect 616 2408 648 2440
rect 688 2408 720 2440
rect 760 2408 792 2440
rect 832 2408 864 2440
rect 904 2408 936 2440
rect 976 2408 1008 2440
rect 1048 2408 1080 2440
rect 1120 2408 1152 2440
rect 1192 2408 1224 2440
rect 1264 2408 1296 2440
rect 1336 2408 1368 2440
rect 1408 2408 1440 2440
rect 1480 2408 1512 2440
rect 1552 2408 1584 2440
rect 1624 2408 1656 2440
rect 1696 2408 1728 2440
rect 1768 2408 1800 2440
rect 1840 2408 1872 2440
rect 1912 2408 1944 2440
rect 1984 2408 2016 2440
rect 2056 2408 2088 2440
rect 2128 2408 2160 2440
rect 2200 2408 2232 2440
rect 2272 2408 2304 2440
rect 2344 2408 2376 2440
rect 2416 2408 2448 2440
rect 2488 2408 2520 2440
rect 2560 2408 2592 2440
rect 2632 2408 2664 2440
rect 2704 2408 2736 2440
rect 2776 2408 2808 2440
rect 2848 2408 2880 2440
rect 2920 2408 2952 2440
rect 2992 2408 3024 2440
rect 3064 2408 3096 2440
rect 3136 2408 3168 2440
rect 3208 2408 3240 2440
rect 3280 2408 3312 2440
rect 3352 2408 3384 2440
rect 3424 2408 3456 2440
rect 3496 2408 3528 2440
rect 3568 2408 3600 2440
rect 3640 2408 3672 2440
rect 3712 2408 3744 2440
rect 3784 2408 3816 2440
rect 3856 2408 3888 2440
rect 3928 2408 3960 2440
rect 40 2336 72 2368
rect 112 2336 144 2368
rect 184 2336 216 2368
rect 256 2336 288 2368
rect 328 2336 360 2368
rect 400 2336 432 2368
rect 472 2336 504 2368
rect 544 2336 576 2368
rect 616 2336 648 2368
rect 688 2336 720 2368
rect 760 2336 792 2368
rect 832 2336 864 2368
rect 904 2336 936 2368
rect 976 2336 1008 2368
rect 1048 2336 1080 2368
rect 1120 2336 1152 2368
rect 1192 2336 1224 2368
rect 1264 2336 1296 2368
rect 1336 2336 1368 2368
rect 1408 2336 1440 2368
rect 1480 2336 1512 2368
rect 1552 2336 1584 2368
rect 1624 2336 1656 2368
rect 1696 2336 1728 2368
rect 1768 2336 1800 2368
rect 1840 2336 1872 2368
rect 1912 2336 1944 2368
rect 1984 2336 2016 2368
rect 2056 2336 2088 2368
rect 2128 2336 2160 2368
rect 2200 2336 2232 2368
rect 2272 2336 2304 2368
rect 2344 2336 2376 2368
rect 2416 2336 2448 2368
rect 2488 2336 2520 2368
rect 2560 2336 2592 2368
rect 2632 2336 2664 2368
rect 2704 2336 2736 2368
rect 2776 2336 2808 2368
rect 2848 2336 2880 2368
rect 2920 2336 2952 2368
rect 2992 2336 3024 2368
rect 3064 2336 3096 2368
rect 3136 2336 3168 2368
rect 3208 2336 3240 2368
rect 3280 2336 3312 2368
rect 3352 2336 3384 2368
rect 3424 2336 3456 2368
rect 3496 2336 3528 2368
rect 3568 2336 3600 2368
rect 3640 2336 3672 2368
rect 3712 2336 3744 2368
rect 3784 2336 3816 2368
rect 3856 2336 3888 2368
rect 3928 2336 3960 2368
rect 40 2264 72 2296
rect 112 2264 144 2296
rect 184 2264 216 2296
rect 256 2264 288 2296
rect 328 2264 360 2296
rect 400 2264 432 2296
rect 472 2264 504 2296
rect 544 2264 576 2296
rect 616 2264 648 2296
rect 688 2264 720 2296
rect 760 2264 792 2296
rect 832 2264 864 2296
rect 904 2264 936 2296
rect 976 2264 1008 2296
rect 1048 2264 1080 2296
rect 1120 2264 1152 2296
rect 1192 2264 1224 2296
rect 1264 2264 1296 2296
rect 1336 2264 1368 2296
rect 1408 2264 1440 2296
rect 1480 2264 1512 2296
rect 1552 2264 1584 2296
rect 1624 2264 1656 2296
rect 1696 2264 1728 2296
rect 1768 2264 1800 2296
rect 1840 2264 1872 2296
rect 1912 2264 1944 2296
rect 1984 2264 2016 2296
rect 2056 2264 2088 2296
rect 2128 2264 2160 2296
rect 2200 2264 2232 2296
rect 2272 2264 2304 2296
rect 2344 2264 2376 2296
rect 2416 2264 2448 2296
rect 2488 2264 2520 2296
rect 2560 2264 2592 2296
rect 2632 2264 2664 2296
rect 2704 2264 2736 2296
rect 2776 2264 2808 2296
rect 2848 2264 2880 2296
rect 2920 2264 2952 2296
rect 2992 2264 3024 2296
rect 3064 2264 3096 2296
rect 3136 2264 3168 2296
rect 3208 2264 3240 2296
rect 3280 2264 3312 2296
rect 3352 2264 3384 2296
rect 3424 2264 3456 2296
rect 3496 2264 3528 2296
rect 3568 2264 3600 2296
rect 3640 2264 3672 2296
rect 3712 2264 3744 2296
rect 3784 2264 3816 2296
rect 3856 2264 3888 2296
rect 3928 2264 3960 2296
rect 40 2192 72 2224
rect 112 2192 144 2224
rect 184 2192 216 2224
rect 256 2192 288 2224
rect 328 2192 360 2224
rect 400 2192 432 2224
rect 472 2192 504 2224
rect 544 2192 576 2224
rect 616 2192 648 2224
rect 688 2192 720 2224
rect 760 2192 792 2224
rect 832 2192 864 2224
rect 904 2192 936 2224
rect 976 2192 1008 2224
rect 1048 2192 1080 2224
rect 1120 2192 1152 2224
rect 1192 2192 1224 2224
rect 1264 2192 1296 2224
rect 1336 2192 1368 2224
rect 1408 2192 1440 2224
rect 1480 2192 1512 2224
rect 1552 2192 1584 2224
rect 1624 2192 1656 2224
rect 1696 2192 1728 2224
rect 1768 2192 1800 2224
rect 1840 2192 1872 2224
rect 1912 2192 1944 2224
rect 1984 2192 2016 2224
rect 2056 2192 2088 2224
rect 2128 2192 2160 2224
rect 2200 2192 2232 2224
rect 2272 2192 2304 2224
rect 2344 2192 2376 2224
rect 2416 2192 2448 2224
rect 2488 2192 2520 2224
rect 2560 2192 2592 2224
rect 2632 2192 2664 2224
rect 2704 2192 2736 2224
rect 2776 2192 2808 2224
rect 2848 2192 2880 2224
rect 2920 2192 2952 2224
rect 2992 2192 3024 2224
rect 3064 2192 3096 2224
rect 3136 2192 3168 2224
rect 3208 2192 3240 2224
rect 3280 2192 3312 2224
rect 3352 2192 3384 2224
rect 3424 2192 3456 2224
rect 3496 2192 3528 2224
rect 3568 2192 3600 2224
rect 3640 2192 3672 2224
rect 3712 2192 3744 2224
rect 3784 2192 3816 2224
rect 3856 2192 3888 2224
rect 3928 2192 3960 2224
rect 40 2120 72 2152
rect 112 2120 144 2152
rect 184 2120 216 2152
rect 256 2120 288 2152
rect 328 2120 360 2152
rect 400 2120 432 2152
rect 472 2120 504 2152
rect 544 2120 576 2152
rect 616 2120 648 2152
rect 688 2120 720 2152
rect 760 2120 792 2152
rect 832 2120 864 2152
rect 904 2120 936 2152
rect 976 2120 1008 2152
rect 1048 2120 1080 2152
rect 1120 2120 1152 2152
rect 1192 2120 1224 2152
rect 1264 2120 1296 2152
rect 1336 2120 1368 2152
rect 1408 2120 1440 2152
rect 1480 2120 1512 2152
rect 1552 2120 1584 2152
rect 1624 2120 1656 2152
rect 1696 2120 1728 2152
rect 1768 2120 1800 2152
rect 1840 2120 1872 2152
rect 1912 2120 1944 2152
rect 1984 2120 2016 2152
rect 2056 2120 2088 2152
rect 2128 2120 2160 2152
rect 2200 2120 2232 2152
rect 2272 2120 2304 2152
rect 2344 2120 2376 2152
rect 2416 2120 2448 2152
rect 2488 2120 2520 2152
rect 2560 2120 2592 2152
rect 2632 2120 2664 2152
rect 2704 2120 2736 2152
rect 2776 2120 2808 2152
rect 2848 2120 2880 2152
rect 2920 2120 2952 2152
rect 2992 2120 3024 2152
rect 3064 2120 3096 2152
rect 3136 2120 3168 2152
rect 3208 2120 3240 2152
rect 3280 2120 3312 2152
rect 3352 2120 3384 2152
rect 3424 2120 3456 2152
rect 3496 2120 3528 2152
rect 3568 2120 3600 2152
rect 3640 2120 3672 2152
rect 3712 2120 3744 2152
rect 3784 2120 3816 2152
rect 3856 2120 3888 2152
rect 3928 2120 3960 2152
rect 40 2048 72 2080
rect 112 2048 144 2080
rect 184 2048 216 2080
rect 256 2048 288 2080
rect 328 2048 360 2080
rect 400 2048 432 2080
rect 472 2048 504 2080
rect 544 2048 576 2080
rect 616 2048 648 2080
rect 688 2048 720 2080
rect 760 2048 792 2080
rect 832 2048 864 2080
rect 904 2048 936 2080
rect 976 2048 1008 2080
rect 1048 2048 1080 2080
rect 1120 2048 1152 2080
rect 1192 2048 1224 2080
rect 1264 2048 1296 2080
rect 1336 2048 1368 2080
rect 1408 2048 1440 2080
rect 1480 2048 1512 2080
rect 1552 2048 1584 2080
rect 1624 2048 1656 2080
rect 1696 2048 1728 2080
rect 1768 2048 1800 2080
rect 1840 2048 1872 2080
rect 1912 2048 1944 2080
rect 1984 2048 2016 2080
rect 2056 2048 2088 2080
rect 2128 2048 2160 2080
rect 2200 2048 2232 2080
rect 2272 2048 2304 2080
rect 2344 2048 2376 2080
rect 2416 2048 2448 2080
rect 2488 2048 2520 2080
rect 2560 2048 2592 2080
rect 2632 2048 2664 2080
rect 2704 2048 2736 2080
rect 2776 2048 2808 2080
rect 2848 2048 2880 2080
rect 2920 2048 2952 2080
rect 2992 2048 3024 2080
rect 3064 2048 3096 2080
rect 3136 2048 3168 2080
rect 3208 2048 3240 2080
rect 3280 2048 3312 2080
rect 3352 2048 3384 2080
rect 3424 2048 3456 2080
rect 3496 2048 3528 2080
rect 3568 2048 3600 2080
rect 3640 2048 3672 2080
rect 3712 2048 3744 2080
rect 3784 2048 3816 2080
rect 3856 2048 3888 2080
rect 3928 2048 3960 2080
rect 40 1976 72 2008
rect 112 1976 144 2008
rect 184 1976 216 2008
rect 256 1976 288 2008
rect 328 1976 360 2008
rect 400 1976 432 2008
rect 472 1976 504 2008
rect 544 1976 576 2008
rect 616 1976 648 2008
rect 688 1976 720 2008
rect 760 1976 792 2008
rect 832 1976 864 2008
rect 904 1976 936 2008
rect 976 1976 1008 2008
rect 1048 1976 1080 2008
rect 1120 1976 1152 2008
rect 1192 1976 1224 2008
rect 1264 1976 1296 2008
rect 1336 1976 1368 2008
rect 1408 1976 1440 2008
rect 1480 1976 1512 2008
rect 1552 1976 1584 2008
rect 1624 1976 1656 2008
rect 1696 1976 1728 2008
rect 1768 1976 1800 2008
rect 1840 1976 1872 2008
rect 1912 1976 1944 2008
rect 1984 1976 2016 2008
rect 2056 1976 2088 2008
rect 2128 1976 2160 2008
rect 2200 1976 2232 2008
rect 2272 1976 2304 2008
rect 2344 1976 2376 2008
rect 2416 1976 2448 2008
rect 2488 1976 2520 2008
rect 2560 1976 2592 2008
rect 2632 1976 2664 2008
rect 2704 1976 2736 2008
rect 2776 1976 2808 2008
rect 2848 1976 2880 2008
rect 2920 1976 2952 2008
rect 2992 1976 3024 2008
rect 3064 1976 3096 2008
rect 3136 1976 3168 2008
rect 3208 1976 3240 2008
rect 3280 1976 3312 2008
rect 3352 1976 3384 2008
rect 3424 1976 3456 2008
rect 3496 1976 3528 2008
rect 3568 1976 3600 2008
rect 3640 1976 3672 2008
rect 3712 1976 3744 2008
rect 3784 1976 3816 2008
rect 3856 1976 3888 2008
rect 3928 1976 3960 2008
rect 40 1904 72 1936
rect 112 1904 144 1936
rect 184 1904 216 1936
rect 256 1904 288 1936
rect 328 1904 360 1936
rect 400 1904 432 1936
rect 472 1904 504 1936
rect 544 1904 576 1936
rect 616 1904 648 1936
rect 688 1904 720 1936
rect 760 1904 792 1936
rect 832 1904 864 1936
rect 904 1904 936 1936
rect 976 1904 1008 1936
rect 1048 1904 1080 1936
rect 1120 1904 1152 1936
rect 1192 1904 1224 1936
rect 1264 1904 1296 1936
rect 1336 1904 1368 1936
rect 1408 1904 1440 1936
rect 1480 1904 1512 1936
rect 1552 1904 1584 1936
rect 1624 1904 1656 1936
rect 1696 1904 1728 1936
rect 1768 1904 1800 1936
rect 1840 1904 1872 1936
rect 1912 1904 1944 1936
rect 1984 1904 2016 1936
rect 2056 1904 2088 1936
rect 2128 1904 2160 1936
rect 2200 1904 2232 1936
rect 2272 1904 2304 1936
rect 2344 1904 2376 1936
rect 2416 1904 2448 1936
rect 2488 1904 2520 1936
rect 2560 1904 2592 1936
rect 2632 1904 2664 1936
rect 2704 1904 2736 1936
rect 2776 1904 2808 1936
rect 2848 1904 2880 1936
rect 2920 1904 2952 1936
rect 2992 1904 3024 1936
rect 3064 1904 3096 1936
rect 3136 1904 3168 1936
rect 3208 1904 3240 1936
rect 3280 1904 3312 1936
rect 3352 1904 3384 1936
rect 3424 1904 3456 1936
rect 3496 1904 3528 1936
rect 3568 1904 3600 1936
rect 3640 1904 3672 1936
rect 3712 1904 3744 1936
rect 3784 1904 3816 1936
rect 3856 1904 3888 1936
rect 3928 1904 3960 1936
rect 40 1832 72 1864
rect 112 1832 144 1864
rect 184 1832 216 1864
rect 256 1832 288 1864
rect 328 1832 360 1864
rect 400 1832 432 1864
rect 472 1832 504 1864
rect 544 1832 576 1864
rect 616 1832 648 1864
rect 688 1832 720 1864
rect 760 1832 792 1864
rect 832 1832 864 1864
rect 904 1832 936 1864
rect 976 1832 1008 1864
rect 1048 1832 1080 1864
rect 1120 1832 1152 1864
rect 1192 1832 1224 1864
rect 1264 1832 1296 1864
rect 1336 1832 1368 1864
rect 1408 1832 1440 1864
rect 1480 1832 1512 1864
rect 1552 1832 1584 1864
rect 1624 1832 1656 1864
rect 1696 1832 1728 1864
rect 1768 1832 1800 1864
rect 1840 1832 1872 1864
rect 1912 1832 1944 1864
rect 1984 1832 2016 1864
rect 2056 1832 2088 1864
rect 2128 1832 2160 1864
rect 2200 1832 2232 1864
rect 2272 1832 2304 1864
rect 2344 1832 2376 1864
rect 2416 1832 2448 1864
rect 2488 1832 2520 1864
rect 2560 1832 2592 1864
rect 2632 1832 2664 1864
rect 2704 1832 2736 1864
rect 2776 1832 2808 1864
rect 2848 1832 2880 1864
rect 2920 1832 2952 1864
rect 2992 1832 3024 1864
rect 3064 1832 3096 1864
rect 3136 1832 3168 1864
rect 3208 1832 3240 1864
rect 3280 1832 3312 1864
rect 3352 1832 3384 1864
rect 3424 1832 3456 1864
rect 3496 1832 3528 1864
rect 3568 1832 3600 1864
rect 3640 1832 3672 1864
rect 3712 1832 3744 1864
rect 3784 1832 3816 1864
rect 3856 1832 3888 1864
rect 3928 1832 3960 1864
rect 40 1760 72 1792
rect 112 1760 144 1792
rect 184 1760 216 1792
rect 256 1760 288 1792
rect 328 1760 360 1792
rect 400 1760 432 1792
rect 472 1760 504 1792
rect 544 1760 576 1792
rect 616 1760 648 1792
rect 688 1760 720 1792
rect 760 1760 792 1792
rect 832 1760 864 1792
rect 904 1760 936 1792
rect 976 1760 1008 1792
rect 1048 1760 1080 1792
rect 1120 1760 1152 1792
rect 1192 1760 1224 1792
rect 1264 1760 1296 1792
rect 1336 1760 1368 1792
rect 1408 1760 1440 1792
rect 1480 1760 1512 1792
rect 1552 1760 1584 1792
rect 1624 1760 1656 1792
rect 1696 1760 1728 1792
rect 1768 1760 1800 1792
rect 1840 1760 1872 1792
rect 1912 1760 1944 1792
rect 1984 1760 2016 1792
rect 2056 1760 2088 1792
rect 2128 1760 2160 1792
rect 2200 1760 2232 1792
rect 2272 1760 2304 1792
rect 2344 1760 2376 1792
rect 2416 1760 2448 1792
rect 2488 1760 2520 1792
rect 2560 1760 2592 1792
rect 2632 1760 2664 1792
rect 2704 1760 2736 1792
rect 2776 1760 2808 1792
rect 2848 1760 2880 1792
rect 2920 1760 2952 1792
rect 2992 1760 3024 1792
rect 3064 1760 3096 1792
rect 3136 1760 3168 1792
rect 3208 1760 3240 1792
rect 3280 1760 3312 1792
rect 3352 1760 3384 1792
rect 3424 1760 3456 1792
rect 3496 1760 3528 1792
rect 3568 1760 3600 1792
rect 3640 1760 3672 1792
rect 3712 1760 3744 1792
rect 3784 1760 3816 1792
rect 3856 1760 3888 1792
rect 3928 1760 3960 1792
rect 40 1688 72 1720
rect 112 1688 144 1720
rect 184 1688 216 1720
rect 256 1688 288 1720
rect 328 1688 360 1720
rect 400 1688 432 1720
rect 472 1688 504 1720
rect 544 1688 576 1720
rect 616 1688 648 1720
rect 688 1688 720 1720
rect 760 1688 792 1720
rect 832 1688 864 1720
rect 904 1688 936 1720
rect 976 1688 1008 1720
rect 1048 1688 1080 1720
rect 1120 1688 1152 1720
rect 1192 1688 1224 1720
rect 1264 1688 1296 1720
rect 1336 1688 1368 1720
rect 1408 1688 1440 1720
rect 1480 1688 1512 1720
rect 1552 1688 1584 1720
rect 1624 1688 1656 1720
rect 1696 1688 1728 1720
rect 1768 1688 1800 1720
rect 1840 1688 1872 1720
rect 1912 1688 1944 1720
rect 1984 1688 2016 1720
rect 2056 1688 2088 1720
rect 2128 1688 2160 1720
rect 2200 1688 2232 1720
rect 2272 1688 2304 1720
rect 2344 1688 2376 1720
rect 2416 1688 2448 1720
rect 2488 1688 2520 1720
rect 2560 1688 2592 1720
rect 2632 1688 2664 1720
rect 2704 1688 2736 1720
rect 2776 1688 2808 1720
rect 2848 1688 2880 1720
rect 2920 1688 2952 1720
rect 2992 1688 3024 1720
rect 3064 1688 3096 1720
rect 3136 1688 3168 1720
rect 3208 1688 3240 1720
rect 3280 1688 3312 1720
rect 3352 1688 3384 1720
rect 3424 1688 3456 1720
rect 3496 1688 3528 1720
rect 3568 1688 3600 1720
rect 3640 1688 3672 1720
rect 3712 1688 3744 1720
rect 3784 1688 3816 1720
rect 3856 1688 3888 1720
rect 3928 1688 3960 1720
rect 40 1616 72 1648
rect 112 1616 144 1648
rect 184 1616 216 1648
rect 256 1616 288 1648
rect 328 1616 360 1648
rect 400 1616 432 1648
rect 472 1616 504 1648
rect 544 1616 576 1648
rect 616 1616 648 1648
rect 688 1616 720 1648
rect 760 1616 792 1648
rect 832 1616 864 1648
rect 904 1616 936 1648
rect 976 1616 1008 1648
rect 1048 1616 1080 1648
rect 1120 1616 1152 1648
rect 1192 1616 1224 1648
rect 1264 1616 1296 1648
rect 1336 1616 1368 1648
rect 1408 1616 1440 1648
rect 1480 1616 1512 1648
rect 1552 1616 1584 1648
rect 1624 1616 1656 1648
rect 1696 1616 1728 1648
rect 1768 1616 1800 1648
rect 1840 1616 1872 1648
rect 1912 1616 1944 1648
rect 1984 1616 2016 1648
rect 2056 1616 2088 1648
rect 2128 1616 2160 1648
rect 2200 1616 2232 1648
rect 2272 1616 2304 1648
rect 2344 1616 2376 1648
rect 2416 1616 2448 1648
rect 2488 1616 2520 1648
rect 2560 1616 2592 1648
rect 2632 1616 2664 1648
rect 2704 1616 2736 1648
rect 2776 1616 2808 1648
rect 2848 1616 2880 1648
rect 2920 1616 2952 1648
rect 2992 1616 3024 1648
rect 3064 1616 3096 1648
rect 3136 1616 3168 1648
rect 3208 1616 3240 1648
rect 3280 1616 3312 1648
rect 3352 1616 3384 1648
rect 3424 1616 3456 1648
rect 3496 1616 3528 1648
rect 3568 1616 3600 1648
rect 3640 1616 3672 1648
rect 3712 1616 3744 1648
rect 3784 1616 3816 1648
rect 3856 1616 3888 1648
rect 3928 1616 3960 1648
rect 40 1544 72 1576
rect 112 1544 144 1576
rect 184 1544 216 1576
rect 256 1544 288 1576
rect 328 1544 360 1576
rect 400 1544 432 1576
rect 472 1544 504 1576
rect 544 1544 576 1576
rect 616 1544 648 1576
rect 688 1544 720 1576
rect 760 1544 792 1576
rect 832 1544 864 1576
rect 904 1544 936 1576
rect 976 1544 1008 1576
rect 1048 1544 1080 1576
rect 1120 1544 1152 1576
rect 1192 1544 1224 1576
rect 1264 1544 1296 1576
rect 1336 1544 1368 1576
rect 1408 1544 1440 1576
rect 1480 1544 1512 1576
rect 1552 1544 1584 1576
rect 1624 1544 1656 1576
rect 1696 1544 1728 1576
rect 1768 1544 1800 1576
rect 1840 1544 1872 1576
rect 1912 1544 1944 1576
rect 1984 1544 2016 1576
rect 2056 1544 2088 1576
rect 2128 1544 2160 1576
rect 2200 1544 2232 1576
rect 2272 1544 2304 1576
rect 2344 1544 2376 1576
rect 2416 1544 2448 1576
rect 2488 1544 2520 1576
rect 2560 1544 2592 1576
rect 2632 1544 2664 1576
rect 2704 1544 2736 1576
rect 2776 1544 2808 1576
rect 2848 1544 2880 1576
rect 2920 1544 2952 1576
rect 2992 1544 3024 1576
rect 3064 1544 3096 1576
rect 3136 1544 3168 1576
rect 3208 1544 3240 1576
rect 3280 1544 3312 1576
rect 3352 1544 3384 1576
rect 3424 1544 3456 1576
rect 3496 1544 3528 1576
rect 3568 1544 3600 1576
rect 3640 1544 3672 1576
rect 3712 1544 3744 1576
rect 3784 1544 3816 1576
rect 3856 1544 3888 1576
rect 3928 1544 3960 1576
rect 40 1472 72 1504
rect 112 1472 144 1504
rect 184 1472 216 1504
rect 256 1472 288 1504
rect 328 1472 360 1504
rect 400 1472 432 1504
rect 472 1472 504 1504
rect 544 1472 576 1504
rect 616 1472 648 1504
rect 688 1472 720 1504
rect 760 1472 792 1504
rect 832 1472 864 1504
rect 904 1472 936 1504
rect 976 1472 1008 1504
rect 1048 1472 1080 1504
rect 1120 1472 1152 1504
rect 1192 1472 1224 1504
rect 1264 1472 1296 1504
rect 1336 1472 1368 1504
rect 1408 1472 1440 1504
rect 1480 1472 1512 1504
rect 1552 1472 1584 1504
rect 1624 1472 1656 1504
rect 1696 1472 1728 1504
rect 1768 1472 1800 1504
rect 1840 1472 1872 1504
rect 1912 1472 1944 1504
rect 1984 1472 2016 1504
rect 2056 1472 2088 1504
rect 2128 1472 2160 1504
rect 2200 1472 2232 1504
rect 2272 1472 2304 1504
rect 2344 1472 2376 1504
rect 2416 1472 2448 1504
rect 2488 1472 2520 1504
rect 2560 1472 2592 1504
rect 2632 1472 2664 1504
rect 2704 1472 2736 1504
rect 2776 1472 2808 1504
rect 2848 1472 2880 1504
rect 2920 1472 2952 1504
rect 2992 1472 3024 1504
rect 3064 1472 3096 1504
rect 3136 1472 3168 1504
rect 3208 1472 3240 1504
rect 3280 1472 3312 1504
rect 3352 1472 3384 1504
rect 3424 1472 3456 1504
rect 3496 1472 3528 1504
rect 3568 1472 3600 1504
rect 3640 1472 3672 1504
rect 3712 1472 3744 1504
rect 3784 1472 3816 1504
rect 3856 1472 3888 1504
rect 3928 1472 3960 1504
rect 40 1400 72 1432
rect 112 1400 144 1432
rect 184 1400 216 1432
rect 256 1400 288 1432
rect 328 1400 360 1432
rect 400 1400 432 1432
rect 472 1400 504 1432
rect 544 1400 576 1432
rect 616 1400 648 1432
rect 688 1400 720 1432
rect 760 1400 792 1432
rect 832 1400 864 1432
rect 904 1400 936 1432
rect 976 1400 1008 1432
rect 1048 1400 1080 1432
rect 1120 1400 1152 1432
rect 1192 1400 1224 1432
rect 1264 1400 1296 1432
rect 1336 1400 1368 1432
rect 1408 1400 1440 1432
rect 1480 1400 1512 1432
rect 1552 1400 1584 1432
rect 1624 1400 1656 1432
rect 1696 1400 1728 1432
rect 1768 1400 1800 1432
rect 1840 1400 1872 1432
rect 1912 1400 1944 1432
rect 1984 1400 2016 1432
rect 2056 1400 2088 1432
rect 2128 1400 2160 1432
rect 2200 1400 2232 1432
rect 2272 1400 2304 1432
rect 2344 1400 2376 1432
rect 2416 1400 2448 1432
rect 2488 1400 2520 1432
rect 2560 1400 2592 1432
rect 2632 1400 2664 1432
rect 2704 1400 2736 1432
rect 2776 1400 2808 1432
rect 2848 1400 2880 1432
rect 2920 1400 2952 1432
rect 2992 1400 3024 1432
rect 3064 1400 3096 1432
rect 3136 1400 3168 1432
rect 3208 1400 3240 1432
rect 3280 1400 3312 1432
rect 3352 1400 3384 1432
rect 3424 1400 3456 1432
rect 3496 1400 3528 1432
rect 3568 1400 3600 1432
rect 3640 1400 3672 1432
rect 3712 1400 3744 1432
rect 3784 1400 3816 1432
rect 3856 1400 3888 1432
rect 3928 1400 3960 1432
rect 40 1328 72 1360
rect 112 1328 144 1360
rect 184 1328 216 1360
rect 256 1328 288 1360
rect 328 1328 360 1360
rect 400 1328 432 1360
rect 472 1328 504 1360
rect 544 1328 576 1360
rect 616 1328 648 1360
rect 688 1328 720 1360
rect 760 1328 792 1360
rect 832 1328 864 1360
rect 904 1328 936 1360
rect 976 1328 1008 1360
rect 1048 1328 1080 1360
rect 1120 1328 1152 1360
rect 1192 1328 1224 1360
rect 1264 1328 1296 1360
rect 1336 1328 1368 1360
rect 1408 1328 1440 1360
rect 1480 1328 1512 1360
rect 1552 1328 1584 1360
rect 1624 1328 1656 1360
rect 1696 1328 1728 1360
rect 1768 1328 1800 1360
rect 1840 1328 1872 1360
rect 1912 1328 1944 1360
rect 1984 1328 2016 1360
rect 2056 1328 2088 1360
rect 2128 1328 2160 1360
rect 2200 1328 2232 1360
rect 2272 1328 2304 1360
rect 2344 1328 2376 1360
rect 2416 1328 2448 1360
rect 2488 1328 2520 1360
rect 2560 1328 2592 1360
rect 2632 1328 2664 1360
rect 2704 1328 2736 1360
rect 2776 1328 2808 1360
rect 2848 1328 2880 1360
rect 2920 1328 2952 1360
rect 2992 1328 3024 1360
rect 3064 1328 3096 1360
rect 3136 1328 3168 1360
rect 3208 1328 3240 1360
rect 3280 1328 3312 1360
rect 3352 1328 3384 1360
rect 3424 1328 3456 1360
rect 3496 1328 3528 1360
rect 3568 1328 3600 1360
rect 3640 1328 3672 1360
rect 3712 1328 3744 1360
rect 3784 1328 3816 1360
rect 3856 1328 3888 1360
rect 3928 1328 3960 1360
rect 40 1256 72 1288
rect 112 1256 144 1288
rect 184 1256 216 1288
rect 256 1256 288 1288
rect 328 1256 360 1288
rect 400 1256 432 1288
rect 472 1256 504 1288
rect 544 1256 576 1288
rect 616 1256 648 1288
rect 688 1256 720 1288
rect 760 1256 792 1288
rect 832 1256 864 1288
rect 904 1256 936 1288
rect 976 1256 1008 1288
rect 1048 1256 1080 1288
rect 1120 1256 1152 1288
rect 1192 1256 1224 1288
rect 1264 1256 1296 1288
rect 1336 1256 1368 1288
rect 1408 1256 1440 1288
rect 1480 1256 1512 1288
rect 1552 1256 1584 1288
rect 1624 1256 1656 1288
rect 1696 1256 1728 1288
rect 1768 1256 1800 1288
rect 1840 1256 1872 1288
rect 1912 1256 1944 1288
rect 1984 1256 2016 1288
rect 2056 1256 2088 1288
rect 2128 1256 2160 1288
rect 2200 1256 2232 1288
rect 2272 1256 2304 1288
rect 2344 1256 2376 1288
rect 2416 1256 2448 1288
rect 2488 1256 2520 1288
rect 2560 1256 2592 1288
rect 2632 1256 2664 1288
rect 2704 1256 2736 1288
rect 2776 1256 2808 1288
rect 2848 1256 2880 1288
rect 2920 1256 2952 1288
rect 2992 1256 3024 1288
rect 3064 1256 3096 1288
rect 3136 1256 3168 1288
rect 3208 1256 3240 1288
rect 3280 1256 3312 1288
rect 3352 1256 3384 1288
rect 3424 1256 3456 1288
rect 3496 1256 3528 1288
rect 3568 1256 3600 1288
rect 3640 1256 3672 1288
rect 3712 1256 3744 1288
rect 3784 1256 3816 1288
rect 3856 1256 3888 1288
rect 3928 1256 3960 1288
rect 184 31384 216 31416
rect 256 31384 288 31416
rect 328 31384 360 31416
rect 400 31384 432 31416
rect 472 31384 504 31416
rect 544 31384 576 31416
rect 616 31384 648 31416
rect 688 31384 720 31416
rect 760 31384 792 31416
rect 832 31384 864 31416
rect 904 31384 936 31416
rect 976 31384 1008 31416
rect 1048 31384 1080 31416
rect 1120 31384 1152 31416
rect 1192 31384 1224 31416
rect 1264 31384 1296 31416
rect 1336 31384 1368 31416
rect 1408 31384 1440 31416
rect 1480 31384 1512 31416
rect 1552 31384 1584 31416
rect 1624 31384 1656 31416
rect 1696 31384 1728 31416
rect 1768 31384 1800 31416
rect 1840 31384 1872 31416
rect 1912 31384 1944 31416
rect 1984 31384 2016 31416
rect 2056 31384 2088 31416
rect 2128 31384 2160 31416
rect 2200 31384 2232 31416
rect 2272 31384 2304 31416
rect 2344 31384 2376 31416
rect 2416 31384 2448 31416
rect 2488 31384 2520 31416
rect 2560 31384 2592 31416
rect 2632 31384 2664 31416
rect 2704 31384 2736 31416
rect 2776 31384 2808 31416
rect 2848 31384 2880 31416
rect 2920 31384 2952 31416
rect 2992 31384 3024 31416
rect 3064 31384 3096 31416
rect 3136 31384 3168 31416
rect 3208 31384 3240 31416
rect 3280 31384 3312 31416
rect 3352 31384 3384 31416
rect 3424 31384 3456 31416
rect 3496 31384 3528 31416
rect 3568 31384 3600 31416
rect 3640 31384 3672 31416
rect 3712 31384 3744 31416
rect 3784 31384 3816 31416
rect 3856 31384 3888 31416
rect 184 27939 216 27971
rect 256 27939 288 27971
rect 328 27939 360 27971
rect 400 27939 432 27971
rect 472 27939 504 27971
rect 544 27939 576 27971
rect 616 27939 648 27971
rect 688 27939 720 27971
rect 760 27939 792 27971
rect 832 27939 864 27971
rect 904 27939 936 27971
rect 976 27939 1008 27971
rect 1048 27939 1080 27971
rect 1120 27939 1152 27971
rect 1192 27939 1224 27971
rect 1264 27939 1296 27971
rect 1336 27939 1368 27971
rect 1408 27939 1440 27971
rect 1480 27939 1512 27971
rect 1552 27939 1584 27971
rect 1624 27939 1656 27971
rect 1696 27939 1728 27971
rect 1768 27939 1800 27971
rect 1840 27939 1872 27971
rect 1912 27939 1944 27971
rect 1984 27939 2016 27971
rect 2056 27939 2088 27971
rect 2128 27939 2160 27971
rect 2200 27939 2232 27971
rect 2272 27939 2304 27971
rect 2344 27939 2376 27971
rect 2416 27939 2448 27971
rect 2488 27939 2520 27971
rect 2560 27939 2592 27971
rect 2632 27939 2664 27971
rect 2704 27939 2736 27971
rect 2776 27939 2808 27971
rect 2848 27939 2880 27971
rect 2920 27939 2952 27971
rect 2992 27939 3024 27971
rect 3064 27939 3096 27971
rect 3136 27939 3168 27971
rect 3208 27939 3240 27971
rect 3280 27939 3312 27971
rect 3352 27939 3384 27971
rect 3424 27939 3456 27971
rect 3496 27939 3528 27971
rect 3568 27939 3600 27971
rect 3640 27939 3672 27971
rect 3712 27939 3744 27971
rect 3784 27939 3816 27971
rect 3856 27939 3888 27971
rect 112 27867 144 27899
rect 184 27867 216 27899
rect 256 27867 288 27899
rect 328 27867 360 27899
rect 400 27867 432 27899
rect 472 27867 504 27899
rect 544 27867 576 27899
rect 616 27867 648 27899
rect 688 27867 720 27899
rect 760 27867 792 27899
rect 832 27867 864 27899
rect 904 27867 936 27899
rect 976 27867 1008 27899
rect 1048 27867 1080 27899
rect 1120 27867 1152 27899
rect 1192 27867 1224 27899
rect 1264 27867 1296 27899
rect 1336 27867 1368 27899
rect 1408 27867 1440 27899
rect 1480 27867 1512 27899
rect 1552 27867 1584 27899
rect 1624 27867 1656 27899
rect 1696 27867 1728 27899
rect 1768 27867 1800 27899
rect 1840 27867 1872 27899
rect 1912 27867 1944 27899
rect 1984 27867 2016 27899
rect 2056 27867 2088 27899
rect 2128 27867 2160 27899
rect 2200 27867 2232 27899
rect 2272 27867 2304 27899
rect 2344 27867 2376 27899
rect 2416 27867 2448 27899
rect 2488 27867 2520 27899
rect 2560 27867 2592 27899
rect 2632 27867 2664 27899
rect 2704 27867 2736 27899
rect 2776 27867 2808 27899
rect 2848 27867 2880 27899
rect 2920 27867 2952 27899
rect 2992 27867 3024 27899
rect 3064 27867 3096 27899
rect 3136 27867 3168 27899
rect 3208 27867 3240 27899
rect 3280 27867 3312 27899
rect 3352 27867 3384 27899
rect 3424 27867 3456 27899
rect 3496 27867 3528 27899
rect 3568 27867 3600 27899
rect 3640 27867 3672 27899
rect 3712 27867 3744 27899
rect 3784 27867 3816 27899
rect 3856 27867 3888 27899
rect 112 27795 144 27827
rect 184 27795 216 27827
rect 256 27795 288 27827
rect 328 27795 360 27827
rect 400 27795 432 27827
rect 472 27795 504 27827
rect 544 27795 576 27827
rect 616 27795 648 27827
rect 688 27795 720 27827
rect 760 27795 792 27827
rect 832 27795 864 27827
rect 904 27795 936 27827
rect 976 27795 1008 27827
rect 1048 27795 1080 27827
rect 1120 27795 1152 27827
rect 1192 27795 1224 27827
rect 1264 27795 1296 27827
rect 1336 27795 1368 27827
rect 1408 27795 1440 27827
rect 1480 27795 1512 27827
rect 1552 27795 1584 27827
rect 1624 27795 1656 27827
rect 1696 27795 1728 27827
rect 1768 27795 1800 27827
rect 1840 27795 1872 27827
rect 1912 27795 1944 27827
rect 1984 27795 2016 27827
rect 2056 27795 2088 27827
rect 2128 27795 2160 27827
rect 2200 27795 2232 27827
rect 2272 27795 2304 27827
rect 2344 27795 2376 27827
rect 2416 27795 2448 27827
rect 2488 27795 2520 27827
rect 2560 27795 2592 27827
rect 2632 27795 2664 27827
rect 2704 27795 2736 27827
rect 2776 27795 2808 27827
rect 2848 27795 2880 27827
rect 2920 27795 2952 27827
rect 2992 27795 3024 27827
rect 3064 27795 3096 27827
rect 3136 27795 3168 27827
rect 3208 27795 3240 27827
rect 3280 27795 3312 27827
rect 3352 27795 3384 27827
rect 3424 27795 3456 27827
rect 3496 27795 3528 27827
rect 3568 27795 3600 27827
rect 3640 27795 3672 27827
rect 3712 27795 3744 27827
rect 3784 27795 3816 27827
rect 3856 27795 3888 27827
rect 112 27723 144 27755
rect 184 27723 216 27755
rect 256 27723 288 27755
rect 328 27723 360 27755
rect 400 27723 432 27755
rect 472 27723 504 27755
rect 544 27723 576 27755
rect 616 27723 648 27755
rect 688 27723 720 27755
rect 760 27723 792 27755
rect 832 27723 864 27755
rect 904 27723 936 27755
rect 976 27723 1008 27755
rect 1048 27723 1080 27755
rect 1120 27723 1152 27755
rect 1192 27723 1224 27755
rect 1264 27723 1296 27755
rect 1336 27723 1368 27755
rect 1408 27723 1440 27755
rect 1480 27723 1512 27755
rect 1552 27723 1584 27755
rect 1624 27723 1656 27755
rect 1696 27723 1728 27755
rect 1768 27723 1800 27755
rect 1840 27723 1872 27755
rect 1912 27723 1944 27755
rect 1984 27723 2016 27755
rect 2056 27723 2088 27755
rect 2128 27723 2160 27755
rect 2200 27723 2232 27755
rect 2272 27723 2304 27755
rect 2344 27723 2376 27755
rect 2416 27723 2448 27755
rect 2488 27723 2520 27755
rect 2560 27723 2592 27755
rect 2632 27723 2664 27755
rect 2704 27723 2736 27755
rect 2776 27723 2808 27755
rect 2848 27723 2880 27755
rect 2920 27723 2952 27755
rect 2992 27723 3024 27755
rect 3064 27723 3096 27755
rect 3136 27723 3168 27755
rect 3208 27723 3240 27755
rect 3280 27723 3312 27755
rect 3352 27723 3384 27755
rect 3424 27723 3456 27755
rect 3496 27723 3528 27755
rect 3568 27723 3600 27755
rect 3640 27723 3672 27755
rect 3712 27723 3744 27755
rect 3784 27723 3816 27755
rect 3856 27723 3888 27755
rect 112 27651 144 27683
rect 184 27651 216 27683
rect 256 27651 288 27683
rect 328 27651 360 27683
rect 400 27651 432 27683
rect 472 27651 504 27683
rect 544 27651 576 27683
rect 616 27651 648 27683
rect 688 27651 720 27683
rect 760 27651 792 27683
rect 832 27651 864 27683
rect 904 27651 936 27683
rect 976 27651 1008 27683
rect 1048 27651 1080 27683
rect 1120 27651 1152 27683
rect 1192 27651 1224 27683
rect 1264 27651 1296 27683
rect 1336 27651 1368 27683
rect 1408 27651 1440 27683
rect 1480 27651 1512 27683
rect 1552 27651 1584 27683
rect 1624 27651 1656 27683
rect 1696 27651 1728 27683
rect 1768 27651 1800 27683
rect 1840 27651 1872 27683
rect 1912 27651 1944 27683
rect 1984 27651 2016 27683
rect 2056 27651 2088 27683
rect 2128 27651 2160 27683
rect 2200 27651 2232 27683
rect 2272 27651 2304 27683
rect 2344 27651 2376 27683
rect 2416 27651 2448 27683
rect 2488 27651 2520 27683
rect 2560 27651 2592 27683
rect 2632 27651 2664 27683
rect 2704 27651 2736 27683
rect 2776 27651 2808 27683
rect 2848 27651 2880 27683
rect 2920 27651 2952 27683
rect 2992 27651 3024 27683
rect 3064 27651 3096 27683
rect 3136 27651 3168 27683
rect 3208 27651 3240 27683
rect 3280 27651 3312 27683
rect 3352 27651 3384 27683
rect 3424 27651 3456 27683
rect 3496 27651 3528 27683
rect 3568 27651 3600 27683
rect 3640 27651 3672 27683
rect 3712 27651 3744 27683
rect 3784 27651 3816 27683
rect 3856 27651 3888 27683
rect 112 27579 144 27611
rect 184 27579 216 27611
rect 256 27579 288 27611
rect 328 27579 360 27611
rect 400 27579 432 27611
rect 472 27579 504 27611
rect 544 27579 576 27611
rect 616 27579 648 27611
rect 688 27579 720 27611
rect 760 27579 792 27611
rect 832 27579 864 27611
rect 904 27579 936 27611
rect 976 27579 1008 27611
rect 1048 27579 1080 27611
rect 1120 27579 1152 27611
rect 1192 27579 1224 27611
rect 1264 27579 1296 27611
rect 1336 27579 1368 27611
rect 1408 27579 1440 27611
rect 1480 27579 1512 27611
rect 1552 27579 1584 27611
rect 1624 27579 1656 27611
rect 1696 27579 1728 27611
rect 1768 27579 1800 27611
rect 1840 27579 1872 27611
rect 1912 27579 1944 27611
rect 1984 27579 2016 27611
rect 2056 27579 2088 27611
rect 2128 27579 2160 27611
rect 2200 27579 2232 27611
rect 2272 27579 2304 27611
rect 2344 27579 2376 27611
rect 2416 27579 2448 27611
rect 2488 27579 2520 27611
rect 2560 27579 2592 27611
rect 2632 27579 2664 27611
rect 2704 27579 2736 27611
rect 2776 27579 2808 27611
rect 2848 27579 2880 27611
rect 2920 27579 2952 27611
rect 2992 27579 3024 27611
rect 3064 27579 3096 27611
rect 3136 27579 3168 27611
rect 3208 27579 3240 27611
rect 3280 27579 3312 27611
rect 3352 27579 3384 27611
rect 3424 27579 3456 27611
rect 3496 27579 3528 27611
rect 3568 27579 3600 27611
rect 3640 27579 3672 27611
rect 3712 27579 3744 27611
rect 3784 27579 3816 27611
rect 3856 27579 3888 27611
rect 112 27507 144 27539
rect 184 27507 216 27539
rect 256 27507 288 27539
rect 328 27507 360 27539
rect 400 27507 432 27539
rect 472 27507 504 27539
rect 544 27507 576 27539
rect 616 27507 648 27539
rect 688 27507 720 27539
rect 760 27507 792 27539
rect 832 27507 864 27539
rect 904 27507 936 27539
rect 976 27507 1008 27539
rect 1048 27507 1080 27539
rect 1120 27507 1152 27539
rect 1192 27507 1224 27539
rect 1264 27507 1296 27539
rect 1336 27507 1368 27539
rect 1408 27507 1440 27539
rect 1480 27507 1512 27539
rect 1552 27507 1584 27539
rect 1624 27507 1656 27539
rect 1696 27507 1728 27539
rect 1768 27507 1800 27539
rect 1840 27507 1872 27539
rect 1912 27507 1944 27539
rect 1984 27507 2016 27539
rect 2056 27507 2088 27539
rect 2128 27507 2160 27539
rect 2200 27507 2232 27539
rect 2272 27507 2304 27539
rect 2344 27507 2376 27539
rect 2416 27507 2448 27539
rect 2488 27507 2520 27539
rect 2560 27507 2592 27539
rect 2632 27507 2664 27539
rect 2704 27507 2736 27539
rect 2776 27507 2808 27539
rect 2848 27507 2880 27539
rect 2920 27507 2952 27539
rect 2992 27507 3024 27539
rect 3064 27507 3096 27539
rect 3136 27507 3168 27539
rect 3208 27507 3240 27539
rect 3280 27507 3312 27539
rect 3352 27507 3384 27539
rect 3424 27507 3456 27539
rect 3496 27507 3528 27539
rect 3568 27507 3600 27539
rect 3640 27507 3672 27539
rect 3712 27507 3744 27539
rect 3784 27507 3816 27539
rect 3856 27507 3888 27539
rect 112 27435 144 27467
rect 184 27435 216 27467
rect 256 27435 288 27467
rect 328 27435 360 27467
rect 400 27435 432 27467
rect 472 27435 504 27467
rect 544 27435 576 27467
rect 616 27435 648 27467
rect 688 27435 720 27467
rect 760 27435 792 27467
rect 832 27435 864 27467
rect 904 27435 936 27467
rect 976 27435 1008 27467
rect 1048 27435 1080 27467
rect 1120 27435 1152 27467
rect 1192 27435 1224 27467
rect 1264 27435 1296 27467
rect 1336 27435 1368 27467
rect 1408 27435 1440 27467
rect 1480 27435 1512 27467
rect 1552 27435 1584 27467
rect 1624 27435 1656 27467
rect 1696 27435 1728 27467
rect 1768 27435 1800 27467
rect 1840 27435 1872 27467
rect 1912 27435 1944 27467
rect 1984 27435 2016 27467
rect 2056 27435 2088 27467
rect 2128 27435 2160 27467
rect 2200 27435 2232 27467
rect 2272 27435 2304 27467
rect 2344 27435 2376 27467
rect 2416 27435 2448 27467
rect 2488 27435 2520 27467
rect 2560 27435 2592 27467
rect 2632 27435 2664 27467
rect 2704 27435 2736 27467
rect 2776 27435 2808 27467
rect 2848 27435 2880 27467
rect 2920 27435 2952 27467
rect 2992 27435 3024 27467
rect 3064 27435 3096 27467
rect 3136 27435 3168 27467
rect 3208 27435 3240 27467
rect 3280 27435 3312 27467
rect 3352 27435 3384 27467
rect 3424 27435 3456 27467
rect 3496 27435 3528 27467
rect 3568 27435 3600 27467
rect 3640 27435 3672 27467
rect 3712 27435 3744 27467
rect 3784 27435 3816 27467
rect 3856 27435 3888 27467
rect 112 27363 144 27395
rect 184 27363 216 27395
rect 256 27363 288 27395
rect 328 27363 360 27395
rect 400 27363 432 27395
rect 472 27363 504 27395
rect 544 27363 576 27395
rect 616 27363 648 27395
rect 688 27363 720 27395
rect 760 27363 792 27395
rect 832 27363 864 27395
rect 904 27363 936 27395
rect 976 27363 1008 27395
rect 1048 27363 1080 27395
rect 1120 27363 1152 27395
rect 1192 27363 1224 27395
rect 1264 27363 1296 27395
rect 1336 27363 1368 27395
rect 1408 27363 1440 27395
rect 1480 27363 1512 27395
rect 1552 27363 1584 27395
rect 1624 27363 1656 27395
rect 1696 27363 1728 27395
rect 1768 27363 1800 27395
rect 1840 27363 1872 27395
rect 1912 27363 1944 27395
rect 1984 27363 2016 27395
rect 2056 27363 2088 27395
rect 2128 27363 2160 27395
rect 2200 27363 2232 27395
rect 2272 27363 2304 27395
rect 2344 27363 2376 27395
rect 2416 27363 2448 27395
rect 2488 27363 2520 27395
rect 2560 27363 2592 27395
rect 2632 27363 2664 27395
rect 2704 27363 2736 27395
rect 2776 27363 2808 27395
rect 2848 27363 2880 27395
rect 2920 27363 2952 27395
rect 2992 27363 3024 27395
rect 3064 27363 3096 27395
rect 3136 27363 3168 27395
rect 3208 27363 3240 27395
rect 3280 27363 3312 27395
rect 3352 27363 3384 27395
rect 3424 27363 3456 27395
rect 3496 27363 3528 27395
rect 3568 27363 3600 27395
rect 3640 27363 3672 27395
rect 3712 27363 3744 27395
rect 3784 27363 3816 27395
rect 3856 27363 3888 27395
rect 112 27291 144 27323
rect 184 27291 216 27323
rect 256 27291 288 27323
rect 328 27291 360 27323
rect 400 27291 432 27323
rect 472 27291 504 27323
rect 544 27291 576 27323
rect 616 27291 648 27323
rect 688 27291 720 27323
rect 760 27291 792 27323
rect 832 27291 864 27323
rect 904 27291 936 27323
rect 976 27291 1008 27323
rect 1048 27291 1080 27323
rect 1120 27291 1152 27323
rect 1192 27291 1224 27323
rect 1264 27291 1296 27323
rect 1336 27291 1368 27323
rect 1408 27291 1440 27323
rect 1480 27291 1512 27323
rect 1552 27291 1584 27323
rect 1624 27291 1656 27323
rect 1696 27291 1728 27323
rect 1768 27291 1800 27323
rect 1840 27291 1872 27323
rect 1912 27291 1944 27323
rect 1984 27291 2016 27323
rect 2056 27291 2088 27323
rect 2128 27291 2160 27323
rect 2200 27291 2232 27323
rect 2272 27291 2304 27323
rect 2344 27291 2376 27323
rect 2416 27291 2448 27323
rect 2488 27291 2520 27323
rect 2560 27291 2592 27323
rect 2632 27291 2664 27323
rect 2704 27291 2736 27323
rect 2776 27291 2808 27323
rect 2848 27291 2880 27323
rect 2920 27291 2952 27323
rect 2992 27291 3024 27323
rect 3064 27291 3096 27323
rect 3136 27291 3168 27323
rect 3208 27291 3240 27323
rect 3280 27291 3312 27323
rect 3352 27291 3384 27323
rect 3424 27291 3456 27323
rect 3496 27291 3528 27323
rect 3568 27291 3600 27323
rect 3640 27291 3672 27323
rect 3712 27291 3744 27323
rect 3784 27291 3816 27323
rect 3856 27291 3888 27323
rect 112 27219 144 27251
rect 184 27219 216 27251
rect 256 27219 288 27251
rect 328 27219 360 27251
rect 400 27219 432 27251
rect 472 27219 504 27251
rect 544 27219 576 27251
rect 616 27219 648 27251
rect 688 27219 720 27251
rect 760 27219 792 27251
rect 832 27219 864 27251
rect 904 27219 936 27251
rect 976 27219 1008 27251
rect 1048 27219 1080 27251
rect 1120 27219 1152 27251
rect 1192 27219 1224 27251
rect 1264 27219 1296 27251
rect 1336 27219 1368 27251
rect 1408 27219 1440 27251
rect 1480 27219 1512 27251
rect 1552 27219 1584 27251
rect 1624 27219 1656 27251
rect 1696 27219 1728 27251
rect 1768 27219 1800 27251
rect 1840 27219 1872 27251
rect 1912 27219 1944 27251
rect 1984 27219 2016 27251
rect 2056 27219 2088 27251
rect 2128 27219 2160 27251
rect 2200 27219 2232 27251
rect 2272 27219 2304 27251
rect 2344 27219 2376 27251
rect 2416 27219 2448 27251
rect 2488 27219 2520 27251
rect 2560 27219 2592 27251
rect 2632 27219 2664 27251
rect 2704 27219 2736 27251
rect 2776 27219 2808 27251
rect 2848 27219 2880 27251
rect 2920 27219 2952 27251
rect 2992 27219 3024 27251
rect 3064 27219 3096 27251
rect 3136 27219 3168 27251
rect 3208 27219 3240 27251
rect 3280 27219 3312 27251
rect 3352 27219 3384 27251
rect 3424 27219 3456 27251
rect 3496 27219 3528 27251
rect 3568 27219 3600 27251
rect 3640 27219 3672 27251
rect 3712 27219 3744 27251
rect 3784 27219 3816 27251
rect 3856 27219 3888 27251
rect 112 27147 144 27179
rect 184 27147 216 27179
rect 256 27147 288 27179
rect 328 27147 360 27179
rect 400 27147 432 27179
rect 472 27147 504 27179
rect 544 27147 576 27179
rect 616 27147 648 27179
rect 688 27147 720 27179
rect 760 27147 792 27179
rect 832 27147 864 27179
rect 904 27147 936 27179
rect 976 27147 1008 27179
rect 1048 27147 1080 27179
rect 1120 27147 1152 27179
rect 1192 27147 1224 27179
rect 1264 27147 1296 27179
rect 1336 27147 1368 27179
rect 1408 27147 1440 27179
rect 1480 27147 1512 27179
rect 1552 27147 1584 27179
rect 1624 27147 1656 27179
rect 1696 27147 1728 27179
rect 1768 27147 1800 27179
rect 1840 27147 1872 27179
rect 1912 27147 1944 27179
rect 1984 27147 2016 27179
rect 2056 27147 2088 27179
rect 2128 27147 2160 27179
rect 2200 27147 2232 27179
rect 2272 27147 2304 27179
rect 2344 27147 2376 27179
rect 2416 27147 2448 27179
rect 2488 27147 2520 27179
rect 2560 27147 2592 27179
rect 2632 27147 2664 27179
rect 2704 27147 2736 27179
rect 2776 27147 2808 27179
rect 2848 27147 2880 27179
rect 2920 27147 2952 27179
rect 2992 27147 3024 27179
rect 3064 27147 3096 27179
rect 3136 27147 3168 27179
rect 3208 27147 3240 27179
rect 3280 27147 3312 27179
rect 3352 27147 3384 27179
rect 3424 27147 3456 27179
rect 3496 27147 3528 27179
rect 3568 27147 3600 27179
rect 3640 27147 3672 27179
rect 3712 27147 3744 27179
rect 3784 27147 3816 27179
rect 3856 27147 3888 27179
rect 112 27075 144 27107
rect 184 27075 216 27107
rect 256 27075 288 27107
rect 328 27075 360 27107
rect 400 27075 432 27107
rect 472 27075 504 27107
rect 544 27075 576 27107
rect 616 27075 648 27107
rect 688 27075 720 27107
rect 760 27075 792 27107
rect 832 27075 864 27107
rect 904 27075 936 27107
rect 976 27075 1008 27107
rect 1048 27075 1080 27107
rect 1120 27075 1152 27107
rect 1192 27075 1224 27107
rect 1264 27075 1296 27107
rect 1336 27075 1368 27107
rect 1408 27075 1440 27107
rect 1480 27075 1512 27107
rect 1552 27075 1584 27107
rect 1624 27075 1656 27107
rect 1696 27075 1728 27107
rect 1768 27075 1800 27107
rect 1840 27075 1872 27107
rect 1912 27075 1944 27107
rect 1984 27075 2016 27107
rect 2056 27075 2088 27107
rect 2128 27075 2160 27107
rect 2200 27075 2232 27107
rect 2272 27075 2304 27107
rect 2344 27075 2376 27107
rect 2416 27075 2448 27107
rect 2488 27075 2520 27107
rect 2560 27075 2592 27107
rect 2632 27075 2664 27107
rect 2704 27075 2736 27107
rect 2776 27075 2808 27107
rect 2848 27075 2880 27107
rect 2920 27075 2952 27107
rect 2992 27075 3024 27107
rect 3064 27075 3096 27107
rect 3136 27075 3168 27107
rect 3208 27075 3240 27107
rect 3280 27075 3312 27107
rect 3352 27075 3384 27107
rect 3424 27075 3456 27107
rect 3496 27075 3528 27107
rect 3568 27075 3600 27107
rect 3640 27075 3672 27107
rect 3712 27075 3744 27107
rect 3784 27075 3816 27107
rect 3856 27075 3888 27107
rect 112 27003 144 27035
rect 184 27003 216 27035
rect 256 27003 288 27035
rect 328 27003 360 27035
rect 400 27003 432 27035
rect 472 27003 504 27035
rect 544 27003 576 27035
rect 616 27003 648 27035
rect 688 27003 720 27035
rect 760 27003 792 27035
rect 832 27003 864 27035
rect 904 27003 936 27035
rect 976 27003 1008 27035
rect 1048 27003 1080 27035
rect 1120 27003 1152 27035
rect 1192 27003 1224 27035
rect 1264 27003 1296 27035
rect 1336 27003 1368 27035
rect 1408 27003 1440 27035
rect 1480 27003 1512 27035
rect 1552 27003 1584 27035
rect 1624 27003 1656 27035
rect 1696 27003 1728 27035
rect 1768 27003 1800 27035
rect 1840 27003 1872 27035
rect 1912 27003 1944 27035
rect 1984 27003 2016 27035
rect 2056 27003 2088 27035
rect 2128 27003 2160 27035
rect 2200 27003 2232 27035
rect 2272 27003 2304 27035
rect 2344 27003 2376 27035
rect 2416 27003 2448 27035
rect 2488 27003 2520 27035
rect 2560 27003 2592 27035
rect 2632 27003 2664 27035
rect 2704 27003 2736 27035
rect 2776 27003 2808 27035
rect 2848 27003 2880 27035
rect 2920 27003 2952 27035
rect 2992 27003 3024 27035
rect 3064 27003 3096 27035
rect 3136 27003 3168 27035
rect 3208 27003 3240 27035
rect 3280 27003 3312 27035
rect 3352 27003 3384 27035
rect 3424 27003 3456 27035
rect 3496 27003 3528 27035
rect 3568 27003 3600 27035
rect 3640 27003 3672 27035
rect 3712 27003 3744 27035
rect 3784 27003 3816 27035
rect 3856 27003 3888 27035
rect 112 26931 144 26963
rect 184 26931 216 26963
rect 256 26931 288 26963
rect 328 26931 360 26963
rect 400 26931 432 26963
rect 472 26931 504 26963
rect 544 26931 576 26963
rect 616 26931 648 26963
rect 688 26931 720 26963
rect 760 26931 792 26963
rect 832 26931 864 26963
rect 904 26931 936 26963
rect 976 26931 1008 26963
rect 1048 26931 1080 26963
rect 1120 26931 1152 26963
rect 1192 26931 1224 26963
rect 1264 26931 1296 26963
rect 1336 26931 1368 26963
rect 1408 26931 1440 26963
rect 1480 26931 1512 26963
rect 1552 26931 1584 26963
rect 1624 26931 1656 26963
rect 1696 26931 1728 26963
rect 1768 26931 1800 26963
rect 1840 26931 1872 26963
rect 1912 26931 1944 26963
rect 1984 26931 2016 26963
rect 2056 26931 2088 26963
rect 2128 26931 2160 26963
rect 2200 26931 2232 26963
rect 2272 26931 2304 26963
rect 2344 26931 2376 26963
rect 2416 26931 2448 26963
rect 2488 26931 2520 26963
rect 2560 26931 2592 26963
rect 2632 26931 2664 26963
rect 2704 26931 2736 26963
rect 2776 26931 2808 26963
rect 2848 26931 2880 26963
rect 2920 26931 2952 26963
rect 2992 26931 3024 26963
rect 3064 26931 3096 26963
rect 3136 26931 3168 26963
rect 3208 26931 3240 26963
rect 3280 26931 3312 26963
rect 3352 26931 3384 26963
rect 3424 26931 3456 26963
rect 3496 26931 3528 26963
rect 3568 26931 3600 26963
rect 3640 26931 3672 26963
rect 3712 26931 3744 26963
rect 3784 26931 3816 26963
rect 3856 26931 3888 26963
rect 112 26859 144 26891
rect 184 26859 216 26891
rect 256 26859 288 26891
rect 328 26859 360 26891
rect 400 26859 432 26891
rect 472 26859 504 26891
rect 544 26859 576 26891
rect 616 26859 648 26891
rect 688 26859 720 26891
rect 760 26859 792 26891
rect 832 26859 864 26891
rect 904 26859 936 26891
rect 976 26859 1008 26891
rect 1048 26859 1080 26891
rect 1120 26859 1152 26891
rect 1192 26859 1224 26891
rect 1264 26859 1296 26891
rect 1336 26859 1368 26891
rect 1408 26859 1440 26891
rect 1480 26859 1512 26891
rect 1552 26859 1584 26891
rect 1624 26859 1656 26891
rect 1696 26859 1728 26891
rect 1768 26859 1800 26891
rect 1840 26859 1872 26891
rect 1912 26859 1944 26891
rect 1984 26859 2016 26891
rect 2056 26859 2088 26891
rect 2128 26859 2160 26891
rect 2200 26859 2232 26891
rect 2272 26859 2304 26891
rect 2344 26859 2376 26891
rect 2416 26859 2448 26891
rect 2488 26859 2520 26891
rect 2560 26859 2592 26891
rect 2632 26859 2664 26891
rect 2704 26859 2736 26891
rect 2776 26859 2808 26891
rect 2848 26859 2880 26891
rect 2920 26859 2952 26891
rect 2992 26859 3024 26891
rect 3064 26859 3096 26891
rect 3136 26859 3168 26891
rect 3208 26859 3240 26891
rect 3280 26859 3312 26891
rect 3352 26859 3384 26891
rect 3424 26859 3456 26891
rect 3496 26859 3528 26891
rect 3568 26859 3600 26891
rect 3640 26859 3672 26891
rect 3712 26859 3744 26891
rect 3784 26859 3816 26891
rect 3856 26859 3888 26891
rect 112 26787 144 26819
rect 184 26787 216 26819
rect 256 26787 288 26819
rect 328 26787 360 26819
rect 400 26787 432 26819
rect 472 26787 504 26819
rect 544 26787 576 26819
rect 616 26787 648 26819
rect 688 26787 720 26819
rect 760 26787 792 26819
rect 832 26787 864 26819
rect 904 26787 936 26819
rect 976 26787 1008 26819
rect 1048 26787 1080 26819
rect 1120 26787 1152 26819
rect 1192 26787 1224 26819
rect 1264 26787 1296 26819
rect 1336 26787 1368 26819
rect 1408 26787 1440 26819
rect 1480 26787 1512 26819
rect 1552 26787 1584 26819
rect 1624 26787 1656 26819
rect 1696 26787 1728 26819
rect 1768 26787 1800 26819
rect 1840 26787 1872 26819
rect 1912 26787 1944 26819
rect 1984 26787 2016 26819
rect 2056 26787 2088 26819
rect 2128 26787 2160 26819
rect 2200 26787 2232 26819
rect 2272 26787 2304 26819
rect 2344 26787 2376 26819
rect 2416 26787 2448 26819
rect 2488 26787 2520 26819
rect 2560 26787 2592 26819
rect 2632 26787 2664 26819
rect 2704 26787 2736 26819
rect 2776 26787 2808 26819
rect 2848 26787 2880 26819
rect 2920 26787 2952 26819
rect 2992 26787 3024 26819
rect 3064 26787 3096 26819
rect 3136 26787 3168 26819
rect 3208 26787 3240 26819
rect 3280 26787 3312 26819
rect 3352 26787 3384 26819
rect 3424 26787 3456 26819
rect 3496 26787 3528 26819
rect 3568 26787 3600 26819
rect 3640 26787 3672 26819
rect 3712 26787 3744 26819
rect 3784 26787 3816 26819
rect 3856 26787 3888 26819
rect 112 26715 144 26747
rect 184 26715 216 26747
rect 256 26715 288 26747
rect 328 26715 360 26747
rect 400 26715 432 26747
rect 472 26715 504 26747
rect 544 26715 576 26747
rect 616 26715 648 26747
rect 688 26715 720 26747
rect 760 26715 792 26747
rect 832 26715 864 26747
rect 904 26715 936 26747
rect 976 26715 1008 26747
rect 1048 26715 1080 26747
rect 1120 26715 1152 26747
rect 1192 26715 1224 26747
rect 1264 26715 1296 26747
rect 1336 26715 1368 26747
rect 1408 26715 1440 26747
rect 1480 26715 1512 26747
rect 1552 26715 1584 26747
rect 1624 26715 1656 26747
rect 1696 26715 1728 26747
rect 1768 26715 1800 26747
rect 1840 26715 1872 26747
rect 1912 26715 1944 26747
rect 1984 26715 2016 26747
rect 2056 26715 2088 26747
rect 2128 26715 2160 26747
rect 2200 26715 2232 26747
rect 2272 26715 2304 26747
rect 2344 26715 2376 26747
rect 2416 26715 2448 26747
rect 2488 26715 2520 26747
rect 2560 26715 2592 26747
rect 2632 26715 2664 26747
rect 2704 26715 2736 26747
rect 2776 26715 2808 26747
rect 2848 26715 2880 26747
rect 2920 26715 2952 26747
rect 2992 26715 3024 26747
rect 3064 26715 3096 26747
rect 3136 26715 3168 26747
rect 3208 26715 3240 26747
rect 3280 26715 3312 26747
rect 3352 26715 3384 26747
rect 3424 26715 3456 26747
rect 3496 26715 3528 26747
rect 3568 26715 3600 26747
rect 3640 26715 3672 26747
rect 3712 26715 3744 26747
rect 3784 26715 3816 26747
rect 3856 26715 3888 26747
rect 112 26643 144 26675
rect 184 26643 216 26675
rect 256 26643 288 26675
rect 328 26643 360 26675
rect 400 26643 432 26675
rect 472 26643 504 26675
rect 544 26643 576 26675
rect 616 26643 648 26675
rect 688 26643 720 26675
rect 760 26643 792 26675
rect 832 26643 864 26675
rect 904 26643 936 26675
rect 976 26643 1008 26675
rect 1048 26643 1080 26675
rect 1120 26643 1152 26675
rect 1192 26643 1224 26675
rect 1264 26643 1296 26675
rect 1336 26643 1368 26675
rect 1408 26643 1440 26675
rect 1480 26643 1512 26675
rect 1552 26643 1584 26675
rect 1624 26643 1656 26675
rect 1696 26643 1728 26675
rect 1768 26643 1800 26675
rect 1840 26643 1872 26675
rect 1912 26643 1944 26675
rect 1984 26643 2016 26675
rect 2056 26643 2088 26675
rect 2128 26643 2160 26675
rect 2200 26643 2232 26675
rect 2272 26643 2304 26675
rect 2344 26643 2376 26675
rect 2416 26643 2448 26675
rect 2488 26643 2520 26675
rect 2560 26643 2592 26675
rect 2632 26643 2664 26675
rect 2704 26643 2736 26675
rect 2776 26643 2808 26675
rect 2848 26643 2880 26675
rect 2920 26643 2952 26675
rect 2992 26643 3024 26675
rect 3064 26643 3096 26675
rect 3136 26643 3168 26675
rect 3208 26643 3240 26675
rect 3280 26643 3312 26675
rect 3352 26643 3384 26675
rect 3424 26643 3456 26675
rect 3496 26643 3528 26675
rect 3568 26643 3600 26675
rect 3640 26643 3672 26675
rect 3712 26643 3744 26675
rect 3784 26643 3816 26675
rect 3856 26643 3888 26675
rect 112 26571 144 26603
rect 184 26571 216 26603
rect 256 26571 288 26603
rect 328 26571 360 26603
rect 400 26571 432 26603
rect 472 26571 504 26603
rect 544 26571 576 26603
rect 616 26571 648 26603
rect 688 26571 720 26603
rect 760 26571 792 26603
rect 832 26571 864 26603
rect 904 26571 936 26603
rect 976 26571 1008 26603
rect 1048 26571 1080 26603
rect 1120 26571 1152 26603
rect 1192 26571 1224 26603
rect 1264 26571 1296 26603
rect 1336 26571 1368 26603
rect 1408 26571 1440 26603
rect 1480 26571 1512 26603
rect 1552 26571 1584 26603
rect 1624 26571 1656 26603
rect 1696 26571 1728 26603
rect 1768 26571 1800 26603
rect 1840 26571 1872 26603
rect 1912 26571 1944 26603
rect 1984 26571 2016 26603
rect 2056 26571 2088 26603
rect 2128 26571 2160 26603
rect 2200 26571 2232 26603
rect 2272 26571 2304 26603
rect 2344 26571 2376 26603
rect 2416 26571 2448 26603
rect 2488 26571 2520 26603
rect 2560 26571 2592 26603
rect 2632 26571 2664 26603
rect 2704 26571 2736 26603
rect 2776 26571 2808 26603
rect 2848 26571 2880 26603
rect 2920 26571 2952 26603
rect 2992 26571 3024 26603
rect 3064 26571 3096 26603
rect 3136 26571 3168 26603
rect 3208 26571 3240 26603
rect 3280 26571 3312 26603
rect 3352 26571 3384 26603
rect 3424 26571 3456 26603
rect 3496 26571 3528 26603
rect 3568 26571 3600 26603
rect 3640 26571 3672 26603
rect 3712 26571 3744 26603
rect 3784 26571 3816 26603
rect 3856 26571 3888 26603
rect 112 26499 144 26531
rect 184 26499 216 26531
rect 256 26499 288 26531
rect 328 26499 360 26531
rect 400 26499 432 26531
rect 472 26499 504 26531
rect 544 26499 576 26531
rect 616 26499 648 26531
rect 688 26499 720 26531
rect 760 26499 792 26531
rect 832 26499 864 26531
rect 904 26499 936 26531
rect 976 26499 1008 26531
rect 1048 26499 1080 26531
rect 1120 26499 1152 26531
rect 1192 26499 1224 26531
rect 1264 26499 1296 26531
rect 1336 26499 1368 26531
rect 1408 26499 1440 26531
rect 1480 26499 1512 26531
rect 1552 26499 1584 26531
rect 1624 26499 1656 26531
rect 1696 26499 1728 26531
rect 1768 26499 1800 26531
rect 1840 26499 1872 26531
rect 1912 26499 1944 26531
rect 1984 26499 2016 26531
rect 2056 26499 2088 26531
rect 2128 26499 2160 26531
rect 2200 26499 2232 26531
rect 2272 26499 2304 26531
rect 2344 26499 2376 26531
rect 2416 26499 2448 26531
rect 2488 26499 2520 26531
rect 2560 26499 2592 26531
rect 2632 26499 2664 26531
rect 2704 26499 2736 26531
rect 2776 26499 2808 26531
rect 2848 26499 2880 26531
rect 2920 26499 2952 26531
rect 2992 26499 3024 26531
rect 3064 26499 3096 26531
rect 3136 26499 3168 26531
rect 3208 26499 3240 26531
rect 3280 26499 3312 26531
rect 3352 26499 3384 26531
rect 3424 26499 3456 26531
rect 3496 26499 3528 26531
rect 3568 26499 3600 26531
rect 3640 26499 3672 26531
rect 3712 26499 3744 26531
rect 3784 26499 3816 26531
rect 3856 26499 3888 26531
rect 112 26427 144 26459
rect 184 26427 216 26459
rect 256 26427 288 26459
rect 328 26427 360 26459
rect 400 26427 432 26459
rect 472 26427 504 26459
rect 544 26427 576 26459
rect 616 26427 648 26459
rect 688 26427 720 26459
rect 760 26427 792 26459
rect 832 26427 864 26459
rect 904 26427 936 26459
rect 976 26427 1008 26459
rect 1048 26427 1080 26459
rect 1120 26427 1152 26459
rect 1192 26427 1224 26459
rect 1264 26427 1296 26459
rect 1336 26427 1368 26459
rect 1408 26427 1440 26459
rect 1480 26427 1512 26459
rect 1552 26427 1584 26459
rect 1624 26427 1656 26459
rect 1696 26427 1728 26459
rect 1768 26427 1800 26459
rect 1840 26427 1872 26459
rect 1912 26427 1944 26459
rect 1984 26427 2016 26459
rect 2056 26427 2088 26459
rect 2128 26427 2160 26459
rect 2200 26427 2232 26459
rect 2272 26427 2304 26459
rect 2344 26427 2376 26459
rect 2416 26427 2448 26459
rect 2488 26427 2520 26459
rect 2560 26427 2592 26459
rect 2632 26427 2664 26459
rect 2704 26427 2736 26459
rect 2776 26427 2808 26459
rect 2848 26427 2880 26459
rect 2920 26427 2952 26459
rect 2992 26427 3024 26459
rect 3064 26427 3096 26459
rect 3136 26427 3168 26459
rect 3208 26427 3240 26459
rect 3280 26427 3312 26459
rect 3352 26427 3384 26459
rect 3424 26427 3456 26459
rect 3496 26427 3528 26459
rect 3568 26427 3600 26459
rect 3640 26427 3672 26459
rect 3712 26427 3744 26459
rect 3784 26427 3816 26459
rect 3856 26427 3888 26459
rect 112 26355 144 26387
rect 184 26355 216 26387
rect 256 26355 288 26387
rect 328 26355 360 26387
rect 400 26355 432 26387
rect 472 26355 504 26387
rect 544 26355 576 26387
rect 616 26355 648 26387
rect 688 26355 720 26387
rect 760 26355 792 26387
rect 832 26355 864 26387
rect 904 26355 936 26387
rect 976 26355 1008 26387
rect 1048 26355 1080 26387
rect 1120 26355 1152 26387
rect 1192 26355 1224 26387
rect 1264 26355 1296 26387
rect 1336 26355 1368 26387
rect 1408 26355 1440 26387
rect 1480 26355 1512 26387
rect 1552 26355 1584 26387
rect 1624 26355 1656 26387
rect 1696 26355 1728 26387
rect 1768 26355 1800 26387
rect 1840 26355 1872 26387
rect 1912 26355 1944 26387
rect 1984 26355 2016 26387
rect 2056 26355 2088 26387
rect 2128 26355 2160 26387
rect 2200 26355 2232 26387
rect 2272 26355 2304 26387
rect 2344 26355 2376 26387
rect 2416 26355 2448 26387
rect 2488 26355 2520 26387
rect 2560 26355 2592 26387
rect 2632 26355 2664 26387
rect 2704 26355 2736 26387
rect 2776 26355 2808 26387
rect 2848 26355 2880 26387
rect 2920 26355 2952 26387
rect 2992 26355 3024 26387
rect 3064 26355 3096 26387
rect 3136 26355 3168 26387
rect 3208 26355 3240 26387
rect 3280 26355 3312 26387
rect 3352 26355 3384 26387
rect 3424 26355 3456 26387
rect 3496 26355 3528 26387
rect 3568 26355 3600 26387
rect 3640 26355 3672 26387
rect 3712 26355 3744 26387
rect 3784 26355 3816 26387
rect 3856 26355 3888 26387
rect 112 26283 144 26315
rect 184 26283 216 26315
rect 256 26283 288 26315
rect 328 26283 360 26315
rect 400 26283 432 26315
rect 472 26283 504 26315
rect 544 26283 576 26315
rect 616 26283 648 26315
rect 688 26283 720 26315
rect 760 26283 792 26315
rect 832 26283 864 26315
rect 904 26283 936 26315
rect 976 26283 1008 26315
rect 1048 26283 1080 26315
rect 1120 26283 1152 26315
rect 1192 26283 1224 26315
rect 1264 26283 1296 26315
rect 1336 26283 1368 26315
rect 1408 26283 1440 26315
rect 1480 26283 1512 26315
rect 1552 26283 1584 26315
rect 1624 26283 1656 26315
rect 1696 26283 1728 26315
rect 1768 26283 1800 26315
rect 1840 26283 1872 26315
rect 1912 26283 1944 26315
rect 1984 26283 2016 26315
rect 2056 26283 2088 26315
rect 2128 26283 2160 26315
rect 2200 26283 2232 26315
rect 2272 26283 2304 26315
rect 2344 26283 2376 26315
rect 2416 26283 2448 26315
rect 2488 26283 2520 26315
rect 2560 26283 2592 26315
rect 2632 26283 2664 26315
rect 2704 26283 2736 26315
rect 2776 26283 2808 26315
rect 2848 26283 2880 26315
rect 2920 26283 2952 26315
rect 2992 26283 3024 26315
rect 3064 26283 3096 26315
rect 3136 26283 3168 26315
rect 3208 26283 3240 26315
rect 3280 26283 3312 26315
rect 3352 26283 3384 26315
rect 3424 26283 3456 26315
rect 3496 26283 3528 26315
rect 3568 26283 3600 26315
rect 3640 26283 3672 26315
rect 3712 26283 3744 26315
rect 3784 26283 3816 26315
rect 3856 26283 3888 26315
rect 112 26211 144 26243
rect 184 26211 216 26243
rect 256 26211 288 26243
rect 328 26211 360 26243
rect 400 26211 432 26243
rect 472 26211 504 26243
rect 544 26211 576 26243
rect 616 26211 648 26243
rect 688 26211 720 26243
rect 760 26211 792 26243
rect 832 26211 864 26243
rect 904 26211 936 26243
rect 976 26211 1008 26243
rect 1048 26211 1080 26243
rect 1120 26211 1152 26243
rect 1192 26211 1224 26243
rect 1264 26211 1296 26243
rect 1336 26211 1368 26243
rect 1408 26211 1440 26243
rect 1480 26211 1512 26243
rect 1552 26211 1584 26243
rect 1624 26211 1656 26243
rect 1696 26211 1728 26243
rect 1768 26211 1800 26243
rect 1840 26211 1872 26243
rect 1912 26211 1944 26243
rect 1984 26211 2016 26243
rect 2056 26211 2088 26243
rect 2128 26211 2160 26243
rect 2200 26211 2232 26243
rect 2272 26211 2304 26243
rect 2344 26211 2376 26243
rect 2416 26211 2448 26243
rect 2488 26211 2520 26243
rect 2560 26211 2592 26243
rect 2632 26211 2664 26243
rect 2704 26211 2736 26243
rect 2776 26211 2808 26243
rect 2848 26211 2880 26243
rect 2920 26211 2952 26243
rect 2992 26211 3024 26243
rect 3064 26211 3096 26243
rect 3136 26211 3168 26243
rect 3208 26211 3240 26243
rect 3280 26211 3312 26243
rect 3352 26211 3384 26243
rect 3424 26211 3456 26243
rect 3496 26211 3528 26243
rect 3568 26211 3600 26243
rect 3640 26211 3672 26243
rect 3712 26211 3744 26243
rect 3784 26211 3816 26243
rect 3856 26211 3888 26243
rect 112 26139 144 26171
rect 184 26139 216 26171
rect 256 26139 288 26171
rect 328 26139 360 26171
rect 400 26139 432 26171
rect 472 26139 504 26171
rect 544 26139 576 26171
rect 616 26139 648 26171
rect 688 26139 720 26171
rect 760 26139 792 26171
rect 832 26139 864 26171
rect 904 26139 936 26171
rect 976 26139 1008 26171
rect 1048 26139 1080 26171
rect 1120 26139 1152 26171
rect 1192 26139 1224 26171
rect 1264 26139 1296 26171
rect 1336 26139 1368 26171
rect 1408 26139 1440 26171
rect 1480 26139 1512 26171
rect 1552 26139 1584 26171
rect 1624 26139 1656 26171
rect 1696 26139 1728 26171
rect 1768 26139 1800 26171
rect 1840 26139 1872 26171
rect 1912 26139 1944 26171
rect 1984 26139 2016 26171
rect 2056 26139 2088 26171
rect 2128 26139 2160 26171
rect 2200 26139 2232 26171
rect 2272 26139 2304 26171
rect 2344 26139 2376 26171
rect 2416 26139 2448 26171
rect 2488 26139 2520 26171
rect 2560 26139 2592 26171
rect 2632 26139 2664 26171
rect 2704 26139 2736 26171
rect 2776 26139 2808 26171
rect 2848 26139 2880 26171
rect 2920 26139 2952 26171
rect 2992 26139 3024 26171
rect 3064 26139 3096 26171
rect 3136 26139 3168 26171
rect 3208 26139 3240 26171
rect 3280 26139 3312 26171
rect 3352 26139 3384 26171
rect 3424 26139 3456 26171
rect 3496 26139 3528 26171
rect 3568 26139 3600 26171
rect 3640 26139 3672 26171
rect 3712 26139 3744 26171
rect 3784 26139 3816 26171
rect 3856 26139 3888 26171
rect 112 26067 144 26099
rect 184 26067 216 26099
rect 256 26067 288 26099
rect 328 26067 360 26099
rect 400 26067 432 26099
rect 472 26067 504 26099
rect 544 26067 576 26099
rect 616 26067 648 26099
rect 688 26067 720 26099
rect 760 26067 792 26099
rect 832 26067 864 26099
rect 904 26067 936 26099
rect 976 26067 1008 26099
rect 1048 26067 1080 26099
rect 1120 26067 1152 26099
rect 1192 26067 1224 26099
rect 1264 26067 1296 26099
rect 1336 26067 1368 26099
rect 1408 26067 1440 26099
rect 1480 26067 1512 26099
rect 1552 26067 1584 26099
rect 1624 26067 1656 26099
rect 1696 26067 1728 26099
rect 1768 26067 1800 26099
rect 1840 26067 1872 26099
rect 1912 26067 1944 26099
rect 1984 26067 2016 26099
rect 2056 26067 2088 26099
rect 2128 26067 2160 26099
rect 2200 26067 2232 26099
rect 2272 26067 2304 26099
rect 2344 26067 2376 26099
rect 2416 26067 2448 26099
rect 2488 26067 2520 26099
rect 2560 26067 2592 26099
rect 2632 26067 2664 26099
rect 2704 26067 2736 26099
rect 2776 26067 2808 26099
rect 2848 26067 2880 26099
rect 2920 26067 2952 26099
rect 2992 26067 3024 26099
rect 3064 26067 3096 26099
rect 3136 26067 3168 26099
rect 3208 26067 3240 26099
rect 3280 26067 3312 26099
rect 3352 26067 3384 26099
rect 3424 26067 3456 26099
rect 3496 26067 3528 26099
rect 3568 26067 3600 26099
rect 3640 26067 3672 26099
rect 3712 26067 3744 26099
rect 3784 26067 3816 26099
rect 3856 26067 3888 26099
rect 112 25995 144 26027
rect 184 25995 216 26027
rect 256 25995 288 26027
rect 328 25995 360 26027
rect 400 25995 432 26027
rect 472 25995 504 26027
rect 544 25995 576 26027
rect 616 25995 648 26027
rect 688 25995 720 26027
rect 760 25995 792 26027
rect 832 25995 864 26027
rect 904 25995 936 26027
rect 976 25995 1008 26027
rect 1048 25995 1080 26027
rect 1120 25995 1152 26027
rect 1192 25995 1224 26027
rect 1264 25995 1296 26027
rect 1336 25995 1368 26027
rect 1408 25995 1440 26027
rect 1480 25995 1512 26027
rect 1552 25995 1584 26027
rect 1624 25995 1656 26027
rect 1696 25995 1728 26027
rect 1768 25995 1800 26027
rect 1840 25995 1872 26027
rect 1912 25995 1944 26027
rect 1984 25995 2016 26027
rect 2056 25995 2088 26027
rect 2128 25995 2160 26027
rect 2200 25995 2232 26027
rect 2272 25995 2304 26027
rect 2344 25995 2376 26027
rect 2416 25995 2448 26027
rect 2488 25995 2520 26027
rect 2560 25995 2592 26027
rect 2632 25995 2664 26027
rect 2704 25995 2736 26027
rect 2776 25995 2808 26027
rect 2848 25995 2880 26027
rect 2920 25995 2952 26027
rect 2992 25995 3024 26027
rect 3064 25995 3096 26027
rect 3136 25995 3168 26027
rect 3208 25995 3240 26027
rect 3280 25995 3312 26027
rect 3352 25995 3384 26027
rect 3424 25995 3456 26027
rect 3496 25995 3528 26027
rect 3568 25995 3600 26027
rect 3640 25995 3672 26027
rect 3712 25995 3744 26027
rect 3784 25995 3816 26027
rect 3856 25995 3888 26027
rect 112 25923 144 25955
rect 184 25923 216 25955
rect 256 25923 288 25955
rect 328 25923 360 25955
rect 400 25923 432 25955
rect 472 25923 504 25955
rect 544 25923 576 25955
rect 616 25923 648 25955
rect 688 25923 720 25955
rect 760 25923 792 25955
rect 832 25923 864 25955
rect 904 25923 936 25955
rect 976 25923 1008 25955
rect 1048 25923 1080 25955
rect 1120 25923 1152 25955
rect 1192 25923 1224 25955
rect 1264 25923 1296 25955
rect 1336 25923 1368 25955
rect 1408 25923 1440 25955
rect 1480 25923 1512 25955
rect 1552 25923 1584 25955
rect 1624 25923 1656 25955
rect 1696 25923 1728 25955
rect 1768 25923 1800 25955
rect 1840 25923 1872 25955
rect 1912 25923 1944 25955
rect 1984 25923 2016 25955
rect 2056 25923 2088 25955
rect 2128 25923 2160 25955
rect 2200 25923 2232 25955
rect 2272 25923 2304 25955
rect 2344 25923 2376 25955
rect 2416 25923 2448 25955
rect 2488 25923 2520 25955
rect 2560 25923 2592 25955
rect 2632 25923 2664 25955
rect 2704 25923 2736 25955
rect 2776 25923 2808 25955
rect 2848 25923 2880 25955
rect 2920 25923 2952 25955
rect 2992 25923 3024 25955
rect 3064 25923 3096 25955
rect 3136 25923 3168 25955
rect 3208 25923 3240 25955
rect 3280 25923 3312 25955
rect 3352 25923 3384 25955
rect 3424 25923 3456 25955
rect 3496 25923 3528 25955
rect 3568 25923 3600 25955
rect 3640 25923 3672 25955
rect 3712 25923 3744 25955
rect 3784 25923 3816 25955
rect 3856 25923 3888 25955
rect 112 25851 144 25883
rect 184 25851 216 25883
rect 256 25851 288 25883
rect 328 25851 360 25883
rect 400 25851 432 25883
rect 472 25851 504 25883
rect 544 25851 576 25883
rect 616 25851 648 25883
rect 688 25851 720 25883
rect 760 25851 792 25883
rect 832 25851 864 25883
rect 904 25851 936 25883
rect 976 25851 1008 25883
rect 1048 25851 1080 25883
rect 1120 25851 1152 25883
rect 1192 25851 1224 25883
rect 1264 25851 1296 25883
rect 1336 25851 1368 25883
rect 1408 25851 1440 25883
rect 1480 25851 1512 25883
rect 1552 25851 1584 25883
rect 1624 25851 1656 25883
rect 1696 25851 1728 25883
rect 1768 25851 1800 25883
rect 1840 25851 1872 25883
rect 1912 25851 1944 25883
rect 1984 25851 2016 25883
rect 2056 25851 2088 25883
rect 2128 25851 2160 25883
rect 2200 25851 2232 25883
rect 2272 25851 2304 25883
rect 2344 25851 2376 25883
rect 2416 25851 2448 25883
rect 2488 25851 2520 25883
rect 2560 25851 2592 25883
rect 2632 25851 2664 25883
rect 2704 25851 2736 25883
rect 2776 25851 2808 25883
rect 2848 25851 2880 25883
rect 2920 25851 2952 25883
rect 2992 25851 3024 25883
rect 3064 25851 3096 25883
rect 3136 25851 3168 25883
rect 3208 25851 3240 25883
rect 3280 25851 3312 25883
rect 3352 25851 3384 25883
rect 3424 25851 3456 25883
rect 3496 25851 3528 25883
rect 3568 25851 3600 25883
rect 3640 25851 3672 25883
rect 3712 25851 3744 25883
rect 3784 25851 3816 25883
rect 3856 25851 3888 25883
rect 112 25779 144 25811
rect 184 25779 216 25811
rect 256 25779 288 25811
rect 328 25779 360 25811
rect 400 25779 432 25811
rect 472 25779 504 25811
rect 544 25779 576 25811
rect 616 25779 648 25811
rect 688 25779 720 25811
rect 760 25779 792 25811
rect 832 25779 864 25811
rect 904 25779 936 25811
rect 976 25779 1008 25811
rect 1048 25779 1080 25811
rect 1120 25779 1152 25811
rect 1192 25779 1224 25811
rect 1264 25779 1296 25811
rect 1336 25779 1368 25811
rect 1408 25779 1440 25811
rect 1480 25779 1512 25811
rect 1552 25779 1584 25811
rect 1624 25779 1656 25811
rect 1696 25779 1728 25811
rect 1768 25779 1800 25811
rect 1840 25779 1872 25811
rect 1912 25779 1944 25811
rect 1984 25779 2016 25811
rect 2056 25779 2088 25811
rect 2128 25779 2160 25811
rect 2200 25779 2232 25811
rect 2272 25779 2304 25811
rect 2344 25779 2376 25811
rect 2416 25779 2448 25811
rect 2488 25779 2520 25811
rect 2560 25779 2592 25811
rect 2632 25779 2664 25811
rect 2704 25779 2736 25811
rect 2776 25779 2808 25811
rect 2848 25779 2880 25811
rect 2920 25779 2952 25811
rect 2992 25779 3024 25811
rect 3064 25779 3096 25811
rect 3136 25779 3168 25811
rect 3208 25779 3240 25811
rect 3280 25779 3312 25811
rect 3352 25779 3384 25811
rect 3424 25779 3456 25811
rect 3496 25779 3528 25811
rect 3568 25779 3600 25811
rect 3640 25779 3672 25811
rect 3712 25779 3744 25811
rect 3784 25779 3816 25811
rect 3856 25779 3888 25811
rect 112 25707 144 25739
rect 184 25707 216 25739
rect 256 25707 288 25739
rect 328 25707 360 25739
rect 400 25707 432 25739
rect 472 25707 504 25739
rect 544 25707 576 25739
rect 616 25707 648 25739
rect 688 25707 720 25739
rect 760 25707 792 25739
rect 832 25707 864 25739
rect 904 25707 936 25739
rect 976 25707 1008 25739
rect 1048 25707 1080 25739
rect 1120 25707 1152 25739
rect 1192 25707 1224 25739
rect 1264 25707 1296 25739
rect 1336 25707 1368 25739
rect 1408 25707 1440 25739
rect 1480 25707 1512 25739
rect 1552 25707 1584 25739
rect 1624 25707 1656 25739
rect 1696 25707 1728 25739
rect 1768 25707 1800 25739
rect 1840 25707 1872 25739
rect 1912 25707 1944 25739
rect 1984 25707 2016 25739
rect 2056 25707 2088 25739
rect 2128 25707 2160 25739
rect 2200 25707 2232 25739
rect 2272 25707 2304 25739
rect 2344 25707 2376 25739
rect 2416 25707 2448 25739
rect 2488 25707 2520 25739
rect 2560 25707 2592 25739
rect 2632 25707 2664 25739
rect 2704 25707 2736 25739
rect 2776 25707 2808 25739
rect 2848 25707 2880 25739
rect 2920 25707 2952 25739
rect 2992 25707 3024 25739
rect 3064 25707 3096 25739
rect 3136 25707 3168 25739
rect 3208 25707 3240 25739
rect 3280 25707 3312 25739
rect 3352 25707 3384 25739
rect 3424 25707 3456 25739
rect 3496 25707 3528 25739
rect 3568 25707 3600 25739
rect 3640 25707 3672 25739
rect 3712 25707 3744 25739
rect 3784 25707 3816 25739
rect 3856 25707 3888 25739
rect 112 25635 144 25667
rect 184 25635 216 25667
rect 256 25635 288 25667
rect 328 25635 360 25667
rect 400 25635 432 25667
rect 472 25635 504 25667
rect 544 25635 576 25667
rect 616 25635 648 25667
rect 688 25635 720 25667
rect 760 25635 792 25667
rect 832 25635 864 25667
rect 904 25635 936 25667
rect 976 25635 1008 25667
rect 1048 25635 1080 25667
rect 1120 25635 1152 25667
rect 1192 25635 1224 25667
rect 1264 25635 1296 25667
rect 1336 25635 1368 25667
rect 1408 25635 1440 25667
rect 1480 25635 1512 25667
rect 1552 25635 1584 25667
rect 1624 25635 1656 25667
rect 1696 25635 1728 25667
rect 1768 25635 1800 25667
rect 1840 25635 1872 25667
rect 1912 25635 1944 25667
rect 1984 25635 2016 25667
rect 2056 25635 2088 25667
rect 2128 25635 2160 25667
rect 2200 25635 2232 25667
rect 2272 25635 2304 25667
rect 2344 25635 2376 25667
rect 2416 25635 2448 25667
rect 2488 25635 2520 25667
rect 2560 25635 2592 25667
rect 2632 25635 2664 25667
rect 2704 25635 2736 25667
rect 2776 25635 2808 25667
rect 2848 25635 2880 25667
rect 2920 25635 2952 25667
rect 2992 25635 3024 25667
rect 3064 25635 3096 25667
rect 3136 25635 3168 25667
rect 3208 25635 3240 25667
rect 3280 25635 3312 25667
rect 3352 25635 3384 25667
rect 3424 25635 3456 25667
rect 3496 25635 3528 25667
rect 3568 25635 3600 25667
rect 3640 25635 3672 25667
rect 3712 25635 3744 25667
rect 3784 25635 3816 25667
rect 3856 25635 3888 25667
rect 112 25563 144 25595
rect 184 25563 216 25595
rect 256 25563 288 25595
rect 328 25563 360 25595
rect 400 25563 432 25595
rect 472 25563 504 25595
rect 544 25563 576 25595
rect 616 25563 648 25595
rect 688 25563 720 25595
rect 760 25563 792 25595
rect 832 25563 864 25595
rect 904 25563 936 25595
rect 976 25563 1008 25595
rect 1048 25563 1080 25595
rect 1120 25563 1152 25595
rect 1192 25563 1224 25595
rect 1264 25563 1296 25595
rect 1336 25563 1368 25595
rect 1408 25563 1440 25595
rect 1480 25563 1512 25595
rect 1552 25563 1584 25595
rect 1624 25563 1656 25595
rect 1696 25563 1728 25595
rect 1768 25563 1800 25595
rect 1840 25563 1872 25595
rect 1912 25563 1944 25595
rect 1984 25563 2016 25595
rect 2056 25563 2088 25595
rect 2128 25563 2160 25595
rect 2200 25563 2232 25595
rect 2272 25563 2304 25595
rect 2344 25563 2376 25595
rect 2416 25563 2448 25595
rect 2488 25563 2520 25595
rect 2560 25563 2592 25595
rect 2632 25563 2664 25595
rect 2704 25563 2736 25595
rect 2776 25563 2808 25595
rect 2848 25563 2880 25595
rect 2920 25563 2952 25595
rect 2992 25563 3024 25595
rect 3064 25563 3096 25595
rect 3136 25563 3168 25595
rect 3208 25563 3240 25595
rect 3280 25563 3312 25595
rect 3352 25563 3384 25595
rect 3424 25563 3456 25595
rect 3496 25563 3528 25595
rect 3568 25563 3600 25595
rect 3640 25563 3672 25595
rect 3712 25563 3744 25595
rect 3784 25563 3816 25595
rect 3856 25563 3888 25595
rect 112 25491 144 25523
rect 184 25491 216 25523
rect 256 25491 288 25523
rect 328 25491 360 25523
rect 400 25491 432 25523
rect 472 25491 504 25523
rect 544 25491 576 25523
rect 616 25491 648 25523
rect 688 25491 720 25523
rect 760 25491 792 25523
rect 832 25491 864 25523
rect 904 25491 936 25523
rect 976 25491 1008 25523
rect 1048 25491 1080 25523
rect 1120 25491 1152 25523
rect 1192 25491 1224 25523
rect 1264 25491 1296 25523
rect 1336 25491 1368 25523
rect 1408 25491 1440 25523
rect 1480 25491 1512 25523
rect 1552 25491 1584 25523
rect 1624 25491 1656 25523
rect 1696 25491 1728 25523
rect 1768 25491 1800 25523
rect 1840 25491 1872 25523
rect 1912 25491 1944 25523
rect 1984 25491 2016 25523
rect 2056 25491 2088 25523
rect 2128 25491 2160 25523
rect 2200 25491 2232 25523
rect 2272 25491 2304 25523
rect 2344 25491 2376 25523
rect 2416 25491 2448 25523
rect 2488 25491 2520 25523
rect 2560 25491 2592 25523
rect 2632 25491 2664 25523
rect 2704 25491 2736 25523
rect 2776 25491 2808 25523
rect 2848 25491 2880 25523
rect 2920 25491 2952 25523
rect 2992 25491 3024 25523
rect 3064 25491 3096 25523
rect 3136 25491 3168 25523
rect 3208 25491 3240 25523
rect 3280 25491 3312 25523
rect 3352 25491 3384 25523
rect 3424 25491 3456 25523
rect 3496 25491 3528 25523
rect 3568 25491 3600 25523
rect 3640 25491 3672 25523
rect 3712 25491 3744 25523
rect 3784 25491 3816 25523
rect 3856 25491 3888 25523
rect 112 25419 144 25451
rect 184 25419 216 25451
rect 256 25419 288 25451
rect 328 25419 360 25451
rect 400 25419 432 25451
rect 472 25419 504 25451
rect 544 25419 576 25451
rect 616 25419 648 25451
rect 688 25419 720 25451
rect 760 25419 792 25451
rect 832 25419 864 25451
rect 904 25419 936 25451
rect 976 25419 1008 25451
rect 1048 25419 1080 25451
rect 1120 25419 1152 25451
rect 1192 25419 1224 25451
rect 1264 25419 1296 25451
rect 1336 25419 1368 25451
rect 1408 25419 1440 25451
rect 1480 25419 1512 25451
rect 1552 25419 1584 25451
rect 1624 25419 1656 25451
rect 1696 25419 1728 25451
rect 1768 25419 1800 25451
rect 1840 25419 1872 25451
rect 1912 25419 1944 25451
rect 1984 25419 2016 25451
rect 2056 25419 2088 25451
rect 2128 25419 2160 25451
rect 2200 25419 2232 25451
rect 2272 25419 2304 25451
rect 2344 25419 2376 25451
rect 2416 25419 2448 25451
rect 2488 25419 2520 25451
rect 2560 25419 2592 25451
rect 2632 25419 2664 25451
rect 2704 25419 2736 25451
rect 2776 25419 2808 25451
rect 2848 25419 2880 25451
rect 2920 25419 2952 25451
rect 2992 25419 3024 25451
rect 3064 25419 3096 25451
rect 3136 25419 3168 25451
rect 3208 25419 3240 25451
rect 3280 25419 3312 25451
rect 3352 25419 3384 25451
rect 3424 25419 3456 25451
rect 3496 25419 3528 25451
rect 3568 25419 3600 25451
rect 3640 25419 3672 25451
rect 3712 25419 3744 25451
rect 3784 25419 3816 25451
rect 3856 25419 3888 25451
rect 112 25347 144 25379
rect 184 25347 216 25379
rect 256 25347 288 25379
rect 328 25347 360 25379
rect 400 25347 432 25379
rect 472 25347 504 25379
rect 544 25347 576 25379
rect 616 25347 648 25379
rect 688 25347 720 25379
rect 760 25347 792 25379
rect 832 25347 864 25379
rect 904 25347 936 25379
rect 976 25347 1008 25379
rect 1048 25347 1080 25379
rect 1120 25347 1152 25379
rect 1192 25347 1224 25379
rect 1264 25347 1296 25379
rect 1336 25347 1368 25379
rect 1408 25347 1440 25379
rect 1480 25347 1512 25379
rect 1552 25347 1584 25379
rect 1624 25347 1656 25379
rect 1696 25347 1728 25379
rect 1768 25347 1800 25379
rect 1840 25347 1872 25379
rect 1912 25347 1944 25379
rect 1984 25347 2016 25379
rect 2056 25347 2088 25379
rect 2128 25347 2160 25379
rect 2200 25347 2232 25379
rect 2272 25347 2304 25379
rect 2344 25347 2376 25379
rect 2416 25347 2448 25379
rect 2488 25347 2520 25379
rect 2560 25347 2592 25379
rect 2632 25347 2664 25379
rect 2704 25347 2736 25379
rect 2776 25347 2808 25379
rect 2848 25347 2880 25379
rect 2920 25347 2952 25379
rect 2992 25347 3024 25379
rect 3064 25347 3096 25379
rect 3136 25347 3168 25379
rect 3208 25347 3240 25379
rect 3280 25347 3312 25379
rect 3352 25347 3384 25379
rect 3424 25347 3456 25379
rect 3496 25347 3528 25379
rect 3568 25347 3600 25379
rect 3640 25347 3672 25379
rect 3712 25347 3744 25379
rect 3784 25347 3816 25379
rect 3856 25347 3888 25379
rect 112 25275 144 25307
rect 184 25275 216 25307
rect 256 25275 288 25307
rect 328 25275 360 25307
rect 400 25275 432 25307
rect 472 25275 504 25307
rect 544 25275 576 25307
rect 616 25275 648 25307
rect 688 25275 720 25307
rect 760 25275 792 25307
rect 832 25275 864 25307
rect 904 25275 936 25307
rect 976 25275 1008 25307
rect 1048 25275 1080 25307
rect 1120 25275 1152 25307
rect 1192 25275 1224 25307
rect 1264 25275 1296 25307
rect 1336 25275 1368 25307
rect 1408 25275 1440 25307
rect 1480 25275 1512 25307
rect 1552 25275 1584 25307
rect 1624 25275 1656 25307
rect 1696 25275 1728 25307
rect 1768 25275 1800 25307
rect 1840 25275 1872 25307
rect 1912 25275 1944 25307
rect 1984 25275 2016 25307
rect 2056 25275 2088 25307
rect 2128 25275 2160 25307
rect 2200 25275 2232 25307
rect 2272 25275 2304 25307
rect 2344 25275 2376 25307
rect 2416 25275 2448 25307
rect 2488 25275 2520 25307
rect 2560 25275 2592 25307
rect 2632 25275 2664 25307
rect 2704 25275 2736 25307
rect 2776 25275 2808 25307
rect 2848 25275 2880 25307
rect 2920 25275 2952 25307
rect 2992 25275 3024 25307
rect 3064 25275 3096 25307
rect 3136 25275 3168 25307
rect 3208 25275 3240 25307
rect 3280 25275 3312 25307
rect 3352 25275 3384 25307
rect 3424 25275 3456 25307
rect 3496 25275 3528 25307
rect 3568 25275 3600 25307
rect 3640 25275 3672 25307
rect 3712 25275 3744 25307
rect 3784 25275 3816 25307
rect 3856 25275 3888 25307
rect 112 25203 144 25235
rect 184 25203 216 25235
rect 256 25203 288 25235
rect 328 25203 360 25235
rect 400 25203 432 25235
rect 472 25203 504 25235
rect 544 25203 576 25235
rect 616 25203 648 25235
rect 688 25203 720 25235
rect 760 25203 792 25235
rect 832 25203 864 25235
rect 904 25203 936 25235
rect 976 25203 1008 25235
rect 1048 25203 1080 25235
rect 1120 25203 1152 25235
rect 1192 25203 1224 25235
rect 1264 25203 1296 25235
rect 1336 25203 1368 25235
rect 1408 25203 1440 25235
rect 1480 25203 1512 25235
rect 1552 25203 1584 25235
rect 1624 25203 1656 25235
rect 1696 25203 1728 25235
rect 1768 25203 1800 25235
rect 1840 25203 1872 25235
rect 1912 25203 1944 25235
rect 1984 25203 2016 25235
rect 2056 25203 2088 25235
rect 2128 25203 2160 25235
rect 2200 25203 2232 25235
rect 2272 25203 2304 25235
rect 2344 25203 2376 25235
rect 2416 25203 2448 25235
rect 2488 25203 2520 25235
rect 2560 25203 2592 25235
rect 2632 25203 2664 25235
rect 2704 25203 2736 25235
rect 2776 25203 2808 25235
rect 2848 25203 2880 25235
rect 2920 25203 2952 25235
rect 2992 25203 3024 25235
rect 3064 25203 3096 25235
rect 3136 25203 3168 25235
rect 3208 25203 3240 25235
rect 3280 25203 3312 25235
rect 3352 25203 3384 25235
rect 3424 25203 3456 25235
rect 3496 25203 3528 25235
rect 3568 25203 3600 25235
rect 3640 25203 3672 25235
rect 3712 25203 3744 25235
rect 3784 25203 3816 25235
rect 3856 25203 3888 25235
rect 112 25131 144 25163
rect 184 25131 216 25163
rect 256 25131 288 25163
rect 328 25131 360 25163
rect 400 25131 432 25163
rect 472 25131 504 25163
rect 544 25131 576 25163
rect 616 25131 648 25163
rect 688 25131 720 25163
rect 760 25131 792 25163
rect 832 25131 864 25163
rect 904 25131 936 25163
rect 976 25131 1008 25163
rect 1048 25131 1080 25163
rect 1120 25131 1152 25163
rect 1192 25131 1224 25163
rect 1264 25131 1296 25163
rect 1336 25131 1368 25163
rect 1408 25131 1440 25163
rect 1480 25131 1512 25163
rect 1552 25131 1584 25163
rect 1624 25131 1656 25163
rect 1696 25131 1728 25163
rect 1768 25131 1800 25163
rect 1840 25131 1872 25163
rect 1912 25131 1944 25163
rect 1984 25131 2016 25163
rect 2056 25131 2088 25163
rect 2128 25131 2160 25163
rect 2200 25131 2232 25163
rect 2272 25131 2304 25163
rect 2344 25131 2376 25163
rect 2416 25131 2448 25163
rect 2488 25131 2520 25163
rect 2560 25131 2592 25163
rect 2632 25131 2664 25163
rect 2704 25131 2736 25163
rect 2776 25131 2808 25163
rect 2848 25131 2880 25163
rect 2920 25131 2952 25163
rect 2992 25131 3024 25163
rect 3064 25131 3096 25163
rect 3136 25131 3168 25163
rect 3208 25131 3240 25163
rect 3280 25131 3312 25163
rect 3352 25131 3384 25163
rect 3424 25131 3456 25163
rect 3496 25131 3528 25163
rect 3568 25131 3600 25163
rect 3640 25131 3672 25163
rect 3712 25131 3744 25163
rect 3784 25131 3816 25163
rect 3856 25131 3888 25163
rect 112 25059 144 25091
rect 184 25059 216 25091
rect 256 25059 288 25091
rect 328 25059 360 25091
rect 400 25059 432 25091
rect 472 25059 504 25091
rect 544 25059 576 25091
rect 616 25059 648 25091
rect 688 25059 720 25091
rect 760 25059 792 25091
rect 832 25059 864 25091
rect 904 25059 936 25091
rect 976 25059 1008 25091
rect 1048 25059 1080 25091
rect 1120 25059 1152 25091
rect 1192 25059 1224 25091
rect 1264 25059 1296 25091
rect 1336 25059 1368 25091
rect 1408 25059 1440 25091
rect 1480 25059 1512 25091
rect 1552 25059 1584 25091
rect 1624 25059 1656 25091
rect 1696 25059 1728 25091
rect 1768 25059 1800 25091
rect 1840 25059 1872 25091
rect 1912 25059 1944 25091
rect 1984 25059 2016 25091
rect 2056 25059 2088 25091
rect 2128 25059 2160 25091
rect 2200 25059 2232 25091
rect 2272 25059 2304 25091
rect 2344 25059 2376 25091
rect 2416 25059 2448 25091
rect 2488 25059 2520 25091
rect 2560 25059 2592 25091
rect 2632 25059 2664 25091
rect 2704 25059 2736 25091
rect 2776 25059 2808 25091
rect 2848 25059 2880 25091
rect 2920 25059 2952 25091
rect 2992 25059 3024 25091
rect 3064 25059 3096 25091
rect 3136 25059 3168 25091
rect 3208 25059 3240 25091
rect 3280 25059 3312 25091
rect 3352 25059 3384 25091
rect 3424 25059 3456 25091
rect 3496 25059 3528 25091
rect 3568 25059 3600 25091
rect 3640 25059 3672 25091
rect 3712 25059 3744 25091
rect 3784 25059 3816 25091
rect 3856 25059 3888 25091
rect 112 24987 144 25019
rect 184 24987 216 25019
rect 256 24987 288 25019
rect 328 24987 360 25019
rect 400 24987 432 25019
rect 472 24987 504 25019
rect 544 24987 576 25019
rect 616 24987 648 25019
rect 688 24987 720 25019
rect 760 24987 792 25019
rect 832 24987 864 25019
rect 904 24987 936 25019
rect 976 24987 1008 25019
rect 1048 24987 1080 25019
rect 1120 24987 1152 25019
rect 1192 24987 1224 25019
rect 1264 24987 1296 25019
rect 1336 24987 1368 25019
rect 1408 24987 1440 25019
rect 1480 24987 1512 25019
rect 1552 24987 1584 25019
rect 1624 24987 1656 25019
rect 1696 24987 1728 25019
rect 1768 24987 1800 25019
rect 1840 24987 1872 25019
rect 1912 24987 1944 25019
rect 1984 24987 2016 25019
rect 2056 24987 2088 25019
rect 2128 24987 2160 25019
rect 2200 24987 2232 25019
rect 2272 24987 2304 25019
rect 2344 24987 2376 25019
rect 2416 24987 2448 25019
rect 2488 24987 2520 25019
rect 2560 24987 2592 25019
rect 2632 24987 2664 25019
rect 2704 24987 2736 25019
rect 2776 24987 2808 25019
rect 2848 24987 2880 25019
rect 2920 24987 2952 25019
rect 2992 24987 3024 25019
rect 3064 24987 3096 25019
rect 3136 24987 3168 25019
rect 3208 24987 3240 25019
rect 3280 24987 3312 25019
rect 3352 24987 3384 25019
rect 3424 24987 3456 25019
rect 3496 24987 3528 25019
rect 3568 24987 3600 25019
rect 3640 24987 3672 25019
rect 3712 24987 3744 25019
rect 3784 24987 3816 25019
rect 3856 24987 3888 25019
rect 112 24915 144 24947
rect 184 24915 216 24947
rect 256 24915 288 24947
rect 328 24915 360 24947
rect 400 24915 432 24947
rect 472 24915 504 24947
rect 544 24915 576 24947
rect 616 24915 648 24947
rect 688 24915 720 24947
rect 760 24915 792 24947
rect 832 24915 864 24947
rect 904 24915 936 24947
rect 976 24915 1008 24947
rect 1048 24915 1080 24947
rect 1120 24915 1152 24947
rect 1192 24915 1224 24947
rect 1264 24915 1296 24947
rect 1336 24915 1368 24947
rect 1408 24915 1440 24947
rect 1480 24915 1512 24947
rect 1552 24915 1584 24947
rect 1624 24915 1656 24947
rect 1696 24915 1728 24947
rect 1768 24915 1800 24947
rect 1840 24915 1872 24947
rect 1912 24915 1944 24947
rect 1984 24915 2016 24947
rect 2056 24915 2088 24947
rect 2128 24915 2160 24947
rect 2200 24915 2232 24947
rect 2272 24915 2304 24947
rect 2344 24915 2376 24947
rect 2416 24915 2448 24947
rect 2488 24915 2520 24947
rect 2560 24915 2592 24947
rect 2632 24915 2664 24947
rect 2704 24915 2736 24947
rect 2776 24915 2808 24947
rect 2848 24915 2880 24947
rect 2920 24915 2952 24947
rect 2992 24915 3024 24947
rect 3064 24915 3096 24947
rect 3136 24915 3168 24947
rect 3208 24915 3240 24947
rect 3280 24915 3312 24947
rect 3352 24915 3384 24947
rect 3424 24915 3456 24947
rect 3496 24915 3528 24947
rect 3568 24915 3600 24947
rect 3640 24915 3672 24947
rect 3712 24915 3744 24947
rect 3784 24915 3816 24947
rect 3856 24915 3888 24947
rect 112 24843 144 24875
rect 184 24843 216 24875
rect 256 24843 288 24875
rect 328 24843 360 24875
rect 400 24843 432 24875
rect 472 24843 504 24875
rect 544 24843 576 24875
rect 616 24843 648 24875
rect 688 24843 720 24875
rect 760 24843 792 24875
rect 832 24843 864 24875
rect 904 24843 936 24875
rect 976 24843 1008 24875
rect 1048 24843 1080 24875
rect 1120 24843 1152 24875
rect 1192 24843 1224 24875
rect 1264 24843 1296 24875
rect 1336 24843 1368 24875
rect 1408 24843 1440 24875
rect 1480 24843 1512 24875
rect 1552 24843 1584 24875
rect 1624 24843 1656 24875
rect 1696 24843 1728 24875
rect 1768 24843 1800 24875
rect 1840 24843 1872 24875
rect 1912 24843 1944 24875
rect 1984 24843 2016 24875
rect 2056 24843 2088 24875
rect 2128 24843 2160 24875
rect 2200 24843 2232 24875
rect 2272 24843 2304 24875
rect 2344 24843 2376 24875
rect 2416 24843 2448 24875
rect 2488 24843 2520 24875
rect 2560 24843 2592 24875
rect 2632 24843 2664 24875
rect 2704 24843 2736 24875
rect 2776 24843 2808 24875
rect 2848 24843 2880 24875
rect 2920 24843 2952 24875
rect 2992 24843 3024 24875
rect 3064 24843 3096 24875
rect 3136 24843 3168 24875
rect 3208 24843 3240 24875
rect 3280 24843 3312 24875
rect 3352 24843 3384 24875
rect 3424 24843 3456 24875
rect 3496 24843 3528 24875
rect 3568 24843 3600 24875
rect 3640 24843 3672 24875
rect 3712 24843 3744 24875
rect 3784 24843 3816 24875
rect 3856 24843 3888 24875
rect 112 24771 144 24803
rect 184 24771 216 24803
rect 256 24771 288 24803
rect 328 24771 360 24803
rect 400 24771 432 24803
rect 472 24771 504 24803
rect 544 24771 576 24803
rect 616 24771 648 24803
rect 688 24771 720 24803
rect 760 24771 792 24803
rect 832 24771 864 24803
rect 904 24771 936 24803
rect 976 24771 1008 24803
rect 1048 24771 1080 24803
rect 1120 24771 1152 24803
rect 1192 24771 1224 24803
rect 1264 24771 1296 24803
rect 1336 24771 1368 24803
rect 1408 24771 1440 24803
rect 1480 24771 1512 24803
rect 1552 24771 1584 24803
rect 1624 24771 1656 24803
rect 1696 24771 1728 24803
rect 1768 24771 1800 24803
rect 1840 24771 1872 24803
rect 1912 24771 1944 24803
rect 1984 24771 2016 24803
rect 2056 24771 2088 24803
rect 2128 24771 2160 24803
rect 2200 24771 2232 24803
rect 2272 24771 2304 24803
rect 2344 24771 2376 24803
rect 2416 24771 2448 24803
rect 2488 24771 2520 24803
rect 2560 24771 2592 24803
rect 2632 24771 2664 24803
rect 2704 24771 2736 24803
rect 2776 24771 2808 24803
rect 2848 24771 2880 24803
rect 2920 24771 2952 24803
rect 2992 24771 3024 24803
rect 3064 24771 3096 24803
rect 3136 24771 3168 24803
rect 3208 24771 3240 24803
rect 3280 24771 3312 24803
rect 3352 24771 3384 24803
rect 3424 24771 3456 24803
rect 3496 24771 3528 24803
rect 3568 24771 3600 24803
rect 3640 24771 3672 24803
rect 3712 24771 3744 24803
rect 3784 24771 3816 24803
rect 3856 24771 3888 24803
rect 112 24699 144 24731
rect 184 24699 216 24731
rect 256 24699 288 24731
rect 328 24699 360 24731
rect 400 24699 432 24731
rect 472 24699 504 24731
rect 544 24699 576 24731
rect 616 24699 648 24731
rect 688 24699 720 24731
rect 760 24699 792 24731
rect 832 24699 864 24731
rect 904 24699 936 24731
rect 976 24699 1008 24731
rect 1048 24699 1080 24731
rect 1120 24699 1152 24731
rect 1192 24699 1224 24731
rect 1264 24699 1296 24731
rect 1336 24699 1368 24731
rect 1408 24699 1440 24731
rect 1480 24699 1512 24731
rect 1552 24699 1584 24731
rect 1624 24699 1656 24731
rect 1696 24699 1728 24731
rect 1768 24699 1800 24731
rect 1840 24699 1872 24731
rect 1912 24699 1944 24731
rect 1984 24699 2016 24731
rect 2056 24699 2088 24731
rect 2128 24699 2160 24731
rect 2200 24699 2232 24731
rect 2272 24699 2304 24731
rect 2344 24699 2376 24731
rect 2416 24699 2448 24731
rect 2488 24699 2520 24731
rect 2560 24699 2592 24731
rect 2632 24699 2664 24731
rect 2704 24699 2736 24731
rect 2776 24699 2808 24731
rect 2848 24699 2880 24731
rect 2920 24699 2952 24731
rect 2992 24699 3024 24731
rect 3064 24699 3096 24731
rect 3136 24699 3168 24731
rect 3208 24699 3240 24731
rect 3280 24699 3312 24731
rect 3352 24699 3384 24731
rect 3424 24699 3456 24731
rect 3496 24699 3528 24731
rect 3568 24699 3600 24731
rect 3640 24699 3672 24731
rect 3712 24699 3744 24731
rect 3784 24699 3816 24731
rect 3856 24699 3888 24731
rect 112 24627 144 24659
rect 184 24627 216 24659
rect 256 24627 288 24659
rect 328 24627 360 24659
rect 400 24627 432 24659
rect 472 24627 504 24659
rect 544 24627 576 24659
rect 616 24627 648 24659
rect 688 24627 720 24659
rect 760 24627 792 24659
rect 832 24627 864 24659
rect 904 24627 936 24659
rect 976 24627 1008 24659
rect 1048 24627 1080 24659
rect 1120 24627 1152 24659
rect 1192 24627 1224 24659
rect 1264 24627 1296 24659
rect 1336 24627 1368 24659
rect 1408 24627 1440 24659
rect 1480 24627 1512 24659
rect 1552 24627 1584 24659
rect 1624 24627 1656 24659
rect 1696 24627 1728 24659
rect 1768 24627 1800 24659
rect 1840 24627 1872 24659
rect 1912 24627 1944 24659
rect 1984 24627 2016 24659
rect 2056 24627 2088 24659
rect 2128 24627 2160 24659
rect 2200 24627 2232 24659
rect 2272 24627 2304 24659
rect 2344 24627 2376 24659
rect 2416 24627 2448 24659
rect 2488 24627 2520 24659
rect 2560 24627 2592 24659
rect 2632 24627 2664 24659
rect 2704 24627 2736 24659
rect 2776 24627 2808 24659
rect 2848 24627 2880 24659
rect 2920 24627 2952 24659
rect 2992 24627 3024 24659
rect 3064 24627 3096 24659
rect 3136 24627 3168 24659
rect 3208 24627 3240 24659
rect 3280 24627 3312 24659
rect 3352 24627 3384 24659
rect 3424 24627 3456 24659
rect 3496 24627 3528 24659
rect 3568 24627 3600 24659
rect 3640 24627 3672 24659
rect 3712 24627 3744 24659
rect 3784 24627 3816 24659
rect 3856 24627 3888 24659
rect 112 24555 144 24587
rect 184 24555 216 24587
rect 256 24555 288 24587
rect 328 24555 360 24587
rect 400 24555 432 24587
rect 472 24555 504 24587
rect 544 24555 576 24587
rect 616 24555 648 24587
rect 688 24555 720 24587
rect 760 24555 792 24587
rect 832 24555 864 24587
rect 904 24555 936 24587
rect 976 24555 1008 24587
rect 1048 24555 1080 24587
rect 1120 24555 1152 24587
rect 1192 24555 1224 24587
rect 1264 24555 1296 24587
rect 1336 24555 1368 24587
rect 1408 24555 1440 24587
rect 1480 24555 1512 24587
rect 1552 24555 1584 24587
rect 1624 24555 1656 24587
rect 1696 24555 1728 24587
rect 1768 24555 1800 24587
rect 1840 24555 1872 24587
rect 1912 24555 1944 24587
rect 1984 24555 2016 24587
rect 2056 24555 2088 24587
rect 2128 24555 2160 24587
rect 2200 24555 2232 24587
rect 2272 24555 2304 24587
rect 2344 24555 2376 24587
rect 2416 24555 2448 24587
rect 2488 24555 2520 24587
rect 2560 24555 2592 24587
rect 2632 24555 2664 24587
rect 2704 24555 2736 24587
rect 2776 24555 2808 24587
rect 2848 24555 2880 24587
rect 2920 24555 2952 24587
rect 2992 24555 3024 24587
rect 3064 24555 3096 24587
rect 3136 24555 3168 24587
rect 3208 24555 3240 24587
rect 3280 24555 3312 24587
rect 3352 24555 3384 24587
rect 3424 24555 3456 24587
rect 3496 24555 3528 24587
rect 3568 24555 3600 24587
rect 3640 24555 3672 24587
rect 3712 24555 3744 24587
rect 3784 24555 3816 24587
rect 3856 24555 3888 24587
rect 112 24483 144 24515
rect 184 24483 216 24515
rect 256 24483 288 24515
rect 328 24483 360 24515
rect 400 24483 432 24515
rect 472 24483 504 24515
rect 544 24483 576 24515
rect 616 24483 648 24515
rect 688 24483 720 24515
rect 760 24483 792 24515
rect 832 24483 864 24515
rect 904 24483 936 24515
rect 976 24483 1008 24515
rect 1048 24483 1080 24515
rect 1120 24483 1152 24515
rect 1192 24483 1224 24515
rect 1264 24483 1296 24515
rect 1336 24483 1368 24515
rect 1408 24483 1440 24515
rect 1480 24483 1512 24515
rect 1552 24483 1584 24515
rect 1624 24483 1656 24515
rect 1696 24483 1728 24515
rect 1768 24483 1800 24515
rect 1840 24483 1872 24515
rect 1912 24483 1944 24515
rect 1984 24483 2016 24515
rect 2056 24483 2088 24515
rect 2128 24483 2160 24515
rect 2200 24483 2232 24515
rect 2272 24483 2304 24515
rect 2344 24483 2376 24515
rect 2416 24483 2448 24515
rect 2488 24483 2520 24515
rect 2560 24483 2592 24515
rect 2632 24483 2664 24515
rect 2704 24483 2736 24515
rect 2776 24483 2808 24515
rect 2848 24483 2880 24515
rect 2920 24483 2952 24515
rect 2992 24483 3024 24515
rect 3064 24483 3096 24515
rect 3136 24483 3168 24515
rect 3208 24483 3240 24515
rect 3280 24483 3312 24515
rect 3352 24483 3384 24515
rect 3424 24483 3456 24515
rect 3496 24483 3528 24515
rect 3568 24483 3600 24515
rect 3640 24483 3672 24515
rect 3712 24483 3744 24515
rect 3784 24483 3816 24515
rect 3856 24483 3888 24515
rect 112 24411 144 24443
rect 184 24411 216 24443
rect 256 24411 288 24443
rect 328 24411 360 24443
rect 400 24411 432 24443
rect 472 24411 504 24443
rect 544 24411 576 24443
rect 616 24411 648 24443
rect 688 24411 720 24443
rect 760 24411 792 24443
rect 832 24411 864 24443
rect 904 24411 936 24443
rect 976 24411 1008 24443
rect 1048 24411 1080 24443
rect 1120 24411 1152 24443
rect 1192 24411 1224 24443
rect 1264 24411 1296 24443
rect 1336 24411 1368 24443
rect 1408 24411 1440 24443
rect 1480 24411 1512 24443
rect 1552 24411 1584 24443
rect 1624 24411 1656 24443
rect 1696 24411 1728 24443
rect 1768 24411 1800 24443
rect 1840 24411 1872 24443
rect 1912 24411 1944 24443
rect 1984 24411 2016 24443
rect 2056 24411 2088 24443
rect 2128 24411 2160 24443
rect 2200 24411 2232 24443
rect 2272 24411 2304 24443
rect 2344 24411 2376 24443
rect 2416 24411 2448 24443
rect 2488 24411 2520 24443
rect 2560 24411 2592 24443
rect 2632 24411 2664 24443
rect 2704 24411 2736 24443
rect 2776 24411 2808 24443
rect 2848 24411 2880 24443
rect 2920 24411 2952 24443
rect 2992 24411 3024 24443
rect 3064 24411 3096 24443
rect 3136 24411 3168 24443
rect 3208 24411 3240 24443
rect 3280 24411 3312 24443
rect 3352 24411 3384 24443
rect 3424 24411 3456 24443
rect 3496 24411 3528 24443
rect 3568 24411 3600 24443
rect 3640 24411 3672 24443
rect 3712 24411 3744 24443
rect 3784 24411 3816 24443
rect 3856 24411 3888 24443
rect 112 24339 144 24371
rect 184 24339 216 24371
rect 256 24339 288 24371
rect 328 24339 360 24371
rect 400 24339 432 24371
rect 472 24339 504 24371
rect 544 24339 576 24371
rect 616 24339 648 24371
rect 688 24339 720 24371
rect 760 24339 792 24371
rect 832 24339 864 24371
rect 904 24339 936 24371
rect 976 24339 1008 24371
rect 1048 24339 1080 24371
rect 1120 24339 1152 24371
rect 1192 24339 1224 24371
rect 1264 24339 1296 24371
rect 1336 24339 1368 24371
rect 1408 24339 1440 24371
rect 1480 24339 1512 24371
rect 1552 24339 1584 24371
rect 1624 24339 1656 24371
rect 1696 24339 1728 24371
rect 1768 24339 1800 24371
rect 1840 24339 1872 24371
rect 1912 24339 1944 24371
rect 1984 24339 2016 24371
rect 2056 24339 2088 24371
rect 2128 24339 2160 24371
rect 2200 24339 2232 24371
rect 2272 24339 2304 24371
rect 2344 24339 2376 24371
rect 2416 24339 2448 24371
rect 2488 24339 2520 24371
rect 2560 24339 2592 24371
rect 2632 24339 2664 24371
rect 2704 24339 2736 24371
rect 2776 24339 2808 24371
rect 2848 24339 2880 24371
rect 2920 24339 2952 24371
rect 2992 24339 3024 24371
rect 3064 24339 3096 24371
rect 3136 24339 3168 24371
rect 3208 24339 3240 24371
rect 3280 24339 3312 24371
rect 3352 24339 3384 24371
rect 3424 24339 3456 24371
rect 3496 24339 3528 24371
rect 3568 24339 3600 24371
rect 3640 24339 3672 24371
rect 3712 24339 3744 24371
rect 3784 24339 3816 24371
rect 3856 24339 3888 24371
rect 112 24267 144 24299
rect 184 24267 216 24299
rect 256 24267 288 24299
rect 328 24267 360 24299
rect 400 24267 432 24299
rect 472 24267 504 24299
rect 544 24267 576 24299
rect 616 24267 648 24299
rect 688 24267 720 24299
rect 760 24267 792 24299
rect 832 24267 864 24299
rect 904 24267 936 24299
rect 976 24267 1008 24299
rect 1048 24267 1080 24299
rect 1120 24267 1152 24299
rect 1192 24267 1224 24299
rect 1264 24267 1296 24299
rect 1336 24267 1368 24299
rect 1408 24267 1440 24299
rect 1480 24267 1512 24299
rect 1552 24267 1584 24299
rect 1624 24267 1656 24299
rect 1696 24267 1728 24299
rect 1768 24267 1800 24299
rect 1840 24267 1872 24299
rect 1912 24267 1944 24299
rect 1984 24267 2016 24299
rect 2056 24267 2088 24299
rect 2128 24267 2160 24299
rect 2200 24267 2232 24299
rect 2272 24267 2304 24299
rect 2344 24267 2376 24299
rect 2416 24267 2448 24299
rect 2488 24267 2520 24299
rect 2560 24267 2592 24299
rect 2632 24267 2664 24299
rect 2704 24267 2736 24299
rect 2776 24267 2808 24299
rect 2848 24267 2880 24299
rect 2920 24267 2952 24299
rect 2992 24267 3024 24299
rect 3064 24267 3096 24299
rect 3136 24267 3168 24299
rect 3208 24267 3240 24299
rect 3280 24267 3312 24299
rect 3352 24267 3384 24299
rect 3424 24267 3456 24299
rect 3496 24267 3528 24299
rect 3568 24267 3600 24299
rect 3640 24267 3672 24299
rect 3712 24267 3744 24299
rect 3784 24267 3816 24299
rect 3856 24267 3888 24299
rect 112 24195 144 24227
rect 184 24195 216 24227
rect 256 24195 288 24227
rect 328 24195 360 24227
rect 400 24195 432 24227
rect 472 24195 504 24227
rect 544 24195 576 24227
rect 616 24195 648 24227
rect 688 24195 720 24227
rect 760 24195 792 24227
rect 832 24195 864 24227
rect 904 24195 936 24227
rect 976 24195 1008 24227
rect 1048 24195 1080 24227
rect 1120 24195 1152 24227
rect 1192 24195 1224 24227
rect 1264 24195 1296 24227
rect 1336 24195 1368 24227
rect 1408 24195 1440 24227
rect 1480 24195 1512 24227
rect 1552 24195 1584 24227
rect 1624 24195 1656 24227
rect 1696 24195 1728 24227
rect 1768 24195 1800 24227
rect 1840 24195 1872 24227
rect 1912 24195 1944 24227
rect 1984 24195 2016 24227
rect 2056 24195 2088 24227
rect 2128 24195 2160 24227
rect 2200 24195 2232 24227
rect 2272 24195 2304 24227
rect 2344 24195 2376 24227
rect 2416 24195 2448 24227
rect 2488 24195 2520 24227
rect 2560 24195 2592 24227
rect 2632 24195 2664 24227
rect 2704 24195 2736 24227
rect 2776 24195 2808 24227
rect 2848 24195 2880 24227
rect 2920 24195 2952 24227
rect 2992 24195 3024 24227
rect 3064 24195 3096 24227
rect 3136 24195 3168 24227
rect 3208 24195 3240 24227
rect 3280 24195 3312 24227
rect 3352 24195 3384 24227
rect 3424 24195 3456 24227
rect 3496 24195 3528 24227
rect 3568 24195 3600 24227
rect 3640 24195 3672 24227
rect 3712 24195 3744 24227
rect 3784 24195 3816 24227
rect 3856 24195 3888 24227
rect 112 24123 144 24155
rect 184 24123 216 24155
rect 256 24123 288 24155
rect 328 24123 360 24155
rect 400 24123 432 24155
rect 472 24123 504 24155
rect 544 24123 576 24155
rect 616 24123 648 24155
rect 688 24123 720 24155
rect 760 24123 792 24155
rect 832 24123 864 24155
rect 904 24123 936 24155
rect 976 24123 1008 24155
rect 1048 24123 1080 24155
rect 1120 24123 1152 24155
rect 1192 24123 1224 24155
rect 1264 24123 1296 24155
rect 1336 24123 1368 24155
rect 1408 24123 1440 24155
rect 1480 24123 1512 24155
rect 1552 24123 1584 24155
rect 1624 24123 1656 24155
rect 1696 24123 1728 24155
rect 1768 24123 1800 24155
rect 1840 24123 1872 24155
rect 1912 24123 1944 24155
rect 1984 24123 2016 24155
rect 2056 24123 2088 24155
rect 2128 24123 2160 24155
rect 2200 24123 2232 24155
rect 2272 24123 2304 24155
rect 2344 24123 2376 24155
rect 2416 24123 2448 24155
rect 2488 24123 2520 24155
rect 2560 24123 2592 24155
rect 2632 24123 2664 24155
rect 2704 24123 2736 24155
rect 2776 24123 2808 24155
rect 2848 24123 2880 24155
rect 2920 24123 2952 24155
rect 2992 24123 3024 24155
rect 3064 24123 3096 24155
rect 3136 24123 3168 24155
rect 3208 24123 3240 24155
rect 3280 24123 3312 24155
rect 3352 24123 3384 24155
rect 3424 24123 3456 24155
rect 3496 24123 3528 24155
rect 3568 24123 3600 24155
rect 3640 24123 3672 24155
rect 3712 24123 3744 24155
rect 3784 24123 3816 24155
rect 3856 24123 3888 24155
rect 112 24051 144 24083
rect 184 24051 216 24083
rect 256 24051 288 24083
rect 328 24051 360 24083
rect 400 24051 432 24083
rect 472 24051 504 24083
rect 544 24051 576 24083
rect 616 24051 648 24083
rect 688 24051 720 24083
rect 760 24051 792 24083
rect 832 24051 864 24083
rect 904 24051 936 24083
rect 976 24051 1008 24083
rect 1048 24051 1080 24083
rect 1120 24051 1152 24083
rect 1192 24051 1224 24083
rect 1264 24051 1296 24083
rect 1336 24051 1368 24083
rect 1408 24051 1440 24083
rect 1480 24051 1512 24083
rect 1552 24051 1584 24083
rect 1624 24051 1656 24083
rect 1696 24051 1728 24083
rect 1768 24051 1800 24083
rect 1840 24051 1872 24083
rect 1912 24051 1944 24083
rect 1984 24051 2016 24083
rect 2056 24051 2088 24083
rect 2128 24051 2160 24083
rect 2200 24051 2232 24083
rect 2272 24051 2304 24083
rect 2344 24051 2376 24083
rect 2416 24051 2448 24083
rect 2488 24051 2520 24083
rect 2560 24051 2592 24083
rect 2632 24051 2664 24083
rect 2704 24051 2736 24083
rect 2776 24051 2808 24083
rect 2848 24051 2880 24083
rect 2920 24051 2952 24083
rect 2992 24051 3024 24083
rect 3064 24051 3096 24083
rect 3136 24051 3168 24083
rect 3208 24051 3240 24083
rect 3280 24051 3312 24083
rect 3352 24051 3384 24083
rect 3424 24051 3456 24083
rect 3496 24051 3528 24083
rect 3568 24051 3600 24083
rect 3640 24051 3672 24083
rect 3712 24051 3744 24083
rect 3784 24051 3816 24083
rect 3856 24051 3888 24083
rect 112 23979 144 24011
rect 184 23979 216 24011
rect 256 23979 288 24011
rect 328 23979 360 24011
rect 400 23979 432 24011
rect 472 23979 504 24011
rect 544 23979 576 24011
rect 616 23979 648 24011
rect 688 23979 720 24011
rect 760 23979 792 24011
rect 832 23979 864 24011
rect 904 23979 936 24011
rect 976 23979 1008 24011
rect 1048 23979 1080 24011
rect 1120 23979 1152 24011
rect 1192 23979 1224 24011
rect 1264 23979 1296 24011
rect 1336 23979 1368 24011
rect 1408 23979 1440 24011
rect 1480 23979 1512 24011
rect 1552 23979 1584 24011
rect 1624 23979 1656 24011
rect 1696 23979 1728 24011
rect 1768 23979 1800 24011
rect 1840 23979 1872 24011
rect 1912 23979 1944 24011
rect 1984 23979 2016 24011
rect 2056 23979 2088 24011
rect 2128 23979 2160 24011
rect 2200 23979 2232 24011
rect 2272 23979 2304 24011
rect 2344 23979 2376 24011
rect 2416 23979 2448 24011
rect 2488 23979 2520 24011
rect 2560 23979 2592 24011
rect 2632 23979 2664 24011
rect 2704 23979 2736 24011
rect 2776 23979 2808 24011
rect 2848 23979 2880 24011
rect 2920 23979 2952 24011
rect 2992 23979 3024 24011
rect 3064 23979 3096 24011
rect 3136 23979 3168 24011
rect 3208 23979 3240 24011
rect 3280 23979 3312 24011
rect 3352 23979 3384 24011
rect 3424 23979 3456 24011
rect 3496 23979 3528 24011
rect 3568 23979 3600 24011
rect 3640 23979 3672 24011
rect 3712 23979 3744 24011
rect 3784 23979 3816 24011
rect 3856 23979 3888 24011
rect 112 23907 144 23939
rect 184 23907 216 23939
rect 256 23907 288 23939
rect 328 23907 360 23939
rect 400 23907 432 23939
rect 472 23907 504 23939
rect 544 23907 576 23939
rect 616 23907 648 23939
rect 688 23907 720 23939
rect 760 23907 792 23939
rect 832 23907 864 23939
rect 904 23907 936 23939
rect 976 23907 1008 23939
rect 1048 23907 1080 23939
rect 1120 23907 1152 23939
rect 1192 23907 1224 23939
rect 1264 23907 1296 23939
rect 1336 23907 1368 23939
rect 1408 23907 1440 23939
rect 1480 23907 1512 23939
rect 1552 23907 1584 23939
rect 1624 23907 1656 23939
rect 1696 23907 1728 23939
rect 1768 23907 1800 23939
rect 1840 23907 1872 23939
rect 1912 23907 1944 23939
rect 1984 23907 2016 23939
rect 2056 23907 2088 23939
rect 2128 23907 2160 23939
rect 2200 23907 2232 23939
rect 2272 23907 2304 23939
rect 2344 23907 2376 23939
rect 2416 23907 2448 23939
rect 2488 23907 2520 23939
rect 2560 23907 2592 23939
rect 2632 23907 2664 23939
rect 2704 23907 2736 23939
rect 2776 23907 2808 23939
rect 2848 23907 2880 23939
rect 2920 23907 2952 23939
rect 2992 23907 3024 23939
rect 3064 23907 3096 23939
rect 3136 23907 3168 23939
rect 3208 23907 3240 23939
rect 3280 23907 3312 23939
rect 3352 23907 3384 23939
rect 3424 23907 3456 23939
rect 3496 23907 3528 23939
rect 3568 23907 3600 23939
rect 3640 23907 3672 23939
rect 3712 23907 3744 23939
rect 3784 23907 3816 23939
rect 3856 23907 3888 23939
rect 112 23835 144 23867
rect 184 23835 216 23867
rect 256 23835 288 23867
rect 328 23835 360 23867
rect 400 23835 432 23867
rect 472 23835 504 23867
rect 544 23835 576 23867
rect 616 23835 648 23867
rect 688 23835 720 23867
rect 760 23835 792 23867
rect 832 23835 864 23867
rect 904 23835 936 23867
rect 976 23835 1008 23867
rect 1048 23835 1080 23867
rect 1120 23835 1152 23867
rect 1192 23835 1224 23867
rect 1264 23835 1296 23867
rect 1336 23835 1368 23867
rect 1408 23835 1440 23867
rect 1480 23835 1512 23867
rect 1552 23835 1584 23867
rect 1624 23835 1656 23867
rect 1696 23835 1728 23867
rect 1768 23835 1800 23867
rect 1840 23835 1872 23867
rect 1912 23835 1944 23867
rect 1984 23835 2016 23867
rect 2056 23835 2088 23867
rect 2128 23835 2160 23867
rect 2200 23835 2232 23867
rect 2272 23835 2304 23867
rect 2344 23835 2376 23867
rect 2416 23835 2448 23867
rect 2488 23835 2520 23867
rect 2560 23835 2592 23867
rect 2632 23835 2664 23867
rect 2704 23835 2736 23867
rect 2776 23835 2808 23867
rect 2848 23835 2880 23867
rect 2920 23835 2952 23867
rect 2992 23835 3024 23867
rect 3064 23835 3096 23867
rect 3136 23835 3168 23867
rect 3208 23835 3240 23867
rect 3280 23835 3312 23867
rect 3352 23835 3384 23867
rect 3424 23835 3456 23867
rect 3496 23835 3528 23867
rect 3568 23835 3600 23867
rect 3640 23835 3672 23867
rect 3712 23835 3744 23867
rect 3784 23835 3816 23867
rect 3856 23835 3888 23867
rect 112 23763 144 23795
rect 184 23763 216 23795
rect 256 23763 288 23795
rect 328 23763 360 23795
rect 400 23763 432 23795
rect 472 23763 504 23795
rect 544 23763 576 23795
rect 616 23763 648 23795
rect 688 23763 720 23795
rect 760 23763 792 23795
rect 832 23763 864 23795
rect 904 23763 936 23795
rect 976 23763 1008 23795
rect 1048 23763 1080 23795
rect 1120 23763 1152 23795
rect 1192 23763 1224 23795
rect 1264 23763 1296 23795
rect 1336 23763 1368 23795
rect 1408 23763 1440 23795
rect 1480 23763 1512 23795
rect 1552 23763 1584 23795
rect 1624 23763 1656 23795
rect 1696 23763 1728 23795
rect 1768 23763 1800 23795
rect 1840 23763 1872 23795
rect 1912 23763 1944 23795
rect 1984 23763 2016 23795
rect 2056 23763 2088 23795
rect 2128 23763 2160 23795
rect 2200 23763 2232 23795
rect 2272 23763 2304 23795
rect 2344 23763 2376 23795
rect 2416 23763 2448 23795
rect 2488 23763 2520 23795
rect 2560 23763 2592 23795
rect 2632 23763 2664 23795
rect 2704 23763 2736 23795
rect 2776 23763 2808 23795
rect 2848 23763 2880 23795
rect 2920 23763 2952 23795
rect 2992 23763 3024 23795
rect 3064 23763 3096 23795
rect 3136 23763 3168 23795
rect 3208 23763 3240 23795
rect 3280 23763 3312 23795
rect 3352 23763 3384 23795
rect 3424 23763 3456 23795
rect 3496 23763 3528 23795
rect 3568 23763 3600 23795
rect 3640 23763 3672 23795
rect 3712 23763 3744 23795
rect 3784 23763 3816 23795
rect 3856 23763 3888 23795
rect 112 23691 144 23723
rect 184 23691 216 23723
rect 256 23691 288 23723
rect 328 23691 360 23723
rect 400 23691 432 23723
rect 472 23691 504 23723
rect 544 23691 576 23723
rect 616 23691 648 23723
rect 688 23691 720 23723
rect 760 23691 792 23723
rect 832 23691 864 23723
rect 904 23691 936 23723
rect 976 23691 1008 23723
rect 1048 23691 1080 23723
rect 1120 23691 1152 23723
rect 1192 23691 1224 23723
rect 1264 23691 1296 23723
rect 1336 23691 1368 23723
rect 1408 23691 1440 23723
rect 1480 23691 1512 23723
rect 1552 23691 1584 23723
rect 1624 23691 1656 23723
rect 1696 23691 1728 23723
rect 1768 23691 1800 23723
rect 1840 23691 1872 23723
rect 1912 23691 1944 23723
rect 1984 23691 2016 23723
rect 2056 23691 2088 23723
rect 2128 23691 2160 23723
rect 2200 23691 2232 23723
rect 2272 23691 2304 23723
rect 2344 23691 2376 23723
rect 2416 23691 2448 23723
rect 2488 23691 2520 23723
rect 2560 23691 2592 23723
rect 2632 23691 2664 23723
rect 2704 23691 2736 23723
rect 2776 23691 2808 23723
rect 2848 23691 2880 23723
rect 2920 23691 2952 23723
rect 2992 23691 3024 23723
rect 3064 23691 3096 23723
rect 3136 23691 3168 23723
rect 3208 23691 3240 23723
rect 3280 23691 3312 23723
rect 3352 23691 3384 23723
rect 3424 23691 3456 23723
rect 3496 23691 3528 23723
rect 3568 23691 3600 23723
rect 3640 23691 3672 23723
rect 3712 23691 3744 23723
rect 3784 23691 3816 23723
rect 3856 23691 3888 23723
rect 112 23619 144 23651
rect 184 23619 216 23651
rect 256 23619 288 23651
rect 328 23619 360 23651
rect 400 23619 432 23651
rect 472 23619 504 23651
rect 544 23619 576 23651
rect 616 23619 648 23651
rect 688 23619 720 23651
rect 760 23619 792 23651
rect 832 23619 864 23651
rect 904 23619 936 23651
rect 976 23619 1008 23651
rect 1048 23619 1080 23651
rect 1120 23619 1152 23651
rect 1192 23619 1224 23651
rect 1264 23619 1296 23651
rect 1336 23619 1368 23651
rect 1408 23619 1440 23651
rect 1480 23619 1512 23651
rect 1552 23619 1584 23651
rect 1624 23619 1656 23651
rect 1696 23619 1728 23651
rect 1768 23619 1800 23651
rect 1840 23619 1872 23651
rect 1912 23619 1944 23651
rect 1984 23619 2016 23651
rect 2056 23619 2088 23651
rect 2128 23619 2160 23651
rect 2200 23619 2232 23651
rect 2272 23619 2304 23651
rect 2344 23619 2376 23651
rect 2416 23619 2448 23651
rect 2488 23619 2520 23651
rect 2560 23619 2592 23651
rect 2632 23619 2664 23651
rect 2704 23619 2736 23651
rect 2776 23619 2808 23651
rect 2848 23619 2880 23651
rect 2920 23619 2952 23651
rect 2992 23619 3024 23651
rect 3064 23619 3096 23651
rect 3136 23619 3168 23651
rect 3208 23619 3240 23651
rect 3280 23619 3312 23651
rect 3352 23619 3384 23651
rect 3424 23619 3456 23651
rect 3496 23619 3528 23651
rect 3568 23619 3600 23651
rect 3640 23619 3672 23651
rect 3712 23619 3744 23651
rect 3784 23619 3816 23651
rect 3856 23619 3888 23651
rect 112 23547 144 23579
rect 184 23547 216 23579
rect 256 23547 288 23579
rect 328 23547 360 23579
rect 400 23547 432 23579
rect 472 23547 504 23579
rect 544 23547 576 23579
rect 616 23547 648 23579
rect 688 23547 720 23579
rect 760 23547 792 23579
rect 832 23547 864 23579
rect 904 23547 936 23579
rect 976 23547 1008 23579
rect 1048 23547 1080 23579
rect 1120 23547 1152 23579
rect 1192 23547 1224 23579
rect 1264 23547 1296 23579
rect 1336 23547 1368 23579
rect 1408 23547 1440 23579
rect 1480 23547 1512 23579
rect 1552 23547 1584 23579
rect 1624 23547 1656 23579
rect 1696 23547 1728 23579
rect 1768 23547 1800 23579
rect 1840 23547 1872 23579
rect 1912 23547 1944 23579
rect 1984 23547 2016 23579
rect 2056 23547 2088 23579
rect 2128 23547 2160 23579
rect 2200 23547 2232 23579
rect 2272 23547 2304 23579
rect 2344 23547 2376 23579
rect 2416 23547 2448 23579
rect 2488 23547 2520 23579
rect 2560 23547 2592 23579
rect 2632 23547 2664 23579
rect 2704 23547 2736 23579
rect 2776 23547 2808 23579
rect 2848 23547 2880 23579
rect 2920 23547 2952 23579
rect 2992 23547 3024 23579
rect 3064 23547 3096 23579
rect 3136 23547 3168 23579
rect 3208 23547 3240 23579
rect 3280 23547 3312 23579
rect 3352 23547 3384 23579
rect 3424 23547 3456 23579
rect 3496 23547 3528 23579
rect 3568 23547 3600 23579
rect 3640 23547 3672 23579
rect 3712 23547 3744 23579
rect 3784 23547 3816 23579
rect 3856 23547 3888 23579
rect 112 23475 144 23507
rect 184 23475 216 23507
rect 256 23475 288 23507
rect 328 23475 360 23507
rect 400 23475 432 23507
rect 472 23475 504 23507
rect 544 23475 576 23507
rect 616 23475 648 23507
rect 688 23475 720 23507
rect 760 23475 792 23507
rect 832 23475 864 23507
rect 904 23475 936 23507
rect 976 23475 1008 23507
rect 1048 23475 1080 23507
rect 1120 23475 1152 23507
rect 1192 23475 1224 23507
rect 1264 23475 1296 23507
rect 1336 23475 1368 23507
rect 1408 23475 1440 23507
rect 1480 23475 1512 23507
rect 1552 23475 1584 23507
rect 1624 23475 1656 23507
rect 1696 23475 1728 23507
rect 1768 23475 1800 23507
rect 1840 23475 1872 23507
rect 1912 23475 1944 23507
rect 1984 23475 2016 23507
rect 2056 23475 2088 23507
rect 2128 23475 2160 23507
rect 2200 23475 2232 23507
rect 2272 23475 2304 23507
rect 2344 23475 2376 23507
rect 2416 23475 2448 23507
rect 2488 23475 2520 23507
rect 2560 23475 2592 23507
rect 2632 23475 2664 23507
rect 2704 23475 2736 23507
rect 2776 23475 2808 23507
rect 2848 23475 2880 23507
rect 2920 23475 2952 23507
rect 2992 23475 3024 23507
rect 3064 23475 3096 23507
rect 3136 23475 3168 23507
rect 3208 23475 3240 23507
rect 3280 23475 3312 23507
rect 3352 23475 3384 23507
rect 3424 23475 3456 23507
rect 3496 23475 3528 23507
rect 3568 23475 3600 23507
rect 3640 23475 3672 23507
rect 3712 23475 3744 23507
rect 3784 23475 3816 23507
rect 3856 23475 3888 23507
rect 112 23403 144 23435
rect 184 23403 216 23435
rect 256 23403 288 23435
rect 328 23403 360 23435
rect 400 23403 432 23435
rect 472 23403 504 23435
rect 544 23403 576 23435
rect 616 23403 648 23435
rect 688 23403 720 23435
rect 760 23403 792 23435
rect 832 23403 864 23435
rect 904 23403 936 23435
rect 976 23403 1008 23435
rect 1048 23403 1080 23435
rect 1120 23403 1152 23435
rect 1192 23403 1224 23435
rect 1264 23403 1296 23435
rect 1336 23403 1368 23435
rect 1408 23403 1440 23435
rect 1480 23403 1512 23435
rect 1552 23403 1584 23435
rect 1624 23403 1656 23435
rect 1696 23403 1728 23435
rect 1768 23403 1800 23435
rect 1840 23403 1872 23435
rect 1912 23403 1944 23435
rect 1984 23403 2016 23435
rect 2056 23403 2088 23435
rect 2128 23403 2160 23435
rect 2200 23403 2232 23435
rect 2272 23403 2304 23435
rect 2344 23403 2376 23435
rect 2416 23403 2448 23435
rect 2488 23403 2520 23435
rect 2560 23403 2592 23435
rect 2632 23403 2664 23435
rect 2704 23403 2736 23435
rect 2776 23403 2808 23435
rect 2848 23403 2880 23435
rect 2920 23403 2952 23435
rect 2992 23403 3024 23435
rect 3064 23403 3096 23435
rect 3136 23403 3168 23435
rect 3208 23403 3240 23435
rect 3280 23403 3312 23435
rect 3352 23403 3384 23435
rect 3424 23403 3456 23435
rect 3496 23403 3528 23435
rect 3568 23403 3600 23435
rect 3640 23403 3672 23435
rect 3712 23403 3744 23435
rect 3784 23403 3816 23435
rect 3856 23403 3888 23435
rect 112 23331 144 23363
rect 184 23331 216 23363
rect 256 23331 288 23363
rect 328 23331 360 23363
rect 400 23331 432 23363
rect 472 23331 504 23363
rect 544 23331 576 23363
rect 616 23331 648 23363
rect 688 23331 720 23363
rect 760 23331 792 23363
rect 832 23331 864 23363
rect 904 23331 936 23363
rect 976 23331 1008 23363
rect 1048 23331 1080 23363
rect 1120 23331 1152 23363
rect 1192 23331 1224 23363
rect 1264 23331 1296 23363
rect 1336 23331 1368 23363
rect 1408 23331 1440 23363
rect 1480 23331 1512 23363
rect 1552 23331 1584 23363
rect 1624 23331 1656 23363
rect 1696 23331 1728 23363
rect 1768 23331 1800 23363
rect 1840 23331 1872 23363
rect 1912 23331 1944 23363
rect 1984 23331 2016 23363
rect 2056 23331 2088 23363
rect 2128 23331 2160 23363
rect 2200 23331 2232 23363
rect 2272 23331 2304 23363
rect 2344 23331 2376 23363
rect 2416 23331 2448 23363
rect 2488 23331 2520 23363
rect 2560 23331 2592 23363
rect 2632 23331 2664 23363
rect 2704 23331 2736 23363
rect 2776 23331 2808 23363
rect 2848 23331 2880 23363
rect 2920 23331 2952 23363
rect 2992 23331 3024 23363
rect 3064 23331 3096 23363
rect 3136 23331 3168 23363
rect 3208 23331 3240 23363
rect 3280 23331 3312 23363
rect 3352 23331 3384 23363
rect 3424 23331 3456 23363
rect 3496 23331 3528 23363
rect 3568 23331 3600 23363
rect 3640 23331 3672 23363
rect 3712 23331 3744 23363
rect 3784 23331 3816 23363
rect 3856 23331 3888 23363
rect 112 23259 144 23291
rect 184 23259 216 23291
rect 256 23259 288 23291
rect 328 23259 360 23291
rect 400 23259 432 23291
rect 472 23259 504 23291
rect 544 23259 576 23291
rect 616 23259 648 23291
rect 688 23259 720 23291
rect 760 23259 792 23291
rect 832 23259 864 23291
rect 904 23259 936 23291
rect 976 23259 1008 23291
rect 1048 23259 1080 23291
rect 1120 23259 1152 23291
rect 1192 23259 1224 23291
rect 1264 23259 1296 23291
rect 1336 23259 1368 23291
rect 1408 23259 1440 23291
rect 1480 23259 1512 23291
rect 1552 23259 1584 23291
rect 1624 23259 1656 23291
rect 1696 23259 1728 23291
rect 1768 23259 1800 23291
rect 1840 23259 1872 23291
rect 1912 23259 1944 23291
rect 1984 23259 2016 23291
rect 2056 23259 2088 23291
rect 2128 23259 2160 23291
rect 2200 23259 2232 23291
rect 2272 23259 2304 23291
rect 2344 23259 2376 23291
rect 2416 23259 2448 23291
rect 2488 23259 2520 23291
rect 2560 23259 2592 23291
rect 2632 23259 2664 23291
rect 2704 23259 2736 23291
rect 2776 23259 2808 23291
rect 2848 23259 2880 23291
rect 2920 23259 2952 23291
rect 2992 23259 3024 23291
rect 3064 23259 3096 23291
rect 3136 23259 3168 23291
rect 3208 23259 3240 23291
rect 3280 23259 3312 23291
rect 3352 23259 3384 23291
rect 3424 23259 3456 23291
rect 3496 23259 3528 23291
rect 3568 23259 3600 23291
rect 3640 23259 3672 23291
rect 3712 23259 3744 23291
rect 3784 23259 3816 23291
rect 3856 23259 3888 23291
rect 112 23187 144 23219
rect 184 23187 216 23219
rect 256 23187 288 23219
rect 328 23187 360 23219
rect 400 23187 432 23219
rect 472 23187 504 23219
rect 544 23187 576 23219
rect 616 23187 648 23219
rect 688 23187 720 23219
rect 760 23187 792 23219
rect 832 23187 864 23219
rect 904 23187 936 23219
rect 976 23187 1008 23219
rect 1048 23187 1080 23219
rect 1120 23187 1152 23219
rect 1192 23187 1224 23219
rect 1264 23187 1296 23219
rect 1336 23187 1368 23219
rect 1408 23187 1440 23219
rect 1480 23187 1512 23219
rect 1552 23187 1584 23219
rect 1624 23187 1656 23219
rect 1696 23187 1728 23219
rect 1768 23187 1800 23219
rect 1840 23187 1872 23219
rect 1912 23187 1944 23219
rect 1984 23187 2016 23219
rect 2056 23187 2088 23219
rect 2128 23187 2160 23219
rect 2200 23187 2232 23219
rect 2272 23187 2304 23219
rect 2344 23187 2376 23219
rect 2416 23187 2448 23219
rect 2488 23187 2520 23219
rect 2560 23187 2592 23219
rect 2632 23187 2664 23219
rect 2704 23187 2736 23219
rect 2776 23187 2808 23219
rect 2848 23187 2880 23219
rect 2920 23187 2952 23219
rect 2992 23187 3024 23219
rect 3064 23187 3096 23219
rect 3136 23187 3168 23219
rect 3208 23187 3240 23219
rect 3280 23187 3312 23219
rect 3352 23187 3384 23219
rect 3424 23187 3456 23219
rect 3496 23187 3528 23219
rect 3568 23187 3600 23219
rect 3640 23187 3672 23219
rect 3712 23187 3744 23219
rect 3784 23187 3816 23219
rect 3856 23187 3888 23219
rect 184 22842 216 22874
rect 256 22842 288 22874
rect 328 22842 360 22874
rect 400 22842 432 22874
rect 472 22842 504 22874
rect 544 22842 576 22874
rect 616 22842 648 22874
rect 688 22842 720 22874
rect 760 22842 792 22874
rect 832 22842 864 22874
rect 904 22842 936 22874
rect 976 22842 1008 22874
rect 1048 22842 1080 22874
rect 1120 22842 1152 22874
rect 1192 22842 1224 22874
rect 1264 22842 1296 22874
rect 1336 22842 1368 22874
rect 1408 22842 1440 22874
rect 1480 22842 1512 22874
rect 1552 22842 1584 22874
rect 1624 22842 1656 22874
rect 1696 22842 1728 22874
rect 1768 22842 1800 22874
rect 1840 22842 1872 22874
rect 1912 22842 1944 22874
rect 1984 22842 2016 22874
rect 2056 22842 2088 22874
rect 2128 22842 2160 22874
rect 2200 22842 2232 22874
rect 2272 22842 2304 22874
rect 2344 22842 2376 22874
rect 2416 22842 2448 22874
rect 2488 22842 2520 22874
rect 2560 22842 2592 22874
rect 2632 22842 2664 22874
rect 2704 22842 2736 22874
rect 2776 22842 2808 22874
rect 2848 22842 2880 22874
rect 2920 22842 2952 22874
rect 2992 22842 3024 22874
rect 3064 22842 3096 22874
rect 3136 22842 3168 22874
rect 3208 22842 3240 22874
rect 3280 22842 3312 22874
rect 3352 22842 3384 22874
rect 3424 22842 3456 22874
rect 3496 22842 3528 22874
rect 3568 22842 3600 22874
rect 3640 22842 3672 22874
rect 3712 22842 3744 22874
rect 3784 22842 3816 22874
rect 3856 22842 3888 22874
rect 112 22770 144 22802
rect 184 22770 216 22802
rect 256 22770 288 22802
rect 328 22770 360 22802
rect 400 22770 432 22802
rect 472 22770 504 22802
rect 544 22770 576 22802
rect 616 22770 648 22802
rect 688 22770 720 22802
rect 760 22770 792 22802
rect 832 22770 864 22802
rect 904 22770 936 22802
rect 976 22770 1008 22802
rect 1048 22770 1080 22802
rect 1120 22770 1152 22802
rect 1192 22770 1224 22802
rect 1264 22770 1296 22802
rect 1336 22770 1368 22802
rect 1408 22770 1440 22802
rect 1480 22770 1512 22802
rect 1552 22770 1584 22802
rect 1624 22770 1656 22802
rect 1696 22770 1728 22802
rect 1768 22770 1800 22802
rect 1840 22770 1872 22802
rect 1912 22770 1944 22802
rect 1984 22770 2016 22802
rect 2056 22770 2088 22802
rect 2128 22770 2160 22802
rect 2200 22770 2232 22802
rect 2272 22770 2304 22802
rect 2344 22770 2376 22802
rect 2416 22770 2448 22802
rect 2488 22770 2520 22802
rect 2560 22770 2592 22802
rect 2632 22770 2664 22802
rect 2704 22770 2736 22802
rect 2776 22770 2808 22802
rect 2848 22770 2880 22802
rect 2920 22770 2952 22802
rect 2992 22770 3024 22802
rect 3064 22770 3096 22802
rect 3136 22770 3168 22802
rect 3208 22770 3240 22802
rect 3280 22770 3312 22802
rect 3352 22770 3384 22802
rect 3424 22770 3456 22802
rect 3496 22770 3528 22802
rect 3568 22770 3600 22802
rect 3640 22770 3672 22802
rect 3712 22770 3744 22802
rect 3784 22770 3816 22802
rect 3856 22770 3888 22802
rect 112 22698 144 22730
rect 184 22698 216 22730
rect 256 22698 288 22730
rect 328 22698 360 22730
rect 400 22698 432 22730
rect 472 22698 504 22730
rect 544 22698 576 22730
rect 616 22698 648 22730
rect 688 22698 720 22730
rect 760 22698 792 22730
rect 832 22698 864 22730
rect 904 22698 936 22730
rect 976 22698 1008 22730
rect 1048 22698 1080 22730
rect 1120 22698 1152 22730
rect 1192 22698 1224 22730
rect 1264 22698 1296 22730
rect 1336 22698 1368 22730
rect 1408 22698 1440 22730
rect 1480 22698 1512 22730
rect 1552 22698 1584 22730
rect 1624 22698 1656 22730
rect 1696 22698 1728 22730
rect 1768 22698 1800 22730
rect 1840 22698 1872 22730
rect 1912 22698 1944 22730
rect 1984 22698 2016 22730
rect 2056 22698 2088 22730
rect 2128 22698 2160 22730
rect 2200 22698 2232 22730
rect 2272 22698 2304 22730
rect 2344 22698 2376 22730
rect 2416 22698 2448 22730
rect 2488 22698 2520 22730
rect 2560 22698 2592 22730
rect 2632 22698 2664 22730
rect 2704 22698 2736 22730
rect 2776 22698 2808 22730
rect 2848 22698 2880 22730
rect 2920 22698 2952 22730
rect 2992 22698 3024 22730
rect 3064 22698 3096 22730
rect 3136 22698 3168 22730
rect 3208 22698 3240 22730
rect 3280 22698 3312 22730
rect 3352 22698 3384 22730
rect 3424 22698 3456 22730
rect 3496 22698 3528 22730
rect 3568 22698 3600 22730
rect 3640 22698 3672 22730
rect 3712 22698 3744 22730
rect 3784 22698 3816 22730
rect 3856 22698 3888 22730
rect 112 22626 144 22658
rect 184 22626 216 22658
rect 256 22626 288 22658
rect 328 22626 360 22658
rect 400 22626 432 22658
rect 472 22626 504 22658
rect 544 22626 576 22658
rect 616 22626 648 22658
rect 688 22626 720 22658
rect 760 22626 792 22658
rect 832 22626 864 22658
rect 904 22626 936 22658
rect 976 22626 1008 22658
rect 1048 22626 1080 22658
rect 1120 22626 1152 22658
rect 1192 22626 1224 22658
rect 1264 22626 1296 22658
rect 1336 22626 1368 22658
rect 1408 22626 1440 22658
rect 1480 22626 1512 22658
rect 1552 22626 1584 22658
rect 1624 22626 1656 22658
rect 1696 22626 1728 22658
rect 1768 22626 1800 22658
rect 1840 22626 1872 22658
rect 1912 22626 1944 22658
rect 1984 22626 2016 22658
rect 2056 22626 2088 22658
rect 2128 22626 2160 22658
rect 2200 22626 2232 22658
rect 2272 22626 2304 22658
rect 2344 22626 2376 22658
rect 2416 22626 2448 22658
rect 2488 22626 2520 22658
rect 2560 22626 2592 22658
rect 2632 22626 2664 22658
rect 2704 22626 2736 22658
rect 2776 22626 2808 22658
rect 2848 22626 2880 22658
rect 2920 22626 2952 22658
rect 2992 22626 3024 22658
rect 3064 22626 3096 22658
rect 3136 22626 3168 22658
rect 3208 22626 3240 22658
rect 3280 22626 3312 22658
rect 3352 22626 3384 22658
rect 3424 22626 3456 22658
rect 3496 22626 3528 22658
rect 3568 22626 3600 22658
rect 3640 22626 3672 22658
rect 3712 22626 3744 22658
rect 3784 22626 3816 22658
rect 3856 22626 3888 22658
rect 112 22554 144 22586
rect 184 22554 216 22586
rect 256 22554 288 22586
rect 328 22554 360 22586
rect 400 22554 432 22586
rect 472 22554 504 22586
rect 544 22554 576 22586
rect 616 22554 648 22586
rect 688 22554 720 22586
rect 760 22554 792 22586
rect 832 22554 864 22586
rect 904 22554 936 22586
rect 976 22554 1008 22586
rect 1048 22554 1080 22586
rect 1120 22554 1152 22586
rect 1192 22554 1224 22586
rect 1264 22554 1296 22586
rect 1336 22554 1368 22586
rect 1408 22554 1440 22586
rect 1480 22554 1512 22586
rect 1552 22554 1584 22586
rect 1624 22554 1656 22586
rect 1696 22554 1728 22586
rect 1768 22554 1800 22586
rect 1840 22554 1872 22586
rect 1912 22554 1944 22586
rect 1984 22554 2016 22586
rect 2056 22554 2088 22586
rect 2128 22554 2160 22586
rect 2200 22554 2232 22586
rect 2272 22554 2304 22586
rect 2344 22554 2376 22586
rect 2416 22554 2448 22586
rect 2488 22554 2520 22586
rect 2560 22554 2592 22586
rect 2632 22554 2664 22586
rect 2704 22554 2736 22586
rect 2776 22554 2808 22586
rect 2848 22554 2880 22586
rect 2920 22554 2952 22586
rect 2992 22554 3024 22586
rect 3064 22554 3096 22586
rect 3136 22554 3168 22586
rect 3208 22554 3240 22586
rect 3280 22554 3312 22586
rect 3352 22554 3384 22586
rect 3424 22554 3456 22586
rect 3496 22554 3528 22586
rect 3568 22554 3600 22586
rect 3640 22554 3672 22586
rect 3712 22554 3744 22586
rect 3784 22554 3816 22586
rect 3856 22554 3888 22586
rect 112 22482 144 22514
rect 184 22482 216 22514
rect 256 22482 288 22514
rect 328 22482 360 22514
rect 400 22482 432 22514
rect 472 22482 504 22514
rect 544 22482 576 22514
rect 616 22482 648 22514
rect 688 22482 720 22514
rect 760 22482 792 22514
rect 832 22482 864 22514
rect 904 22482 936 22514
rect 976 22482 1008 22514
rect 1048 22482 1080 22514
rect 1120 22482 1152 22514
rect 1192 22482 1224 22514
rect 1264 22482 1296 22514
rect 1336 22482 1368 22514
rect 1408 22482 1440 22514
rect 1480 22482 1512 22514
rect 1552 22482 1584 22514
rect 1624 22482 1656 22514
rect 1696 22482 1728 22514
rect 1768 22482 1800 22514
rect 1840 22482 1872 22514
rect 1912 22482 1944 22514
rect 1984 22482 2016 22514
rect 2056 22482 2088 22514
rect 2128 22482 2160 22514
rect 2200 22482 2232 22514
rect 2272 22482 2304 22514
rect 2344 22482 2376 22514
rect 2416 22482 2448 22514
rect 2488 22482 2520 22514
rect 2560 22482 2592 22514
rect 2632 22482 2664 22514
rect 2704 22482 2736 22514
rect 2776 22482 2808 22514
rect 2848 22482 2880 22514
rect 2920 22482 2952 22514
rect 2992 22482 3024 22514
rect 3064 22482 3096 22514
rect 3136 22482 3168 22514
rect 3208 22482 3240 22514
rect 3280 22482 3312 22514
rect 3352 22482 3384 22514
rect 3424 22482 3456 22514
rect 3496 22482 3528 22514
rect 3568 22482 3600 22514
rect 3640 22482 3672 22514
rect 3712 22482 3744 22514
rect 3784 22482 3816 22514
rect 3856 22482 3888 22514
rect 112 22410 144 22442
rect 184 22410 216 22442
rect 256 22410 288 22442
rect 328 22410 360 22442
rect 400 22410 432 22442
rect 472 22410 504 22442
rect 544 22410 576 22442
rect 616 22410 648 22442
rect 688 22410 720 22442
rect 760 22410 792 22442
rect 832 22410 864 22442
rect 904 22410 936 22442
rect 976 22410 1008 22442
rect 1048 22410 1080 22442
rect 1120 22410 1152 22442
rect 1192 22410 1224 22442
rect 1264 22410 1296 22442
rect 1336 22410 1368 22442
rect 1408 22410 1440 22442
rect 1480 22410 1512 22442
rect 1552 22410 1584 22442
rect 1624 22410 1656 22442
rect 1696 22410 1728 22442
rect 1768 22410 1800 22442
rect 1840 22410 1872 22442
rect 1912 22410 1944 22442
rect 1984 22410 2016 22442
rect 2056 22410 2088 22442
rect 2128 22410 2160 22442
rect 2200 22410 2232 22442
rect 2272 22410 2304 22442
rect 2344 22410 2376 22442
rect 2416 22410 2448 22442
rect 2488 22410 2520 22442
rect 2560 22410 2592 22442
rect 2632 22410 2664 22442
rect 2704 22410 2736 22442
rect 2776 22410 2808 22442
rect 2848 22410 2880 22442
rect 2920 22410 2952 22442
rect 2992 22410 3024 22442
rect 3064 22410 3096 22442
rect 3136 22410 3168 22442
rect 3208 22410 3240 22442
rect 3280 22410 3312 22442
rect 3352 22410 3384 22442
rect 3424 22410 3456 22442
rect 3496 22410 3528 22442
rect 3568 22410 3600 22442
rect 3640 22410 3672 22442
rect 3712 22410 3744 22442
rect 3784 22410 3816 22442
rect 3856 22410 3888 22442
rect 112 22338 144 22370
rect 184 22338 216 22370
rect 256 22338 288 22370
rect 328 22338 360 22370
rect 400 22338 432 22370
rect 472 22338 504 22370
rect 544 22338 576 22370
rect 616 22338 648 22370
rect 688 22338 720 22370
rect 760 22338 792 22370
rect 832 22338 864 22370
rect 904 22338 936 22370
rect 976 22338 1008 22370
rect 1048 22338 1080 22370
rect 1120 22338 1152 22370
rect 1192 22338 1224 22370
rect 1264 22338 1296 22370
rect 1336 22338 1368 22370
rect 1408 22338 1440 22370
rect 1480 22338 1512 22370
rect 1552 22338 1584 22370
rect 1624 22338 1656 22370
rect 1696 22338 1728 22370
rect 1768 22338 1800 22370
rect 1840 22338 1872 22370
rect 1912 22338 1944 22370
rect 1984 22338 2016 22370
rect 2056 22338 2088 22370
rect 2128 22338 2160 22370
rect 2200 22338 2232 22370
rect 2272 22338 2304 22370
rect 2344 22338 2376 22370
rect 2416 22338 2448 22370
rect 2488 22338 2520 22370
rect 2560 22338 2592 22370
rect 2632 22338 2664 22370
rect 2704 22338 2736 22370
rect 2776 22338 2808 22370
rect 2848 22338 2880 22370
rect 2920 22338 2952 22370
rect 2992 22338 3024 22370
rect 3064 22338 3096 22370
rect 3136 22338 3168 22370
rect 3208 22338 3240 22370
rect 3280 22338 3312 22370
rect 3352 22338 3384 22370
rect 3424 22338 3456 22370
rect 3496 22338 3528 22370
rect 3568 22338 3600 22370
rect 3640 22338 3672 22370
rect 3712 22338 3744 22370
rect 3784 22338 3816 22370
rect 3856 22338 3888 22370
rect 112 22266 144 22298
rect 184 22266 216 22298
rect 256 22266 288 22298
rect 328 22266 360 22298
rect 400 22266 432 22298
rect 472 22266 504 22298
rect 544 22266 576 22298
rect 616 22266 648 22298
rect 688 22266 720 22298
rect 760 22266 792 22298
rect 832 22266 864 22298
rect 904 22266 936 22298
rect 976 22266 1008 22298
rect 1048 22266 1080 22298
rect 1120 22266 1152 22298
rect 1192 22266 1224 22298
rect 1264 22266 1296 22298
rect 1336 22266 1368 22298
rect 1408 22266 1440 22298
rect 1480 22266 1512 22298
rect 1552 22266 1584 22298
rect 1624 22266 1656 22298
rect 1696 22266 1728 22298
rect 1768 22266 1800 22298
rect 1840 22266 1872 22298
rect 1912 22266 1944 22298
rect 1984 22266 2016 22298
rect 2056 22266 2088 22298
rect 2128 22266 2160 22298
rect 2200 22266 2232 22298
rect 2272 22266 2304 22298
rect 2344 22266 2376 22298
rect 2416 22266 2448 22298
rect 2488 22266 2520 22298
rect 2560 22266 2592 22298
rect 2632 22266 2664 22298
rect 2704 22266 2736 22298
rect 2776 22266 2808 22298
rect 2848 22266 2880 22298
rect 2920 22266 2952 22298
rect 2992 22266 3024 22298
rect 3064 22266 3096 22298
rect 3136 22266 3168 22298
rect 3208 22266 3240 22298
rect 3280 22266 3312 22298
rect 3352 22266 3384 22298
rect 3424 22266 3456 22298
rect 3496 22266 3528 22298
rect 3568 22266 3600 22298
rect 3640 22266 3672 22298
rect 3712 22266 3744 22298
rect 3784 22266 3816 22298
rect 3856 22266 3888 22298
rect 112 22194 144 22226
rect 184 22194 216 22226
rect 256 22194 288 22226
rect 328 22194 360 22226
rect 400 22194 432 22226
rect 472 22194 504 22226
rect 544 22194 576 22226
rect 616 22194 648 22226
rect 688 22194 720 22226
rect 760 22194 792 22226
rect 832 22194 864 22226
rect 904 22194 936 22226
rect 976 22194 1008 22226
rect 1048 22194 1080 22226
rect 1120 22194 1152 22226
rect 1192 22194 1224 22226
rect 1264 22194 1296 22226
rect 1336 22194 1368 22226
rect 1408 22194 1440 22226
rect 1480 22194 1512 22226
rect 1552 22194 1584 22226
rect 1624 22194 1656 22226
rect 1696 22194 1728 22226
rect 1768 22194 1800 22226
rect 1840 22194 1872 22226
rect 1912 22194 1944 22226
rect 1984 22194 2016 22226
rect 2056 22194 2088 22226
rect 2128 22194 2160 22226
rect 2200 22194 2232 22226
rect 2272 22194 2304 22226
rect 2344 22194 2376 22226
rect 2416 22194 2448 22226
rect 2488 22194 2520 22226
rect 2560 22194 2592 22226
rect 2632 22194 2664 22226
rect 2704 22194 2736 22226
rect 2776 22194 2808 22226
rect 2848 22194 2880 22226
rect 2920 22194 2952 22226
rect 2992 22194 3024 22226
rect 3064 22194 3096 22226
rect 3136 22194 3168 22226
rect 3208 22194 3240 22226
rect 3280 22194 3312 22226
rect 3352 22194 3384 22226
rect 3424 22194 3456 22226
rect 3496 22194 3528 22226
rect 3568 22194 3600 22226
rect 3640 22194 3672 22226
rect 3712 22194 3744 22226
rect 3784 22194 3816 22226
rect 3856 22194 3888 22226
rect 112 22122 144 22154
rect 184 22122 216 22154
rect 256 22122 288 22154
rect 328 22122 360 22154
rect 400 22122 432 22154
rect 472 22122 504 22154
rect 544 22122 576 22154
rect 616 22122 648 22154
rect 688 22122 720 22154
rect 760 22122 792 22154
rect 832 22122 864 22154
rect 904 22122 936 22154
rect 976 22122 1008 22154
rect 1048 22122 1080 22154
rect 1120 22122 1152 22154
rect 1192 22122 1224 22154
rect 1264 22122 1296 22154
rect 1336 22122 1368 22154
rect 1408 22122 1440 22154
rect 1480 22122 1512 22154
rect 1552 22122 1584 22154
rect 1624 22122 1656 22154
rect 1696 22122 1728 22154
rect 1768 22122 1800 22154
rect 1840 22122 1872 22154
rect 1912 22122 1944 22154
rect 1984 22122 2016 22154
rect 2056 22122 2088 22154
rect 2128 22122 2160 22154
rect 2200 22122 2232 22154
rect 2272 22122 2304 22154
rect 2344 22122 2376 22154
rect 2416 22122 2448 22154
rect 2488 22122 2520 22154
rect 2560 22122 2592 22154
rect 2632 22122 2664 22154
rect 2704 22122 2736 22154
rect 2776 22122 2808 22154
rect 2848 22122 2880 22154
rect 2920 22122 2952 22154
rect 2992 22122 3024 22154
rect 3064 22122 3096 22154
rect 3136 22122 3168 22154
rect 3208 22122 3240 22154
rect 3280 22122 3312 22154
rect 3352 22122 3384 22154
rect 3424 22122 3456 22154
rect 3496 22122 3528 22154
rect 3568 22122 3600 22154
rect 3640 22122 3672 22154
rect 3712 22122 3744 22154
rect 3784 22122 3816 22154
rect 3856 22122 3888 22154
rect 112 22050 144 22082
rect 184 22050 216 22082
rect 256 22050 288 22082
rect 328 22050 360 22082
rect 400 22050 432 22082
rect 472 22050 504 22082
rect 544 22050 576 22082
rect 616 22050 648 22082
rect 688 22050 720 22082
rect 760 22050 792 22082
rect 832 22050 864 22082
rect 904 22050 936 22082
rect 976 22050 1008 22082
rect 1048 22050 1080 22082
rect 1120 22050 1152 22082
rect 1192 22050 1224 22082
rect 1264 22050 1296 22082
rect 1336 22050 1368 22082
rect 1408 22050 1440 22082
rect 1480 22050 1512 22082
rect 1552 22050 1584 22082
rect 1624 22050 1656 22082
rect 1696 22050 1728 22082
rect 1768 22050 1800 22082
rect 1840 22050 1872 22082
rect 1912 22050 1944 22082
rect 1984 22050 2016 22082
rect 2056 22050 2088 22082
rect 2128 22050 2160 22082
rect 2200 22050 2232 22082
rect 2272 22050 2304 22082
rect 2344 22050 2376 22082
rect 2416 22050 2448 22082
rect 2488 22050 2520 22082
rect 2560 22050 2592 22082
rect 2632 22050 2664 22082
rect 2704 22050 2736 22082
rect 2776 22050 2808 22082
rect 2848 22050 2880 22082
rect 2920 22050 2952 22082
rect 2992 22050 3024 22082
rect 3064 22050 3096 22082
rect 3136 22050 3168 22082
rect 3208 22050 3240 22082
rect 3280 22050 3312 22082
rect 3352 22050 3384 22082
rect 3424 22050 3456 22082
rect 3496 22050 3528 22082
rect 3568 22050 3600 22082
rect 3640 22050 3672 22082
rect 3712 22050 3744 22082
rect 3784 22050 3816 22082
rect 3856 22050 3888 22082
rect 112 21978 144 22010
rect 184 21978 216 22010
rect 256 21978 288 22010
rect 328 21978 360 22010
rect 400 21978 432 22010
rect 472 21978 504 22010
rect 544 21978 576 22010
rect 616 21978 648 22010
rect 688 21978 720 22010
rect 760 21978 792 22010
rect 832 21978 864 22010
rect 904 21978 936 22010
rect 976 21978 1008 22010
rect 1048 21978 1080 22010
rect 1120 21978 1152 22010
rect 1192 21978 1224 22010
rect 1264 21978 1296 22010
rect 1336 21978 1368 22010
rect 1408 21978 1440 22010
rect 1480 21978 1512 22010
rect 1552 21978 1584 22010
rect 1624 21978 1656 22010
rect 1696 21978 1728 22010
rect 1768 21978 1800 22010
rect 1840 21978 1872 22010
rect 1912 21978 1944 22010
rect 1984 21978 2016 22010
rect 2056 21978 2088 22010
rect 2128 21978 2160 22010
rect 2200 21978 2232 22010
rect 2272 21978 2304 22010
rect 2344 21978 2376 22010
rect 2416 21978 2448 22010
rect 2488 21978 2520 22010
rect 2560 21978 2592 22010
rect 2632 21978 2664 22010
rect 2704 21978 2736 22010
rect 2776 21978 2808 22010
rect 2848 21978 2880 22010
rect 2920 21978 2952 22010
rect 2992 21978 3024 22010
rect 3064 21978 3096 22010
rect 3136 21978 3168 22010
rect 3208 21978 3240 22010
rect 3280 21978 3312 22010
rect 3352 21978 3384 22010
rect 3424 21978 3456 22010
rect 3496 21978 3528 22010
rect 3568 21978 3600 22010
rect 3640 21978 3672 22010
rect 3712 21978 3744 22010
rect 3784 21978 3816 22010
rect 3856 21978 3888 22010
rect 112 21906 144 21938
rect 184 21906 216 21938
rect 256 21906 288 21938
rect 328 21906 360 21938
rect 400 21906 432 21938
rect 472 21906 504 21938
rect 544 21906 576 21938
rect 616 21906 648 21938
rect 688 21906 720 21938
rect 760 21906 792 21938
rect 832 21906 864 21938
rect 904 21906 936 21938
rect 976 21906 1008 21938
rect 1048 21906 1080 21938
rect 1120 21906 1152 21938
rect 1192 21906 1224 21938
rect 1264 21906 1296 21938
rect 1336 21906 1368 21938
rect 1408 21906 1440 21938
rect 1480 21906 1512 21938
rect 1552 21906 1584 21938
rect 1624 21906 1656 21938
rect 1696 21906 1728 21938
rect 1768 21906 1800 21938
rect 1840 21906 1872 21938
rect 1912 21906 1944 21938
rect 1984 21906 2016 21938
rect 2056 21906 2088 21938
rect 2128 21906 2160 21938
rect 2200 21906 2232 21938
rect 2272 21906 2304 21938
rect 2344 21906 2376 21938
rect 2416 21906 2448 21938
rect 2488 21906 2520 21938
rect 2560 21906 2592 21938
rect 2632 21906 2664 21938
rect 2704 21906 2736 21938
rect 2776 21906 2808 21938
rect 2848 21906 2880 21938
rect 2920 21906 2952 21938
rect 2992 21906 3024 21938
rect 3064 21906 3096 21938
rect 3136 21906 3168 21938
rect 3208 21906 3240 21938
rect 3280 21906 3312 21938
rect 3352 21906 3384 21938
rect 3424 21906 3456 21938
rect 3496 21906 3528 21938
rect 3568 21906 3600 21938
rect 3640 21906 3672 21938
rect 3712 21906 3744 21938
rect 3784 21906 3816 21938
rect 3856 21906 3888 21938
rect 112 21834 144 21866
rect 184 21834 216 21866
rect 256 21834 288 21866
rect 328 21834 360 21866
rect 400 21834 432 21866
rect 472 21834 504 21866
rect 544 21834 576 21866
rect 616 21834 648 21866
rect 688 21834 720 21866
rect 760 21834 792 21866
rect 832 21834 864 21866
rect 904 21834 936 21866
rect 976 21834 1008 21866
rect 1048 21834 1080 21866
rect 1120 21834 1152 21866
rect 1192 21834 1224 21866
rect 1264 21834 1296 21866
rect 1336 21834 1368 21866
rect 1408 21834 1440 21866
rect 1480 21834 1512 21866
rect 1552 21834 1584 21866
rect 1624 21834 1656 21866
rect 1696 21834 1728 21866
rect 1768 21834 1800 21866
rect 1840 21834 1872 21866
rect 1912 21834 1944 21866
rect 1984 21834 2016 21866
rect 2056 21834 2088 21866
rect 2128 21834 2160 21866
rect 2200 21834 2232 21866
rect 2272 21834 2304 21866
rect 2344 21834 2376 21866
rect 2416 21834 2448 21866
rect 2488 21834 2520 21866
rect 2560 21834 2592 21866
rect 2632 21834 2664 21866
rect 2704 21834 2736 21866
rect 2776 21834 2808 21866
rect 2848 21834 2880 21866
rect 2920 21834 2952 21866
rect 2992 21834 3024 21866
rect 3064 21834 3096 21866
rect 3136 21834 3168 21866
rect 3208 21834 3240 21866
rect 3280 21834 3312 21866
rect 3352 21834 3384 21866
rect 3424 21834 3456 21866
rect 3496 21834 3528 21866
rect 3568 21834 3600 21866
rect 3640 21834 3672 21866
rect 3712 21834 3744 21866
rect 3784 21834 3816 21866
rect 3856 21834 3888 21866
rect 112 21762 144 21794
rect 184 21762 216 21794
rect 256 21762 288 21794
rect 328 21762 360 21794
rect 400 21762 432 21794
rect 472 21762 504 21794
rect 544 21762 576 21794
rect 616 21762 648 21794
rect 688 21762 720 21794
rect 760 21762 792 21794
rect 832 21762 864 21794
rect 904 21762 936 21794
rect 976 21762 1008 21794
rect 1048 21762 1080 21794
rect 1120 21762 1152 21794
rect 1192 21762 1224 21794
rect 1264 21762 1296 21794
rect 1336 21762 1368 21794
rect 1408 21762 1440 21794
rect 1480 21762 1512 21794
rect 1552 21762 1584 21794
rect 1624 21762 1656 21794
rect 1696 21762 1728 21794
rect 1768 21762 1800 21794
rect 1840 21762 1872 21794
rect 1912 21762 1944 21794
rect 1984 21762 2016 21794
rect 2056 21762 2088 21794
rect 2128 21762 2160 21794
rect 2200 21762 2232 21794
rect 2272 21762 2304 21794
rect 2344 21762 2376 21794
rect 2416 21762 2448 21794
rect 2488 21762 2520 21794
rect 2560 21762 2592 21794
rect 2632 21762 2664 21794
rect 2704 21762 2736 21794
rect 2776 21762 2808 21794
rect 2848 21762 2880 21794
rect 2920 21762 2952 21794
rect 2992 21762 3024 21794
rect 3064 21762 3096 21794
rect 3136 21762 3168 21794
rect 3208 21762 3240 21794
rect 3280 21762 3312 21794
rect 3352 21762 3384 21794
rect 3424 21762 3456 21794
rect 3496 21762 3528 21794
rect 3568 21762 3600 21794
rect 3640 21762 3672 21794
rect 3712 21762 3744 21794
rect 3784 21762 3816 21794
rect 3856 21762 3888 21794
rect 112 21690 144 21722
rect 184 21690 216 21722
rect 256 21690 288 21722
rect 328 21690 360 21722
rect 400 21690 432 21722
rect 472 21690 504 21722
rect 544 21690 576 21722
rect 616 21690 648 21722
rect 688 21690 720 21722
rect 760 21690 792 21722
rect 832 21690 864 21722
rect 904 21690 936 21722
rect 976 21690 1008 21722
rect 1048 21690 1080 21722
rect 1120 21690 1152 21722
rect 1192 21690 1224 21722
rect 1264 21690 1296 21722
rect 1336 21690 1368 21722
rect 1408 21690 1440 21722
rect 1480 21690 1512 21722
rect 1552 21690 1584 21722
rect 1624 21690 1656 21722
rect 1696 21690 1728 21722
rect 1768 21690 1800 21722
rect 1840 21690 1872 21722
rect 1912 21690 1944 21722
rect 1984 21690 2016 21722
rect 2056 21690 2088 21722
rect 2128 21690 2160 21722
rect 2200 21690 2232 21722
rect 2272 21690 2304 21722
rect 2344 21690 2376 21722
rect 2416 21690 2448 21722
rect 2488 21690 2520 21722
rect 2560 21690 2592 21722
rect 2632 21690 2664 21722
rect 2704 21690 2736 21722
rect 2776 21690 2808 21722
rect 2848 21690 2880 21722
rect 2920 21690 2952 21722
rect 2992 21690 3024 21722
rect 3064 21690 3096 21722
rect 3136 21690 3168 21722
rect 3208 21690 3240 21722
rect 3280 21690 3312 21722
rect 3352 21690 3384 21722
rect 3424 21690 3456 21722
rect 3496 21690 3528 21722
rect 3568 21690 3600 21722
rect 3640 21690 3672 21722
rect 3712 21690 3744 21722
rect 3784 21690 3816 21722
rect 3856 21690 3888 21722
rect 112 21618 144 21650
rect 184 21618 216 21650
rect 256 21618 288 21650
rect 328 21618 360 21650
rect 400 21618 432 21650
rect 472 21618 504 21650
rect 544 21618 576 21650
rect 616 21618 648 21650
rect 688 21618 720 21650
rect 760 21618 792 21650
rect 832 21618 864 21650
rect 904 21618 936 21650
rect 976 21618 1008 21650
rect 1048 21618 1080 21650
rect 1120 21618 1152 21650
rect 1192 21618 1224 21650
rect 1264 21618 1296 21650
rect 1336 21618 1368 21650
rect 1408 21618 1440 21650
rect 1480 21618 1512 21650
rect 1552 21618 1584 21650
rect 1624 21618 1656 21650
rect 1696 21618 1728 21650
rect 1768 21618 1800 21650
rect 1840 21618 1872 21650
rect 1912 21618 1944 21650
rect 1984 21618 2016 21650
rect 2056 21618 2088 21650
rect 2128 21618 2160 21650
rect 2200 21618 2232 21650
rect 2272 21618 2304 21650
rect 2344 21618 2376 21650
rect 2416 21618 2448 21650
rect 2488 21618 2520 21650
rect 2560 21618 2592 21650
rect 2632 21618 2664 21650
rect 2704 21618 2736 21650
rect 2776 21618 2808 21650
rect 2848 21618 2880 21650
rect 2920 21618 2952 21650
rect 2992 21618 3024 21650
rect 3064 21618 3096 21650
rect 3136 21618 3168 21650
rect 3208 21618 3240 21650
rect 3280 21618 3312 21650
rect 3352 21618 3384 21650
rect 3424 21618 3456 21650
rect 3496 21618 3528 21650
rect 3568 21618 3600 21650
rect 3640 21618 3672 21650
rect 3712 21618 3744 21650
rect 3784 21618 3816 21650
rect 3856 21618 3888 21650
rect 112 21546 144 21578
rect 184 21546 216 21578
rect 256 21546 288 21578
rect 328 21546 360 21578
rect 400 21546 432 21578
rect 472 21546 504 21578
rect 544 21546 576 21578
rect 616 21546 648 21578
rect 688 21546 720 21578
rect 760 21546 792 21578
rect 832 21546 864 21578
rect 904 21546 936 21578
rect 976 21546 1008 21578
rect 1048 21546 1080 21578
rect 1120 21546 1152 21578
rect 1192 21546 1224 21578
rect 1264 21546 1296 21578
rect 1336 21546 1368 21578
rect 1408 21546 1440 21578
rect 1480 21546 1512 21578
rect 1552 21546 1584 21578
rect 1624 21546 1656 21578
rect 1696 21546 1728 21578
rect 1768 21546 1800 21578
rect 1840 21546 1872 21578
rect 1912 21546 1944 21578
rect 1984 21546 2016 21578
rect 2056 21546 2088 21578
rect 2128 21546 2160 21578
rect 2200 21546 2232 21578
rect 2272 21546 2304 21578
rect 2344 21546 2376 21578
rect 2416 21546 2448 21578
rect 2488 21546 2520 21578
rect 2560 21546 2592 21578
rect 2632 21546 2664 21578
rect 2704 21546 2736 21578
rect 2776 21546 2808 21578
rect 2848 21546 2880 21578
rect 2920 21546 2952 21578
rect 2992 21546 3024 21578
rect 3064 21546 3096 21578
rect 3136 21546 3168 21578
rect 3208 21546 3240 21578
rect 3280 21546 3312 21578
rect 3352 21546 3384 21578
rect 3424 21546 3456 21578
rect 3496 21546 3528 21578
rect 3568 21546 3600 21578
rect 3640 21546 3672 21578
rect 3712 21546 3744 21578
rect 3784 21546 3816 21578
rect 3856 21546 3888 21578
rect 112 21474 144 21506
rect 184 21474 216 21506
rect 256 21474 288 21506
rect 328 21474 360 21506
rect 400 21474 432 21506
rect 472 21474 504 21506
rect 544 21474 576 21506
rect 616 21474 648 21506
rect 688 21474 720 21506
rect 760 21474 792 21506
rect 832 21474 864 21506
rect 904 21474 936 21506
rect 976 21474 1008 21506
rect 1048 21474 1080 21506
rect 1120 21474 1152 21506
rect 1192 21474 1224 21506
rect 1264 21474 1296 21506
rect 1336 21474 1368 21506
rect 1408 21474 1440 21506
rect 1480 21474 1512 21506
rect 1552 21474 1584 21506
rect 1624 21474 1656 21506
rect 1696 21474 1728 21506
rect 1768 21474 1800 21506
rect 1840 21474 1872 21506
rect 1912 21474 1944 21506
rect 1984 21474 2016 21506
rect 2056 21474 2088 21506
rect 2128 21474 2160 21506
rect 2200 21474 2232 21506
rect 2272 21474 2304 21506
rect 2344 21474 2376 21506
rect 2416 21474 2448 21506
rect 2488 21474 2520 21506
rect 2560 21474 2592 21506
rect 2632 21474 2664 21506
rect 2704 21474 2736 21506
rect 2776 21474 2808 21506
rect 2848 21474 2880 21506
rect 2920 21474 2952 21506
rect 2992 21474 3024 21506
rect 3064 21474 3096 21506
rect 3136 21474 3168 21506
rect 3208 21474 3240 21506
rect 3280 21474 3312 21506
rect 3352 21474 3384 21506
rect 3424 21474 3456 21506
rect 3496 21474 3528 21506
rect 3568 21474 3600 21506
rect 3640 21474 3672 21506
rect 3712 21474 3744 21506
rect 3784 21474 3816 21506
rect 3856 21474 3888 21506
rect 112 21402 144 21434
rect 184 21402 216 21434
rect 256 21402 288 21434
rect 328 21402 360 21434
rect 400 21402 432 21434
rect 472 21402 504 21434
rect 544 21402 576 21434
rect 616 21402 648 21434
rect 688 21402 720 21434
rect 760 21402 792 21434
rect 832 21402 864 21434
rect 904 21402 936 21434
rect 976 21402 1008 21434
rect 1048 21402 1080 21434
rect 1120 21402 1152 21434
rect 1192 21402 1224 21434
rect 1264 21402 1296 21434
rect 1336 21402 1368 21434
rect 1408 21402 1440 21434
rect 1480 21402 1512 21434
rect 1552 21402 1584 21434
rect 1624 21402 1656 21434
rect 1696 21402 1728 21434
rect 1768 21402 1800 21434
rect 1840 21402 1872 21434
rect 1912 21402 1944 21434
rect 1984 21402 2016 21434
rect 2056 21402 2088 21434
rect 2128 21402 2160 21434
rect 2200 21402 2232 21434
rect 2272 21402 2304 21434
rect 2344 21402 2376 21434
rect 2416 21402 2448 21434
rect 2488 21402 2520 21434
rect 2560 21402 2592 21434
rect 2632 21402 2664 21434
rect 2704 21402 2736 21434
rect 2776 21402 2808 21434
rect 2848 21402 2880 21434
rect 2920 21402 2952 21434
rect 2992 21402 3024 21434
rect 3064 21402 3096 21434
rect 3136 21402 3168 21434
rect 3208 21402 3240 21434
rect 3280 21402 3312 21434
rect 3352 21402 3384 21434
rect 3424 21402 3456 21434
rect 3496 21402 3528 21434
rect 3568 21402 3600 21434
rect 3640 21402 3672 21434
rect 3712 21402 3744 21434
rect 3784 21402 3816 21434
rect 3856 21402 3888 21434
rect 112 21330 144 21362
rect 184 21330 216 21362
rect 256 21330 288 21362
rect 328 21330 360 21362
rect 400 21330 432 21362
rect 472 21330 504 21362
rect 544 21330 576 21362
rect 616 21330 648 21362
rect 688 21330 720 21362
rect 760 21330 792 21362
rect 832 21330 864 21362
rect 904 21330 936 21362
rect 976 21330 1008 21362
rect 1048 21330 1080 21362
rect 1120 21330 1152 21362
rect 1192 21330 1224 21362
rect 1264 21330 1296 21362
rect 1336 21330 1368 21362
rect 1408 21330 1440 21362
rect 1480 21330 1512 21362
rect 1552 21330 1584 21362
rect 1624 21330 1656 21362
rect 1696 21330 1728 21362
rect 1768 21330 1800 21362
rect 1840 21330 1872 21362
rect 1912 21330 1944 21362
rect 1984 21330 2016 21362
rect 2056 21330 2088 21362
rect 2128 21330 2160 21362
rect 2200 21330 2232 21362
rect 2272 21330 2304 21362
rect 2344 21330 2376 21362
rect 2416 21330 2448 21362
rect 2488 21330 2520 21362
rect 2560 21330 2592 21362
rect 2632 21330 2664 21362
rect 2704 21330 2736 21362
rect 2776 21330 2808 21362
rect 2848 21330 2880 21362
rect 2920 21330 2952 21362
rect 2992 21330 3024 21362
rect 3064 21330 3096 21362
rect 3136 21330 3168 21362
rect 3208 21330 3240 21362
rect 3280 21330 3312 21362
rect 3352 21330 3384 21362
rect 3424 21330 3456 21362
rect 3496 21330 3528 21362
rect 3568 21330 3600 21362
rect 3640 21330 3672 21362
rect 3712 21330 3744 21362
rect 3784 21330 3816 21362
rect 3856 21330 3888 21362
rect 112 21258 144 21290
rect 184 21258 216 21290
rect 256 21258 288 21290
rect 328 21258 360 21290
rect 400 21258 432 21290
rect 472 21258 504 21290
rect 544 21258 576 21290
rect 616 21258 648 21290
rect 688 21258 720 21290
rect 760 21258 792 21290
rect 832 21258 864 21290
rect 904 21258 936 21290
rect 976 21258 1008 21290
rect 1048 21258 1080 21290
rect 1120 21258 1152 21290
rect 1192 21258 1224 21290
rect 1264 21258 1296 21290
rect 1336 21258 1368 21290
rect 1408 21258 1440 21290
rect 1480 21258 1512 21290
rect 1552 21258 1584 21290
rect 1624 21258 1656 21290
rect 1696 21258 1728 21290
rect 1768 21258 1800 21290
rect 1840 21258 1872 21290
rect 1912 21258 1944 21290
rect 1984 21258 2016 21290
rect 2056 21258 2088 21290
rect 2128 21258 2160 21290
rect 2200 21258 2232 21290
rect 2272 21258 2304 21290
rect 2344 21258 2376 21290
rect 2416 21258 2448 21290
rect 2488 21258 2520 21290
rect 2560 21258 2592 21290
rect 2632 21258 2664 21290
rect 2704 21258 2736 21290
rect 2776 21258 2808 21290
rect 2848 21258 2880 21290
rect 2920 21258 2952 21290
rect 2992 21258 3024 21290
rect 3064 21258 3096 21290
rect 3136 21258 3168 21290
rect 3208 21258 3240 21290
rect 3280 21258 3312 21290
rect 3352 21258 3384 21290
rect 3424 21258 3456 21290
rect 3496 21258 3528 21290
rect 3568 21258 3600 21290
rect 3640 21258 3672 21290
rect 3712 21258 3744 21290
rect 3784 21258 3816 21290
rect 3856 21258 3888 21290
rect 112 21186 144 21218
rect 184 21186 216 21218
rect 256 21186 288 21218
rect 328 21186 360 21218
rect 400 21186 432 21218
rect 472 21186 504 21218
rect 544 21186 576 21218
rect 616 21186 648 21218
rect 688 21186 720 21218
rect 760 21186 792 21218
rect 832 21186 864 21218
rect 904 21186 936 21218
rect 976 21186 1008 21218
rect 1048 21186 1080 21218
rect 1120 21186 1152 21218
rect 1192 21186 1224 21218
rect 1264 21186 1296 21218
rect 1336 21186 1368 21218
rect 1408 21186 1440 21218
rect 1480 21186 1512 21218
rect 1552 21186 1584 21218
rect 1624 21186 1656 21218
rect 1696 21186 1728 21218
rect 1768 21186 1800 21218
rect 1840 21186 1872 21218
rect 1912 21186 1944 21218
rect 1984 21186 2016 21218
rect 2056 21186 2088 21218
rect 2128 21186 2160 21218
rect 2200 21186 2232 21218
rect 2272 21186 2304 21218
rect 2344 21186 2376 21218
rect 2416 21186 2448 21218
rect 2488 21186 2520 21218
rect 2560 21186 2592 21218
rect 2632 21186 2664 21218
rect 2704 21186 2736 21218
rect 2776 21186 2808 21218
rect 2848 21186 2880 21218
rect 2920 21186 2952 21218
rect 2992 21186 3024 21218
rect 3064 21186 3096 21218
rect 3136 21186 3168 21218
rect 3208 21186 3240 21218
rect 3280 21186 3312 21218
rect 3352 21186 3384 21218
rect 3424 21186 3456 21218
rect 3496 21186 3528 21218
rect 3568 21186 3600 21218
rect 3640 21186 3672 21218
rect 3712 21186 3744 21218
rect 3784 21186 3816 21218
rect 3856 21186 3888 21218
rect 112 21114 144 21146
rect 184 21114 216 21146
rect 256 21114 288 21146
rect 328 21114 360 21146
rect 400 21114 432 21146
rect 472 21114 504 21146
rect 544 21114 576 21146
rect 616 21114 648 21146
rect 688 21114 720 21146
rect 760 21114 792 21146
rect 832 21114 864 21146
rect 904 21114 936 21146
rect 976 21114 1008 21146
rect 1048 21114 1080 21146
rect 1120 21114 1152 21146
rect 1192 21114 1224 21146
rect 1264 21114 1296 21146
rect 1336 21114 1368 21146
rect 1408 21114 1440 21146
rect 1480 21114 1512 21146
rect 1552 21114 1584 21146
rect 1624 21114 1656 21146
rect 1696 21114 1728 21146
rect 1768 21114 1800 21146
rect 1840 21114 1872 21146
rect 1912 21114 1944 21146
rect 1984 21114 2016 21146
rect 2056 21114 2088 21146
rect 2128 21114 2160 21146
rect 2200 21114 2232 21146
rect 2272 21114 2304 21146
rect 2344 21114 2376 21146
rect 2416 21114 2448 21146
rect 2488 21114 2520 21146
rect 2560 21114 2592 21146
rect 2632 21114 2664 21146
rect 2704 21114 2736 21146
rect 2776 21114 2808 21146
rect 2848 21114 2880 21146
rect 2920 21114 2952 21146
rect 2992 21114 3024 21146
rect 3064 21114 3096 21146
rect 3136 21114 3168 21146
rect 3208 21114 3240 21146
rect 3280 21114 3312 21146
rect 3352 21114 3384 21146
rect 3424 21114 3456 21146
rect 3496 21114 3528 21146
rect 3568 21114 3600 21146
rect 3640 21114 3672 21146
rect 3712 21114 3744 21146
rect 3784 21114 3816 21146
rect 3856 21114 3888 21146
rect 112 21042 144 21074
rect 184 21042 216 21074
rect 256 21042 288 21074
rect 328 21042 360 21074
rect 400 21042 432 21074
rect 472 21042 504 21074
rect 544 21042 576 21074
rect 616 21042 648 21074
rect 688 21042 720 21074
rect 760 21042 792 21074
rect 832 21042 864 21074
rect 904 21042 936 21074
rect 976 21042 1008 21074
rect 1048 21042 1080 21074
rect 1120 21042 1152 21074
rect 1192 21042 1224 21074
rect 1264 21042 1296 21074
rect 1336 21042 1368 21074
rect 1408 21042 1440 21074
rect 1480 21042 1512 21074
rect 1552 21042 1584 21074
rect 1624 21042 1656 21074
rect 1696 21042 1728 21074
rect 1768 21042 1800 21074
rect 1840 21042 1872 21074
rect 1912 21042 1944 21074
rect 1984 21042 2016 21074
rect 2056 21042 2088 21074
rect 2128 21042 2160 21074
rect 2200 21042 2232 21074
rect 2272 21042 2304 21074
rect 2344 21042 2376 21074
rect 2416 21042 2448 21074
rect 2488 21042 2520 21074
rect 2560 21042 2592 21074
rect 2632 21042 2664 21074
rect 2704 21042 2736 21074
rect 2776 21042 2808 21074
rect 2848 21042 2880 21074
rect 2920 21042 2952 21074
rect 2992 21042 3024 21074
rect 3064 21042 3096 21074
rect 3136 21042 3168 21074
rect 3208 21042 3240 21074
rect 3280 21042 3312 21074
rect 3352 21042 3384 21074
rect 3424 21042 3456 21074
rect 3496 21042 3528 21074
rect 3568 21042 3600 21074
rect 3640 21042 3672 21074
rect 3712 21042 3744 21074
rect 3784 21042 3816 21074
rect 3856 21042 3888 21074
rect 112 20970 144 21002
rect 184 20970 216 21002
rect 256 20970 288 21002
rect 328 20970 360 21002
rect 400 20970 432 21002
rect 472 20970 504 21002
rect 544 20970 576 21002
rect 616 20970 648 21002
rect 688 20970 720 21002
rect 760 20970 792 21002
rect 832 20970 864 21002
rect 904 20970 936 21002
rect 976 20970 1008 21002
rect 1048 20970 1080 21002
rect 1120 20970 1152 21002
rect 1192 20970 1224 21002
rect 1264 20970 1296 21002
rect 1336 20970 1368 21002
rect 1408 20970 1440 21002
rect 1480 20970 1512 21002
rect 1552 20970 1584 21002
rect 1624 20970 1656 21002
rect 1696 20970 1728 21002
rect 1768 20970 1800 21002
rect 1840 20970 1872 21002
rect 1912 20970 1944 21002
rect 1984 20970 2016 21002
rect 2056 20970 2088 21002
rect 2128 20970 2160 21002
rect 2200 20970 2232 21002
rect 2272 20970 2304 21002
rect 2344 20970 2376 21002
rect 2416 20970 2448 21002
rect 2488 20970 2520 21002
rect 2560 20970 2592 21002
rect 2632 20970 2664 21002
rect 2704 20970 2736 21002
rect 2776 20970 2808 21002
rect 2848 20970 2880 21002
rect 2920 20970 2952 21002
rect 2992 20970 3024 21002
rect 3064 20970 3096 21002
rect 3136 20970 3168 21002
rect 3208 20970 3240 21002
rect 3280 20970 3312 21002
rect 3352 20970 3384 21002
rect 3424 20970 3456 21002
rect 3496 20970 3528 21002
rect 3568 20970 3600 21002
rect 3640 20970 3672 21002
rect 3712 20970 3744 21002
rect 3784 20970 3816 21002
rect 3856 20970 3888 21002
rect 112 20898 144 20930
rect 184 20898 216 20930
rect 256 20898 288 20930
rect 328 20898 360 20930
rect 400 20898 432 20930
rect 472 20898 504 20930
rect 544 20898 576 20930
rect 616 20898 648 20930
rect 688 20898 720 20930
rect 760 20898 792 20930
rect 832 20898 864 20930
rect 904 20898 936 20930
rect 976 20898 1008 20930
rect 1048 20898 1080 20930
rect 1120 20898 1152 20930
rect 1192 20898 1224 20930
rect 1264 20898 1296 20930
rect 1336 20898 1368 20930
rect 1408 20898 1440 20930
rect 1480 20898 1512 20930
rect 1552 20898 1584 20930
rect 1624 20898 1656 20930
rect 1696 20898 1728 20930
rect 1768 20898 1800 20930
rect 1840 20898 1872 20930
rect 1912 20898 1944 20930
rect 1984 20898 2016 20930
rect 2056 20898 2088 20930
rect 2128 20898 2160 20930
rect 2200 20898 2232 20930
rect 2272 20898 2304 20930
rect 2344 20898 2376 20930
rect 2416 20898 2448 20930
rect 2488 20898 2520 20930
rect 2560 20898 2592 20930
rect 2632 20898 2664 20930
rect 2704 20898 2736 20930
rect 2776 20898 2808 20930
rect 2848 20898 2880 20930
rect 2920 20898 2952 20930
rect 2992 20898 3024 20930
rect 3064 20898 3096 20930
rect 3136 20898 3168 20930
rect 3208 20898 3240 20930
rect 3280 20898 3312 20930
rect 3352 20898 3384 20930
rect 3424 20898 3456 20930
rect 3496 20898 3528 20930
rect 3568 20898 3600 20930
rect 3640 20898 3672 20930
rect 3712 20898 3744 20930
rect 3784 20898 3816 20930
rect 3856 20898 3888 20930
rect 112 20826 144 20858
rect 184 20826 216 20858
rect 256 20826 288 20858
rect 328 20826 360 20858
rect 400 20826 432 20858
rect 472 20826 504 20858
rect 544 20826 576 20858
rect 616 20826 648 20858
rect 688 20826 720 20858
rect 760 20826 792 20858
rect 832 20826 864 20858
rect 904 20826 936 20858
rect 976 20826 1008 20858
rect 1048 20826 1080 20858
rect 1120 20826 1152 20858
rect 1192 20826 1224 20858
rect 1264 20826 1296 20858
rect 1336 20826 1368 20858
rect 1408 20826 1440 20858
rect 1480 20826 1512 20858
rect 1552 20826 1584 20858
rect 1624 20826 1656 20858
rect 1696 20826 1728 20858
rect 1768 20826 1800 20858
rect 1840 20826 1872 20858
rect 1912 20826 1944 20858
rect 1984 20826 2016 20858
rect 2056 20826 2088 20858
rect 2128 20826 2160 20858
rect 2200 20826 2232 20858
rect 2272 20826 2304 20858
rect 2344 20826 2376 20858
rect 2416 20826 2448 20858
rect 2488 20826 2520 20858
rect 2560 20826 2592 20858
rect 2632 20826 2664 20858
rect 2704 20826 2736 20858
rect 2776 20826 2808 20858
rect 2848 20826 2880 20858
rect 2920 20826 2952 20858
rect 2992 20826 3024 20858
rect 3064 20826 3096 20858
rect 3136 20826 3168 20858
rect 3208 20826 3240 20858
rect 3280 20826 3312 20858
rect 3352 20826 3384 20858
rect 3424 20826 3456 20858
rect 3496 20826 3528 20858
rect 3568 20826 3600 20858
rect 3640 20826 3672 20858
rect 3712 20826 3744 20858
rect 3784 20826 3816 20858
rect 3856 20826 3888 20858
rect 112 20754 144 20786
rect 184 20754 216 20786
rect 256 20754 288 20786
rect 328 20754 360 20786
rect 400 20754 432 20786
rect 472 20754 504 20786
rect 544 20754 576 20786
rect 616 20754 648 20786
rect 688 20754 720 20786
rect 760 20754 792 20786
rect 832 20754 864 20786
rect 904 20754 936 20786
rect 976 20754 1008 20786
rect 1048 20754 1080 20786
rect 1120 20754 1152 20786
rect 1192 20754 1224 20786
rect 1264 20754 1296 20786
rect 1336 20754 1368 20786
rect 1408 20754 1440 20786
rect 1480 20754 1512 20786
rect 1552 20754 1584 20786
rect 1624 20754 1656 20786
rect 1696 20754 1728 20786
rect 1768 20754 1800 20786
rect 1840 20754 1872 20786
rect 1912 20754 1944 20786
rect 1984 20754 2016 20786
rect 2056 20754 2088 20786
rect 2128 20754 2160 20786
rect 2200 20754 2232 20786
rect 2272 20754 2304 20786
rect 2344 20754 2376 20786
rect 2416 20754 2448 20786
rect 2488 20754 2520 20786
rect 2560 20754 2592 20786
rect 2632 20754 2664 20786
rect 2704 20754 2736 20786
rect 2776 20754 2808 20786
rect 2848 20754 2880 20786
rect 2920 20754 2952 20786
rect 2992 20754 3024 20786
rect 3064 20754 3096 20786
rect 3136 20754 3168 20786
rect 3208 20754 3240 20786
rect 3280 20754 3312 20786
rect 3352 20754 3384 20786
rect 3424 20754 3456 20786
rect 3496 20754 3528 20786
rect 3568 20754 3600 20786
rect 3640 20754 3672 20786
rect 3712 20754 3744 20786
rect 3784 20754 3816 20786
rect 3856 20754 3888 20786
rect 112 20682 144 20714
rect 184 20682 216 20714
rect 256 20682 288 20714
rect 328 20682 360 20714
rect 400 20682 432 20714
rect 472 20682 504 20714
rect 544 20682 576 20714
rect 616 20682 648 20714
rect 688 20682 720 20714
rect 760 20682 792 20714
rect 832 20682 864 20714
rect 904 20682 936 20714
rect 976 20682 1008 20714
rect 1048 20682 1080 20714
rect 1120 20682 1152 20714
rect 1192 20682 1224 20714
rect 1264 20682 1296 20714
rect 1336 20682 1368 20714
rect 1408 20682 1440 20714
rect 1480 20682 1512 20714
rect 1552 20682 1584 20714
rect 1624 20682 1656 20714
rect 1696 20682 1728 20714
rect 1768 20682 1800 20714
rect 1840 20682 1872 20714
rect 1912 20682 1944 20714
rect 1984 20682 2016 20714
rect 2056 20682 2088 20714
rect 2128 20682 2160 20714
rect 2200 20682 2232 20714
rect 2272 20682 2304 20714
rect 2344 20682 2376 20714
rect 2416 20682 2448 20714
rect 2488 20682 2520 20714
rect 2560 20682 2592 20714
rect 2632 20682 2664 20714
rect 2704 20682 2736 20714
rect 2776 20682 2808 20714
rect 2848 20682 2880 20714
rect 2920 20682 2952 20714
rect 2992 20682 3024 20714
rect 3064 20682 3096 20714
rect 3136 20682 3168 20714
rect 3208 20682 3240 20714
rect 3280 20682 3312 20714
rect 3352 20682 3384 20714
rect 3424 20682 3456 20714
rect 3496 20682 3528 20714
rect 3568 20682 3600 20714
rect 3640 20682 3672 20714
rect 3712 20682 3744 20714
rect 3784 20682 3816 20714
rect 3856 20682 3888 20714
rect 112 20610 144 20642
rect 184 20610 216 20642
rect 256 20610 288 20642
rect 328 20610 360 20642
rect 400 20610 432 20642
rect 472 20610 504 20642
rect 544 20610 576 20642
rect 616 20610 648 20642
rect 688 20610 720 20642
rect 760 20610 792 20642
rect 832 20610 864 20642
rect 904 20610 936 20642
rect 976 20610 1008 20642
rect 1048 20610 1080 20642
rect 1120 20610 1152 20642
rect 1192 20610 1224 20642
rect 1264 20610 1296 20642
rect 1336 20610 1368 20642
rect 1408 20610 1440 20642
rect 1480 20610 1512 20642
rect 1552 20610 1584 20642
rect 1624 20610 1656 20642
rect 1696 20610 1728 20642
rect 1768 20610 1800 20642
rect 1840 20610 1872 20642
rect 1912 20610 1944 20642
rect 1984 20610 2016 20642
rect 2056 20610 2088 20642
rect 2128 20610 2160 20642
rect 2200 20610 2232 20642
rect 2272 20610 2304 20642
rect 2344 20610 2376 20642
rect 2416 20610 2448 20642
rect 2488 20610 2520 20642
rect 2560 20610 2592 20642
rect 2632 20610 2664 20642
rect 2704 20610 2736 20642
rect 2776 20610 2808 20642
rect 2848 20610 2880 20642
rect 2920 20610 2952 20642
rect 2992 20610 3024 20642
rect 3064 20610 3096 20642
rect 3136 20610 3168 20642
rect 3208 20610 3240 20642
rect 3280 20610 3312 20642
rect 3352 20610 3384 20642
rect 3424 20610 3456 20642
rect 3496 20610 3528 20642
rect 3568 20610 3600 20642
rect 3640 20610 3672 20642
rect 3712 20610 3744 20642
rect 3784 20610 3816 20642
rect 3856 20610 3888 20642
rect 112 20538 144 20570
rect 184 20538 216 20570
rect 256 20538 288 20570
rect 328 20538 360 20570
rect 400 20538 432 20570
rect 472 20538 504 20570
rect 544 20538 576 20570
rect 616 20538 648 20570
rect 688 20538 720 20570
rect 760 20538 792 20570
rect 832 20538 864 20570
rect 904 20538 936 20570
rect 976 20538 1008 20570
rect 1048 20538 1080 20570
rect 1120 20538 1152 20570
rect 1192 20538 1224 20570
rect 1264 20538 1296 20570
rect 1336 20538 1368 20570
rect 1408 20538 1440 20570
rect 1480 20538 1512 20570
rect 1552 20538 1584 20570
rect 1624 20538 1656 20570
rect 1696 20538 1728 20570
rect 1768 20538 1800 20570
rect 1840 20538 1872 20570
rect 1912 20538 1944 20570
rect 1984 20538 2016 20570
rect 2056 20538 2088 20570
rect 2128 20538 2160 20570
rect 2200 20538 2232 20570
rect 2272 20538 2304 20570
rect 2344 20538 2376 20570
rect 2416 20538 2448 20570
rect 2488 20538 2520 20570
rect 2560 20538 2592 20570
rect 2632 20538 2664 20570
rect 2704 20538 2736 20570
rect 2776 20538 2808 20570
rect 2848 20538 2880 20570
rect 2920 20538 2952 20570
rect 2992 20538 3024 20570
rect 3064 20538 3096 20570
rect 3136 20538 3168 20570
rect 3208 20538 3240 20570
rect 3280 20538 3312 20570
rect 3352 20538 3384 20570
rect 3424 20538 3456 20570
rect 3496 20538 3528 20570
rect 3568 20538 3600 20570
rect 3640 20538 3672 20570
rect 3712 20538 3744 20570
rect 3784 20538 3816 20570
rect 3856 20538 3888 20570
rect 112 20466 144 20498
rect 184 20466 216 20498
rect 256 20466 288 20498
rect 328 20466 360 20498
rect 400 20466 432 20498
rect 472 20466 504 20498
rect 544 20466 576 20498
rect 616 20466 648 20498
rect 688 20466 720 20498
rect 760 20466 792 20498
rect 832 20466 864 20498
rect 904 20466 936 20498
rect 976 20466 1008 20498
rect 1048 20466 1080 20498
rect 1120 20466 1152 20498
rect 1192 20466 1224 20498
rect 1264 20466 1296 20498
rect 1336 20466 1368 20498
rect 1408 20466 1440 20498
rect 1480 20466 1512 20498
rect 1552 20466 1584 20498
rect 1624 20466 1656 20498
rect 1696 20466 1728 20498
rect 1768 20466 1800 20498
rect 1840 20466 1872 20498
rect 1912 20466 1944 20498
rect 1984 20466 2016 20498
rect 2056 20466 2088 20498
rect 2128 20466 2160 20498
rect 2200 20466 2232 20498
rect 2272 20466 2304 20498
rect 2344 20466 2376 20498
rect 2416 20466 2448 20498
rect 2488 20466 2520 20498
rect 2560 20466 2592 20498
rect 2632 20466 2664 20498
rect 2704 20466 2736 20498
rect 2776 20466 2808 20498
rect 2848 20466 2880 20498
rect 2920 20466 2952 20498
rect 2992 20466 3024 20498
rect 3064 20466 3096 20498
rect 3136 20466 3168 20498
rect 3208 20466 3240 20498
rect 3280 20466 3312 20498
rect 3352 20466 3384 20498
rect 3424 20466 3456 20498
rect 3496 20466 3528 20498
rect 3568 20466 3600 20498
rect 3640 20466 3672 20498
rect 3712 20466 3744 20498
rect 3784 20466 3816 20498
rect 3856 20466 3888 20498
rect 112 20394 144 20426
rect 184 20394 216 20426
rect 256 20394 288 20426
rect 328 20394 360 20426
rect 400 20394 432 20426
rect 472 20394 504 20426
rect 544 20394 576 20426
rect 616 20394 648 20426
rect 688 20394 720 20426
rect 760 20394 792 20426
rect 832 20394 864 20426
rect 904 20394 936 20426
rect 976 20394 1008 20426
rect 1048 20394 1080 20426
rect 1120 20394 1152 20426
rect 1192 20394 1224 20426
rect 1264 20394 1296 20426
rect 1336 20394 1368 20426
rect 1408 20394 1440 20426
rect 1480 20394 1512 20426
rect 1552 20394 1584 20426
rect 1624 20394 1656 20426
rect 1696 20394 1728 20426
rect 1768 20394 1800 20426
rect 1840 20394 1872 20426
rect 1912 20394 1944 20426
rect 1984 20394 2016 20426
rect 2056 20394 2088 20426
rect 2128 20394 2160 20426
rect 2200 20394 2232 20426
rect 2272 20394 2304 20426
rect 2344 20394 2376 20426
rect 2416 20394 2448 20426
rect 2488 20394 2520 20426
rect 2560 20394 2592 20426
rect 2632 20394 2664 20426
rect 2704 20394 2736 20426
rect 2776 20394 2808 20426
rect 2848 20394 2880 20426
rect 2920 20394 2952 20426
rect 2992 20394 3024 20426
rect 3064 20394 3096 20426
rect 3136 20394 3168 20426
rect 3208 20394 3240 20426
rect 3280 20394 3312 20426
rect 3352 20394 3384 20426
rect 3424 20394 3456 20426
rect 3496 20394 3528 20426
rect 3568 20394 3600 20426
rect 3640 20394 3672 20426
rect 3712 20394 3744 20426
rect 3784 20394 3816 20426
rect 3856 20394 3888 20426
rect 112 20322 144 20354
rect 184 20322 216 20354
rect 256 20322 288 20354
rect 328 20322 360 20354
rect 400 20322 432 20354
rect 472 20322 504 20354
rect 544 20322 576 20354
rect 616 20322 648 20354
rect 688 20322 720 20354
rect 760 20322 792 20354
rect 832 20322 864 20354
rect 904 20322 936 20354
rect 976 20322 1008 20354
rect 1048 20322 1080 20354
rect 1120 20322 1152 20354
rect 1192 20322 1224 20354
rect 1264 20322 1296 20354
rect 1336 20322 1368 20354
rect 1408 20322 1440 20354
rect 1480 20322 1512 20354
rect 1552 20322 1584 20354
rect 1624 20322 1656 20354
rect 1696 20322 1728 20354
rect 1768 20322 1800 20354
rect 1840 20322 1872 20354
rect 1912 20322 1944 20354
rect 1984 20322 2016 20354
rect 2056 20322 2088 20354
rect 2128 20322 2160 20354
rect 2200 20322 2232 20354
rect 2272 20322 2304 20354
rect 2344 20322 2376 20354
rect 2416 20322 2448 20354
rect 2488 20322 2520 20354
rect 2560 20322 2592 20354
rect 2632 20322 2664 20354
rect 2704 20322 2736 20354
rect 2776 20322 2808 20354
rect 2848 20322 2880 20354
rect 2920 20322 2952 20354
rect 2992 20322 3024 20354
rect 3064 20322 3096 20354
rect 3136 20322 3168 20354
rect 3208 20322 3240 20354
rect 3280 20322 3312 20354
rect 3352 20322 3384 20354
rect 3424 20322 3456 20354
rect 3496 20322 3528 20354
rect 3568 20322 3600 20354
rect 3640 20322 3672 20354
rect 3712 20322 3744 20354
rect 3784 20322 3816 20354
rect 3856 20322 3888 20354
rect 112 20250 144 20282
rect 184 20250 216 20282
rect 256 20250 288 20282
rect 328 20250 360 20282
rect 400 20250 432 20282
rect 472 20250 504 20282
rect 544 20250 576 20282
rect 616 20250 648 20282
rect 688 20250 720 20282
rect 760 20250 792 20282
rect 832 20250 864 20282
rect 904 20250 936 20282
rect 976 20250 1008 20282
rect 1048 20250 1080 20282
rect 1120 20250 1152 20282
rect 1192 20250 1224 20282
rect 1264 20250 1296 20282
rect 1336 20250 1368 20282
rect 1408 20250 1440 20282
rect 1480 20250 1512 20282
rect 1552 20250 1584 20282
rect 1624 20250 1656 20282
rect 1696 20250 1728 20282
rect 1768 20250 1800 20282
rect 1840 20250 1872 20282
rect 1912 20250 1944 20282
rect 1984 20250 2016 20282
rect 2056 20250 2088 20282
rect 2128 20250 2160 20282
rect 2200 20250 2232 20282
rect 2272 20250 2304 20282
rect 2344 20250 2376 20282
rect 2416 20250 2448 20282
rect 2488 20250 2520 20282
rect 2560 20250 2592 20282
rect 2632 20250 2664 20282
rect 2704 20250 2736 20282
rect 2776 20250 2808 20282
rect 2848 20250 2880 20282
rect 2920 20250 2952 20282
rect 2992 20250 3024 20282
rect 3064 20250 3096 20282
rect 3136 20250 3168 20282
rect 3208 20250 3240 20282
rect 3280 20250 3312 20282
rect 3352 20250 3384 20282
rect 3424 20250 3456 20282
rect 3496 20250 3528 20282
rect 3568 20250 3600 20282
rect 3640 20250 3672 20282
rect 3712 20250 3744 20282
rect 3784 20250 3816 20282
rect 3856 20250 3888 20282
rect 112 20178 144 20210
rect 184 20178 216 20210
rect 256 20178 288 20210
rect 328 20178 360 20210
rect 400 20178 432 20210
rect 472 20178 504 20210
rect 544 20178 576 20210
rect 616 20178 648 20210
rect 688 20178 720 20210
rect 760 20178 792 20210
rect 832 20178 864 20210
rect 904 20178 936 20210
rect 976 20178 1008 20210
rect 1048 20178 1080 20210
rect 1120 20178 1152 20210
rect 1192 20178 1224 20210
rect 1264 20178 1296 20210
rect 1336 20178 1368 20210
rect 1408 20178 1440 20210
rect 1480 20178 1512 20210
rect 1552 20178 1584 20210
rect 1624 20178 1656 20210
rect 1696 20178 1728 20210
rect 1768 20178 1800 20210
rect 1840 20178 1872 20210
rect 1912 20178 1944 20210
rect 1984 20178 2016 20210
rect 2056 20178 2088 20210
rect 2128 20178 2160 20210
rect 2200 20178 2232 20210
rect 2272 20178 2304 20210
rect 2344 20178 2376 20210
rect 2416 20178 2448 20210
rect 2488 20178 2520 20210
rect 2560 20178 2592 20210
rect 2632 20178 2664 20210
rect 2704 20178 2736 20210
rect 2776 20178 2808 20210
rect 2848 20178 2880 20210
rect 2920 20178 2952 20210
rect 2992 20178 3024 20210
rect 3064 20178 3096 20210
rect 3136 20178 3168 20210
rect 3208 20178 3240 20210
rect 3280 20178 3312 20210
rect 3352 20178 3384 20210
rect 3424 20178 3456 20210
rect 3496 20178 3528 20210
rect 3568 20178 3600 20210
rect 3640 20178 3672 20210
rect 3712 20178 3744 20210
rect 3784 20178 3816 20210
rect 3856 20178 3888 20210
rect 112 20106 144 20138
rect 184 20106 216 20138
rect 256 20106 288 20138
rect 328 20106 360 20138
rect 400 20106 432 20138
rect 472 20106 504 20138
rect 544 20106 576 20138
rect 616 20106 648 20138
rect 688 20106 720 20138
rect 760 20106 792 20138
rect 832 20106 864 20138
rect 904 20106 936 20138
rect 976 20106 1008 20138
rect 1048 20106 1080 20138
rect 1120 20106 1152 20138
rect 1192 20106 1224 20138
rect 1264 20106 1296 20138
rect 1336 20106 1368 20138
rect 1408 20106 1440 20138
rect 1480 20106 1512 20138
rect 1552 20106 1584 20138
rect 1624 20106 1656 20138
rect 1696 20106 1728 20138
rect 1768 20106 1800 20138
rect 1840 20106 1872 20138
rect 1912 20106 1944 20138
rect 1984 20106 2016 20138
rect 2056 20106 2088 20138
rect 2128 20106 2160 20138
rect 2200 20106 2232 20138
rect 2272 20106 2304 20138
rect 2344 20106 2376 20138
rect 2416 20106 2448 20138
rect 2488 20106 2520 20138
rect 2560 20106 2592 20138
rect 2632 20106 2664 20138
rect 2704 20106 2736 20138
rect 2776 20106 2808 20138
rect 2848 20106 2880 20138
rect 2920 20106 2952 20138
rect 2992 20106 3024 20138
rect 3064 20106 3096 20138
rect 3136 20106 3168 20138
rect 3208 20106 3240 20138
rect 3280 20106 3312 20138
rect 3352 20106 3384 20138
rect 3424 20106 3456 20138
rect 3496 20106 3528 20138
rect 3568 20106 3600 20138
rect 3640 20106 3672 20138
rect 3712 20106 3744 20138
rect 3784 20106 3816 20138
rect 3856 20106 3888 20138
rect 112 20034 144 20066
rect 184 20034 216 20066
rect 256 20034 288 20066
rect 328 20034 360 20066
rect 400 20034 432 20066
rect 472 20034 504 20066
rect 544 20034 576 20066
rect 616 20034 648 20066
rect 688 20034 720 20066
rect 760 20034 792 20066
rect 832 20034 864 20066
rect 904 20034 936 20066
rect 976 20034 1008 20066
rect 1048 20034 1080 20066
rect 1120 20034 1152 20066
rect 1192 20034 1224 20066
rect 1264 20034 1296 20066
rect 1336 20034 1368 20066
rect 1408 20034 1440 20066
rect 1480 20034 1512 20066
rect 1552 20034 1584 20066
rect 1624 20034 1656 20066
rect 1696 20034 1728 20066
rect 1768 20034 1800 20066
rect 1840 20034 1872 20066
rect 1912 20034 1944 20066
rect 1984 20034 2016 20066
rect 2056 20034 2088 20066
rect 2128 20034 2160 20066
rect 2200 20034 2232 20066
rect 2272 20034 2304 20066
rect 2344 20034 2376 20066
rect 2416 20034 2448 20066
rect 2488 20034 2520 20066
rect 2560 20034 2592 20066
rect 2632 20034 2664 20066
rect 2704 20034 2736 20066
rect 2776 20034 2808 20066
rect 2848 20034 2880 20066
rect 2920 20034 2952 20066
rect 2992 20034 3024 20066
rect 3064 20034 3096 20066
rect 3136 20034 3168 20066
rect 3208 20034 3240 20066
rect 3280 20034 3312 20066
rect 3352 20034 3384 20066
rect 3424 20034 3456 20066
rect 3496 20034 3528 20066
rect 3568 20034 3600 20066
rect 3640 20034 3672 20066
rect 3712 20034 3744 20066
rect 3784 20034 3816 20066
rect 3856 20034 3888 20066
rect 112 19962 144 19994
rect 184 19962 216 19994
rect 256 19962 288 19994
rect 328 19962 360 19994
rect 400 19962 432 19994
rect 472 19962 504 19994
rect 544 19962 576 19994
rect 616 19962 648 19994
rect 688 19962 720 19994
rect 760 19962 792 19994
rect 832 19962 864 19994
rect 904 19962 936 19994
rect 976 19962 1008 19994
rect 1048 19962 1080 19994
rect 1120 19962 1152 19994
rect 1192 19962 1224 19994
rect 1264 19962 1296 19994
rect 1336 19962 1368 19994
rect 1408 19962 1440 19994
rect 1480 19962 1512 19994
rect 1552 19962 1584 19994
rect 1624 19962 1656 19994
rect 1696 19962 1728 19994
rect 1768 19962 1800 19994
rect 1840 19962 1872 19994
rect 1912 19962 1944 19994
rect 1984 19962 2016 19994
rect 2056 19962 2088 19994
rect 2128 19962 2160 19994
rect 2200 19962 2232 19994
rect 2272 19962 2304 19994
rect 2344 19962 2376 19994
rect 2416 19962 2448 19994
rect 2488 19962 2520 19994
rect 2560 19962 2592 19994
rect 2632 19962 2664 19994
rect 2704 19962 2736 19994
rect 2776 19962 2808 19994
rect 2848 19962 2880 19994
rect 2920 19962 2952 19994
rect 2992 19962 3024 19994
rect 3064 19962 3096 19994
rect 3136 19962 3168 19994
rect 3208 19962 3240 19994
rect 3280 19962 3312 19994
rect 3352 19962 3384 19994
rect 3424 19962 3456 19994
rect 3496 19962 3528 19994
rect 3568 19962 3600 19994
rect 3640 19962 3672 19994
rect 3712 19962 3744 19994
rect 3784 19962 3816 19994
rect 3856 19962 3888 19994
rect 112 19890 144 19922
rect 184 19890 216 19922
rect 256 19890 288 19922
rect 328 19890 360 19922
rect 400 19890 432 19922
rect 472 19890 504 19922
rect 544 19890 576 19922
rect 616 19890 648 19922
rect 688 19890 720 19922
rect 760 19890 792 19922
rect 832 19890 864 19922
rect 904 19890 936 19922
rect 976 19890 1008 19922
rect 1048 19890 1080 19922
rect 1120 19890 1152 19922
rect 1192 19890 1224 19922
rect 1264 19890 1296 19922
rect 1336 19890 1368 19922
rect 1408 19890 1440 19922
rect 1480 19890 1512 19922
rect 1552 19890 1584 19922
rect 1624 19890 1656 19922
rect 1696 19890 1728 19922
rect 1768 19890 1800 19922
rect 1840 19890 1872 19922
rect 1912 19890 1944 19922
rect 1984 19890 2016 19922
rect 2056 19890 2088 19922
rect 2128 19890 2160 19922
rect 2200 19890 2232 19922
rect 2272 19890 2304 19922
rect 2344 19890 2376 19922
rect 2416 19890 2448 19922
rect 2488 19890 2520 19922
rect 2560 19890 2592 19922
rect 2632 19890 2664 19922
rect 2704 19890 2736 19922
rect 2776 19890 2808 19922
rect 2848 19890 2880 19922
rect 2920 19890 2952 19922
rect 2992 19890 3024 19922
rect 3064 19890 3096 19922
rect 3136 19890 3168 19922
rect 3208 19890 3240 19922
rect 3280 19890 3312 19922
rect 3352 19890 3384 19922
rect 3424 19890 3456 19922
rect 3496 19890 3528 19922
rect 3568 19890 3600 19922
rect 3640 19890 3672 19922
rect 3712 19890 3744 19922
rect 3784 19890 3816 19922
rect 3856 19890 3888 19922
rect 112 19818 144 19850
rect 184 19818 216 19850
rect 256 19818 288 19850
rect 328 19818 360 19850
rect 400 19818 432 19850
rect 472 19818 504 19850
rect 544 19818 576 19850
rect 616 19818 648 19850
rect 688 19818 720 19850
rect 760 19818 792 19850
rect 832 19818 864 19850
rect 904 19818 936 19850
rect 976 19818 1008 19850
rect 1048 19818 1080 19850
rect 1120 19818 1152 19850
rect 1192 19818 1224 19850
rect 1264 19818 1296 19850
rect 1336 19818 1368 19850
rect 1408 19818 1440 19850
rect 1480 19818 1512 19850
rect 1552 19818 1584 19850
rect 1624 19818 1656 19850
rect 1696 19818 1728 19850
rect 1768 19818 1800 19850
rect 1840 19818 1872 19850
rect 1912 19818 1944 19850
rect 1984 19818 2016 19850
rect 2056 19818 2088 19850
rect 2128 19818 2160 19850
rect 2200 19818 2232 19850
rect 2272 19818 2304 19850
rect 2344 19818 2376 19850
rect 2416 19818 2448 19850
rect 2488 19818 2520 19850
rect 2560 19818 2592 19850
rect 2632 19818 2664 19850
rect 2704 19818 2736 19850
rect 2776 19818 2808 19850
rect 2848 19818 2880 19850
rect 2920 19818 2952 19850
rect 2992 19818 3024 19850
rect 3064 19818 3096 19850
rect 3136 19818 3168 19850
rect 3208 19818 3240 19850
rect 3280 19818 3312 19850
rect 3352 19818 3384 19850
rect 3424 19818 3456 19850
rect 3496 19818 3528 19850
rect 3568 19818 3600 19850
rect 3640 19818 3672 19850
rect 3712 19818 3744 19850
rect 3784 19818 3816 19850
rect 3856 19818 3888 19850
rect 112 19746 144 19778
rect 184 19746 216 19778
rect 256 19746 288 19778
rect 328 19746 360 19778
rect 400 19746 432 19778
rect 472 19746 504 19778
rect 544 19746 576 19778
rect 616 19746 648 19778
rect 688 19746 720 19778
rect 760 19746 792 19778
rect 832 19746 864 19778
rect 904 19746 936 19778
rect 976 19746 1008 19778
rect 1048 19746 1080 19778
rect 1120 19746 1152 19778
rect 1192 19746 1224 19778
rect 1264 19746 1296 19778
rect 1336 19746 1368 19778
rect 1408 19746 1440 19778
rect 1480 19746 1512 19778
rect 1552 19746 1584 19778
rect 1624 19746 1656 19778
rect 1696 19746 1728 19778
rect 1768 19746 1800 19778
rect 1840 19746 1872 19778
rect 1912 19746 1944 19778
rect 1984 19746 2016 19778
rect 2056 19746 2088 19778
rect 2128 19746 2160 19778
rect 2200 19746 2232 19778
rect 2272 19746 2304 19778
rect 2344 19746 2376 19778
rect 2416 19746 2448 19778
rect 2488 19746 2520 19778
rect 2560 19746 2592 19778
rect 2632 19746 2664 19778
rect 2704 19746 2736 19778
rect 2776 19746 2808 19778
rect 2848 19746 2880 19778
rect 2920 19746 2952 19778
rect 2992 19746 3024 19778
rect 3064 19746 3096 19778
rect 3136 19746 3168 19778
rect 3208 19746 3240 19778
rect 3280 19746 3312 19778
rect 3352 19746 3384 19778
rect 3424 19746 3456 19778
rect 3496 19746 3528 19778
rect 3568 19746 3600 19778
rect 3640 19746 3672 19778
rect 3712 19746 3744 19778
rect 3784 19746 3816 19778
rect 3856 19746 3888 19778
rect 112 19674 144 19706
rect 184 19674 216 19706
rect 256 19674 288 19706
rect 328 19674 360 19706
rect 400 19674 432 19706
rect 472 19674 504 19706
rect 544 19674 576 19706
rect 616 19674 648 19706
rect 688 19674 720 19706
rect 760 19674 792 19706
rect 832 19674 864 19706
rect 904 19674 936 19706
rect 976 19674 1008 19706
rect 1048 19674 1080 19706
rect 1120 19674 1152 19706
rect 1192 19674 1224 19706
rect 1264 19674 1296 19706
rect 1336 19674 1368 19706
rect 1408 19674 1440 19706
rect 1480 19674 1512 19706
rect 1552 19674 1584 19706
rect 1624 19674 1656 19706
rect 1696 19674 1728 19706
rect 1768 19674 1800 19706
rect 1840 19674 1872 19706
rect 1912 19674 1944 19706
rect 1984 19674 2016 19706
rect 2056 19674 2088 19706
rect 2128 19674 2160 19706
rect 2200 19674 2232 19706
rect 2272 19674 2304 19706
rect 2344 19674 2376 19706
rect 2416 19674 2448 19706
rect 2488 19674 2520 19706
rect 2560 19674 2592 19706
rect 2632 19674 2664 19706
rect 2704 19674 2736 19706
rect 2776 19674 2808 19706
rect 2848 19674 2880 19706
rect 2920 19674 2952 19706
rect 2992 19674 3024 19706
rect 3064 19674 3096 19706
rect 3136 19674 3168 19706
rect 3208 19674 3240 19706
rect 3280 19674 3312 19706
rect 3352 19674 3384 19706
rect 3424 19674 3456 19706
rect 3496 19674 3528 19706
rect 3568 19674 3600 19706
rect 3640 19674 3672 19706
rect 3712 19674 3744 19706
rect 3784 19674 3816 19706
rect 3856 19674 3888 19706
rect 112 19602 144 19634
rect 184 19602 216 19634
rect 256 19602 288 19634
rect 328 19602 360 19634
rect 400 19602 432 19634
rect 472 19602 504 19634
rect 544 19602 576 19634
rect 616 19602 648 19634
rect 688 19602 720 19634
rect 760 19602 792 19634
rect 832 19602 864 19634
rect 904 19602 936 19634
rect 976 19602 1008 19634
rect 1048 19602 1080 19634
rect 1120 19602 1152 19634
rect 1192 19602 1224 19634
rect 1264 19602 1296 19634
rect 1336 19602 1368 19634
rect 1408 19602 1440 19634
rect 1480 19602 1512 19634
rect 1552 19602 1584 19634
rect 1624 19602 1656 19634
rect 1696 19602 1728 19634
rect 1768 19602 1800 19634
rect 1840 19602 1872 19634
rect 1912 19602 1944 19634
rect 1984 19602 2016 19634
rect 2056 19602 2088 19634
rect 2128 19602 2160 19634
rect 2200 19602 2232 19634
rect 2272 19602 2304 19634
rect 2344 19602 2376 19634
rect 2416 19602 2448 19634
rect 2488 19602 2520 19634
rect 2560 19602 2592 19634
rect 2632 19602 2664 19634
rect 2704 19602 2736 19634
rect 2776 19602 2808 19634
rect 2848 19602 2880 19634
rect 2920 19602 2952 19634
rect 2992 19602 3024 19634
rect 3064 19602 3096 19634
rect 3136 19602 3168 19634
rect 3208 19602 3240 19634
rect 3280 19602 3312 19634
rect 3352 19602 3384 19634
rect 3424 19602 3456 19634
rect 3496 19602 3528 19634
rect 3568 19602 3600 19634
rect 3640 19602 3672 19634
rect 3712 19602 3744 19634
rect 3784 19602 3816 19634
rect 3856 19602 3888 19634
rect 112 19530 144 19562
rect 184 19530 216 19562
rect 256 19530 288 19562
rect 328 19530 360 19562
rect 400 19530 432 19562
rect 472 19530 504 19562
rect 544 19530 576 19562
rect 616 19530 648 19562
rect 688 19530 720 19562
rect 760 19530 792 19562
rect 832 19530 864 19562
rect 904 19530 936 19562
rect 976 19530 1008 19562
rect 1048 19530 1080 19562
rect 1120 19530 1152 19562
rect 1192 19530 1224 19562
rect 1264 19530 1296 19562
rect 1336 19530 1368 19562
rect 1408 19530 1440 19562
rect 1480 19530 1512 19562
rect 1552 19530 1584 19562
rect 1624 19530 1656 19562
rect 1696 19530 1728 19562
rect 1768 19530 1800 19562
rect 1840 19530 1872 19562
rect 1912 19530 1944 19562
rect 1984 19530 2016 19562
rect 2056 19530 2088 19562
rect 2128 19530 2160 19562
rect 2200 19530 2232 19562
rect 2272 19530 2304 19562
rect 2344 19530 2376 19562
rect 2416 19530 2448 19562
rect 2488 19530 2520 19562
rect 2560 19530 2592 19562
rect 2632 19530 2664 19562
rect 2704 19530 2736 19562
rect 2776 19530 2808 19562
rect 2848 19530 2880 19562
rect 2920 19530 2952 19562
rect 2992 19530 3024 19562
rect 3064 19530 3096 19562
rect 3136 19530 3168 19562
rect 3208 19530 3240 19562
rect 3280 19530 3312 19562
rect 3352 19530 3384 19562
rect 3424 19530 3456 19562
rect 3496 19530 3528 19562
rect 3568 19530 3600 19562
rect 3640 19530 3672 19562
rect 3712 19530 3744 19562
rect 3784 19530 3816 19562
rect 3856 19530 3888 19562
rect 112 19458 144 19490
rect 184 19458 216 19490
rect 256 19458 288 19490
rect 328 19458 360 19490
rect 400 19458 432 19490
rect 472 19458 504 19490
rect 544 19458 576 19490
rect 616 19458 648 19490
rect 688 19458 720 19490
rect 760 19458 792 19490
rect 832 19458 864 19490
rect 904 19458 936 19490
rect 976 19458 1008 19490
rect 1048 19458 1080 19490
rect 1120 19458 1152 19490
rect 1192 19458 1224 19490
rect 1264 19458 1296 19490
rect 1336 19458 1368 19490
rect 1408 19458 1440 19490
rect 1480 19458 1512 19490
rect 1552 19458 1584 19490
rect 1624 19458 1656 19490
rect 1696 19458 1728 19490
rect 1768 19458 1800 19490
rect 1840 19458 1872 19490
rect 1912 19458 1944 19490
rect 1984 19458 2016 19490
rect 2056 19458 2088 19490
rect 2128 19458 2160 19490
rect 2200 19458 2232 19490
rect 2272 19458 2304 19490
rect 2344 19458 2376 19490
rect 2416 19458 2448 19490
rect 2488 19458 2520 19490
rect 2560 19458 2592 19490
rect 2632 19458 2664 19490
rect 2704 19458 2736 19490
rect 2776 19458 2808 19490
rect 2848 19458 2880 19490
rect 2920 19458 2952 19490
rect 2992 19458 3024 19490
rect 3064 19458 3096 19490
rect 3136 19458 3168 19490
rect 3208 19458 3240 19490
rect 3280 19458 3312 19490
rect 3352 19458 3384 19490
rect 3424 19458 3456 19490
rect 3496 19458 3528 19490
rect 3568 19458 3600 19490
rect 3640 19458 3672 19490
rect 3712 19458 3744 19490
rect 3784 19458 3816 19490
rect 3856 19458 3888 19490
rect 112 19386 144 19418
rect 184 19386 216 19418
rect 256 19386 288 19418
rect 328 19386 360 19418
rect 400 19386 432 19418
rect 472 19386 504 19418
rect 544 19386 576 19418
rect 616 19386 648 19418
rect 688 19386 720 19418
rect 760 19386 792 19418
rect 832 19386 864 19418
rect 904 19386 936 19418
rect 976 19386 1008 19418
rect 1048 19386 1080 19418
rect 1120 19386 1152 19418
rect 1192 19386 1224 19418
rect 1264 19386 1296 19418
rect 1336 19386 1368 19418
rect 1408 19386 1440 19418
rect 1480 19386 1512 19418
rect 1552 19386 1584 19418
rect 1624 19386 1656 19418
rect 1696 19386 1728 19418
rect 1768 19386 1800 19418
rect 1840 19386 1872 19418
rect 1912 19386 1944 19418
rect 1984 19386 2016 19418
rect 2056 19386 2088 19418
rect 2128 19386 2160 19418
rect 2200 19386 2232 19418
rect 2272 19386 2304 19418
rect 2344 19386 2376 19418
rect 2416 19386 2448 19418
rect 2488 19386 2520 19418
rect 2560 19386 2592 19418
rect 2632 19386 2664 19418
rect 2704 19386 2736 19418
rect 2776 19386 2808 19418
rect 2848 19386 2880 19418
rect 2920 19386 2952 19418
rect 2992 19386 3024 19418
rect 3064 19386 3096 19418
rect 3136 19386 3168 19418
rect 3208 19386 3240 19418
rect 3280 19386 3312 19418
rect 3352 19386 3384 19418
rect 3424 19386 3456 19418
rect 3496 19386 3528 19418
rect 3568 19386 3600 19418
rect 3640 19386 3672 19418
rect 3712 19386 3744 19418
rect 3784 19386 3816 19418
rect 3856 19386 3888 19418
rect 112 19314 144 19346
rect 184 19314 216 19346
rect 256 19314 288 19346
rect 328 19314 360 19346
rect 400 19314 432 19346
rect 472 19314 504 19346
rect 544 19314 576 19346
rect 616 19314 648 19346
rect 688 19314 720 19346
rect 760 19314 792 19346
rect 832 19314 864 19346
rect 904 19314 936 19346
rect 976 19314 1008 19346
rect 1048 19314 1080 19346
rect 1120 19314 1152 19346
rect 1192 19314 1224 19346
rect 1264 19314 1296 19346
rect 1336 19314 1368 19346
rect 1408 19314 1440 19346
rect 1480 19314 1512 19346
rect 1552 19314 1584 19346
rect 1624 19314 1656 19346
rect 1696 19314 1728 19346
rect 1768 19314 1800 19346
rect 1840 19314 1872 19346
rect 1912 19314 1944 19346
rect 1984 19314 2016 19346
rect 2056 19314 2088 19346
rect 2128 19314 2160 19346
rect 2200 19314 2232 19346
rect 2272 19314 2304 19346
rect 2344 19314 2376 19346
rect 2416 19314 2448 19346
rect 2488 19314 2520 19346
rect 2560 19314 2592 19346
rect 2632 19314 2664 19346
rect 2704 19314 2736 19346
rect 2776 19314 2808 19346
rect 2848 19314 2880 19346
rect 2920 19314 2952 19346
rect 2992 19314 3024 19346
rect 3064 19314 3096 19346
rect 3136 19314 3168 19346
rect 3208 19314 3240 19346
rect 3280 19314 3312 19346
rect 3352 19314 3384 19346
rect 3424 19314 3456 19346
rect 3496 19314 3528 19346
rect 3568 19314 3600 19346
rect 3640 19314 3672 19346
rect 3712 19314 3744 19346
rect 3784 19314 3816 19346
rect 3856 19314 3888 19346
rect 112 19242 144 19274
rect 184 19242 216 19274
rect 256 19242 288 19274
rect 328 19242 360 19274
rect 400 19242 432 19274
rect 472 19242 504 19274
rect 544 19242 576 19274
rect 616 19242 648 19274
rect 688 19242 720 19274
rect 760 19242 792 19274
rect 832 19242 864 19274
rect 904 19242 936 19274
rect 976 19242 1008 19274
rect 1048 19242 1080 19274
rect 1120 19242 1152 19274
rect 1192 19242 1224 19274
rect 1264 19242 1296 19274
rect 1336 19242 1368 19274
rect 1408 19242 1440 19274
rect 1480 19242 1512 19274
rect 1552 19242 1584 19274
rect 1624 19242 1656 19274
rect 1696 19242 1728 19274
rect 1768 19242 1800 19274
rect 1840 19242 1872 19274
rect 1912 19242 1944 19274
rect 1984 19242 2016 19274
rect 2056 19242 2088 19274
rect 2128 19242 2160 19274
rect 2200 19242 2232 19274
rect 2272 19242 2304 19274
rect 2344 19242 2376 19274
rect 2416 19242 2448 19274
rect 2488 19242 2520 19274
rect 2560 19242 2592 19274
rect 2632 19242 2664 19274
rect 2704 19242 2736 19274
rect 2776 19242 2808 19274
rect 2848 19242 2880 19274
rect 2920 19242 2952 19274
rect 2992 19242 3024 19274
rect 3064 19242 3096 19274
rect 3136 19242 3168 19274
rect 3208 19242 3240 19274
rect 3280 19242 3312 19274
rect 3352 19242 3384 19274
rect 3424 19242 3456 19274
rect 3496 19242 3528 19274
rect 3568 19242 3600 19274
rect 3640 19242 3672 19274
rect 3712 19242 3744 19274
rect 3784 19242 3816 19274
rect 3856 19242 3888 19274
rect 112 19170 144 19202
rect 184 19170 216 19202
rect 256 19170 288 19202
rect 328 19170 360 19202
rect 400 19170 432 19202
rect 472 19170 504 19202
rect 544 19170 576 19202
rect 616 19170 648 19202
rect 688 19170 720 19202
rect 760 19170 792 19202
rect 832 19170 864 19202
rect 904 19170 936 19202
rect 976 19170 1008 19202
rect 1048 19170 1080 19202
rect 1120 19170 1152 19202
rect 1192 19170 1224 19202
rect 1264 19170 1296 19202
rect 1336 19170 1368 19202
rect 1408 19170 1440 19202
rect 1480 19170 1512 19202
rect 1552 19170 1584 19202
rect 1624 19170 1656 19202
rect 1696 19170 1728 19202
rect 1768 19170 1800 19202
rect 1840 19170 1872 19202
rect 1912 19170 1944 19202
rect 1984 19170 2016 19202
rect 2056 19170 2088 19202
rect 2128 19170 2160 19202
rect 2200 19170 2232 19202
rect 2272 19170 2304 19202
rect 2344 19170 2376 19202
rect 2416 19170 2448 19202
rect 2488 19170 2520 19202
rect 2560 19170 2592 19202
rect 2632 19170 2664 19202
rect 2704 19170 2736 19202
rect 2776 19170 2808 19202
rect 2848 19170 2880 19202
rect 2920 19170 2952 19202
rect 2992 19170 3024 19202
rect 3064 19170 3096 19202
rect 3136 19170 3168 19202
rect 3208 19170 3240 19202
rect 3280 19170 3312 19202
rect 3352 19170 3384 19202
rect 3424 19170 3456 19202
rect 3496 19170 3528 19202
rect 3568 19170 3600 19202
rect 3640 19170 3672 19202
rect 3712 19170 3744 19202
rect 3784 19170 3816 19202
rect 3856 19170 3888 19202
rect 112 19098 144 19130
rect 184 19098 216 19130
rect 256 19098 288 19130
rect 328 19098 360 19130
rect 400 19098 432 19130
rect 472 19098 504 19130
rect 544 19098 576 19130
rect 616 19098 648 19130
rect 688 19098 720 19130
rect 760 19098 792 19130
rect 832 19098 864 19130
rect 904 19098 936 19130
rect 976 19098 1008 19130
rect 1048 19098 1080 19130
rect 1120 19098 1152 19130
rect 1192 19098 1224 19130
rect 1264 19098 1296 19130
rect 1336 19098 1368 19130
rect 1408 19098 1440 19130
rect 1480 19098 1512 19130
rect 1552 19098 1584 19130
rect 1624 19098 1656 19130
rect 1696 19098 1728 19130
rect 1768 19098 1800 19130
rect 1840 19098 1872 19130
rect 1912 19098 1944 19130
rect 1984 19098 2016 19130
rect 2056 19098 2088 19130
rect 2128 19098 2160 19130
rect 2200 19098 2232 19130
rect 2272 19098 2304 19130
rect 2344 19098 2376 19130
rect 2416 19098 2448 19130
rect 2488 19098 2520 19130
rect 2560 19098 2592 19130
rect 2632 19098 2664 19130
rect 2704 19098 2736 19130
rect 2776 19098 2808 19130
rect 2848 19098 2880 19130
rect 2920 19098 2952 19130
rect 2992 19098 3024 19130
rect 3064 19098 3096 19130
rect 3136 19098 3168 19130
rect 3208 19098 3240 19130
rect 3280 19098 3312 19130
rect 3352 19098 3384 19130
rect 3424 19098 3456 19130
rect 3496 19098 3528 19130
rect 3568 19098 3600 19130
rect 3640 19098 3672 19130
rect 3712 19098 3744 19130
rect 3784 19098 3816 19130
rect 3856 19098 3888 19130
rect 112 19026 144 19058
rect 184 19026 216 19058
rect 256 19026 288 19058
rect 328 19026 360 19058
rect 400 19026 432 19058
rect 472 19026 504 19058
rect 544 19026 576 19058
rect 616 19026 648 19058
rect 688 19026 720 19058
rect 760 19026 792 19058
rect 832 19026 864 19058
rect 904 19026 936 19058
rect 976 19026 1008 19058
rect 1048 19026 1080 19058
rect 1120 19026 1152 19058
rect 1192 19026 1224 19058
rect 1264 19026 1296 19058
rect 1336 19026 1368 19058
rect 1408 19026 1440 19058
rect 1480 19026 1512 19058
rect 1552 19026 1584 19058
rect 1624 19026 1656 19058
rect 1696 19026 1728 19058
rect 1768 19026 1800 19058
rect 1840 19026 1872 19058
rect 1912 19026 1944 19058
rect 1984 19026 2016 19058
rect 2056 19026 2088 19058
rect 2128 19026 2160 19058
rect 2200 19026 2232 19058
rect 2272 19026 2304 19058
rect 2344 19026 2376 19058
rect 2416 19026 2448 19058
rect 2488 19026 2520 19058
rect 2560 19026 2592 19058
rect 2632 19026 2664 19058
rect 2704 19026 2736 19058
rect 2776 19026 2808 19058
rect 2848 19026 2880 19058
rect 2920 19026 2952 19058
rect 2992 19026 3024 19058
rect 3064 19026 3096 19058
rect 3136 19026 3168 19058
rect 3208 19026 3240 19058
rect 3280 19026 3312 19058
rect 3352 19026 3384 19058
rect 3424 19026 3456 19058
rect 3496 19026 3528 19058
rect 3568 19026 3600 19058
rect 3640 19026 3672 19058
rect 3712 19026 3744 19058
rect 3784 19026 3816 19058
rect 3856 19026 3888 19058
rect 112 18954 144 18986
rect 184 18954 216 18986
rect 256 18954 288 18986
rect 328 18954 360 18986
rect 400 18954 432 18986
rect 472 18954 504 18986
rect 544 18954 576 18986
rect 616 18954 648 18986
rect 688 18954 720 18986
rect 760 18954 792 18986
rect 832 18954 864 18986
rect 904 18954 936 18986
rect 976 18954 1008 18986
rect 1048 18954 1080 18986
rect 1120 18954 1152 18986
rect 1192 18954 1224 18986
rect 1264 18954 1296 18986
rect 1336 18954 1368 18986
rect 1408 18954 1440 18986
rect 1480 18954 1512 18986
rect 1552 18954 1584 18986
rect 1624 18954 1656 18986
rect 1696 18954 1728 18986
rect 1768 18954 1800 18986
rect 1840 18954 1872 18986
rect 1912 18954 1944 18986
rect 1984 18954 2016 18986
rect 2056 18954 2088 18986
rect 2128 18954 2160 18986
rect 2200 18954 2232 18986
rect 2272 18954 2304 18986
rect 2344 18954 2376 18986
rect 2416 18954 2448 18986
rect 2488 18954 2520 18986
rect 2560 18954 2592 18986
rect 2632 18954 2664 18986
rect 2704 18954 2736 18986
rect 2776 18954 2808 18986
rect 2848 18954 2880 18986
rect 2920 18954 2952 18986
rect 2992 18954 3024 18986
rect 3064 18954 3096 18986
rect 3136 18954 3168 18986
rect 3208 18954 3240 18986
rect 3280 18954 3312 18986
rect 3352 18954 3384 18986
rect 3424 18954 3456 18986
rect 3496 18954 3528 18986
rect 3568 18954 3600 18986
rect 3640 18954 3672 18986
rect 3712 18954 3744 18986
rect 3784 18954 3816 18986
rect 3856 18954 3888 18986
rect 112 18882 144 18914
rect 184 18882 216 18914
rect 256 18882 288 18914
rect 328 18882 360 18914
rect 400 18882 432 18914
rect 472 18882 504 18914
rect 544 18882 576 18914
rect 616 18882 648 18914
rect 688 18882 720 18914
rect 760 18882 792 18914
rect 832 18882 864 18914
rect 904 18882 936 18914
rect 976 18882 1008 18914
rect 1048 18882 1080 18914
rect 1120 18882 1152 18914
rect 1192 18882 1224 18914
rect 1264 18882 1296 18914
rect 1336 18882 1368 18914
rect 1408 18882 1440 18914
rect 1480 18882 1512 18914
rect 1552 18882 1584 18914
rect 1624 18882 1656 18914
rect 1696 18882 1728 18914
rect 1768 18882 1800 18914
rect 1840 18882 1872 18914
rect 1912 18882 1944 18914
rect 1984 18882 2016 18914
rect 2056 18882 2088 18914
rect 2128 18882 2160 18914
rect 2200 18882 2232 18914
rect 2272 18882 2304 18914
rect 2344 18882 2376 18914
rect 2416 18882 2448 18914
rect 2488 18882 2520 18914
rect 2560 18882 2592 18914
rect 2632 18882 2664 18914
rect 2704 18882 2736 18914
rect 2776 18882 2808 18914
rect 2848 18882 2880 18914
rect 2920 18882 2952 18914
rect 2992 18882 3024 18914
rect 3064 18882 3096 18914
rect 3136 18882 3168 18914
rect 3208 18882 3240 18914
rect 3280 18882 3312 18914
rect 3352 18882 3384 18914
rect 3424 18882 3456 18914
rect 3496 18882 3528 18914
rect 3568 18882 3600 18914
rect 3640 18882 3672 18914
rect 3712 18882 3744 18914
rect 3784 18882 3816 18914
rect 3856 18882 3888 18914
rect 112 18810 144 18842
rect 184 18810 216 18842
rect 256 18810 288 18842
rect 328 18810 360 18842
rect 400 18810 432 18842
rect 472 18810 504 18842
rect 544 18810 576 18842
rect 616 18810 648 18842
rect 688 18810 720 18842
rect 760 18810 792 18842
rect 832 18810 864 18842
rect 904 18810 936 18842
rect 976 18810 1008 18842
rect 1048 18810 1080 18842
rect 1120 18810 1152 18842
rect 1192 18810 1224 18842
rect 1264 18810 1296 18842
rect 1336 18810 1368 18842
rect 1408 18810 1440 18842
rect 1480 18810 1512 18842
rect 1552 18810 1584 18842
rect 1624 18810 1656 18842
rect 1696 18810 1728 18842
rect 1768 18810 1800 18842
rect 1840 18810 1872 18842
rect 1912 18810 1944 18842
rect 1984 18810 2016 18842
rect 2056 18810 2088 18842
rect 2128 18810 2160 18842
rect 2200 18810 2232 18842
rect 2272 18810 2304 18842
rect 2344 18810 2376 18842
rect 2416 18810 2448 18842
rect 2488 18810 2520 18842
rect 2560 18810 2592 18842
rect 2632 18810 2664 18842
rect 2704 18810 2736 18842
rect 2776 18810 2808 18842
rect 2848 18810 2880 18842
rect 2920 18810 2952 18842
rect 2992 18810 3024 18842
rect 3064 18810 3096 18842
rect 3136 18810 3168 18842
rect 3208 18810 3240 18842
rect 3280 18810 3312 18842
rect 3352 18810 3384 18842
rect 3424 18810 3456 18842
rect 3496 18810 3528 18842
rect 3568 18810 3600 18842
rect 3640 18810 3672 18842
rect 3712 18810 3744 18842
rect 3784 18810 3816 18842
rect 3856 18810 3888 18842
rect 112 18738 144 18770
rect 184 18738 216 18770
rect 256 18738 288 18770
rect 328 18738 360 18770
rect 400 18738 432 18770
rect 472 18738 504 18770
rect 544 18738 576 18770
rect 616 18738 648 18770
rect 688 18738 720 18770
rect 760 18738 792 18770
rect 832 18738 864 18770
rect 904 18738 936 18770
rect 976 18738 1008 18770
rect 1048 18738 1080 18770
rect 1120 18738 1152 18770
rect 1192 18738 1224 18770
rect 1264 18738 1296 18770
rect 1336 18738 1368 18770
rect 1408 18738 1440 18770
rect 1480 18738 1512 18770
rect 1552 18738 1584 18770
rect 1624 18738 1656 18770
rect 1696 18738 1728 18770
rect 1768 18738 1800 18770
rect 1840 18738 1872 18770
rect 1912 18738 1944 18770
rect 1984 18738 2016 18770
rect 2056 18738 2088 18770
rect 2128 18738 2160 18770
rect 2200 18738 2232 18770
rect 2272 18738 2304 18770
rect 2344 18738 2376 18770
rect 2416 18738 2448 18770
rect 2488 18738 2520 18770
rect 2560 18738 2592 18770
rect 2632 18738 2664 18770
rect 2704 18738 2736 18770
rect 2776 18738 2808 18770
rect 2848 18738 2880 18770
rect 2920 18738 2952 18770
rect 2992 18738 3024 18770
rect 3064 18738 3096 18770
rect 3136 18738 3168 18770
rect 3208 18738 3240 18770
rect 3280 18738 3312 18770
rect 3352 18738 3384 18770
rect 3424 18738 3456 18770
rect 3496 18738 3528 18770
rect 3568 18738 3600 18770
rect 3640 18738 3672 18770
rect 3712 18738 3744 18770
rect 3784 18738 3816 18770
rect 3856 18738 3888 18770
rect 112 18666 144 18698
rect 184 18666 216 18698
rect 256 18666 288 18698
rect 328 18666 360 18698
rect 400 18666 432 18698
rect 472 18666 504 18698
rect 544 18666 576 18698
rect 616 18666 648 18698
rect 688 18666 720 18698
rect 760 18666 792 18698
rect 832 18666 864 18698
rect 904 18666 936 18698
rect 976 18666 1008 18698
rect 1048 18666 1080 18698
rect 1120 18666 1152 18698
rect 1192 18666 1224 18698
rect 1264 18666 1296 18698
rect 1336 18666 1368 18698
rect 1408 18666 1440 18698
rect 1480 18666 1512 18698
rect 1552 18666 1584 18698
rect 1624 18666 1656 18698
rect 1696 18666 1728 18698
rect 1768 18666 1800 18698
rect 1840 18666 1872 18698
rect 1912 18666 1944 18698
rect 1984 18666 2016 18698
rect 2056 18666 2088 18698
rect 2128 18666 2160 18698
rect 2200 18666 2232 18698
rect 2272 18666 2304 18698
rect 2344 18666 2376 18698
rect 2416 18666 2448 18698
rect 2488 18666 2520 18698
rect 2560 18666 2592 18698
rect 2632 18666 2664 18698
rect 2704 18666 2736 18698
rect 2776 18666 2808 18698
rect 2848 18666 2880 18698
rect 2920 18666 2952 18698
rect 2992 18666 3024 18698
rect 3064 18666 3096 18698
rect 3136 18666 3168 18698
rect 3208 18666 3240 18698
rect 3280 18666 3312 18698
rect 3352 18666 3384 18698
rect 3424 18666 3456 18698
rect 3496 18666 3528 18698
rect 3568 18666 3600 18698
rect 3640 18666 3672 18698
rect 3712 18666 3744 18698
rect 3784 18666 3816 18698
rect 3856 18666 3888 18698
rect 112 18594 144 18626
rect 184 18594 216 18626
rect 256 18594 288 18626
rect 328 18594 360 18626
rect 400 18594 432 18626
rect 472 18594 504 18626
rect 544 18594 576 18626
rect 616 18594 648 18626
rect 688 18594 720 18626
rect 760 18594 792 18626
rect 832 18594 864 18626
rect 904 18594 936 18626
rect 976 18594 1008 18626
rect 1048 18594 1080 18626
rect 1120 18594 1152 18626
rect 1192 18594 1224 18626
rect 1264 18594 1296 18626
rect 1336 18594 1368 18626
rect 1408 18594 1440 18626
rect 1480 18594 1512 18626
rect 1552 18594 1584 18626
rect 1624 18594 1656 18626
rect 1696 18594 1728 18626
rect 1768 18594 1800 18626
rect 1840 18594 1872 18626
rect 1912 18594 1944 18626
rect 1984 18594 2016 18626
rect 2056 18594 2088 18626
rect 2128 18594 2160 18626
rect 2200 18594 2232 18626
rect 2272 18594 2304 18626
rect 2344 18594 2376 18626
rect 2416 18594 2448 18626
rect 2488 18594 2520 18626
rect 2560 18594 2592 18626
rect 2632 18594 2664 18626
rect 2704 18594 2736 18626
rect 2776 18594 2808 18626
rect 2848 18594 2880 18626
rect 2920 18594 2952 18626
rect 2992 18594 3024 18626
rect 3064 18594 3096 18626
rect 3136 18594 3168 18626
rect 3208 18594 3240 18626
rect 3280 18594 3312 18626
rect 3352 18594 3384 18626
rect 3424 18594 3456 18626
rect 3496 18594 3528 18626
rect 3568 18594 3600 18626
rect 3640 18594 3672 18626
rect 3712 18594 3744 18626
rect 3784 18594 3816 18626
rect 3856 18594 3888 18626
rect 112 18522 144 18554
rect 184 18522 216 18554
rect 256 18522 288 18554
rect 328 18522 360 18554
rect 400 18522 432 18554
rect 472 18522 504 18554
rect 544 18522 576 18554
rect 616 18522 648 18554
rect 688 18522 720 18554
rect 760 18522 792 18554
rect 832 18522 864 18554
rect 904 18522 936 18554
rect 976 18522 1008 18554
rect 1048 18522 1080 18554
rect 1120 18522 1152 18554
rect 1192 18522 1224 18554
rect 1264 18522 1296 18554
rect 1336 18522 1368 18554
rect 1408 18522 1440 18554
rect 1480 18522 1512 18554
rect 1552 18522 1584 18554
rect 1624 18522 1656 18554
rect 1696 18522 1728 18554
rect 1768 18522 1800 18554
rect 1840 18522 1872 18554
rect 1912 18522 1944 18554
rect 1984 18522 2016 18554
rect 2056 18522 2088 18554
rect 2128 18522 2160 18554
rect 2200 18522 2232 18554
rect 2272 18522 2304 18554
rect 2344 18522 2376 18554
rect 2416 18522 2448 18554
rect 2488 18522 2520 18554
rect 2560 18522 2592 18554
rect 2632 18522 2664 18554
rect 2704 18522 2736 18554
rect 2776 18522 2808 18554
rect 2848 18522 2880 18554
rect 2920 18522 2952 18554
rect 2992 18522 3024 18554
rect 3064 18522 3096 18554
rect 3136 18522 3168 18554
rect 3208 18522 3240 18554
rect 3280 18522 3312 18554
rect 3352 18522 3384 18554
rect 3424 18522 3456 18554
rect 3496 18522 3528 18554
rect 3568 18522 3600 18554
rect 3640 18522 3672 18554
rect 3712 18522 3744 18554
rect 3784 18522 3816 18554
rect 3856 18522 3888 18554
rect 112 18450 144 18482
rect 184 18450 216 18482
rect 256 18450 288 18482
rect 328 18450 360 18482
rect 400 18450 432 18482
rect 472 18450 504 18482
rect 544 18450 576 18482
rect 616 18450 648 18482
rect 688 18450 720 18482
rect 760 18450 792 18482
rect 832 18450 864 18482
rect 904 18450 936 18482
rect 976 18450 1008 18482
rect 1048 18450 1080 18482
rect 1120 18450 1152 18482
rect 1192 18450 1224 18482
rect 1264 18450 1296 18482
rect 1336 18450 1368 18482
rect 1408 18450 1440 18482
rect 1480 18450 1512 18482
rect 1552 18450 1584 18482
rect 1624 18450 1656 18482
rect 1696 18450 1728 18482
rect 1768 18450 1800 18482
rect 1840 18450 1872 18482
rect 1912 18450 1944 18482
rect 1984 18450 2016 18482
rect 2056 18450 2088 18482
rect 2128 18450 2160 18482
rect 2200 18450 2232 18482
rect 2272 18450 2304 18482
rect 2344 18450 2376 18482
rect 2416 18450 2448 18482
rect 2488 18450 2520 18482
rect 2560 18450 2592 18482
rect 2632 18450 2664 18482
rect 2704 18450 2736 18482
rect 2776 18450 2808 18482
rect 2848 18450 2880 18482
rect 2920 18450 2952 18482
rect 2992 18450 3024 18482
rect 3064 18450 3096 18482
rect 3136 18450 3168 18482
rect 3208 18450 3240 18482
rect 3280 18450 3312 18482
rect 3352 18450 3384 18482
rect 3424 18450 3456 18482
rect 3496 18450 3528 18482
rect 3568 18450 3600 18482
rect 3640 18450 3672 18482
rect 3712 18450 3744 18482
rect 3784 18450 3816 18482
rect 3856 18450 3888 18482
rect 112 18378 144 18410
rect 184 18378 216 18410
rect 256 18378 288 18410
rect 328 18378 360 18410
rect 400 18378 432 18410
rect 472 18378 504 18410
rect 544 18378 576 18410
rect 616 18378 648 18410
rect 688 18378 720 18410
rect 760 18378 792 18410
rect 832 18378 864 18410
rect 904 18378 936 18410
rect 976 18378 1008 18410
rect 1048 18378 1080 18410
rect 1120 18378 1152 18410
rect 1192 18378 1224 18410
rect 1264 18378 1296 18410
rect 1336 18378 1368 18410
rect 1408 18378 1440 18410
rect 1480 18378 1512 18410
rect 1552 18378 1584 18410
rect 1624 18378 1656 18410
rect 1696 18378 1728 18410
rect 1768 18378 1800 18410
rect 1840 18378 1872 18410
rect 1912 18378 1944 18410
rect 1984 18378 2016 18410
rect 2056 18378 2088 18410
rect 2128 18378 2160 18410
rect 2200 18378 2232 18410
rect 2272 18378 2304 18410
rect 2344 18378 2376 18410
rect 2416 18378 2448 18410
rect 2488 18378 2520 18410
rect 2560 18378 2592 18410
rect 2632 18378 2664 18410
rect 2704 18378 2736 18410
rect 2776 18378 2808 18410
rect 2848 18378 2880 18410
rect 2920 18378 2952 18410
rect 2992 18378 3024 18410
rect 3064 18378 3096 18410
rect 3136 18378 3168 18410
rect 3208 18378 3240 18410
rect 3280 18378 3312 18410
rect 3352 18378 3384 18410
rect 3424 18378 3456 18410
rect 3496 18378 3528 18410
rect 3568 18378 3600 18410
rect 3640 18378 3672 18410
rect 3712 18378 3744 18410
rect 3784 18378 3816 18410
rect 3856 18378 3888 18410
rect 112 18306 144 18338
rect 184 18306 216 18338
rect 256 18306 288 18338
rect 328 18306 360 18338
rect 400 18306 432 18338
rect 472 18306 504 18338
rect 544 18306 576 18338
rect 616 18306 648 18338
rect 688 18306 720 18338
rect 760 18306 792 18338
rect 832 18306 864 18338
rect 904 18306 936 18338
rect 976 18306 1008 18338
rect 1048 18306 1080 18338
rect 1120 18306 1152 18338
rect 1192 18306 1224 18338
rect 1264 18306 1296 18338
rect 1336 18306 1368 18338
rect 1408 18306 1440 18338
rect 1480 18306 1512 18338
rect 1552 18306 1584 18338
rect 1624 18306 1656 18338
rect 1696 18306 1728 18338
rect 1768 18306 1800 18338
rect 1840 18306 1872 18338
rect 1912 18306 1944 18338
rect 1984 18306 2016 18338
rect 2056 18306 2088 18338
rect 2128 18306 2160 18338
rect 2200 18306 2232 18338
rect 2272 18306 2304 18338
rect 2344 18306 2376 18338
rect 2416 18306 2448 18338
rect 2488 18306 2520 18338
rect 2560 18306 2592 18338
rect 2632 18306 2664 18338
rect 2704 18306 2736 18338
rect 2776 18306 2808 18338
rect 2848 18306 2880 18338
rect 2920 18306 2952 18338
rect 2992 18306 3024 18338
rect 3064 18306 3096 18338
rect 3136 18306 3168 18338
rect 3208 18306 3240 18338
rect 3280 18306 3312 18338
rect 3352 18306 3384 18338
rect 3424 18306 3456 18338
rect 3496 18306 3528 18338
rect 3568 18306 3600 18338
rect 3640 18306 3672 18338
rect 3712 18306 3744 18338
rect 3784 18306 3816 18338
rect 3856 18306 3888 18338
rect 112 18234 144 18266
rect 184 18234 216 18266
rect 256 18234 288 18266
rect 328 18234 360 18266
rect 400 18234 432 18266
rect 472 18234 504 18266
rect 544 18234 576 18266
rect 616 18234 648 18266
rect 688 18234 720 18266
rect 760 18234 792 18266
rect 832 18234 864 18266
rect 904 18234 936 18266
rect 976 18234 1008 18266
rect 1048 18234 1080 18266
rect 1120 18234 1152 18266
rect 1192 18234 1224 18266
rect 1264 18234 1296 18266
rect 1336 18234 1368 18266
rect 1408 18234 1440 18266
rect 1480 18234 1512 18266
rect 1552 18234 1584 18266
rect 1624 18234 1656 18266
rect 1696 18234 1728 18266
rect 1768 18234 1800 18266
rect 1840 18234 1872 18266
rect 1912 18234 1944 18266
rect 1984 18234 2016 18266
rect 2056 18234 2088 18266
rect 2128 18234 2160 18266
rect 2200 18234 2232 18266
rect 2272 18234 2304 18266
rect 2344 18234 2376 18266
rect 2416 18234 2448 18266
rect 2488 18234 2520 18266
rect 2560 18234 2592 18266
rect 2632 18234 2664 18266
rect 2704 18234 2736 18266
rect 2776 18234 2808 18266
rect 2848 18234 2880 18266
rect 2920 18234 2952 18266
rect 2992 18234 3024 18266
rect 3064 18234 3096 18266
rect 3136 18234 3168 18266
rect 3208 18234 3240 18266
rect 3280 18234 3312 18266
rect 3352 18234 3384 18266
rect 3424 18234 3456 18266
rect 3496 18234 3528 18266
rect 3568 18234 3600 18266
rect 3640 18234 3672 18266
rect 3712 18234 3744 18266
rect 3784 18234 3816 18266
rect 3856 18234 3888 18266
rect 112 18162 144 18194
rect 184 18162 216 18194
rect 256 18162 288 18194
rect 328 18162 360 18194
rect 400 18162 432 18194
rect 472 18162 504 18194
rect 544 18162 576 18194
rect 616 18162 648 18194
rect 688 18162 720 18194
rect 760 18162 792 18194
rect 832 18162 864 18194
rect 904 18162 936 18194
rect 976 18162 1008 18194
rect 1048 18162 1080 18194
rect 1120 18162 1152 18194
rect 1192 18162 1224 18194
rect 1264 18162 1296 18194
rect 1336 18162 1368 18194
rect 1408 18162 1440 18194
rect 1480 18162 1512 18194
rect 1552 18162 1584 18194
rect 1624 18162 1656 18194
rect 1696 18162 1728 18194
rect 1768 18162 1800 18194
rect 1840 18162 1872 18194
rect 1912 18162 1944 18194
rect 1984 18162 2016 18194
rect 2056 18162 2088 18194
rect 2128 18162 2160 18194
rect 2200 18162 2232 18194
rect 2272 18162 2304 18194
rect 2344 18162 2376 18194
rect 2416 18162 2448 18194
rect 2488 18162 2520 18194
rect 2560 18162 2592 18194
rect 2632 18162 2664 18194
rect 2704 18162 2736 18194
rect 2776 18162 2808 18194
rect 2848 18162 2880 18194
rect 2920 18162 2952 18194
rect 2992 18162 3024 18194
rect 3064 18162 3096 18194
rect 3136 18162 3168 18194
rect 3208 18162 3240 18194
rect 3280 18162 3312 18194
rect 3352 18162 3384 18194
rect 3424 18162 3456 18194
rect 3496 18162 3528 18194
rect 3568 18162 3600 18194
rect 3640 18162 3672 18194
rect 3712 18162 3744 18194
rect 3784 18162 3816 18194
rect 3856 18162 3888 18194
rect 184 17816 216 17848
rect 256 17816 288 17848
rect 328 17816 360 17848
rect 400 17816 432 17848
rect 472 17816 504 17848
rect 544 17816 576 17848
rect 616 17816 648 17848
rect 688 17816 720 17848
rect 760 17816 792 17848
rect 832 17816 864 17848
rect 904 17816 936 17848
rect 976 17816 1008 17848
rect 1048 17816 1080 17848
rect 1120 17816 1152 17848
rect 1192 17816 1224 17848
rect 1264 17816 1296 17848
rect 1336 17816 1368 17848
rect 1408 17816 1440 17848
rect 1480 17816 1512 17848
rect 1552 17816 1584 17848
rect 1624 17816 1656 17848
rect 1696 17816 1728 17848
rect 1768 17816 1800 17848
rect 1840 17816 1872 17848
rect 1912 17816 1944 17848
rect 1984 17816 2016 17848
rect 2056 17816 2088 17848
rect 2128 17816 2160 17848
rect 2200 17816 2232 17848
rect 2272 17816 2304 17848
rect 2344 17816 2376 17848
rect 2416 17816 2448 17848
rect 2488 17816 2520 17848
rect 2560 17816 2592 17848
rect 2632 17816 2664 17848
rect 2704 17816 2736 17848
rect 2776 17816 2808 17848
rect 2848 17816 2880 17848
rect 2920 17816 2952 17848
rect 2992 17816 3024 17848
rect 3064 17816 3096 17848
rect 3136 17816 3168 17848
rect 3208 17816 3240 17848
rect 3280 17816 3312 17848
rect 3352 17816 3384 17848
rect 3424 17816 3456 17848
rect 3496 17816 3528 17848
rect 3568 17816 3600 17848
rect 3640 17816 3672 17848
rect 3712 17816 3744 17848
rect 3784 17816 3816 17848
rect 3856 17816 3888 17848
rect 112 17744 144 17776
rect 184 17744 216 17776
rect 256 17744 288 17776
rect 328 17744 360 17776
rect 400 17744 432 17776
rect 472 17744 504 17776
rect 544 17744 576 17776
rect 616 17744 648 17776
rect 688 17744 720 17776
rect 760 17744 792 17776
rect 832 17744 864 17776
rect 904 17744 936 17776
rect 976 17744 1008 17776
rect 1048 17744 1080 17776
rect 1120 17744 1152 17776
rect 1192 17744 1224 17776
rect 1264 17744 1296 17776
rect 1336 17744 1368 17776
rect 1408 17744 1440 17776
rect 1480 17744 1512 17776
rect 1552 17744 1584 17776
rect 1624 17744 1656 17776
rect 1696 17744 1728 17776
rect 1768 17744 1800 17776
rect 1840 17744 1872 17776
rect 1912 17744 1944 17776
rect 1984 17744 2016 17776
rect 2056 17744 2088 17776
rect 2128 17744 2160 17776
rect 2200 17744 2232 17776
rect 2272 17744 2304 17776
rect 2344 17744 2376 17776
rect 2416 17744 2448 17776
rect 2488 17744 2520 17776
rect 2560 17744 2592 17776
rect 2632 17744 2664 17776
rect 2704 17744 2736 17776
rect 2776 17744 2808 17776
rect 2848 17744 2880 17776
rect 2920 17744 2952 17776
rect 2992 17744 3024 17776
rect 3064 17744 3096 17776
rect 3136 17744 3168 17776
rect 3208 17744 3240 17776
rect 3280 17744 3312 17776
rect 3352 17744 3384 17776
rect 3424 17744 3456 17776
rect 3496 17744 3528 17776
rect 3568 17744 3600 17776
rect 3640 17744 3672 17776
rect 3712 17744 3744 17776
rect 3784 17744 3816 17776
rect 3856 17744 3888 17776
rect 112 17672 144 17704
rect 184 17672 216 17704
rect 256 17672 288 17704
rect 328 17672 360 17704
rect 400 17672 432 17704
rect 472 17672 504 17704
rect 544 17672 576 17704
rect 616 17672 648 17704
rect 688 17672 720 17704
rect 760 17672 792 17704
rect 832 17672 864 17704
rect 904 17672 936 17704
rect 976 17672 1008 17704
rect 1048 17672 1080 17704
rect 1120 17672 1152 17704
rect 1192 17672 1224 17704
rect 1264 17672 1296 17704
rect 1336 17672 1368 17704
rect 1408 17672 1440 17704
rect 1480 17672 1512 17704
rect 1552 17672 1584 17704
rect 1624 17672 1656 17704
rect 1696 17672 1728 17704
rect 1768 17672 1800 17704
rect 1840 17672 1872 17704
rect 1912 17672 1944 17704
rect 1984 17672 2016 17704
rect 2056 17672 2088 17704
rect 2128 17672 2160 17704
rect 2200 17672 2232 17704
rect 2272 17672 2304 17704
rect 2344 17672 2376 17704
rect 2416 17672 2448 17704
rect 2488 17672 2520 17704
rect 2560 17672 2592 17704
rect 2632 17672 2664 17704
rect 2704 17672 2736 17704
rect 2776 17672 2808 17704
rect 2848 17672 2880 17704
rect 2920 17672 2952 17704
rect 2992 17672 3024 17704
rect 3064 17672 3096 17704
rect 3136 17672 3168 17704
rect 3208 17672 3240 17704
rect 3280 17672 3312 17704
rect 3352 17672 3384 17704
rect 3424 17672 3456 17704
rect 3496 17672 3528 17704
rect 3568 17672 3600 17704
rect 3640 17672 3672 17704
rect 3712 17672 3744 17704
rect 3784 17672 3816 17704
rect 3856 17672 3888 17704
rect 112 17600 144 17632
rect 184 17600 216 17632
rect 256 17600 288 17632
rect 328 17600 360 17632
rect 400 17600 432 17632
rect 472 17600 504 17632
rect 544 17600 576 17632
rect 616 17600 648 17632
rect 688 17600 720 17632
rect 760 17600 792 17632
rect 832 17600 864 17632
rect 904 17600 936 17632
rect 976 17600 1008 17632
rect 1048 17600 1080 17632
rect 1120 17600 1152 17632
rect 1192 17600 1224 17632
rect 1264 17600 1296 17632
rect 1336 17600 1368 17632
rect 1408 17600 1440 17632
rect 1480 17600 1512 17632
rect 1552 17600 1584 17632
rect 1624 17600 1656 17632
rect 1696 17600 1728 17632
rect 1768 17600 1800 17632
rect 1840 17600 1872 17632
rect 1912 17600 1944 17632
rect 1984 17600 2016 17632
rect 2056 17600 2088 17632
rect 2128 17600 2160 17632
rect 2200 17600 2232 17632
rect 2272 17600 2304 17632
rect 2344 17600 2376 17632
rect 2416 17600 2448 17632
rect 2488 17600 2520 17632
rect 2560 17600 2592 17632
rect 2632 17600 2664 17632
rect 2704 17600 2736 17632
rect 2776 17600 2808 17632
rect 2848 17600 2880 17632
rect 2920 17600 2952 17632
rect 2992 17600 3024 17632
rect 3064 17600 3096 17632
rect 3136 17600 3168 17632
rect 3208 17600 3240 17632
rect 3280 17600 3312 17632
rect 3352 17600 3384 17632
rect 3424 17600 3456 17632
rect 3496 17600 3528 17632
rect 3568 17600 3600 17632
rect 3640 17600 3672 17632
rect 3712 17600 3744 17632
rect 3784 17600 3816 17632
rect 3856 17600 3888 17632
rect 112 17528 144 17560
rect 184 17528 216 17560
rect 256 17528 288 17560
rect 328 17528 360 17560
rect 400 17528 432 17560
rect 472 17528 504 17560
rect 544 17528 576 17560
rect 616 17528 648 17560
rect 688 17528 720 17560
rect 760 17528 792 17560
rect 832 17528 864 17560
rect 904 17528 936 17560
rect 976 17528 1008 17560
rect 1048 17528 1080 17560
rect 1120 17528 1152 17560
rect 1192 17528 1224 17560
rect 1264 17528 1296 17560
rect 1336 17528 1368 17560
rect 1408 17528 1440 17560
rect 1480 17528 1512 17560
rect 1552 17528 1584 17560
rect 1624 17528 1656 17560
rect 1696 17528 1728 17560
rect 1768 17528 1800 17560
rect 1840 17528 1872 17560
rect 1912 17528 1944 17560
rect 1984 17528 2016 17560
rect 2056 17528 2088 17560
rect 2128 17528 2160 17560
rect 2200 17528 2232 17560
rect 2272 17528 2304 17560
rect 2344 17528 2376 17560
rect 2416 17528 2448 17560
rect 2488 17528 2520 17560
rect 2560 17528 2592 17560
rect 2632 17528 2664 17560
rect 2704 17528 2736 17560
rect 2776 17528 2808 17560
rect 2848 17528 2880 17560
rect 2920 17528 2952 17560
rect 2992 17528 3024 17560
rect 3064 17528 3096 17560
rect 3136 17528 3168 17560
rect 3208 17528 3240 17560
rect 3280 17528 3312 17560
rect 3352 17528 3384 17560
rect 3424 17528 3456 17560
rect 3496 17528 3528 17560
rect 3568 17528 3600 17560
rect 3640 17528 3672 17560
rect 3712 17528 3744 17560
rect 3784 17528 3816 17560
rect 3856 17528 3888 17560
rect 112 17456 144 17488
rect 184 17456 216 17488
rect 256 17456 288 17488
rect 328 17456 360 17488
rect 400 17456 432 17488
rect 472 17456 504 17488
rect 544 17456 576 17488
rect 616 17456 648 17488
rect 688 17456 720 17488
rect 760 17456 792 17488
rect 832 17456 864 17488
rect 904 17456 936 17488
rect 976 17456 1008 17488
rect 1048 17456 1080 17488
rect 1120 17456 1152 17488
rect 1192 17456 1224 17488
rect 1264 17456 1296 17488
rect 1336 17456 1368 17488
rect 1408 17456 1440 17488
rect 1480 17456 1512 17488
rect 1552 17456 1584 17488
rect 1624 17456 1656 17488
rect 1696 17456 1728 17488
rect 1768 17456 1800 17488
rect 1840 17456 1872 17488
rect 1912 17456 1944 17488
rect 1984 17456 2016 17488
rect 2056 17456 2088 17488
rect 2128 17456 2160 17488
rect 2200 17456 2232 17488
rect 2272 17456 2304 17488
rect 2344 17456 2376 17488
rect 2416 17456 2448 17488
rect 2488 17456 2520 17488
rect 2560 17456 2592 17488
rect 2632 17456 2664 17488
rect 2704 17456 2736 17488
rect 2776 17456 2808 17488
rect 2848 17456 2880 17488
rect 2920 17456 2952 17488
rect 2992 17456 3024 17488
rect 3064 17456 3096 17488
rect 3136 17456 3168 17488
rect 3208 17456 3240 17488
rect 3280 17456 3312 17488
rect 3352 17456 3384 17488
rect 3424 17456 3456 17488
rect 3496 17456 3528 17488
rect 3568 17456 3600 17488
rect 3640 17456 3672 17488
rect 3712 17456 3744 17488
rect 3784 17456 3816 17488
rect 3856 17456 3888 17488
rect 112 17384 144 17416
rect 184 17384 216 17416
rect 256 17384 288 17416
rect 328 17384 360 17416
rect 400 17384 432 17416
rect 472 17384 504 17416
rect 544 17384 576 17416
rect 616 17384 648 17416
rect 688 17384 720 17416
rect 760 17384 792 17416
rect 832 17384 864 17416
rect 904 17384 936 17416
rect 976 17384 1008 17416
rect 1048 17384 1080 17416
rect 1120 17384 1152 17416
rect 1192 17384 1224 17416
rect 1264 17384 1296 17416
rect 1336 17384 1368 17416
rect 1408 17384 1440 17416
rect 1480 17384 1512 17416
rect 1552 17384 1584 17416
rect 1624 17384 1656 17416
rect 1696 17384 1728 17416
rect 1768 17384 1800 17416
rect 1840 17384 1872 17416
rect 1912 17384 1944 17416
rect 1984 17384 2016 17416
rect 2056 17384 2088 17416
rect 2128 17384 2160 17416
rect 2200 17384 2232 17416
rect 2272 17384 2304 17416
rect 2344 17384 2376 17416
rect 2416 17384 2448 17416
rect 2488 17384 2520 17416
rect 2560 17384 2592 17416
rect 2632 17384 2664 17416
rect 2704 17384 2736 17416
rect 2776 17384 2808 17416
rect 2848 17384 2880 17416
rect 2920 17384 2952 17416
rect 2992 17384 3024 17416
rect 3064 17384 3096 17416
rect 3136 17384 3168 17416
rect 3208 17384 3240 17416
rect 3280 17384 3312 17416
rect 3352 17384 3384 17416
rect 3424 17384 3456 17416
rect 3496 17384 3528 17416
rect 3568 17384 3600 17416
rect 3640 17384 3672 17416
rect 3712 17384 3744 17416
rect 3784 17384 3816 17416
rect 3856 17384 3888 17416
rect 112 17312 144 17344
rect 184 17312 216 17344
rect 256 17312 288 17344
rect 328 17312 360 17344
rect 400 17312 432 17344
rect 472 17312 504 17344
rect 544 17312 576 17344
rect 616 17312 648 17344
rect 688 17312 720 17344
rect 760 17312 792 17344
rect 832 17312 864 17344
rect 904 17312 936 17344
rect 976 17312 1008 17344
rect 1048 17312 1080 17344
rect 1120 17312 1152 17344
rect 1192 17312 1224 17344
rect 1264 17312 1296 17344
rect 1336 17312 1368 17344
rect 1408 17312 1440 17344
rect 1480 17312 1512 17344
rect 1552 17312 1584 17344
rect 1624 17312 1656 17344
rect 1696 17312 1728 17344
rect 1768 17312 1800 17344
rect 1840 17312 1872 17344
rect 1912 17312 1944 17344
rect 1984 17312 2016 17344
rect 2056 17312 2088 17344
rect 2128 17312 2160 17344
rect 2200 17312 2232 17344
rect 2272 17312 2304 17344
rect 2344 17312 2376 17344
rect 2416 17312 2448 17344
rect 2488 17312 2520 17344
rect 2560 17312 2592 17344
rect 2632 17312 2664 17344
rect 2704 17312 2736 17344
rect 2776 17312 2808 17344
rect 2848 17312 2880 17344
rect 2920 17312 2952 17344
rect 2992 17312 3024 17344
rect 3064 17312 3096 17344
rect 3136 17312 3168 17344
rect 3208 17312 3240 17344
rect 3280 17312 3312 17344
rect 3352 17312 3384 17344
rect 3424 17312 3456 17344
rect 3496 17312 3528 17344
rect 3568 17312 3600 17344
rect 3640 17312 3672 17344
rect 3712 17312 3744 17344
rect 3784 17312 3816 17344
rect 3856 17312 3888 17344
rect 112 17240 144 17272
rect 184 17240 216 17272
rect 256 17240 288 17272
rect 328 17240 360 17272
rect 400 17240 432 17272
rect 472 17240 504 17272
rect 544 17240 576 17272
rect 616 17240 648 17272
rect 688 17240 720 17272
rect 760 17240 792 17272
rect 832 17240 864 17272
rect 904 17240 936 17272
rect 976 17240 1008 17272
rect 1048 17240 1080 17272
rect 1120 17240 1152 17272
rect 1192 17240 1224 17272
rect 1264 17240 1296 17272
rect 1336 17240 1368 17272
rect 1408 17240 1440 17272
rect 1480 17240 1512 17272
rect 1552 17240 1584 17272
rect 1624 17240 1656 17272
rect 1696 17240 1728 17272
rect 1768 17240 1800 17272
rect 1840 17240 1872 17272
rect 1912 17240 1944 17272
rect 1984 17240 2016 17272
rect 2056 17240 2088 17272
rect 2128 17240 2160 17272
rect 2200 17240 2232 17272
rect 2272 17240 2304 17272
rect 2344 17240 2376 17272
rect 2416 17240 2448 17272
rect 2488 17240 2520 17272
rect 2560 17240 2592 17272
rect 2632 17240 2664 17272
rect 2704 17240 2736 17272
rect 2776 17240 2808 17272
rect 2848 17240 2880 17272
rect 2920 17240 2952 17272
rect 2992 17240 3024 17272
rect 3064 17240 3096 17272
rect 3136 17240 3168 17272
rect 3208 17240 3240 17272
rect 3280 17240 3312 17272
rect 3352 17240 3384 17272
rect 3424 17240 3456 17272
rect 3496 17240 3528 17272
rect 3568 17240 3600 17272
rect 3640 17240 3672 17272
rect 3712 17240 3744 17272
rect 3784 17240 3816 17272
rect 3856 17240 3888 17272
rect 112 17168 144 17200
rect 184 17168 216 17200
rect 256 17168 288 17200
rect 328 17168 360 17200
rect 400 17168 432 17200
rect 472 17168 504 17200
rect 544 17168 576 17200
rect 616 17168 648 17200
rect 688 17168 720 17200
rect 760 17168 792 17200
rect 832 17168 864 17200
rect 904 17168 936 17200
rect 976 17168 1008 17200
rect 1048 17168 1080 17200
rect 1120 17168 1152 17200
rect 1192 17168 1224 17200
rect 1264 17168 1296 17200
rect 1336 17168 1368 17200
rect 1408 17168 1440 17200
rect 1480 17168 1512 17200
rect 1552 17168 1584 17200
rect 1624 17168 1656 17200
rect 1696 17168 1728 17200
rect 1768 17168 1800 17200
rect 1840 17168 1872 17200
rect 1912 17168 1944 17200
rect 1984 17168 2016 17200
rect 2056 17168 2088 17200
rect 2128 17168 2160 17200
rect 2200 17168 2232 17200
rect 2272 17168 2304 17200
rect 2344 17168 2376 17200
rect 2416 17168 2448 17200
rect 2488 17168 2520 17200
rect 2560 17168 2592 17200
rect 2632 17168 2664 17200
rect 2704 17168 2736 17200
rect 2776 17168 2808 17200
rect 2848 17168 2880 17200
rect 2920 17168 2952 17200
rect 2992 17168 3024 17200
rect 3064 17168 3096 17200
rect 3136 17168 3168 17200
rect 3208 17168 3240 17200
rect 3280 17168 3312 17200
rect 3352 17168 3384 17200
rect 3424 17168 3456 17200
rect 3496 17168 3528 17200
rect 3568 17168 3600 17200
rect 3640 17168 3672 17200
rect 3712 17168 3744 17200
rect 3784 17168 3816 17200
rect 3856 17168 3888 17200
rect 112 17096 144 17128
rect 184 17096 216 17128
rect 256 17096 288 17128
rect 328 17096 360 17128
rect 400 17096 432 17128
rect 472 17096 504 17128
rect 544 17096 576 17128
rect 616 17096 648 17128
rect 688 17096 720 17128
rect 760 17096 792 17128
rect 832 17096 864 17128
rect 904 17096 936 17128
rect 976 17096 1008 17128
rect 1048 17096 1080 17128
rect 1120 17096 1152 17128
rect 1192 17096 1224 17128
rect 1264 17096 1296 17128
rect 1336 17096 1368 17128
rect 1408 17096 1440 17128
rect 1480 17096 1512 17128
rect 1552 17096 1584 17128
rect 1624 17096 1656 17128
rect 1696 17096 1728 17128
rect 1768 17096 1800 17128
rect 1840 17096 1872 17128
rect 1912 17096 1944 17128
rect 1984 17096 2016 17128
rect 2056 17096 2088 17128
rect 2128 17096 2160 17128
rect 2200 17096 2232 17128
rect 2272 17096 2304 17128
rect 2344 17096 2376 17128
rect 2416 17096 2448 17128
rect 2488 17096 2520 17128
rect 2560 17096 2592 17128
rect 2632 17096 2664 17128
rect 2704 17096 2736 17128
rect 2776 17096 2808 17128
rect 2848 17096 2880 17128
rect 2920 17096 2952 17128
rect 2992 17096 3024 17128
rect 3064 17096 3096 17128
rect 3136 17096 3168 17128
rect 3208 17096 3240 17128
rect 3280 17096 3312 17128
rect 3352 17096 3384 17128
rect 3424 17096 3456 17128
rect 3496 17096 3528 17128
rect 3568 17096 3600 17128
rect 3640 17096 3672 17128
rect 3712 17096 3744 17128
rect 3784 17096 3816 17128
rect 3856 17096 3888 17128
rect 112 17024 144 17056
rect 184 17024 216 17056
rect 256 17024 288 17056
rect 328 17024 360 17056
rect 400 17024 432 17056
rect 472 17024 504 17056
rect 544 17024 576 17056
rect 616 17024 648 17056
rect 688 17024 720 17056
rect 760 17024 792 17056
rect 832 17024 864 17056
rect 904 17024 936 17056
rect 976 17024 1008 17056
rect 1048 17024 1080 17056
rect 1120 17024 1152 17056
rect 1192 17024 1224 17056
rect 1264 17024 1296 17056
rect 1336 17024 1368 17056
rect 1408 17024 1440 17056
rect 1480 17024 1512 17056
rect 1552 17024 1584 17056
rect 1624 17024 1656 17056
rect 1696 17024 1728 17056
rect 1768 17024 1800 17056
rect 1840 17024 1872 17056
rect 1912 17024 1944 17056
rect 1984 17024 2016 17056
rect 2056 17024 2088 17056
rect 2128 17024 2160 17056
rect 2200 17024 2232 17056
rect 2272 17024 2304 17056
rect 2344 17024 2376 17056
rect 2416 17024 2448 17056
rect 2488 17024 2520 17056
rect 2560 17024 2592 17056
rect 2632 17024 2664 17056
rect 2704 17024 2736 17056
rect 2776 17024 2808 17056
rect 2848 17024 2880 17056
rect 2920 17024 2952 17056
rect 2992 17024 3024 17056
rect 3064 17024 3096 17056
rect 3136 17024 3168 17056
rect 3208 17024 3240 17056
rect 3280 17024 3312 17056
rect 3352 17024 3384 17056
rect 3424 17024 3456 17056
rect 3496 17024 3528 17056
rect 3568 17024 3600 17056
rect 3640 17024 3672 17056
rect 3712 17024 3744 17056
rect 3784 17024 3816 17056
rect 3856 17024 3888 17056
rect 112 16952 144 16984
rect 184 16952 216 16984
rect 256 16952 288 16984
rect 328 16952 360 16984
rect 400 16952 432 16984
rect 472 16952 504 16984
rect 544 16952 576 16984
rect 616 16952 648 16984
rect 688 16952 720 16984
rect 760 16952 792 16984
rect 832 16952 864 16984
rect 904 16952 936 16984
rect 976 16952 1008 16984
rect 1048 16952 1080 16984
rect 1120 16952 1152 16984
rect 1192 16952 1224 16984
rect 1264 16952 1296 16984
rect 1336 16952 1368 16984
rect 1408 16952 1440 16984
rect 1480 16952 1512 16984
rect 1552 16952 1584 16984
rect 1624 16952 1656 16984
rect 1696 16952 1728 16984
rect 1768 16952 1800 16984
rect 1840 16952 1872 16984
rect 1912 16952 1944 16984
rect 1984 16952 2016 16984
rect 2056 16952 2088 16984
rect 2128 16952 2160 16984
rect 2200 16952 2232 16984
rect 2272 16952 2304 16984
rect 2344 16952 2376 16984
rect 2416 16952 2448 16984
rect 2488 16952 2520 16984
rect 2560 16952 2592 16984
rect 2632 16952 2664 16984
rect 2704 16952 2736 16984
rect 2776 16952 2808 16984
rect 2848 16952 2880 16984
rect 2920 16952 2952 16984
rect 2992 16952 3024 16984
rect 3064 16952 3096 16984
rect 3136 16952 3168 16984
rect 3208 16952 3240 16984
rect 3280 16952 3312 16984
rect 3352 16952 3384 16984
rect 3424 16952 3456 16984
rect 3496 16952 3528 16984
rect 3568 16952 3600 16984
rect 3640 16952 3672 16984
rect 3712 16952 3744 16984
rect 3784 16952 3816 16984
rect 3856 16952 3888 16984
rect 112 16880 144 16912
rect 184 16880 216 16912
rect 256 16880 288 16912
rect 328 16880 360 16912
rect 400 16880 432 16912
rect 472 16880 504 16912
rect 544 16880 576 16912
rect 616 16880 648 16912
rect 688 16880 720 16912
rect 760 16880 792 16912
rect 832 16880 864 16912
rect 904 16880 936 16912
rect 976 16880 1008 16912
rect 1048 16880 1080 16912
rect 1120 16880 1152 16912
rect 1192 16880 1224 16912
rect 1264 16880 1296 16912
rect 1336 16880 1368 16912
rect 1408 16880 1440 16912
rect 1480 16880 1512 16912
rect 1552 16880 1584 16912
rect 1624 16880 1656 16912
rect 1696 16880 1728 16912
rect 1768 16880 1800 16912
rect 1840 16880 1872 16912
rect 1912 16880 1944 16912
rect 1984 16880 2016 16912
rect 2056 16880 2088 16912
rect 2128 16880 2160 16912
rect 2200 16880 2232 16912
rect 2272 16880 2304 16912
rect 2344 16880 2376 16912
rect 2416 16880 2448 16912
rect 2488 16880 2520 16912
rect 2560 16880 2592 16912
rect 2632 16880 2664 16912
rect 2704 16880 2736 16912
rect 2776 16880 2808 16912
rect 2848 16880 2880 16912
rect 2920 16880 2952 16912
rect 2992 16880 3024 16912
rect 3064 16880 3096 16912
rect 3136 16880 3168 16912
rect 3208 16880 3240 16912
rect 3280 16880 3312 16912
rect 3352 16880 3384 16912
rect 3424 16880 3456 16912
rect 3496 16880 3528 16912
rect 3568 16880 3600 16912
rect 3640 16880 3672 16912
rect 3712 16880 3744 16912
rect 3784 16880 3816 16912
rect 3856 16880 3888 16912
rect 112 16808 144 16840
rect 184 16808 216 16840
rect 256 16808 288 16840
rect 328 16808 360 16840
rect 400 16808 432 16840
rect 472 16808 504 16840
rect 544 16808 576 16840
rect 616 16808 648 16840
rect 688 16808 720 16840
rect 760 16808 792 16840
rect 832 16808 864 16840
rect 904 16808 936 16840
rect 976 16808 1008 16840
rect 1048 16808 1080 16840
rect 1120 16808 1152 16840
rect 1192 16808 1224 16840
rect 1264 16808 1296 16840
rect 1336 16808 1368 16840
rect 1408 16808 1440 16840
rect 1480 16808 1512 16840
rect 1552 16808 1584 16840
rect 1624 16808 1656 16840
rect 1696 16808 1728 16840
rect 1768 16808 1800 16840
rect 1840 16808 1872 16840
rect 1912 16808 1944 16840
rect 1984 16808 2016 16840
rect 2056 16808 2088 16840
rect 2128 16808 2160 16840
rect 2200 16808 2232 16840
rect 2272 16808 2304 16840
rect 2344 16808 2376 16840
rect 2416 16808 2448 16840
rect 2488 16808 2520 16840
rect 2560 16808 2592 16840
rect 2632 16808 2664 16840
rect 2704 16808 2736 16840
rect 2776 16808 2808 16840
rect 2848 16808 2880 16840
rect 2920 16808 2952 16840
rect 2992 16808 3024 16840
rect 3064 16808 3096 16840
rect 3136 16808 3168 16840
rect 3208 16808 3240 16840
rect 3280 16808 3312 16840
rect 3352 16808 3384 16840
rect 3424 16808 3456 16840
rect 3496 16808 3528 16840
rect 3568 16808 3600 16840
rect 3640 16808 3672 16840
rect 3712 16808 3744 16840
rect 3784 16808 3816 16840
rect 3856 16808 3888 16840
rect 112 16736 144 16768
rect 184 16736 216 16768
rect 256 16736 288 16768
rect 328 16736 360 16768
rect 400 16736 432 16768
rect 472 16736 504 16768
rect 544 16736 576 16768
rect 616 16736 648 16768
rect 688 16736 720 16768
rect 760 16736 792 16768
rect 832 16736 864 16768
rect 904 16736 936 16768
rect 976 16736 1008 16768
rect 1048 16736 1080 16768
rect 1120 16736 1152 16768
rect 1192 16736 1224 16768
rect 1264 16736 1296 16768
rect 1336 16736 1368 16768
rect 1408 16736 1440 16768
rect 1480 16736 1512 16768
rect 1552 16736 1584 16768
rect 1624 16736 1656 16768
rect 1696 16736 1728 16768
rect 1768 16736 1800 16768
rect 1840 16736 1872 16768
rect 1912 16736 1944 16768
rect 1984 16736 2016 16768
rect 2056 16736 2088 16768
rect 2128 16736 2160 16768
rect 2200 16736 2232 16768
rect 2272 16736 2304 16768
rect 2344 16736 2376 16768
rect 2416 16736 2448 16768
rect 2488 16736 2520 16768
rect 2560 16736 2592 16768
rect 2632 16736 2664 16768
rect 2704 16736 2736 16768
rect 2776 16736 2808 16768
rect 2848 16736 2880 16768
rect 2920 16736 2952 16768
rect 2992 16736 3024 16768
rect 3064 16736 3096 16768
rect 3136 16736 3168 16768
rect 3208 16736 3240 16768
rect 3280 16736 3312 16768
rect 3352 16736 3384 16768
rect 3424 16736 3456 16768
rect 3496 16736 3528 16768
rect 3568 16736 3600 16768
rect 3640 16736 3672 16768
rect 3712 16736 3744 16768
rect 3784 16736 3816 16768
rect 3856 16736 3888 16768
rect 112 16664 144 16696
rect 184 16664 216 16696
rect 256 16664 288 16696
rect 328 16664 360 16696
rect 400 16664 432 16696
rect 472 16664 504 16696
rect 544 16664 576 16696
rect 616 16664 648 16696
rect 688 16664 720 16696
rect 760 16664 792 16696
rect 832 16664 864 16696
rect 904 16664 936 16696
rect 976 16664 1008 16696
rect 1048 16664 1080 16696
rect 1120 16664 1152 16696
rect 1192 16664 1224 16696
rect 1264 16664 1296 16696
rect 1336 16664 1368 16696
rect 1408 16664 1440 16696
rect 1480 16664 1512 16696
rect 1552 16664 1584 16696
rect 1624 16664 1656 16696
rect 1696 16664 1728 16696
rect 1768 16664 1800 16696
rect 1840 16664 1872 16696
rect 1912 16664 1944 16696
rect 1984 16664 2016 16696
rect 2056 16664 2088 16696
rect 2128 16664 2160 16696
rect 2200 16664 2232 16696
rect 2272 16664 2304 16696
rect 2344 16664 2376 16696
rect 2416 16664 2448 16696
rect 2488 16664 2520 16696
rect 2560 16664 2592 16696
rect 2632 16664 2664 16696
rect 2704 16664 2736 16696
rect 2776 16664 2808 16696
rect 2848 16664 2880 16696
rect 2920 16664 2952 16696
rect 2992 16664 3024 16696
rect 3064 16664 3096 16696
rect 3136 16664 3168 16696
rect 3208 16664 3240 16696
rect 3280 16664 3312 16696
rect 3352 16664 3384 16696
rect 3424 16664 3456 16696
rect 3496 16664 3528 16696
rect 3568 16664 3600 16696
rect 3640 16664 3672 16696
rect 3712 16664 3744 16696
rect 3784 16664 3816 16696
rect 3856 16664 3888 16696
rect 112 16592 144 16624
rect 184 16592 216 16624
rect 256 16592 288 16624
rect 328 16592 360 16624
rect 400 16592 432 16624
rect 472 16592 504 16624
rect 544 16592 576 16624
rect 616 16592 648 16624
rect 688 16592 720 16624
rect 760 16592 792 16624
rect 832 16592 864 16624
rect 904 16592 936 16624
rect 976 16592 1008 16624
rect 1048 16592 1080 16624
rect 1120 16592 1152 16624
rect 1192 16592 1224 16624
rect 1264 16592 1296 16624
rect 1336 16592 1368 16624
rect 1408 16592 1440 16624
rect 1480 16592 1512 16624
rect 1552 16592 1584 16624
rect 1624 16592 1656 16624
rect 1696 16592 1728 16624
rect 1768 16592 1800 16624
rect 1840 16592 1872 16624
rect 1912 16592 1944 16624
rect 1984 16592 2016 16624
rect 2056 16592 2088 16624
rect 2128 16592 2160 16624
rect 2200 16592 2232 16624
rect 2272 16592 2304 16624
rect 2344 16592 2376 16624
rect 2416 16592 2448 16624
rect 2488 16592 2520 16624
rect 2560 16592 2592 16624
rect 2632 16592 2664 16624
rect 2704 16592 2736 16624
rect 2776 16592 2808 16624
rect 2848 16592 2880 16624
rect 2920 16592 2952 16624
rect 2992 16592 3024 16624
rect 3064 16592 3096 16624
rect 3136 16592 3168 16624
rect 3208 16592 3240 16624
rect 3280 16592 3312 16624
rect 3352 16592 3384 16624
rect 3424 16592 3456 16624
rect 3496 16592 3528 16624
rect 3568 16592 3600 16624
rect 3640 16592 3672 16624
rect 3712 16592 3744 16624
rect 3784 16592 3816 16624
rect 3856 16592 3888 16624
rect 112 16520 144 16552
rect 184 16520 216 16552
rect 256 16520 288 16552
rect 328 16520 360 16552
rect 400 16520 432 16552
rect 472 16520 504 16552
rect 544 16520 576 16552
rect 616 16520 648 16552
rect 688 16520 720 16552
rect 760 16520 792 16552
rect 832 16520 864 16552
rect 904 16520 936 16552
rect 976 16520 1008 16552
rect 1048 16520 1080 16552
rect 1120 16520 1152 16552
rect 1192 16520 1224 16552
rect 1264 16520 1296 16552
rect 1336 16520 1368 16552
rect 1408 16520 1440 16552
rect 1480 16520 1512 16552
rect 1552 16520 1584 16552
rect 1624 16520 1656 16552
rect 1696 16520 1728 16552
rect 1768 16520 1800 16552
rect 1840 16520 1872 16552
rect 1912 16520 1944 16552
rect 1984 16520 2016 16552
rect 2056 16520 2088 16552
rect 2128 16520 2160 16552
rect 2200 16520 2232 16552
rect 2272 16520 2304 16552
rect 2344 16520 2376 16552
rect 2416 16520 2448 16552
rect 2488 16520 2520 16552
rect 2560 16520 2592 16552
rect 2632 16520 2664 16552
rect 2704 16520 2736 16552
rect 2776 16520 2808 16552
rect 2848 16520 2880 16552
rect 2920 16520 2952 16552
rect 2992 16520 3024 16552
rect 3064 16520 3096 16552
rect 3136 16520 3168 16552
rect 3208 16520 3240 16552
rect 3280 16520 3312 16552
rect 3352 16520 3384 16552
rect 3424 16520 3456 16552
rect 3496 16520 3528 16552
rect 3568 16520 3600 16552
rect 3640 16520 3672 16552
rect 3712 16520 3744 16552
rect 3784 16520 3816 16552
rect 3856 16520 3888 16552
rect 112 16448 144 16480
rect 184 16448 216 16480
rect 256 16448 288 16480
rect 328 16448 360 16480
rect 400 16448 432 16480
rect 472 16448 504 16480
rect 544 16448 576 16480
rect 616 16448 648 16480
rect 688 16448 720 16480
rect 760 16448 792 16480
rect 832 16448 864 16480
rect 904 16448 936 16480
rect 976 16448 1008 16480
rect 1048 16448 1080 16480
rect 1120 16448 1152 16480
rect 1192 16448 1224 16480
rect 1264 16448 1296 16480
rect 1336 16448 1368 16480
rect 1408 16448 1440 16480
rect 1480 16448 1512 16480
rect 1552 16448 1584 16480
rect 1624 16448 1656 16480
rect 1696 16448 1728 16480
rect 1768 16448 1800 16480
rect 1840 16448 1872 16480
rect 1912 16448 1944 16480
rect 1984 16448 2016 16480
rect 2056 16448 2088 16480
rect 2128 16448 2160 16480
rect 2200 16448 2232 16480
rect 2272 16448 2304 16480
rect 2344 16448 2376 16480
rect 2416 16448 2448 16480
rect 2488 16448 2520 16480
rect 2560 16448 2592 16480
rect 2632 16448 2664 16480
rect 2704 16448 2736 16480
rect 2776 16448 2808 16480
rect 2848 16448 2880 16480
rect 2920 16448 2952 16480
rect 2992 16448 3024 16480
rect 3064 16448 3096 16480
rect 3136 16448 3168 16480
rect 3208 16448 3240 16480
rect 3280 16448 3312 16480
rect 3352 16448 3384 16480
rect 3424 16448 3456 16480
rect 3496 16448 3528 16480
rect 3568 16448 3600 16480
rect 3640 16448 3672 16480
rect 3712 16448 3744 16480
rect 3784 16448 3816 16480
rect 3856 16448 3888 16480
rect 112 16376 144 16408
rect 184 16376 216 16408
rect 256 16376 288 16408
rect 328 16376 360 16408
rect 400 16376 432 16408
rect 472 16376 504 16408
rect 544 16376 576 16408
rect 616 16376 648 16408
rect 688 16376 720 16408
rect 760 16376 792 16408
rect 832 16376 864 16408
rect 904 16376 936 16408
rect 976 16376 1008 16408
rect 1048 16376 1080 16408
rect 1120 16376 1152 16408
rect 1192 16376 1224 16408
rect 1264 16376 1296 16408
rect 1336 16376 1368 16408
rect 1408 16376 1440 16408
rect 1480 16376 1512 16408
rect 1552 16376 1584 16408
rect 1624 16376 1656 16408
rect 1696 16376 1728 16408
rect 1768 16376 1800 16408
rect 1840 16376 1872 16408
rect 1912 16376 1944 16408
rect 1984 16376 2016 16408
rect 2056 16376 2088 16408
rect 2128 16376 2160 16408
rect 2200 16376 2232 16408
rect 2272 16376 2304 16408
rect 2344 16376 2376 16408
rect 2416 16376 2448 16408
rect 2488 16376 2520 16408
rect 2560 16376 2592 16408
rect 2632 16376 2664 16408
rect 2704 16376 2736 16408
rect 2776 16376 2808 16408
rect 2848 16376 2880 16408
rect 2920 16376 2952 16408
rect 2992 16376 3024 16408
rect 3064 16376 3096 16408
rect 3136 16376 3168 16408
rect 3208 16376 3240 16408
rect 3280 16376 3312 16408
rect 3352 16376 3384 16408
rect 3424 16376 3456 16408
rect 3496 16376 3528 16408
rect 3568 16376 3600 16408
rect 3640 16376 3672 16408
rect 3712 16376 3744 16408
rect 3784 16376 3816 16408
rect 3856 16376 3888 16408
rect 112 16304 144 16336
rect 184 16304 216 16336
rect 256 16304 288 16336
rect 328 16304 360 16336
rect 400 16304 432 16336
rect 472 16304 504 16336
rect 544 16304 576 16336
rect 616 16304 648 16336
rect 688 16304 720 16336
rect 760 16304 792 16336
rect 832 16304 864 16336
rect 904 16304 936 16336
rect 976 16304 1008 16336
rect 1048 16304 1080 16336
rect 1120 16304 1152 16336
rect 1192 16304 1224 16336
rect 1264 16304 1296 16336
rect 1336 16304 1368 16336
rect 1408 16304 1440 16336
rect 1480 16304 1512 16336
rect 1552 16304 1584 16336
rect 1624 16304 1656 16336
rect 1696 16304 1728 16336
rect 1768 16304 1800 16336
rect 1840 16304 1872 16336
rect 1912 16304 1944 16336
rect 1984 16304 2016 16336
rect 2056 16304 2088 16336
rect 2128 16304 2160 16336
rect 2200 16304 2232 16336
rect 2272 16304 2304 16336
rect 2344 16304 2376 16336
rect 2416 16304 2448 16336
rect 2488 16304 2520 16336
rect 2560 16304 2592 16336
rect 2632 16304 2664 16336
rect 2704 16304 2736 16336
rect 2776 16304 2808 16336
rect 2848 16304 2880 16336
rect 2920 16304 2952 16336
rect 2992 16304 3024 16336
rect 3064 16304 3096 16336
rect 3136 16304 3168 16336
rect 3208 16304 3240 16336
rect 3280 16304 3312 16336
rect 3352 16304 3384 16336
rect 3424 16304 3456 16336
rect 3496 16304 3528 16336
rect 3568 16304 3600 16336
rect 3640 16304 3672 16336
rect 3712 16304 3744 16336
rect 3784 16304 3816 16336
rect 3856 16304 3888 16336
rect 112 16232 144 16264
rect 184 16232 216 16264
rect 256 16232 288 16264
rect 328 16232 360 16264
rect 400 16232 432 16264
rect 472 16232 504 16264
rect 544 16232 576 16264
rect 616 16232 648 16264
rect 688 16232 720 16264
rect 760 16232 792 16264
rect 832 16232 864 16264
rect 904 16232 936 16264
rect 976 16232 1008 16264
rect 1048 16232 1080 16264
rect 1120 16232 1152 16264
rect 1192 16232 1224 16264
rect 1264 16232 1296 16264
rect 1336 16232 1368 16264
rect 1408 16232 1440 16264
rect 1480 16232 1512 16264
rect 1552 16232 1584 16264
rect 1624 16232 1656 16264
rect 1696 16232 1728 16264
rect 1768 16232 1800 16264
rect 1840 16232 1872 16264
rect 1912 16232 1944 16264
rect 1984 16232 2016 16264
rect 2056 16232 2088 16264
rect 2128 16232 2160 16264
rect 2200 16232 2232 16264
rect 2272 16232 2304 16264
rect 2344 16232 2376 16264
rect 2416 16232 2448 16264
rect 2488 16232 2520 16264
rect 2560 16232 2592 16264
rect 2632 16232 2664 16264
rect 2704 16232 2736 16264
rect 2776 16232 2808 16264
rect 2848 16232 2880 16264
rect 2920 16232 2952 16264
rect 2992 16232 3024 16264
rect 3064 16232 3096 16264
rect 3136 16232 3168 16264
rect 3208 16232 3240 16264
rect 3280 16232 3312 16264
rect 3352 16232 3384 16264
rect 3424 16232 3456 16264
rect 3496 16232 3528 16264
rect 3568 16232 3600 16264
rect 3640 16232 3672 16264
rect 3712 16232 3744 16264
rect 3784 16232 3816 16264
rect 3856 16232 3888 16264
rect 112 16160 144 16192
rect 184 16160 216 16192
rect 256 16160 288 16192
rect 328 16160 360 16192
rect 400 16160 432 16192
rect 472 16160 504 16192
rect 544 16160 576 16192
rect 616 16160 648 16192
rect 688 16160 720 16192
rect 760 16160 792 16192
rect 832 16160 864 16192
rect 904 16160 936 16192
rect 976 16160 1008 16192
rect 1048 16160 1080 16192
rect 1120 16160 1152 16192
rect 1192 16160 1224 16192
rect 1264 16160 1296 16192
rect 1336 16160 1368 16192
rect 1408 16160 1440 16192
rect 1480 16160 1512 16192
rect 1552 16160 1584 16192
rect 1624 16160 1656 16192
rect 1696 16160 1728 16192
rect 1768 16160 1800 16192
rect 1840 16160 1872 16192
rect 1912 16160 1944 16192
rect 1984 16160 2016 16192
rect 2056 16160 2088 16192
rect 2128 16160 2160 16192
rect 2200 16160 2232 16192
rect 2272 16160 2304 16192
rect 2344 16160 2376 16192
rect 2416 16160 2448 16192
rect 2488 16160 2520 16192
rect 2560 16160 2592 16192
rect 2632 16160 2664 16192
rect 2704 16160 2736 16192
rect 2776 16160 2808 16192
rect 2848 16160 2880 16192
rect 2920 16160 2952 16192
rect 2992 16160 3024 16192
rect 3064 16160 3096 16192
rect 3136 16160 3168 16192
rect 3208 16160 3240 16192
rect 3280 16160 3312 16192
rect 3352 16160 3384 16192
rect 3424 16160 3456 16192
rect 3496 16160 3528 16192
rect 3568 16160 3600 16192
rect 3640 16160 3672 16192
rect 3712 16160 3744 16192
rect 3784 16160 3816 16192
rect 3856 16160 3888 16192
rect 112 16088 144 16120
rect 184 16088 216 16120
rect 256 16088 288 16120
rect 328 16088 360 16120
rect 400 16088 432 16120
rect 472 16088 504 16120
rect 544 16088 576 16120
rect 616 16088 648 16120
rect 688 16088 720 16120
rect 760 16088 792 16120
rect 832 16088 864 16120
rect 904 16088 936 16120
rect 976 16088 1008 16120
rect 1048 16088 1080 16120
rect 1120 16088 1152 16120
rect 1192 16088 1224 16120
rect 1264 16088 1296 16120
rect 1336 16088 1368 16120
rect 1408 16088 1440 16120
rect 1480 16088 1512 16120
rect 1552 16088 1584 16120
rect 1624 16088 1656 16120
rect 1696 16088 1728 16120
rect 1768 16088 1800 16120
rect 1840 16088 1872 16120
rect 1912 16088 1944 16120
rect 1984 16088 2016 16120
rect 2056 16088 2088 16120
rect 2128 16088 2160 16120
rect 2200 16088 2232 16120
rect 2272 16088 2304 16120
rect 2344 16088 2376 16120
rect 2416 16088 2448 16120
rect 2488 16088 2520 16120
rect 2560 16088 2592 16120
rect 2632 16088 2664 16120
rect 2704 16088 2736 16120
rect 2776 16088 2808 16120
rect 2848 16088 2880 16120
rect 2920 16088 2952 16120
rect 2992 16088 3024 16120
rect 3064 16088 3096 16120
rect 3136 16088 3168 16120
rect 3208 16088 3240 16120
rect 3280 16088 3312 16120
rect 3352 16088 3384 16120
rect 3424 16088 3456 16120
rect 3496 16088 3528 16120
rect 3568 16088 3600 16120
rect 3640 16088 3672 16120
rect 3712 16088 3744 16120
rect 3784 16088 3816 16120
rect 3856 16088 3888 16120
rect 112 16016 144 16048
rect 184 16016 216 16048
rect 256 16016 288 16048
rect 328 16016 360 16048
rect 400 16016 432 16048
rect 472 16016 504 16048
rect 544 16016 576 16048
rect 616 16016 648 16048
rect 688 16016 720 16048
rect 760 16016 792 16048
rect 832 16016 864 16048
rect 904 16016 936 16048
rect 976 16016 1008 16048
rect 1048 16016 1080 16048
rect 1120 16016 1152 16048
rect 1192 16016 1224 16048
rect 1264 16016 1296 16048
rect 1336 16016 1368 16048
rect 1408 16016 1440 16048
rect 1480 16016 1512 16048
rect 1552 16016 1584 16048
rect 1624 16016 1656 16048
rect 1696 16016 1728 16048
rect 1768 16016 1800 16048
rect 1840 16016 1872 16048
rect 1912 16016 1944 16048
rect 1984 16016 2016 16048
rect 2056 16016 2088 16048
rect 2128 16016 2160 16048
rect 2200 16016 2232 16048
rect 2272 16016 2304 16048
rect 2344 16016 2376 16048
rect 2416 16016 2448 16048
rect 2488 16016 2520 16048
rect 2560 16016 2592 16048
rect 2632 16016 2664 16048
rect 2704 16016 2736 16048
rect 2776 16016 2808 16048
rect 2848 16016 2880 16048
rect 2920 16016 2952 16048
rect 2992 16016 3024 16048
rect 3064 16016 3096 16048
rect 3136 16016 3168 16048
rect 3208 16016 3240 16048
rect 3280 16016 3312 16048
rect 3352 16016 3384 16048
rect 3424 16016 3456 16048
rect 3496 16016 3528 16048
rect 3568 16016 3600 16048
rect 3640 16016 3672 16048
rect 3712 16016 3744 16048
rect 3784 16016 3816 16048
rect 3856 16016 3888 16048
rect 112 15944 144 15976
rect 184 15944 216 15976
rect 256 15944 288 15976
rect 328 15944 360 15976
rect 400 15944 432 15976
rect 472 15944 504 15976
rect 544 15944 576 15976
rect 616 15944 648 15976
rect 688 15944 720 15976
rect 760 15944 792 15976
rect 832 15944 864 15976
rect 904 15944 936 15976
rect 976 15944 1008 15976
rect 1048 15944 1080 15976
rect 1120 15944 1152 15976
rect 1192 15944 1224 15976
rect 1264 15944 1296 15976
rect 1336 15944 1368 15976
rect 1408 15944 1440 15976
rect 1480 15944 1512 15976
rect 1552 15944 1584 15976
rect 1624 15944 1656 15976
rect 1696 15944 1728 15976
rect 1768 15944 1800 15976
rect 1840 15944 1872 15976
rect 1912 15944 1944 15976
rect 1984 15944 2016 15976
rect 2056 15944 2088 15976
rect 2128 15944 2160 15976
rect 2200 15944 2232 15976
rect 2272 15944 2304 15976
rect 2344 15944 2376 15976
rect 2416 15944 2448 15976
rect 2488 15944 2520 15976
rect 2560 15944 2592 15976
rect 2632 15944 2664 15976
rect 2704 15944 2736 15976
rect 2776 15944 2808 15976
rect 2848 15944 2880 15976
rect 2920 15944 2952 15976
rect 2992 15944 3024 15976
rect 3064 15944 3096 15976
rect 3136 15944 3168 15976
rect 3208 15944 3240 15976
rect 3280 15944 3312 15976
rect 3352 15944 3384 15976
rect 3424 15944 3456 15976
rect 3496 15944 3528 15976
rect 3568 15944 3600 15976
rect 3640 15944 3672 15976
rect 3712 15944 3744 15976
rect 3784 15944 3816 15976
rect 3856 15944 3888 15976
rect 112 15872 144 15904
rect 184 15872 216 15904
rect 256 15872 288 15904
rect 328 15872 360 15904
rect 400 15872 432 15904
rect 472 15872 504 15904
rect 544 15872 576 15904
rect 616 15872 648 15904
rect 688 15872 720 15904
rect 760 15872 792 15904
rect 832 15872 864 15904
rect 904 15872 936 15904
rect 976 15872 1008 15904
rect 1048 15872 1080 15904
rect 1120 15872 1152 15904
rect 1192 15872 1224 15904
rect 1264 15872 1296 15904
rect 1336 15872 1368 15904
rect 1408 15872 1440 15904
rect 1480 15872 1512 15904
rect 1552 15872 1584 15904
rect 1624 15872 1656 15904
rect 1696 15872 1728 15904
rect 1768 15872 1800 15904
rect 1840 15872 1872 15904
rect 1912 15872 1944 15904
rect 1984 15872 2016 15904
rect 2056 15872 2088 15904
rect 2128 15872 2160 15904
rect 2200 15872 2232 15904
rect 2272 15872 2304 15904
rect 2344 15872 2376 15904
rect 2416 15872 2448 15904
rect 2488 15872 2520 15904
rect 2560 15872 2592 15904
rect 2632 15872 2664 15904
rect 2704 15872 2736 15904
rect 2776 15872 2808 15904
rect 2848 15872 2880 15904
rect 2920 15872 2952 15904
rect 2992 15872 3024 15904
rect 3064 15872 3096 15904
rect 3136 15872 3168 15904
rect 3208 15872 3240 15904
rect 3280 15872 3312 15904
rect 3352 15872 3384 15904
rect 3424 15872 3456 15904
rect 3496 15872 3528 15904
rect 3568 15872 3600 15904
rect 3640 15872 3672 15904
rect 3712 15872 3744 15904
rect 3784 15872 3816 15904
rect 3856 15872 3888 15904
rect 112 15800 144 15832
rect 184 15800 216 15832
rect 256 15800 288 15832
rect 328 15800 360 15832
rect 400 15800 432 15832
rect 472 15800 504 15832
rect 544 15800 576 15832
rect 616 15800 648 15832
rect 688 15800 720 15832
rect 760 15800 792 15832
rect 832 15800 864 15832
rect 904 15800 936 15832
rect 976 15800 1008 15832
rect 1048 15800 1080 15832
rect 1120 15800 1152 15832
rect 1192 15800 1224 15832
rect 1264 15800 1296 15832
rect 1336 15800 1368 15832
rect 1408 15800 1440 15832
rect 1480 15800 1512 15832
rect 1552 15800 1584 15832
rect 1624 15800 1656 15832
rect 1696 15800 1728 15832
rect 1768 15800 1800 15832
rect 1840 15800 1872 15832
rect 1912 15800 1944 15832
rect 1984 15800 2016 15832
rect 2056 15800 2088 15832
rect 2128 15800 2160 15832
rect 2200 15800 2232 15832
rect 2272 15800 2304 15832
rect 2344 15800 2376 15832
rect 2416 15800 2448 15832
rect 2488 15800 2520 15832
rect 2560 15800 2592 15832
rect 2632 15800 2664 15832
rect 2704 15800 2736 15832
rect 2776 15800 2808 15832
rect 2848 15800 2880 15832
rect 2920 15800 2952 15832
rect 2992 15800 3024 15832
rect 3064 15800 3096 15832
rect 3136 15800 3168 15832
rect 3208 15800 3240 15832
rect 3280 15800 3312 15832
rect 3352 15800 3384 15832
rect 3424 15800 3456 15832
rect 3496 15800 3528 15832
rect 3568 15800 3600 15832
rect 3640 15800 3672 15832
rect 3712 15800 3744 15832
rect 3784 15800 3816 15832
rect 3856 15800 3888 15832
rect 112 15728 144 15760
rect 184 15728 216 15760
rect 256 15728 288 15760
rect 328 15728 360 15760
rect 400 15728 432 15760
rect 472 15728 504 15760
rect 544 15728 576 15760
rect 616 15728 648 15760
rect 688 15728 720 15760
rect 760 15728 792 15760
rect 832 15728 864 15760
rect 904 15728 936 15760
rect 976 15728 1008 15760
rect 1048 15728 1080 15760
rect 1120 15728 1152 15760
rect 1192 15728 1224 15760
rect 1264 15728 1296 15760
rect 1336 15728 1368 15760
rect 1408 15728 1440 15760
rect 1480 15728 1512 15760
rect 1552 15728 1584 15760
rect 1624 15728 1656 15760
rect 1696 15728 1728 15760
rect 1768 15728 1800 15760
rect 1840 15728 1872 15760
rect 1912 15728 1944 15760
rect 1984 15728 2016 15760
rect 2056 15728 2088 15760
rect 2128 15728 2160 15760
rect 2200 15728 2232 15760
rect 2272 15728 2304 15760
rect 2344 15728 2376 15760
rect 2416 15728 2448 15760
rect 2488 15728 2520 15760
rect 2560 15728 2592 15760
rect 2632 15728 2664 15760
rect 2704 15728 2736 15760
rect 2776 15728 2808 15760
rect 2848 15728 2880 15760
rect 2920 15728 2952 15760
rect 2992 15728 3024 15760
rect 3064 15728 3096 15760
rect 3136 15728 3168 15760
rect 3208 15728 3240 15760
rect 3280 15728 3312 15760
rect 3352 15728 3384 15760
rect 3424 15728 3456 15760
rect 3496 15728 3528 15760
rect 3568 15728 3600 15760
rect 3640 15728 3672 15760
rect 3712 15728 3744 15760
rect 3784 15728 3816 15760
rect 3856 15728 3888 15760
rect 112 15656 144 15688
rect 184 15656 216 15688
rect 256 15656 288 15688
rect 328 15656 360 15688
rect 400 15656 432 15688
rect 472 15656 504 15688
rect 544 15656 576 15688
rect 616 15656 648 15688
rect 688 15656 720 15688
rect 760 15656 792 15688
rect 832 15656 864 15688
rect 904 15656 936 15688
rect 976 15656 1008 15688
rect 1048 15656 1080 15688
rect 1120 15656 1152 15688
rect 1192 15656 1224 15688
rect 1264 15656 1296 15688
rect 1336 15656 1368 15688
rect 1408 15656 1440 15688
rect 1480 15656 1512 15688
rect 1552 15656 1584 15688
rect 1624 15656 1656 15688
rect 1696 15656 1728 15688
rect 1768 15656 1800 15688
rect 1840 15656 1872 15688
rect 1912 15656 1944 15688
rect 1984 15656 2016 15688
rect 2056 15656 2088 15688
rect 2128 15656 2160 15688
rect 2200 15656 2232 15688
rect 2272 15656 2304 15688
rect 2344 15656 2376 15688
rect 2416 15656 2448 15688
rect 2488 15656 2520 15688
rect 2560 15656 2592 15688
rect 2632 15656 2664 15688
rect 2704 15656 2736 15688
rect 2776 15656 2808 15688
rect 2848 15656 2880 15688
rect 2920 15656 2952 15688
rect 2992 15656 3024 15688
rect 3064 15656 3096 15688
rect 3136 15656 3168 15688
rect 3208 15656 3240 15688
rect 3280 15656 3312 15688
rect 3352 15656 3384 15688
rect 3424 15656 3456 15688
rect 3496 15656 3528 15688
rect 3568 15656 3600 15688
rect 3640 15656 3672 15688
rect 3712 15656 3744 15688
rect 3784 15656 3816 15688
rect 3856 15656 3888 15688
rect 112 15584 144 15616
rect 184 15584 216 15616
rect 256 15584 288 15616
rect 328 15584 360 15616
rect 400 15584 432 15616
rect 472 15584 504 15616
rect 544 15584 576 15616
rect 616 15584 648 15616
rect 688 15584 720 15616
rect 760 15584 792 15616
rect 832 15584 864 15616
rect 904 15584 936 15616
rect 976 15584 1008 15616
rect 1048 15584 1080 15616
rect 1120 15584 1152 15616
rect 1192 15584 1224 15616
rect 1264 15584 1296 15616
rect 1336 15584 1368 15616
rect 1408 15584 1440 15616
rect 1480 15584 1512 15616
rect 1552 15584 1584 15616
rect 1624 15584 1656 15616
rect 1696 15584 1728 15616
rect 1768 15584 1800 15616
rect 1840 15584 1872 15616
rect 1912 15584 1944 15616
rect 1984 15584 2016 15616
rect 2056 15584 2088 15616
rect 2128 15584 2160 15616
rect 2200 15584 2232 15616
rect 2272 15584 2304 15616
rect 2344 15584 2376 15616
rect 2416 15584 2448 15616
rect 2488 15584 2520 15616
rect 2560 15584 2592 15616
rect 2632 15584 2664 15616
rect 2704 15584 2736 15616
rect 2776 15584 2808 15616
rect 2848 15584 2880 15616
rect 2920 15584 2952 15616
rect 2992 15584 3024 15616
rect 3064 15584 3096 15616
rect 3136 15584 3168 15616
rect 3208 15584 3240 15616
rect 3280 15584 3312 15616
rect 3352 15584 3384 15616
rect 3424 15584 3456 15616
rect 3496 15584 3528 15616
rect 3568 15584 3600 15616
rect 3640 15584 3672 15616
rect 3712 15584 3744 15616
rect 3784 15584 3816 15616
rect 3856 15584 3888 15616
rect 112 15512 144 15544
rect 184 15512 216 15544
rect 256 15512 288 15544
rect 328 15512 360 15544
rect 400 15512 432 15544
rect 472 15512 504 15544
rect 544 15512 576 15544
rect 616 15512 648 15544
rect 688 15512 720 15544
rect 760 15512 792 15544
rect 832 15512 864 15544
rect 904 15512 936 15544
rect 976 15512 1008 15544
rect 1048 15512 1080 15544
rect 1120 15512 1152 15544
rect 1192 15512 1224 15544
rect 1264 15512 1296 15544
rect 1336 15512 1368 15544
rect 1408 15512 1440 15544
rect 1480 15512 1512 15544
rect 1552 15512 1584 15544
rect 1624 15512 1656 15544
rect 1696 15512 1728 15544
rect 1768 15512 1800 15544
rect 1840 15512 1872 15544
rect 1912 15512 1944 15544
rect 1984 15512 2016 15544
rect 2056 15512 2088 15544
rect 2128 15512 2160 15544
rect 2200 15512 2232 15544
rect 2272 15512 2304 15544
rect 2344 15512 2376 15544
rect 2416 15512 2448 15544
rect 2488 15512 2520 15544
rect 2560 15512 2592 15544
rect 2632 15512 2664 15544
rect 2704 15512 2736 15544
rect 2776 15512 2808 15544
rect 2848 15512 2880 15544
rect 2920 15512 2952 15544
rect 2992 15512 3024 15544
rect 3064 15512 3096 15544
rect 3136 15512 3168 15544
rect 3208 15512 3240 15544
rect 3280 15512 3312 15544
rect 3352 15512 3384 15544
rect 3424 15512 3456 15544
rect 3496 15512 3528 15544
rect 3568 15512 3600 15544
rect 3640 15512 3672 15544
rect 3712 15512 3744 15544
rect 3784 15512 3816 15544
rect 3856 15512 3888 15544
rect 112 15440 144 15472
rect 184 15440 216 15472
rect 256 15440 288 15472
rect 328 15440 360 15472
rect 400 15440 432 15472
rect 472 15440 504 15472
rect 544 15440 576 15472
rect 616 15440 648 15472
rect 688 15440 720 15472
rect 760 15440 792 15472
rect 832 15440 864 15472
rect 904 15440 936 15472
rect 976 15440 1008 15472
rect 1048 15440 1080 15472
rect 1120 15440 1152 15472
rect 1192 15440 1224 15472
rect 1264 15440 1296 15472
rect 1336 15440 1368 15472
rect 1408 15440 1440 15472
rect 1480 15440 1512 15472
rect 1552 15440 1584 15472
rect 1624 15440 1656 15472
rect 1696 15440 1728 15472
rect 1768 15440 1800 15472
rect 1840 15440 1872 15472
rect 1912 15440 1944 15472
rect 1984 15440 2016 15472
rect 2056 15440 2088 15472
rect 2128 15440 2160 15472
rect 2200 15440 2232 15472
rect 2272 15440 2304 15472
rect 2344 15440 2376 15472
rect 2416 15440 2448 15472
rect 2488 15440 2520 15472
rect 2560 15440 2592 15472
rect 2632 15440 2664 15472
rect 2704 15440 2736 15472
rect 2776 15440 2808 15472
rect 2848 15440 2880 15472
rect 2920 15440 2952 15472
rect 2992 15440 3024 15472
rect 3064 15440 3096 15472
rect 3136 15440 3168 15472
rect 3208 15440 3240 15472
rect 3280 15440 3312 15472
rect 3352 15440 3384 15472
rect 3424 15440 3456 15472
rect 3496 15440 3528 15472
rect 3568 15440 3600 15472
rect 3640 15440 3672 15472
rect 3712 15440 3744 15472
rect 3784 15440 3816 15472
rect 3856 15440 3888 15472
rect 112 15368 144 15400
rect 184 15368 216 15400
rect 256 15368 288 15400
rect 328 15368 360 15400
rect 400 15368 432 15400
rect 472 15368 504 15400
rect 544 15368 576 15400
rect 616 15368 648 15400
rect 688 15368 720 15400
rect 760 15368 792 15400
rect 832 15368 864 15400
rect 904 15368 936 15400
rect 976 15368 1008 15400
rect 1048 15368 1080 15400
rect 1120 15368 1152 15400
rect 1192 15368 1224 15400
rect 1264 15368 1296 15400
rect 1336 15368 1368 15400
rect 1408 15368 1440 15400
rect 1480 15368 1512 15400
rect 1552 15368 1584 15400
rect 1624 15368 1656 15400
rect 1696 15368 1728 15400
rect 1768 15368 1800 15400
rect 1840 15368 1872 15400
rect 1912 15368 1944 15400
rect 1984 15368 2016 15400
rect 2056 15368 2088 15400
rect 2128 15368 2160 15400
rect 2200 15368 2232 15400
rect 2272 15368 2304 15400
rect 2344 15368 2376 15400
rect 2416 15368 2448 15400
rect 2488 15368 2520 15400
rect 2560 15368 2592 15400
rect 2632 15368 2664 15400
rect 2704 15368 2736 15400
rect 2776 15368 2808 15400
rect 2848 15368 2880 15400
rect 2920 15368 2952 15400
rect 2992 15368 3024 15400
rect 3064 15368 3096 15400
rect 3136 15368 3168 15400
rect 3208 15368 3240 15400
rect 3280 15368 3312 15400
rect 3352 15368 3384 15400
rect 3424 15368 3456 15400
rect 3496 15368 3528 15400
rect 3568 15368 3600 15400
rect 3640 15368 3672 15400
rect 3712 15368 3744 15400
rect 3784 15368 3816 15400
rect 3856 15368 3888 15400
rect 112 15296 144 15328
rect 184 15296 216 15328
rect 256 15296 288 15328
rect 328 15296 360 15328
rect 400 15296 432 15328
rect 472 15296 504 15328
rect 544 15296 576 15328
rect 616 15296 648 15328
rect 688 15296 720 15328
rect 760 15296 792 15328
rect 832 15296 864 15328
rect 904 15296 936 15328
rect 976 15296 1008 15328
rect 1048 15296 1080 15328
rect 1120 15296 1152 15328
rect 1192 15296 1224 15328
rect 1264 15296 1296 15328
rect 1336 15296 1368 15328
rect 1408 15296 1440 15328
rect 1480 15296 1512 15328
rect 1552 15296 1584 15328
rect 1624 15296 1656 15328
rect 1696 15296 1728 15328
rect 1768 15296 1800 15328
rect 1840 15296 1872 15328
rect 1912 15296 1944 15328
rect 1984 15296 2016 15328
rect 2056 15296 2088 15328
rect 2128 15296 2160 15328
rect 2200 15296 2232 15328
rect 2272 15296 2304 15328
rect 2344 15296 2376 15328
rect 2416 15296 2448 15328
rect 2488 15296 2520 15328
rect 2560 15296 2592 15328
rect 2632 15296 2664 15328
rect 2704 15296 2736 15328
rect 2776 15296 2808 15328
rect 2848 15296 2880 15328
rect 2920 15296 2952 15328
rect 2992 15296 3024 15328
rect 3064 15296 3096 15328
rect 3136 15296 3168 15328
rect 3208 15296 3240 15328
rect 3280 15296 3312 15328
rect 3352 15296 3384 15328
rect 3424 15296 3456 15328
rect 3496 15296 3528 15328
rect 3568 15296 3600 15328
rect 3640 15296 3672 15328
rect 3712 15296 3744 15328
rect 3784 15296 3816 15328
rect 3856 15296 3888 15328
rect 112 15224 144 15256
rect 184 15224 216 15256
rect 256 15224 288 15256
rect 328 15224 360 15256
rect 400 15224 432 15256
rect 472 15224 504 15256
rect 544 15224 576 15256
rect 616 15224 648 15256
rect 688 15224 720 15256
rect 760 15224 792 15256
rect 832 15224 864 15256
rect 904 15224 936 15256
rect 976 15224 1008 15256
rect 1048 15224 1080 15256
rect 1120 15224 1152 15256
rect 1192 15224 1224 15256
rect 1264 15224 1296 15256
rect 1336 15224 1368 15256
rect 1408 15224 1440 15256
rect 1480 15224 1512 15256
rect 1552 15224 1584 15256
rect 1624 15224 1656 15256
rect 1696 15224 1728 15256
rect 1768 15224 1800 15256
rect 1840 15224 1872 15256
rect 1912 15224 1944 15256
rect 1984 15224 2016 15256
rect 2056 15224 2088 15256
rect 2128 15224 2160 15256
rect 2200 15224 2232 15256
rect 2272 15224 2304 15256
rect 2344 15224 2376 15256
rect 2416 15224 2448 15256
rect 2488 15224 2520 15256
rect 2560 15224 2592 15256
rect 2632 15224 2664 15256
rect 2704 15224 2736 15256
rect 2776 15224 2808 15256
rect 2848 15224 2880 15256
rect 2920 15224 2952 15256
rect 2992 15224 3024 15256
rect 3064 15224 3096 15256
rect 3136 15224 3168 15256
rect 3208 15224 3240 15256
rect 3280 15224 3312 15256
rect 3352 15224 3384 15256
rect 3424 15224 3456 15256
rect 3496 15224 3528 15256
rect 3568 15224 3600 15256
rect 3640 15224 3672 15256
rect 3712 15224 3744 15256
rect 3784 15224 3816 15256
rect 3856 15224 3888 15256
rect 112 15152 144 15184
rect 184 15152 216 15184
rect 256 15152 288 15184
rect 328 15152 360 15184
rect 400 15152 432 15184
rect 472 15152 504 15184
rect 544 15152 576 15184
rect 616 15152 648 15184
rect 688 15152 720 15184
rect 760 15152 792 15184
rect 832 15152 864 15184
rect 904 15152 936 15184
rect 976 15152 1008 15184
rect 1048 15152 1080 15184
rect 1120 15152 1152 15184
rect 1192 15152 1224 15184
rect 1264 15152 1296 15184
rect 1336 15152 1368 15184
rect 1408 15152 1440 15184
rect 1480 15152 1512 15184
rect 1552 15152 1584 15184
rect 1624 15152 1656 15184
rect 1696 15152 1728 15184
rect 1768 15152 1800 15184
rect 1840 15152 1872 15184
rect 1912 15152 1944 15184
rect 1984 15152 2016 15184
rect 2056 15152 2088 15184
rect 2128 15152 2160 15184
rect 2200 15152 2232 15184
rect 2272 15152 2304 15184
rect 2344 15152 2376 15184
rect 2416 15152 2448 15184
rect 2488 15152 2520 15184
rect 2560 15152 2592 15184
rect 2632 15152 2664 15184
rect 2704 15152 2736 15184
rect 2776 15152 2808 15184
rect 2848 15152 2880 15184
rect 2920 15152 2952 15184
rect 2992 15152 3024 15184
rect 3064 15152 3096 15184
rect 3136 15152 3168 15184
rect 3208 15152 3240 15184
rect 3280 15152 3312 15184
rect 3352 15152 3384 15184
rect 3424 15152 3456 15184
rect 3496 15152 3528 15184
rect 3568 15152 3600 15184
rect 3640 15152 3672 15184
rect 3712 15152 3744 15184
rect 3784 15152 3816 15184
rect 3856 15152 3888 15184
rect 112 15080 144 15112
rect 184 15080 216 15112
rect 256 15080 288 15112
rect 328 15080 360 15112
rect 400 15080 432 15112
rect 472 15080 504 15112
rect 544 15080 576 15112
rect 616 15080 648 15112
rect 688 15080 720 15112
rect 760 15080 792 15112
rect 832 15080 864 15112
rect 904 15080 936 15112
rect 976 15080 1008 15112
rect 1048 15080 1080 15112
rect 1120 15080 1152 15112
rect 1192 15080 1224 15112
rect 1264 15080 1296 15112
rect 1336 15080 1368 15112
rect 1408 15080 1440 15112
rect 1480 15080 1512 15112
rect 1552 15080 1584 15112
rect 1624 15080 1656 15112
rect 1696 15080 1728 15112
rect 1768 15080 1800 15112
rect 1840 15080 1872 15112
rect 1912 15080 1944 15112
rect 1984 15080 2016 15112
rect 2056 15080 2088 15112
rect 2128 15080 2160 15112
rect 2200 15080 2232 15112
rect 2272 15080 2304 15112
rect 2344 15080 2376 15112
rect 2416 15080 2448 15112
rect 2488 15080 2520 15112
rect 2560 15080 2592 15112
rect 2632 15080 2664 15112
rect 2704 15080 2736 15112
rect 2776 15080 2808 15112
rect 2848 15080 2880 15112
rect 2920 15080 2952 15112
rect 2992 15080 3024 15112
rect 3064 15080 3096 15112
rect 3136 15080 3168 15112
rect 3208 15080 3240 15112
rect 3280 15080 3312 15112
rect 3352 15080 3384 15112
rect 3424 15080 3456 15112
rect 3496 15080 3528 15112
rect 3568 15080 3600 15112
rect 3640 15080 3672 15112
rect 3712 15080 3744 15112
rect 3784 15080 3816 15112
rect 3856 15080 3888 15112
rect 112 15008 144 15040
rect 184 15008 216 15040
rect 256 15008 288 15040
rect 328 15008 360 15040
rect 400 15008 432 15040
rect 472 15008 504 15040
rect 544 15008 576 15040
rect 616 15008 648 15040
rect 688 15008 720 15040
rect 760 15008 792 15040
rect 832 15008 864 15040
rect 904 15008 936 15040
rect 976 15008 1008 15040
rect 1048 15008 1080 15040
rect 1120 15008 1152 15040
rect 1192 15008 1224 15040
rect 1264 15008 1296 15040
rect 1336 15008 1368 15040
rect 1408 15008 1440 15040
rect 1480 15008 1512 15040
rect 1552 15008 1584 15040
rect 1624 15008 1656 15040
rect 1696 15008 1728 15040
rect 1768 15008 1800 15040
rect 1840 15008 1872 15040
rect 1912 15008 1944 15040
rect 1984 15008 2016 15040
rect 2056 15008 2088 15040
rect 2128 15008 2160 15040
rect 2200 15008 2232 15040
rect 2272 15008 2304 15040
rect 2344 15008 2376 15040
rect 2416 15008 2448 15040
rect 2488 15008 2520 15040
rect 2560 15008 2592 15040
rect 2632 15008 2664 15040
rect 2704 15008 2736 15040
rect 2776 15008 2808 15040
rect 2848 15008 2880 15040
rect 2920 15008 2952 15040
rect 2992 15008 3024 15040
rect 3064 15008 3096 15040
rect 3136 15008 3168 15040
rect 3208 15008 3240 15040
rect 3280 15008 3312 15040
rect 3352 15008 3384 15040
rect 3424 15008 3456 15040
rect 3496 15008 3528 15040
rect 3568 15008 3600 15040
rect 3640 15008 3672 15040
rect 3712 15008 3744 15040
rect 3784 15008 3816 15040
rect 3856 15008 3888 15040
rect 112 14936 144 14968
rect 184 14936 216 14968
rect 256 14936 288 14968
rect 328 14936 360 14968
rect 400 14936 432 14968
rect 472 14936 504 14968
rect 544 14936 576 14968
rect 616 14936 648 14968
rect 688 14936 720 14968
rect 760 14936 792 14968
rect 832 14936 864 14968
rect 904 14936 936 14968
rect 976 14936 1008 14968
rect 1048 14936 1080 14968
rect 1120 14936 1152 14968
rect 1192 14936 1224 14968
rect 1264 14936 1296 14968
rect 1336 14936 1368 14968
rect 1408 14936 1440 14968
rect 1480 14936 1512 14968
rect 1552 14936 1584 14968
rect 1624 14936 1656 14968
rect 1696 14936 1728 14968
rect 1768 14936 1800 14968
rect 1840 14936 1872 14968
rect 1912 14936 1944 14968
rect 1984 14936 2016 14968
rect 2056 14936 2088 14968
rect 2128 14936 2160 14968
rect 2200 14936 2232 14968
rect 2272 14936 2304 14968
rect 2344 14936 2376 14968
rect 2416 14936 2448 14968
rect 2488 14936 2520 14968
rect 2560 14936 2592 14968
rect 2632 14936 2664 14968
rect 2704 14936 2736 14968
rect 2776 14936 2808 14968
rect 2848 14936 2880 14968
rect 2920 14936 2952 14968
rect 2992 14936 3024 14968
rect 3064 14936 3096 14968
rect 3136 14936 3168 14968
rect 3208 14936 3240 14968
rect 3280 14936 3312 14968
rect 3352 14936 3384 14968
rect 3424 14936 3456 14968
rect 3496 14936 3528 14968
rect 3568 14936 3600 14968
rect 3640 14936 3672 14968
rect 3712 14936 3744 14968
rect 3784 14936 3816 14968
rect 3856 14936 3888 14968
rect 112 14864 144 14896
rect 184 14864 216 14896
rect 256 14864 288 14896
rect 328 14864 360 14896
rect 400 14864 432 14896
rect 472 14864 504 14896
rect 544 14864 576 14896
rect 616 14864 648 14896
rect 688 14864 720 14896
rect 760 14864 792 14896
rect 832 14864 864 14896
rect 904 14864 936 14896
rect 976 14864 1008 14896
rect 1048 14864 1080 14896
rect 1120 14864 1152 14896
rect 1192 14864 1224 14896
rect 1264 14864 1296 14896
rect 1336 14864 1368 14896
rect 1408 14864 1440 14896
rect 1480 14864 1512 14896
rect 1552 14864 1584 14896
rect 1624 14864 1656 14896
rect 1696 14864 1728 14896
rect 1768 14864 1800 14896
rect 1840 14864 1872 14896
rect 1912 14864 1944 14896
rect 1984 14864 2016 14896
rect 2056 14864 2088 14896
rect 2128 14864 2160 14896
rect 2200 14864 2232 14896
rect 2272 14864 2304 14896
rect 2344 14864 2376 14896
rect 2416 14864 2448 14896
rect 2488 14864 2520 14896
rect 2560 14864 2592 14896
rect 2632 14864 2664 14896
rect 2704 14864 2736 14896
rect 2776 14864 2808 14896
rect 2848 14864 2880 14896
rect 2920 14864 2952 14896
rect 2992 14864 3024 14896
rect 3064 14864 3096 14896
rect 3136 14864 3168 14896
rect 3208 14864 3240 14896
rect 3280 14864 3312 14896
rect 3352 14864 3384 14896
rect 3424 14864 3456 14896
rect 3496 14864 3528 14896
rect 3568 14864 3600 14896
rect 3640 14864 3672 14896
rect 3712 14864 3744 14896
rect 3784 14864 3816 14896
rect 3856 14864 3888 14896
rect 112 14792 144 14824
rect 184 14792 216 14824
rect 256 14792 288 14824
rect 328 14792 360 14824
rect 400 14792 432 14824
rect 472 14792 504 14824
rect 544 14792 576 14824
rect 616 14792 648 14824
rect 688 14792 720 14824
rect 760 14792 792 14824
rect 832 14792 864 14824
rect 904 14792 936 14824
rect 976 14792 1008 14824
rect 1048 14792 1080 14824
rect 1120 14792 1152 14824
rect 1192 14792 1224 14824
rect 1264 14792 1296 14824
rect 1336 14792 1368 14824
rect 1408 14792 1440 14824
rect 1480 14792 1512 14824
rect 1552 14792 1584 14824
rect 1624 14792 1656 14824
rect 1696 14792 1728 14824
rect 1768 14792 1800 14824
rect 1840 14792 1872 14824
rect 1912 14792 1944 14824
rect 1984 14792 2016 14824
rect 2056 14792 2088 14824
rect 2128 14792 2160 14824
rect 2200 14792 2232 14824
rect 2272 14792 2304 14824
rect 2344 14792 2376 14824
rect 2416 14792 2448 14824
rect 2488 14792 2520 14824
rect 2560 14792 2592 14824
rect 2632 14792 2664 14824
rect 2704 14792 2736 14824
rect 2776 14792 2808 14824
rect 2848 14792 2880 14824
rect 2920 14792 2952 14824
rect 2992 14792 3024 14824
rect 3064 14792 3096 14824
rect 3136 14792 3168 14824
rect 3208 14792 3240 14824
rect 3280 14792 3312 14824
rect 3352 14792 3384 14824
rect 3424 14792 3456 14824
rect 3496 14792 3528 14824
rect 3568 14792 3600 14824
rect 3640 14792 3672 14824
rect 3712 14792 3744 14824
rect 3784 14792 3816 14824
rect 3856 14792 3888 14824
rect 112 14720 144 14752
rect 184 14720 216 14752
rect 256 14720 288 14752
rect 328 14720 360 14752
rect 400 14720 432 14752
rect 472 14720 504 14752
rect 544 14720 576 14752
rect 616 14720 648 14752
rect 688 14720 720 14752
rect 760 14720 792 14752
rect 832 14720 864 14752
rect 904 14720 936 14752
rect 976 14720 1008 14752
rect 1048 14720 1080 14752
rect 1120 14720 1152 14752
rect 1192 14720 1224 14752
rect 1264 14720 1296 14752
rect 1336 14720 1368 14752
rect 1408 14720 1440 14752
rect 1480 14720 1512 14752
rect 1552 14720 1584 14752
rect 1624 14720 1656 14752
rect 1696 14720 1728 14752
rect 1768 14720 1800 14752
rect 1840 14720 1872 14752
rect 1912 14720 1944 14752
rect 1984 14720 2016 14752
rect 2056 14720 2088 14752
rect 2128 14720 2160 14752
rect 2200 14720 2232 14752
rect 2272 14720 2304 14752
rect 2344 14720 2376 14752
rect 2416 14720 2448 14752
rect 2488 14720 2520 14752
rect 2560 14720 2592 14752
rect 2632 14720 2664 14752
rect 2704 14720 2736 14752
rect 2776 14720 2808 14752
rect 2848 14720 2880 14752
rect 2920 14720 2952 14752
rect 2992 14720 3024 14752
rect 3064 14720 3096 14752
rect 3136 14720 3168 14752
rect 3208 14720 3240 14752
rect 3280 14720 3312 14752
rect 3352 14720 3384 14752
rect 3424 14720 3456 14752
rect 3496 14720 3528 14752
rect 3568 14720 3600 14752
rect 3640 14720 3672 14752
rect 3712 14720 3744 14752
rect 3784 14720 3816 14752
rect 3856 14720 3888 14752
rect 112 14648 144 14680
rect 184 14648 216 14680
rect 256 14648 288 14680
rect 328 14648 360 14680
rect 400 14648 432 14680
rect 472 14648 504 14680
rect 544 14648 576 14680
rect 616 14648 648 14680
rect 688 14648 720 14680
rect 760 14648 792 14680
rect 832 14648 864 14680
rect 904 14648 936 14680
rect 976 14648 1008 14680
rect 1048 14648 1080 14680
rect 1120 14648 1152 14680
rect 1192 14648 1224 14680
rect 1264 14648 1296 14680
rect 1336 14648 1368 14680
rect 1408 14648 1440 14680
rect 1480 14648 1512 14680
rect 1552 14648 1584 14680
rect 1624 14648 1656 14680
rect 1696 14648 1728 14680
rect 1768 14648 1800 14680
rect 1840 14648 1872 14680
rect 1912 14648 1944 14680
rect 1984 14648 2016 14680
rect 2056 14648 2088 14680
rect 2128 14648 2160 14680
rect 2200 14648 2232 14680
rect 2272 14648 2304 14680
rect 2344 14648 2376 14680
rect 2416 14648 2448 14680
rect 2488 14648 2520 14680
rect 2560 14648 2592 14680
rect 2632 14648 2664 14680
rect 2704 14648 2736 14680
rect 2776 14648 2808 14680
rect 2848 14648 2880 14680
rect 2920 14648 2952 14680
rect 2992 14648 3024 14680
rect 3064 14648 3096 14680
rect 3136 14648 3168 14680
rect 3208 14648 3240 14680
rect 3280 14648 3312 14680
rect 3352 14648 3384 14680
rect 3424 14648 3456 14680
rect 3496 14648 3528 14680
rect 3568 14648 3600 14680
rect 3640 14648 3672 14680
rect 3712 14648 3744 14680
rect 3784 14648 3816 14680
rect 3856 14648 3888 14680
rect 112 14576 144 14608
rect 184 14576 216 14608
rect 256 14576 288 14608
rect 328 14576 360 14608
rect 400 14576 432 14608
rect 472 14576 504 14608
rect 544 14576 576 14608
rect 616 14576 648 14608
rect 688 14576 720 14608
rect 760 14576 792 14608
rect 832 14576 864 14608
rect 904 14576 936 14608
rect 976 14576 1008 14608
rect 1048 14576 1080 14608
rect 1120 14576 1152 14608
rect 1192 14576 1224 14608
rect 1264 14576 1296 14608
rect 1336 14576 1368 14608
rect 1408 14576 1440 14608
rect 1480 14576 1512 14608
rect 1552 14576 1584 14608
rect 1624 14576 1656 14608
rect 1696 14576 1728 14608
rect 1768 14576 1800 14608
rect 1840 14576 1872 14608
rect 1912 14576 1944 14608
rect 1984 14576 2016 14608
rect 2056 14576 2088 14608
rect 2128 14576 2160 14608
rect 2200 14576 2232 14608
rect 2272 14576 2304 14608
rect 2344 14576 2376 14608
rect 2416 14576 2448 14608
rect 2488 14576 2520 14608
rect 2560 14576 2592 14608
rect 2632 14576 2664 14608
rect 2704 14576 2736 14608
rect 2776 14576 2808 14608
rect 2848 14576 2880 14608
rect 2920 14576 2952 14608
rect 2992 14576 3024 14608
rect 3064 14576 3096 14608
rect 3136 14576 3168 14608
rect 3208 14576 3240 14608
rect 3280 14576 3312 14608
rect 3352 14576 3384 14608
rect 3424 14576 3456 14608
rect 3496 14576 3528 14608
rect 3568 14576 3600 14608
rect 3640 14576 3672 14608
rect 3712 14576 3744 14608
rect 3784 14576 3816 14608
rect 3856 14576 3888 14608
rect 112 14504 144 14536
rect 184 14504 216 14536
rect 256 14504 288 14536
rect 328 14504 360 14536
rect 400 14504 432 14536
rect 472 14504 504 14536
rect 544 14504 576 14536
rect 616 14504 648 14536
rect 688 14504 720 14536
rect 760 14504 792 14536
rect 832 14504 864 14536
rect 904 14504 936 14536
rect 976 14504 1008 14536
rect 1048 14504 1080 14536
rect 1120 14504 1152 14536
rect 1192 14504 1224 14536
rect 1264 14504 1296 14536
rect 1336 14504 1368 14536
rect 1408 14504 1440 14536
rect 1480 14504 1512 14536
rect 1552 14504 1584 14536
rect 1624 14504 1656 14536
rect 1696 14504 1728 14536
rect 1768 14504 1800 14536
rect 1840 14504 1872 14536
rect 1912 14504 1944 14536
rect 1984 14504 2016 14536
rect 2056 14504 2088 14536
rect 2128 14504 2160 14536
rect 2200 14504 2232 14536
rect 2272 14504 2304 14536
rect 2344 14504 2376 14536
rect 2416 14504 2448 14536
rect 2488 14504 2520 14536
rect 2560 14504 2592 14536
rect 2632 14504 2664 14536
rect 2704 14504 2736 14536
rect 2776 14504 2808 14536
rect 2848 14504 2880 14536
rect 2920 14504 2952 14536
rect 2992 14504 3024 14536
rect 3064 14504 3096 14536
rect 3136 14504 3168 14536
rect 3208 14504 3240 14536
rect 3280 14504 3312 14536
rect 3352 14504 3384 14536
rect 3424 14504 3456 14536
rect 3496 14504 3528 14536
rect 3568 14504 3600 14536
rect 3640 14504 3672 14536
rect 3712 14504 3744 14536
rect 3784 14504 3816 14536
rect 3856 14504 3888 14536
rect 112 14432 144 14464
rect 184 14432 216 14464
rect 256 14432 288 14464
rect 328 14432 360 14464
rect 400 14432 432 14464
rect 472 14432 504 14464
rect 544 14432 576 14464
rect 616 14432 648 14464
rect 688 14432 720 14464
rect 760 14432 792 14464
rect 832 14432 864 14464
rect 904 14432 936 14464
rect 976 14432 1008 14464
rect 1048 14432 1080 14464
rect 1120 14432 1152 14464
rect 1192 14432 1224 14464
rect 1264 14432 1296 14464
rect 1336 14432 1368 14464
rect 1408 14432 1440 14464
rect 1480 14432 1512 14464
rect 1552 14432 1584 14464
rect 1624 14432 1656 14464
rect 1696 14432 1728 14464
rect 1768 14432 1800 14464
rect 1840 14432 1872 14464
rect 1912 14432 1944 14464
rect 1984 14432 2016 14464
rect 2056 14432 2088 14464
rect 2128 14432 2160 14464
rect 2200 14432 2232 14464
rect 2272 14432 2304 14464
rect 2344 14432 2376 14464
rect 2416 14432 2448 14464
rect 2488 14432 2520 14464
rect 2560 14432 2592 14464
rect 2632 14432 2664 14464
rect 2704 14432 2736 14464
rect 2776 14432 2808 14464
rect 2848 14432 2880 14464
rect 2920 14432 2952 14464
rect 2992 14432 3024 14464
rect 3064 14432 3096 14464
rect 3136 14432 3168 14464
rect 3208 14432 3240 14464
rect 3280 14432 3312 14464
rect 3352 14432 3384 14464
rect 3424 14432 3456 14464
rect 3496 14432 3528 14464
rect 3568 14432 3600 14464
rect 3640 14432 3672 14464
rect 3712 14432 3744 14464
rect 3784 14432 3816 14464
rect 3856 14432 3888 14464
rect 112 14360 144 14392
rect 184 14360 216 14392
rect 256 14360 288 14392
rect 328 14360 360 14392
rect 400 14360 432 14392
rect 472 14360 504 14392
rect 544 14360 576 14392
rect 616 14360 648 14392
rect 688 14360 720 14392
rect 760 14360 792 14392
rect 832 14360 864 14392
rect 904 14360 936 14392
rect 976 14360 1008 14392
rect 1048 14360 1080 14392
rect 1120 14360 1152 14392
rect 1192 14360 1224 14392
rect 1264 14360 1296 14392
rect 1336 14360 1368 14392
rect 1408 14360 1440 14392
rect 1480 14360 1512 14392
rect 1552 14360 1584 14392
rect 1624 14360 1656 14392
rect 1696 14360 1728 14392
rect 1768 14360 1800 14392
rect 1840 14360 1872 14392
rect 1912 14360 1944 14392
rect 1984 14360 2016 14392
rect 2056 14360 2088 14392
rect 2128 14360 2160 14392
rect 2200 14360 2232 14392
rect 2272 14360 2304 14392
rect 2344 14360 2376 14392
rect 2416 14360 2448 14392
rect 2488 14360 2520 14392
rect 2560 14360 2592 14392
rect 2632 14360 2664 14392
rect 2704 14360 2736 14392
rect 2776 14360 2808 14392
rect 2848 14360 2880 14392
rect 2920 14360 2952 14392
rect 2992 14360 3024 14392
rect 3064 14360 3096 14392
rect 3136 14360 3168 14392
rect 3208 14360 3240 14392
rect 3280 14360 3312 14392
rect 3352 14360 3384 14392
rect 3424 14360 3456 14392
rect 3496 14360 3528 14392
rect 3568 14360 3600 14392
rect 3640 14360 3672 14392
rect 3712 14360 3744 14392
rect 3784 14360 3816 14392
rect 3856 14360 3888 14392
rect 112 14288 144 14320
rect 184 14288 216 14320
rect 256 14288 288 14320
rect 328 14288 360 14320
rect 400 14288 432 14320
rect 472 14288 504 14320
rect 544 14288 576 14320
rect 616 14288 648 14320
rect 688 14288 720 14320
rect 760 14288 792 14320
rect 832 14288 864 14320
rect 904 14288 936 14320
rect 976 14288 1008 14320
rect 1048 14288 1080 14320
rect 1120 14288 1152 14320
rect 1192 14288 1224 14320
rect 1264 14288 1296 14320
rect 1336 14288 1368 14320
rect 1408 14288 1440 14320
rect 1480 14288 1512 14320
rect 1552 14288 1584 14320
rect 1624 14288 1656 14320
rect 1696 14288 1728 14320
rect 1768 14288 1800 14320
rect 1840 14288 1872 14320
rect 1912 14288 1944 14320
rect 1984 14288 2016 14320
rect 2056 14288 2088 14320
rect 2128 14288 2160 14320
rect 2200 14288 2232 14320
rect 2272 14288 2304 14320
rect 2344 14288 2376 14320
rect 2416 14288 2448 14320
rect 2488 14288 2520 14320
rect 2560 14288 2592 14320
rect 2632 14288 2664 14320
rect 2704 14288 2736 14320
rect 2776 14288 2808 14320
rect 2848 14288 2880 14320
rect 2920 14288 2952 14320
rect 2992 14288 3024 14320
rect 3064 14288 3096 14320
rect 3136 14288 3168 14320
rect 3208 14288 3240 14320
rect 3280 14288 3312 14320
rect 3352 14288 3384 14320
rect 3424 14288 3456 14320
rect 3496 14288 3528 14320
rect 3568 14288 3600 14320
rect 3640 14288 3672 14320
rect 3712 14288 3744 14320
rect 3784 14288 3816 14320
rect 3856 14288 3888 14320
rect 112 14216 144 14248
rect 184 14216 216 14248
rect 256 14216 288 14248
rect 328 14216 360 14248
rect 400 14216 432 14248
rect 472 14216 504 14248
rect 544 14216 576 14248
rect 616 14216 648 14248
rect 688 14216 720 14248
rect 760 14216 792 14248
rect 832 14216 864 14248
rect 904 14216 936 14248
rect 976 14216 1008 14248
rect 1048 14216 1080 14248
rect 1120 14216 1152 14248
rect 1192 14216 1224 14248
rect 1264 14216 1296 14248
rect 1336 14216 1368 14248
rect 1408 14216 1440 14248
rect 1480 14216 1512 14248
rect 1552 14216 1584 14248
rect 1624 14216 1656 14248
rect 1696 14216 1728 14248
rect 1768 14216 1800 14248
rect 1840 14216 1872 14248
rect 1912 14216 1944 14248
rect 1984 14216 2016 14248
rect 2056 14216 2088 14248
rect 2128 14216 2160 14248
rect 2200 14216 2232 14248
rect 2272 14216 2304 14248
rect 2344 14216 2376 14248
rect 2416 14216 2448 14248
rect 2488 14216 2520 14248
rect 2560 14216 2592 14248
rect 2632 14216 2664 14248
rect 2704 14216 2736 14248
rect 2776 14216 2808 14248
rect 2848 14216 2880 14248
rect 2920 14216 2952 14248
rect 2992 14216 3024 14248
rect 3064 14216 3096 14248
rect 3136 14216 3168 14248
rect 3208 14216 3240 14248
rect 3280 14216 3312 14248
rect 3352 14216 3384 14248
rect 3424 14216 3456 14248
rect 3496 14216 3528 14248
rect 3568 14216 3600 14248
rect 3640 14216 3672 14248
rect 3712 14216 3744 14248
rect 3784 14216 3816 14248
rect 3856 14216 3888 14248
rect 112 14144 144 14176
rect 184 14144 216 14176
rect 256 14144 288 14176
rect 328 14144 360 14176
rect 400 14144 432 14176
rect 472 14144 504 14176
rect 544 14144 576 14176
rect 616 14144 648 14176
rect 688 14144 720 14176
rect 760 14144 792 14176
rect 832 14144 864 14176
rect 904 14144 936 14176
rect 976 14144 1008 14176
rect 1048 14144 1080 14176
rect 1120 14144 1152 14176
rect 1192 14144 1224 14176
rect 1264 14144 1296 14176
rect 1336 14144 1368 14176
rect 1408 14144 1440 14176
rect 1480 14144 1512 14176
rect 1552 14144 1584 14176
rect 1624 14144 1656 14176
rect 1696 14144 1728 14176
rect 1768 14144 1800 14176
rect 1840 14144 1872 14176
rect 1912 14144 1944 14176
rect 1984 14144 2016 14176
rect 2056 14144 2088 14176
rect 2128 14144 2160 14176
rect 2200 14144 2232 14176
rect 2272 14144 2304 14176
rect 2344 14144 2376 14176
rect 2416 14144 2448 14176
rect 2488 14144 2520 14176
rect 2560 14144 2592 14176
rect 2632 14144 2664 14176
rect 2704 14144 2736 14176
rect 2776 14144 2808 14176
rect 2848 14144 2880 14176
rect 2920 14144 2952 14176
rect 2992 14144 3024 14176
rect 3064 14144 3096 14176
rect 3136 14144 3168 14176
rect 3208 14144 3240 14176
rect 3280 14144 3312 14176
rect 3352 14144 3384 14176
rect 3424 14144 3456 14176
rect 3496 14144 3528 14176
rect 3568 14144 3600 14176
rect 3640 14144 3672 14176
rect 3712 14144 3744 14176
rect 3784 14144 3816 14176
rect 3856 14144 3888 14176
rect 112 14072 144 14104
rect 184 14072 216 14104
rect 256 14072 288 14104
rect 328 14072 360 14104
rect 400 14072 432 14104
rect 472 14072 504 14104
rect 544 14072 576 14104
rect 616 14072 648 14104
rect 688 14072 720 14104
rect 760 14072 792 14104
rect 832 14072 864 14104
rect 904 14072 936 14104
rect 976 14072 1008 14104
rect 1048 14072 1080 14104
rect 1120 14072 1152 14104
rect 1192 14072 1224 14104
rect 1264 14072 1296 14104
rect 1336 14072 1368 14104
rect 1408 14072 1440 14104
rect 1480 14072 1512 14104
rect 1552 14072 1584 14104
rect 1624 14072 1656 14104
rect 1696 14072 1728 14104
rect 1768 14072 1800 14104
rect 1840 14072 1872 14104
rect 1912 14072 1944 14104
rect 1984 14072 2016 14104
rect 2056 14072 2088 14104
rect 2128 14072 2160 14104
rect 2200 14072 2232 14104
rect 2272 14072 2304 14104
rect 2344 14072 2376 14104
rect 2416 14072 2448 14104
rect 2488 14072 2520 14104
rect 2560 14072 2592 14104
rect 2632 14072 2664 14104
rect 2704 14072 2736 14104
rect 2776 14072 2808 14104
rect 2848 14072 2880 14104
rect 2920 14072 2952 14104
rect 2992 14072 3024 14104
rect 3064 14072 3096 14104
rect 3136 14072 3168 14104
rect 3208 14072 3240 14104
rect 3280 14072 3312 14104
rect 3352 14072 3384 14104
rect 3424 14072 3456 14104
rect 3496 14072 3528 14104
rect 3568 14072 3600 14104
rect 3640 14072 3672 14104
rect 3712 14072 3744 14104
rect 3784 14072 3816 14104
rect 3856 14072 3888 14104
rect 112 14000 144 14032
rect 184 14000 216 14032
rect 256 14000 288 14032
rect 328 14000 360 14032
rect 400 14000 432 14032
rect 472 14000 504 14032
rect 544 14000 576 14032
rect 616 14000 648 14032
rect 688 14000 720 14032
rect 760 14000 792 14032
rect 832 14000 864 14032
rect 904 14000 936 14032
rect 976 14000 1008 14032
rect 1048 14000 1080 14032
rect 1120 14000 1152 14032
rect 1192 14000 1224 14032
rect 1264 14000 1296 14032
rect 1336 14000 1368 14032
rect 1408 14000 1440 14032
rect 1480 14000 1512 14032
rect 1552 14000 1584 14032
rect 1624 14000 1656 14032
rect 1696 14000 1728 14032
rect 1768 14000 1800 14032
rect 1840 14000 1872 14032
rect 1912 14000 1944 14032
rect 1984 14000 2016 14032
rect 2056 14000 2088 14032
rect 2128 14000 2160 14032
rect 2200 14000 2232 14032
rect 2272 14000 2304 14032
rect 2344 14000 2376 14032
rect 2416 14000 2448 14032
rect 2488 14000 2520 14032
rect 2560 14000 2592 14032
rect 2632 14000 2664 14032
rect 2704 14000 2736 14032
rect 2776 14000 2808 14032
rect 2848 14000 2880 14032
rect 2920 14000 2952 14032
rect 2992 14000 3024 14032
rect 3064 14000 3096 14032
rect 3136 14000 3168 14032
rect 3208 14000 3240 14032
rect 3280 14000 3312 14032
rect 3352 14000 3384 14032
rect 3424 14000 3456 14032
rect 3496 14000 3528 14032
rect 3568 14000 3600 14032
rect 3640 14000 3672 14032
rect 3712 14000 3744 14032
rect 3784 14000 3816 14032
rect 3856 14000 3888 14032
rect 112 13928 144 13960
rect 184 13928 216 13960
rect 256 13928 288 13960
rect 328 13928 360 13960
rect 400 13928 432 13960
rect 472 13928 504 13960
rect 544 13928 576 13960
rect 616 13928 648 13960
rect 688 13928 720 13960
rect 760 13928 792 13960
rect 832 13928 864 13960
rect 904 13928 936 13960
rect 976 13928 1008 13960
rect 1048 13928 1080 13960
rect 1120 13928 1152 13960
rect 1192 13928 1224 13960
rect 1264 13928 1296 13960
rect 1336 13928 1368 13960
rect 1408 13928 1440 13960
rect 1480 13928 1512 13960
rect 1552 13928 1584 13960
rect 1624 13928 1656 13960
rect 1696 13928 1728 13960
rect 1768 13928 1800 13960
rect 1840 13928 1872 13960
rect 1912 13928 1944 13960
rect 1984 13928 2016 13960
rect 2056 13928 2088 13960
rect 2128 13928 2160 13960
rect 2200 13928 2232 13960
rect 2272 13928 2304 13960
rect 2344 13928 2376 13960
rect 2416 13928 2448 13960
rect 2488 13928 2520 13960
rect 2560 13928 2592 13960
rect 2632 13928 2664 13960
rect 2704 13928 2736 13960
rect 2776 13928 2808 13960
rect 2848 13928 2880 13960
rect 2920 13928 2952 13960
rect 2992 13928 3024 13960
rect 3064 13928 3096 13960
rect 3136 13928 3168 13960
rect 3208 13928 3240 13960
rect 3280 13928 3312 13960
rect 3352 13928 3384 13960
rect 3424 13928 3456 13960
rect 3496 13928 3528 13960
rect 3568 13928 3600 13960
rect 3640 13928 3672 13960
rect 3712 13928 3744 13960
rect 3784 13928 3816 13960
rect 3856 13928 3888 13960
rect 112 13856 144 13888
rect 184 13856 216 13888
rect 256 13856 288 13888
rect 328 13856 360 13888
rect 400 13856 432 13888
rect 472 13856 504 13888
rect 544 13856 576 13888
rect 616 13856 648 13888
rect 688 13856 720 13888
rect 760 13856 792 13888
rect 832 13856 864 13888
rect 904 13856 936 13888
rect 976 13856 1008 13888
rect 1048 13856 1080 13888
rect 1120 13856 1152 13888
rect 1192 13856 1224 13888
rect 1264 13856 1296 13888
rect 1336 13856 1368 13888
rect 1408 13856 1440 13888
rect 1480 13856 1512 13888
rect 1552 13856 1584 13888
rect 1624 13856 1656 13888
rect 1696 13856 1728 13888
rect 1768 13856 1800 13888
rect 1840 13856 1872 13888
rect 1912 13856 1944 13888
rect 1984 13856 2016 13888
rect 2056 13856 2088 13888
rect 2128 13856 2160 13888
rect 2200 13856 2232 13888
rect 2272 13856 2304 13888
rect 2344 13856 2376 13888
rect 2416 13856 2448 13888
rect 2488 13856 2520 13888
rect 2560 13856 2592 13888
rect 2632 13856 2664 13888
rect 2704 13856 2736 13888
rect 2776 13856 2808 13888
rect 2848 13856 2880 13888
rect 2920 13856 2952 13888
rect 2992 13856 3024 13888
rect 3064 13856 3096 13888
rect 3136 13856 3168 13888
rect 3208 13856 3240 13888
rect 3280 13856 3312 13888
rect 3352 13856 3384 13888
rect 3424 13856 3456 13888
rect 3496 13856 3528 13888
rect 3568 13856 3600 13888
rect 3640 13856 3672 13888
rect 3712 13856 3744 13888
rect 3784 13856 3816 13888
rect 3856 13856 3888 13888
rect 112 13784 144 13816
rect 184 13784 216 13816
rect 256 13784 288 13816
rect 328 13784 360 13816
rect 400 13784 432 13816
rect 472 13784 504 13816
rect 544 13784 576 13816
rect 616 13784 648 13816
rect 688 13784 720 13816
rect 760 13784 792 13816
rect 832 13784 864 13816
rect 904 13784 936 13816
rect 976 13784 1008 13816
rect 1048 13784 1080 13816
rect 1120 13784 1152 13816
rect 1192 13784 1224 13816
rect 1264 13784 1296 13816
rect 1336 13784 1368 13816
rect 1408 13784 1440 13816
rect 1480 13784 1512 13816
rect 1552 13784 1584 13816
rect 1624 13784 1656 13816
rect 1696 13784 1728 13816
rect 1768 13784 1800 13816
rect 1840 13784 1872 13816
rect 1912 13784 1944 13816
rect 1984 13784 2016 13816
rect 2056 13784 2088 13816
rect 2128 13784 2160 13816
rect 2200 13784 2232 13816
rect 2272 13784 2304 13816
rect 2344 13784 2376 13816
rect 2416 13784 2448 13816
rect 2488 13784 2520 13816
rect 2560 13784 2592 13816
rect 2632 13784 2664 13816
rect 2704 13784 2736 13816
rect 2776 13784 2808 13816
rect 2848 13784 2880 13816
rect 2920 13784 2952 13816
rect 2992 13784 3024 13816
rect 3064 13784 3096 13816
rect 3136 13784 3168 13816
rect 3208 13784 3240 13816
rect 3280 13784 3312 13816
rect 3352 13784 3384 13816
rect 3424 13784 3456 13816
rect 3496 13784 3528 13816
rect 3568 13784 3600 13816
rect 3640 13784 3672 13816
rect 3712 13784 3744 13816
rect 3784 13784 3816 13816
rect 3856 13784 3888 13816
rect 112 13712 144 13744
rect 184 13712 216 13744
rect 256 13712 288 13744
rect 328 13712 360 13744
rect 400 13712 432 13744
rect 472 13712 504 13744
rect 544 13712 576 13744
rect 616 13712 648 13744
rect 688 13712 720 13744
rect 760 13712 792 13744
rect 832 13712 864 13744
rect 904 13712 936 13744
rect 976 13712 1008 13744
rect 1048 13712 1080 13744
rect 1120 13712 1152 13744
rect 1192 13712 1224 13744
rect 1264 13712 1296 13744
rect 1336 13712 1368 13744
rect 1408 13712 1440 13744
rect 1480 13712 1512 13744
rect 1552 13712 1584 13744
rect 1624 13712 1656 13744
rect 1696 13712 1728 13744
rect 1768 13712 1800 13744
rect 1840 13712 1872 13744
rect 1912 13712 1944 13744
rect 1984 13712 2016 13744
rect 2056 13712 2088 13744
rect 2128 13712 2160 13744
rect 2200 13712 2232 13744
rect 2272 13712 2304 13744
rect 2344 13712 2376 13744
rect 2416 13712 2448 13744
rect 2488 13712 2520 13744
rect 2560 13712 2592 13744
rect 2632 13712 2664 13744
rect 2704 13712 2736 13744
rect 2776 13712 2808 13744
rect 2848 13712 2880 13744
rect 2920 13712 2952 13744
rect 2992 13712 3024 13744
rect 3064 13712 3096 13744
rect 3136 13712 3168 13744
rect 3208 13712 3240 13744
rect 3280 13712 3312 13744
rect 3352 13712 3384 13744
rect 3424 13712 3456 13744
rect 3496 13712 3528 13744
rect 3568 13712 3600 13744
rect 3640 13712 3672 13744
rect 3712 13712 3744 13744
rect 3784 13712 3816 13744
rect 3856 13712 3888 13744
rect 112 13640 144 13672
rect 184 13640 216 13672
rect 256 13640 288 13672
rect 328 13640 360 13672
rect 400 13640 432 13672
rect 472 13640 504 13672
rect 544 13640 576 13672
rect 616 13640 648 13672
rect 688 13640 720 13672
rect 760 13640 792 13672
rect 832 13640 864 13672
rect 904 13640 936 13672
rect 976 13640 1008 13672
rect 1048 13640 1080 13672
rect 1120 13640 1152 13672
rect 1192 13640 1224 13672
rect 1264 13640 1296 13672
rect 1336 13640 1368 13672
rect 1408 13640 1440 13672
rect 1480 13640 1512 13672
rect 1552 13640 1584 13672
rect 1624 13640 1656 13672
rect 1696 13640 1728 13672
rect 1768 13640 1800 13672
rect 1840 13640 1872 13672
rect 1912 13640 1944 13672
rect 1984 13640 2016 13672
rect 2056 13640 2088 13672
rect 2128 13640 2160 13672
rect 2200 13640 2232 13672
rect 2272 13640 2304 13672
rect 2344 13640 2376 13672
rect 2416 13640 2448 13672
rect 2488 13640 2520 13672
rect 2560 13640 2592 13672
rect 2632 13640 2664 13672
rect 2704 13640 2736 13672
rect 2776 13640 2808 13672
rect 2848 13640 2880 13672
rect 2920 13640 2952 13672
rect 2992 13640 3024 13672
rect 3064 13640 3096 13672
rect 3136 13640 3168 13672
rect 3208 13640 3240 13672
rect 3280 13640 3312 13672
rect 3352 13640 3384 13672
rect 3424 13640 3456 13672
rect 3496 13640 3528 13672
rect 3568 13640 3600 13672
rect 3640 13640 3672 13672
rect 3712 13640 3744 13672
rect 3784 13640 3816 13672
rect 3856 13640 3888 13672
rect 112 13568 144 13600
rect 184 13568 216 13600
rect 256 13568 288 13600
rect 328 13568 360 13600
rect 400 13568 432 13600
rect 472 13568 504 13600
rect 544 13568 576 13600
rect 616 13568 648 13600
rect 688 13568 720 13600
rect 760 13568 792 13600
rect 832 13568 864 13600
rect 904 13568 936 13600
rect 976 13568 1008 13600
rect 1048 13568 1080 13600
rect 1120 13568 1152 13600
rect 1192 13568 1224 13600
rect 1264 13568 1296 13600
rect 1336 13568 1368 13600
rect 1408 13568 1440 13600
rect 1480 13568 1512 13600
rect 1552 13568 1584 13600
rect 1624 13568 1656 13600
rect 1696 13568 1728 13600
rect 1768 13568 1800 13600
rect 1840 13568 1872 13600
rect 1912 13568 1944 13600
rect 1984 13568 2016 13600
rect 2056 13568 2088 13600
rect 2128 13568 2160 13600
rect 2200 13568 2232 13600
rect 2272 13568 2304 13600
rect 2344 13568 2376 13600
rect 2416 13568 2448 13600
rect 2488 13568 2520 13600
rect 2560 13568 2592 13600
rect 2632 13568 2664 13600
rect 2704 13568 2736 13600
rect 2776 13568 2808 13600
rect 2848 13568 2880 13600
rect 2920 13568 2952 13600
rect 2992 13568 3024 13600
rect 3064 13568 3096 13600
rect 3136 13568 3168 13600
rect 3208 13568 3240 13600
rect 3280 13568 3312 13600
rect 3352 13568 3384 13600
rect 3424 13568 3456 13600
rect 3496 13568 3528 13600
rect 3568 13568 3600 13600
rect 3640 13568 3672 13600
rect 3712 13568 3744 13600
rect 3784 13568 3816 13600
rect 3856 13568 3888 13600
rect 112 13496 144 13528
rect 184 13496 216 13528
rect 256 13496 288 13528
rect 328 13496 360 13528
rect 400 13496 432 13528
rect 472 13496 504 13528
rect 544 13496 576 13528
rect 616 13496 648 13528
rect 688 13496 720 13528
rect 760 13496 792 13528
rect 832 13496 864 13528
rect 904 13496 936 13528
rect 976 13496 1008 13528
rect 1048 13496 1080 13528
rect 1120 13496 1152 13528
rect 1192 13496 1224 13528
rect 1264 13496 1296 13528
rect 1336 13496 1368 13528
rect 1408 13496 1440 13528
rect 1480 13496 1512 13528
rect 1552 13496 1584 13528
rect 1624 13496 1656 13528
rect 1696 13496 1728 13528
rect 1768 13496 1800 13528
rect 1840 13496 1872 13528
rect 1912 13496 1944 13528
rect 1984 13496 2016 13528
rect 2056 13496 2088 13528
rect 2128 13496 2160 13528
rect 2200 13496 2232 13528
rect 2272 13496 2304 13528
rect 2344 13496 2376 13528
rect 2416 13496 2448 13528
rect 2488 13496 2520 13528
rect 2560 13496 2592 13528
rect 2632 13496 2664 13528
rect 2704 13496 2736 13528
rect 2776 13496 2808 13528
rect 2848 13496 2880 13528
rect 2920 13496 2952 13528
rect 2992 13496 3024 13528
rect 3064 13496 3096 13528
rect 3136 13496 3168 13528
rect 3208 13496 3240 13528
rect 3280 13496 3312 13528
rect 3352 13496 3384 13528
rect 3424 13496 3456 13528
rect 3496 13496 3528 13528
rect 3568 13496 3600 13528
rect 3640 13496 3672 13528
rect 3712 13496 3744 13528
rect 3784 13496 3816 13528
rect 3856 13496 3888 13528
rect 112 13424 144 13456
rect 184 13424 216 13456
rect 256 13424 288 13456
rect 328 13424 360 13456
rect 400 13424 432 13456
rect 472 13424 504 13456
rect 544 13424 576 13456
rect 616 13424 648 13456
rect 688 13424 720 13456
rect 760 13424 792 13456
rect 832 13424 864 13456
rect 904 13424 936 13456
rect 976 13424 1008 13456
rect 1048 13424 1080 13456
rect 1120 13424 1152 13456
rect 1192 13424 1224 13456
rect 1264 13424 1296 13456
rect 1336 13424 1368 13456
rect 1408 13424 1440 13456
rect 1480 13424 1512 13456
rect 1552 13424 1584 13456
rect 1624 13424 1656 13456
rect 1696 13424 1728 13456
rect 1768 13424 1800 13456
rect 1840 13424 1872 13456
rect 1912 13424 1944 13456
rect 1984 13424 2016 13456
rect 2056 13424 2088 13456
rect 2128 13424 2160 13456
rect 2200 13424 2232 13456
rect 2272 13424 2304 13456
rect 2344 13424 2376 13456
rect 2416 13424 2448 13456
rect 2488 13424 2520 13456
rect 2560 13424 2592 13456
rect 2632 13424 2664 13456
rect 2704 13424 2736 13456
rect 2776 13424 2808 13456
rect 2848 13424 2880 13456
rect 2920 13424 2952 13456
rect 2992 13424 3024 13456
rect 3064 13424 3096 13456
rect 3136 13424 3168 13456
rect 3208 13424 3240 13456
rect 3280 13424 3312 13456
rect 3352 13424 3384 13456
rect 3424 13424 3456 13456
rect 3496 13424 3528 13456
rect 3568 13424 3600 13456
rect 3640 13424 3672 13456
rect 3712 13424 3744 13456
rect 3784 13424 3816 13456
rect 3856 13424 3888 13456
rect 112 13352 144 13384
rect 184 13352 216 13384
rect 256 13352 288 13384
rect 328 13352 360 13384
rect 400 13352 432 13384
rect 472 13352 504 13384
rect 544 13352 576 13384
rect 616 13352 648 13384
rect 688 13352 720 13384
rect 760 13352 792 13384
rect 832 13352 864 13384
rect 904 13352 936 13384
rect 976 13352 1008 13384
rect 1048 13352 1080 13384
rect 1120 13352 1152 13384
rect 1192 13352 1224 13384
rect 1264 13352 1296 13384
rect 1336 13352 1368 13384
rect 1408 13352 1440 13384
rect 1480 13352 1512 13384
rect 1552 13352 1584 13384
rect 1624 13352 1656 13384
rect 1696 13352 1728 13384
rect 1768 13352 1800 13384
rect 1840 13352 1872 13384
rect 1912 13352 1944 13384
rect 1984 13352 2016 13384
rect 2056 13352 2088 13384
rect 2128 13352 2160 13384
rect 2200 13352 2232 13384
rect 2272 13352 2304 13384
rect 2344 13352 2376 13384
rect 2416 13352 2448 13384
rect 2488 13352 2520 13384
rect 2560 13352 2592 13384
rect 2632 13352 2664 13384
rect 2704 13352 2736 13384
rect 2776 13352 2808 13384
rect 2848 13352 2880 13384
rect 2920 13352 2952 13384
rect 2992 13352 3024 13384
rect 3064 13352 3096 13384
rect 3136 13352 3168 13384
rect 3208 13352 3240 13384
rect 3280 13352 3312 13384
rect 3352 13352 3384 13384
rect 3424 13352 3456 13384
rect 3496 13352 3528 13384
rect 3568 13352 3600 13384
rect 3640 13352 3672 13384
rect 3712 13352 3744 13384
rect 3784 13352 3816 13384
rect 3856 13352 3888 13384
rect 112 13280 144 13312
rect 184 13280 216 13312
rect 256 13280 288 13312
rect 328 13280 360 13312
rect 400 13280 432 13312
rect 472 13280 504 13312
rect 544 13280 576 13312
rect 616 13280 648 13312
rect 688 13280 720 13312
rect 760 13280 792 13312
rect 832 13280 864 13312
rect 904 13280 936 13312
rect 976 13280 1008 13312
rect 1048 13280 1080 13312
rect 1120 13280 1152 13312
rect 1192 13280 1224 13312
rect 1264 13280 1296 13312
rect 1336 13280 1368 13312
rect 1408 13280 1440 13312
rect 1480 13280 1512 13312
rect 1552 13280 1584 13312
rect 1624 13280 1656 13312
rect 1696 13280 1728 13312
rect 1768 13280 1800 13312
rect 1840 13280 1872 13312
rect 1912 13280 1944 13312
rect 1984 13280 2016 13312
rect 2056 13280 2088 13312
rect 2128 13280 2160 13312
rect 2200 13280 2232 13312
rect 2272 13280 2304 13312
rect 2344 13280 2376 13312
rect 2416 13280 2448 13312
rect 2488 13280 2520 13312
rect 2560 13280 2592 13312
rect 2632 13280 2664 13312
rect 2704 13280 2736 13312
rect 2776 13280 2808 13312
rect 2848 13280 2880 13312
rect 2920 13280 2952 13312
rect 2992 13280 3024 13312
rect 3064 13280 3096 13312
rect 3136 13280 3168 13312
rect 3208 13280 3240 13312
rect 3280 13280 3312 13312
rect 3352 13280 3384 13312
rect 3424 13280 3456 13312
rect 3496 13280 3528 13312
rect 3568 13280 3600 13312
rect 3640 13280 3672 13312
rect 3712 13280 3744 13312
rect 3784 13280 3816 13312
rect 3856 13280 3888 13312
rect 112 13208 144 13240
rect 184 13208 216 13240
rect 256 13208 288 13240
rect 328 13208 360 13240
rect 400 13208 432 13240
rect 472 13208 504 13240
rect 544 13208 576 13240
rect 616 13208 648 13240
rect 688 13208 720 13240
rect 760 13208 792 13240
rect 832 13208 864 13240
rect 904 13208 936 13240
rect 976 13208 1008 13240
rect 1048 13208 1080 13240
rect 1120 13208 1152 13240
rect 1192 13208 1224 13240
rect 1264 13208 1296 13240
rect 1336 13208 1368 13240
rect 1408 13208 1440 13240
rect 1480 13208 1512 13240
rect 1552 13208 1584 13240
rect 1624 13208 1656 13240
rect 1696 13208 1728 13240
rect 1768 13208 1800 13240
rect 1840 13208 1872 13240
rect 1912 13208 1944 13240
rect 1984 13208 2016 13240
rect 2056 13208 2088 13240
rect 2128 13208 2160 13240
rect 2200 13208 2232 13240
rect 2272 13208 2304 13240
rect 2344 13208 2376 13240
rect 2416 13208 2448 13240
rect 2488 13208 2520 13240
rect 2560 13208 2592 13240
rect 2632 13208 2664 13240
rect 2704 13208 2736 13240
rect 2776 13208 2808 13240
rect 2848 13208 2880 13240
rect 2920 13208 2952 13240
rect 2992 13208 3024 13240
rect 3064 13208 3096 13240
rect 3136 13208 3168 13240
rect 3208 13208 3240 13240
rect 3280 13208 3312 13240
rect 3352 13208 3384 13240
rect 3424 13208 3456 13240
rect 3496 13208 3528 13240
rect 3568 13208 3600 13240
rect 3640 13208 3672 13240
rect 3712 13208 3744 13240
rect 3784 13208 3816 13240
rect 3856 13208 3888 13240
rect 112 13136 144 13168
rect 184 13136 216 13168
rect 256 13136 288 13168
rect 328 13136 360 13168
rect 400 13136 432 13168
rect 472 13136 504 13168
rect 544 13136 576 13168
rect 616 13136 648 13168
rect 688 13136 720 13168
rect 760 13136 792 13168
rect 832 13136 864 13168
rect 904 13136 936 13168
rect 976 13136 1008 13168
rect 1048 13136 1080 13168
rect 1120 13136 1152 13168
rect 1192 13136 1224 13168
rect 1264 13136 1296 13168
rect 1336 13136 1368 13168
rect 1408 13136 1440 13168
rect 1480 13136 1512 13168
rect 1552 13136 1584 13168
rect 1624 13136 1656 13168
rect 1696 13136 1728 13168
rect 1768 13136 1800 13168
rect 1840 13136 1872 13168
rect 1912 13136 1944 13168
rect 1984 13136 2016 13168
rect 2056 13136 2088 13168
rect 2128 13136 2160 13168
rect 2200 13136 2232 13168
rect 2272 13136 2304 13168
rect 2344 13136 2376 13168
rect 2416 13136 2448 13168
rect 2488 13136 2520 13168
rect 2560 13136 2592 13168
rect 2632 13136 2664 13168
rect 2704 13136 2736 13168
rect 2776 13136 2808 13168
rect 2848 13136 2880 13168
rect 2920 13136 2952 13168
rect 2992 13136 3024 13168
rect 3064 13136 3096 13168
rect 3136 13136 3168 13168
rect 3208 13136 3240 13168
rect 3280 13136 3312 13168
rect 3352 13136 3384 13168
rect 3424 13136 3456 13168
rect 3496 13136 3528 13168
rect 3568 13136 3600 13168
rect 3640 13136 3672 13168
rect 3712 13136 3744 13168
rect 3784 13136 3816 13168
rect 3856 13136 3888 13168
rect 112 13064 144 13096
rect 184 13064 216 13096
rect 256 13064 288 13096
rect 328 13064 360 13096
rect 400 13064 432 13096
rect 472 13064 504 13096
rect 544 13064 576 13096
rect 616 13064 648 13096
rect 688 13064 720 13096
rect 760 13064 792 13096
rect 832 13064 864 13096
rect 904 13064 936 13096
rect 976 13064 1008 13096
rect 1048 13064 1080 13096
rect 1120 13064 1152 13096
rect 1192 13064 1224 13096
rect 1264 13064 1296 13096
rect 1336 13064 1368 13096
rect 1408 13064 1440 13096
rect 1480 13064 1512 13096
rect 1552 13064 1584 13096
rect 1624 13064 1656 13096
rect 1696 13064 1728 13096
rect 1768 13064 1800 13096
rect 1840 13064 1872 13096
rect 1912 13064 1944 13096
rect 1984 13064 2016 13096
rect 2056 13064 2088 13096
rect 2128 13064 2160 13096
rect 2200 13064 2232 13096
rect 2272 13064 2304 13096
rect 2344 13064 2376 13096
rect 2416 13064 2448 13096
rect 2488 13064 2520 13096
rect 2560 13064 2592 13096
rect 2632 13064 2664 13096
rect 2704 13064 2736 13096
rect 2776 13064 2808 13096
rect 2848 13064 2880 13096
rect 2920 13064 2952 13096
rect 2992 13064 3024 13096
rect 3064 13064 3096 13096
rect 3136 13064 3168 13096
rect 3208 13064 3240 13096
rect 3280 13064 3312 13096
rect 3352 13064 3384 13096
rect 3424 13064 3456 13096
rect 3496 13064 3528 13096
rect 3568 13064 3600 13096
rect 3640 13064 3672 13096
rect 3712 13064 3744 13096
rect 3784 13064 3816 13096
rect 3856 13064 3888 13096
rect 0 33384 112 33416
rect 144 33384 184 33416
rect 216 33384 256 33416
rect 288 33384 328 33416
rect 360 33384 400 33416
rect 432 33384 472 33416
rect 504 33384 544 33416
rect 576 33384 616 33416
rect 648 33384 688 33416
rect 720 33384 760 33416
rect 792 33384 832 33416
rect 864 33384 904 33416
rect 936 33384 976 33416
rect 1008 33384 1048 33416
rect 1080 33384 1120 33416
rect 1152 33384 1192 33416
rect 1224 33384 1264 33416
rect 1296 33384 1336 33416
rect 1368 33384 1408 33416
rect 1440 33384 1480 33416
rect 1512 33384 1552 33416
rect 1584 33384 1624 33416
rect 1656 33384 1696 33416
rect 1728 33384 1768 33416
rect 1800 33384 1840 33416
rect 1872 33384 1912 33416
rect 1944 33384 1984 33416
rect 2016 33384 2056 33416
rect 2088 33384 2128 33416
rect 2160 33384 2200 33416
rect 2232 33384 2272 33416
rect 2304 33384 2344 33416
rect 2376 33384 2416 33416
rect 2448 33384 2488 33416
rect 2520 33384 2560 33416
rect 2592 33384 2632 33416
rect 2664 33384 2704 33416
rect 2736 33384 2776 33416
rect 2808 33384 2848 33416
rect 2880 33384 2920 33416
rect 2952 33384 2992 33416
rect 3024 33384 3064 33416
rect 3096 33384 3136 33416
rect 3168 33384 3208 33416
rect 3240 33384 3280 33416
rect 3312 33384 3352 33416
rect 3384 33384 3424 33416
rect 3456 33384 3496 33416
rect 3528 33384 3568 33416
rect 3600 33384 3640 33416
rect 3672 33384 3712 33416
rect 3744 33384 3784 33416
rect 3816 33384 3856 33416
rect 3888 33384 4000 33416
rect 0 31384 112 31416
rect 144 31384 184 31416
rect 216 31384 256 31416
rect 288 31384 328 31416
rect 360 31384 400 31416
rect 432 31384 472 31416
rect 504 31384 544 31416
rect 576 31384 616 31416
rect 648 31384 688 31416
rect 720 31384 760 31416
rect 792 31384 832 31416
rect 864 31384 904 31416
rect 936 31384 976 31416
rect 1008 31384 1048 31416
rect 1080 31384 1120 31416
rect 1152 31384 1192 31416
rect 1224 31384 1264 31416
rect 1296 31384 1336 31416
rect 1368 31384 1408 31416
rect 1440 31384 1480 31416
rect 1512 31384 1552 31416
rect 1584 31384 1624 31416
rect 1656 31384 1696 31416
rect 1728 31384 1768 31416
rect 1800 31384 1840 31416
rect 1872 31384 1912 31416
rect 1944 31384 1984 31416
rect 2016 31384 2056 31416
rect 2088 31384 2128 31416
rect 2160 31384 2200 31416
rect 2232 31384 2272 31416
rect 2304 31384 2344 31416
rect 2376 31384 2416 31416
rect 2448 31384 2488 31416
rect 2520 31384 2560 31416
rect 2592 31384 2632 31416
rect 2664 31384 2704 31416
rect 2736 31384 2776 31416
rect 2808 31384 2848 31416
rect 2880 31384 2920 31416
rect 2952 31384 2992 31416
rect 3024 31384 3064 31416
rect 3096 31384 3136 31416
rect 3168 31384 3208 31416
rect 3240 31384 3280 31416
rect 3312 31384 3352 31416
rect 3384 31384 3424 31416
rect 3456 31384 3496 31416
rect 3528 31384 3568 31416
rect 3600 31384 3640 31416
rect 3672 31384 3712 31416
rect 3744 31384 3784 31416
rect 3816 31384 3856 31416
rect 3888 31384 4000 31416
rect 0 29684 112 29716
rect 144 29684 184 29716
rect 216 29684 256 29716
rect 288 29684 328 29716
rect 360 29684 400 29716
rect 432 29684 472 29716
rect 504 29684 544 29716
rect 576 29684 616 29716
rect 648 29684 688 29716
rect 720 29684 760 29716
rect 792 29684 832 29716
rect 864 29684 904 29716
rect 936 29684 976 29716
rect 1008 29684 1048 29716
rect 1080 29684 1120 29716
rect 1152 29684 1192 29716
rect 1224 29684 1264 29716
rect 1296 29684 1336 29716
rect 1368 29684 1408 29716
rect 1440 29684 1480 29716
rect 1512 29684 1552 29716
rect 1584 29684 1624 29716
rect 1656 29684 1696 29716
rect 1728 29684 1768 29716
rect 1800 29684 1840 29716
rect 1872 29684 1912 29716
rect 1944 29684 1984 29716
rect 2016 29684 2056 29716
rect 2088 29684 2128 29716
rect 2160 29684 2200 29716
rect 2232 29684 2272 29716
rect 2304 29684 2344 29716
rect 2376 29684 2416 29716
rect 2448 29684 2488 29716
rect 2520 29684 2560 29716
rect 2592 29684 2632 29716
rect 2664 29684 2704 29716
rect 2736 29684 2776 29716
rect 2808 29684 2848 29716
rect 2880 29684 2920 29716
rect 2952 29684 2992 29716
rect 3024 29684 3064 29716
rect 3096 29684 3136 29716
rect 3168 29684 3208 29716
rect 3240 29684 3280 29716
rect 3312 29684 3352 29716
rect 3384 29684 3424 29716
rect 3456 29684 3496 29716
rect 3528 29684 3568 29716
rect 3600 29684 3640 29716
rect 3672 29684 3712 29716
rect 3744 29684 3784 29716
rect 3816 29684 3856 29716
rect 3888 29684 4000 29716
rect 0 27971 4000 28034
rect 0 27939 112 27971
rect 144 27939 184 27971
rect 216 27939 256 27971
rect 288 27939 328 27971
rect 360 27939 400 27971
rect 432 27939 472 27971
rect 504 27939 544 27971
rect 576 27939 616 27971
rect 648 27939 688 27971
rect 720 27939 760 27971
rect 792 27939 832 27971
rect 864 27939 904 27971
rect 936 27939 976 27971
rect 1008 27939 1048 27971
rect 1080 27939 1120 27971
rect 1152 27939 1192 27971
rect 1224 27939 1264 27971
rect 1296 27939 1336 27971
rect 1368 27939 1408 27971
rect 1440 27939 1480 27971
rect 1512 27939 1552 27971
rect 1584 27939 1624 27971
rect 1656 27939 1696 27971
rect 1728 27939 1768 27971
rect 1800 27939 1840 27971
rect 1872 27939 1912 27971
rect 1944 27939 1984 27971
rect 2016 27939 2056 27971
rect 2088 27939 2128 27971
rect 2160 27939 2200 27971
rect 2232 27939 2272 27971
rect 2304 27939 2344 27971
rect 2376 27939 2416 27971
rect 2448 27939 2488 27971
rect 2520 27939 2560 27971
rect 2592 27939 2632 27971
rect 2664 27939 2704 27971
rect 2736 27939 2776 27971
rect 2808 27939 2848 27971
rect 2880 27939 2920 27971
rect 2952 27939 2992 27971
rect 3024 27939 3064 27971
rect 3096 27939 3136 27971
rect 3168 27939 3208 27971
rect 3240 27939 3280 27971
rect 3312 27939 3352 27971
rect 3384 27939 3424 27971
rect 3456 27939 3496 27971
rect 3528 27939 3568 27971
rect 3600 27939 3640 27971
rect 3672 27939 3712 27971
rect 3744 27939 3784 27971
rect 3816 27939 3856 27971
rect 3888 27939 4000 27971
rect 0 27899 4000 27939
rect 0 27867 112 27899
rect 144 27867 184 27899
rect 216 27867 256 27899
rect 288 27867 328 27899
rect 360 27867 400 27899
rect 432 27867 472 27899
rect 504 27867 544 27899
rect 576 27867 616 27899
rect 648 27867 688 27899
rect 720 27867 760 27899
rect 792 27867 832 27899
rect 864 27867 904 27899
rect 936 27867 976 27899
rect 1008 27867 1048 27899
rect 1080 27867 1120 27899
rect 1152 27867 1192 27899
rect 1224 27867 1264 27899
rect 1296 27867 1336 27899
rect 1368 27867 1408 27899
rect 1440 27867 1480 27899
rect 1512 27867 1552 27899
rect 1584 27867 1624 27899
rect 1656 27867 1696 27899
rect 1728 27867 1768 27899
rect 1800 27867 1840 27899
rect 1872 27867 1912 27899
rect 1944 27867 1984 27899
rect 2016 27867 2056 27899
rect 2088 27867 2128 27899
rect 2160 27867 2200 27899
rect 2232 27867 2272 27899
rect 2304 27867 2344 27899
rect 2376 27867 2416 27899
rect 2448 27867 2488 27899
rect 2520 27867 2560 27899
rect 2592 27867 2632 27899
rect 2664 27867 2704 27899
rect 2736 27867 2776 27899
rect 2808 27867 2848 27899
rect 2880 27867 2920 27899
rect 2952 27867 2992 27899
rect 3024 27867 3064 27899
rect 3096 27867 3136 27899
rect 3168 27867 3208 27899
rect 3240 27867 3280 27899
rect 3312 27867 3352 27899
rect 3384 27867 3424 27899
rect 3456 27867 3496 27899
rect 3528 27867 3568 27899
rect 3600 27867 3640 27899
rect 3672 27867 3712 27899
rect 3744 27867 3784 27899
rect 3816 27867 3856 27899
rect 3888 27867 4000 27899
rect 0 27827 4000 27867
rect 0 27795 112 27827
rect 144 27795 184 27827
rect 216 27795 256 27827
rect 288 27795 328 27827
rect 360 27795 400 27827
rect 432 27795 472 27827
rect 504 27795 544 27827
rect 576 27795 616 27827
rect 648 27795 688 27827
rect 720 27795 760 27827
rect 792 27795 832 27827
rect 864 27795 904 27827
rect 936 27795 976 27827
rect 1008 27795 1048 27827
rect 1080 27795 1120 27827
rect 1152 27795 1192 27827
rect 1224 27795 1264 27827
rect 1296 27795 1336 27827
rect 1368 27795 1408 27827
rect 1440 27795 1480 27827
rect 1512 27795 1552 27827
rect 1584 27795 1624 27827
rect 1656 27795 1696 27827
rect 1728 27795 1768 27827
rect 1800 27795 1840 27827
rect 1872 27795 1912 27827
rect 1944 27795 1984 27827
rect 2016 27795 2056 27827
rect 2088 27795 2128 27827
rect 2160 27795 2200 27827
rect 2232 27795 2272 27827
rect 2304 27795 2344 27827
rect 2376 27795 2416 27827
rect 2448 27795 2488 27827
rect 2520 27795 2560 27827
rect 2592 27795 2632 27827
rect 2664 27795 2704 27827
rect 2736 27795 2776 27827
rect 2808 27795 2848 27827
rect 2880 27795 2920 27827
rect 2952 27795 2992 27827
rect 3024 27795 3064 27827
rect 3096 27795 3136 27827
rect 3168 27795 3208 27827
rect 3240 27795 3280 27827
rect 3312 27795 3352 27827
rect 3384 27795 3424 27827
rect 3456 27795 3496 27827
rect 3528 27795 3568 27827
rect 3600 27795 3640 27827
rect 3672 27795 3712 27827
rect 3744 27795 3784 27827
rect 3816 27795 3856 27827
rect 3888 27795 4000 27827
rect 0 27755 4000 27795
rect 0 27723 112 27755
rect 144 27723 184 27755
rect 216 27723 256 27755
rect 288 27723 328 27755
rect 360 27723 400 27755
rect 432 27723 472 27755
rect 504 27723 544 27755
rect 576 27723 616 27755
rect 648 27723 688 27755
rect 720 27723 760 27755
rect 792 27723 832 27755
rect 864 27723 904 27755
rect 936 27723 976 27755
rect 1008 27723 1048 27755
rect 1080 27723 1120 27755
rect 1152 27723 1192 27755
rect 1224 27723 1264 27755
rect 1296 27723 1336 27755
rect 1368 27723 1408 27755
rect 1440 27723 1480 27755
rect 1512 27723 1552 27755
rect 1584 27723 1624 27755
rect 1656 27723 1696 27755
rect 1728 27723 1768 27755
rect 1800 27723 1840 27755
rect 1872 27723 1912 27755
rect 1944 27723 1984 27755
rect 2016 27723 2056 27755
rect 2088 27723 2128 27755
rect 2160 27723 2200 27755
rect 2232 27723 2272 27755
rect 2304 27723 2344 27755
rect 2376 27723 2416 27755
rect 2448 27723 2488 27755
rect 2520 27723 2560 27755
rect 2592 27723 2632 27755
rect 2664 27723 2704 27755
rect 2736 27723 2776 27755
rect 2808 27723 2848 27755
rect 2880 27723 2920 27755
rect 2952 27723 2992 27755
rect 3024 27723 3064 27755
rect 3096 27723 3136 27755
rect 3168 27723 3208 27755
rect 3240 27723 3280 27755
rect 3312 27723 3352 27755
rect 3384 27723 3424 27755
rect 3456 27723 3496 27755
rect 3528 27723 3568 27755
rect 3600 27723 3640 27755
rect 3672 27723 3712 27755
rect 3744 27723 3784 27755
rect 3816 27723 3856 27755
rect 3888 27723 4000 27755
rect 0 27683 4000 27723
rect 0 27651 112 27683
rect 144 27651 184 27683
rect 216 27651 256 27683
rect 288 27651 328 27683
rect 360 27651 400 27683
rect 432 27651 472 27683
rect 504 27651 544 27683
rect 576 27651 616 27683
rect 648 27651 688 27683
rect 720 27651 760 27683
rect 792 27651 832 27683
rect 864 27651 904 27683
rect 936 27651 976 27683
rect 1008 27651 1048 27683
rect 1080 27651 1120 27683
rect 1152 27651 1192 27683
rect 1224 27651 1264 27683
rect 1296 27651 1336 27683
rect 1368 27651 1408 27683
rect 1440 27651 1480 27683
rect 1512 27651 1552 27683
rect 1584 27651 1624 27683
rect 1656 27651 1696 27683
rect 1728 27651 1768 27683
rect 1800 27651 1840 27683
rect 1872 27651 1912 27683
rect 1944 27651 1984 27683
rect 2016 27651 2056 27683
rect 2088 27651 2128 27683
rect 2160 27651 2200 27683
rect 2232 27651 2272 27683
rect 2304 27651 2344 27683
rect 2376 27651 2416 27683
rect 2448 27651 2488 27683
rect 2520 27651 2560 27683
rect 2592 27651 2632 27683
rect 2664 27651 2704 27683
rect 2736 27651 2776 27683
rect 2808 27651 2848 27683
rect 2880 27651 2920 27683
rect 2952 27651 2992 27683
rect 3024 27651 3064 27683
rect 3096 27651 3136 27683
rect 3168 27651 3208 27683
rect 3240 27651 3280 27683
rect 3312 27651 3352 27683
rect 3384 27651 3424 27683
rect 3456 27651 3496 27683
rect 3528 27651 3568 27683
rect 3600 27651 3640 27683
rect 3672 27651 3712 27683
rect 3744 27651 3784 27683
rect 3816 27651 3856 27683
rect 3888 27651 4000 27683
rect 0 27611 4000 27651
rect 0 27579 112 27611
rect 144 27579 184 27611
rect 216 27579 256 27611
rect 288 27579 328 27611
rect 360 27579 400 27611
rect 432 27579 472 27611
rect 504 27579 544 27611
rect 576 27579 616 27611
rect 648 27579 688 27611
rect 720 27579 760 27611
rect 792 27579 832 27611
rect 864 27579 904 27611
rect 936 27579 976 27611
rect 1008 27579 1048 27611
rect 1080 27579 1120 27611
rect 1152 27579 1192 27611
rect 1224 27579 1264 27611
rect 1296 27579 1336 27611
rect 1368 27579 1408 27611
rect 1440 27579 1480 27611
rect 1512 27579 1552 27611
rect 1584 27579 1624 27611
rect 1656 27579 1696 27611
rect 1728 27579 1768 27611
rect 1800 27579 1840 27611
rect 1872 27579 1912 27611
rect 1944 27579 1984 27611
rect 2016 27579 2056 27611
rect 2088 27579 2128 27611
rect 2160 27579 2200 27611
rect 2232 27579 2272 27611
rect 2304 27579 2344 27611
rect 2376 27579 2416 27611
rect 2448 27579 2488 27611
rect 2520 27579 2560 27611
rect 2592 27579 2632 27611
rect 2664 27579 2704 27611
rect 2736 27579 2776 27611
rect 2808 27579 2848 27611
rect 2880 27579 2920 27611
rect 2952 27579 2992 27611
rect 3024 27579 3064 27611
rect 3096 27579 3136 27611
rect 3168 27579 3208 27611
rect 3240 27579 3280 27611
rect 3312 27579 3352 27611
rect 3384 27579 3424 27611
rect 3456 27579 3496 27611
rect 3528 27579 3568 27611
rect 3600 27579 3640 27611
rect 3672 27579 3712 27611
rect 3744 27579 3784 27611
rect 3816 27579 3856 27611
rect 3888 27579 4000 27611
rect 0 27539 4000 27579
rect 0 27507 112 27539
rect 144 27507 184 27539
rect 216 27507 256 27539
rect 288 27507 328 27539
rect 360 27507 400 27539
rect 432 27507 472 27539
rect 504 27507 544 27539
rect 576 27507 616 27539
rect 648 27507 688 27539
rect 720 27507 760 27539
rect 792 27507 832 27539
rect 864 27507 904 27539
rect 936 27507 976 27539
rect 1008 27507 1048 27539
rect 1080 27507 1120 27539
rect 1152 27507 1192 27539
rect 1224 27507 1264 27539
rect 1296 27507 1336 27539
rect 1368 27507 1408 27539
rect 1440 27507 1480 27539
rect 1512 27507 1552 27539
rect 1584 27507 1624 27539
rect 1656 27507 1696 27539
rect 1728 27507 1768 27539
rect 1800 27507 1840 27539
rect 1872 27507 1912 27539
rect 1944 27507 1984 27539
rect 2016 27507 2056 27539
rect 2088 27507 2128 27539
rect 2160 27507 2200 27539
rect 2232 27507 2272 27539
rect 2304 27507 2344 27539
rect 2376 27507 2416 27539
rect 2448 27507 2488 27539
rect 2520 27507 2560 27539
rect 2592 27507 2632 27539
rect 2664 27507 2704 27539
rect 2736 27507 2776 27539
rect 2808 27507 2848 27539
rect 2880 27507 2920 27539
rect 2952 27507 2992 27539
rect 3024 27507 3064 27539
rect 3096 27507 3136 27539
rect 3168 27507 3208 27539
rect 3240 27507 3280 27539
rect 3312 27507 3352 27539
rect 3384 27507 3424 27539
rect 3456 27507 3496 27539
rect 3528 27507 3568 27539
rect 3600 27507 3640 27539
rect 3672 27507 3712 27539
rect 3744 27507 3784 27539
rect 3816 27507 3856 27539
rect 3888 27507 4000 27539
rect 0 27467 4000 27507
rect 0 27435 112 27467
rect 144 27435 184 27467
rect 216 27435 256 27467
rect 288 27435 328 27467
rect 360 27435 400 27467
rect 432 27435 472 27467
rect 504 27435 544 27467
rect 576 27435 616 27467
rect 648 27435 688 27467
rect 720 27435 760 27467
rect 792 27435 832 27467
rect 864 27435 904 27467
rect 936 27435 976 27467
rect 1008 27435 1048 27467
rect 1080 27435 1120 27467
rect 1152 27435 1192 27467
rect 1224 27435 1264 27467
rect 1296 27435 1336 27467
rect 1368 27435 1408 27467
rect 1440 27435 1480 27467
rect 1512 27435 1552 27467
rect 1584 27435 1624 27467
rect 1656 27435 1696 27467
rect 1728 27435 1768 27467
rect 1800 27435 1840 27467
rect 1872 27435 1912 27467
rect 1944 27435 1984 27467
rect 2016 27435 2056 27467
rect 2088 27435 2128 27467
rect 2160 27435 2200 27467
rect 2232 27435 2272 27467
rect 2304 27435 2344 27467
rect 2376 27435 2416 27467
rect 2448 27435 2488 27467
rect 2520 27435 2560 27467
rect 2592 27435 2632 27467
rect 2664 27435 2704 27467
rect 2736 27435 2776 27467
rect 2808 27435 2848 27467
rect 2880 27435 2920 27467
rect 2952 27435 2992 27467
rect 3024 27435 3064 27467
rect 3096 27435 3136 27467
rect 3168 27435 3208 27467
rect 3240 27435 3280 27467
rect 3312 27435 3352 27467
rect 3384 27435 3424 27467
rect 3456 27435 3496 27467
rect 3528 27435 3568 27467
rect 3600 27435 3640 27467
rect 3672 27435 3712 27467
rect 3744 27435 3784 27467
rect 3816 27435 3856 27467
rect 3888 27435 4000 27467
rect 0 27395 4000 27435
rect 0 27363 112 27395
rect 144 27363 184 27395
rect 216 27363 256 27395
rect 288 27363 328 27395
rect 360 27363 400 27395
rect 432 27363 472 27395
rect 504 27363 544 27395
rect 576 27363 616 27395
rect 648 27363 688 27395
rect 720 27363 760 27395
rect 792 27363 832 27395
rect 864 27363 904 27395
rect 936 27363 976 27395
rect 1008 27363 1048 27395
rect 1080 27363 1120 27395
rect 1152 27363 1192 27395
rect 1224 27363 1264 27395
rect 1296 27363 1336 27395
rect 1368 27363 1408 27395
rect 1440 27363 1480 27395
rect 1512 27363 1552 27395
rect 1584 27363 1624 27395
rect 1656 27363 1696 27395
rect 1728 27363 1768 27395
rect 1800 27363 1840 27395
rect 1872 27363 1912 27395
rect 1944 27363 1984 27395
rect 2016 27363 2056 27395
rect 2088 27363 2128 27395
rect 2160 27363 2200 27395
rect 2232 27363 2272 27395
rect 2304 27363 2344 27395
rect 2376 27363 2416 27395
rect 2448 27363 2488 27395
rect 2520 27363 2560 27395
rect 2592 27363 2632 27395
rect 2664 27363 2704 27395
rect 2736 27363 2776 27395
rect 2808 27363 2848 27395
rect 2880 27363 2920 27395
rect 2952 27363 2992 27395
rect 3024 27363 3064 27395
rect 3096 27363 3136 27395
rect 3168 27363 3208 27395
rect 3240 27363 3280 27395
rect 3312 27363 3352 27395
rect 3384 27363 3424 27395
rect 3456 27363 3496 27395
rect 3528 27363 3568 27395
rect 3600 27363 3640 27395
rect 3672 27363 3712 27395
rect 3744 27363 3784 27395
rect 3816 27363 3856 27395
rect 3888 27363 4000 27395
rect 0 27323 4000 27363
rect 0 27291 112 27323
rect 144 27291 184 27323
rect 216 27291 256 27323
rect 288 27291 328 27323
rect 360 27291 400 27323
rect 432 27291 472 27323
rect 504 27291 544 27323
rect 576 27291 616 27323
rect 648 27291 688 27323
rect 720 27291 760 27323
rect 792 27291 832 27323
rect 864 27291 904 27323
rect 936 27291 976 27323
rect 1008 27291 1048 27323
rect 1080 27291 1120 27323
rect 1152 27291 1192 27323
rect 1224 27291 1264 27323
rect 1296 27291 1336 27323
rect 1368 27291 1408 27323
rect 1440 27291 1480 27323
rect 1512 27291 1552 27323
rect 1584 27291 1624 27323
rect 1656 27291 1696 27323
rect 1728 27291 1768 27323
rect 1800 27291 1840 27323
rect 1872 27291 1912 27323
rect 1944 27291 1984 27323
rect 2016 27291 2056 27323
rect 2088 27291 2128 27323
rect 2160 27291 2200 27323
rect 2232 27291 2272 27323
rect 2304 27291 2344 27323
rect 2376 27291 2416 27323
rect 2448 27291 2488 27323
rect 2520 27291 2560 27323
rect 2592 27291 2632 27323
rect 2664 27291 2704 27323
rect 2736 27291 2776 27323
rect 2808 27291 2848 27323
rect 2880 27291 2920 27323
rect 2952 27291 2992 27323
rect 3024 27291 3064 27323
rect 3096 27291 3136 27323
rect 3168 27291 3208 27323
rect 3240 27291 3280 27323
rect 3312 27291 3352 27323
rect 3384 27291 3424 27323
rect 3456 27291 3496 27323
rect 3528 27291 3568 27323
rect 3600 27291 3640 27323
rect 3672 27291 3712 27323
rect 3744 27291 3784 27323
rect 3816 27291 3856 27323
rect 3888 27291 4000 27323
rect 0 27251 4000 27291
rect 0 27219 112 27251
rect 144 27219 184 27251
rect 216 27219 256 27251
rect 288 27219 328 27251
rect 360 27219 400 27251
rect 432 27219 472 27251
rect 504 27219 544 27251
rect 576 27219 616 27251
rect 648 27219 688 27251
rect 720 27219 760 27251
rect 792 27219 832 27251
rect 864 27219 904 27251
rect 936 27219 976 27251
rect 1008 27219 1048 27251
rect 1080 27219 1120 27251
rect 1152 27219 1192 27251
rect 1224 27219 1264 27251
rect 1296 27219 1336 27251
rect 1368 27219 1408 27251
rect 1440 27219 1480 27251
rect 1512 27219 1552 27251
rect 1584 27219 1624 27251
rect 1656 27219 1696 27251
rect 1728 27219 1768 27251
rect 1800 27219 1840 27251
rect 1872 27219 1912 27251
rect 1944 27219 1984 27251
rect 2016 27219 2056 27251
rect 2088 27219 2128 27251
rect 2160 27219 2200 27251
rect 2232 27219 2272 27251
rect 2304 27219 2344 27251
rect 2376 27219 2416 27251
rect 2448 27219 2488 27251
rect 2520 27219 2560 27251
rect 2592 27219 2632 27251
rect 2664 27219 2704 27251
rect 2736 27219 2776 27251
rect 2808 27219 2848 27251
rect 2880 27219 2920 27251
rect 2952 27219 2992 27251
rect 3024 27219 3064 27251
rect 3096 27219 3136 27251
rect 3168 27219 3208 27251
rect 3240 27219 3280 27251
rect 3312 27219 3352 27251
rect 3384 27219 3424 27251
rect 3456 27219 3496 27251
rect 3528 27219 3568 27251
rect 3600 27219 3640 27251
rect 3672 27219 3712 27251
rect 3744 27219 3784 27251
rect 3816 27219 3856 27251
rect 3888 27219 4000 27251
rect 0 27179 4000 27219
rect 0 27147 112 27179
rect 144 27147 184 27179
rect 216 27147 256 27179
rect 288 27147 328 27179
rect 360 27147 400 27179
rect 432 27147 472 27179
rect 504 27147 544 27179
rect 576 27147 616 27179
rect 648 27147 688 27179
rect 720 27147 760 27179
rect 792 27147 832 27179
rect 864 27147 904 27179
rect 936 27147 976 27179
rect 1008 27147 1048 27179
rect 1080 27147 1120 27179
rect 1152 27147 1192 27179
rect 1224 27147 1264 27179
rect 1296 27147 1336 27179
rect 1368 27147 1408 27179
rect 1440 27147 1480 27179
rect 1512 27147 1552 27179
rect 1584 27147 1624 27179
rect 1656 27147 1696 27179
rect 1728 27147 1768 27179
rect 1800 27147 1840 27179
rect 1872 27147 1912 27179
rect 1944 27147 1984 27179
rect 2016 27147 2056 27179
rect 2088 27147 2128 27179
rect 2160 27147 2200 27179
rect 2232 27147 2272 27179
rect 2304 27147 2344 27179
rect 2376 27147 2416 27179
rect 2448 27147 2488 27179
rect 2520 27147 2560 27179
rect 2592 27147 2632 27179
rect 2664 27147 2704 27179
rect 2736 27147 2776 27179
rect 2808 27147 2848 27179
rect 2880 27147 2920 27179
rect 2952 27147 2992 27179
rect 3024 27147 3064 27179
rect 3096 27147 3136 27179
rect 3168 27147 3208 27179
rect 3240 27147 3280 27179
rect 3312 27147 3352 27179
rect 3384 27147 3424 27179
rect 3456 27147 3496 27179
rect 3528 27147 3568 27179
rect 3600 27147 3640 27179
rect 3672 27147 3712 27179
rect 3744 27147 3784 27179
rect 3816 27147 3856 27179
rect 3888 27147 4000 27179
rect 0 27107 4000 27147
rect 0 27075 112 27107
rect 144 27075 184 27107
rect 216 27075 256 27107
rect 288 27075 328 27107
rect 360 27075 400 27107
rect 432 27075 472 27107
rect 504 27075 544 27107
rect 576 27075 616 27107
rect 648 27075 688 27107
rect 720 27075 760 27107
rect 792 27075 832 27107
rect 864 27075 904 27107
rect 936 27075 976 27107
rect 1008 27075 1048 27107
rect 1080 27075 1120 27107
rect 1152 27075 1192 27107
rect 1224 27075 1264 27107
rect 1296 27075 1336 27107
rect 1368 27075 1408 27107
rect 1440 27075 1480 27107
rect 1512 27075 1552 27107
rect 1584 27075 1624 27107
rect 1656 27075 1696 27107
rect 1728 27075 1768 27107
rect 1800 27075 1840 27107
rect 1872 27075 1912 27107
rect 1944 27075 1984 27107
rect 2016 27075 2056 27107
rect 2088 27075 2128 27107
rect 2160 27075 2200 27107
rect 2232 27075 2272 27107
rect 2304 27075 2344 27107
rect 2376 27075 2416 27107
rect 2448 27075 2488 27107
rect 2520 27075 2560 27107
rect 2592 27075 2632 27107
rect 2664 27075 2704 27107
rect 2736 27075 2776 27107
rect 2808 27075 2848 27107
rect 2880 27075 2920 27107
rect 2952 27075 2992 27107
rect 3024 27075 3064 27107
rect 3096 27075 3136 27107
rect 3168 27075 3208 27107
rect 3240 27075 3280 27107
rect 3312 27075 3352 27107
rect 3384 27075 3424 27107
rect 3456 27075 3496 27107
rect 3528 27075 3568 27107
rect 3600 27075 3640 27107
rect 3672 27075 3712 27107
rect 3744 27075 3784 27107
rect 3816 27075 3856 27107
rect 3888 27075 4000 27107
rect 0 27035 4000 27075
rect 0 27003 112 27035
rect 144 27003 184 27035
rect 216 27003 256 27035
rect 288 27003 328 27035
rect 360 27003 400 27035
rect 432 27003 472 27035
rect 504 27003 544 27035
rect 576 27003 616 27035
rect 648 27003 688 27035
rect 720 27003 760 27035
rect 792 27003 832 27035
rect 864 27003 904 27035
rect 936 27003 976 27035
rect 1008 27003 1048 27035
rect 1080 27003 1120 27035
rect 1152 27003 1192 27035
rect 1224 27003 1264 27035
rect 1296 27003 1336 27035
rect 1368 27003 1408 27035
rect 1440 27003 1480 27035
rect 1512 27003 1552 27035
rect 1584 27003 1624 27035
rect 1656 27003 1696 27035
rect 1728 27003 1768 27035
rect 1800 27003 1840 27035
rect 1872 27003 1912 27035
rect 1944 27003 1984 27035
rect 2016 27003 2056 27035
rect 2088 27003 2128 27035
rect 2160 27003 2200 27035
rect 2232 27003 2272 27035
rect 2304 27003 2344 27035
rect 2376 27003 2416 27035
rect 2448 27003 2488 27035
rect 2520 27003 2560 27035
rect 2592 27003 2632 27035
rect 2664 27003 2704 27035
rect 2736 27003 2776 27035
rect 2808 27003 2848 27035
rect 2880 27003 2920 27035
rect 2952 27003 2992 27035
rect 3024 27003 3064 27035
rect 3096 27003 3136 27035
rect 3168 27003 3208 27035
rect 3240 27003 3280 27035
rect 3312 27003 3352 27035
rect 3384 27003 3424 27035
rect 3456 27003 3496 27035
rect 3528 27003 3568 27035
rect 3600 27003 3640 27035
rect 3672 27003 3712 27035
rect 3744 27003 3784 27035
rect 3816 27003 3856 27035
rect 3888 27003 4000 27035
rect 0 26963 4000 27003
rect 0 26931 112 26963
rect 144 26931 184 26963
rect 216 26931 256 26963
rect 288 26931 328 26963
rect 360 26931 400 26963
rect 432 26931 472 26963
rect 504 26931 544 26963
rect 576 26931 616 26963
rect 648 26931 688 26963
rect 720 26931 760 26963
rect 792 26931 832 26963
rect 864 26931 904 26963
rect 936 26931 976 26963
rect 1008 26931 1048 26963
rect 1080 26931 1120 26963
rect 1152 26931 1192 26963
rect 1224 26931 1264 26963
rect 1296 26931 1336 26963
rect 1368 26931 1408 26963
rect 1440 26931 1480 26963
rect 1512 26931 1552 26963
rect 1584 26931 1624 26963
rect 1656 26931 1696 26963
rect 1728 26931 1768 26963
rect 1800 26931 1840 26963
rect 1872 26931 1912 26963
rect 1944 26931 1984 26963
rect 2016 26931 2056 26963
rect 2088 26931 2128 26963
rect 2160 26931 2200 26963
rect 2232 26931 2272 26963
rect 2304 26931 2344 26963
rect 2376 26931 2416 26963
rect 2448 26931 2488 26963
rect 2520 26931 2560 26963
rect 2592 26931 2632 26963
rect 2664 26931 2704 26963
rect 2736 26931 2776 26963
rect 2808 26931 2848 26963
rect 2880 26931 2920 26963
rect 2952 26931 2992 26963
rect 3024 26931 3064 26963
rect 3096 26931 3136 26963
rect 3168 26931 3208 26963
rect 3240 26931 3280 26963
rect 3312 26931 3352 26963
rect 3384 26931 3424 26963
rect 3456 26931 3496 26963
rect 3528 26931 3568 26963
rect 3600 26931 3640 26963
rect 3672 26931 3712 26963
rect 3744 26931 3784 26963
rect 3816 26931 3856 26963
rect 3888 26931 4000 26963
rect 0 26891 4000 26931
rect 0 26859 112 26891
rect 144 26859 184 26891
rect 216 26859 256 26891
rect 288 26859 328 26891
rect 360 26859 400 26891
rect 432 26859 472 26891
rect 504 26859 544 26891
rect 576 26859 616 26891
rect 648 26859 688 26891
rect 720 26859 760 26891
rect 792 26859 832 26891
rect 864 26859 904 26891
rect 936 26859 976 26891
rect 1008 26859 1048 26891
rect 1080 26859 1120 26891
rect 1152 26859 1192 26891
rect 1224 26859 1264 26891
rect 1296 26859 1336 26891
rect 1368 26859 1408 26891
rect 1440 26859 1480 26891
rect 1512 26859 1552 26891
rect 1584 26859 1624 26891
rect 1656 26859 1696 26891
rect 1728 26859 1768 26891
rect 1800 26859 1840 26891
rect 1872 26859 1912 26891
rect 1944 26859 1984 26891
rect 2016 26859 2056 26891
rect 2088 26859 2128 26891
rect 2160 26859 2200 26891
rect 2232 26859 2272 26891
rect 2304 26859 2344 26891
rect 2376 26859 2416 26891
rect 2448 26859 2488 26891
rect 2520 26859 2560 26891
rect 2592 26859 2632 26891
rect 2664 26859 2704 26891
rect 2736 26859 2776 26891
rect 2808 26859 2848 26891
rect 2880 26859 2920 26891
rect 2952 26859 2992 26891
rect 3024 26859 3064 26891
rect 3096 26859 3136 26891
rect 3168 26859 3208 26891
rect 3240 26859 3280 26891
rect 3312 26859 3352 26891
rect 3384 26859 3424 26891
rect 3456 26859 3496 26891
rect 3528 26859 3568 26891
rect 3600 26859 3640 26891
rect 3672 26859 3712 26891
rect 3744 26859 3784 26891
rect 3816 26859 3856 26891
rect 3888 26859 4000 26891
rect 0 26819 4000 26859
rect 0 26787 112 26819
rect 144 26787 184 26819
rect 216 26787 256 26819
rect 288 26787 328 26819
rect 360 26787 400 26819
rect 432 26787 472 26819
rect 504 26787 544 26819
rect 576 26787 616 26819
rect 648 26787 688 26819
rect 720 26787 760 26819
rect 792 26787 832 26819
rect 864 26787 904 26819
rect 936 26787 976 26819
rect 1008 26787 1048 26819
rect 1080 26787 1120 26819
rect 1152 26787 1192 26819
rect 1224 26787 1264 26819
rect 1296 26787 1336 26819
rect 1368 26787 1408 26819
rect 1440 26787 1480 26819
rect 1512 26787 1552 26819
rect 1584 26787 1624 26819
rect 1656 26787 1696 26819
rect 1728 26787 1768 26819
rect 1800 26787 1840 26819
rect 1872 26787 1912 26819
rect 1944 26787 1984 26819
rect 2016 26787 2056 26819
rect 2088 26787 2128 26819
rect 2160 26787 2200 26819
rect 2232 26787 2272 26819
rect 2304 26787 2344 26819
rect 2376 26787 2416 26819
rect 2448 26787 2488 26819
rect 2520 26787 2560 26819
rect 2592 26787 2632 26819
rect 2664 26787 2704 26819
rect 2736 26787 2776 26819
rect 2808 26787 2848 26819
rect 2880 26787 2920 26819
rect 2952 26787 2992 26819
rect 3024 26787 3064 26819
rect 3096 26787 3136 26819
rect 3168 26787 3208 26819
rect 3240 26787 3280 26819
rect 3312 26787 3352 26819
rect 3384 26787 3424 26819
rect 3456 26787 3496 26819
rect 3528 26787 3568 26819
rect 3600 26787 3640 26819
rect 3672 26787 3712 26819
rect 3744 26787 3784 26819
rect 3816 26787 3856 26819
rect 3888 26787 4000 26819
rect 0 26747 4000 26787
rect 0 26715 112 26747
rect 144 26715 184 26747
rect 216 26715 256 26747
rect 288 26715 328 26747
rect 360 26715 400 26747
rect 432 26715 472 26747
rect 504 26715 544 26747
rect 576 26715 616 26747
rect 648 26715 688 26747
rect 720 26715 760 26747
rect 792 26715 832 26747
rect 864 26715 904 26747
rect 936 26715 976 26747
rect 1008 26715 1048 26747
rect 1080 26715 1120 26747
rect 1152 26715 1192 26747
rect 1224 26715 1264 26747
rect 1296 26715 1336 26747
rect 1368 26715 1408 26747
rect 1440 26715 1480 26747
rect 1512 26715 1552 26747
rect 1584 26715 1624 26747
rect 1656 26715 1696 26747
rect 1728 26715 1768 26747
rect 1800 26715 1840 26747
rect 1872 26715 1912 26747
rect 1944 26715 1984 26747
rect 2016 26715 2056 26747
rect 2088 26715 2128 26747
rect 2160 26715 2200 26747
rect 2232 26715 2272 26747
rect 2304 26715 2344 26747
rect 2376 26715 2416 26747
rect 2448 26715 2488 26747
rect 2520 26715 2560 26747
rect 2592 26715 2632 26747
rect 2664 26715 2704 26747
rect 2736 26715 2776 26747
rect 2808 26715 2848 26747
rect 2880 26715 2920 26747
rect 2952 26715 2992 26747
rect 3024 26715 3064 26747
rect 3096 26715 3136 26747
rect 3168 26715 3208 26747
rect 3240 26715 3280 26747
rect 3312 26715 3352 26747
rect 3384 26715 3424 26747
rect 3456 26715 3496 26747
rect 3528 26715 3568 26747
rect 3600 26715 3640 26747
rect 3672 26715 3712 26747
rect 3744 26715 3784 26747
rect 3816 26715 3856 26747
rect 3888 26715 4000 26747
rect 0 26675 4000 26715
rect 0 26643 112 26675
rect 144 26643 184 26675
rect 216 26643 256 26675
rect 288 26643 328 26675
rect 360 26643 400 26675
rect 432 26643 472 26675
rect 504 26643 544 26675
rect 576 26643 616 26675
rect 648 26643 688 26675
rect 720 26643 760 26675
rect 792 26643 832 26675
rect 864 26643 904 26675
rect 936 26643 976 26675
rect 1008 26643 1048 26675
rect 1080 26643 1120 26675
rect 1152 26643 1192 26675
rect 1224 26643 1264 26675
rect 1296 26643 1336 26675
rect 1368 26643 1408 26675
rect 1440 26643 1480 26675
rect 1512 26643 1552 26675
rect 1584 26643 1624 26675
rect 1656 26643 1696 26675
rect 1728 26643 1768 26675
rect 1800 26643 1840 26675
rect 1872 26643 1912 26675
rect 1944 26643 1984 26675
rect 2016 26643 2056 26675
rect 2088 26643 2128 26675
rect 2160 26643 2200 26675
rect 2232 26643 2272 26675
rect 2304 26643 2344 26675
rect 2376 26643 2416 26675
rect 2448 26643 2488 26675
rect 2520 26643 2560 26675
rect 2592 26643 2632 26675
rect 2664 26643 2704 26675
rect 2736 26643 2776 26675
rect 2808 26643 2848 26675
rect 2880 26643 2920 26675
rect 2952 26643 2992 26675
rect 3024 26643 3064 26675
rect 3096 26643 3136 26675
rect 3168 26643 3208 26675
rect 3240 26643 3280 26675
rect 3312 26643 3352 26675
rect 3384 26643 3424 26675
rect 3456 26643 3496 26675
rect 3528 26643 3568 26675
rect 3600 26643 3640 26675
rect 3672 26643 3712 26675
rect 3744 26643 3784 26675
rect 3816 26643 3856 26675
rect 3888 26643 4000 26675
rect 0 26603 4000 26643
rect 0 26571 112 26603
rect 144 26571 184 26603
rect 216 26571 256 26603
rect 288 26571 328 26603
rect 360 26571 400 26603
rect 432 26571 472 26603
rect 504 26571 544 26603
rect 576 26571 616 26603
rect 648 26571 688 26603
rect 720 26571 760 26603
rect 792 26571 832 26603
rect 864 26571 904 26603
rect 936 26571 976 26603
rect 1008 26571 1048 26603
rect 1080 26571 1120 26603
rect 1152 26571 1192 26603
rect 1224 26571 1264 26603
rect 1296 26571 1336 26603
rect 1368 26571 1408 26603
rect 1440 26571 1480 26603
rect 1512 26571 1552 26603
rect 1584 26571 1624 26603
rect 1656 26571 1696 26603
rect 1728 26571 1768 26603
rect 1800 26571 1840 26603
rect 1872 26571 1912 26603
rect 1944 26571 1984 26603
rect 2016 26571 2056 26603
rect 2088 26571 2128 26603
rect 2160 26571 2200 26603
rect 2232 26571 2272 26603
rect 2304 26571 2344 26603
rect 2376 26571 2416 26603
rect 2448 26571 2488 26603
rect 2520 26571 2560 26603
rect 2592 26571 2632 26603
rect 2664 26571 2704 26603
rect 2736 26571 2776 26603
rect 2808 26571 2848 26603
rect 2880 26571 2920 26603
rect 2952 26571 2992 26603
rect 3024 26571 3064 26603
rect 3096 26571 3136 26603
rect 3168 26571 3208 26603
rect 3240 26571 3280 26603
rect 3312 26571 3352 26603
rect 3384 26571 3424 26603
rect 3456 26571 3496 26603
rect 3528 26571 3568 26603
rect 3600 26571 3640 26603
rect 3672 26571 3712 26603
rect 3744 26571 3784 26603
rect 3816 26571 3856 26603
rect 3888 26571 4000 26603
rect 0 26531 4000 26571
rect 0 26499 112 26531
rect 144 26499 184 26531
rect 216 26499 256 26531
rect 288 26499 328 26531
rect 360 26499 400 26531
rect 432 26499 472 26531
rect 504 26499 544 26531
rect 576 26499 616 26531
rect 648 26499 688 26531
rect 720 26499 760 26531
rect 792 26499 832 26531
rect 864 26499 904 26531
rect 936 26499 976 26531
rect 1008 26499 1048 26531
rect 1080 26499 1120 26531
rect 1152 26499 1192 26531
rect 1224 26499 1264 26531
rect 1296 26499 1336 26531
rect 1368 26499 1408 26531
rect 1440 26499 1480 26531
rect 1512 26499 1552 26531
rect 1584 26499 1624 26531
rect 1656 26499 1696 26531
rect 1728 26499 1768 26531
rect 1800 26499 1840 26531
rect 1872 26499 1912 26531
rect 1944 26499 1984 26531
rect 2016 26499 2056 26531
rect 2088 26499 2128 26531
rect 2160 26499 2200 26531
rect 2232 26499 2272 26531
rect 2304 26499 2344 26531
rect 2376 26499 2416 26531
rect 2448 26499 2488 26531
rect 2520 26499 2560 26531
rect 2592 26499 2632 26531
rect 2664 26499 2704 26531
rect 2736 26499 2776 26531
rect 2808 26499 2848 26531
rect 2880 26499 2920 26531
rect 2952 26499 2992 26531
rect 3024 26499 3064 26531
rect 3096 26499 3136 26531
rect 3168 26499 3208 26531
rect 3240 26499 3280 26531
rect 3312 26499 3352 26531
rect 3384 26499 3424 26531
rect 3456 26499 3496 26531
rect 3528 26499 3568 26531
rect 3600 26499 3640 26531
rect 3672 26499 3712 26531
rect 3744 26499 3784 26531
rect 3816 26499 3856 26531
rect 3888 26499 4000 26531
rect 0 26459 4000 26499
rect 0 26427 112 26459
rect 144 26427 184 26459
rect 216 26427 256 26459
rect 288 26427 328 26459
rect 360 26427 400 26459
rect 432 26427 472 26459
rect 504 26427 544 26459
rect 576 26427 616 26459
rect 648 26427 688 26459
rect 720 26427 760 26459
rect 792 26427 832 26459
rect 864 26427 904 26459
rect 936 26427 976 26459
rect 1008 26427 1048 26459
rect 1080 26427 1120 26459
rect 1152 26427 1192 26459
rect 1224 26427 1264 26459
rect 1296 26427 1336 26459
rect 1368 26427 1408 26459
rect 1440 26427 1480 26459
rect 1512 26427 1552 26459
rect 1584 26427 1624 26459
rect 1656 26427 1696 26459
rect 1728 26427 1768 26459
rect 1800 26427 1840 26459
rect 1872 26427 1912 26459
rect 1944 26427 1984 26459
rect 2016 26427 2056 26459
rect 2088 26427 2128 26459
rect 2160 26427 2200 26459
rect 2232 26427 2272 26459
rect 2304 26427 2344 26459
rect 2376 26427 2416 26459
rect 2448 26427 2488 26459
rect 2520 26427 2560 26459
rect 2592 26427 2632 26459
rect 2664 26427 2704 26459
rect 2736 26427 2776 26459
rect 2808 26427 2848 26459
rect 2880 26427 2920 26459
rect 2952 26427 2992 26459
rect 3024 26427 3064 26459
rect 3096 26427 3136 26459
rect 3168 26427 3208 26459
rect 3240 26427 3280 26459
rect 3312 26427 3352 26459
rect 3384 26427 3424 26459
rect 3456 26427 3496 26459
rect 3528 26427 3568 26459
rect 3600 26427 3640 26459
rect 3672 26427 3712 26459
rect 3744 26427 3784 26459
rect 3816 26427 3856 26459
rect 3888 26427 4000 26459
rect 0 26387 4000 26427
rect 0 26355 112 26387
rect 144 26355 184 26387
rect 216 26355 256 26387
rect 288 26355 328 26387
rect 360 26355 400 26387
rect 432 26355 472 26387
rect 504 26355 544 26387
rect 576 26355 616 26387
rect 648 26355 688 26387
rect 720 26355 760 26387
rect 792 26355 832 26387
rect 864 26355 904 26387
rect 936 26355 976 26387
rect 1008 26355 1048 26387
rect 1080 26355 1120 26387
rect 1152 26355 1192 26387
rect 1224 26355 1264 26387
rect 1296 26355 1336 26387
rect 1368 26355 1408 26387
rect 1440 26355 1480 26387
rect 1512 26355 1552 26387
rect 1584 26355 1624 26387
rect 1656 26355 1696 26387
rect 1728 26355 1768 26387
rect 1800 26355 1840 26387
rect 1872 26355 1912 26387
rect 1944 26355 1984 26387
rect 2016 26355 2056 26387
rect 2088 26355 2128 26387
rect 2160 26355 2200 26387
rect 2232 26355 2272 26387
rect 2304 26355 2344 26387
rect 2376 26355 2416 26387
rect 2448 26355 2488 26387
rect 2520 26355 2560 26387
rect 2592 26355 2632 26387
rect 2664 26355 2704 26387
rect 2736 26355 2776 26387
rect 2808 26355 2848 26387
rect 2880 26355 2920 26387
rect 2952 26355 2992 26387
rect 3024 26355 3064 26387
rect 3096 26355 3136 26387
rect 3168 26355 3208 26387
rect 3240 26355 3280 26387
rect 3312 26355 3352 26387
rect 3384 26355 3424 26387
rect 3456 26355 3496 26387
rect 3528 26355 3568 26387
rect 3600 26355 3640 26387
rect 3672 26355 3712 26387
rect 3744 26355 3784 26387
rect 3816 26355 3856 26387
rect 3888 26355 4000 26387
rect 0 26315 4000 26355
rect 0 26283 112 26315
rect 144 26283 184 26315
rect 216 26283 256 26315
rect 288 26283 328 26315
rect 360 26283 400 26315
rect 432 26283 472 26315
rect 504 26283 544 26315
rect 576 26283 616 26315
rect 648 26283 688 26315
rect 720 26283 760 26315
rect 792 26283 832 26315
rect 864 26283 904 26315
rect 936 26283 976 26315
rect 1008 26283 1048 26315
rect 1080 26283 1120 26315
rect 1152 26283 1192 26315
rect 1224 26283 1264 26315
rect 1296 26283 1336 26315
rect 1368 26283 1408 26315
rect 1440 26283 1480 26315
rect 1512 26283 1552 26315
rect 1584 26283 1624 26315
rect 1656 26283 1696 26315
rect 1728 26283 1768 26315
rect 1800 26283 1840 26315
rect 1872 26283 1912 26315
rect 1944 26283 1984 26315
rect 2016 26283 2056 26315
rect 2088 26283 2128 26315
rect 2160 26283 2200 26315
rect 2232 26283 2272 26315
rect 2304 26283 2344 26315
rect 2376 26283 2416 26315
rect 2448 26283 2488 26315
rect 2520 26283 2560 26315
rect 2592 26283 2632 26315
rect 2664 26283 2704 26315
rect 2736 26283 2776 26315
rect 2808 26283 2848 26315
rect 2880 26283 2920 26315
rect 2952 26283 2992 26315
rect 3024 26283 3064 26315
rect 3096 26283 3136 26315
rect 3168 26283 3208 26315
rect 3240 26283 3280 26315
rect 3312 26283 3352 26315
rect 3384 26283 3424 26315
rect 3456 26283 3496 26315
rect 3528 26283 3568 26315
rect 3600 26283 3640 26315
rect 3672 26283 3712 26315
rect 3744 26283 3784 26315
rect 3816 26283 3856 26315
rect 3888 26283 4000 26315
rect 0 26243 4000 26283
rect 0 26211 112 26243
rect 144 26211 184 26243
rect 216 26211 256 26243
rect 288 26211 328 26243
rect 360 26211 400 26243
rect 432 26211 472 26243
rect 504 26211 544 26243
rect 576 26211 616 26243
rect 648 26211 688 26243
rect 720 26211 760 26243
rect 792 26211 832 26243
rect 864 26211 904 26243
rect 936 26211 976 26243
rect 1008 26211 1048 26243
rect 1080 26211 1120 26243
rect 1152 26211 1192 26243
rect 1224 26211 1264 26243
rect 1296 26211 1336 26243
rect 1368 26211 1408 26243
rect 1440 26211 1480 26243
rect 1512 26211 1552 26243
rect 1584 26211 1624 26243
rect 1656 26211 1696 26243
rect 1728 26211 1768 26243
rect 1800 26211 1840 26243
rect 1872 26211 1912 26243
rect 1944 26211 1984 26243
rect 2016 26211 2056 26243
rect 2088 26211 2128 26243
rect 2160 26211 2200 26243
rect 2232 26211 2272 26243
rect 2304 26211 2344 26243
rect 2376 26211 2416 26243
rect 2448 26211 2488 26243
rect 2520 26211 2560 26243
rect 2592 26211 2632 26243
rect 2664 26211 2704 26243
rect 2736 26211 2776 26243
rect 2808 26211 2848 26243
rect 2880 26211 2920 26243
rect 2952 26211 2992 26243
rect 3024 26211 3064 26243
rect 3096 26211 3136 26243
rect 3168 26211 3208 26243
rect 3240 26211 3280 26243
rect 3312 26211 3352 26243
rect 3384 26211 3424 26243
rect 3456 26211 3496 26243
rect 3528 26211 3568 26243
rect 3600 26211 3640 26243
rect 3672 26211 3712 26243
rect 3744 26211 3784 26243
rect 3816 26211 3856 26243
rect 3888 26211 4000 26243
rect 0 26171 4000 26211
rect 0 26139 112 26171
rect 144 26139 184 26171
rect 216 26139 256 26171
rect 288 26139 328 26171
rect 360 26139 400 26171
rect 432 26139 472 26171
rect 504 26139 544 26171
rect 576 26139 616 26171
rect 648 26139 688 26171
rect 720 26139 760 26171
rect 792 26139 832 26171
rect 864 26139 904 26171
rect 936 26139 976 26171
rect 1008 26139 1048 26171
rect 1080 26139 1120 26171
rect 1152 26139 1192 26171
rect 1224 26139 1264 26171
rect 1296 26139 1336 26171
rect 1368 26139 1408 26171
rect 1440 26139 1480 26171
rect 1512 26139 1552 26171
rect 1584 26139 1624 26171
rect 1656 26139 1696 26171
rect 1728 26139 1768 26171
rect 1800 26139 1840 26171
rect 1872 26139 1912 26171
rect 1944 26139 1984 26171
rect 2016 26139 2056 26171
rect 2088 26139 2128 26171
rect 2160 26139 2200 26171
rect 2232 26139 2272 26171
rect 2304 26139 2344 26171
rect 2376 26139 2416 26171
rect 2448 26139 2488 26171
rect 2520 26139 2560 26171
rect 2592 26139 2632 26171
rect 2664 26139 2704 26171
rect 2736 26139 2776 26171
rect 2808 26139 2848 26171
rect 2880 26139 2920 26171
rect 2952 26139 2992 26171
rect 3024 26139 3064 26171
rect 3096 26139 3136 26171
rect 3168 26139 3208 26171
rect 3240 26139 3280 26171
rect 3312 26139 3352 26171
rect 3384 26139 3424 26171
rect 3456 26139 3496 26171
rect 3528 26139 3568 26171
rect 3600 26139 3640 26171
rect 3672 26139 3712 26171
rect 3744 26139 3784 26171
rect 3816 26139 3856 26171
rect 3888 26139 4000 26171
rect 0 26099 4000 26139
rect 0 26067 112 26099
rect 144 26067 184 26099
rect 216 26067 256 26099
rect 288 26067 328 26099
rect 360 26067 400 26099
rect 432 26067 472 26099
rect 504 26067 544 26099
rect 576 26067 616 26099
rect 648 26067 688 26099
rect 720 26067 760 26099
rect 792 26067 832 26099
rect 864 26067 904 26099
rect 936 26067 976 26099
rect 1008 26067 1048 26099
rect 1080 26067 1120 26099
rect 1152 26067 1192 26099
rect 1224 26067 1264 26099
rect 1296 26067 1336 26099
rect 1368 26067 1408 26099
rect 1440 26067 1480 26099
rect 1512 26067 1552 26099
rect 1584 26067 1624 26099
rect 1656 26067 1696 26099
rect 1728 26067 1768 26099
rect 1800 26067 1840 26099
rect 1872 26067 1912 26099
rect 1944 26067 1984 26099
rect 2016 26067 2056 26099
rect 2088 26067 2128 26099
rect 2160 26067 2200 26099
rect 2232 26067 2272 26099
rect 2304 26067 2344 26099
rect 2376 26067 2416 26099
rect 2448 26067 2488 26099
rect 2520 26067 2560 26099
rect 2592 26067 2632 26099
rect 2664 26067 2704 26099
rect 2736 26067 2776 26099
rect 2808 26067 2848 26099
rect 2880 26067 2920 26099
rect 2952 26067 2992 26099
rect 3024 26067 3064 26099
rect 3096 26067 3136 26099
rect 3168 26067 3208 26099
rect 3240 26067 3280 26099
rect 3312 26067 3352 26099
rect 3384 26067 3424 26099
rect 3456 26067 3496 26099
rect 3528 26067 3568 26099
rect 3600 26067 3640 26099
rect 3672 26067 3712 26099
rect 3744 26067 3784 26099
rect 3816 26067 3856 26099
rect 3888 26067 4000 26099
rect 0 26027 4000 26067
rect 0 25995 112 26027
rect 144 25995 184 26027
rect 216 25995 256 26027
rect 288 25995 328 26027
rect 360 25995 400 26027
rect 432 25995 472 26027
rect 504 25995 544 26027
rect 576 25995 616 26027
rect 648 25995 688 26027
rect 720 25995 760 26027
rect 792 25995 832 26027
rect 864 25995 904 26027
rect 936 25995 976 26027
rect 1008 25995 1048 26027
rect 1080 25995 1120 26027
rect 1152 25995 1192 26027
rect 1224 25995 1264 26027
rect 1296 25995 1336 26027
rect 1368 25995 1408 26027
rect 1440 25995 1480 26027
rect 1512 25995 1552 26027
rect 1584 25995 1624 26027
rect 1656 25995 1696 26027
rect 1728 25995 1768 26027
rect 1800 25995 1840 26027
rect 1872 25995 1912 26027
rect 1944 25995 1984 26027
rect 2016 25995 2056 26027
rect 2088 25995 2128 26027
rect 2160 25995 2200 26027
rect 2232 25995 2272 26027
rect 2304 25995 2344 26027
rect 2376 25995 2416 26027
rect 2448 25995 2488 26027
rect 2520 25995 2560 26027
rect 2592 25995 2632 26027
rect 2664 25995 2704 26027
rect 2736 25995 2776 26027
rect 2808 25995 2848 26027
rect 2880 25995 2920 26027
rect 2952 25995 2992 26027
rect 3024 25995 3064 26027
rect 3096 25995 3136 26027
rect 3168 25995 3208 26027
rect 3240 25995 3280 26027
rect 3312 25995 3352 26027
rect 3384 25995 3424 26027
rect 3456 25995 3496 26027
rect 3528 25995 3568 26027
rect 3600 25995 3640 26027
rect 3672 25995 3712 26027
rect 3744 25995 3784 26027
rect 3816 25995 3856 26027
rect 3888 25995 4000 26027
rect 0 25955 4000 25995
rect 0 25923 112 25955
rect 144 25923 184 25955
rect 216 25923 256 25955
rect 288 25923 328 25955
rect 360 25923 400 25955
rect 432 25923 472 25955
rect 504 25923 544 25955
rect 576 25923 616 25955
rect 648 25923 688 25955
rect 720 25923 760 25955
rect 792 25923 832 25955
rect 864 25923 904 25955
rect 936 25923 976 25955
rect 1008 25923 1048 25955
rect 1080 25923 1120 25955
rect 1152 25923 1192 25955
rect 1224 25923 1264 25955
rect 1296 25923 1336 25955
rect 1368 25923 1408 25955
rect 1440 25923 1480 25955
rect 1512 25923 1552 25955
rect 1584 25923 1624 25955
rect 1656 25923 1696 25955
rect 1728 25923 1768 25955
rect 1800 25923 1840 25955
rect 1872 25923 1912 25955
rect 1944 25923 1984 25955
rect 2016 25923 2056 25955
rect 2088 25923 2128 25955
rect 2160 25923 2200 25955
rect 2232 25923 2272 25955
rect 2304 25923 2344 25955
rect 2376 25923 2416 25955
rect 2448 25923 2488 25955
rect 2520 25923 2560 25955
rect 2592 25923 2632 25955
rect 2664 25923 2704 25955
rect 2736 25923 2776 25955
rect 2808 25923 2848 25955
rect 2880 25923 2920 25955
rect 2952 25923 2992 25955
rect 3024 25923 3064 25955
rect 3096 25923 3136 25955
rect 3168 25923 3208 25955
rect 3240 25923 3280 25955
rect 3312 25923 3352 25955
rect 3384 25923 3424 25955
rect 3456 25923 3496 25955
rect 3528 25923 3568 25955
rect 3600 25923 3640 25955
rect 3672 25923 3712 25955
rect 3744 25923 3784 25955
rect 3816 25923 3856 25955
rect 3888 25923 4000 25955
rect 0 25883 4000 25923
rect 0 25851 112 25883
rect 144 25851 184 25883
rect 216 25851 256 25883
rect 288 25851 328 25883
rect 360 25851 400 25883
rect 432 25851 472 25883
rect 504 25851 544 25883
rect 576 25851 616 25883
rect 648 25851 688 25883
rect 720 25851 760 25883
rect 792 25851 832 25883
rect 864 25851 904 25883
rect 936 25851 976 25883
rect 1008 25851 1048 25883
rect 1080 25851 1120 25883
rect 1152 25851 1192 25883
rect 1224 25851 1264 25883
rect 1296 25851 1336 25883
rect 1368 25851 1408 25883
rect 1440 25851 1480 25883
rect 1512 25851 1552 25883
rect 1584 25851 1624 25883
rect 1656 25851 1696 25883
rect 1728 25851 1768 25883
rect 1800 25851 1840 25883
rect 1872 25851 1912 25883
rect 1944 25851 1984 25883
rect 2016 25851 2056 25883
rect 2088 25851 2128 25883
rect 2160 25851 2200 25883
rect 2232 25851 2272 25883
rect 2304 25851 2344 25883
rect 2376 25851 2416 25883
rect 2448 25851 2488 25883
rect 2520 25851 2560 25883
rect 2592 25851 2632 25883
rect 2664 25851 2704 25883
rect 2736 25851 2776 25883
rect 2808 25851 2848 25883
rect 2880 25851 2920 25883
rect 2952 25851 2992 25883
rect 3024 25851 3064 25883
rect 3096 25851 3136 25883
rect 3168 25851 3208 25883
rect 3240 25851 3280 25883
rect 3312 25851 3352 25883
rect 3384 25851 3424 25883
rect 3456 25851 3496 25883
rect 3528 25851 3568 25883
rect 3600 25851 3640 25883
rect 3672 25851 3712 25883
rect 3744 25851 3784 25883
rect 3816 25851 3856 25883
rect 3888 25851 4000 25883
rect 0 25811 4000 25851
rect 0 25779 112 25811
rect 144 25779 184 25811
rect 216 25779 256 25811
rect 288 25779 328 25811
rect 360 25779 400 25811
rect 432 25779 472 25811
rect 504 25779 544 25811
rect 576 25779 616 25811
rect 648 25779 688 25811
rect 720 25779 760 25811
rect 792 25779 832 25811
rect 864 25779 904 25811
rect 936 25779 976 25811
rect 1008 25779 1048 25811
rect 1080 25779 1120 25811
rect 1152 25779 1192 25811
rect 1224 25779 1264 25811
rect 1296 25779 1336 25811
rect 1368 25779 1408 25811
rect 1440 25779 1480 25811
rect 1512 25779 1552 25811
rect 1584 25779 1624 25811
rect 1656 25779 1696 25811
rect 1728 25779 1768 25811
rect 1800 25779 1840 25811
rect 1872 25779 1912 25811
rect 1944 25779 1984 25811
rect 2016 25779 2056 25811
rect 2088 25779 2128 25811
rect 2160 25779 2200 25811
rect 2232 25779 2272 25811
rect 2304 25779 2344 25811
rect 2376 25779 2416 25811
rect 2448 25779 2488 25811
rect 2520 25779 2560 25811
rect 2592 25779 2632 25811
rect 2664 25779 2704 25811
rect 2736 25779 2776 25811
rect 2808 25779 2848 25811
rect 2880 25779 2920 25811
rect 2952 25779 2992 25811
rect 3024 25779 3064 25811
rect 3096 25779 3136 25811
rect 3168 25779 3208 25811
rect 3240 25779 3280 25811
rect 3312 25779 3352 25811
rect 3384 25779 3424 25811
rect 3456 25779 3496 25811
rect 3528 25779 3568 25811
rect 3600 25779 3640 25811
rect 3672 25779 3712 25811
rect 3744 25779 3784 25811
rect 3816 25779 3856 25811
rect 3888 25779 4000 25811
rect 0 25739 4000 25779
rect 0 25707 112 25739
rect 144 25707 184 25739
rect 216 25707 256 25739
rect 288 25707 328 25739
rect 360 25707 400 25739
rect 432 25707 472 25739
rect 504 25707 544 25739
rect 576 25707 616 25739
rect 648 25707 688 25739
rect 720 25707 760 25739
rect 792 25707 832 25739
rect 864 25707 904 25739
rect 936 25707 976 25739
rect 1008 25707 1048 25739
rect 1080 25707 1120 25739
rect 1152 25707 1192 25739
rect 1224 25707 1264 25739
rect 1296 25707 1336 25739
rect 1368 25707 1408 25739
rect 1440 25707 1480 25739
rect 1512 25707 1552 25739
rect 1584 25707 1624 25739
rect 1656 25707 1696 25739
rect 1728 25707 1768 25739
rect 1800 25707 1840 25739
rect 1872 25707 1912 25739
rect 1944 25707 1984 25739
rect 2016 25707 2056 25739
rect 2088 25707 2128 25739
rect 2160 25707 2200 25739
rect 2232 25707 2272 25739
rect 2304 25707 2344 25739
rect 2376 25707 2416 25739
rect 2448 25707 2488 25739
rect 2520 25707 2560 25739
rect 2592 25707 2632 25739
rect 2664 25707 2704 25739
rect 2736 25707 2776 25739
rect 2808 25707 2848 25739
rect 2880 25707 2920 25739
rect 2952 25707 2992 25739
rect 3024 25707 3064 25739
rect 3096 25707 3136 25739
rect 3168 25707 3208 25739
rect 3240 25707 3280 25739
rect 3312 25707 3352 25739
rect 3384 25707 3424 25739
rect 3456 25707 3496 25739
rect 3528 25707 3568 25739
rect 3600 25707 3640 25739
rect 3672 25707 3712 25739
rect 3744 25707 3784 25739
rect 3816 25707 3856 25739
rect 3888 25707 4000 25739
rect 0 25667 4000 25707
rect 0 25635 112 25667
rect 144 25635 184 25667
rect 216 25635 256 25667
rect 288 25635 328 25667
rect 360 25635 400 25667
rect 432 25635 472 25667
rect 504 25635 544 25667
rect 576 25635 616 25667
rect 648 25635 688 25667
rect 720 25635 760 25667
rect 792 25635 832 25667
rect 864 25635 904 25667
rect 936 25635 976 25667
rect 1008 25635 1048 25667
rect 1080 25635 1120 25667
rect 1152 25635 1192 25667
rect 1224 25635 1264 25667
rect 1296 25635 1336 25667
rect 1368 25635 1408 25667
rect 1440 25635 1480 25667
rect 1512 25635 1552 25667
rect 1584 25635 1624 25667
rect 1656 25635 1696 25667
rect 1728 25635 1768 25667
rect 1800 25635 1840 25667
rect 1872 25635 1912 25667
rect 1944 25635 1984 25667
rect 2016 25635 2056 25667
rect 2088 25635 2128 25667
rect 2160 25635 2200 25667
rect 2232 25635 2272 25667
rect 2304 25635 2344 25667
rect 2376 25635 2416 25667
rect 2448 25635 2488 25667
rect 2520 25635 2560 25667
rect 2592 25635 2632 25667
rect 2664 25635 2704 25667
rect 2736 25635 2776 25667
rect 2808 25635 2848 25667
rect 2880 25635 2920 25667
rect 2952 25635 2992 25667
rect 3024 25635 3064 25667
rect 3096 25635 3136 25667
rect 3168 25635 3208 25667
rect 3240 25635 3280 25667
rect 3312 25635 3352 25667
rect 3384 25635 3424 25667
rect 3456 25635 3496 25667
rect 3528 25635 3568 25667
rect 3600 25635 3640 25667
rect 3672 25635 3712 25667
rect 3744 25635 3784 25667
rect 3816 25635 3856 25667
rect 3888 25635 4000 25667
rect 0 25595 4000 25635
rect 0 25563 112 25595
rect 144 25563 184 25595
rect 216 25563 256 25595
rect 288 25563 328 25595
rect 360 25563 400 25595
rect 432 25563 472 25595
rect 504 25563 544 25595
rect 576 25563 616 25595
rect 648 25563 688 25595
rect 720 25563 760 25595
rect 792 25563 832 25595
rect 864 25563 904 25595
rect 936 25563 976 25595
rect 1008 25563 1048 25595
rect 1080 25563 1120 25595
rect 1152 25563 1192 25595
rect 1224 25563 1264 25595
rect 1296 25563 1336 25595
rect 1368 25563 1408 25595
rect 1440 25563 1480 25595
rect 1512 25563 1552 25595
rect 1584 25563 1624 25595
rect 1656 25563 1696 25595
rect 1728 25563 1768 25595
rect 1800 25563 1840 25595
rect 1872 25563 1912 25595
rect 1944 25563 1984 25595
rect 2016 25563 2056 25595
rect 2088 25563 2128 25595
rect 2160 25563 2200 25595
rect 2232 25563 2272 25595
rect 2304 25563 2344 25595
rect 2376 25563 2416 25595
rect 2448 25563 2488 25595
rect 2520 25563 2560 25595
rect 2592 25563 2632 25595
rect 2664 25563 2704 25595
rect 2736 25563 2776 25595
rect 2808 25563 2848 25595
rect 2880 25563 2920 25595
rect 2952 25563 2992 25595
rect 3024 25563 3064 25595
rect 3096 25563 3136 25595
rect 3168 25563 3208 25595
rect 3240 25563 3280 25595
rect 3312 25563 3352 25595
rect 3384 25563 3424 25595
rect 3456 25563 3496 25595
rect 3528 25563 3568 25595
rect 3600 25563 3640 25595
rect 3672 25563 3712 25595
rect 3744 25563 3784 25595
rect 3816 25563 3856 25595
rect 3888 25563 4000 25595
rect 0 25523 4000 25563
rect 0 25491 112 25523
rect 144 25491 184 25523
rect 216 25491 256 25523
rect 288 25491 328 25523
rect 360 25491 400 25523
rect 432 25491 472 25523
rect 504 25491 544 25523
rect 576 25491 616 25523
rect 648 25491 688 25523
rect 720 25491 760 25523
rect 792 25491 832 25523
rect 864 25491 904 25523
rect 936 25491 976 25523
rect 1008 25491 1048 25523
rect 1080 25491 1120 25523
rect 1152 25491 1192 25523
rect 1224 25491 1264 25523
rect 1296 25491 1336 25523
rect 1368 25491 1408 25523
rect 1440 25491 1480 25523
rect 1512 25491 1552 25523
rect 1584 25491 1624 25523
rect 1656 25491 1696 25523
rect 1728 25491 1768 25523
rect 1800 25491 1840 25523
rect 1872 25491 1912 25523
rect 1944 25491 1984 25523
rect 2016 25491 2056 25523
rect 2088 25491 2128 25523
rect 2160 25491 2200 25523
rect 2232 25491 2272 25523
rect 2304 25491 2344 25523
rect 2376 25491 2416 25523
rect 2448 25491 2488 25523
rect 2520 25491 2560 25523
rect 2592 25491 2632 25523
rect 2664 25491 2704 25523
rect 2736 25491 2776 25523
rect 2808 25491 2848 25523
rect 2880 25491 2920 25523
rect 2952 25491 2992 25523
rect 3024 25491 3064 25523
rect 3096 25491 3136 25523
rect 3168 25491 3208 25523
rect 3240 25491 3280 25523
rect 3312 25491 3352 25523
rect 3384 25491 3424 25523
rect 3456 25491 3496 25523
rect 3528 25491 3568 25523
rect 3600 25491 3640 25523
rect 3672 25491 3712 25523
rect 3744 25491 3784 25523
rect 3816 25491 3856 25523
rect 3888 25491 4000 25523
rect 0 25451 4000 25491
rect 0 25419 112 25451
rect 144 25419 184 25451
rect 216 25419 256 25451
rect 288 25419 328 25451
rect 360 25419 400 25451
rect 432 25419 472 25451
rect 504 25419 544 25451
rect 576 25419 616 25451
rect 648 25419 688 25451
rect 720 25419 760 25451
rect 792 25419 832 25451
rect 864 25419 904 25451
rect 936 25419 976 25451
rect 1008 25419 1048 25451
rect 1080 25419 1120 25451
rect 1152 25419 1192 25451
rect 1224 25419 1264 25451
rect 1296 25419 1336 25451
rect 1368 25419 1408 25451
rect 1440 25419 1480 25451
rect 1512 25419 1552 25451
rect 1584 25419 1624 25451
rect 1656 25419 1696 25451
rect 1728 25419 1768 25451
rect 1800 25419 1840 25451
rect 1872 25419 1912 25451
rect 1944 25419 1984 25451
rect 2016 25419 2056 25451
rect 2088 25419 2128 25451
rect 2160 25419 2200 25451
rect 2232 25419 2272 25451
rect 2304 25419 2344 25451
rect 2376 25419 2416 25451
rect 2448 25419 2488 25451
rect 2520 25419 2560 25451
rect 2592 25419 2632 25451
rect 2664 25419 2704 25451
rect 2736 25419 2776 25451
rect 2808 25419 2848 25451
rect 2880 25419 2920 25451
rect 2952 25419 2992 25451
rect 3024 25419 3064 25451
rect 3096 25419 3136 25451
rect 3168 25419 3208 25451
rect 3240 25419 3280 25451
rect 3312 25419 3352 25451
rect 3384 25419 3424 25451
rect 3456 25419 3496 25451
rect 3528 25419 3568 25451
rect 3600 25419 3640 25451
rect 3672 25419 3712 25451
rect 3744 25419 3784 25451
rect 3816 25419 3856 25451
rect 3888 25419 4000 25451
rect 0 25379 4000 25419
rect 0 25347 112 25379
rect 144 25347 184 25379
rect 216 25347 256 25379
rect 288 25347 328 25379
rect 360 25347 400 25379
rect 432 25347 472 25379
rect 504 25347 544 25379
rect 576 25347 616 25379
rect 648 25347 688 25379
rect 720 25347 760 25379
rect 792 25347 832 25379
rect 864 25347 904 25379
rect 936 25347 976 25379
rect 1008 25347 1048 25379
rect 1080 25347 1120 25379
rect 1152 25347 1192 25379
rect 1224 25347 1264 25379
rect 1296 25347 1336 25379
rect 1368 25347 1408 25379
rect 1440 25347 1480 25379
rect 1512 25347 1552 25379
rect 1584 25347 1624 25379
rect 1656 25347 1696 25379
rect 1728 25347 1768 25379
rect 1800 25347 1840 25379
rect 1872 25347 1912 25379
rect 1944 25347 1984 25379
rect 2016 25347 2056 25379
rect 2088 25347 2128 25379
rect 2160 25347 2200 25379
rect 2232 25347 2272 25379
rect 2304 25347 2344 25379
rect 2376 25347 2416 25379
rect 2448 25347 2488 25379
rect 2520 25347 2560 25379
rect 2592 25347 2632 25379
rect 2664 25347 2704 25379
rect 2736 25347 2776 25379
rect 2808 25347 2848 25379
rect 2880 25347 2920 25379
rect 2952 25347 2992 25379
rect 3024 25347 3064 25379
rect 3096 25347 3136 25379
rect 3168 25347 3208 25379
rect 3240 25347 3280 25379
rect 3312 25347 3352 25379
rect 3384 25347 3424 25379
rect 3456 25347 3496 25379
rect 3528 25347 3568 25379
rect 3600 25347 3640 25379
rect 3672 25347 3712 25379
rect 3744 25347 3784 25379
rect 3816 25347 3856 25379
rect 3888 25347 4000 25379
rect 0 25307 4000 25347
rect 0 25275 112 25307
rect 144 25275 184 25307
rect 216 25275 256 25307
rect 288 25275 328 25307
rect 360 25275 400 25307
rect 432 25275 472 25307
rect 504 25275 544 25307
rect 576 25275 616 25307
rect 648 25275 688 25307
rect 720 25275 760 25307
rect 792 25275 832 25307
rect 864 25275 904 25307
rect 936 25275 976 25307
rect 1008 25275 1048 25307
rect 1080 25275 1120 25307
rect 1152 25275 1192 25307
rect 1224 25275 1264 25307
rect 1296 25275 1336 25307
rect 1368 25275 1408 25307
rect 1440 25275 1480 25307
rect 1512 25275 1552 25307
rect 1584 25275 1624 25307
rect 1656 25275 1696 25307
rect 1728 25275 1768 25307
rect 1800 25275 1840 25307
rect 1872 25275 1912 25307
rect 1944 25275 1984 25307
rect 2016 25275 2056 25307
rect 2088 25275 2128 25307
rect 2160 25275 2200 25307
rect 2232 25275 2272 25307
rect 2304 25275 2344 25307
rect 2376 25275 2416 25307
rect 2448 25275 2488 25307
rect 2520 25275 2560 25307
rect 2592 25275 2632 25307
rect 2664 25275 2704 25307
rect 2736 25275 2776 25307
rect 2808 25275 2848 25307
rect 2880 25275 2920 25307
rect 2952 25275 2992 25307
rect 3024 25275 3064 25307
rect 3096 25275 3136 25307
rect 3168 25275 3208 25307
rect 3240 25275 3280 25307
rect 3312 25275 3352 25307
rect 3384 25275 3424 25307
rect 3456 25275 3496 25307
rect 3528 25275 3568 25307
rect 3600 25275 3640 25307
rect 3672 25275 3712 25307
rect 3744 25275 3784 25307
rect 3816 25275 3856 25307
rect 3888 25275 4000 25307
rect 0 25235 4000 25275
rect 0 25203 112 25235
rect 144 25203 184 25235
rect 216 25203 256 25235
rect 288 25203 328 25235
rect 360 25203 400 25235
rect 432 25203 472 25235
rect 504 25203 544 25235
rect 576 25203 616 25235
rect 648 25203 688 25235
rect 720 25203 760 25235
rect 792 25203 832 25235
rect 864 25203 904 25235
rect 936 25203 976 25235
rect 1008 25203 1048 25235
rect 1080 25203 1120 25235
rect 1152 25203 1192 25235
rect 1224 25203 1264 25235
rect 1296 25203 1336 25235
rect 1368 25203 1408 25235
rect 1440 25203 1480 25235
rect 1512 25203 1552 25235
rect 1584 25203 1624 25235
rect 1656 25203 1696 25235
rect 1728 25203 1768 25235
rect 1800 25203 1840 25235
rect 1872 25203 1912 25235
rect 1944 25203 1984 25235
rect 2016 25203 2056 25235
rect 2088 25203 2128 25235
rect 2160 25203 2200 25235
rect 2232 25203 2272 25235
rect 2304 25203 2344 25235
rect 2376 25203 2416 25235
rect 2448 25203 2488 25235
rect 2520 25203 2560 25235
rect 2592 25203 2632 25235
rect 2664 25203 2704 25235
rect 2736 25203 2776 25235
rect 2808 25203 2848 25235
rect 2880 25203 2920 25235
rect 2952 25203 2992 25235
rect 3024 25203 3064 25235
rect 3096 25203 3136 25235
rect 3168 25203 3208 25235
rect 3240 25203 3280 25235
rect 3312 25203 3352 25235
rect 3384 25203 3424 25235
rect 3456 25203 3496 25235
rect 3528 25203 3568 25235
rect 3600 25203 3640 25235
rect 3672 25203 3712 25235
rect 3744 25203 3784 25235
rect 3816 25203 3856 25235
rect 3888 25203 4000 25235
rect 0 25163 4000 25203
rect 0 25131 112 25163
rect 144 25131 184 25163
rect 216 25131 256 25163
rect 288 25131 328 25163
rect 360 25131 400 25163
rect 432 25131 472 25163
rect 504 25131 544 25163
rect 576 25131 616 25163
rect 648 25131 688 25163
rect 720 25131 760 25163
rect 792 25131 832 25163
rect 864 25131 904 25163
rect 936 25131 976 25163
rect 1008 25131 1048 25163
rect 1080 25131 1120 25163
rect 1152 25131 1192 25163
rect 1224 25131 1264 25163
rect 1296 25131 1336 25163
rect 1368 25131 1408 25163
rect 1440 25131 1480 25163
rect 1512 25131 1552 25163
rect 1584 25131 1624 25163
rect 1656 25131 1696 25163
rect 1728 25131 1768 25163
rect 1800 25131 1840 25163
rect 1872 25131 1912 25163
rect 1944 25131 1984 25163
rect 2016 25131 2056 25163
rect 2088 25131 2128 25163
rect 2160 25131 2200 25163
rect 2232 25131 2272 25163
rect 2304 25131 2344 25163
rect 2376 25131 2416 25163
rect 2448 25131 2488 25163
rect 2520 25131 2560 25163
rect 2592 25131 2632 25163
rect 2664 25131 2704 25163
rect 2736 25131 2776 25163
rect 2808 25131 2848 25163
rect 2880 25131 2920 25163
rect 2952 25131 2992 25163
rect 3024 25131 3064 25163
rect 3096 25131 3136 25163
rect 3168 25131 3208 25163
rect 3240 25131 3280 25163
rect 3312 25131 3352 25163
rect 3384 25131 3424 25163
rect 3456 25131 3496 25163
rect 3528 25131 3568 25163
rect 3600 25131 3640 25163
rect 3672 25131 3712 25163
rect 3744 25131 3784 25163
rect 3816 25131 3856 25163
rect 3888 25131 4000 25163
rect 0 25091 4000 25131
rect 0 25059 112 25091
rect 144 25059 184 25091
rect 216 25059 256 25091
rect 288 25059 328 25091
rect 360 25059 400 25091
rect 432 25059 472 25091
rect 504 25059 544 25091
rect 576 25059 616 25091
rect 648 25059 688 25091
rect 720 25059 760 25091
rect 792 25059 832 25091
rect 864 25059 904 25091
rect 936 25059 976 25091
rect 1008 25059 1048 25091
rect 1080 25059 1120 25091
rect 1152 25059 1192 25091
rect 1224 25059 1264 25091
rect 1296 25059 1336 25091
rect 1368 25059 1408 25091
rect 1440 25059 1480 25091
rect 1512 25059 1552 25091
rect 1584 25059 1624 25091
rect 1656 25059 1696 25091
rect 1728 25059 1768 25091
rect 1800 25059 1840 25091
rect 1872 25059 1912 25091
rect 1944 25059 1984 25091
rect 2016 25059 2056 25091
rect 2088 25059 2128 25091
rect 2160 25059 2200 25091
rect 2232 25059 2272 25091
rect 2304 25059 2344 25091
rect 2376 25059 2416 25091
rect 2448 25059 2488 25091
rect 2520 25059 2560 25091
rect 2592 25059 2632 25091
rect 2664 25059 2704 25091
rect 2736 25059 2776 25091
rect 2808 25059 2848 25091
rect 2880 25059 2920 25091
rect 2952 25059 2992 25091
rect 3024 25059 3064 25091
rect 3096 25059 3136 25091
rect 3168 25059 3208 25091
rect 3240 25059 3280 25091
rect 3312 25059 3352 25091
rect 3384 25059 3424 25091
rect 3456 25059 3496 25091
rect 3528 25059 3568 25091
rect 3600 25059 3640 25091
rect 3672 25059 3712 25091
rect 3744 25059 3784 25091
rect 3816 25059 3856 25091
rect 3888 25059 4000 25091
rect 0 25019 4000 25059
rect 0 24987 112 25019
rect 144 24987 184 25019
rect 216 24987 256 25019
rect 288 24987 328 25019
rect 360 24987 400 25019
rect 432 24987 472 25019
rect 504 24987 544 25019
rect 576 24987 616 25019
rect 648 24987 688 25019
rect 720 24987 760 25019
rect 792 24987 832 25019
rect 864 24987 904 25019
rect 936 24987 976 25019
rect 1008 24987 1048 25019
rect 1080 24987 1120 25019
rect 1152 24987 1192 25019
rect 1224 24987 1264 25019
rect 1296 24987 1336 25019
rect 1368 24987 1408 25019
rect 1440 24987 1480 25019
rect 1512 24987 1552 25019
rect 1584 24987 1624 25019
rect 1656 24987 1696 25019
rect 1728 24987 1768 25019
rect 1800 24987 1840 25019
rect 1872 24987 1912 25019
rect 1944 24987 1984 25019
rect 2016 24987 2056 25019
rect 2088 24987 2128 25019
rect 2160 24987 2200 25019
rect 2232 24987 2272 25019
rect 2304 24987 2344 25019
rect 2376 24987 2416 25019
rect 2448 24987 2488 25019
rect 2520 24987 2560 25019
rect 2592 24987 2632 25019
rect 2664 24987 2704 25019
rect 2736 24987 2776 25019
rect 2808 24987 2848 25019
rect 2880 24987 2920 25019
rect 2952 24987 2992 25019
rect 3024 24987 3064 25019
rect 3096 24987 3136 25019
rect 3168 24987 3208 25019
rect 3240 24987 3280 25019
rect 3312 24987 3352 25019
rect 3384 24987 3424 25019
rect 3456 24987 3496 25019
rect 3528 24987 3568 25019
rect 3600 24987 3640 25019
rect 3672 24987 3712 25019
rect 3744 24987 3784 25019
rect 3816 24987 3856 25019
rect 3888 24987 4000 25019
rect 0 24947 4000 24987
rect 0 24915 112 24947
rect 144 24915 184 24947
rect 216 24915 256 24947
rect 288 24915 328 24947
rect 360 24915 400 24947
rect 432 24915 472 24947
rect 504 24915 544 24947
rect 576 24915 616 24947
rect 648 24915 688 24947
rect 720 24915 760 24947
rect 792 24915 832 24947
rect 864 24915 904 24947
rect 936 24915 976 24947
rect 1008 24915 1048 24947
rect 1080 24915 1120 24947
rect 1152 24915 1192 24947
rect 1224 24915 1264 24947
rect 1296 24915 1336 24947
rect 1368 24915 1408 24947
rect 1440 24915 1480 24947
rect 1512 24915 1552 24947
rect 1584 24915 1624 24947
rect 1656 24915 1696 24947
rect 1728 24915 1768 24947
rect 1800 24915 1840 24947
rect 1872 24915 1912 24947
rect 1944 24915 1984 24947
rect 2016 24915 2056 24947
rect 2088 24915 2128 24947
rect 2160 24915 2200 24947
rect 2232 24915 2272 24947
rect 2304 24915 2344 24947
rect 2376 24915 2416 24947
rect 2448 24915 2488 24947
rect 2520 24915 2560 24947
rect 2592 24915 2632 24947
rect 2664 24915 2704 24947
rect 2736 24915 2776 24947
rect 2808 24915 2848 24947
rect 2880 24915 2920 24947
rect 2952 24915 2992 24947
rect 3024 24915 3064 24947
rect 3096 24915 3136 24947
rect 3168 24915 3208 24947
rect 3240 24915 3280 24947
rect 3312 24915 3352 24947
rect 3384 24915 3424 24947
rect 3456 24915 3496 24947
rect 3528 24915 3568 24947
rect 3600 24915 3640 24947
rect 3672 24915 3712 24947
rect 3744 24915 3784 24947
rect 3816 24915 3856 24947
rect 3888 24915 4000 24947
rect 0 24875 4000 24915
rect 0 24843 112 24875
rect 144 24843 184 24875
rect 216 24843 256 24875
rect 288 24843 328 24875
rect 360 24843 400 24875
rect 432 24843 472 24875
rect 504 24843 544 24875
rect 576 24843 616 24875
rect 648 24843 688 24875
rect 720 24843 760 24875
rect 792 24843 832 24875
rect 864 24843 904 24875
rect 936 24843 976 24875
rect 1008 24843 1048 24875
rect 1080 24843 1120 24875
rect 1152 24843 1192 24875
rect 1224 24843 1264 24875
rect 1296 24843 1336 24875
rect 1368 24843 1408 24875
rect 1440 24843 1480 24875
rect 1512 24843 1552 24875
rect 1584 24843 1624 24875
rect 1656 24843 1696 24875
rect 1728 24843 1768 24875
rect 1800 24843 1840 24875
rect 1872 24843 1912 24875
rect 1944 24843 1984 24875
rect 2016 24843 2056 24875
rect 2088 24843 2128 24875
rect 2160 24843 2200 24875
rect 2232 24843 2272 24875
rect 2304 24843 2344 24875
rect 2376 24843 2416 24875
rect 2448 24843 2488 24875
rect 2520 24843 2560 24875
rect 2592 24843 2632 24875
rect 2664 24843 2704 24875
rect 2736 24843 2776 24875
rect 2808 24843 2848 24875
rect 2880 24843 2920 24875
rect 2952 24843 2992 24875
rect 3024 24843 3064 24875
rect 3096 24843 3136 24875
rect 3168 24843 3208 24875
rect 3240 24843 3280 24875
rect 3312 24843 3352 24875
rect 3384 24843 3424 24875
rect 3456 24843 3496 24875
rect 3528 24843 3568 24875
rect 3600 24843 3640 24875
rect 3672 24843 3712 24875
rect 3744 24843 3784 24875
rect 3816 24843 3856 24875
rect 3888 24843 4000 24875
rect 0 24803 4000 24843
rect 0 24771 112 24803
rect 144 24771 184 24803
rect 216 24771 256 24803
rect 288 24771 328 24803
rect 360 24771 400 24803
rect 432 24771 472 24803
rect 504 24771 544 24803
rect 576 24771 616 24803
rect 648 24771 688 24803
rect 720 24771 760 24803
rect 792 24771 832 24803
rect 864 24771 904 24803
rect 936 24771 976 24803
rect 1008 24771 1048 24803
rect 1080 24771 1120 24803
rect 1152 24771 1192 24803
rect 1224 24771 1264 24803
rect 1296 24771 1336 24803
rect 1368 24771 1408 24803
rect 1440 24771 1480 24803
rect 1512 24771 1552 24803
rect 1584 24771 1624 24803
rect 1656 24771 1696 24803
rect 1728 24771 1768 24803
rect 1800 24771 1840 24803
rect 1872 24771 1912 24803
rect 1944 24771 1984 24803
rect 2016 24771 2056 24803
rect 2088 24771 2128 24803
rect 2160 24771 2200 24803
rect 2232 24771 2272 24803
rect 2304 24771 2344 24803
rect 2376 24771 2416 24803
rect 2448 24771 2488 24803
rect 2520 24771 2560 24803
rect 2592 24771 2632 24803
rect 2664 24771 2704 24803
rect 2736 24771 2776 24803
rect 2808 24771 2848 24803
rect 2880 24771 2920 24803
rect 2952 24771 2992 24803
rect 3024 24771 3064 24803
rect 3096 24771 3136 24803
rect 3168 24771 3208 24803
rect 3240 24771 3280 24803
rect 3312 24771 3352 24803
rect 3384 24771 3424 24803
rect 3456 24771 3496 24803
rect 3528 24771 3568 24803
rect 3600 24771 3640 24803
rect 3672 24771 3712 24803
rect 3744 24771 3784 24803
rect 3816 24771 3856 24803
rect 3888 24771 4000 24803
rect 0 24731 4000 24771
rect 0 24699 112 24731
rect 144 24699 184 24731
rect 216 24699 256 24731
rect 288 24699 328 24731
rect 360 24699 400 24731
rect 432 24699 472 24731
rect 504 24699 544 24731
rect 576 24699 616 24731
rect 648 24699 688 24731
rect 720 24699 760 24731
rect 792 24699 832 24731
rect 864 24699 904 24731
rect 936 24699 976 24731
rect 1008 24699 1048 24731
rect 1080 24699 1120 24731
rect 1152 24699 1192 24731
rect 1224 24699 1264 24731
rect 1296 24699 1336 24731
rect 1368 24699 1408 24731
rect 1440 24699 1480 24731
rect 1512 24699 1552 24731
rect 1584 24699 1624 24731
rect 1656 24699 1696 24731
rect 1728 24699 1768 24731
rect 1800 24699 1840 24731
rect 1872 24699 1912 24731
rect 1944 24699 1984 24731
rect 2016 24699 2056 24731
rect 2088 24699 2128 24731
rect 2160 24699 2200 24731
rect 2232 24699 2272 24731
rect 2304 24699 2344 24731
rect 2376 24699 2416 24731
rect 2448 24699 2488 24731
rect 2520 24699 2560 24731
rect 2592 24699 2632 24731
rect 2664 24699 2704 24731
rect 2736 24699 2776 24731
rect 2808 24699 2848 24731
rect 2880 24699 2920 24731
rect 2952 24699 2992 24731
rect 3024 24699 3064 24731
rect 3096 24699 3136 24731
rect 3168 24699 3208 24731
rect 3240 24699 3280 24731
rect 3312 24699 3352 24731
rect 3384 24699 3424 24731
rect 3456 24699 3496 24731
rect 3528 24699 3568 24731
rect 3600 24699 3640 24731
rect 3672 24699 3712 24731
rect 3744 24699 3784 24731
rect 3816 24699 3856 24731
rect 3888 24699 4000 24731
rect 0 24659 4000 24699
rect 0 24627 112 24659
rect 144 24627 184 24659
rect 216 24627 256 24659
rect 288 24627 328 24659
rect 360 24627 400 24659
rect 432 24627 472 24659
rect 504 24627 544 24659
rect 576 24627 616 24659
rect 648 24627 688 24659
rect 720 24627 760 24659
rect 792 24627 832 24659
rect 864 24627 904 24659
rect 936 24627 976 24659
rect 1008 24627 1048 24659
rect 1080 24627 1120 24659
rect 1152 24627 1192 24659
rect 1224 24627 1264 24659
rect 1296 24627 1336 24659
rect 1368 24627 1408 24659
rect 1440 24627 1480 24659
rect 1512 24627 1552 24659
rect 1584 24627 1624 24659
rect 1656 24627 1696 24659
rect 1728 24627 1768 24659
rect 1800 24627 1840 24659
rect 1872 24627 1912 24659
rect 1944 24627 1984 24659
rect 2016 24627 2056 24659
rect 2088 24627 2128 24659
rect 2160 24627 2200 24659
rect 2232 24627 2272 24659
rect 2304 24627 2344 24659
rect 2376 24627 2416 24659
rect 2448 24627 2488 24659
rect 2520 24627 2560 24659
rect 2592 24627 2632 24659
rect 2664 24627 2704 24659
rect 2736 24627 2776 24659
rect 2808 24627 2848 24659
rect 2880 24627 2920 24659
rect 2952 24627 2992 24659
rect 3024 24627 3064 24659
rect 3096 24627 3136 24659
rect 3168 24627 3208 24659
rect 3240 24627 3280 24659
rect 3312 24627 3352 24659
rect 3384 24627 3424 24659
rect 3456 24627 3496 24659
rect 3528 24627 3568 24659
rect 3600 24627 3640 24659
rect 3672 24627 3712 24659
rect 3744 24627 3784 24659
rect 3816 24627 3856 24659
rect 3888 24627 4000 24659
rect 0 24587 4000 24627
rect 0 24555 112 24587
rect 144 24555 184 24587
rect 216 24555 256 24587
rect 288 24555 328 24587
rect 360 24555 400 24587
rect 432 24555 472 24587
rect 504 24555 544 24587
rect 576 24555 616 24587
rect 648 24555 688 24587
rect 720 24555 760 24587
rect 792 24555 832 24587
rect 864 24555 904 24587
rect 936 24555 976 24587
rect 1008 24555 1048 24587
rect 1080 24555 1120 24587
rect 1152 24555 1192 24587
rect 1224 24555 1264 24587
rect 1296 24555 1336 24587
rect 1368 24555 1408 24587
rect 1440 24555 1480 24587
rect 1512 24555 1552 24587
rect 1584 24555 1624 24587
rect 1656 24555 1696 24587
rect 1728 24555 1768 24587
rect 1800 24555 1840 24587
rect 1872 24555 1912 24587
rect 1944 24555 1984 24587
rect 2016 24555 2056 24587
rect 2088 24555 2128 24587
rect 2160 24555 2200 24587
rect 2232 24555 2272 24587
rect 2304 24555 2344 24587
rect 2376 24555 2416 24587
rect 2448 24555 2488 24587
rect 2520 24555 2560 24587
rect 2592 24555 2632 24587
rect 2664 24555 2704 24587
rect 2736 24555 2776 24587
rect 2808 24555 2848 24587
rect 2880 24555 2920 24587
rect 2952 24555 2992 24587
rect 3024 24555 3064 24587
rect 3096 24555 3136 24587
rect 3168 24555 3208 24587
rect 3240 24555 3280 24587
rect 3312 24555 3352 24587
rect 3384 24555 3424 24587
rect 3456 24555 3496 24587
rect 3528 24555 3568 24587
rect 3600 24555 3640 24587
rect 3672 24555 3712 24587
rect 3744 24555 3784 24587
rect 3816 24555 3856 24587
rect 3888 24555 4000 24587
rect 0 24515 4000 24555
rect 0 24483 112 24515
rect 144 24483 184 24515
rect 216 24483 256 24515
rect 288 24483 328 24515
rect 360 24483 400 24515
rect 432 24483 472 24515
rect 504 24483 544 24515
rect 576 24483 616 24515
rect 648 24483 688 24515
rect 720 24483 760 24515
rect 792 24483 832 24515
rect 864 24483 904 24515
rect 936 24483 976 24515
rect 1008 24483 1048 24515
rect 1080 24483 1120 24515
rect 1152 24483 1192 24515
rect 1224 24483 1264 24515
rect 1296 24483 1336 24515
rect 1368 24483 1408 24515
rect 1440 24483 1480 24515
rect 1512 24483 1552 24515
rect 1584 24483 1624 24515
rect 1656 24483 1696 24515
rect 1728 24483 1768 24515
rect 1800 24483 1840 24515
rect 1872 24483 1912 24515
rect 1944 24483 1984 24515
rect 2016 24483 2056 24515
rect 2088 24483 2128 24515
rect 2160 24483 2200 24515
rect 2232 24483 2272 24515
rect 2304 24483 2344 24515
rect 2376 24483 2416 24515
rect 2448 24483 2488 24515
rect 2520 24483 2560 24515
rect 2592 24483 2632 24515
rect 2664 24483 2704 24515
rect 2736 24483 2776 24515
rect 2808 24483 2848 24515
rect 2880 24483 2920 24515
rect 2952 24483 2992 24515
rect 3024 24483 3064 24515
rect 3096 24483 3136 24515
rect 3168 24483 3208 24515
rect 3240 24483 3280 24515
rect 3312 24483 3352 24515
rect 3384 24483 3424 24515
rect 3456 24483 3496 24515
rect 3528 24483 3568 24515
rect 3600 24483 3640 24515
rect 3672 24483 3712 24515
rect 3744 24483 3784 24515
rect 3816 24483 3856 24515
rect 3888 24483 4000 24515
rect 0 24443 4000 24483
rect 0 24411 112 24443
rect 144 24411 184 24443
rect 216 24411 256 24443
rect 288 24411 328 24443
rect 360 24411 400 24443
rect 432 24411 472 24443
rect 504 24411 544 24443
rect 576 24411 616 24443
rect 648 24411 688 24443
rect 720 24411 760 24443
rect 792 24411 832 24443
rect 864 24411 904 24443
rect 936 24411 976 24443
rect 1008 24411 1048 24443
rect 1080 24411 1120 24443
rect 1152 24411 1192 24443
rect 1224 24411 1264 24443
rect 1296 24411 1336 24443
rect 1368 24411 1408 24443
rect 1440 24411 1480 24443
rect 1512 24411 1552 24443
rect 1584 24411 1624 24443
rect 1656 24411 1696 24443
rect 1728 24411 1768 24443
rect 1800 24411 1840 24443
rect 1872 24411 1912 24443
rect 1944 24411 1984 24443
rect 2016 24411 2056 24443
rect 2088 24411 2128 24443
rect 2160 24411 2200 24443
rect 2232 24411 2272 24443
rect 2304 24411 2344 24443
rect 2376 24411 2416 24443
rect 2448 24411 2488 24443
rect 2520 24411 2560 24443
rect 2592 24411 2632 24443
rect 2664 24411 2704 24443
rect 2736 24411 2776 24443
rect 2808 24411 2848 24443
rect 2880 24411 2920 24443
rect 2952 24411 2992 24443
rect 3024 24411 3064 24443
rect 3096 24411 3136 24443
rect 3168 24411 3208 24443
rect 3240 24411 3280 24443
rect 3312 24411 3352 24443
rect 3384 24411 3424 24443
rect 3456 24411 3496 24443
rect 3528 24411 3568 24443
rect 3600 24411 3640 24443
rect 3672 24411 3712 24443
rect 3744 24411 3784 24443
rect 3816 24411 3856 24443
rect 3888 24411 4000 24443
rect 0 24371 4000 24411
rect 0 24339 112 24371
rect 144 24339 184 24371
rect 216 24339 256 24371
rect 288 24339 328 24371
rect 360 24339 400 24371
rect 432 24339 472 24371
rect 504 24339 544 24371
rect 576 24339 616 24371
rect 648 24339 688 24371
rect 720 24339 760 24371
rect 792 24339 832 24371
rect 864 24339 904 24371
rect 936 24339 976 24371
rect 1008 24339 1048 24371
rect 1080 24339 1120 24371
rect 1152 24339 1192 24371
rect 1224 24339 1264 24371
rect 1296 24339 1336 24371
rect 1368 24339 1408 24371
rect 1440 24339 1480 24371
rect 1512 24339 1552 24371
rect 1584 24339 1624 24371
rect 1656 24339 1696 24371
rect 1728 24339 1768 24371
rect 1800 24339 1840 24371
rect 1872 24339 1912 24371
rect 1944 24339 1984 24371
rect 2016 24339 2056 24371
rect 2088 24339 2128 24371
rect 2160 24339 2200 24371
rect 2232 24339 2272 24371
rect 2304 24339 2344 24371
rect 2376 24339 2416 24371
rect 2448 24339 2488 24371
rect 2520 24339 2560 24371
rect 2592 24339 2632 24371
rect 2664 24339 2704 24371
rect 2736 24339 2776 24371
rect 2808 24339 2848 24371
rect 2880 24339 2920 24371
rect 2952 24339 2992 24371
rect 3024 24339 3064 24371
rect 3096 24339 3136 24371
rect 3168 24339 3208 24371
rect 3240 24339 3280 24371
rect 3312 24339 3352 24371
rect 3384 24339 3424 24371
rect 3456 24339 3496 24371
rect 3528 24339 3568 24371
rect 3600 24339 3640 24371
rect 3672 24339 3712 24371
rect 3744 24339 3784 24371
rect 3816 24339 3856 24371
rect 3888 24339 4000 24371
rect 0 24299 4000 24339
rect 0 24267 112 24299
rect 144 24267 184 24299
rect 216 24267 256 24299
rect 288 24267 328 24299
rect 360 24267 400 24299
rect 432 24267 472 24299
rect 504 24267 544 24299
rect 576 24267 616 24299
rect 648 24267 688 24299
rect 720 24267 760 24299
rect 792 24267 832 24299
rect 864 24267 904 24299
rect 936 24267 976 24299
rect 1008 24267 1048 24299
rect 1080 24267 1120 24299
rect 1152 24267 1192 24299
rect 1224 24267 1264 24299
rect 1296 24267 1336 24299
rect 1368 24267 1408 24299
rect 1440 24267 1480 24299
rect 1512 24267 1552 24299
rect 1584 24267 1624 24299
rect 1656 24267 1696 24299
rect 1728 24267 1768 24299
rect 1800 24267 1840 24299
rect 1872 24267 1912 24299
rect 1944 24267 1984 24299
rect 2016 24267 2056 24299
rect 2088 24267 2128 24299
rect 2160 24267 2200 24299
rect 2232 24267 2272 24299
rect 2304 24267 2344 24299
rect 2376 24267 2416 24299
rect 2448 24267 2488 24299
rect 2520 24267 2560 24299
rect 2592 24267 2632 24299
rect 2664 24267 2704 24299
rect 2736 24267 2776 24299
rect 2808 24267 2848 24299
rect 2880 24267 2920 24299
rect 2952 24267 2992 24299
rect 3024 24267 3064 24299
rect 3096 24267 3136 24299
rect 3168 24267 3208 24299
rect 3240 24267 3280 24299
rect 3312 24267 3352 24299
rect 3384 24267 3424 24299
rect 3456 24267 3496 24299
rect 3528 24267 3568 24299
rect 3600 24267 3640 24299
rect 3672 24267 3712 24299
rect 3744 24267 3784 24299
rect 3816 24267 3856 24299
rect 3888 24267 4000 24299
rect 0 24227 4000 24267
rect 0 24195 112 24227
rect 144 24195 184 24227
rect 216 24195 256 24227
rect 288 24195 328 24227
rect 360 24195 400 24227
rect 432 24195 472 24227
rect 504 24195 544 24227
rect 576 24195 616 24227
rect 648 24195 688 24227
rect 720 24195 760 24227
rect 792 24195 832 24227
rect 864 24195 904 24227
rect 936 24195 976 24227
rect 1008 24195 1048 24227
rect 1080 24195 1120 24227
rect 1152 24195 1192 24227
rect 1224 24195 1264 24227
rect 1296 24195 1336 24227
rect 1368 24195 1408 24227
rect 1440 24195 1480 24227
rect 1512 24195 1552 24227
rect 1584 24195 1624 24227
rect 1656 24195 1696 24227
rect 1728 24195 1768 24227
rect 1800 24195 1840 24227
rect 1872 24195 1912 24227
rect 1944 24195 1984 24227
rect 2016 24195 2056 24227
rect 2088 24195 2128 24227
rect 2160 24195 2200 24227
rect 2232 24195 2272 24227
rect 2304 24195 2344 24227
rect 2376 24195 2416 24227
rect 2448 24195 2488 24227
rect 2520 24195 2560 24227
rect 2592 24195 2632 24227
rect 2664 24195 2704 24227
rect 2736 24195 2776 24227
rect 2808 24195 2848 24227
rect 2880 24195 2920 24227
rect 2952 24195 2992 24227
rect 3024 24195 3064 24227
rect 3096 24195 3136 24227
rect 3168 24195 3208 24227
rect 3240 24195 3280 24227
rect 3312 24195 3352 24227
rect 3384 24195 3424 24227
rect 3456 24195 3496 24227
rect 3528 24195 3568 24227
rect 3600 24195 3640 24227
rect 3672 24195 3712 24227
rect 3744 24195 3784 24227
rect 3816 24195 3856 24227
rect 3888 24195 4000 24227
rect 0 24155 4000 24195
rect 0 24123 112 24155
rect 144 24123 184 24155
rect 216 24123 256 24155
rect 288 24123 328 24155
rect 360 24123 400 24155
rect 432 24123 472 24155
rect 504 24123 544 24155
rect 576 24123 616 24155
rect 648 24123 688 24155
rect 720 24123 760 24155
rect 792 24123 832 24155
rect 864 24123 904 24155
rect 936 24123 976 24155
rect 1008 24123 1048 24155
rect 1080 24123 1120 24155
rect 1152 24123 1192 24155
rect 1224 24123 1264 24155
rect 1296 24123 1336 24155
rect 1368 24123 1408 24155
rect 1440 24123 1480 24155
rect 1512 24123 1552 24155
rect 1584 24123 1624 24155
rect 1656 24123 1696 24155
rect 1728 24123 1768 24155
rect 1800 24123 1840 24155
rect 1872 24123 1912 24155
rect 1944 24123 1984 24155
rect 2016 24123 2056 24155
rect 2088 24123 2128 24155
rect 2160 24123 2200 24155
rect 2232 24123 2272 24155
rect 2304 24123 2344 24155
rect 2376 24123 2416 24155
rect 2448 24123 2488 24155
rect 2520 24123 2560 24155
rect 2592 24123 2632 24155
rect 2664 24123 2704 24155
rect 2736 24123 2776 24155
rect 2808 24123 2848 24155
rect 2880 24123 2920 24155
rect 2952 24123 2992 24155
rect 3024 24123 3064 24155
rect 3096 24123 3136 24155
rect 3168 24123 3208 24155
rect 3240 24123 3280 24155
rect 3312 24123 3352 24155
rect 3384 24123 3424 24155
rect 3456 24123 3496 24155
rect 3528 24123 3568 24155
rect 3600 24123 3640 24155
rect 3672 24123 3712 24155
rect 3744 24123 3784 24155
rect 3816 24123 3856 24155
rect 3888 24123 4000 24155
rect 0 24083 4000 24123
rect 0 24051 112 24083
rect 144 24051 184 24083
rect 216 24051 256 24083
rect 288 24051 328 24083
rect 360 24051 400 24083
rect 432 24051 472 24083
rect 504 24051 544 24083
rect 576 24051 616 24083
rect 648 24051 688 24083
rect 720 24051 760 24083
rect 792 24051 832 24083
rect 864 24051 904 24083
rect 936 24051 976 24083
rect 1008 24051 1048 24083
rect 1080 24051 1120 24083
rect 1152 24051 1192 24083
rect 1224 24051 1264 24083
rect 1296 24051 1336 24083
rect 1368 24051 1408 24083
rect 1440 24051 1480 24083
rect 1512 24051 1552 24083
rect 1584 24051 1624 24083
rect 1656 24051 1696 24083
rect 1728 24051 1768 24083
rect 1800 24051 1840 24083
rect 1872 24051 1912 24083
rect 1944 24051 1984 24083
rect 2016 24051 2056 24083
rect 2088 24051 2128 24083
rect 2160 24051 2200 24083
rect 2232 24051 2272 24083
rect 2304 24051 2344 24083
rect 2376 24051 2416 24083
rect 2448 24051 2488 24083
rect 2520 24051 2560 24083
rect 2592 24051 2632 24083
rect 2664 24051 2704 24083
rect 2736 24051 2776 24083
rect 2808 24051 2848 24083
rect 2880 24051 2920 24083
rect 2952 24051 2992 24083
rect 3024 24051 3064 24083
rect 3096 24051 3136 24083
rect 3168 24051 3208 24083
rect 3240 24051 3280 24083
rect 3312 24051 3352 24083
rect 3384 24051 3424 24083
rect 3456 24051 3496 24083
rect 3528 24051 3568 24083
rect 3600 24051 3640 24083
rect 3672 24051 3712 24083
rect 3744 24051 3784 24083
rect 3816 24051 3856 24083
rect 3888 24051 4000 24083
rect 0 24011 4000 24051
rect 0 23979 112 24011
rect 144 23979 184 24011
rect 216 23979 256 24011
rect 288 23979 328 24011
rect 360 23979 400 24011
rect 432 23979 472 24011
rect 504 23979 544 24011
rect 576 23979 616 24011
rect 648 23979 688 24011
rect 720 23979 760 24011
rect 792 23979 832 24011
rect 864 23979 904 24011
rect 936 23979 976 24011
rect 1008 23979 1048 24011
rect 1080 23979 1120 24011
rect 1152 23979 1192 24011
rect 1224 23979 1264 24011
rect 1296 23979 1336 24011
rect 1368 23979 1408 24011
rect 1440 23979 1480 24011
rect 1512 23979 1552 24011
rect 1584 23979 1624 24011
rect 1656 23979 1696 24011
rect 1728 23979 1768 24011
rect 1800 23979 1840 24011
rect 1872 23979 1912 24011
rect 1944 23979 1984 24011
rect 2016 23979 2056 24011
rect 2088 23979 2128 24011
rect 2160 23979 2200 24011
rect 2232 23979 2272 24011
rect 2304 23979 2344 24011
rect 2376 23979 2416 24011
rect 2448 23979 2488 24011
rect 2520 23979 2560 24011
rect 2592 23979 2632 24011
rect 2664 23979 2704 24011
rect 2736 23979 2776 24011
rect 2808 23979 2848 24011
rect 2880 23979 2920 24011
rect 2952 23979 2992 24011
rect 3024 23979 3064 24011
rect 3096 23979 3136 24011
rect 3168 23979 3208 24011
rect 3240 23979 3280 24011
rect 3312 23979 3352 24011
rect 3384 23979 3424 24011
rect 3456 23979 3496 24011
rect 3528 23979 3568 24011
rect 3600 23979 3640 24011
rect 3672 23979 3712 24011
rect 3744 23979 3784 24011
rect 3816 23979 3856 24011
rect 3888 23979 4000 24011
rect 0 23939 4000 23979
rect 0 23907 112 23939
rect 144 23907 184 23939
rect 216 23907 256 23939
rect 288 23907 328 23939
rect 360 23907 400 23939
rect 432 23907 472 23939
rect 504 23907 544 23939
rect 576 23907 616 23939
rect 648 23907 688 23939
rect 720 23907 760 23939
rect 792 23907 832 23939
rect 864 23907 904 23939
rect 936 23907 976 23939
rect 1008 23907 1048 23939
rect 1080 23907 1120 23939
rect 1152 23907 1192 23939
rect 1224 23907 1264 23939
rect 1296 23907 1336 23939
rect 1368 23907 1408 23939
rect 1440 23907 1480 23939
rect 1512 23907 1552 23939
rect 1584 23907 1624 23939
rect 1656 23907 1696 23939
rect 1728 23907 1768 23939
rect 1800 23907 1840 23939
rect 1872 23907 1912 23939
rect 1944 23907 1984 23939
rect 2016 23907 2056 23939
rect 2088 23907 2128 23939
rect 2160 23907 2200 23939
rect 2232 23907 2272 23939
rect 2304 23907 2344 23939
rect 2376 23907 2416 23939
rect 2448 23907 2488 23939
rect 2520 23907 2560 23939
rect 2592 23907 2632 23939
rect 2664 23907 2704 23939
rect 2736 23907 2776 23939
rect 2808 23907 2848 23939
rect 2880 23907 2920 23939
rect 2952 23907 2992 23939
rect 3024 23907 3064 23939
rect 3096 23907 3136 23939
rect 3168 23907 3208 23939
rect 3240 23907 3280 23939
rect 3312 23907 3352 23939
rect 3384 23907 3424 23939
rect 3456 23907 3496 23939
rect 3528 23907 3568 23939
rect 3600 23907 3640 23939
rect 3672 23907 3712 23939
rect 3744 23907 3784 23939
rect 3816 23907 3856 23939
rect 3888 23907 4000 23939
rect 0 23867 4000 23907
rect 0 23835 112 23867
rect 144 23835 184 23867
rect 216 23835 256 23867
rect 288 23835 328 23867
rect 360 23835 400 23867
rect 432 23835 472 23867
rect 504 23835 544 23867
rect 576 23835 616 23867
rect 648 23835 688 23867
rect 720 23835 760 23867
rect 792 23835 832 23867
rect 864 23835 904 23867
rect 936 23835 976 23867
rect 1008 23835 1048 23867
rect 1080 23835 1120 23867
rect 1152 23835 1192 23867
rect 1224 23835 1264 23867
rect 1296 23835 1336 23867
rect 1368 23835 1408 23867
rect 1440 23835 1480 23867
rect 1512 23835 1552 23867
rect 1584 23835 1624 23867
rect 1656 23835 1696 23867
rect 1728 23835 1768 23867
rect 1800 23835 1840 23867
rect 1872 23835 1912 23867
rect 1944 23835 1984 23867
rect 2016 23835 2056 23867
rect 2088 23835 2128 23867
rect 2160 23835 2200 23867
rect 2232 23835 2272 23867
rect 2304 23835 2344 23867
rect 2376 23835 2416 23867
rect 2448 23835 2488 23867
rect 2520 23835 2560 23867
rect 2592 23835 2632 23867
rect 2664 23835 2704 23867
rect 2736 23835 2776 23867
rect 2808 23835 2848 23867
rect 2880 23835 2920 23867
rect 2952 23835 2992 23867
rect 3024 23835 3064 23867
rect 3096 23835 3136 23867
rect 3168 23835 3208 23867
rect 3240 23835 3280 23867
rect 3312 23835 3352 23867
rect 3384 23835 3424 23867
rect 3456 23835 3496 23867
rect 3528 23835 3568 23867
rect 3600 23835 3640 23867
rect 3672 23835 3712 23867
rect 3744 23835 3784 23867
rect 3816 23835 3856 23867
rect 3888 23835 4000 23867
rect 0 23795 4000 23835
rect 0 23763 112 23795
rect 144 23763 184 23795
rect 216 23763 256 23795
rect 288 23763 328 23795
rect 360 23763 400 23795
rect 432 23763 472 23795
rect 504 23763 544 23795
rect 576 23763 616 23795
rect 648 23763 688 23795
rect 720 23763 760 23795
rect 792 23763 832 23795
rect 864 23763 904 23795
rect 936 23763 976 23795
rect 1008 23763 1048 23795
rect 1080 23763 1120 23795
rect 1152 23763 1192 23795
rect 1224 23763 1264 23795
rect 1296 23763 1336 23795
rect 1368 23763 1408 23795
rect 1440 23763 1480 23795
rect 1512 23763 1552 23795
rect 1584 23763 1624 23795
rect 1656 23763 1696 23795
rect 1728 23763 1768 23795
rect 1800 23763 1840 23795
rect 1872 23763 1912 23795
rect 1944 23763 1984 23795
rect 2016 23763 2056 23795
rect 2088 23763 2128 23795
rect 2160 23763 2200 23795
rect 2232 23763 2272 23795
rect 2304 23763 2344 23795
rect 2376 23763 2416 23795
rect 2448 23763 2488 23795
rect 2520 23763 2560 23795
rect 2592 23763 2632 23795
rect 2664 23763 2704 23795
rect 2736 23763 2776 23795
rect 2808 23763 2848 23795
rect 2880 23763 2920 23795
rect 2952 23763 2992 23795
rect 3024 23763 3064 23795
rect 3096 23763 3136 23795
rect 3168 23763 3208 23795
rect 3240 23763 3280 23795
rect 3312 23763 3352 23795
rect 3384 23763 3424 23795
rect 3456 23763 3496 23795
rect 3528 23763 3568 23795
rect 3600 23763 3640 23795
rect 3672 23763 3712 23795
rect 3744 23763 3784 23795
rect 3816 23763 3856 23795
rect 3888 23763 4000 23795
rect 0 23723 4000 23763
rect 0 23691 112 23723
rect 144 23691 184 23723
rect 216 23691 256 23723
rect 288 23691 328 23723
rect 360 23691 400 23723
rect 432 23691 472 23723
rect 504 23691 544 23723
rect 576 23691 616 23723
rect 648 23691 688 23723
rect 720 23691 760 23723
rect 792 23691 832 23723
rect 864 23691 904 23723
rect 936 23691 976 23723
rect 1008 23691 1048 23723
rect 1080 23691 1120 23723
rect 1152 23691 1192 23723
rect 1224 23691 1264 23723
rect 1296 23691 1336 23723
rect 1368 23691 1408 23723
rect 1440 23691 1480 23723
rect 1512 23691 1552 23723
rect 1584 23691 1624 23723
rect 1656 23691 1696 23723
rect 1728 23691 1768 23723
rect 1800 23691 1840 23723
rect 1872 23691 1912 23723
rect 1944 23691 1984 23723
rect 2016 23691 2056 23723
rect 2088 23691 2128 23723
rect 2160 23691 2200 23723
rect 2232 23691 2272 23723
rect 2304 23691 2344 23723
rect 2376 23691 2416 23723
rect 2448 23691 2488 23723
rect 2520 23691 2560 23723
rect 2592 23691 2632 23723
rect 2664 23691 2704 23723
rect 2736 23691 2776 23723
rect 2808 23691 2848 23723
rect 2880 23691 2920 23723
rect 2952 23691 2992 23723
rect 3024 23691 3064 23723
rect 3096 23691 3136 23723
rect 3168 23691 3208 23723
rect 3240 23691 3280 23723
rect 3312 23691 3352 23723
rect 3384 23691 3424 23723
rect 3456 23691 3496 23723
rect 3528 23691 3568 23723
rect 3600 23691 3640 23723
rect 3672 23691 3712 23723
rect 3744 23691 3784 23723
rect 3816 23691 3856 23723
rect 3888 23691 4000 23723
rect 0 23651 4000 23691
rect 0 23619 112 23651
rect 144 23619 184 23651
rect 216 23619 256 23651
rect 288 23619 328 23651
rect 360 23619 400 23651
rect 432 23619 472 23651
rect 504 23619 544 23651
rect 576 23619 616 23651
rect 648 23619 688 23651
rect 720 23619 760 23651
rect 792 23619 832 23651
rect 864 23619 904 23651
rect 936 23619 976 23651
rect 1008 23619 1048 23651
rect 1080 23619 1120 23651
rect 1152 23619 1192 23651
rect 1224 23619 1264 23651
rect 1296 23619 1336 23651
rect 1368 23619 1408 23651
rect 1440 23619 1480 23651
rect 1512 23619 1552 23651
rect 1584 23619 1624 23651
rect 1656 23619 1696 23651
rect 1728 23619 1768 23651
rect 1800 23619 1840 23651
rect 1872 23619 1912 23651
rect 1944 23619 1984 23651
rect 2016 23619 2056 23651
rect 2088 23619 2128 23651
rect 2160 23619 2200 23651
rect 2232 23619 2272 23651
rect 2304 23619 2344 23651
rect 2376 23619 2416 23651
rect 2448 23619 2488 23651
rect 2520 23619 2560 23651
rect 2592 23619 2632 23651
rect 2664 23619 2704 23651
rect 2736 23619 2776 23651
rect 2808 23619 2848 23651
rect 2880 23619 2920 23651
rect 2952 23619 2992 23651
rect 3024 23619 3064 23651
rect 3096 23619 3136 23651
rect 3168 23619 3208 23651
rect 3240 23619 3280 23651
rect 3312 23619 3352 23651
rect 3384 23619 3424 23651
rect 3456 23619 3496 23651
rect 3528 23619 3568 23651
rect 3600 23619 3640 23651
rect 3672 23619 3712 23651
rect 3744 23619 3784 23651
rect 3816 23619 3856 23651
rect 3888 23619 4000 23651
rect 0 23579 4000 23619
rect 0 23547 112 23579
rect 144 23547 184 23579
rect 216 23547 256 23579
rect 288 23547 328 23579
rect 360 23547 400 23579
rect 432 23547 472 23579
rect 504 23547 544 23579
rect 576 23547 616 23579
rect 648 23547 688 23579
rect 720 23547 760 23579
rect 792 23547 832 23579
rect 864 23547 904 23579
rect 936 23547 976 23579
rect 1008 23547 1048 23579
rect 1080 23547 1120 23579
rect 1152 23547 1192 23579
rect 1224 23547 1264 23579
rect 1296 23547 1336 23579
rect 1368 23547 1408 23579
rect 1440 23547 1480 23579
rect 1512 23547 1552 23579
rect 1584 23547 1624 23579
rect 1656 23547 1696 23579
rect 1728 23547 1768 23579
rect 1800 23547 1840 23579
rect 1872 23547 1912 23579
rect 1944 23547 1984 23579
rect 2016 23547 2056 23579
rect 2088 23547 2128 23579
rect 2160 23547 2200 23579
rect 2232 23547 2272 23579
rect 2304 23547 2344 23579
rect 2376 23547 2416 23579
rect 2448 23547 2488 23579
rect 2520 23547 2560 23579
rect 2592 23547 2632 23579
rect 2664 23547 2704 23579
rect 2736 23547 2776 23579
rect 2808 23547 2848 23579
rect 2880 23547 2920 23579
rect 2952 23547 2992 23579
rect 3024 23547 3064 23579
rect 3096 23547 3136 23579
rect 3168 23547 3208 23579
rect 3240 23547 3280 23579
rect 3312 23547 3352 23579
rect 3384 23547 3424 23579
rect 3456 23547 3496 23579
rect 3528 23547 3568 23579
rect 3600 23547 3640 23579
rect 3672 23547 3712 23579
rect 3744 23547 3784 23579
rect 3816 23547 3856 23579
rect 3888 23547 4000 23579
rect 0 23507 4000 23547
rect 0 23475 112 23507
rect 144 23475 184 23507
rect 216 23475 256 23507
rect 288 23475 328 23507
rect 360 23475 400 23507
rect 432 23475 472 23507
rect 504 23475 544 23507
rect 576 23475 616 23507
rect 648 23475 688 23507
rect 720 23475 760 23507
rect 792 23475 832 23507
rect 864 23475 904 23507
rect 936 23475 976 23507
rect 1008 23475 1048 23507
rect 1080 23475 1120 23507
rect 1152 23475 1192 23507
rect 1224 23475 1264 23507
rect 1296 23475 1336 23507
rect 1368 23475 1408 23507
rect 1440 23475 1480 23507
rect 1512 23475 1552 23507
rect 1584 23475 1624 23507
rect 1656 23475 1696 23507
rect 1728 23475 1768 23507
rect 1800 23475 1840 23507
rect 1872 23475 1912 23507
rect 1944 23475 1984 23507
rect 2016 23475 2056 23507
rect 2088 23475 2128 23507
rect 2160 23475 2200 23507
rect 2232 23475 2272 23507
rect 2304 23475 2344 23507
rect 2376 23475 2416 23507
rect 2448 23475 2488 23507
rect 2520 23475 2560 23507
rect 2592 23475 2632 23507
rect 2664 23475 2704 23507
rect 2736 23475 2776 23507
rect 2808 23475 2848 23507
rect 2880 23475 2920 23507
rect 2952 23475 2992 23507
rect 3024 23475 3064 23507
rect 3096 23475 3136 23507
rect 3168 23475 3208 23507
rect 3240 23475 3280 23507
rect 3312 23475 3352 23507
rect 3384 23475 3424 23507
rect 3456 23475 3496 23507
rect 3528 23475 3568 23507
rect 3600 23475 3640 23507
rect 3672 23475 3712 23507
rect 3744 23475 3784 23507
rect 3816 23475 3856 23507
rect 3888 23475 4000 23507
rect 0 23435 4000 23475
rect 0 23403 112 23435
rect 144 23403 184 23435
rect 216 23403 256 23435
rect 288 23403 328 23435
rect 360 23403 400 23435
rect 432 23403 472 23435
rect 504 23403 544 23435
rect 576 23403 616 23435
rect 648 23403 688 23435
rect 720 23403 760 23435
rect 792 23403 832 23435
rect 864 23403 904 23435
rect 936 23403 976 23435
rect 1008 23403 1048 23435
rect 1080 23403 1120 23435
rect 1152 23403 1192 23435
rect 1224 23403 1264 23435
rect 1296 23403 1336 23435
rect 1368 23403 1408 23435
rect 1440 23403 1480 23435
rect 1512 23403 1552 23435
rect 1584 23403 1624 23435
rect 1656 23403 1696 23435
rect 1728 23403 1768 23435
rect 1800 23403 1840 23435
rect 1872 23403 1912 23435
rect 1944 23403 1984 23435
rect 2016 23403 2056 23435
rect 2088 23403 2128 23435
rect 2160 23403 2200 23435
rect 2232 23403 2272 23435
rect 2304 23403 2344 23435
rect 2376 23403 2416 23435
rect 2448 23403 2488 23435
rect 2520 23403 2560 23435
rect 2592 23403 2632 23435
rect 2664 23403 2704 23435
rect 2736 23403 2776 23435
rect 2808 23403 2848 23435
rect 2880 23403 2920 23435
rect 2952 23403 2992 23435
rect 3024 23403 3064 23435
rect 3096 23403 3136 23435
rect 3168 23403 3208 23435
rect 3240 23403 3280 23435
rect 3312 23403 3352 23435
rect 3384 23403 3424 23435
rect 3456 23403 3496 23435
rect 3528 23403 3568 23435
rect 3600 23403 3640 23435
rect 3672 23403 3712 23435
rect 3744 23403 3784 23435
rect 3816 23403 3856 23435
rect 3888 23403 4000 23435
rect 0 23363 4000 23403
rect 0 23331 112 23363
rect 144 23331 184 23363
rect 216 23331 256 23363
rect 288 23331 328 23363
rect 360 23331 400 23363
rect 432 23331 472 23363
rect 504 23331 544 23363
rect 576 23331 616 23363
rect 648 23331 688 23363
rect 720 23331 760 23363
rect 792 23331 832 23363
rect 864 23331 904 23363
rect 936 23331 976 23363
rect 1008 23331 1048 23363
rect 1080 23331 1120 23363
rect 1152 23331 1192 23363
rect 1224 23331 1264 23363
rect 1296 23331 1336 23363
rect 1368 23331 1408 23363
rect 1440 23331 1480 23363
rect 1512 23331 1552 23363
rect 1584 23331 1624 23363
rect 1656 23331 1696 23363
rect 1728 23331 1768 23363
rect 1800 23331 1840 23363
rect 1872 23331 1912 23363
rect 1944 23331 1984 23363
rect 2016 23331 2056 23363
rect 2088 23331 2128 23363
rect 2160 23331 2200 23363
rect 2232 23331 2272 23363
rect 2304 23331 2344 23363
rect 2376 23331 2416 23363
rect 2448 23331 2488 23363
rect 2520 23331 2560 23363
rect 2592 23331 2632 23363
rect 2664 23331 2704 23363
rect 2736 23331 2776 23363
rect 2808 23331 2848 23363
rect 2880 23331 2920 23363
rect 2952 23331 2992 23363
rect 3024 23331 3064 23363
rect 3096 23331 3136 23363
rect 3168 23331 3208 23363
rect 3240 23331 3280 23363
rect 3312 23331 3352 23363
rect 3384 23331 3424 23363
rect 3456 23331 3496 23363
rect 3528 23331 3568 23363
rect 3600 23331 3640 23363
rect 3672 23331 3712 23363
rect 3744 23331 3784 23363
rect 3816 23331 3856 23363
rect 3888 23331 4000 23363
rect 0 23291 4000 23331
rect 0 23259 112 23291
rect 144 23259 184 23291
rect 216 23259 256 23291
rect 288 23259 328 23291
rect 360 23259 400 23291
rect 432 23259 472 23291
rect 504 23259 544 23291
rect 576 23259 616 23291
rect 648 23259 688 23291
rect 720 23259 760 23291
rect 792 23259 832 23291
rect 864 23259 904 23291
rect 936 23259 976 23291
rect 1008 23259 1048 23291
rect 1080 23259 1120 23291
rect 1152 23259 1192 23291
rect 1224 23259 1264 23291
rect 1296 23259 1336 23291
rect 1368 23259 1408 23291
rect 1440 23259 1480 23291
rect 1512 23259 1552 23291
rect 1584 23259 1624 23291
rect 1656 23259 1696 23291
rect 1728 23259 1768 23291
rect 1800 23259 1840 23291
rect 1872 23259 1912 23291
rect 1944 23259 1984 23291
rect 2016 23259 2056 23291
rect 2088 23259 2128 23291
rect 2160 23259 2200 23291
rect 2232 23259 2272 23291
rect 2304 23259 2344 23291
rect 2376 23259 2416 23291
rect 2448 23259 2488 23291
rect 2520 23259 2560 23291
rect 2592 23259 2632 23291
rect 2664 23259 2704 23291
rect 2736 23259 2776 23291
rect 2808 23259 2848 23291
rect 2880 23259 2920 23291
rect 2952 23259 2992 23291
rect 3024 23259 3064 23291
rect 3096 23259 3136 23291
rect 3168 23259 3208 23291
rect 3240 23259 3280 23291
rect 3312 23259 3352 23291
rect 3384 23259 3424 23291
rect 3456 23259 3496 23291
rect 3528 23259 3568 23291
rect 3600 23259 3640 23291
rect 3672 23259 3712 23291
rect 3744 23259 3784 23291
rect 3816 23259 3856 23291
rect 3888 23259 4000 23291
rect 0 23219 4000 23259
rect 0 23187 112 23219
rect 144 23187 184 23219
rect 216 23187 256 23219
rect 288 23187 328 23219
rect 360 23187 400 23219
rect 432 23187 472 23219
rect 504 23187 544 23219
rect 576 23187 616 23219
rect 648 23187 688 23219
rect 720 23187 760 23219
rect 792 23187 832 23219
rect 864 23187 904 23219
rect 936 23187 976 23219
rect 1008 23187 1048 23219
rect 1080 23187 1120 23219
rect 1152 23187 1192 23219
rect 1224 23187 1264 23219
rect 1296 23187 1336 23219
rect 1368 23187 1408 23219
rect 1440 23187 1480 23219
rect 1512 23187 1552 23219
rect 1584 23187 1624 23219
rect 1656 23187 1696 23219
rect 1728 23187 1768 23219
rect 1800 23187 1840 23219
rect 1872 23187 1912 23219
rect 1944 23187 1984 23219
rect 2016 23187 2056 23219
rect 2088 23187 2128 23219
rect 2160 23187 2200 23219
rect 2232 23187 2272 23219
rect 2304 23187 2344 23219
rect 2376 23187 2416 23219
rect 2448 23187 2488 23219
rect 2520 23187 2560 23219
rect 2592 23187 2632 23219
rect 2664 23187 2704 23219
rect 2736 23187 2776 23219
rect 2808 23187 2848 23219
rect 2880 23187 2920 23219
rect 2952 23187 2992 23219
rect 3024 23187 3064 23219
rect 3096 23187 3136 23219
rect 3168 23187 3208 23219
rect 3240 23187 3280 23219
rect 3312 23187 3352 23219
rect 3384 23187 3424 23219
rect 3456 23187 3496 23219
rect 3528 23187 3568 23219
rect 3600 23187 3640 23219
rect 3672 23187 3712 23219
rect 3744 23187 3784 23219
rect 3816 23187 3856 23219
rect 3888 23187 4000 23219
rect 0 23124 4000 23187
rect 0 22874 4000 22924
rect 0 22842 112 22874
rect 144 22842 184 22874
rect 216 22842 256 22874
rect 288 22842 328 22874
rect 360 22842 400 22874
rect 432 22842 472 22874
rect 504 22842 544 22874
rect 576 22842 616 22874
rect 648 22842 688 22874
rect 720 22842 760 22874
rect 792 22842 832 22874
rect 864 22842 904 22874
rect 936 22842 976 22874
rect 1008 22842 1048 22874
rect 1080 22842 1120 22874
rect 1152 22842 1192 22874
rect 1224 22842 1264 22874
rect 1296 22842 1336 22874
rect 1368 22842 1408 22874
rect 1440 22842 1480 22874
rect 1512 22842 1552 22874
rect 1584 22842 1624 22874
rect 1656 22842 1696 22874
rect 1728 22842 1768 22874
rect 1800 22842 1840 22874
rect 1872 22842 1912 22874
rect 1944 22842 1984 22874
rect 2016 22842 2056 22874
rect 2088 22842 2128 22874
rect 2160 22842 2200 22874
rect 2232 22842 2272 22874
rect 2304 22842 2344 22874
rect 2376 22842 2416 22874
rect 2448 22842 2488 22874
rect 2520 22842 2560 22874
rect 2592 22842 2632 22874
rect 2664 22842 2704 22874
rect 2736 22842 2776 22874
rect 2808 22842 2848 22874
rect 2880 22842 2920 22874
rect 2952 22842 2992 22874
rect 3024 22842 3064 22874
rect 3096 22842 3136 22874
rect 3168 22842 3208 22874
rect 3240 22842 3280 22874
rect 3312 22842 3352 22874
rect 3384 22842 3424 22874
rect 3456 22842 3496 22874
rect 3528 22842 3568 22874
rect 3600 22842 3640 22874
rect 3672 22842 3712 22874
rect 3744 22842 3784 22874
rect 3816 22842 3856 22874
rect 3888 22842 4000 22874
rect 0 22802 4000 22842
rect 0 22770 112 22802
rect 144 22770 184 22802
rect 216 22770 256 22802
rect 288 22770 328 22802
rect 360 22770 400 22802
rect 432 22770 472 22802
rect 504 22770 544 22802
rect 576 22770 616 22802
rect 648 22770 688 22802
rect 720 22770 760 22802
rect 792 22770 832 22802
rect 864 22770 904 22802
rect 936 22770 976 22802
rect 1008 22770 1048 22802
rect 1080 22770 1120 22802
rect 1152 22770 1192 22802
rect 1224 22770 1264 22802
rect 1296 22770 1336 22802
rect 1368 22770 1408 22802
rect 1440 22770 1480 22802
rect 1512 22770 1552 22802
rect 1584 22770 1624 22802
rect 1656 22770 1696 22802
rect 1728 22770 1768 22802
rect 1800 22770 1840 22802
rect 1872 22770 1912 22802
rect 1944 22770 1984 22802
rect 2016 22770 2056 22802
rect 2088 22770 2128 22802
rect 2160 22770 2200 22802
rect 2232 22770 2272 22802
rect 2304 22770 2344 22802
rect 2376 22770 2416 22802
rect 2448 22770 2488 22802
rect 2520 22770 2560 22802
rect 2592 22770 2632 22802
rect 2664 22770 2704 22802
rect 2736 22770 2776 22802
rect 2808 22770 2848 22802
rect 2880 22770 2920 22802
rect 2952 22770 2992 22802
rect 3024 22770 3064 22802
rect 3096 22770 3136 22802
rect 3168 22770 3208 22802
rect 3240 22770 3280 22802
rect 3312 22770 3352 22802
rect 3384 22770 3424 22802
rect 3456 22770 3496 22802
rect 3528 22770 3568 22802
rect 3600 22770 3640 22802
rect 3672 22770 3712 22802
rect 3744 22770 3784 22802
rect 3816 22770 3856 22802
rect 3888 22770 4000 22802
rect 0 22730 4000 22770
rect 0 22698 112 22730
rect 144 22698 184 22730
rect 216 22698 256 22730
rect 288 22698 328 22730
rect 360 22698 400 22730
rect 432 22698 472 22730
rect 504 22698 544 22730
rect 576 22698 616 22730
rect 648 22698 688 22730
rect 720 22698 760 22730
rect 792 22698 832 22730
rect 864 22698 904 22730
rect 936 22698 976 22730
rect 1008 22698 1048 22730
rect 1080 22698 1120 22730
rect 1152 22698 1192 22730
rect 1224 22698 1264 22730
rect 1296 22698 1336 22730
rect 1368 22698 1408 22730
rect 1440 22698 1480 22730
rect 1512 22698 1552 22730
rect 1584 22698 1624 22730
rect 1656 22698 1696 22730
rect 1728 22698 1768 22730
rect 1800 22698 1840 22730
rect 1872 22698 1912 22730
rect 1944 22698 1984 22730
rect 2016 22698 2056 22730
rect 2088 22698 2128 22730
rect 2160 22698 2200 22730
rect 2232 22698 2272 22730
rect 2304 22698 2344 22730
rect 2376 22698 2416 22730
rect 2448 22698 2488 22730
rect 2520 22698 2560 22730
rect 2592 22698 2632 22730
rect 2664 22698 2704 22730
rect 2736 22698 2776 22730
rect 2808 22698 2848 22730
rect 2880 22698 2920 22730
rect 2952 22698 2992 22730
rect 3024 22698 3064 22730
rect 3096 22698 3136 22730
rect 3168 22698 3208 22730
rect 3240 22698 3280 22730
rect 3312 22698 3352 22730
rect 3384 22698 3424 22730
rect 3456 22698 3496 22730
rect 3528 22698 3568 22730
rect 3600 22698 3640 22730
rect 3672 22698 3712 22730
rect 3744 22698 3784 22730
rect 3816 22698 3856 22730
rect 3888 22698 4000 22730
rect 0 22658 4000 22698
rect 0 22626 112 22658
rect 144 22626 184 22658
rect 216 22626 256 22658
rect 288 22626 328 22658
rect 360 22626 400 22658
rect 432 22626 472 22658
rect 504 22626 544 22658
rect 576 22626 616 22658
rect 648 22626 688 22658
rect 720 22626 760 22658
rect 792 22626 832 22658
rect 864 22626 904 22658
rect 936 22626 976 22658
rect 1008 22626 1048 22658
rect 1080 22626 1120 22658
rect 1152 22626 1192 22658
rect 1224 22626 1264 22658
rect 1296 22626 1336 22658
rect 1368 22626 1408 22658
rect 1440 22626 1480 22658
rect 1512 22626 1552 22658
rect 1584 22626 1624 22658
rect 1656 22626 1696 22658
rect 1728 22626 1768 22658
rect 1800 22626 1840 22658
rect 1872 22626 1912 22658
rect 1944 22626 1984 22658
rect 2016 22626 2056 22658
rect 2088 22626 2128 22658
rect 2160 22626 2200 22658
rect 2232 22626 2272 22658
rect 2304 22626 2344 22658
rect 2376 22626 2416 22658
rect 2448 22626 2488 22658
rect 2520 22626 2560 22658
rect 2592 22626 2632 22658
rect 2664 22626 2704 22658
rect 2736 22626 2776 22658
rect 2808 22626 2848 22658
rect 2880 22626 2920 22658
rect 2952 22626 2992 22658
rect 3024 22626 3064 22658
rect 3096 22626 3136 22658
rect 3168 22626 3208 22658
rect 3240 22626 3280 22658
rect 3312 22626 3352 22658
rect 3384 22626 3424 22658
rect 3456 22626 3496 22658
rect 3528 22626 3568 22658
rect 3600 22626 3640 22658
rect 3672 22626 3712 22658
rect 3744 22626 3784 22658
rect 3816 22626 3856 22658
rect 3888 22626 4000 22658
rect 0 22586 4000 22626
rect 0 22554 112 22586
rect 144 22554 184 22586
rect 216 22554 256 22586
rect 288 22554 328 22586
rect 360 22554 400 22586
rect 432 22554 472 22586
rect 504 22554 544 22586
rect 576 22554 616 22586
rect 648 22554 688 22586
rect 720 22554 760 22586
rect 792 22554 832 22586
rect 864 22554 904 22586
rect 936 22554 976 22586
rect 1008 22554 1048 22586
rect 1080 22554 1120 22586
rect 1152 22554 1192 22586
rect 1224 22554 1264 22586
rect 1296 22554 1336 22586
rect 1368 22554 1408 22586
rect 1440 22554 1480 22586
rect 1512 22554 1552 22586
rect 1584 22554 1624 22586
rect 1656 22554 1696 22586
rect 1728 22554 1768 22586
rect 1800 22554 1840 22586
rect 1872 22554 1912 22586
rect 1944 22554 1984 22586
rect 2016 22554 2056 22586
rect 2088 22554 2128 22586
rect 2160 22554 2200 22586
rect 2232 22554 2272 22586
rect 2304 22554 2344 22586
rect 2376 22554 2416 22586
rect 2448 22554 2488 22586
rect 2520 22554 2560 22586
rect 2592 22554 2632 22586
rect 2664 22554 2704 22586
rect 2736 22554 2776 22586
rect 2808 22554 2848 22586
rect 2880 22554 2920 22586
rect 2952 22554 2992 22586
rect 3024 22554 3064 22586
rect 3096 22554 3136 22586
rect 3168 22554 3208 22586
rect 3240 22554 3280 22586
rect 3312 22554 3352 22586
rect 3384 22554 3424 22586
rect 3456 22554 3496 22586
rect 3528 22554 3568 22586
rect 3600 22554 3640 22586
rect 3672 22554 3712 22586
rect 3744 22554 3784 22586
rect 3816 22554 3856 22586
rect 3888 22554 4000 22586
rect 0 22514 4000 22554
rect 0 22482 112 22514
rect 144 22482 184 22514
rect 216 22482 256 22514
rect 288 22482 328 22514
rect 360 22482 400 22514
rect 432 22482 472 22514
rect 504 22482 544 22514
rect 576 22482 616 22514
rect 648 22482 688 22514
rect 720 22482 760 22514
rect 792 22482 832 22514
rect 864 22482 904 22514
rect 936 22482 976 22514
rect 1008 22482 1048 22514
rect 1080 22482 1120 22514
rect 1152 22482 1192 22514
rect 1224 22482 1264 22514
rect 1296 22482 1336 22514
rect 1368 22482 1408 22514
rect 1440 22482 1480 22514
rect 1512 22482 1552 22514
rect 1584 22482 1624 22514
rect 1656 22482 1696 22514
rect 1728 22482 1768 22514
rect 1800 22482 1840 22514
rect 1872 22482 1912 22514
rect 1944 22482 1984 22514
rect 2016 22482 2056 22514
rect 2088 22482 2128 22514
rect 2160 22482 2200 22514
rect 2232 22482 2272 22514
rect 2304 22482 2344 22514
rect 2376 22482 2416 22514
rect 2448 22482 2488 22514
rect 2520 22482 2560 22514
rect 2592 22482 2632 22514
rect 2664 22482 2704 22514
rect 2736 22482 2776 22514
rect 2808 22482 2848 22514
rect 2880 22482 2920 22514
rect 2952 22482 2992 22514
rect 3024 22482 3064 22514
rect 3096 22482 3136 22514
rect 3168 22482 3208 22514
rect 3240 22482 3280 22514
rect 3312 22482 3352 22514
rect 3384 22482 3424 22514
rect 3456 22482 3496 22514
rect 3528 22482 3568 22514
rect 3600 22482 3640 22514
rect 3672 22482 3712 22514
rect 3744 22482 3784 22514
rect 3816 22482 3856 22514
rect 3888 22482 4000 22514
rect 0 22442 4000 22482
rect 0 22410 112 22442
rect 144 22410 184 22442
rect 216 22410 256 22442
rect 288 22410 328 22442
rect 360 22410 400 22442
rect 432 22410 472 22442
rect 504 22410 544 22442
rect 576 22410 616 22442
rect 648 22410 688 22442
rect 720 22410 760 22442
rect 792 22410 832 22442
rect 864 22410 904 22442
rect 936 22410 976 22442
rect 1008 22410 1048 22442
rect 1080 22410 1120 22442
rect 1152 22410 1192 22442
rect 1224 22410 1264 22442
rect 1296 22410 1336 22442
rect 1368 22410 1408 22442
rect 1440 22410 1480 22442
rect 1512 22410 1552 22442
rect 1584 22410 1624 22442
rect 1656 22410 1696 22442
rect 1728 22410 1768 22442
rect 1800 22410 1840 22442
rect 1872 22410 1912 22442
rect 1944 22410 1984 22442
rect 2016 22410 2056 22442
rect 2088 22410 2128 22442
rect 2160 22410 2200 22442
rect 2232 22410 2272 22442
rect 2304 22410 2344 22442
rect 2376 22410 2416 22442
rect 2448 22410 2488 22442
rect 2520 22410 2560 22442
rect 2592 22410 2632 22442
rect 2664 22410 2704 22442
rect 2736 22410 2776 22442
rect 2808 22410 2848 22442
rect 2880 22410 2920 22442
rect 2952 22410 2992 22442
rect 3024 22410 3064 22442
rect 3096 22410 3136 22442
rect 3168 22410 3208 22442
rect 3240 22410 3280 22442
rect 3312 22410 3352 22442
rect 3384 22410 3424 22442
rect 3456 22410 3496 22442
rect 3528 22410 3568 22442
rect 3600 22410 3640 22442
rect 3672 22410 3712 22442
rect 3744 22410 3784 22442
rect 3816 22410 3856 22442
rect 3888 22410 4000 22442
rect 0 22370 4000 22410
rect 0 22338 112 22370
rect 144 22338 184 22370
rect 216 22338 256 22370
rect 288 22338 328 22370
rect 360 22338 400 22370
rect 432 22338 472 22370
rect 504 22338 544 22370
rect 576 22338 616 22370
rect 648 22338 688 22370
rect 720 22338 760 22370
rect 792 22338 832 22370
rect 864 22338 904 22370
rect 936 22338 976 22370
rect 1008 22338 1048 22370
rect 1080 22338 1120 22370
rect 1152 22338 1192 22370
rect 1224 22338 1264 22370
rect 1296 22338 1336 22370
rect 1368 22338 1408 22370
rect 1440 22338 1480 22370
rect 1512 22338 1552 22370
rect 1584 22338 1624 22370
rect 1656 22338 1696 22370
rect 1728 22338 1768 22370
rect 1800 22338 1840 22370
rect 1872 22338 1912 22370
rect 1944 22338 1984 22370
rect 2016 22338 2056 22370
rect 2088 22338 2128 22370
rect 2160 22338 2200 22370
rect 2232 22338 2272 22370
rect 2304 22338 2344 22370
rect 2376 22338 2416 22370
rect 2448 22338 2488 22370
rect 2520 22338 2560 22370
rect 2592 22338 2632 22370
rect 2664 22338 2704 22370
rect 2736 22338 2776 22370
rect 2808 22338 2848 22370
rect 2880 22338 2920 22370
rect 2952 22338 2992 22370
rect 3024 22338 3064 22370
rect 3096 22338 3136 22370
rect 3168 22338 3208 22370
rect 3240 22338 3280 22370
rect 3312 22338 3352 22370
rect 3384 22338 3424 22370
rect 3456 22338 3496 22370
rect 3528 22338 3568 22370
rect 3600 22338 3640 22370
rect 3672 22338 3712 22370
rect 3744 22338 3784 22370
rect 3816 22338 3856 22370
rect 3888 22338 4000 22370
rect 0 22298 4000 22338
rect 0 22266 112 22298
rect 144 22266 184 22298
rect 216 22266 256 22298
rect 288 22266 328 22298
rect 360 22266 400 22298
rect 432 22266 472 22298
rect 504 22266 544 22298
rect 576 22266 616 22298
rect 648 22266 688 22298
rect 720 22266 760 22298
rect 792 22266 832 22298
rect 864 22266 904 22298
rect 936 22266 976 22298
rect 1008 22266 1048 22298
rect 1080 22266 1120 22298
rect 1152 22266 1192 22298
rect 1224 22266 1264 22298
rect 1296 22266 1336 22298
rect 1368 22266 1408 22298
rect 1440 22266 1480 22298
rect 1512 22266 1552 22298
rect 1584 22266 1624 22298
rect 1656 22266 1696 22298
rect 1728 22266 1768 22298
rect 1800 22266 1840 22298
rect 1872 22266 1912 22298
rect 1944 22266 1984 22298
rect 2016 22266 2056 22298
rect 2088 22266 2128 22298
rect 2160 22266 2200 22298
rect 2232 22266 2272 22298
rect 2304 22266 2344 22298
rect 2376 22266 2416 22298
rect 2448 22266 2488 22298
rect 2520 22266 2560 22298
rect 2592 22266 2632 22298
rect 2664 22266 2704 22298
rect 2736 22266 2776 22298
rect 2808 22266 2848 22298
rect 2880 22266 2920 22298
rect 2952 22266 2992 22298
rect 3024 22266 3064 22298
rect 3096 22266 3136 22298
rect 3168 22266 3208 22298
rect 3240 22266 3280 22298
rect 3312 22266 3352 22298
rect 3384 22266 3424 22298
rect 3456 22266 3496 22298
rect 3528 22266 3568 22298
rect 3600 22266 3640 22298
rect 3672 22266 3712 22298
rect 3744 22266 3784 22298
rect 3816 22266 3856 22298
rect 3888 22266 4000 22298
rect 0 22226 4000 22266
rect 0 22194 112 22226
rect 144 22194 184 22226
rect 216 22194 256 22226
rect 288 22194 328 22226
rect 360 22194 400 22226
rect 432 22194 472 22226
rect 504 22194 544 22226
rect 576 22194 616 22226
rect 648 22194 688 22226
rect 720 22194 760 22226
rect 792 22194 832 22226
rect 864 22194 904 22226
rect 936 22194 976 22226
rect 1008 22194 1048 22226
rect 1080 22194 1120 22226
rect 1152 22194 1192 22226
rect 1224 22194 1264 22226
rect 1296 22194 1336 22226
rect 1368 22194 1408 22226
rect 1440 22194 1480 22226
rect 1512 22194 1552 22226
rect 1584 22194 1624 22226
rect 1656 22194 1696 22226
rect 1728 22194 1768 22226
rect 1800 22194 1840 22226
rect 1872 22194 1912 22226
rect 1944 22194 1984 22226
rect 2016 22194 2056 22226
rect 2088 22194 2128 22226
rect 2160 22194 2200 22226
rect 2232 22194 2272 22226
rect 2304 22194 2344 22226
rect 2376 22194 2416 22226
rect 2448 22194 2488 22226
rect 2520 22194 2560 22226
rect 2592 22194 2632 22226
rect 2664 22194 2704 22226
rect 2736 22194 2776 22226
rect 2808 22194 2848 22226
rect 2880 22194 2920 22226
rect 2952 22194 2992 22226
rect 3024 22194 3064 22226
rect 3096 22194 3136 22226
rect 3168 22194 3208 22226
rect 3240 22194 3280 22226
rect 3312 22194 3352 22226
rect 3384 22194 3424 22226
rect 3456 22194 3496 22226
rect 3528 22194 3568 22226
rect 3600 22194 3640 22226
rect 3672 22194 3712 22226
rect 3744 22194 3784 22226
rect 3816 22194 3856 22226
rect 3888 22194 4000 22226
rect 0 22154 4000 22194
rect 0 22122 112 22154
rect 144 22122 184 22154
rect 216 22122 256 22154
rect 288 22122 328 22154
rect 360 22122 400 22154
rect 432 22122 472 22154
rect 504 22122 544 22154
rect 576 22122 616 22154
rect 648 22122 688 22154
rect 720 22122 760 22154
rect 792 22122 832 22154
rect 864 22122 904 22154
rect 936 22122 976 22154
rect 1008 22122 1048 22154
rect 1080 22122 1120 22154
rect 1152 22122 1192 22154
rect 1224 22122 1264 22154
rect 1296 22122 1336 22154
rect 1368 22122 1408 22154
rect 1440 22122 1480 22154
rect 1512 22122 1552 22154
rect 1584 22122 1624 22154
rect 1656 22122 1696 22154
rect 1728 22122 1768 22154
rect 1800 22122 1840 22154
rect 1872 22122 1912 22154
rect 1944 22122 1984 22154
rect 2016 22122 2056 22154
rect 2088 22122 2128 22154
rect 2160 22122 2200 22154
rect 2232 22122 2272 22154
rect 2304 22122 2344 22154
rect 2376 22122 2416 22154
rect 2448 22122 2488 22154
rect 2520 22122 2560 22154
rect 2592 22122 2632 22154
rect 2664 22122 2704 22154
rect 2736 22122 2776 22154
rect 2808 22122 2848 22154
rect 2880 22122 2920 22154
rect 2952 22122 2992 22154
rect 3024 22122 3064 22154
rect 3096 22122 3136 22154
rect 3168 22122 3208 22154
rect 3240 22122 3280 22154
rect 3312 22122 3352 22154
rect 3384 22122 3424 22154
rect 3456 22122 3496 22154
rect 3528 22122 3568 22154
rect 3600 22122 3640 22154
rect 3672 22122 3712 22154
rect 3744 22122 3784 22154
rect 3816 22122 3856 22154
rect 3888 22122 4000 22154
rect 0 22082 4000 22122
rect 0 22050 112 22082
rect 144 22050 184 22082
rect 216 22050 256 22082
rect 288 22050 328 22082
rect 360 22050 400 22082
rect 432 22050 472 22082
rect 504 22050 544 22082
rect 576 22050 616 22082
rect 648 22050 688 22082
rect 720 22050 760 22082
rect 792 22050 832 22082
rect 864 22050 904 22082
rect 936 22050 976 22082
rect 1008 22050 1048 22082
rect 1080 22050 1120 22082
rect 1152 22050 1192 22082
rect 1224 22050 1264 22082
rect 1296 22050 1336 22082
rect 1368 22050 1408 22082
rect 1440 22050 1480 22082
rect 1512 22050 1552 22082
rect 1584 22050 1624 22082
rect 1656 22050 1696 22082
rect 1728 22050 1768 22082
rect 1800 22050 1840 22082
rect 1872 22050 1912 22082
rect 1944 22050 1984 22082
rect 2016 22050 2056 22082
rect 2088 22050 2128 22082
rect 2160 22050 2200 22082
rect 2232 22050 2272 22082
rect 2304 22050 2344 22082
rect 2376 22050 2416 22082
rect 2448 22050 2488 22082
rect 2520 22050 2560 22082
rect 2592 22050 2632 22082
rect 2664 22050 2704 22082
rect 2736 22050 2776 22082
rect 2808 22050 2848 22082
rect 2880 22050 2920 22082
rect 2952 22050 2992 22082
rect 3024 22050 3064 22082
rect 3096 22050 3136 22082
rect 3168 22050 3208 22082
rect 3240 22050 3280 22082
rect 3312 22050 3352 22082
rect 3384 22050 3424 22082
rect 3456 22050 3496 22082
rect 3528 22050 3568 22082
rect 3600 22050 3640 22082
rect 3672 22050 3712 22082
rect 3744 22050 3784 22082
rect 3816 22050 3856 22082
rect 3888 22050 4000 22082
rect 0 22010 4000 22050
rect 0 21978 112 22010
rect 144 21978 184 22010
rect 216 21978 256 22010
rect 288 21978 328 22010
rect 360 21978 400 22010
rect 432 21978 472 22010
rect 504 21978 544 22010
rect 576 21978 616 22010
rect 648 21978 688 22010
rect 720 21978 760 22010
rect 792 21978 832 22010
rect 864 21978 904 22010
rect 936 21978 976 22010
rect 1008 21978 1048 22010
rect 1080 21978 1120 22010
rect 1152 21978 1192 22010
rect 1224 21978 1264 22010
rect 1296 21978 1336 22010
rect 1368 21978 1408 22010
rect 1440 21978 1480 22010
rect 1512 21978 1552 22010
rect 1584 21978 1624 22010
rect 1656 21978 1696 22010
rect 1728 21978 1768 22010
rect 1800 21978 1840 22010
rect 1872 21978 1912 22010
rect 1944 21978 1984 22010
rect 2016 21978 2056 22010
rect 2088 21978 2128 22010
rect 2160 21978 2200 22010
rect 2232 21978 2272 22010
rect 2304 21978 2344 22010
rect 2376 21978 2416 22010
rect 2448 21978 2488 22010
rect 2520 21978 2560 22010
rect 2592 21978 2632 22010
rect 2664 21978 2704 22010
rect 2736 21978 2776 22010
rect 2808 21978 2848 22010
rect 2880 21978 2920 22010
rect 2952 21978 2992 22010
rect 3024 21978 3064 22010
rect 3096 21978 3136 22010
rect 3168 21978 3208 22010
rect 3240 21978 3280 22010
rect 3312 21978 3352 22010
rect 3384 21978 3424 22010
rect 3456 21978 3496 22010
rect 3528 21978 3568 22010
rect 3600 21978 3640 22010
rect 3672 21978 3712 22010
rect 3744 21978 3784 22010
rect 3816 21978 3856 22010
rect 3888 21978 4000 22010
rect 0 21938 4000 21978
rect 0 21906 112 21938
rect 144 21906 184 21938
rect 216 21906 256 21938
rect 288 21906 328 21938
rect 360 21906 400 21938
rect 432 21906 472 21938
rect 504 21906 544 21938
rect 576 21906 616 21938
rect 648 21906 688 21938
rect 720 21906 760 21938
rect 792 21906 832 21938
rect 864 21906 904 21938
rect 936 21906 976 21938
rect 1008 21906 1048 21938
rect 1080 21906 1120 21938
rect 1152 21906 1192 21938
rect 1224 21906 1264 21938
rect 1296 21906 1336 21938
rect 1368 21906 1408 21938
rect 1440 21906 1480 21938
rect 1512 21906 1552 21938
rect 1584 21906 1624 21938
rect 1656 21906 1696 21938
rect 1728 21906 1768 21938
rect 1800 21906 1840 21938
rect 1872 21906 1912 21938
rect 1944 21906 1984 21938
rect 2016 21906 2056 21938
rect 2088 21906 2128 21938
rect 2160 21906 2200 21938
rect 2232 21906 2272 21938
rect 2304 21906 2344 21938
rect 2376 21906 2416 21938
rect 2448 21906 2488 21938
rect 2520 21906 2560 21938
rect 2592 21906 2632 21938
rect 2664 21906 2704 21938
rect 2736 21906 2776 21938
rect 2808 21906 2848 21938
rect 2880 21906 2920 21938
rect 2952 21906 2992 21938
rect 3024 21906 3064 21938
rect 3096 21906 3136 21938
rect 3168 21906 3208 21938
rect 3240 21906 3280 21938
rect 3312 21906 3352 21938
rect 3384 21906 3424 21938
rect 3456 21906 3496 21938
rect 3528 21906 3568 21938
rect 3600 21906 3640 21938
rect 3672 21906 3712 21938
rect 3744 21906 3784 21938
rect 3816 21906 3856 21938
rect 3888 21906 4000 21938
rect 0 21866 4000 21906
rect 0 21834 112 21866
rect 144 21834 184 21866
rect 216 21834 256 21866
rect 288 21834 328 21866
rect 360 21834 400 21866
rect 432 21834 472 21866
rect 504 21834 544 21866
rect 576 21834 616 21866
rect 648 21834 688 21866
rect 720 21834 760 21866
rect 792 21834 832 21866
rect 864 21834 904 21866
rect 936 21834 976 21866
rect 1008 21834 1048 21866
rect 1080 21834 1120 21866
rect 1152 21834 1192 21866
rect 1224 21834 1264 21866
rect 1296 21834 1336 21866
rect 1368 21834 1408 21866
rect 1440 21834 1480 21866
rect 1512 21834 1552 21866
rect 1584 21834 1624 21866
rect 1656 21834 1696 21866
rect 1728 21834 1768 21866
rect 1800 21834 1840 21866
rect 1872 21834 1912 21866
rect 1944 21834 1984 21866
rect 2016 21834 2056 21866
rect 2088 21834 2128 21866
rect 2160 21834 2200 21866
rect 2232 21834 2272 21866
rect 2304 21834 2344 21866
rect 2376 21834 2416 21866
rect 2448 21834 2488 21866
rect 2520 21834 2560 21866
rect 2592 21834 2632 21866
rect 2664 21834 2704 21866
rect 2736 21834 2776 21866
rect 2808 21834 2848 21866
rect 2880 21834 2920 21866
rect 2952 21834 2992 21866
rect 3024 21834 3064 21866
rect 3096 21834 3136 21866
rect 3168 21834 3208 21866
rect 3240 21834 3280 21866
rect 3312 21834 3352 21866
rect 3384 21834 3424 21866
rect 3456 21834 3496 21866
rect 3528 21834 3568 21866
rect 3600 21834 3640 21866
rect 3672 21834 3712 21866
rect 3744 21834 3784 21866
rect 3816 21834 3856 21866
rect 3888 21834 4000 21866
rect 0 21794 4000 21834
rect 0 21762 112 21794
rect 144 21762 184 21794
rect 216 21762 256 21794
rect 288 21762 328 21794
rect 360 21762 400 21794
rect 432 21762 472 21794
rect 504 21762 544 21794
rect 576 21762 616 21794
rect 648 21762 688 21794
rect 720 21762 760 21794
rect 792 21762 832 21794
rect 864 21762 904 21794
rect 936 21762 976 21794
rect 1008 21762 1048 21794
rect 1080 21762 1120 21794
rect 1152 21762 1192 21794
rect 1224 21762 1264 21794
rect 1296 21762 1336 21794
rect 1368 21762 1408 21794
rect 1440 21762 1480 21794
rect 1512 21762 1552 21794
rect 1584 21762 1624 21794
rect 1656 21762 1696 21794
rect 1728 21762 1768 21794
rect 1800 21762 1840 21794
rect 1872 21762 1912 21794
rect 1944 21762 1984 21794
rect 2016 21762 2056 21794
rect 2088 21762 2128 21794
rect 2160 21762 2200 21794
rect 2232 21762 2272 21794
rect 2304 21762 2344 21794
rect 2376 21762 2416 21794
rect 2448 21762 2488 21794
rect 2520 21762 2560 21794
rect 2592 21762 2632 21794
rect 2664 21762 2704 21794
rect 2736 21762 2776 21794
rect 2808 21762 2848 21794
rect 2880 21762 2920 21794
rect 2952 21762 2992 21794
rect 3024 21762 3064 21794
rect 3096 21762 3136 21794
rect 3168 21762 3208 21794
rect 3240 21762 3280 21794
rect 3312 21762 3352 21794
rect 3384 21762 3424 21794
rect 3456 21762 3496 21794
rect 3528 21762 3568 21794
rect 3600 21762 3640 21794
rect 3672 21762 3712 21794
rect 3744 21762 3784 21794
rect 3816 21762 3856 21794
rect 3888 21762 4000 21794
rect 0 21722 4000 21762
rect 0 21690 112 21722
rect 144 21690 184 21722
rect 216 21690 256 21722
rect 288 21690 328 21722
rect 360 21690 400 21722
rect 432 21690 472 21722
rect 504 21690 544 21722
rect 576 21690 616 21722
rect 648 21690 688 21722
rect 720 21690 760 21722
rect 792 21690 832 21722
rect 864 21690 904 21722
rect 936 21690 976 21722
rect 1008 21690 1048 21722
rect 1080 21690 1120 21722
rect 1152 21690 1192 21722
rect 1224 21690 1264 21722
rect 1296 21690 1336 21722
rect 1368 21690 1408 21722
rect 1440 21690 1480 21722
rect 1512 21690 1552 21722
rect 1584 21690 1624 21722
rect 1656 21690 1696 21722
rect 1728 21690 1768 21722
rect 1800 21690 1840 21722
rect 1872 21690 1912 21722
rect 1944 21690 1984 21722
rect 2016 21690 2056 21722
rect 2088 21690 2128 21722
rect 2160 21690 2200 21722
rect 2232 21690 2272 21722
rect 2304 21690 2344 21722
rect 2376 21690 2416 21722
rect 2448 21690 2488 21722
rect 2520 21690 2560 21722
rect 2592 21690 2632 21722
rect 2664 21690 2704 21722
rect 2736 21690 2776 21722
rect 2808 21690 2848 21722
rect 2880 21690 2920 21722
rect 2952 21690 2992 21722
rect 3024 21690 3064 21722
rect 3096 21690 3136 21722
rect 3168 21690 3208 21722
rect 3240 21690 3280 21722
rect 3312 21690 3352 21722
rect 3384 21690 3424 21722
rect 3456 21690 3496 21722
rect 3528 21690 3568 21722
rect 3600 21690 3640 21722
rect 3672 21690 3712 21722
rect 3744 21690 3784 21722
rect 3816 21690 3856 21722
rect 3888 21690 4000 21722
rect 0 21650 4000 21690
rect 0 21618 112 21650
rect 144 21618 184 21650
rect 216 21618 256 21650
rect 288 21618 328 21650
rect 360 21618 400 21650
rect 432 21618 472 21650
rect 504 21618 544 21650
rect 576 21618 616 21650
rect 648 21618 688 21650
rect 720 21618 760 21650
rect 792 21618 832 21650
rect 864 21618 904 21650
rect 936 21618 976 21650
rect 1008 21618 1048 21650
rect 1080 21618 1120 21650
rect 1152 21618 1192 21650
rect 1224 21618 1264 21650
rect 1296 21618 1336 21650
rect 1368 21618 1408 21650
rect 1440 21618 1480 21650
rect 1512 21618 1552 21650
rect 1584 21618 1624 21650
rect 1656 21618 1696 21650
rect 1728 21618 1768 21650
rect 1800 21618 1840 21650
rect 1872 21618 1912 21650
rect 1944 21618 1984 21650
rect 2016 21618 2056 21650
rect 2088 21618 2128 21650
rect 2160 21618 2200 21650
rect 2232 21618 2272 21650
rect 2304 21618 2344 21650
rect 2376 21618 2416 21650
rect 2448 21618 2488 21650
rect 2520 21618 2560 21650
rect 2592 21618 2632 21650
rect 2664 21618 2704 21650
rect 2736 21618 2776 21650
rect 2808 21618 2848 21650
rect 2880 21618 2920 21650
rect 2952 21618 2992 21650
rect 3024 21618 3064 21650
rect 3096 21618 3136 21650
rect 3168 21618 3208 21650
rect 3240 21618 3280 21650
rect 3312 21618 3352 21650
rect 3384 21618 3424 21650
rect 3456 21618 3496 21650
rect 3528 21618 3568 21650
rect 3600 21618 3640 21650
rect 3672 21618 3712 21650
rect 3744 21618 3784 21650
rect 3816 21618 3856 21650
rect 3888 21618 4000 21650
rect 0 21578 4000 21618
rect 0 21546 112 21578
rect 144 21546 184 21578
rect 216 21546 256 21578
rect 288 21546 328 21578
rect 360 21546 400 21578
rect 432 21546 472 21578
rect 504 21546 544 21578
rect 576 21546 616 21578
rect 648 21546 688 21578
rect 720 21546 760 21578
rect 792 21546 832 21578
rect 864 21546 904 21578
rect 936 21546 976 21578
rect 1008 21546 1048 21578
rect 1080 21546 1120 21578
rect 1152 21546 1192 21578
rect 1224 21546 1264 21578
rect 1296 21546 1336 21578
rect 1368 21546 1408 21578
rect 1440 21546 1480 21578
rect 1512 21546 1552 21578
rect 1584 21546 1624 21578
rect 1656 21546 1696 21578
rect 1728 21546 1768 21578
rect 1800 21546 1840 21578
rect 1872 21546 1912 21578
rect 1944 21546 1984 21578
rect 2016 21546 2056 21578
rect 2088 21546 2128 21578
rect 2160 21546 2200 21578
rect 2232 21546 2272 21578
rect 2304 21546 2344 21578
rect 2376 21546 2416 21578
rect 2448 21546 2488 21578
rect 2520 21546 2560 21578
rect 2592 21546 2632 21578
rect 2664 21546 2704 21578
rect 2736 21546 2776 21578
rect 2808 21546 2848 21578
rect 2880 21546 2920 21578
rect 2952 21546 2992 21578
rect 3024 21546 3064 21578
rect 3096 21546 3136 21578
rect 3168 21546 3208 21578
rect 3240 21546 3280 21578
rect 3312 21546 3352 21578
rect 3384 21546 3424 21578
rect 3456 21546 3496 21578
rect 3528 21546 3568 21578
rect 3600 21546 3640 21578
rect 3672 21546 3712 21578
rect 3744 21546 3784 21578
rect 3816 21546 3856 21578
rect 3888 21546 4000 21578
rect 0 21506 4000 21546
rect 0 21474 112 21506
rect 144 21474 184 21506
rect 216 21474 256 21506
rect 288 21474 328 21506
rect 360 21474 400 21506
rect 432 21474 472 21506
rect 504 21474 544 21506
rect 576 21474 616 21506
rect 648 21474 688 21506
rect 720 21474 760 21506
rect 792 21474 832 21506
rect 864 21474 904 21506
rect 936 21474 976 21506
rect 1008 21474 1048 21506
rect 1080 21474 1120 21506
rect 1152 21474 1192 21506
rect 1224 21474 1264 21506
rect 1296 21474 1336 21506
rect 1368 21474 1408 21506
rect 1440 21474 1480 21506
rect 1512 21474 1552 21506
rect 1584 21474 1624 21506
rect 1656 21474 1696 21506
rect 1728 21474 1768 21506
rect 1800 21474 1840 21506
rect 1872 21474 1912 21506
rect 1944 21474 1984 21506
rect 2016 21474 2056 21506
rect 2088 21474 2128 21506
rect 2160 21474 2200 21506
rect 2232 21474 2272 21506
rect 2304 21474 2344 21506
rect 2376 21474 2416 21506
rect 2448 21474 2488 21506
rect 2520 21474 2560 21506
rect 2592 21474 2632 21506
rect 2664 21474 2704 21506
rect 2736 21474 2776 21506
rect 2808 21474 2848 21506
rect 2880 21474 2920 21506
rect 2952 21474 2992 21506
rect 3024 21474 3064 21506
rect 3096 21474 3136 21506
rect 3168 21474 3208 21506
rect 3240 21474 3280 21506
rect 3312 21474 3352 21506
rect 3384 21474 3424 21506
rect 3456 21474 3496 21506
rect 3528 21474 3568 21506
rect 3600 21474 3640 21506
rect 3672 21474 3712 21506
rect 3744 21474 3784 21506
rect 3816 21474 3856 21506
rect 3888 21474 4000 21506
rect 0 21434 4000 21474
rect 0 21402 112 21434
rect 144 21402 184 21434
rect 216 21402 256 21434
rect 288 21402 328 21434
rect 360 21402 400 21434
rect 432 21402 472 21434
rect 504 21402 544 21434
rect 576 21402 616 21434
rect 648 21402 688 21434
rect 720 21402 760 21434
rect 792 21402 832 21434
rect 864 21402 904 21434
rect 936 21402 976 21434
rect 1008 21402 1048 21434
rect 1080 21402 1120 21434
rect 1152 21402 1192 21434
rect 1224 21402 1264 21434
rect 1296 21402 1336 21434
rect 1368 21402 1408 21434
rect 1440 21402 1480 21434
rect 1512 21402 1552 21434
rect 1584 21402 1624 21434
rect 1656 21402 1696 21434
rect 1728 21402 1768 21434
rect 1800 21402 1840 21434
rect 1872 21402 1912 21434
rect 1944 21402 1984 21434
rect 2016 21402 2056 21434
rect 2088 21402 2128 21434
rect 2160 21402 2200 21434
rect 2232 21402 2272 21434
rect 2304 21402 2344 21434
rect 2376 21402 2416 21434
rect 2448 21402 2488 21434
rect 2520 21402 2560 21434
rect 2592 21402 2632 21434
rect 2664 21402 2704 21434
rect 2736 21402 2776 21434
rect 2808 21402 2848 21434
rect 2880 21402 2920 21434
rect 2952 21402 2992 21434
rect 3024 21402 3064 21434
rect 3096 21402 3136 21434
rect 3168 21402 3208 21434
rect 3240 21402 3280 21434
rect 3312 21402 3352 21434
rect 3384 21402 3424 21434
rect 3456 21402 3496 21434
rect 3528 21402 3568 21434
rect 3600 21402 3640 21434
rect 3672 21402 3712 21434
rect 3744 21402 3784 21434
rect 3816 21402 3856 21434
rect 3888 21402 4000 21434
rect 0 21362 4000 21402
rect 0 21330 112 21362
rect 144 21330 184 21362
rect 216 21330 256 21362
rect 288 21330 328 21362
rect 360 21330 400 21362
rect 432 21330 472 21362
rect 504 21330 544 21362
rect 576 21330 616 21362
rect 648 21330 688 21362
rect 720 21330 760 21362
rect 792 21330 832 21362
rect 864 21330 904 21362
rect 936 21330 976 21362
rect 1008 21330 1048 21362
rect 1080 21330 1120 21362
rect 1152 21330 1192 21362
rect 1224 21330 1264 21362
rect 1296 21330 1336 21362
rect 1368 21330 1408 21362
rect 1440 21330 1480 21362
rect 1512 21330 1552 21362
rect 1584 21330 1624 21362
rect 1656 21330 1696 21362
rect 1728 21330 1768 21362
rect 1800 21330 1840 21362
rect 1872 21330 1912 21362
rect 1944 21330 1984 21362
rect 2016 21330 2056 21362
rect 2088 21330 2128 21362
rect 2160 21330 2200 21362
rect 2232 21330 2272 21362
rect 2304 21330 2344 21362
rect 2376 21330 2416 21362
rect 2448 21330 2488 21362
rect 2520 21330 2560 21362
rect 2592 21330 2632 21362
rect 2664 21330 2704 21362
rect 2736 21330 2776 21362
rect 2808 21330 2848 21362
rect 2880 21330 2920 21362
rect 2952 21330 2992 21362
rect 3024 21330 3064 21362
rect 3096 21330 3136 21362
rect 3168 21330 3208 21362
rect 3240 21330 3280 21362
rect 3312 21330 3352 21362
rect 3384 21330 3424 21362
rect 3456 21330 3496 21362
rect 3528 21330 3568 21362
rect 3600 21330 3640 21362
rect 3672 21330 3712 21362
rect 3744 21330 3784 21362
rect 3816 21330 3856 21362
rect 3888 21330 4000 21362
rect 0 21290 4000 21330
rect 0 21258 112 21290
rect 144 21258 184 21290
rect 216 21258 256 21290
rect 288 21258 328 21290
rect 360 21258 400 21290
rect 432 21258 472 21290
rect 504 21258 544 21290
rect 576 21258 616 21290
rect 648 21258 688 21290
rect 720 21258 760 21290
rect 792 21258 832 21290
rect 864 21258 904 21290
rect 936 21258 976 21290
rect 1008 21258 1048 21290
rect 1080 21258 1120 21290
rect 1152 21258 1192 21290
rect 1224 21258 1264 21290
rect 1296 21258 1336 21290
rect 1368 21258 1408 21290
rect 1440 21258 1480 21290
rect 1512 21258 1552 21290
rect 1584 21258 1624 21290
rect 1656 21258 1696 21290
rect 1728 21258 1768 21290
rect 1800 21258 1840 21290
rect 1872 21258 1912 21290
rect 1944 21258 1984 21290
rect 2016 21258 2056 21290
rect 2088 21258 2128 21290
rect 2160 21258 2200 21290
rect 2232 21258 2272 21290
rect 2304 21258 2344 21290
rect 2376 21258 2416 21290
rect 2448 21258 2488 21290
rect 2520 21258 2560 21290
rect 2592 21258 2632 21290
rect 2664 21258 2704 21290
rect 2736 21258 2776 21290
rect 2808 21258 2848 21290
rect 2880 21258 2920 21290
rect 2952 21258 2992 21290
rect 3024 21258 3064 21290
rect 3096 21258 3136 21290
rect 3168 21258 3208 21290
rect 3240 21258 3280 21290
rect 3312 21258 3352 21290
rect 3384 21258 3424 21290
rect 3456 21258 3496 21290
rect 3528 21258 3568 21290
rect 3600 21258 3640 21290
rect 3672 21258 3712 21290
rect 3744 21258 3784 21290
rect 3816 21258 3856 21290
rect 3888 21258 4000 21290
rect 0 21218 4000 21258
rect 0 21186 112 21218
rect 144 21186 184 21218
rect 216 21186 256 21218
rect 288 21186 328 21218
rect 360 21186 400 21218
rect 432 21186 472 21218
rect 504 21186 544 21218
rect 576 21186 616 21218
rect 648 21186 688 21218
rect 720 21186 760 21218
rect 792 21186 832 21218
rect 864 21186 904 21218
rect 936 21186 976 21218
rect 1008 21186 1048 21218
rect 1080 21186 1120 21218
rect 1152 21186 1192 21218
rect 1224 21186 1264 21218
rect 1296 21186 1336 21218
rect 1368 21186 1408 21218
rect 1440 21186 1480 21218
rect 1512 21186 1552 21218
rect 1584 21186 1624 21218
rect 1656 21186 1696 21218
rect 1728 21186 1768 21218
rect 1800 21186 1840 21218
rect 1872 21186 1912 21218
rect 1944 21186 1984 21218
rect 2016 21186 2056 21218
rect 2088 21186 2128 21218
rect 2160 21186 2200 21218
rect 2232 21186 2272 21218
rect 2304 21186 2344 21218
rect 2376 21186 2416 21218
rect 2448 21186 2488 21218
rect 2520 21186 2560 21218
rect 2592 21186 2632 21218
rect 2664 21186 2704 21218
rect 2736 21186 2776 21218
rect 2808 21186 2848 21218
rect 2880 21186 2920 21218
rect 2952 21186 2992 21218
rect 3024 21186 3064 21218
rect 3096 21186 3136 21218
rect 3168 21186 3208 21218
rect 3240 21186 3280 21218
rect 3312 21186 3352 21218
rect 3384 21186 3424 21218
rect 3456 21186 3496 21218
rect 3528 21186 3568 21218
rect 3600 21186 3640 21218
rect 3672 21186 3712 21218
rect 3744 21186 3784 21218
rect 3816 21186 3856 21218
rect 3888 21186 4000 21218
rect 0 21146 4000 21186
rect 0 21114 112 21146
rect 144 21114 184 21146
rect 216 21114 256 21146
rect 288 21114 328 21146
rect 360 21114 400 21146
rect 432 21114 472 21146
rect 504 21114 544 21146
rect 576 21114 616 21146
rect 648 21114 688 21146
rect 720 21114 760 21146
rect 792 21114 832 21146
rect 864 21114 904 21146
rect 936 21114 976 21146
rect 1008 21114 1048 21146
rect 1080 21114 1120 21146
rect 1152 21114 1192 21146
rect 1224 21114 1264 21146
rect 1296 21114 1336 21146
rect 1368 21114 1408 21146
rect 1440 21114 1480 21146
rect 1512 21114 1552 21146
rect 1584 21114 1624 21146
rect 1656 21114 1696 21146
rect 1728 21114 1768 21146
rect 1800 21114 1840 21146
rect 1872 21114 1912 21146
rect 1944 21114 1984 21146
rect 2016 21114 2056 21146
rect 2088 21114 2128 21146
rect 2160 21114 2200 21146
rect 2232 21114 2272 21146
rect 2304 21114 2344 21146
rect 2376 21114 2416 21146
rect 2448 21114 2488 21146
rect 2520 21114 2560 21146
rect 2592 21114 2632 21146
rect 2664 21114 2704 21146
rect 2736 21114 2776 21146
rect 2808 21114 2848 21146
rect 2880 21114 2920 21146
rect 2952 21114 2992 21146
rect 3024 21114 3064 21146
rect 3096 21114 3136 21146
rect 3168 21114 3208 21146
rect 3240 21114 3280 21146
rect 3312 21114 3352 21146
rect 3384 21114 3424 21146
rect 3456 21114 3496 21146
rect 3528 21114 3568 21146
rect 3600 21114 3640 21146
rect 3672 21114 3712 21146
rect 3744 21114 3784 21146
rect 3816 21114 3856 21146
rect 3888 21114 4000 21146
rect 0 21074 4000 21114
rect 0 21042 112 21074
rect 144 21042 184 21074
rect 216 21042 256 21074
rect 288 21042 328 21074
rect 360 21042 400 21074
rect 432 21042 472 21074
rect 504 21042 544 21074
rect 576 21042 616 21074
rect 648 21042 688 21074
rect 720 21042 760 21074
rect 792 21042 832 21074
rect 864 21042 904 21074
rect 936 21042 976 21074
rect 1008 21042 1048 21074
rect 1080 21042 1120 21074
rect 1152 21042 1192 21074
rect 1224 21042 1264 21074
rect 1296 21042 1336 21074
rect 1368 21042 1408 21074
rect 1440 21042 1480 21074
rect 1512 21042 1552 21074
rect 1584 21042 1624 21074
rect 1656 21042 1696 21074
rect 1728 21042 1768 21074
rect 1800 21042 1840 21074
rect 1872 21042 1912 21074
rect 1944 21042 1984 21074
rect 2016 21042 2056 21074
rect 2088 21042 2128 21074
rect 2160 21042 2200 21074
rect 2232 21042 2272 21074
rect 2304 21042 2344 21074
rect 2376 21042 2416 21074
rect 2448 21042 2488 21074
rect 2520 21042 2560 21074
rect 2592 21042 2632 21074
rect 2664 21042 2704 21074
rect 2736 21042 2776 21074
rect 2808 21042 2848 21074
rect 2880 21042 2920 21074
rect 2952 21042 2992 21074
rect 3024 21042 3064 21074
rect 3096 21042 3136 21074
rect 3168 21042 3208 21074
rect 3240 21042 3280 21074
rect 3312 21042 3352 21074
rect 3384 21042 3424 21074
rect 3456 21042 3496 21074
rect 3528 21042 3568 21074
rect 3600 21042 3640 21074
rect 3672 21042 3712 21074
rect 3744 21042 3784 21074
rect 3816 21042 3856 21074
rect 3888 21042 4000 21074
rect 0 21002 4000 21042
rect 0 20970 112 21002
rect 144 20970 184 21002
rect 216 20970 256 21002
rect 288 20970 328 21002
rect 360 20970 400 21002
rect 432 20970 472 21002
rect 504 20970 544 21002
rect 576 20970 616 21002
rect 648 20970 688 21002
rect 720 20970 760 21002
rect 792 20970 832 21002
rect 864 20970 904 21002
rect 936 20970 976 21002
rect 1008 20970 1048 21002
rect 1080 20970 1120 21002
rect 1152 20970 1192 21002
rect 1224 20970 1264 21002
rect 1296 20970 1336 21002
rect 1368 20970 1408 21002
rect 1440 20970 1480 21002
rect 1512 20970 1552 21002
rect 1584 20970 1624 21002
rect 1656 20970 1696 21002
rect 1728 20970 1768 21002
rect 1800 20970 1840 21002
rect 1872 20970 1912 21002
rect 1944 20970 1984 21002
rect 2016 20970 2056 21002
rect 2088 20970 2128 21002
rect 2160 20970 2200 21002
rect 2232 20970 2272 21002
rect 2304 20970 2344 21002
rect 2376 20970 2416 21002
rect 2448 20970 2488 21002
rect 2520 20970 2560 21002
rect 2592 20970 2632 21002
rect 2664 20970 2704 21002
rect 2736 20970 2776 21002
rect 2808 20970 2848 21002
rect 2880 20970 2920 21002
rect 2952 20970 2992 21002
rect 3024 20970 3064 21002
rect 3096 20970 3136 21002
rect 3168 20970 3208 21002
rect 3240 20970 3280 21002
rect 3312 20970 3352 21002
rect 3384 20970 3424 21002
rect 3456 20970 3496 21002
rect 3528 20970 3568 21002
rect 3600 20970 3640 21002
rect 3672 20970 3712 21002
rect 3744 20970 3784 21002
rect 3816 20970 3856 21002
rect 3888 20970 4000 21002
rect 0 20930 4000 20970
rect 0 20898 112 20930
rect 144 20898 184 20930
rect 216 20898 256 20930
rect 288 20898 328 20930
rect 360 20898 400 20930
rect 432 20898 472 20930
rect 504 20898 544 20930
rect 576 20898 616 20930
rect 648 20898 688 20930
rect 720 20898 760 20930
rect 792 20898 832 20930
rect 864 20898 904 20930
rect 936 20898 976 20930
rect 1008 20898 1048 20930
rect 1080 20898 1120 20930
rect 1152 20898 1192 20930
rect 1224 20898 1264 20930
rect 1296 20898 1336 20930
rect 1368 20898 1408 20930
rect 1440 20898 1480 20930
rect 1512 20898 1552 20930
rect 1584 20898 1624 20930
rect 1656 20898 1696 20930
rect 1728 20898 1768 20930
rect 1800 20898 1840 20930
rect 1872 20898 1912 20930
rect 1944 20898 1984 20930
rect 2016 20898 2056 20930
rect 2088 20898 2128 20930
rect 2160 20898 2200 20930
rect 2232 20898 2272 20930
rect 2304 20898 2344 20930
rect 2376 20898 2416 20930
rect 2448 20898 2488 20930
rect 2520 20898 2560 20930
rect 2592 20898 2632 20930
rect 2664 20898 2704 20930
rect 2736 20898 2776 20930
rect 2808 20898 2848 20930
rect 2880 20898 2920 20930
rect 2952 20898 2992 20930
rect 3024 20898 3064 20930
rect 3096 20898 3136 20930
rect 3168 20898 3208 20930
rect 3240 20898 3280 20930
rect 3312 20898 3352 20930
rect 3384 20898 3424 20930
rect 3456 20898 3496 20930
rect 3528 20898 3568 20930
rect 3600 20898 3640 20930
rect 3672 20898 3712 20930
rect 3744 20898 3784 20930
rect 3816 20898 3856 20930
rect 3888 20898 4000 20930
rect 0 20858 4000 20898
rect 0 20826 112 20858
rect 144 20826 184 20858
rect 216 20826 256 20858
rect 288 20826 328 20858
rect 360 20826 400 20858
rect 432 20826 472 20858
rect 504 20826 544 20858
rect 576 20826 616 20858
rect 648 20826 688 20858
rect 720 20826 760 20858
rect 792 20826 832 20858
rect 864 20826 904 20858
rect 936 20826 976 20858
rect 1008 20826 1048 20858
rect 1080 20826 1120 20858
rect 1152 20826 1192 20858
rect 1224 20826 1264 20858
rect 1296 20826 1336 20858
rect 1368 20826 1408 20858
rect 1440 20826 1480 20858
rect 1512 20826 1552 20858
rect 1584 20826 1624 20858
rect 1656 20826 1696 20858
rect 1728 20826 1768 20858
rect 1800 20826 1840 20858
rect 1872 20826 1912 20858
rect 1944 20826 1984 20858
rect 2016 20826 2056 20858
rect 2088 20826 2128 20858
rect 2160 20826 2200 20858
rect 2232 20826 2272 20858
rect 2304 20826 2344 20858
rect 2376 20826 2416 20858
rect 2448 20826 2488 20858
rect 2520 20826 2560 20858
rect 2592 20826 2632 20858
rect 2664 20826 2704 20858
rect 2736 20826 2776 20858
rect 2808 20826 2848 20858
rect 2880 20826 2920 20858
rect 2952 20826 2992 20858
rect 3024 20826 3064 20858
rect 3096 20826 3136 20858
rect 3168 20826 3208 20858
rect 3240 20826 3280 20858
rect 3312 20826 3352 20858
rect 3384 20826 3424 20858
rect 3456 20826 3496 20858
rect 3528 20826 3568 20858
rect 3600 20826 3640 20858
rect 3672 20826 3712 20858
rect 3744 20826 3784 20858
rect 3816 20826 3856 20858
rect 3888 20826 4000 20858
rect 0 20786 4000 20826
rect 0 20754 112 20786
rect 144 20754 184 20786
rect 216 20754 256 20786
rect 288 20754 328 20786
rect 360 20754 400 20786
rect 432 20754 472 20786
rect 504 20754 544 20786
rect 576 20754 616 20786
rect 648 20754 688 20786
rect 720 20754 760 20786
rect 792 20754 832 20786
rect 864 20754 904 20786
rect 936 20754 976 20786
rect 1008 20754 1048 20786
rect 1080 20754 1120 20786
rect 1152 20754 1192 20786
rect 1224 20754 1264 20786
rect 1296 20754 1336 20786
rect 1368 20754 1408 20786
rect 1440 20754 1480 20786
rect 1512 20754 1552 20786
rect 1584 20754 1624 20786
rect 1656 20754 1696 20786
rect 1728 20754 1768 20786
rect 1800 20754 1840 20786
rect 1872 20754 1912 20786
rect 1944 20754 1984 20786
rect 2016 20754 2056 20786
rect 2088 20754 2128 20786
rect 2160 20754 2200 20786
rect 2232 20754 2272 20786
rect 2304 20754 2344 20786
rect 2376 20754 2416 20786
rect 2448 20754 2488 20786
rect 2520 20754 2560 20786
rect 2592 20754 2632 20786
rect 2664 20754 2704 20786
rect 2736 20754 2776 20786
rect 2808 20754 2848 20786
rect 2880 20754 2920 20786
rect 2952 20754 2992 20786
rect 3024 20754 3064 20786
rect 3096 20754 3136 20786
rect 3168 20754 3208 20786
rect 3240 20754 3280 20786
rect 3312 20754 3352 20786
rect 3384 20754 3424 20786
rect 3456 20754 3496 20786
rect 3528 20754 3568 20786
rect 3600 20754 3640 20786
rect 3672 20754 3712 20786
rect 3744 20754 3784 20786
rect 3816 20754 3856 20786
rect 3888 20754 4000 20786
rect 0 20714 4000 20754
rect 0 20682 112 20714
rect 144 20682 184 20714
rect 216 20682 256 20714
rect 288 20682 328 20714
rect 360 20682 400 20714
rect 432 20682 472 20714
rect 504 20682 544 20714
rect 576 20682 616 20714
rect 648 20682 688 20714
rect 720 20682 760 20714
rect 792 20682 832 20714
rect 864 20682 904 20714
rect 936 20682 976 20714
rect 1008 20682 1048 20714
rect 1080 20682 1120 20714
rect 1152 20682 1192 20714
rect 1224 20682 1264 20714
rect 1296 20682 1336 20714
rect 1368 20682 1408 20714
rect 1440 20682 1480 20714
rect 1512 20682 1552 20714
rect 1584 20682 1624 20714
rect 1656 20682 1696 20714
rect 1728 20682 1768 20714
rect 1800 20682 1840 20714
rect 1872 20682 1912 20714
rect 1944 20682 1984 20714
rect 2016 20682 2056 20714
rect 2088 20682 2128 20714
rect 2160 20682 2200 20714
rect 2232 20682 2272 20714
rect 2304 20682 2344 20714
rect 2376 20682 2416 20714
rect 2448 20682 2488 20714
rect 2520 20682 2560 20714
rect 2592 20682 2632 20714
rect 2664 20682 2704 20714
rect 2736 20682 2776 20714
rect 2808 20682 2848 20714
rect 2880 20682 2920 20714
rect 2952 20682 2992 20714
rect 3024 20682 3064 20714
rect 3096 20682 3136 20714
rect 3168 20682 3208 20714
rect 3240 20682 3280 20714
rect 3312 20682 3352 20714
rect 3384 20682 3424 20714
rect 3456 20682 3496 20714
rect 3528 20682 3568 20714
rect 3600 20682 3640 20714
rect 3672 20682 3712 20714
rect 3744 20682 3784 20714
rect 3816 20682 3856 20714
rect 3888 20682 4000 20714
rect 0 20642 4000 20682
rect 0 20610 112 20642
rect 144 20610 184 20642
rect 216 20610 256 20642
rect 288 20610 328 20642
rect 360 20610 400 20642
rect 432 20610 472 20642
rect 504 20610 544 20642
rect 576 20610 616 20642
rect 648 20610 688 20642
rect 720 20610 760 20642
rect 792 20610 832 20642
rect 864 20610 904 20642
rect 936 20610 976 20642
rect 1008 20610 1048 20642
rect 1080 20610 1120 20642
rect 1152 20610 1192 20642
rect 1224 20610 1264 20642
rect 1296 20610 1336 20642
rect 1368 20610 1408 20642
rect 1440 20610 1480 20642
rect 1512 20610 1552 20642
rect 1584 20610 1624 20642
rect 1656 20610 1696 20642
rect 1728 20610 1768 20642
rect 1800 20610 1840 20642
rect 1872 20610 1912 20642
rect 1944 20610 1984 20642
rect 2016 20610 2056 20642
rect 2088 20610 2128 20642
rect 2160 20610 2200 20642
rect 2232 20610 2272 20642
rect 2304 20610 2344 20642
rect 2376 20610 2416 20642
rect 2448 20610 2488 20642
rect 2520 20610 2560 20642
rect 2592 20610 2632 20642
rect 2664 20610 2704 20642
rect 2736 20610 2776 20642
rect 2808 20610 2848 20642
rect 2880 20610 2920 20642
rect 2952 20610 2992 20642
rect 3024 20610 3064 20642
rect 3096 20610 3136 20642
rect 3168 20610 3208 20642
rect 3240 20610 3280 20642
rect 3312 20610 3352 20642
rect 3384 20610 3424 20642
rect 3456 20610 3496 20642
rect 3528 20610 3568 20642
rect 3600 20610 3640 20642
rect 3672 20610 3712 20642
rect 3744 20610 3784 20642
rect 3816 20610 3856 20642
rect 3888 20610 4000 20642
rect 0 20570 4000 20610
rect 0 20538 112 20570
rect 144 20538 184 20570
rect 216 20538 256 20570
rect 288 20538 328 20570
rect 360 20538 400 20570
rect 432 20538 472 20570
rect 504 20538 544 20570
rect 576 20538 616 20570
rect 648 20538 688 20570
rect 720 20538 760 20570
rect 792 20538 832 20570
rect 864 20538 904 20570
rect 936 20538 976 20570
rect 1008 20538 1048 20570
rect 1080 20538 1120 20570
rect 1152 20538 1192 20570
rect 1224 20538 1264 20570
rect 1296 20538 1336 20570
rect 1368 20538 1408 20570
rect 1440 20538 1480 20570
rect 1512 20538 1552 20570
rect 1584 20538 1624 20570
rect 1656 20538 1696 20570
rect 1728 20538 1768 20570
rect 1800 20538 1840 20570
rect 1872 20538 1912 20570
rect 1944 20538 1984 20570
rect 2016 20538 2056 20570
rect 2088 20538 2128 20570
rect 2160 20538 2200 20570
rect 2232 20538 2272 20570
rect 2304 20538 2344 20570
rect 2376 20538 2416 20570
rect 2448 20538 2488 20570
rect 2520 20538 2560 20570
rect 2592 20538 2632 20570
rect 2664 20538 2704 20570
rect 2736 20538 2776 20570
rect 2808 20538 2848 20570
rect 2880 20538 2920 20570
rect 2952 20538 2992 20570
rect 3024 20538 3064 20570
rect 3096 20538 3136 20570
rect 3168 20538 3208 20570
rect 3240 20538 3280 20570
rect 3312 20538 3352 20570
rect 3384 20538 3424 20570
rect 3456 20538 3496 20570
rect 3528 20538 3568 20570
rect 3600 20538 3640 20570
rect 3672 20538 3712 20570
rect 3744 20538 3784 20570
rect 3816 20538 3856 20570
rect 3888 20538 4000 20570
rect 0 20498 4000 20538
rect 0 20466 112 20498
rect 144 20466 184 20498
rect 216 20466 256 20498
rect 288 20466 328 20498
rect 360 20466 400 20498
rect 432 20466 472 20498
rect 504 20466 544 20498
rect 576 20466 616 20498
rect 648 20466 688 20498
rect 720 20466 760 20498
rect 792 20466 832 20498
rect 864 20466 904 20498
rect 936 20466 976 20498
rect 1008 20466 1048 20498
rect 1080 20466 1120 20498
rect 1152 20466 1192 20498
rect 1224 20466 1264 20498
rect 1296 20466 1336 20498
rect 1368 20466 1408 20498
rect 1440 20466 1480 20498
rect 1512 20466 1552 20498
rect 1584 20466 1624 20498
rect 1656 20466 1696 20498
rect 1728 20466 1768 20498
rect 1800 20466 1840 20498
rect 1872 20466 1912 20498
rect 1944 20466 1984 20498
rect 2016 20466 2056 20498
rect 2088 20466 2128 20498
rect 2160 20466 2200 20498
rect 2232 20466 2272 20498
rect 2304 20466 2344 20498
rect 2376 20466 2416 20498
rect 2448 20466 2488 20498
rect 2520 20466 2560 20498
rect 2592 20466 2632 20498
rect 2664 20466 2704 20498
rect 2736 20466 2776 20498
rect 2808 20466 2848 20498
rect 2880 20466 2920 20498
rect 2952 20466 2992 20498
rect 3024 20466 3064 20498
rect 3096 20466 3136 20498
rect 3168 20466 3208 20498
rect 3240 20466 3280 20498
rect 3312 20466 3352 20498
rect 3384 20466 3424 20498
rect 3456 20466 3496 20498
rect 3528 20466 3568 20498
rect 3600 20466 3640 20498
rect 3672 20466 3712 20498
rect 3744 20466 3784 20498
rect 3816 20466 3856 20498
rect 3888 20466 4000 20498
rect 0 20426 4000 20466
rect 0 20394 112 20426
rect 144 20394 184 20426
rect 216 20394 256 20426
rect 288 20394 328 20426
rect 360 20394 400 20426
rect 432 20394 472 20426
rect 504 20394 544 20426
rect 576 20394 616 20426
rect 648 20394 688 20426
rect 720 20394 760 20426
rect 792 20394 832 20426
rect 864 20394 904 20426
rect 936 20394 976 20426
rect 1008 20394 1048 20426
rect 1080 20394 1120 20426
rect 1152 20394 1192 20426
rect 1224 20394 1264 20426
rect 1296 20394 1336 20426
rect 1368 20394 1408 20426
rect 1440 20394 1480 20426
rect 1512 20394 1552 20426
rect 1584 20394 1624 20426
rect 1656 20394 1696 20426
rect 1728 20394 1768 20426
rect 1800 20394 1840 20426
rect 1872 20394 1912 20426
rect 1944 20394 1984 20426
rect 2016 20394 2056 20426
rect 2088 20394 2128 20426
rect 2160 20394 2200 20426
rect 2232 20394 2272 20426
rect 2304 20394 2344 20426
rect 2376 20394 2416 20426
rect 2448 20394 2488 20426
rect 2520 20394 2560 20426
rect 2592 20394 2632 20426
rect 2664 20394 2704 20426
rect 2736 20394 2776 20426
rect 2808 20394 2848 20426
rect 2880 20394 2920 20426
rect 2952 20394 2992 20426
rect 3024 20394 3064 20426
rect 3096 20394 3136 20426
rect 3168 20394 3208 20426
rect 3240 20394 3280 20426
rect 3312 20394 3352 20426
rect 3384 20394 3424 20426
rect 3456 20394 3496 20426
rect 3528 20394 3568 20426
rect 3600 20394 3640 20426
rect 3672 20394 3712 20426
rect 3744 20394 3784 20426
rect 3816 20394 3856 20426
rect 3888 20394 4000 20426
rect 0 20354 4000 20394
rect 0 20322 112 20354
rect 144 20322 184 20354
rect 216 20322 256 20354
rect 288 20322 328 20354
rect 360 20322 400 20354
rect 432 20322 472 20354
rect 504 20322 544 20354
rect 576 20322 616 20354
rect 648 20322 688 20354
rect 720 20322 760 20354
rect 792 20322 832 20354
rect 864 20322 904 20354
rect 936 20322 976 20354
rect 1008 20322 1048 20354
rect 1080 20322 1120 20354
rect 1152 20322 1192 20354
rect 1224 20322 1264 20354
rect 1296 20322 1336 20354
rect 1368 20322 1408 20354
rect 1440 20322 1480 20354
rect 1512 20322 1552 20354
rect 1584 20322 1624 20354
rect 1656 20322 1696 20354
rect 1728 20322 1768 20354
rect 1800 20322 1840 20354
rect 1872 20322 1912 20354
rect 1944 20322 1984 20354
rect 2016 20322 2056 20354
rect 2088 20322 2128 20354
rect 2160 20322 2200 20354
rect 2232 20322 2272 20354
rect 2304 20322 2344 20354
rect 2376 20322 2416 20354
rect 2448 20322 2488 20354
rect 2520 20322 2560 20354
rect 2592 20322 2632 20354
rect 2664 20322 2704 20354
rect 2736 20322 2776 20354
rect 2808 20322 2848 20354
rect 2880 20322 2920 20354
rect 2952 20322 2992 20354
rect 3024 20322 3064 20354
rect 3096 20322 3136 20354
rect 3168 20322 3208 20354
rect 3240 20322 3280 20354
rect 3312 20322 3352 20354
rect 3384 20322 3424 20354
rect 3456 20322 3496 20354
rect 3528 20322 3568 20354
rect 3600 20322 3640 20354
rect 3672 20322 3712 20354
rect 3744 20322 3784 20354
rect 3816 20322 3856 20354
rect 3888 20322 4000 20354
rect 0 20282 4000 20322
rect 0 20250 112 20282
rect 144 20250 184 20282
rect 216 20250 256 20282
rect 288 20250 328 20282
rect 360 20250 400 20282
rect 432 20250 472 20282
rect 504 20250 544 20282
rect 576 20250 616 20282
rect 648 20250 688 20282
rect 720 20250 760 20282
rect 792 20250 832 20282
rect 864 20250 904 20282
rect 936 20250 976 20282
rect 1008 20250 1048 20282
rect 1080 20250 1120 20282
rect 1152 20250 1192 20282
rect 1224 20250 1264 20282
rect 1296 20250 1336 20282
rect 1368 20250 1408 20282
rect 1440 20250 1480 20282
rect 1512 20250 1552 20282
rect 1584 20250 1624 20282
rect 1656 20250 1696 20282
rect 1728 20250 1768 20282
rect 1800 20250 1840 20282
rect 1872 20250 1912 20282
rect 1944 20250 1984 20282
rect 2016 20250 2056 20282
rect 2088 20250 2128 20282
rect 2160 20250 2200 20282
rect 2232 20250 2272 20282
rect 2304 20250 2344 20282
rect 2376 20250 2416 20282
rect 2448 20250 2488 20282
rect 2520 20250 2560 20282
rect 2592 20250 2632 20282
rect 2664 20250 2704 20282
rect 2736 20250 2776 20282
rect 2808 20250 2848 20282
rect 2880 20250 2920 20282
rect 2952 20250 2992 20282
rect 3024 20250 3064 20282
rect 3096 20250 3136 20282
rect 3168 20250 3208 20282
rect 3240 20250 3280 20282
rect 3312 20250 3352 20282
rect 3384 20250 3424 20282
rect 3456 20250 3496 20282
rect 3528 20250 3568 20282
rect 3600 20250 3640 20282
rect 3672 20250 3712 20282
rect 3744 20250 3784 20282
rect 3816 20250 3856 20282
rect 3888 20250 4000 20282
rect 0 20210 4000 20250
rect 0 20178 112 20210
rect 144 20178 184 20210
rect 216 20178 256 20210
rect 288 20178 328 20210
rect 360 20178 400 20210
rect 432 20178 472 20210
rect 504 20178 544 20210
rect 576 20178 616 20210
rect 648 20178 688 20210
rect 720 20178 760 20210
rect 792 20178 832 20210
rect 864 20178 904 20210
rect 936 20178 976 20210
rect 1008 20178 1048 20210
rect 1080 20178 1120 20210
rect 1152 20178 1192 20210
rect 1224 20178 1264 20210
rect 1296 20178 1336 20210
rect 1368 20178 1408 20210
rect 1440 20178 1480 20210
rect 1512 20178 1552 20210
rect 1584 20178 1624 20210
rect 1656 20178 1696 20210
rect 1728 20178 1768 20210
rect 1800 20178 1840 20210
rect 1872 20178 1912 20210
rect 1944 20178 1984 20210
rect 2016 20178 2056 20210
rect 2088 20178 2128 20210
rect 2160 20178 2200 20210
rect 2232 20178 2272 20210
rect 2304 20178 2344 20210
rect 2376 20178 2416 20210
rect 2448 20178 2488 20210
rect 2520 20178 2560 20210
rect 2592 20178 2632 20210
rect 2664 20178 2704 20210
rect 2736 20178 2776 20210
rect 2808 20178 2848 20210
rect 2880 20178 2920 20210
rect 2952 20178 2992 20210
rect 3024 20178 3064 20210
rect 3096 20178 3136 20210
rect 3168 20178 3208 20210
rect 3240 20178 3280 20210
rect 3312 20178 3352 20210
rect 3384 20178 3424 20210
rect 3456 20178 3496 20210
rect 3528 20178 3568 20210
rect 3600 20178 3640 20210
rect 3672 20178 3712 20210
rect 3744 20178 3784 20210
rect 3816 20178 3856 20210
rect 3888 20178 4000 20210
rect 0 20138 4000 20178
rect 0 20106 112 20138
rect 144 20106 184 20138
rect 216 20106 256 20138
rect 288 20106 328 20138
rect 360 20106 400 20138
rect 432 20106 472 20138
rect 504 20106 544 20138
rect 576 20106 616 20138
rect 648 20106 688 20138
rect 720 20106 760 20138
rect 792 20106 832 20138
rect 864 20106 904 20138
rect 936 20106 976 20138
rect 1008 20106 1048 20138
rect 1080 20106 1120 20138
rect 1152 20106 1192 20138
rect 1224 20106 1264 20138
rect 1296 20106 1336 20138
rect 1368 20106 1408 20138
rect 1440 20106 1480 20138
rect 1512 20106 1552 20138
rect 1584 20106 1624 20138
rect 1656 20106 1696 20138
rect 1728 20106 1768 20138
rect 1800 20106 1840 20138
rect 1872 20106 1912 20138
rect 1944 20106 1984 20138
rect 2016 20106 2056 20138
rect 2088 20106 2128 20138
rect 2160 20106 2200 20138
rect 2232 20106 2272 20138
rect 2304 20106 2344 20138
rect 2376 20106 2416 20138
rect 2448 20106 2488 20138
rect 2520 20106 2560 20138
rect 2592 20106 2632 20138
rect 2664 20106 2704 20138
rect 2736 20106 2776 20138
rect 2808 20106 2848 20138
rect 2880 20106 2920 20138
rect 2952 20106 2992 20138
rect 3024 20106 3064 20138
rect 3096 20106 3136 20138
rect 3168 20106 3208 20138
rect 3240 20106 3280 20138
rect 3312 20106 3352 20138
rect 3384 20106 3424 20138
rect 3456 20106 3496 20138
rect 3528 20106 3568 20138
rect 3600 20106 3640 20138
rect 3672 20106 3712 20138
rect 3744 20106 3784 20138
rect 3816 20106 3856 20138
rect 3888 20106 4000 20138
rect 0 20066 4000 20106
rect 0 20034 112 20066
rect 144 20034 184 20066
rect 216 20034 256 20066
rect 288 20034 328 20066
rect 360 20034 400 20066
rect 432 20034 472 20066
rect 504 20034 544 20066
rect 576 20034 616 20066
rect 648 20034 688 20066
rect 720 20034 760 20066
rect 792 20034 832 20066
rect 864 20034 904 20066
rect 936 20034 976 20066
rect 1008 20034 1048 20066
rect 1080 20034 1120 20066
rect 1152 20034 1192 20066
rect 1224 20034 1264 20066
rect 1296 20034 1336 20066
rect 1368 20034 1408 20066
rect 1440 20034 1480 20066
rect 1512 20034 1552 20066
rect 1584 20034 1624 20066
rect 1656 20034 1696 20066
rect 1728 20034 1768 20066
rect 1800 20034 1840 20066
rect 1872 20034 1912 20066
rect 1944 20034 1984 20066
rect 2016 20034 2056 20066
rect 2088 20034 2128 20066
rect 2160 20034 2200 20066
rect 2232 20034 2272 20066
rect 2304 20034 2344 20066
rect 2376 20034 2416 20066
rect 2448 20034 2488 20066
rect 2520 20034 2560 20066
rect 2592 20034 2632 20066
rect 2664 20034 2704 20066
rect 2736 20034 2776 20066
rect 2808 20034 2848 20066
rect 2880 20034 2920 20066
rect 2952 20034 2992 20066
rect 3024 20034 3064 20066
rect 3096 20034 3136 20066
rect 3168 20034 3208 20066
rect 3240 20034 3280 20066
rect 3312 20034 3352 20066
rect 3384 20034 3424 20066
rect 3456 20034 3496 20066
rect 3528 20034 3568 20066
rect 3600 20034 3640 20066
rect 3672 20034 3712 20066
rect 3744 20034 3784 20066
rect 3816 20034 3856 20066
rect 3888 20034 4000 20066
rect 0 19994 4000 20034
rect 0 19962 112 19994
rect 144 19962 184 19994
rect 216 19962 256 19994
rect 288 19962 328 19994
rect 360 19962 400 19994
rect 432 19962 472 19994
rect 504 19962 544 19994
rect 576 19962 616 19994
rect 648 19962 688 19994
rect 720 19962 760 19994
rect 792 19962 832 19994
rect 864 19962 904 19994
rect 936 19962 976 19994
rect 1008 19962 1048 19994
rect 1080 19962 1120 19994
rect 1152 19962 1192 19994
rect 1224 19962 1264 19994
rect 1296 19962 1336 19994
rect 1368 19962 1408 19994
rect 1440 19962 1480 19994
rect 1512 19962 1552 19994
rect 1584 19962 1624 19994
rect 1656 19962 1696 19994
rect 1728 19962 1768 19994
rect 1800 19962 1840 19994
rect 1872 19962 1912 19994
rect 1944 19962 1984 19994
rect 2016 19962 2056 19994
rect 2088 19962 2128 19994
rect 2160 19962 2200 19994
rect 2232 19962 2272 19994
rect 2304 19962 2344 19994
rect 2376 19962 2416 19994
rect 2448 19962 2488 19994
rect 2520 19962 2560 19994
rect 2592 19962 2632 19994
rect 2664 19962 2704 19994
rect 2736 19962 2776 19994
rect 2808 19962 2848 19994
rect 2880 19962 2920 19994
rect 2952 19962 2992 19994
rect 3024 19962 3064 19994
rect 3096 19962 3136 19994
rect 3168 19962 3208 19994
rect 3240 19962 3280 19994
rect 3312 19962 3352 19994
rect 3384 19962 3424 19994
rect 3456 19962 3496 19994
rect 3528 19962 3568 19994
rect 3600 19962 3640 19994
rect 3672 19962 3712 19994
rect 3744 19962 3784 19994
rect 3816 19962 3856 19994
rect 3888 19962 4000 19994
rect 0 19922 4000 19962
rect 0 19890 112 19922
rect 144 19890 184 19922
rect 216 19890 256 19922
rect 288 19890 328 19922
rect 360 19890 400 19922
rect 432 19890 472 19922
rect 504 19890 544 19922
rect 576 19890 616 19922
rect 648 19890 688 19922
rect 720 19890 760 19922
rect 792 19890 832 19922
rect 864 19890 904 19922
rect 936 19890 976 19922
rect 1008 19890 1048 19922
rect 1080 19890 1120 19922
rect 1152 19890 1192 19922
rect 1224 19890 1264 19922
rect 1296 19890 1336 19922
rect 1368 19890 1408 19922
rect 1440 19890 1480 19922
rect 1512 19890 1552 19922
rect 1584 19890 1624 19922
rect 1656 19890 1696 19922
rect 1728 19890 1768 19922
rect 1800 19890 1840 19922
rect 1872 19890 1912 19922
rect 1944 19890 1984 19922
rect 2016 19890 2056 19922
rect 2088 19890 2128 19922
rect 2160 19890 2200 19922
rect 2232 19890 2272 19922
rect 2304 19890 2344 19922
rect 2376 19890 2416 19922
rect 2448 19890 2488 19922
rect 2520 19890 2560 19922
rect 2592 19890 2632 19922
rect 2664 19890 2704 19922
rect 2736 19890 2776 19922
rect 2808 19890 2848 19922
rect 2880 19890 2920 19922
rect 2952 19890 2992 19922
rect 3024 19890 3064 19922
rect 3096 19890 3136 19922
rect 3168 19890 3208 19922
rect 3240 19890 3280 19922
rect 3312 19890 3352 19922
rect 3384 19890 3424 19922
rect 3456 19890 3496 19922
rect 3528 19890 3568 19922
rect 3600 19890 3640 19922
rect 3672 19890 3712 19922
rect 3744 19890 3784 19922
rect 3816 19890 3856 19922
rect 3888 19890 4000 19922
rect 0 19850 4000 19890
rect 0 19818 112 19850
rect 144 19818 184 19850
rect 216 19818 256 19850
rect 288 19818 328 19850
rect 360 19818 400 19850
rect 432 19818 472 19850
rect 504 19818 544 19850
rect 576 19818 616 19850
rect 648 19818 688 19850
rect 720 19818 760 19850
rect 792 19818 832 19850
rect 864 19818 904 19850
rect 936 19818 976 19850
rect 1008 19818 1048 19850
rect 1080 19818 1120 19850
rect 1152 19818 1192 19850
rect 1224 19818 1264 19850
rect 1296 19818 1336 19850
rect 1368 19818 1408 19850
rect 1440 19818 1480 19850
rect 1512 19818 1552 19850
rect 1584 19818 1624 19850
rect 1656 19818 1696 19850
rect 1728 19818 1768 19850
rect 1800 19818 1840 19850
rect 1872 19818 1912 19850
rect 1944 19818 1984 19850
rect 2016 19818 2056 19850
rect 2088 19818 2128 19850
rect 2160 19818 2200 19850
rect 2232 19818 2272 19850
rect 2304 19818 2344 19850
rect 2376 19818 2416 19850
rect 2448 19818 2488 19850
rect 2520 19818 2560 19850
rect 2592 19818 2632 19850
rect 2664 19818 2704 19850
rect 2736 19818 2776 19850
rect 2808 19818 2848 19850
rect 2880 19818 2920 19850
rect 2952 19818 2992 19850
rect 3024 19818 3064 19850
rect 3096 19818 3136 19850
rect 3168 19818 3208 19850
rect 3240 19818 3280 19850
rect 3312 19818 3352 19850
rect 3384 19818 3424 19850
rect 3456 19818 3496 19850
rect 3528 19818 3568 19850
rect 3600 19818 3640 19850
rect 3672 19818 3712 19850
rect 3744 19818 3784 19850
rect 3816 19818 3856 19850
rect 3888 19818 4000 19850
rect 0 19778 4000 19818
rect 0 19746 112 19778
rect 144 19746 184 19778
rect 216 19746 256 19778
rect 288 19746 328 19778
rect 360 19746 400 19778
rect 432 19746 472 19778
rect 504 19746 544 19778
rect 576 19746 616 19778
rect 648 19746 688 19778
rect 720 19746 760 19778
rect 792 19746 832 19778
rect 864 19746 904 19778
rect 936 19746 976 19778
rect 1008 19746 1048 19778
rect 1080 19746 1120 19778
rect 1152 19746 1192 19778
rect 1224 19746 1264 19778
rect 1296 19746 1336 19778
rect 1368 19746 1408 19778
rect 1440 19746 1480 19778
rect 1512 19746 1552 19778
rect 1584 19746 1624 19778
rect 1656 19746 1696 19778
rect 1728 19746 1768 19778
rect 1800 19746 1840 19778
rect 1872 19746 1912 19778
rect 1944 19746 1984 19778
rect 2016 19746 2056 19778
rect 2088 19746 2128 19778
rect 2160 19746 2200 19778
rect 2232 19746 2272 19778
rect 2304 19746 2344 19778
rect 2376 19746 2416 19778
rect 2448 19746 2488 19778
rect 2520 19746 2560 19778
rect 2592 19746 2632 19778
rect 2664 19746 2704 19778
rect 2736 19746 2776 19778
rect 2808 19746 2848 19778
rect 2880 19746 2920 19778
rect 2952 19746 2992 19778
rect 3024 19746 3064 19778
rect 3096 19746 3136 19778
rect 3168 19746 3208 19778
rect 3240 19746 3280 19778
rect 3312 19746 3352 19778
rect 3384 19746 3424 19778
rect 3456 19746 3496 19778
rect 3528 19746 3568 19778
rect 3600 19746 3640 19778
rect 3672 19746 3712 19778
rect 3744 19746 3784 19778
rect 3816 19746 3856 19778
rect 3888 19746 4000 19778
rect 0 19706 4000 19746
rect 0 19674 112 19706
rect 144 19674 184 19706
rect 216 19674 256 19706
rect 288 19674 328 19706
rect 360 19674 400 19706
rect 432 19674 472 19706
rect 504 19674 544 19706
rect 576 19674 616 19706
rect 648 19674 688 19706
rect 720 19674 760 19706
rect 792 19674 832 19706
rect 864 19674 904 19706
rect 936 19674 976 19706
rect 1008 19674 1048 19706
rect 1080 19674 1120 19706
rect 1152 19674 1192 19706
rect 1224 19674 1264 19706
rect 1296 19674 1336 19706
rect 1368 19674 1408 19706
rect 1440 19674 1480 19706
rect 1512 19674 1552 19706
rect 1584 19674 1624 19706
rect 1656 19674 1696 19706
rect 1728 19674 1768 19706
rect 1800 19674 1840 19706
rect 1872 19674 1912 19706
rect 1944 19674 1984 19706
rect 2016 19674 2056 19706
rect 2088 19674 2128 19706
rect 2160 19674 2200 19706
rect 2232 19674 2272 19706
rect 2304 19674 2344 19706
rect 2376 19674 2416 19706
rect 2448 19674 2488 19706
rect 2520 19674 2560 19706
rect 2592 19674 2632 19706
rect 2664 19674 2704 19706
rect 2736 19674 2776 19706
rect 2808 19674 2848 19706
rect 2880 19674 2920 19706
rect 2952 19674 2992 19706
rect 3024 19674 3064 19706
rect 3096 19674 3136 19706
rect 3168 19674 3208 19706
rect 3240 19674 3280 19706
rect 3312 19674 3352 19706
rect 3384 19674 3424 19706
rect 3456 19674 3496 19706
rect 3528 19674 3568 19706
rect 3600 19674 3640 19706
rect 3672 19674 3712 19706
rect 3744 19674 3784 19706
rect 3816 19674 3856 19706
rect 3888 19674 4000 19706
rect 0 19634 4000 19674
rect 0 19602 112 19634
rect 144 19602 184 19634
rect 216 19602 256 19634
rect 288 19602 328 19634
rect 360 19602 400 19634
rect 432 19602 472 19634
rect 504 19602 544 19634
rect 576 19602 616 19634
rect 648 19602 688 19634
rect 720 19602 760 19634
rect 792 19602 832 19634
rect 864 19602 904 19634
rect 936 19602 976 19634
rect 1008 19602 1048 19634
rect 1080 19602 1120 19634
rect 1152 19602 1192 19634
rect 1224 19602 1264 19634
rect 1296 19602 1336 19634
rect 1368 19602 1408 19634
rect 1440 19602 1480 19634
rect 1512 19602 1552 19634
rect 1584 19602 1624 19634
rect 1656 19602 1696 19634
rect 1728 19602 1768 19634
rect 1800 19602 1840 19634
rect 1872 19602 1912 19634
rect 1944 19602 1984 19634
rect 2016 19602 2056 19634
rect 2088 19602 2128 19634
rect 2160 19602 2200 19634
rect 2232 19602 2272 19634
rect 2304 19602 2344 19634
rect 2376 19602 2416 19634
rect 2448 19602 2488 19634
rect 2520 19602 2560 19634
rect 2592 19602 2632 19634
rect 2664 19602 2704 19634
rect 2736 19602 2776 19634
rect 2808 19602 2848 19634
rect 2880 19602 2920 19634
rect 2952 19602 2992 19634
rect 3024 19602 3064 19634
rect 3096 19602 3136 19634
rect 3168 19602 3208 19634
rect 3240 19602 3280 19634
rect 3312 19602 3352 19634
rect 3384 19602 3424 19634
rect 3456 19602 3496 19634
rect 3528 19602 3568 19634
rect 3600 19602 3640 19634
rect 3672 19602 3712 19634
rect 3744 19602 3784 19634
rect 3816 19602 3856 19634
rect 3888 19602 4000 19634
rect 0 19562 4000 19602
rect 0 19530 112 19562
rect 144 19530 184 19562
rect 216 19530 256 19562
rect 288 19530 328 19562
rect 360 19530 400 19562
rect 432 19530 472 19562
rect 504 19530 544 19562
rect 576 19530 616 19562
rect 648 19530 688 19562
rect 720 19530 760 19562
rect 792 19530 832 19562
rect 864 19530 904 19562
rect 936 19530 976 19562
rect 1008 19530 1048 19562
rect 1080 19530 1120 19562
rect 1152 19530 1192 19562
rect 1224 19530 1264 19562
rect 1296 19530 1336 19562
rect 1368 19530 1408 19562
rect 1440 19530 1480 19562
rect 1512 19530 1552 19562
rect 1584 19530 1624 19562
rect 1656 19530 1696 19562
rect 1728 19530 1768 19562
rect 1800 19530 1840 19562
rect 1872 19530 1912 19562
rect 1944 19530 1984 19562
rect 2016 19530 2056 19562
rect 2088 19530 2128 19562
rect 2160 19530 2200 19562
rect 2232 19530 2272 19562
rect 2304 19530 2344 19562
rect 2376 19530 2416 19562
rect 2448 19530 2488 19562
rect 2520 19530 2560 19562
rect 2592 19530 2632 19562
rect 2664 19530 2704 19562
rect 2736 19530 2776 19562
rect 2808 19530 2848 19562
rect 2880 19530 2920 19562
rect 2952 19530 2992 19562
rect 3024 19530 3064 19562
rect 3096 19530 3136 19562
rect 3168 19530 3208 19562
rect 3240 19530 3280 19562
rect 3312 19530 3352 19562
rect 3384 19530 3424 19562
rect 3456 19530 3496 19562
rect 3528 19530 3568 19562
rect 3600 19530 3640 19562
rect 3672 19530 3712 19562
rect 3744 19530 3784 19562
rect 3816 19530 3856 19562
rect 3888 19530 4000 19562
rect 0 19490 4000 19530
rect 0 19458 112 19490
rect 144 19458 184 19490
rect 216 19458 256 19490
rect 288 19458 328 19490
rect 360 19458 400 19490
rect 432 19458 472 19490
rect 504 19458 544 19490
rect 576 19458 616 19490
rect 648 19458 688 19490
rect 720 19458 760 19490
rect 792 19458 832 19490
rect 864 19458 904 19490
rect 936 19458 976 19490
rect 1008 19458 1048 19490
rect 1080 19458 1120 19490
rect 1152 19458 1192 19490
rect 1224 19458 1264 19490
rect 1296 19458 1336 19490
rect 1368 19458 1408 19490
rect 1440 19458 1480 19490
rect 1512 19458 1552 19490
rect 1584 19458 1624 19490
rect 1656 19458 1696 19490
rect 1728 19458 1768 19490
rect 1800 19458 1840 19490
rect 1872 19458 1912 19490
rect 1944 19458 1984 19490
rect 2016 19458 2056 19490
rect 2088 19458 2128 19490
rect 2160 19458 2200 19490
rect 2232 19458 2272 19490
rect 2304 19458 2344 19490
rect 2376 19458 2416 19490
rect 2448 19458 2488 19490
rect 2520 19458 2560 19490
rect 2592 19458 2632 19490
rect 2664 19458 2704 19490
rect 2736 19458 2776 19490
rect 2808 19458 2848 19490
rect 2880 19458 2920 19490
rect 2952 19458 2992 19490
rect 3024 19458 3064 19490
rect 3096 19458 3136 19490
rect 3168 19458 3208 19490
rect 3240 19458 3280 19490
rect 3312 19458 3352 19490
rect 3384 19458 3424 19490
rect 3456 19458 3496 19490
rect 3528 19458 3568 19490
rect 3600 19458 3640 19490
rect 3672 19458 3712 19490
rect 3744 19458 3784 19490
rect 3816 19458 3856 19490
rect 3888 19458 4000 19490
rect 0 19418 4000 19458
rect 0 19386 112 19418
rect 144 19386 184 19418
rect 216 19386 256 19418
rect 288 19386 328 19418
rect 360 19386 400 19418
rect 432 19386 472 19418
rect 504 19386 544 19418
rect 576 19386 616 19418
rect 648 19386 688 19418
rect 720 19386 760 19418
rect 792 19386 832 19418
rect 864 19386 904 19418
rect 936 19386 976 19418
rect 1008 19386 1048 19418
rect 1080 19386 1120 19418
rect 1152 19386 1192 19418
rect 1224 19386 1264 19418
rect 1296 19386 1336 19418
rect 1368 19386 1408 19418
rect 1440 19386 1480 19418
rect 1512 19386 1552 19418
rect 1584 19386 1624 19418
rect 1656 19386 1696 19418
rect 1728 19386 1768 19418
rect 1800 19386 1840 19418
rect 1872 19386 1912 19418
rect 1944 19386 1984 19418
rect 2016 19386 2056 19418
rect 2088 19386 2128 19418
rect 2160 19386 2200 19418
rect 2232 19386 2272 19418
rect 2304 19386 2344 19418
rect 2376 19386 2416 19418
rect 2448 19386 2488 19418
rect 2520 19386 2560 19418
rect 2592 19386 2632 19418
rect 2664 19386 2704 19418
rect 2736 19386 2776 19418
rect 2808 19386 2848 19418
rect 2880 19386 2920 19418
rect 2952 19386 2992 19418
rect 3024 19386 3064 19418
rect 3096 19386 3136 19418
rect 3168 19386 3208 19418
rect 3240 19386 3280 19418
rect 3312 19386 3352 19418
rect 3384 19386 3424 19418
rect 3456 19386 3496 19418
rect 3528 19386 3568 19418
rect 3600 19386 3640 19418
rect 3672 19386 3712 19418
rect 3744 19386 3784 19418
rect 3816 19386 3856 19418
rect 3888 19386 4000 19418
rect 0 19346 4000 19386
rect 0 19314 112 19346
rect 144 19314 184 19346
rect 216 19314 256 19346
rect 288 19314 328 19346
rect 360 19314 400 19346
rect 432 19314 472 19346
rect 504 19314 544 19346
rect 576 19314 616 19346
rect 648 19314 688 19346
rect 720 19314 760 19346
rect 792 19314 832 19346
rect 864 19314 904 19346
rect 936 19314 976 19346
rect 1008 19314 1048 19346
rect 1080 19314 1120 19346
rect 1152 19314 1192 19346
rect 1224 19314 1264 19346
rect 1296 19314 1336 19346
rect 1368 19314 1408 19346
rect 1440 19314 1480 19346
rect 1512 19314 1552 19346
rect 1584 19314 1624 19346
rect 1656 19314 1696 19346
rect 1728 19314 1768 19346
rect 1800 19314 1840 19346
rect 1872 19314 1912 19346
rect 1944 19314 1984 19346
rect 2016 19314 2056 19346
rect 2088 19314 2128 19346
rect 2160 19314 2200 19346
rect 2232 19314 2272 19346
rect 2304 19314 2344 19346
rect 2376 19314 2416 19346
rect 2448 19314 2488 19346
rect 2520 19314 2560 19346
rect 2592 19314 2632 19346
rect 2664 19314 2704 19346
rect 2736 19314 2776 19346
rect 2808 19314 2848 19346
rect 2880 19314 2920 19346
rect 2952 19314 2992 19346
rect 3024 19314 3064 19346
rect 3096 19314 3136 19346
rect 3168 19314 3208 19346
rect 3240 19314 3280 19346
rect 3312 19314 3352 19346
rect 3384 19314 3424 19346
rect 3456 19314 3496 19346
rect 3528 19314 3568 19346
rect 3600 19314 3640 19346
rect 3672 19314 3712 19346
rect 3744 19314 3784 19346
rect 3816 19314 3856 19346
rect 3888 19314 4000 19346
rect 0 19274 4000 19314
rect 0 19242 112 19274
rect 144 19242 184 19274
rect 216 19242 256 19274
rect 288 19242 328 19274
rect 360 19242 400 19274
rect 432 19242 472 19274
rect 504 19242 544 19274
rect 576 19242 616 19274
rect 648 19242 688 19274
rect 720 19242 760 19274
rect 792 19242 832 19274
rect 864 19242 904 19274
rect 936 19242 976 19274
rect 1008 19242 1048 19274
rect 1080 19242 1120 19274
rect 1152 19242 1192 19274
rect 1224 19242 1264 19274
rect 1296 19242 1336 19274
rect 1368 19242 1408 19274
rect 1440 19242 1480 19274
rect 1512 19242 1552 19274
rect 1584 19242 1624 19274
rect 1656 19242 1696 19274
rect 1728 19242 1768 19274
rect 1800 19242 1840 19274
rect 1872 19242 1912 19274
rect 1944 19242 1984 19274
rect 2016 19242 2056 19274
rect 2088 19242 2128 19274
rect 2160 19242 2200 19274
rect 2232 19242 2272 19274
rect 2304 19242 2344 19274
rect 2376 19242 2416 19274
rect 2448 19242 2488 19274
rect 2520 19242 2560 19274
rect 2592 19242 2632 19274
rect 2664 19242 2704 19274
rect 2736 19242 2776 19274
rect 2808 19242 2848 19274
rect 2880 19242 2920 19274
rect 2952 19242 2992 19274
rect 3024 19242 3064 19274
rect 3096 19242 3136 19274
rect 3168 19242 3208 19274
rect 3240 19242 3280 19274
rect 3312 19242 3352 19274
rect 3384 19242 3424 19274
rect 3456 19242 3496 19274
rect 3528 19242 3568 19274
rect 3600 19242 3640 19274
rect 3672 19242 3712 19274
rect 3744 19242 3784 19274
rect 3816 19242 3856 19274
rect 3888 19242 4000 19274
rect 0 19202 4000 19242
rect 0 19170 112 19202
rect 144 19170 184 19202
rect 216 19170 256 19202
rect 288 19170 328 19202
rect 360 19170 400 19202
rect 432 19170 472 19202
rect 504 19170 544 19202
rect 576 19170 616 19202
rect 648 19170 688 19202
rect 720 19170 760 19202
rect 792 19170 832 19202
rect 864 19170 904 19202
rect 936 19170 976 19202
rect 1008 19170 1048 19202
rect 1080 19170 1120 19202
rect 1152 19170 1192 19202
rect 1224 19170 1264 19202
rect 1296 19170 1336 19202
rect 1368 19170 1408 19202
rect 1440 19170 1480 19202
rect 1512 19170 1552 19202
rect 1584 19170 1624 19202
rect 1656 19170 1696 19202
rect 1728 19170 1768 19202
rect 1800 19170 1840 19202
rect 1872 19170 1912 19202
rect 1944 19170 1984 19202
rect 2016 19170 2056 19202
rect 2088 19170 2128 19202
rect 2160 19170 2200 19202
rect 2232 19170 2272 19202
rect 2304 19170 2344 19202
rect 2376 19170 2416 19202
rect 2448 19170 2488 19202
rect 2520 19170 2560 19202
rect 2592 19170 2632 19202
rect 2664 19170 2704 19202
rect 2736 19170 2776 19202
rect 2808 19170 2848 19202
rect 2880 19170 2920 19202
rect 2952 19170 2992 19202
rect 3024 19170 3064 19202
rect 3096 19170 3136 19202
rect 3168 19170 3208 19202
rect 3240 19170 3280 19202
rect 3312 19170 3352 19202
rect 3384 19170 3424 19202
rect 3456 19170 3496 19202
rect 3528 19170 3568 19202
rect 3600 19170 3640 19202
rect 3672 19170 3712 19202
rect 3744 19170 3784 19202
rect 3816 19170 3856 19202
rect 3888 19170 4000 19202
rect 0 19130 4000 19170
rect 0 19098 112 19130
rect 144 19098 184 19130
rect 216 19098 256 19130
rect 288 19098 328 19130
rect 360 19098 400 19130
rect 432 19098 472 19130
rect 504 19098 544 19130
rect 576 19098 616 19130
rect 648 19098 688 19130
rect 720 19098 760 19130
rect 792 19098 832 19130
rect 864 19098 904 19130
rect 936 19098 976 19130
rect 1008 19098 1048 19130
rect 1080 19098 1120 19130
rect 1152 19098 1192 19130
rect 1224 19098 1264 19130
rect 1296 19098 1336 19130
rect 1368 19098 1408 19130
rect 1440 19098 1480 19130
rect 1512 19098 1552 19130
rect 1584 19098 1624 19130
rect 1656 19098 1696 19130
rect 1728 19098 1768 19130
rect 1800 19098 1840 19130
rect 1872 19098 1912 19130
rect 1944 19098 1984 19130
rect 2016 19098 2056 19130
rect 2088 19098 2128 19130
rect 2160 19098 2200 19130
rect 2232 19098 2272 19130
rect 2304 19098 2344 19130
rect 2376 19098 2416 19130
rect 2448 19098 2488 19130
rect 2520 19098 2560 19130
rect 2592 19098 2632 19130
rect 2664 19098 2704 19130
rect 2736 19098 2776 19130
rect 2808 19098 2848 19130
rect 2880 19098 2920 19130
rect 2952 19098 2992 19130
rect 3024 19098 3064 19130
rect 3096 19098 3136 19130
rect 3168 19098 3208 19130
rect 3240 19098 3280 19130
rect 3312 19098 3352 19130
rect 3384 19098 3424 19130
rect 3456 19098 3496 19130
rect 3528 19098 3568 19130
rect 3600 19098 3640 19130
rect 3672 19098 3712 19130
rect 3744 19098 3784 19130
rect 3816 19098 3856 19130
rect 3888 19098 4000 19130
rect 0 19058 4000 19098
rect 0 19026 112 19058
rect 144 19026 184 19058
rect 216 19026 256 19058
rect 288 19026 328 19058
rect 360 19026 400 19058
rect 432 19026 472 19058
rect 504 19026 544 19058
rect 576 19026 616 19058
rect 648 19026 688 19058
rect 720 19026 760 19058
rect 792 19026 832 19058
rect 864 19026 904 19058
rect 936 19026 976 19058
rect 1008 19026 1048 19058
rect 1080 19026 1120 19058
rect 1152 19026 1192 19058
rect 1224 19026 1264 19058
rect 1296 19026 1336 19058
rect 1368 19026 1408 19058
rect 1440 19026 1480 19058
rect 1512 19026 1552 19058
rect 1584 19026 1624 19058
rect 1656 19026 1696 19058
rect 1728 19026 1768 19058
rect 1800 19026 1840 19058
rect 1872 19026 1912 19058
rect 1944 19026 1984 19058
rect 2016 19026 2056 19058
rect 2088 19026 2128 19058
rect 2160 19026 2200 19058
rect 2232 19026 2272 19058
rect 2304 19026 2344 19058
rect 2376 19026 2416 19058
rect 2448 19026 2488 19058
rect 2520 19026 2560 19058
rect 2592 19026 2632 19058
rect 2664 19026 2704 19058
rect 2736 19026 2776 19058
rect 2808 19026 2848 19058
rect 2880 19026 2920 19058
rect 2952 19026 2992 19058
rect 3024 19026 3064 19058
rect 3096 19026 3136 19058
rect 3168 19026 3208 19058
rect 3240 19026 3280 19058
rect 3312 19026 3352 19058
rect 3384 19026 3424 19058
rect 3456 19026 3496 19058
rect 3528 19026 3568 19058
rect 3600 19026 3640 19058
rect 3672 19026 3712 19058
rect 3744 19026 3784 19058
rect 3816 19026 3856 19058
rect 3888 19026 4000 19058
rect 0 18986 4000 19026
rect 0 18954 112 18986
rect 144 18954 184 18986
rect 216 18954 256 18986
rect 288 18954 328 18986
rect 360 18954 400 18986
rect 432 18954 472 18986
rect 504 18954 544 18986
rect 576 18954 616 18986
rect 648 18954 688 18986
rect 720 18954 760 18986
rect 792 18954 832 18986
rect 864 18954 904 18986
rect 936 18954 976 18986
rect 1008 18954 1048 18986
rect 1080 18954 1120 18986
rect 1152 18954 1192 18986
rect 1224 18954 1264 18986
rect 1296 18954 1336 18986
rect 1368 18954 1408 18986
rect 1440 18954 1480 18986
rect 1512 18954 1552 18986
rect 1584 18954 1624 18986
rect 1656 18954 1696 18986
rect 1728 18954 1768 18986
rect 1800 18954 1840 18986
rect 1872 18954 1912 18986
rect 1944 18954 1984 18986
rect 2016 18954 2056 18986
rect 2088 18954 2128 18986
rect 2160 18954 2200 18986
rect 2232 18954 2272 18986
rect 2304 18954 2344 18986
rect 2376 18954 2416 18986
rect 2448 18954 2488 18986
rect 2520 18954 2560 18986
rect 2592 18954 2632 18986
rect 2664 18954 2704 18986
rect 2736 18954 2776 18986
rect 2808 18954 2848 18986
rect 2880 18954 2920 18986
rect 2952 18954 2992 18986
rect 3024 18954 3064 18986
rect 3096 18954 3136 18986
rect 3168 18954 3208 18986
rect 3240 18954 3280 18986
rect 3312 18954 3352 18986
rect 3384 18954 3424 18986
rect 3456 18954 3496 18986
rect 3528 18954 3568 18986
rect 3600 18954 3640 18986
rect 3672 18954 3712 18986
rect 3744 18954 3784 18986
rect 3816 18954 3856 18986
rect 3888 18954 4000 18986
rect 0 18914 4000 18954
rect 0 18882 112 18914
rect 144 18882 184 18914
rect 216 18882 256 18914
rect 288 18882 328 18914
rect 360 18882 400 18914
rect 432 18882 472 18914
rect 504 18882 544 18914
rect 576 18882 616 18914
rect 648 18882 688 18914
rect 720 18882 760 18914
rect 792 18882 832 18914
rect 864 18882 904 18914
rect 936 18882 976 18914
rect 1008 18882 1048 18914
rect 1080 18882 1120 18914
rect 1152 18882 1192 18914
rect 1224 18882 1264 18914
rect 1296 18882 1336 18914
rect 1368 18882 1408 18914
rect 1440 18882 1480 18914
rect 1512 18882 1552 18914
rect 1584 18882 1624 18914
rect 1656 18882 1696 18914
rect 1728 18882 1768 18914
rect 1800 18882 1840 18914
rect 1872 18882 1912 18914
rect 1944 18882 1984 18914
rect 2016 18882 2056 18914
rect 2088 18882 2128 18914
rect 2160 18882 2200 18914
rect 2232 18882 2272 18914
rect 2304 18882 2344 18914
rect 2376 18882 2416 18914
rect 2448 18882 2488 18914
rect 2520 18882 2560 18914
rect 2592 18882 2632 18914
rect 2664 18882 2704 18914
rect 2736 18882 2776 18914
rect 2808 18882 2848 18914
rect 2880 18882 2920 18914
rect 2952 18882 2992 18914
rect 3024 18882 3064 18914
rect 3096 18882 3136 18914
rect 3168 18882 3208 18914
rect 3240 18882 3280 18914
rect 3312 18882 3352 18914
rect 3384 18882 3424 18914
rect 3456 18882 3496 18914
rect 3528 18882 3568 18914
rect 3600 18882 3640 18914
rect 3672 18882 3712 18914
rect 3744 18882 3784 18914
rect 3816 18882 3856 18914
rect 3888 18882 4000 18914
rect 0 18842 4000 18882
rect 0 18810 112 18842
rect 144 18810 184 18842
rect 216 18810 256 18842
rect 288 18810 328 18842
rect 360 18810 400 18842
rect 432 18810 472 18842
rect 504 18810 544 18842
rect 576 18810 616 18842
rect 648 18810 688 18842
rect 720 18810 760 18842
rect 792 18810 832 18842
rect 864 18810 904 18842
rect 936 18810 976 18842
rect 1008 18810 1048 18842
rect 1080 18810 1120 18842
rect 1152 18810 1192 18842
rect 1224 18810 1264 18842
rect 1296 18810 1336 18842
rect 1368 18810 1408 18842
rect 1440 18810 1480 18842
rect 1512 18810 1552 18842
rect 1584 18810 1624 18842
rect 1656 18810 1696 18842
rect 1728 18810 1768 18842
rect 1800 18810 1840 18842
rect 1872 18810 1912 18842
rect 1944 18810 1984 18842
rect 2016 18810 2056 18842
rect 2088 18810 2128 18842
rect 2160 18810 2200 18842
rect 2232 18810 2272 18842
rect 2304 18810 2344 18842
rect 2376 18810 2416 18842
rect 2448 18810 2488 18842
rect 2520 18810 2560 18842
rect 2592 18810 2632 18842
rect 2664 18810 2704 18842
rect 2736 18810 2776 18842
rect 2808 18810 2848 18842
rect 2880 18810 2920 18842
rect 2952 18810 2992 18842
rect 3024 18810 3064 18842
rect 3096 18810 3136 18842
rect 3168 18810 3208 18842
rect 3240 18810 3280 18842
rect 3312 18810 3352 18842
rect 3384 18810 3424 18842
rect 3456 18810 3496 18842
rect 3528 18810 3568 18842
rect 3600 18810 3640 18842
rect 3672 18810 3712 18842
rect 3744 18810 3784 18842
rect 3816 18810 3856 18842
rect 3888 18810 4000 18842
rect 0 18770 4000 18810
rect 0 18738 112 18770
rect 144 18738 184 18770
rect 216 18738 256 18770
rect 288 18738 328 18770
rect 360 18738 400 18770
rect 432 18738 472 18770
rect 504 18738 544 18770
rect 576 18738 616 18770
rect 648 18738 688 18770
rect 720 18738 760 18770
rect 792 18738 832 18770
rect 864 18738 904 18770
rect 936 18738 976 18770
rect 1008 18738 1048 18770
rect 1080 18738 1120 18770
rect 1152 18738 1192 18770
rect 1224 18738 1264 18770
rect 1296 18738 1336 18770
rect 1368 18738 1408 18770
rect 1440 18738 1480 18770
rect 1512 18738 1552 18770
rect 1584 18738 1624 18770
rect 1656 18738 1696 18770
rect 1728 18738 1768 18770
rect 1800 18738 1840 18770
rect 1872 18738 1912 18770
rect 1944 18738 1984 18770
rect 2016 18738 2056 18770
rect 2088 18738 2128 18770
rect 2160 18738 2200 18770
rect 2232 18738 2272 18770
rect 2304 18738 2344 18770
rect 2376 18738 2416 18770
rect 2448 18738 2488 18770
rect 2520 18738 2560 18770
rect 2592 18738 2632 18770
rect 2664 18738 2704 18770
rect 2736 18738 2776 18770
rect 2808 18738 2848 18770
rect 2880 18738 2920 18770
rect 2952 18738 2992 18770
rect 3024 18738 3064 18770
rect 3096 18738 3136 18770
rect 3168 18738 3208 18770
rect 3240 18738 3280 18770
rect 3312 18738 3352 18770
rect 3384 18738 3424 18770
rect 3456 18738 3496 18770
rect 3528 18738 3568 18770
rect 3600 18738 3640 18770
rect 3672 18738 3712 18770
rect 3744 18738 3784 18770
rect 3816 18738 3856 18770
rect 3888 18738 4000 18770
rect 0 18698 4000 18738
rect 0 18666 112 18698
rect 144 18666 184 18698
rect 216 18666 256 18698
rect 288 18666 328 18698
rect 360 18666 400 18698
rect 432 18666 472 18698
rect 504 18666 544 18698
rect 576 18666 616 18698
rect 648 18666 688 18698
rect 720 18666 760 18698
rect 792 18666 832 18698
rect 864 18666 904 18698
rect 936 18666 976 18698
rect 1008 18666 1048 18698
rect 1080 18666 1120 18698
rect 1152 18666 1192 18698
rect 1224 18666 1264 18698
rect 1296 18666 1336 18698
rect 1368 18666 1408 18698
rect 1440 18666 1480 18698
rect 1512 18666 1552 18698
rect 1584 18666 1624 18698
rect 1656 18666 1696 18698
rect 1728 18666 1768 18698
rect 1800 18666 1840 18698
rect 1872 18666 1912 18698
rect 1944 18666 1984 18698
rect 2016 18666 2056 18698
rect 2088 18666 2128 18698
rect 2160 18666 2200 18698
rect 2232 18666 2272 18698
rect 2304 18666 2344 18698
rect 2376 18666 2416 18698
rect 2448 18666 2488 18698
rect 2520 18666 2560 18698
rect 2592 18666 2632 18698
rect 2664 18666 2704 18698
rect 2736 18666 2776 18698
rect 2808 18666 2848 18698
rect 2880 18666 2920 18698
rect 2952 18666 2992 18698
rect 3024 18666 3064 18698
rect 3096 18666 3136 18698
rect 3168 18666 3208 18698
rect 3240 18666 3280 18698
rect 3312 18666 3352 18698
rect 3384 18666 3424 18698
rect 3456 18666 3496 18698
rect 3528 18666 3568 18698
rect 3600 18666 3640 18698
rect 3672 18666 3712 18698
rect 3744 18666 3784 18698
rect 3816 18666 3856 18698
rect 3888 18666 4000 18698
rect 0 18626 4000 18666
rect 0 18594 112 18626
rect 144 18594 184 18626
rect 216 18594 256 18626
rect 288 18594 328 18626
rect 360 18594 400 18626
rect 432 18594 472 18626
rect 504 18594 544 18626
rect 576 18594 616 18626
rect 648 18594 688 18626
rect 720 18594 760 18626
rect 792 18594 832 18626
rect 864 18594 904 18626
rect 936 18594 976 18626
rect 1008 18594 1048 18626
rect 1080 18594 1120 18626
rect 1152 18594 1192 18626
rect 1224 18594 1264 18626
rect 1296 18594 1336 18626
rect 1368 18594 1408 18626
rect 1440 18594 1480 18626
rect 1512 18594 1552 18626
rect 1584 18594 1624 18626
rect 1656 18594 1696 18626
rect 1728 18594 1768 18626
rect 1800 18594 1840 18626
rect 1872 18594 1912 18626
rect 1944 18594 1984 18626
rect 2016 18594 2056 18626
rect 2088 18594 2128 18626
rect 2160 18594 2200 18626
rect 2232 18594 2272 18626
rect 2304 18594 2344 18626
rect 2376 18594 2416 18626
rect 2448 18594 2488 18626
rect 2520 18594 2560 18626
rect 2592 18594 2632 18626
rect 2664 18594 2704 18626
rect 2736 18594 2776 18626
rect 2808 18594 2848 18626
rect 2880 18594 2920 18626
rect 2952 18594 2992 18626
rect 3024 18594 3064 18626
rect 3096 18594 3136 18626
rect 3168 18594 3208 18626
rect 3240 18594 3280 18626
rect 3312 18594 3352 18626
rect 3384 18594 3424 18626
rect 3456 18594 3496 18626
rect 3528 18594 3568 18626
rect 3600 18594 3640 18626
rect 3672 18594 3712 18626
rect 3744 18594 3784 18626
rect 3816 18594 3856 18626
rect 3888 18594 4000 18626
rect 0 18554 4000 18594
rect 0 18522 112 18554
rect 144 18522 184 18554
rect 216 18522 256 18554
rect 288 18522 328 18554
rect 360 18522 400 18554
rect 432 18522 472 18554
rect 504 18522 544 18554
rect 576 18522 616 18554
rect 648 18522 688 18554
rect 720 18522 760 18554
rect 792 18522 832 18554
rect 864 18522 904 18554
rect 936 18522 976 18554
rect 1008 18522 1048 18554
rect 1080 18522 1120 18554
rect 1152 18522 1192 18554
rect 1224 18522 1264 18554
rect 1296 18522 1336 18554
rect 1368 18522 1408 18554
rect 1440 18522 1480 18554
rect 1512 18522 1552 18554
rect 1584 18522 1624 18554
rect 1656 18522 1696 18554
rect 1728 18522 1768 18554
rect 1800 18522 1840 18554
rect 1872 18522 1912 18554
rect 1944 18522 1984 18554
rect 2016 18522 2056 18554
rect 2088 18522 2128 18554
rect 2160 18522 2200 18554
rect 2232 18522 2272 18554
rect 2304 18522 2344 18554
rect 2376 18522 2416 18554
rect 2448 18522 2488 18554
rect 2520 18522 2560 18554
rect 2592 18522 2632 18554
rect 2664 18522 2704 18554
rect 2736 18522 2776 18554
rect 2808 18522 2848 18554
rect 2880 18522 2920 18554
rect 2952 18522 2992 18554
rect 3024 18522 3064 18554
rect 3096 18522 3136 18554
rect 3168 18522 3208 18554
rect 3240 18522 3280 18554
rect 3312 18522 3352 18554
rect 3384 18522 3424 18554
rect 3456 18522 3496 18554
rect 3528 18522 3568 18554
rect 3600 18522 3640 18554
rect 3672 18522 3712 18554
rect 3744 18522 3784 18554
rect 3816 18522 3856 18554
rect 3888 18522 4000 18554
rect 0 18482 4000 18522
rect 0 18450 112 18482
rect 144 18450 184 18482
rect 216 18450 256 18482
rect 288 18450 328 18482
rect 360 18450 400 18482
rect 432 18450 472 18482
rect 504 18450 544 18482
rect 576 18450 616 18482
rect 648 18450 688 18482
rect 720 18450 760 18482
rect 792 18450 832 18482
rect 864 18450 904 18482
rect 936 18450 976 18482
rect 1008 18450 1048 18482
rect 1080 18450 1120 18482
rect 1152 18450 1192 18482
rect 1224 18450 1264 18482
rect 1296 18450 1336 18482
rect 1368 18450 1408 18482
rect 1440 18450 1480 18482
rect 1512 18450 1552 18482
rect 1584 18450 1624 18482
rect 1656 18450 1696 18482
rect 1728 18450 1768 18482
rect 1800 18450 1840 18482
rect 1872 18450 1912 18482
rect 1944 18450 1984 18482
rect 2016 18450 2056 18482
rect 2088 18450 2128 18482
rect 2160 18450 2200 18482
rect 2232 18450 2272 18482
rect 2304 18450 2344 18482
rect 2376 18450 2416 18482
rect 2448 18450 2488 18482
rect 2520 18450 2560 18482
rect 2592 18450 2632 18482
rect 2664 18450 2704 18482
rect 2736 18450 2776 18482
rect 2808 18450 2848 18482
rect 2880 18450 2920 18482
rect 2952 18450 2992 18482
rect 3024 18450 3064 18482
rect 3096 18450 3136 18482
rect 3168 18450 3208 18482
rect 3240 18450 3280 18482
rect 3312 18450 3352 18482
rect 3384 18450 3424 18482
rect 3456 18450 3496 18482
rect 3528 18450 3568 18482
rect 3600 18450 3640 18482
rect 3672 18450 3712 18482
rect 3744 18450 3784 18482
rect 3816 18450 3856 18482
rect 3888 18450 4000 18482
rect 0 18410 4000 18450
rect 0 18378 112 18410
rect 144 18378 184 18410
rect 216 18378 256 18410
rect 288 18378 328 18410
rect 360 18378 400 18410
rect 432 18378 472 18410
rect 504 18378 544 18410
rect 576 18378 616 18410
rect 648 18378 688 18410
rect 720 18378 760 18410
rect 792 18378 832 18410
rect 864 18378 904 18410
rect 936 18378 976 18410
rect 1008 18378 1048 18410
rect 1080 18378 1120 18410
rect 1152 18378 1192 18410
rect 1224 18378 1264 18410
rect 1296 18378 1336 18410
rect 1368 18378 1408 18410
rect 1440 18378 1480 18410
rect 1512 18378 1552 18410
rect 1584 18378 1624 18410
rect 1656 18378 1696 18410
rect 1728 18378 1768 18410
rect 1800 18378 1840 18410
rect 1872 18378 1912 18410
rect 1944 18378 1984 18410
rect 2016 18378 2056 18410
rect 2088 18378 2128 18410
rect 2160 18378 2200 18410
rect 2232 18378 2272 18410
rect 2304 18378 2344 18410
rect 2376 18378 2416 18410
rect 2448 18378 2488 18410
rect 2520 18378 2560 18410
rect 2592 18378 2632 18410
rect 2664 18378 2704 18410
rect 2736 18378 2776 18410
rect 2808 18378 2848 18410
rect 2880 18378 2920 18410
rect 2952 18378 2992 18410
rect 3024 18378 3064 18410
rect 3096 18378 3136 18410
rect 3168 18378 3208 18410
rect 3240 18378 3280 18410
rect 3312 18378 3352 18410
rect 3384 18378 3424 18410
rect 3456 18378 3496 18410
rect 3528 18378 3568 18410
rect 3600 18378 3640 18410
rect 3672 18378 3712 18410
rect 3744 18378 3784 18410
rect 3816 18378 3856 18410
rect 3888 18378 4000 18410
rect 0 18338 4000 18378
rect 0 18306 112 18338
rect 144 18306 184 18338
rect 216 18306 256 18338
rect 288 18306 328 18338
rect 360 18306 400 18338
rect 432 18306 472 18338
rect 504 18306 544 18338
rect 576 18306 616 18338
rect 648 18306 688 18338
rect 720 18306 760 18338
rect 792 18306 832 18338
rect 864 18306 904 18338
rect 936 18306 976 18338
rect 1008 18306 1048 18338
rect 1080 18306 1120 18338
rect 1152 18306 1192 18338
rect 1224 18306 1264 18338
rect 1296 18306 1336 18338
rect 1368 18306 1408 18338
rect 1440 18306 1480 18338
rect 1512 18306 1552 18338
rect 1584 18306 1624 18338
rect 1656 18306 1696 18338
rect 1728 18306 1768 18338
rect 1800 18306 1840 18338
rect 1872 18306 1912 18338
rect 1944 18306 1984 18338
rect 2016 18306 2056 18338
rect 2088 18306 2128 18338
rect 2160 18306 2200 18338
rect 2232 18306 2272 18338
rect 2304 18306 2344 18338
rect 2376 18306 2416 18338
rect 2448 18306 2488 18338
rect 2520 18306 2560 18338
rect 2592 18306 2632 18338
rect 2664 18306 2704 18338
rect 2736 18306 2776 18338
rect 2808 18306 2848 18338
rect 2880 18306 2920 18338
rect 2952 18306 2992 18338
rect 3024 18306 3064 18338
rect 3096 18306 3136 18338
rect 3168 18306 3208 18338
rect 3240 18306 3280 18338
rect 3312 18306 3352 18338
rect 3384 18306 3424 18338
rect 3456 18306 3496 18338
rect 3528 18306 3568 18338
rect 3600 18306 3640 18338
rect 3672 18306 3712 18338
rect 3744 18306 3784 18338
rect 3816 18306 3856 18338
rect 3888 18306 4000 18338
rect 0 18266 4000 18306
rect 0 18234 112 18266
rect 144 18234 184 18266
rect 216 18234 256 18266
rect 288 18234 328 18266
rect 360 18234 400 18266
rect 432 18234 472 18266
rect 504 18234 544 18266
rect 576 18234 616 18266
rect 648 18234 688 18266
rect 720 18234 760 18266
rect 792 18234 832 18266
rect 864 18234 904 18266
rect 936 18234 976 18266
rect 1008 18234 1048 18266
rect 1080 18234 1120 18266
rect 1152 18234 1192 18266
rect 1224 18234 1264 18266
rect 1296 18234 1336 18266
rect 1368 18234 1408 18266
rect 1440 18234 1480 18266
rect 1512 18234 1552 18266
rect 1584 18234 1624 18266
rect 1656 18234 1696 18266
rect 1728 18234 1768 18266
rect 1800 18234 1840 18266
rect 1872 18234 1912 18266
rect 1944 18234 1984 18266
rect 2016 18234 2056 18266
rect 2088 18234 2128 18266
rect 2160 18234 2200 18266
rect 2232 18234 2272 18266
rect 2304 18234 2344 18266
rect 2376 18234 2416 18266
rect 2448 18234 2488 18266
rect 2520 18234 2560 18266
rect 2592 18234 2632 18266
rect 2664 18234 2704 18266
rect 2736 18234 2776 18266
rect 2808 18234 2848 18266
rect 2880 18234 2920 18266
rect 2952 18234 2992 18266
rect 3024 18234 3064 18266
rect 3096 18234 3136 18266
rect 3168 18234 3208 18266
rect 3240 18234 3280 18266
rect 3312 18234 3352 18266
rect 3384 18234 3424 18266
rect 3456 18234 3496 18266
rect 3528 18234 3568 18266
rect 3600 18234 3640 18266
rect 3672 18234 3712 18266
rect 3744 18234 3784 18266
rect 3816 18234 3856 18266
rect 3888 18234 4000 18266
rect 0 18194 4000 18234
rect 0 18162 112 18194
rect 144 18162 184 18194
rect 216 18162 256 18194
rect 288 18162 328 18194
rect 360 18162 400 18194
rect 432 18162 472 18194
rect 504 18162 544 18194
rect 576 18162 616 18194
rect 648 18162 688 18194
rect 720 18162 760 18194
rect 792 18162 832 18194
rect 864 18162 904 18194
rect 936 18162 976 18194
rect 1008 18162 1048 18194
rect 1080 18162 1120 18194
rect 1152 18162 1192 18194
rect 1224 18162 1264 18194
rect 1296 18162 1336 18194
rect 1368 18162 1408 18194
rect 1440 18162 1480 18194
rect 1512 18162 1552 18194
rect 1584 18162 1624 18194
rect 1656 18162 1696 18194
rect 1728 18162 1768 18194
rect 1800 18162 1840 18194
rect 1872 18162 1912 18194
rect 1944 18162 1984 18194
rect 2016 18162 2056 18194
rect 2088 18162 2128 18194
rect 2160 18162 2200 18194
rect 2232 18162 2272 18194
rect 2304 18162 2344 18194
rect 2376 18162 2416 18194
rect 2448 18162 2488 18194
rect 2520 18162 2560 18194
rect 2592 18162 2632 18194
rect 2664 18162 2704 18194
rect 2736 18162 2776 18194
rect 2808 18162 2848 18194
rect 2880 18162 2920 18194
rect 2952 18162 2992 18194
rect 3024 18162 3064 18194
rect 3096 18162 3136 18194
rect 3168 18162 3208 18194
rect 3240 18162 3280 18194
rect 3312 18162 3352 18194
rect 3384 18162 3424 18194
rect 3456 18162 3496 18194
rect 3528 18162 3568 18194
rect 3600 18162 3640 18194
rect 3672 18162 3712 18194
rect 3744 18162 3784 18194
rect 3816 18162 3856 18194
rect 3888 18162 4000 18194
rect 0 18112 4000 18162
rect 0 17848 4000 17912
rect 0 17816 112 17848
rect 144 17816 184 17848
rect 216 17816 256 17848
rect 288 17816 328 17848
rect 360 17816 400 17848
rect 432 17816 472 17848
rect 504 17816 544 17848
rect 576 17816 616 17848
rect 648 17816 688 17848
rect 720 17816 760 17848
rect 792 17816 832 17848
rect 864 17816 904 17848
rect 936 17816 976 17848
rect 1008 17816 1048 17848
rect 1080 17816 1120 17848
rect 1152 17816 1192 17848
rect 1224 17816 1264 17848
rect 1296 17816 1336 17848
rect 1368 17816 1408 17848
rect 1440 17816 1480 17848
rect 1512 17816 1552 17848
rect 1584 17816 1624 17848
rect 1656 17816 1696 17848
rect 1728 17816 1768 17848
rect 1800 17816 1840 17848
rect 1872 17816 1912 17848
rect 1944 17816 1984 17848
rect 2016 17816 2056 17848
rect 2088 17816 2128 17848
rect 2160 17816 2200 17848
rect 2232 17816 2272 17848
rect 2304 17816 2344 17848
rect 2376 17816 2416 17848
rect 2448 17816 2488 17848
rect 2520 17816 2560 17848
rect 2592 17816 2632 17848
rect 2664 17816 2704 17848
rect 2736 17816 2776 17848
rect 2808 17816 2848 17848
rect 2880 17816 2920 17848
rect 2952 17816 2992 17848
rect 3024 17816 3064 17848
rect 3096 17816 3136 17848
rect 3168 17816 3208 17848
rect 3240 17816 3280 17848
rect 3312 17816 3352 17848
rect 3384 17816 3424 17848
rect 3456 17816 3496 17848
rect 3528 17816 3568 17848
rect 3600 17816 3640 17848
rect 3672 17816 3712 17848
rect 3744 17816 3784 17848
rect 3816 17816 3856 17848
rect 3888 17816 4000 17848
rect 0 17776 4000 17816
rect 0 17744 112 17776
rect 144 17744 184 17776
rect 216 17744 256 17776
rect 288 17744 328 17776
rect 360 17744 400 17776
rect 432 17744 472 17776
rect 504 17744 544 17776
rect 576 17744 616 17776
rect 648 17744 688 17776
rect 720 17744 760 17776
rect 792 17744 832 17776
rect 864 17744 904 17776
rect 936 17744 976 17776
rect 1008 17744 1048 17776
rect 1080 17744 1120 17776
rect 1152 17744 1192 17776
rect 1224 17744 1264 17776
rect 1296 17744 1336 17776
rect 1368 17744 1408 17776
rect 1440 17744 1480 17776
rect 1512 17744 1552 17776
rect 1584 17744 1624 17776
rect 1656 17744 1696 17776
rect 1728 17744 1768 17776
rect 1800 17744 1840 17776
rect 1872 17744 1912 17776
rect 1944 17744 1984 17776
rect 2016 17744 2056 17776
rect 2088 17744 2128 17776
rect 2160 17744 2200 17776
rect 2232 17744 2272 17776
rect 2304 17744 2344 17776
rect 2376 17744 2416 17776
rect 2448 17744 2488 17776
rect 2520 17744 2560 17776
rect 2592 17744 2632 17776
rect 2664 17744 2704 17776
rect 2736 17744 2776 17776
rect 2808 17744 2848 17776
rect 2880 17744 2920 17776
rect 2952 17744 2992 17776
rect 3024 17744 3064 17776
rect 3096 17744 3136 17776
rect 3168 17744 3208 17776
rect 3240 17744 3280 17776
rect 3312 17744 3352 17776
rect 3384 17744 3424 17776
rect 3456 17744 3496 17776
rect 3528 17744 3568 17776
rect 3600 17744 3640 17776
rect 3672 17744 3712 17776
rect 3744 17744 3784 17776
rect 3816 17744 3856 17776
rect 3888 17744 4000 17776
rect 0 17704 4000 17744
rect 0 17672 112 17704
rect 144 17672 184 17704
rect 216 17672 256 17704
rect 288 17672 328 17704
rect 360 17672 400 17704
rect 432 17672 472 17704
rect 504 17672 544 17704
rect 576 17672 616 17704
rect 648 17672 688 17704
rect 720 17672 760 17704
rect 792 17672 832 17704
rect 864 17672 904 17704
rect 936 17672 976 17704
rect 1008 17672 1048 17704
rect 1080 17672 1120 17704
rect 1152 17672 1192 17704
rect 1224 17672 1264 17704
rect 1296 17672 1336 17704
rect 1368 17672 1408 17704
rect 1440 17672 1480 17704
rect 1512 17672 1552 17704
rect 1584 17672 1624 17704
rect 1656 17672 1696 17704
rect 1728 17672 1768 17704
rect 1800 17672 1840 17704
rect 1872 17672 1912 17704
rect 1944 17672 1984 17704
rect 2016 17672 2056 17704
rect 2088 17672 2128 17704
rect 2160 17672 2200 17704
rect 2232 17672 2272 17704
rect 2304 17672 2344 17704
rect 2376 17672 2416 17704
rect 2448 17672 2488 17704
rect 2520 17672 2560 17704
rect 2592 17672 2632 17704
rect 2664 17672 2704 17704
rect 2736 17672 2776 17704
rect 2808 17672 2848 17704
rect 2880 17672 2920 17704
rect 2952 17672 2992 17704
rect 3024 17672 3064 17704
rect 3096 17672 3136 17704
rect 3168 17672 3208 17704
rect 3240 17672 3280 17704
rect 3312 17672 3352 17704
rect 3384 17672 3424 17704
rect 3456 17672 3496 17704
rect 3528 17672 3568 17704
rect 3600 17672 3640 17704
rect 3672 17672 3712 17704
rect 3744 17672 3784 17704
rect 3816 17672 3856 17704
rect 3888 17672 4000 17704
rect 0 17632 4000 17672
rect 0 17600 112 17632
rect 144 17600 184 17632
rect 216 17600 256 17632
rect 288 17600 328 17632
rect 360 17600 400 17632
rect 432 17600 472 17632
rect 504 17600 544 17632
rect 576 17600 616 17632
rect 648 17600 688 17632
rect 720 17600 760 17632
rect 792 17600 832 17632
rect 864 17600 904 17632
rect 936 17600 976 17632
rect 1008 17600 1048 17632
rect 1080 17600 1120 17632
rect 1152 17600 1192 17632
rect 1224 17600 1264 17632
rect 1296 17600 1336 17632
rect 1368 17600 1408 17632
rect 1440 17600 1480 17632
rect 1512 17600 1552 17632
rect 1584 17600 1624 17632
rect 1656 17600 1696 17632
rect 1728 17600 1768 17632
rect 1800 17600 1840 17632
rect 1872 17600 1912 17632
rect 1944 17600 1984 17632
rect 2016 17600 2056 17632
rect 2088 17600 2128 17632
rect 2160 17600 2200 17632
rect 2232 17600 2272 17632
rect 2304 17600 2344 17632
rect 2376 17600 2416 17632
rect 2448 17600 2488 17632
rect 2520 17600 2560 17632
rect 2592 17600 2632 17632
rect 2664 17600 2704 17632
rect 2736 17600 2776 17632
rect 2808 17600 2848 17632
rect 2880 17600 2920 17632
rect 2952 17600 2992 17632
rect 3024 17600 3064 17632
rect 3096 17600 3136 17632
rect 3168 17600 3208 17632
rect 3240 17600 3280 17632
rect 3312 17600 3352 17632
rect 3384 17600 3424 17632
rect 3456 17600 3496 17632
rect 3528 17600 3568 17632
rect 3600 17600 3640 17632
rect 3672 17600 3712 17632
rect 3744 17600 3784 17632
rect 3816 17600 3856 17632
rect 3888 17600 4000 17632
rect 0 17560 4000 17600
rect 0 17528 112 17560
rect 144 17528 184 17560
rect 216 17528 256 17560
rect 288 17528 328 17560
rect 360 17528 400 17560
rect 432 17528 472 17560
rect 504 17528 544 17560
rect 576 17528 616 17560
rect 648 17528 688 17560
rect 720 17528 760 17560
rect 792 17528 832 17560
rect 864 17528 904 17560
rect 936 17528 976 17560
rect 1008 17528 1048 17560
rect 1080 17528 1120 17560
rect 1152 17528 1192 17560
rect 1224 17528 1264 17560
rect 1296 17528 1336 17560
rect 1368 17528 1408 17560
rect 1440 17528 1480 17560
rect 1512 17528 1552 17560
rect 1584 17528 1624 17560
rect 1656 17528 1696 17560
rect 1728 17528 1768 17560
rect 1800 17528 1840 17560
rect 1872 17528 1912 17560
rect 1944 17528 1984 17560
rect 2016 17528 2056 17560
rect 2088 17528 2128 17560
rect 2160 17528 2200 17560
rect 2232 17528 2272 17560
rect 2304 17528 2344 17560
rect 2376 17528 2416 17560
rect 2448 17528 2488 17560
rect 2520 17528 2560 17560
rect 2592 17528 2632 17560
rect 2664 17528 2704 17560
rect 2736 17528 2776 17560
rect 2808 17528 2848 17560
rect 2880 17528 2920 17560
rect 2952 17528 2992 17560
rect 3024 17528 3064 17560
rect 3096 17528 3136 17560
rect 3168 17528 3208 17560
rect 3240 17528 3280 17560
rect 3312 17528 3352 17560
rect 3384 17528 3424 17560
rect 3456 17528 3496 17560
rect 3528 17528 3568 17560
rect 3600 17528 3640 17560
rect 3672 17528 3712 17560
rect 3744 17528 3784 17560
rect 3816 17528 3856 17560
rect 3888 17528 4000 17560
rect 0 17488 4000 17528
rect 0 17456 112 17488
rect 144 17456 184 17488
rect 216 17456 256 17488
rect 288 17456 328 17488
rect 360 17456 400 17488
rect 432 17456 472 17488
rect 504 17456 544 17488
rect 576 17456 616 17488
rect 648 17456 688 17488
rect 720 17456 760 17488
rect 792 17456 832 17488
rect 864 17456 904 17488
rect 936 17456 976 17488
rect 1008 17456 1048 17488
rect 1080 17456 1120 17488
rect 1152 17456 1192 17488
rect 1224 17456 1264 17488
rect 1296 17456 1336 17488
rect 1368 17456 1408 17488
rect 1440 17456 1480 17488
rect 1512 17456 1552 17488
rect 1584 17456 1624 17488
rect 1656 17456 1696 17488
rect 1728 17456 1768 17488
rect 1800 17456 1840 17488
rect 1872 17456 1912 17488
rect 1944 17456 1984 17488
rect 2016 17456 2056 17488
rect 2088 17456 2128 17488
rect 2160 17456 2200 17488
rect 2232 17456 2272 17488
rect 2304 17456 2344 17488
rect 2376 17456 2416 17488
rect 2448 17456 2488 17488
rect 2520 17456 2560 17488
rect 2592 17456 2632 17488
rect 2664 17456 2704 17488
rect 2736 17456 2776 17488
rect 2808 17456 2848 17488
rect 2880 17456 2920 17488
rect 2952 17456 2992 17488
rect 3024 17456 3064 17488
rect 3096 17456 3136 17488
rect 3168 17456 3208 17488
rect 3240 17456 3280 17488
rect 3312 17456 3352 17488
rect 3384 17456 3424 17488
rect 3456 17456 3496 17488
rect 3528 17456 3568 17488
rect 3600 17456 3640 17488
rect 3672 17456 3712 17488
rect 3744 17456 3784 17488
rect 3816 17456 3856 17488
rect 3888 17456 4000 17488
rect 0 17416 4000 17456
rect 0 17384 112 17416
rect 144 17384 184 17416
rect 216 17384 256 17416
rect 288 17384 328 17416
rect 360 17384 400 17416
rect 432 17384 472 17416
rect 504 17384 544 17416
rect 576 17384 616 17416
rect 648 17384 688 17416
rect 720 17384 760 17416
rect 792 17384 832 17416
rect 864 17384 904 17416
rect 936 17384 976 17416
rect 1008 17384 1048 17416
rect 1080 17384 1120 17416
rect 1152 17384 1192 17416
rect 1224 17384 1264 17416
rect 1296 17384 1336 17416
rect 1368 17384 1408 17416
rect 1440 17384 1480 17416
rect 1512 17384 1552 17416
rect 1584 17384 1624 17416
rect 1656 17384 1696 17416
rect 1728 17384 1768 17416
rect 1800 17384 1840 17416
rect 1872 17384 1912 17416
rect 1944 17384 1984 17416
rect 2016 17384 2056 17416
rect 2088 17384 2128 17416
rect 2160 17384 2200 17416
rect 2232 17384 2272 17416
rect 2304 17384 2344 17416
rect 2376 17384 2416 17416
rect 2448 17384 2488 17416
rect 2520 17384 2560 17416
rect 2592 17384 2632 17416
rect 2664 17384 2704 17416
rect 2736 17384 2776 17416
rect 2808 17384 2848 17416
rect 2880 17384 2920 17416
rect 2952 17384 2992 17416
rect 3024 17384 3064 17416
rect 3096 17384 3136 17416
rect 3168 17384 3208 17416
rect 3240 17384 3280 17416
rect 3312 17384 3352 17416
rect 3384 17384 3424 17416
rect 3456 17384 3496 17416
rect 3528 17384 3568 17416
rect 3600 17384 3640 17416
rect 3672 17384 3712 17416
rect 3744 17384 3784 17416
rect 3816 17384 3856 17416
rect 3888 17384 4000 17416
rect 0 17344 4000 17384
rect 0 17312 112 17344
rect 144 17312 184 17344
rect 216 17312 256 17344
rect 288 17312 328 17344
rect 360 17312 400 17344
rect 432 17312 472 17344
rect 504 17312 544 17344
rect 576 17312 616 17344
rect 648 17312 688 17344
rect 720 17312 760 17344
rect 792 17312 832 17344
rect 864 17312 904 17344
rect 936 17312 976 17344
rect 1008 17312 1048 17344
rect 1080 17312 1120 17344
rect 1152 17312 1192 17344
rect 1224 17312 1264 17344
rect 1296 17312 1336 17344
rect 1368 17312 1408 17344
rect 1440 17312 1480 17344
rect 1512 17312 1552 17344
rect 1584 17312 1624 17344
rect 1656 17312 1696 17344
rect 1728 17312 1768 17344
rect 1800 17312 1840 17344
rect 1872 17312 1912 17344
rect 1944 17312 1984 17344
rect 2016 17312 2056 17344
rect 2088 17312 2128 17344
rect 2160 17312 2200 17344
rect 2232 17312 2272 17344
rect 2304 17312 2344 17344
rect 2376 17312 2416 17344
rect 2448 17312 2488 17344
rect 2520 17312 2560 17344
rect 2592 17312 2632 17344
rect 2664 17312 2704 17344
rect 2736 17312 2776 17344
rect 2808 17312 2848 17344
rect 2880 17312 2920 17344
rect 2952 17312 2992 17344
rect 3024 17312 3064 17344
rect 3096 17312 3136 17344
rect 3168 17312 3208 17344
rect 3240 17312 3280 17344
rect 3312 17312 3352 17344
rect 3384 17312 3424 17344
rect 3456 17312 3496 17344
rect 3528 17312 3568 17344
rect 3600 17312 3640 17344
rect 3672 17312 3712 17344
rect 3744 17312 3784 17344
rect 3816 17312 3856 17344
rect 3888 17312 4000 17344
rect 0 17272 4000 17312
rect 0 17240 112 17272
rect 144 17240 184 17272
rect 216 17240 256 17272
rect 288 17240 328 17272
rect 360 17240 400 17272
rect 432 17240 472 17272
rect 504 17240 544 17272
rect 576 17240 616 17272
rect 648 17240 688 17272
rect 720 17240 760 17272
rect 792 17240 832 17272
rect 864 17240 904 17272
rect 936 17240 976 17272
rect 1008 17240 1048 17272
rect 1080 17240 1120 17272
rect 1152 17240 1192 17272
rect 1224 17240 1264 17272
rect 1296 17240 1336 17272
rect 1368 17240 1408 17272
rect 1440 17240 1480 17272
rect 1512 17240 1552 17272
rect 1584 17240 1624 17272
rect 1656 17240 1696 17272
rect 1728 17240 1768 17272
rect 1800 17240 1840 17272
rect 1872 17240 1912 17272
rect 1944 17240 1984 17272
rect 2016 17240 2056 17272
rect 2088 17240 2128 17272
rect 2160 17240 2200 17272
rect 2232 17240 2272 17272
rect 2304 17240 2344 17272
rect 2376 17240 2416 17272
rect 2448 17240 2488 17272
rect 2520 17240 2560 17272
rect 2592 17240 2632 17272
rect 2664 17240 2704 17272
rect 2736 17240 2776 17272
rect 2808 17240 2848 17272
rect 2880 17240 2920 17272
rect 2952 17240 2992 17272
rect 3024 17240 3064 17272
rect 3096 17240 3136 17272
rect 3168 17240 3208 17272
rect 3240 17240 3280 17272
rect 3312 17240 3352 17272
rect 3384 17240 3424 17272
rect 3456 17240 3496 17272
rect 3528 17240 3568 17272
rect 3600 17240 3640 17272
rect 3672 17240 3712 17272
rect 3744 17240 3784 17272
rect 3816 17240 3856 17272
rect 3888 17240 4000 17272
rect 0 17200 4000 17240
rect 0 17168 112 17200
rect 144 17168 184 17200
rect 216 17168 256 17200
rect 288 17168 328 17200
rect 360 17168 400 17200
rect 432 17168 472 17200
rect 504 17168 544 17200
rect 576 17168 616 17200
rect 648 17168 688 17200
rect 720 17168 760 17200
rect 792 17168 832 17200
rect 864 17168 904 17200
rect 936 17168 976 17200
rect 1008 17168 1048 17200
rect 1080 17168 1120 17200
rect 1152 17168 1192 17200
rect 1224 17168 1264 17200
rect 1296 17168 1336 17200
rect 1368 17168 1408 17200
rect 1440 17168 1480 17200
rect 1512 17168 1552 17200
rect 1584 17168 1624 17200
rect 1656 17168 1696 17200
rect 1728 17168 1768 17200
rect 1800 17168 1840 17200
rect 1872 17168 1912 17200
rect 1944 17168 1984 17200
rect 2016 17168 2056 17200
rect 2088 17168 2128 17200
rect 2160 17168 2200 17200
rect 2232 17168 2272 17200
rect 2304 17168 2344 17200
rect 2376 17168 2416 17200
rect 2448 17168 2488 17200
rect 2520 17168 2560 17200
rect 2592 17168 2632 17200
rect 2664 17168 2704 17200
rect 2736 17168 2776 17200
rect 2808 17168 2848 17200
rect 2880 17168 2920 17200
rect 2952 17168 2992 17200
rect 3024 17168 3064 17200
rect 3096 17168 3136 17200
rect 3168 17168 3208 17200
rect 3240 17168 3280 17200
rect 3312 17168 3352 17200
rect 3384 17168 3424 17200
rect 3456 17168 3496 17200
rect 3528 17168 3568 17200
rect 3600 17168 3640 17200
rect 3672 17168 3712 17200
rect 3744 17168 3784 17200
rect 3816 17168 3856 17200
rect 3888 17168 4000 17200
rect 0 17128 4000 17168
rect 0 17096 112 17128
rect 144 17096 184 17128
rect 216 17096 256 17128
rect 288 17096 328 17128
rect 360 17096 400 17128
rect 432 17096 472 17128
rect 504 17096 544 17128
rect 576 17096 616 17128
rect 648 17096 688 17128
rect 720 17096 760 17128
rect 792 17096 832 17128
rect 864 17096 904 17128
rect 936 17096 976 17128
rect 1008 17096 1048 17128
rect 1080 17096 1120 17128
rect 1152 17096 1192 17128
rect 1224 17096 1264 17128
rect 1296 17096 1336 17128
rect 1368 17096 1408 17128
rect 1440 17096 1480 17128
rect 1512 17096 1552 17128
rect 1584 17096 1624 17128
rect 1656 17096 1696 17128
rect 1728 17096 1768 17128
rect 1800 17096 1840 17128
rect 1872 17096 1912 17128
rect 1944 17096 1984 17128
rect 2016 17096 2056 17128
rect 2088 17096 2128 17128
rect 2160 17096 2200 17128
rect 2232 17096 2272 17128
rect 2304 17096 2344 17128
rect 2376 17096 2416 17128
rect 2448 17096 2488 17128
rect 2520 17096 2560 17128
rect 2592 17096 2632 17128
rect 2664 17096 2704 17128
rect 2736 17096 2776 17128
rect 2808 17096 2848 17128
rect 2880 17096 2920 17128
rect 2952 17096 2992 17128
rect 3024 17096 3064 17128
rect 3096 17096 3136 17128
rect 3168 17096 3208 17128
rect 3240 17096 3280 17128
rect 3312 17096 3352 17128
rect 3384 17096 3424 17128
rect 3456 17096 3496 17128
rect 3528 17096 3568 17128
rect 3600 17096 3640 17128
rect 3672 17096 3712 17128
rect 3744 17096 3784 17128
rect 3816 17096 3856 17128
rect 3888 17096 4000 17128
rect 0 17056 4000 17096
rect 0 17024 112 17056
rect 144 17024 184 17056
rect 216 17024 256 17056
rect 288 17024 328 17056
rect 360 17024 400 17056
rect 432 17024 472 17056
rect 504 17024 544 17056
rect 576 17024 616 17056
rect 648 17024 688 17056
rect 720 17024 760 17056
rect 792 17024 832 17056
rect 864 17024 904 17056
rect 936 17024 976 17056
rect 1008 17024 1048 17056
rect 1080 17024 1120 17056
rect 1152 17024 1192 17056
rect 1224 17024 1264 17056
rect 1296 17024 1336 17056
rect 1368 17024 1408 17056
rect 1440 17024 1480 17056
rect 1512 17024 1552 17056
rect 1584 17024 1624 17056
rect 1656 17024 1696 17056
rect 1728 17024 1768 17056
rect 1800 17024 1840 17056
rect 1872 17024 1912 17056
rect 1944 17024 1984 17056
rect 2016 17024 2056 17056
rect 2088 17024 2128 17056
rect 2160 17024 2200 17056
rect 2232 17024 2272 17056
rect 2304 17024 2344 17056
rect 2376 17024 2416 17056
rect 2448 17024 2488 17056
rect 2520 17024 2560 17056
rect 2592 17024 2632 17056
rect 2664 17024 2704 17056
rect 2736 17024 2776 17056
rect 2808 17024 2848 17056
rect 2880 17024 2920 17056
rect 2952 17024 2992 17056
rect 3024 17024 3064 17056
rect 3096 17024 3136 17056
rect 3168 17024 3208 17056
rect 3240 17024 3280 17056
rect 3312 17024 3352 17056
rect 3384 17024 3424 17056
rect 3456 17024 3496 17056
rect 3528 17024 3568 17056
rect 3600 17024 3640 17056
rect 3672 17024 3712 17056
rect 3744 17024 3784 17056
rect 3816 17024 3856 17056
rect 3888 17024 4000 17056
rect 0 16984 4000 17024
rect 0 16952 112 16984
rect 144 16952 184 16984
rect 216 16952 256 16984
rect 288 16952 328 16984
rect 360 16952 400 16984
rect 432 16952 472 16984
rect 504 16952 544 16984
rect 576 16952 616 16984
rect 648 16952 688 16984
rect 720 16952 760 16984
rect 792 16952 832 16984
rect 864 16952 904 16984
rect 936 16952 976 16984
rect 1008 16952 1048 16984
rect 1080 16952 1120 16984
rect 1152 16952 1192 16984
rect 1224 16952 1264 16984
rect 1296 16952 1336 16984
rect 1368 16952 1408 16984
rect 1440 16952 1480 16984
rect 1512 16952 1552 16984
rect 1584 16952 1624 16984
rect 1656 16952 1696 16984
rect 1728 16952 1768 16984
rect 1800 16952 1840 16984
rect 1872 16952 1912 16984
rect 1944 16952 1984 16984
rect 2016 16952 2056 16984
rect 2088 16952 2128 16984
rect 2160 16952 2200 16984
rect 2232 16952 2272 16984
rect 2304 16952 2344 16984
rect 2376 16952 2416 16984
rect 2448 16952 2488 16984
rect 2520 16952 2560 16984
rect 2592 16952 2632 16984
rect 2664 16952 2704 16984
rect 2736 16952 2776 16984
rect 2808 16952 2848 16984
rect 2880 16952 2920 16984
rect 2952 16952 2992 16984
rect 3024 16952 3064 16984
rect 3096 16952 3136 16984
rect 3168 16952 3208 16984
rect 3240 16952 3280 16984
rect 3312 16952 3352 16984
rect 3384 16952 3424 16984
rect 3456 16952 3496 16984
rect 3528 16952 3568 16984
rect 3600 16952 3640 16984
rect 3672 16952 3712 16984
rect 3744 16952 3784 16984
rect 3816 16952 3856 16984
rect 3888 16952 4000 16984
rect 0 16912 4000 16952
rect 0 16880 112 16912
rect 144 16880 184 16912
rect 216 16880 256 16912
rect 288 16880 328 16912
rect 360 16880 400 16912
rect 432 16880 472 16912
rect 504 16880 544 16912
rect 576 16880 616 16912
rect 648 16880 688 16912
rect 720 16880 760 16912
rect 792 16880 832 16912
rect 864 16880 904 16912
rect 936 16880 976 16912
rect 1008 16880 1048 16912
rect 1080 16880 1120 16912
rect 1152 16880 1192 16912
rect 1224 16880 1264 16912
rect 1296 16880 1336 16912
rect 1368 16880 1408 16912
rect 1440 16880 1480 16912
rect 1512 16880 1552 16912
rect 1584 16880 1624 16912
rect 1656 16880 1696 16912
rect 1728 16880 1768 16912
rect 1800 16880 1840 16912
rect 1872 16880 1912 16912
rect 1944 16880 1984 16912
rect 2016 16880 2056 16912
rect 2088 16880 2128 16912
rect 2160 16880 2200 16912
rect 2232 16880 2272 16912
rect 2304 16880 2344 16912
rect 2376 16880 2416 16912
rect 2448 16880 2488 16912
rect 2520 16880 2560 16912
rect 2592 16880 2632 16912
rect 2664 16880 2704 16912
rect 2736 16880 2776 16912
rect 2808 16880 2848 16912
rect 2880 16880 2920 16912
rect 2952 16880 2992 16912
rect 3024 16880 3064 16912
rect 3096 16880 3136 16912
rect 3168 16880 3208 16912
rect 3240 16880 3280 16912
rect 3312 16880 3352 16912
rect 3384 16880 3424 16912
rect 3456 16880 3496 16912
rect 3528 16880 3568 16912
rect 3600 16880 3640 16912
rect 3672 16880 3712 16912
rect 3744 16880 3784 16912
rect 3816 16880 3856 16912
rect 3888 16880 4000 16912
rect 0 16840 4000 16880
rect 0 16808 112 16840
rect 144 16808 184 16840
rect 216 16808 256 16840
rect 288 16808 328 16840
rect 360 16808 400 16840
rect 432 16808 472 16840
rect 504 16808 544 16840
rect 576 16808 616 16840
rect 648 16808 688 16840
rect 720 16808 760 16840
rect 792 16808 832 16840
rect 864 16808 904 16840
rect 936 16808 976 16840
rect 1008 16808 1048 16840
rect 1080 16808 1120 16840
rect 1152 16808 1192 16840
rect 1224 16808 1264 16840
rect 1296 16808 1336 16840
rect 1368 16808 1408 16840
rect 1440 16808 1480 16840
rect 1512 16808 1552 16840
rect 1584 16808 1624 16840
rect 1656 16808 1696 16840
rect 1728 16808 1768 16840
rect 1800 16808 1840 16840
rect 1872 16808 1912 16840
rect 1944 16808 1984 16840
rect 2016 16808 2056 16840
rect 2088 16808 2128 16840
rect 2160 16808 2200 16840
rect 2232 16808 2272 16840
rect 2304 16808 2344 16840
rect 2376 16808 2416 16840
rect 2448 16808 2488 16840
rect 2520 16808 2560 16840
rect 2592 16808 2632 16840
rect 2664 16808 2704 16840
rect 2736 16808 2776 16840
rect 2808 16808 2848 16840
rect 2880 16808 2920 16840
rect 2952 16808 2992 16840
rect 3024 16808 3064 16840
rect 3096 16808 3136 16840
rect 3168 16808 3208 16840
rect 3240 16808 3280 16840
rect 3312 16808 3352 16840
rect 3384 16808 3424 16840
rect 3456 16808 3496 16840
rect 3528 16808 3568 16840
rect 3600 16808 3640 16840
rect 3672 16808 3712 16840
rect 3744 16808 3784 16840
rect 3816 16808 3856 16840
rect 3888 16808 4000 16840
rect 0 16768 4000 16808
rect 0 16736 112 16768
rect 144 16736 184 16768
rect 216 16736 256 16768
rect 288 16736 328 16768
rect 360 16736 400 16768
rect 432 16736 472 16768
rect 504 16736 544 16768
rect 576 16736 616 16768
rect 648 16736 688 16768
rect 720 16736 760 16768
rect 792 16736 832 16768
rect 864 16736 904 16768
rect 936 16736 976 16768
rect 1008 16736 1048 16768
rect 1080 16736 1120 16768
rect 1152 16736 1192 16768
rect 1224 16736 1264 16768
rect 1296 16736 1336 16768
rect 1368 16736 1408 16768
rect 1440 16736 1480 16768
rect 1512 16736 1552 16768
rect 1584 16736 1624 16768
rect 1656 16736 1696 16768
rect 1728 16736 1768 16768
rect 1800 16736 1840 16768
rect 1872 16736 1912 16768
rect 1944 16736 1984 16768
rect 2016 16736 2056 16768
rect 2088 16736 2128 16768
rect 2160 16736 2200 16768
rect 2232 16736 2272 16768
rect 2304 16736 2344 16768
rect 2376 16736 2416 16768
rect 2448 16736 2488 16768
rect 2520 16736 2560 16768
rect 2592 16736 2632 16768
rect 2664 16736 2704 16768
rect 2736 16736 2776 16768
rect 2808 16736 2848 16768
rect 2880 16736 2920 16768
rect 2952 16736 2992 16768
rect 3024 16736 3064 16768
rect 3096 16736 3136 16768
rect 3168 16736 3208 16768
rect 3240 16736 3280 16768
rect 3312 16736 3352 16768
rect 3384 16736 3424 16768
rect 3456 16736 3496 16768
rect 3528 16736 3568 16768
rect 3600 16736 3640 16768
rect 3672 16736 3712 16768
rect 3744 16736 3784 16768
rect 3816 16736 3856 16768
rect 3888 16736 4000 16768
rect 0 16696 4000 16736
rect 0 16664 112 16696
rect 144 16664 184 16696
rect 216 16664 256 16696
rect 288 16664 328 16696
rect 360 16664 400 16696
rect 432 16664 472 16696
rect 504 16664 544 16696
rect 576 16664 616 16696
rect 648 16664 688 16696
rect 720 16664 760 16696
rect 792 16664 832 16696
rect 864 16664 904 16696
rect 936 16664 976 16696
rect 1008 16664 1048 16696
rect 1080 16664 1120 16696
rect 1152 16664 1192 16696
rect 1224 16664 1264 16696
rect 1296 16664 1336 16696
rect 1368 16664 1408 16696
rect 1440 16664 1480 16696
rect 1512 16664 1552 16696
rect 1584 16664 1624 16696
rect 1656 16664 1696 16696
rect 1728 16664 1768 16696
rect 1800 16664 1840 16696
rect 1872 16664 1912 16696
rect 1944 16664 1984 16696
rect 2016 16664 2056 16696
rect 2088 16664 2128 16696
rect 2160 16664 2200 16696
rect 2232 16664 2272 16696
rect 2304 16664 2344 16696
rect 2376 16664 2416 16696
rect 2448 16664 2488 16696
rect 2520 16664 2560 16696
rect 2592 16664 2632 16696
rect 2664 16664 2704 16696
rect 2736 16664 2776 16696
rect 2808 16664 2848 16696
rect 2880 16664 2920 16696
rect 2952 16664 2992 16696
rect 3024 16664 3064 16696
rect 3096 16664 3136 16696
rect 3168 16664 3208 16696
rect 3240 16664 3280 16696
rect 3312 16664 3352 16696
rect 3384 16664 3424 16696
rect 3456 16664 3496 16696
rect 3528 16664 3568 16696
rect 3600 16664 3640 16696
rect 3672 16664 3712 16696
rect 3744 16664 3784 16696
rect 3816 16664 3856 16696
rect 3888 16664 4000 16696
rect 0 16624 4000 16664
rect 0 16592 112 16624
rect 144 16592 184 16624
rect 216 16592 256 16624
rect 288 16592 328 16624
rect 360 16592 400 16624
rect 432 16592 472 16624
rect 504 16592 544 16624
rect 576 16592 616 16624
rect 648 16592 688 16624
rect 720 16592 760 16624
rect 792 16592 832 16624
rect 864 16592 904 16624
rect 936 16592 976 16624
rect 1008 16592 1048 16624
rect 1080 16592 1120 16624
rect 1152 16592 1192 16624
rect 1224 16592 1264 16624
rect 1296 16592 1336 16624
rect 1368 16592 1408 16624
rect 1440 16592 1480 16624
rect 1512 16592 1552 16624
rect 1584 16592 1624 16624
rect 1656 16592 1696 16624
rect 1728 16592 1768 16624
rect 1800 16592 1840 16624
rect 1872 16592 1912 16624
rect 1944 16592 1984 16624
rect 2016 16592 2056 16624
rect 2088 16592 2128 16624
rect 2160 16592 2200 16624
rect 2232 16592 2272 16624
rect 2304 16592 2344 16624
rect 2376 16592 2416 16624
rect 2448 16592 2488 16624
rect 2520 16592 2560 16624
rect 2592 16592 2632 16624
rect 2664 16592 2704 16624
rect 2736 16592 2776 16624
rect 2808 16592 2848 16624
rect 2880 16592 2920 16624
rect 2952 16592 2992 16624
rect 3024 16592 3064 16624
rect 3096 16592 3136 16624
rect 3168 16592 3208 16624
rect 3240 16592 3280 16624
rect 3312 16592 3352 16624
rect 3384 16592 3424 16624
rect 3456 16592 3496 16624
rect 3528 16592 3568 16624
rect 3600 16592 3640 16624
rect 3672 16592 3712 16624
rect 3744 16592 3784 16624
rect 3816 16592 3856 16624
rect 3888 16592 4000 16624
rect 0 16552 4000 16592
rect 0 16520 112 16552
rect 144 16520 184 16552
rect 216 16520 256 16552
rect 288 16520 328 16552
rect 360 16520 400 16552
rect 432 16520 472 16552
rect 504 16520 544 16552
rect 576 16520 616 16552
rect 648 16520 688 16552
rect 720 16520 760 16552
rect 792 16520 832 16552
rect 864 16520 904 16552
rect 936 16520 976 16552
rect 1008 16520 1048 16552
rect 1080 16520 1120 16552
rect 1152 16520 1192 16552
rect 1224 16520 1264 16552
rect 1296 16520 1336 16552
rect 1368 16520 1408 16552
rect 1440 16520 1480 16552
rect 1512 16520 1552 16552
rect 1584 16520 1624 16552
rect 1656 16520 1696 16552
rect 1728 16520 1768 16552
rect 1800 16520 1840 16552
rect 1872 16520 1912 16552
rect 1944 16520 1984 16552
rect 2016 16520 2056 16552
rect 2088 16520 2128 16552
rect 2160 16520 2200 16552
rect 2232 16520 2272 16552
rect 2304 16520 2344 16552
rect 2376 16520 2416 16552
rect 2448 16520 2488 16552
rect 2520 16520 2560 16552
rect 2592 16520 2632 16552
rect 2664 16520 2704 16552
rect 2736 16520 2776 16552
rect 2808 16520 2848 16552
rect 2880 16520 2920 16552
rect 2952 16520 2992 16552
rect 3024 16520 3064 16552
rect 3096 16520 3136 16552
rect 3168 16520 3208 16552
rect 3240 16520 3280 16552
rect 3312 16520 3352 16552
rect 3384 16520 3424 16552
rect 3456 16520 3496 16552
rect 3528 16520 3568 16552
rect 3600 16520 3640 16552
rect 3672 16520 3712 16552
rect 3744 16520 3784 16552
rect 3816 16520 3856 16552
rect 3888 16520 4000 16552
rect 0 16480 4000 16520
rect 0 16448 112 16480
rect 144 16448 184 16480
rect 216 16448 256 16480
rect 288 16448 328 16480
rect 360 16448 400 16480
rect 432 16448 472 16480
rect 504 16448 544 16480
rect 576 16448 616 16480
rect 648 16448 688 16480
rect 720 16448 760 16480
rect 792 16448 832 16480
rect 864 16448 904 16480
rect 936 16448 976 16480
rect 1008 16448 1048 16480
rect 1080 16448 1120 16480
rect 1152 16448 1192 16480
rect 1224 16448 1264 16480
rect 1296 16448 1336 16480
rect 1368 16448 1408 16480
rect 1440 16448 1480 16480
rect 1512 16448 1552 16480
rect 1584 16448 1624 16480
rect 1656 16448 1696 16480
rect 1728 16448 1768 16480
rect 1800 16448 1840 16480
rect 1872 16448 1912 16480
rect 1944 16448 1984 16480
rect 2016 16448 2056 16480
rect 2088 16448 2128 16480
rect 2160 16448 2200 16480
rect 2232 16448 2272 16480
rect 2304 16448 2344 16480
rect 2376 16448 2416 16480
rect 2448 16448 2488 16480
rect 2520 16448 2560 16480
rect 2592 16448 2632 16480
rect 2664 16448 2704 16480
rect 2736 16448 2776 16480
rect 2808 16448 2848 16480
rect 2880 16448 2920 16480
rect 2952 16448 2992 16480
rect 3024 16448 3064 16480
rect 3096 16448 3136 16480
rect 3168 16448 3208 16480
rect 3240 16448 3280 16480
rect 3312 16448 3352 16480
rect 3384 16448 3424 16480
rect 3456 16448 3496 16480
rect 3528 16448 3568 16480
rect 3600 16448 3640 16480
rect 3672 16448 3712 16480
rect 3744 16448 3784 16480
rect 3816 16448 3856 16480
rect 3888 16448 4000 16480
rect 0 16408 4000 16448
rect 0 16376 112 16408
rect 144 16376 184 16408
rect 216 16376 256 16408
rect 288 16376 328 16408
rect 360 16376 400 16408
rect 432 16376 472 16408
rect 504 16376 544 16408
rect 576 16376 616 16408
rect 648 16376 688 16408
rect 720 16376 760 16408
rect 792 16376 832 16408
rect 864 16376 904 16408
rect 936 16376 976 16408
rect 1008 16376 1048 16408
rect 1080 16376 1120 16408
rect 1152 16376 1192 16408
rect 1224 16376 1264 16408
rect 1296 16376 1336 16408
rect 1368 16376 1408 16408
rect 1440 16376 1480 16408
rect 1512 16376 1552 16408
rect 1584 16376 1624 16408
rect 1656 16376 1696 16408
rect 1728 16376 1768 16408
rect 1800 16376 1840 16408
rect 1872 16376 1912 16408
rect 1944 16376 1984 16408
rect 2016 16376 2056 16408
rect 2088 16376 2128 16408
rect 2160 16376 2200 16408
rect 2232 16376 2272 16408
rect 2304 16376 2344 16408
rect 2376 16376 2416 16408
rect 2448 16376 2488 16408
rect 2520 16376 2560 16408
rect 2592 16376 2632 16408
rect 2664 16376 2704 16408
rect 2736 16376 2776 16408
rect 2808 16376 2848 16408
rect 2880 16376 2920 16408
rect 2952 16376 2992 16408
rect 3024 16376 3064 16408
rect 3096 16376 3136 16408
rect 3168 16376 3208 16408
rect 3240 16376 3280 16408
rect 3312 16376 3352 16408
rect 3384 16376 3424 16408
rect 3456 16376 3496 16408
rect 3528 16376 3568 16408
rect 3600 16376 3640 16408
rect 3672 16376 3712 16408
rect 3744 16376 3784 16408
rect 3816 16376 3856 16408
rect 3888 16376 4000 16408
rect 0 16336 4000 16376
rect 0 16304 112 16336
rect 144 16304 184 16336
rect 216 16304 256 16336
rect 288 16304 328 16336
rect 360 16304 400 16336
rect 432 16304 472 16336
rect 504 16304 544 16336
rect 576 16304 616 16336
rect 648 16304 688 16336
rect 720 16304 760 16336
rect 792 16304 832 16336
rect 864 16304 904 16336
rect 936 16304 976 16336
rect 1008 16304 1048 16336
rect 1080 16304 1120 16336
rect 1152 16304 1192 16336
rect 1224 16304 1264 16336
rect 1296 16304 1336 16336
rect 1368 16304 1408 16336
rect 1440 16304 1480 16336
rect 1512 16304 1552 16336
rect 1584 16304 1624 16336
rect 1656 16304 1696 16336
rect 1728 16304 1768 16336
rect 1800 16304 1840 16336
rect 1872 16304 1912 16336
rect 1944 16304 1984 16336
rect 2016 16304 2056 16336
rect 2088 16304 2128 16336
rect 2160 16304 2200 16336
rect 2232 16304 2272 16336
rect 2304 16304 2344 16336
rect 2376 16304 2416 16336
rect 2448 16304 2488 16336
rect 2520 16304 2560 16336
rect 2592 16304 2632 16336
rect 2664 16304 2704 16336
rect 2736 16304 2776 16336
rect 2808 16304 2848 16336
rect 2880 16304 2920 16336
rect 2952 16304 2992 16336
rect 3024 16304 3064 16336
rect 3096 16304 3136 16336
rect 3168 16304 3208 16336
rect 3240 16304 3280 16336
rect 3312 16304 3352 16336
rect 3384 16304 3424 16336
rect 3456 16304 3496 16336
rect 3528 16304 3568 16336
rect 3600 16304 3640 16336
rect 3672 16304 3712 16336
rect 3744 16304 3784 16336
rect 3816 16304 3856 16336
rect 3888 16304 4000 16336
rect 0 16264 4000 16304
rect 0 16232 112 16264
rect 144 16232 184 16264
rect 216 16232 256 16264
rect 288 16232 328 16264
rect 360 16232 400 16264
rect 432 16232 472 16264
rect 504 16232 544 16264
rect 576 16232 616 16264
rect 648 16232 688 16264
rect 720 16232 760 16264
rect 792 16232 832 16264
rect 864 16232 904 16264
rect 936 16232 976 16264
rect 1008 16232 1048 16264
rect 1080 16232 1120 16264
rect 1152 16232 1192 16264
rect 1224 16232 1264 16264
rect 1296 16232 1336 16264
rect 1368 16232 1408 16264
rect 1440 16232 1480 16264
rect 1512 16232 1552 16264
rect 1584 16232 1624 16264
rect 1656 16232 1696 16264
rect 1728 16232 1768 16264
rect 1800 16232 1840 16264
rect 1872 16232 1912 16264
rect 1944 16232 1984 16264
rect 2016 16232 2056 16264
rect 2088 16232 2128 16264
rect 2160 16232 2200 16264
rect 2232 16232 2272 16264
rect 2304 16232 2344 16264
rect 2376 16232 2416 16264
rect 2448 16232 2488 16264
rect 2520 16232 2560 16264
rect 2592 16232 2632 16264
rect 2664 16232 2704 16264
rect 2736 16232 2776 16264
rect 2808 16232 2848 16264
rect 2880 16232 2920 16264
rect 2952 16232 2992 16264
rect 3024 16232 3064 16264
rect 3096 16232 3136 16264
rect 3168 16232 3208 16264
rect 3240 16232 3280 16264
rect 3312 16232 3352 16264
rect 3384 16232 3424 16264
rect 3456 16232 3496 16264
rect 3528 16232 3568 16264
rect 3600 16232 3640 16264
rect 3672 16232 3712 16264
rect 3744 16232 3784 16264
rect 3816 16232 3856 16264
rect 3888 16232 4000 16264
rect 0 16192 4000 16232
rect 0 16160 112 16192
rect 144 16160 184 16192
rect 216 16160 256 16192
rect 288 16160 328 16192
rect 360 16160 400 16192
rect 432 16160 472 16192
rect 504 16160 544 16192
rect 576 16160 616 16192
rect 648 16160 688 16192
rect 720 16160 760 16192
rect 792 16160 832 16192
rect 864 16160 904 16192
rect 936 16160 976 16192
rect 1008 16160 1048 16192
rect 1080 16160 1120 16192
rect 1152 16160 1192 16192
rect 1224 16160 1264 16192
rect 1296 16160 1336 16192
rect 1368 16160 1408 16192
rect 1440 16160 1480 16192
rect 1512 16160 1552 16192
rect 1584 16160 1624 16192
rect 1656 16160 1696 16192
rect 1728 16160 1768 16192
rect 1800 16160 1840 16192
rect 1872 16160 1912 16192
rect 1944 16160 1984 16192
rect 2016 16160 2056 16192
rect 2088 16160 2128 16192
rect 2160 16160 2200 16192
rect 2232 16160 2272 16192
rect 2304 16160 2344 16192
rect 2376 16160 2416 16192
rect 2448 16160 2488 16192
rect 2520 16160 2560 16192
rect 2592 16160 2632 16192
rect 2664 16160 2704 16192
rect 2736 16160 2776 16192
rect 2808 16160 2848 16192
rect 2880 16160 2920 16192
rect 2952 16160 2992 16192
rect 3024 16160 3064 16192
rect 3096 16160 3136 16192
rect 3168 16160 3208 16192
rect 3240 16160 3280 16192
rect 3312 16160 3352 16192
rect 3384 16160 3424 16192
rect 3456 16160 3496 16192
rect 3528 16160 3568 16192
rect 3600 16160 3640 16192
rect 3672 16160 3712 16192
rect 3744 16160 3784 16192
rect 3816 16160 3856 16192
rect 3888 16160 4000 16192
rect 0 16120 4000 16160
rect 0 16088 112 16120
rect 144 16088 184 16120
rect 216 16088 256 16120
rect 288 16088 328 16120
rect 360 16088 400 16120
rect 432 16088 472 16120
rect 504 16088 544 16120
rect 576 16088 616 16120
rect 648 16088 688 16120
rect 720 16088 760 16120
rect 792 16088 832 16120
rect 864 16088 904 16120
rect 936 16088 976 16120
rect 1008 16088 1048 16120
rect 1080 16088 1120 16120
rect 1152 16088 1192 16120
rect 1224 16088 1264 16120
rect 1296 16088 1336 16120
rect 1368 16088 1408 16120
rect 1440 16088 1480 16120
rect 1512 16088 1552 16120
rect 1584 16088 1624 16120
rect 1656 16088 1696 16120
rect 1728 16088 1768 16120
rect 1800 16088 1840 16120
rect 1872 16088 1912 16120
rect 1944 16088 1984 16120
rect 2016 16088 2056 16120
rect 2088 16088 2128 16120
rect 2160 16088 2200 16120
rect 2232 16088 2272 16120
rect 2304 16088 2344 16120
rect 2376 16088 2416 16120
rect 2448 16088 2488 16120
rect 2520 16088 2560 16120
rect 2592 16088 2632 16120
rect 2664 16088 2704 16120
rect 2736 16088 2776 16120
rect 2808 16088 2848 16120
rect 2880 16088 2920 16120
rect 2952 16088 2992 16120
rect 3024 16088 3064 16120
rect 3096 16088 3136 16120
rect 3168 16088 3208 16120
rect 3240 16088 3280 16120
rect 3312 16088 3352 16120
rect 3384 16088 3424 16120
rect 3456 16088 3496 16120
rect 3528 16088 3568 16120
rect 3600 16088 3640 16120
rect 3672 16088 3712 16120
rect 3744 16088 3784 16120
rect 3816 16088 3856 16120
rect 3888 16088 4000 16120
rect 0 16048 4000 16088
rect 0 16016 112 16048
rect 144 16016 184 16048
rect 216 16016 256 16048
rect 288 16016 328 16048
rect 360 16016 400 16048
rect 432 16016 472 16048
rect 504 16016 544 16048
rect 576 16016 616 16048
rect 648 16016 688 16048
rect 720 16016 760 16048
rect 792 16016 832 16048
rect 864 16016 904 16048
rect 936 16016 976 16048
rect 1008 16016 1048 16048
rect 1080 16016 1120 16048
rect 1152 16016 1192 16048
rect 1224 16016 1264 16048
rect 1296 16016 1336 16048
rect 1368 16016 1408 16048
rect 1440 16016 1480 16048
rect 1512 16016 1552 16048
rect 1584 16016 1624 16048
rect 1656 16016 1696 16048
rect 1728 16016 1768 16048
rect 1800 16016 1840 16048
rect 1872 16016 1912 16048
rect 1944 16016 1984 16048
rect 2016 16016 2056 16048
rect 2088 16016 2128 16048
rect 2160 16016 2200 16048
rect 2232 16016 2272 16048
rect 2304 16016 2344 16048
rect 2376 16016 2416 16048
rect 2448 16016 2488 16048
rect 2520 16016 2560 16048
rect 2592 16016 2632 16048
rect 2664 16016 2704 16048
rect 2736 16016 2776 16048
rect 2808 16016 2848 16048
rect 2880 16016 2920 16048
rect 2952 16016 2992 16048
rect 3024 16016 3064 16048
rect 3096 16016 3136 16048
rect 3168 16016 3208 16048
rect 3240 16016 3280 16048
rect 3312 16016 3352 16048
rect 3384 16016 3424 16048
rect 3456 16016 3496 16048
rect 3528 16016 3568 16048
rect 3600 16016 3640 16048
rect 3672 16016 3712 16048
rect 3744 16016 3784 16048
rect 3816 16016 3856 16048
rect 3888 16016 4000 16048
rect 0 15976 4000 16016
rect 0 15944 112 15976
rect 144 15944 184 15976
rect 216 15944 256 15976
rect 288 15944 328 15976
rect 360 15944 400 15976
rect 432 15944 472 15976
rect 504 15944 544 15976
rect 576 15944 616 15976
rect 648 15944 688 15976
rect 720 15944 760 15976
rect 792 15944 832 15976
rect 864 15944 904 15976
rect 936 15944 976 15976
rect 1008 15944 1048 15976
rect 1080 15944 1120 15976
rect 1152 15944 1192 15976
rect 1224 15944 1264 15976
rect 1296 15944 1336 15976
rect 1368 15944 1408 15976
rect 1440 15944 1480 15976
rect 1512 15944 1552 15976
rect 1584 15944 1624 15976
rect 1656 15944 1696 15976
rect 1728 15944 1768 15976
rect 1800 15944 1840 15976
rect 1872 15944 1912 15976
rect 1944 15944 1984 15976
rect 2016 15944 2056 15976
rect 2088 15944 2128 15976
rect 2160 15944 2200 15976
rect 2232 15944 2272 15976
rect 2304 15944 2344 15976
rect 2376 15944 2416 15976
rect 2448 15944 2488 15976
rect 2520 15944 2560 15976
rect 2592 15944 2632 15976
rect 2664 15944 2704 15976
rect 2736 15944 2776 15976
rect 2808 15944 2848 15976
rect 2880 15944 2920 15976
rect 2952 15944 2992 15976
rect 3024 15944 3064 15976
rect 3096 15944 3136 15976
rect 3168 15944 3208 15976
rect 3240 15944 3280 15976
rect 3312 15944 3352 15976
rect 3384 15944 3424 15976
rect 3456 15944 3496 15976
rect 3528 15944 3568 15976
rect 3600 15944 3640 15976
rect 3672 15944 3712 15976
rect 3744 15944 3784 15976
rect 3816 15944 3856 15976
rect 3888 15944 4000 15976
rect 0 15904 4000 15944
rect 0 15872 112 15904
rect 144 15872 184 15904
rect 216 15872 256 15904
rect 288 15872 328 15904
rect 360 15872 400 15904
rect 432 15872 472 15904
rect 504 15872 544 15904
rect 576 15872 616 15904
rect 648 15872 688 15904
rect 720 15872 760 15904
rect 792 15872 832 15904
rect 864 15872 904 15904
rect 936 15872 976 15904
rect 1008 15872 1048 15904
rect 1080 15872 1120 15904
rect 1152 15872 1192 15904
rect 1224 15872 1264 15904
rect 1296 15872 1336 15904
rect 1368 15872 1408 15904
rect 1440 15872 1480 15904
rect 1512 15872 1552 15904
rect 1584 15872 1624 15904
rect 1656 15872 1696 15904
rect 1728 15872 1768 15904
rect 1800 15872 1840 15904
rect 1872 15872 1912 15904
rect 1944 15872 1984 15904
rect 2016 15872 2056 15904
rect 2088 15872 2128 15904
rect 2160 15872 2200 15904
rect 2232 15872 2272 15904
rect 2304 15872 2344 15904
rect 2376 15872 2416 15904
rect 2448 15872 2488 15904
rect 2520 15872 2560 15904
rect 2592 15872 2632 15904
rect 2664 15872 2704 15904
rect 2736 15872 2776 15904
rect 2808 15872 2848 15904
rect 2880 15872 2920 15904
rect 2952 15872 2992 15904
rect 3024 15872 3064 15904
rect 3096 15872 3136 15904
rect 3168 15872 3208 15904
rect 3240 15872 3280 15904
rect 3312 15872 3352 15904
rect 3384 15872 3424 15904
rect 3456 15872 3496 15904
rect 3528 15872 3568 15904
rect 3600 15872 3640 15904
rect 3672 15872 3712 15904
rect 3744 15872 3784 15904
rect 3816 15872 3856 15904
rect 3888 15872 4000 15904
rect 0 15832 4000 15872
rect 0 15800 112 15832
rect 144 15800 184 15832
rect 216 15800 256 15832
rect 288 15800 328 15832
rect 360 15800 400 15832
rect 432 15800 472 15832
rect 504 15800 544 15832
rect 576 15800 616 15832
rect 648 15800 688 15832
rect 720 15800 760 15832
rect 792 15800 832 15832
rect 864 15800 904 15832
rect 936 15800 976 15832
rect 1008 15800 1048 15832
rect 1080 15800 1120 15832
rect 1152 15800 1192 15832
rect 1224 15800 1264 15832
rect 1296 15800 1336 15832
rect 1368 15800 1408 15832
rect 1440 15800 1480 15832
rect 1512 15800 1552 15832
rect 1584 15800 1624 15832
rect 1656 15800 1696 15832
rect 1728 15800 1768 15832
rect 1800 15800 1840 15832
rect 1872 15800 1912 15832
rect 1944 15800 1984 15832
rect 2016 15800 2056 15832
rect 2088 15800 2128 15832
rect 2160 15800 2200 15832
rect 2232 15800 2272 15832
rect 2304 15800 2344 15832
rect 2376 15800 2416 15832
rect 2448 15800 2488 15832
rect 2520 15800 2560 15832
rect 2592 15800 2632 15832
rect 2664 15800 2704 15832
rect 2736 15800 2776 15832
rect 2808 15800 2848 15832
rect 2880 15800 2920 15832
rect 2952 15800 2992 15832
rect 3024 15800 3064 15832
rect 3096 15800 3136 15832
rect 3168 15800 3208 15832
rect 3240 15800 3280 15832
rect 3312 15800 3352 15832
rect 3384 15800 3424 15832
rect 3456 15800 3496 15832
rect 3528 15800 3568 15832
rect 3600 15800 3640 15832
rect 3672 15800 3712 15832
rect 3744 15800 3784 15832
rect 3816 15800 3856 15832
rect 3888 15800 4000 15832
rect 0 15760 4000 15800
rect 0 15728 112 15760
rect 144 15728 184 15760
rect 216 15728 256 15760
rect 288 15728 328 15760
rect 360 15728 400 15760
rect 432 15728 472 15760
rect 504 15728 544 15760
rect 576 15728 616 15760
rect 648 15728 688 15760
rect 720 15728 760 15760
rect 792 15728 832 15760
rect 864 15728 904 15760
rect 936 15728 976 15760
rect 1008 15728 1048 15760
rect 1080 15728 1120 15760
rect 1152 15728 1192 15760
rect 1224 15728 1264 15760
rect 1296 15728 1336 15760
rect 1368 15728 1408 15760
rect 1440 15728 1480 15760
rect 1512 15728 1552 15760
rect 1584 15728 1624 15760
rect 1656 15728 1696 15760
rect 1728 15728 1768 15760
rect 1800 15728 1840 15760
rect 1872 15728 1912 15760
rect 1944 15728 1984 15760
rect 2016 15728 2056 15760
rect 2088 15728 2128 15760
rect 2160 15728 2200 15760
rect 2232 15728 2272 15760
rect 2304 15728 2344 15760
rect 2376 15728 2416 15760
rect 2448 15728 2488 15760
rect 2520 15728 2560 15760
rect 2592 15728 2632 15760
rect 2664 15728 2704 15760
rect 2736 15728 2776 15760
rect 2808 15728 2848 15760
rect 2880 15728 2920 15760
rect 2952 15728 2992 15760
rect 3024 15728 3064 15760
rect 3096 15728 3136 15760
rect 3168 15728 3208 15760
rect 3240 15728 3280 15760
rect 3312 15728 3352 15760
rect 3384 15728 3424 15760
rect 3456 15728 3496 15760
rect 3528 15728 3568 15760
rect 3600 15728 3640 15760
rect 3672 15728 3712 15760
rect 3744 15728 3784 15760
rect 3816 15728 3856 15760
rect 3888 15728 4000 15760
rect 0 15688 4000 15728
rect 0 15656 112 15688
rect 144 15656 184 15688
rect 216 15656 256 15688
rect 288 15656 328 15688
rect 360 15656 400 15688
rect 432 15656 472 15688
rect 504 15656 544 15688
rect 576 15656 616 15688
rect 648 15656 688 15688
rect 720 15656 760 15688
rect 792 15656 832 15688
rect 864 15656 904 15688
rect 936 15656 976 15688
rect 1008 15656 1048 15688
rect 1080 15656 1120 15688
rect 1152 15656 1192 15688
rect 1224 15656 1264 15688
rect 1296 15656 1336 15688
rect 1368 15656 1408 15688
rect 1440 15656 1480 15688
rect 1512 15656 1552 15688
rect 1584 15656 1624 15688
rect 1656 15656 1696 15688
rect 1728 15656 1768 15688
rect 1800 15656 1840 15688
rect 1872 15656 1912 15688
rect 1944 15656 1984 15688
rect 2016 15656 2056 15688
rect 2088 15656 2128 15688
rect 2160 15656 2200 15688
rect 2232 15656 2272 15688
rect 2304 15656 2344 15688
rect 2376 15656 2416 15688
rect 2448 15656 2488 15688
rect 2520 15656 2560 15688
rect 2592 15656 2632 15688
rect 2664 15656 2704 15688
rect 2736 15656 2776 15688
rect 2808 15656 2848 15688
rect 2880 15656 2920 15688
rect 2952 15656 2992 15688
rect 3024 15656 3064 15688
rect 3096 15656 3136 15688
rect 3168 15656 3208 15688
rect 3240 15656 3280 15688
rect 3312 15656 3352 15688
rect 3384 15656 3424 15688
rect 3456 15656 3496 15688
rect 3528 15656 3568 15688
rect 3600 15656 3640 15688
rect 3672 15656 3712 15688
rect 3744 15656 3784 15688
rect 3816 15656 3856 15688
rect 3888 15656 4000 15688
rect 0 15616 4000 15656
rect 0 15584 112 15616
rect 144 15584 184 15616
rect 216 15584 256 15616
rect 288 15584 328 15616
rect 360 15584 400 15616
rect 432 15584 472 15616
rect 504 15584 544 15616
rect 576 15584 616 15616
rect 648 15584 688 15616
rect 720 15584 760 15616
rect 792 15584 832 15616
rect 864 15584 904 15616
rect 936 15584 976 15616
rect 1008 15584 1048 15616
rect 1080 15584 1120 15616
rect 1152 15584 1192 15616
rect 1224 15584 1264 15616
rect 1296 15584 1336 15616
rect 1368 15584 1408 15616
rect 1440 15584 1480 15616
rect 1512 15584 1552 15616
rect 1584 15584 1624 15616
rect 1656 15584 1696 15616
rect 1728 15584 1768 15616
rect 1800 15584 1840 15616
rect 1872 15584 1912 15616
rect 1944 15584 1984 15616
rect 2016 15584 2056 15616
rect 2088 15584 2128 15616
rect 2160 15584 2200 15616
rect 2232 15584 2272 15616
rect 2304 15584 2344 15616
rect 2376 15584 2416 15616
rect 2448 15584 2488 15616
rect 2520 15584 2560 15616
rect 2592 15584 2632 15616
rect 2664 15584 2704 15616
rect 2736 15584 2776 15616
rect 2808 15584 2848 15616
rect 2880 15584 2920 15616
rect 2952 15584 2992 15616
rect 3024 15584 3064 15616
rect 3096 15584 3136 15616
rect 3168 15584 3208 15616
rect 3240 15584 3280 15616
rect 3312 15584 3352 15616
rect 3384 15584 3424 15616
rect 3456 15584 3496 15616
rect 3528 15584 3568 15616
rect 3600 15584 3640 15616
rect 3672 15584 3712 15616
rect 3744 15584 3784 15616
rect 3816 15584 3856 15616
rect 3888 15584 4000 15616
rect 0 15544 4000 15584
rect 0 15512 112 15544
rect 144 15512 184 15544
rect 216 15512 256 15544
rect 288 15512 328 15544
rect 360 15512 400 15544
rect 432 15512 472 15544
rect 504 15512 544 15544
rect 576 15512 616 15544
rect 648 15512 688 15544
rect 720 15512 760 15544
rect 792 15512 832 15544
rect 864 15512 904 15544
rect 936 15512 976 15544
rect 1008 15512 1048 15544
rect 1080 15512 1120 15544
rect 1152 15512 1192 15544
rect 1224 15512 1264 15544
rect 1296 15512 1336 15544
rect 1368 15512 1408 15544
rect 1440 15512 1480 15544
rect 1512 15512 1552 15544
rect 1584 15512 1624 15544
rect 1656 15512 1696 15544
rect 1728 15512 1768 15544
rect 1800 15512 1840 15544
rect 1872 15512 1912 15544
rect 1944 15512 1984 15544
rect 2016 15512 2056 15544
rect 2088 15512 2128 15544
rect 2160 15512 2200 15544
rect 2232 15512 2272 15544
rect 2304 15512 2344 15544
rect 2376 15512 2416 15544
rect 2448 15512 2488 15544
rect 2520 15512 2560 15544
rect 2592 15512 2632 15544
rect 2664 15512 2704 15544
rect 2736 15512 2776 15544
rect 2808 15512 2848 15544
rect 2880 15512 2920 15544
rect 2952 15512 2992 15544
rect 3024 15512 3064 15544
rect 3096 15512 3136 15544
rect 3168 15512 3208 15544
rect 3240 15512 3280 15544
rect 3312 15512 3352 15544
rect 3384 15512 3424 15544
rect 3456 15512 3496 15544
rect 3528 15512 3568 15544
rect 3600 15512 3640 15544
rect 3672 15512 3712 15544
rect 3744 15512 3784 15544
rect 3816 15512 3856 15544
rect 3888 15512 4000 15544
rect 0 15472 4000 15512
rect 0 15440 112 15472
rect 144 15440 184 15472
rect 216 15440 256 15472
rect 288 15440 328 15472
rect 360 15440 400 15472
rect 432 15440 472 15472
rect 504 15440 544 15472
rect 576 15440 616 15472
rect 648 15440 688 15472
rect 720 15440 760 15472
rect 792 15440 832 15472
rect 864 15440 904 15472
rect 936 15440 976 15472
rect 1008 15440 1048 15472
rect 1080 15440 1120 15472
rect 1152 15440 1192 15472
rect 1224 15440 1264 15472
rect 1296 15440 1336 15472
rect 1368 15440 1408 15472
rect 1440 15440 1480 15472
rect 1512 15440 1552 15472
rect 1584 15440 1624 15472
rect 1656 15440 1696 15472
rect 1728 15440 1768 15472
rect 1800 15440 1840 15472
rect 1872 15440 1912 15472
rect 1944 15440 1984 15472
rect 2016 15440 2056 15472
rect 2088 15440 2128 15472
rect 2160 15440 2200 15472
rect 2232 15440 2272 15472
rect 2304 15440 2344 15472
rect 2376 15440 2416 15472
rect 2448 15440 2488 15472
rect 2520 15440 2560 15472
rect 2592 15440 2632 15472
rect 2664 15440 2704 15472
rect 2736 15440 2776 15472
rect 2808 15440 2848 15472
rect 2880 15440 2920 15472
rect 2952 15440 2992 15472
rect 3024 15440 3064 15472
rect 3096 15440 3136 15472
rect 3168 15440 3208 15472
rect 3240 15440 3280 15472
rect 3312 15440 3352 15472
rect 3384 15440 3424 15472
rect 3456 15440 3496 15472
rect 3528 15440 3568 15472
rect 3600 15440 3640 15472
rect 3672 15440 3712 15472
rect 3744 15440 3784 15472
rect 3816 15440 3856 15472
rect 3888 15440 4000 15472
rect 0 15400 4000 15440
rect 0 15368 112 15400
rect 144 15368 184 15400
rect 216 15368 256 15400
rect 288 15368 328 15400
rect 360 15368 400 15400
rect 432 15368 472 15400
rect 504 15368 544 15400
rect 576 15368 616 15400
rect 648 15368 688 15400
rect 720 15368 760 15400
rect 792 15368 832 15400
rect 864 15368 904 15400
rect 936 15368 976 15400
rect 1008 15368 1048 15400
rect 1080 15368 1120 15400
rect 1152 15368 1192 15400
rect 1224 15368 1264 15400
rect 1296 15368 1336 15400
rect 1368 15368 1408 15400
rect 1440 15368 1480 15400
rect 1512 15368 1552 15400
rect 1584 15368 1624 15400
rect 1656 15368 1696 15400
rect 1728 15368 1768 15400
rect 1800 15368 1840 15400
rect 1872 15368 1912 15400
rect 1944 15368 1984 15400
rect 2016 15368 2056 15400
rect 2088 15368 2128 15400
rect 2160 15368 2200 15400
rect 2232 15368 2272 15400
rect 2304 15368 2344 15400
rect 2376 15368 2416 15400
rect 2448 15368 2488 15400
rect 2520 15368 2560 15400
rect 2592 15368 2632 15400
rect 2664 15368 2704 15400
rect 2736 15368 2776 15400
rect 2808 15368 2848 15400
rect 2880 15368 2920 15400
rect 2952 15368 2992 15400
rect 3024 15368 3064 15400
rect 3096 15368 3136 15400
rect 3168 15368 3208 15400
rect 3240 15368 3280 15400
rect 3312 15368 3352 15400
rect 3384 15368 3424 15400
rect 3456 15368 3496 15400
rect 3528 15368 3568 15400
rect 3600 15368 3640 15400
rect 3672 15368 3712 15400
rect 3744 15368 3784 15400
rect 3816 15368 3856 15400
rect 3888 15368 4000 15400
rect 0 15328 4000 15368
rect 0 15296 112 15328
rect 144 15296 184 15328
rect 216 15296 256 15328
rect 288 15296 328 15328
rect 360 15296 400 15328
rect 432 15296 472 15328
rect 504 15296 544 15328
rect 576 15296 616 15328
rect 648 15296 688 15328
rect 720 15296 760 15328
rect 792 15296 832 15328
rect 864 15296 904 15328
rect 936 15296 976 15328
rect 1008 15296 1048 15328
rect 1080 15296 1120 15328
rect 1152 15296 1192 15328
rect 1224 15296 1264 15328
rect 1296 15296 1336 15328
rect 1368 15296 1408 15328
rect 1440 15296 1480 15328
rect 1512 15296 1552 15328
rect 1584 15296 1624 15328
rect 1656 15296 1696 15328
rect 1728 15296 1768 15328
rect 1800 15296 1840 15328
rect 1872 15296 1912 15328
rect 1944 15296 1984 15328
rect 2016 15296 2056 15328
rect 2088 15296 2128 15328
rect 2160 15296 2200 15328
rect 2232 15296 2272 15328
rect 2304 15296 2344 15328
rect 2376 15296 2416 15328
rect 2448 15296 2488 15328
rect 2520 15296 2560 15328
rect 2592 15296 2632 15328
rect 2664 15296 2704 15328
rect 2736 15296 2776 15328
rect 2808 15296 2848 15328
rect 2880 15296 2920 15328
rect 2952 15296 2992 15328
rect 3024 15296 3064 15328
rect 3096 15296 3136 15328
rect 3168 15296 3208 15328
rect 3240 15296 3280 15328
rect 3312 15296 3352 15328
rect 3384 15296 3424 15328
rect 3456 15296 3496 15328
rect 3528 15296 3568 15328
rect 3600 15296 3640 15328
rect 3672 15296 3712 15328
rect 3744 15296 3784 15328
rect 3816 15296 3856 15328
rect 3888 15296 4000 15328
rect 0 15256 4000 15296
rect 0 15224 112 15256
rect 144 15224 184 15256
rect 216 15224 256 15256
rect 288 15224 328 15256
rect 360 15224 400 15256
rect 432 15224 472 15256
rect 504 15224 544 15256
rect 576 15224 616 15256
rect 648 15224 688 15256
rect 720 15224 760 15256
rect 792 15224 832 15256
rect 864 15224 904 15256
rect 936 15224 976 15256
rect 1008 15224 1048 15256
rect 1080 15224 1120 15256
rect 1152 15224 1192 15256
rect 1224 15224 1264 15256
rect 1296 15224 1336 15256
rect 1368 15224 1408 15256
rect 1440 15224 1480 15256
rect 1512 15224 1552 15256
rect 1584 15224 1624 15256
rect 1656 15224 1696 15256
rect 1728 15224 1768 15256
rect 1800 15224 1840 15256
rect 1872 15224 1912 15256
rect 1944 15224 1984 15256
rect 2016 15224 2056 15256
rect 2088 15224 2128 15256
rect 2160 15224 2200 15256
rect 2232 15224 2272 15256
rect 2304 15224 2344 15256
rect 2376 15224 2416 15256
rect 2448 15224 2488 15256
rect 2520 15224 2560 15256
rect 2592 15224 2632 15256
rect 2664 15224 2704 15256
rect 2736 15224 2776 15256
rect 2808 15224 2848 15256
rect 2880 15224 2920 15256
rect 2952 15224 2992 15256
rect 3024 15224 3064 15256
rect 3096 15224 3136 15256
rect 3168 15224 3208 15256
rect 3240 15224 3280 15256
rect 3312 15224 3352 15256
rect 3384 15224 3424 15256
rect 3456 15224 3496 15256
rect 3528 15224 3568 15256
rect 3600 15224 3640 15256
rect 3672 15224 3712 15256
rect 3744 15224 3784 15256
rect 3816 15224 3856 15256
rect 3888 15224 4000 15256
rect 0 15184 4000 15224
rect 0 15152 112 15184
rect 144 15152 184 15184
rect 216 15152 256 15184
rect 288 15152 328 15184
rect 360 15152 400 15184
rect 432 15152 472 15184
rect 504 15152 544 15184
rect 576 15152 616 15184
rect 648 15152 688 15184
rect 720 15152 760 15184
rect 792 15152 832 15184
rect 864 15152 904 15184
rect 936 15152 976 15184
rect 1008 15152 1048 15184
rect 1080 15152 1120 15184
rect 1152 15152 1192 15184
rect 1224 15152 1264 15184
rect 1296 15152 1336 15184
rect 1368 15152 1408 15184
rect 1440 15152 1480 15184
rect 1512 15152 1552 15184
rect 1584 15152 1624 15184
rect 1656 15152 1696 15184
rect 1728 15152 1768 15184
rect 1800 15152 1840 15184
rect 1872 15152 1912 15184
rect 1944 15152 1984 15184
rect 2016 15152 2056 15184
rect 2088 15152 2128 15184
rect 2160 15152 2200 15184
rect 2232 15152 2272 15184
rect 2304 15152 2344 15184
rect 2376 15152 2416 15184
rect 2448 15152 2488 15184
rect 2520 15152 2560 15184
rect 2592 15152 2632 15184
rect 2664 15152 2704 15184
rect 2736 15152 2776 15184
rect 2808 15152 2848 15184
rect 2880 15152 2920 15184
rect 2952 15152 2992 15184
rect 3024 15152 3064 15184
rect 3096 15152 3136 15184
rect 3168 15152 3208 15184
rect 3240 15152 3280 15184
rect 3312 15152 3352 15184
rect 3384 15152 3424 15184
rect 3456 15152 3496 15184
rect 3528 15152 3568 15184
rect 3600 15152 3640 15184
rect 3672 15152 3712 15184
rect 3744 15152 3784 15184
rect 3816 15152 3856 15184
rect 3888 15152 4000 15184
rect 0 15112 4000 15152
rect 0 15080 112 15112
rect 144 15080 184 15112
rect 216 15080 256 15112
rect 288 15080 328 15112
rect 360 15080 400 15112
rect 432 15080 472 15112
rect 504 15080 544 15112
rect 576 15080 616 15112
rect 648 15080 688 15112
rect 720 15080 760 15112
rect 792 15080 832 15112
rect 864 15080 904 15112
rect 936 15080 976 15112
rect 1008 15080 1048 15112
rect 1080 15080 1120 15112
rect 1152 15080 1192 15112
rect 1224 15080 1264 15112
rect 1296 15080 1336 15112
rect 1368 15080 1408 15112
rect 1440 15080 1480 15112
rect 1512 15080 1552 15112
rect 1584 15080 1624 15112
rect 1656 15080 1696 15112
rect 1728 15080 1768 15112
rect 1800 15080 1840 15112
rect 1872 15080 1912 15112
rect 1944 15080 1984 15112
rect 2016 15080 2056 15112
rect 2088 15080 2128 15112
rect 2160 15080 2200 15112
rect 2232 15080 2272 15112
rect 2304 15080 2344 15112
rect 2376 15080 2416 15112
rect 2448 15080 2488 15112
rect 2520 15080 2560 15112
rect 2592 15080 2632 15112
rect 2664 15080 2704 15112
rect 2736 15080 2776 15112
rect 2808 15080 2848 15112
rect 2880 15080 2920 15112
rect 2952 15080 2992 15112
rect 3024 15080 3064 15112
rect 3096 15080 3136 15112
rect 3168 15080 3208 15112
rect 3240 15080 3280 15112
rect 3312 15080 3352 15112
rect 3384 15080 3424 15112
rect 3456 15080 3496 15112
rect 3528 15080 3568 15112
rect 3600 15080 3640 15112
rect 3672 15080 3712 15112
rect 3744 15080 3784 15112
rect 3816 15080 3856 15112
rect 3888 15080 4000 15112
rect 0 15040 4000 15080
rect 0 15008 112 15040
rect 144 15008 184 15040
rect 216 15008 256 15040
rect 288 15008 328 15040
rect 360 15008 400 15040
rect 432 15008 472 15040
rect 504 15008 544 15040
rect 576 15008 616 15040
rect 648 15008 688 15040
rect 720 15008 760 15040
rect 792 15008 832 15040
rect 864 15008 904 15040
rect 936 15008 976 15040
rect 1008 15008 1048 15040
rect 1080 15008 1120 15040
rect 1152 15008 1192 15040
rect 1224 15008 1264 15040
rect 1296 15008 1336 15040
rect 1368 15008 1408 15040
rect 1440 15008 1480 15040
rect 1512 15008 1552 15040
rect 1584 15008 1624 15040
rect 1656 15008 1696 15040
rect 1728 15008 1768 15040
rect 1800 15008 1840 15040
rect 1872 15008 1912 15040
rect 1944 15008 1984 15040
rect 2016 15008 2056 15040
rect 2088 15008 2128 15040
rect 2160 15008 2200 15040
rect 2232 15008 2272 15040
rect 2304 15008 2344 15040
rect 2376 15008 2416 15040
rect 2448 15008 2488 15040
rect 2520 15008 2560 15040
rect 2592 15008 2632 15040
rect 2664 15008 2704 15040
rect 2736 15008 2776 15040
rect 2808 15008 2848 15040
rect 2880 15008 2920 15040
rect 2952 15008 2992 15040
rect 3024 15008 3064 15040
rect 3096 15008 3136 15040
rect 3168 15008 3208 15040
rect 3240 15008 3280 15040
rect 3312 15008 3352 15040
rect 3384 15008 3424 15040
rect 3456 15008 3496 15040
rect 3528 15008 3568 15040
rect 3600 15008 3640 15040
rect 3672 15008 3712 15040
rect 3744 15008 3784 15040
rect 3816 15008 3856 15040
rect 3888 15008 4000 15040
rect 0 14968 4000 15008
rect 0 14936 112 14968
rect 144 14936 184 14968
rect 216 14936 256 14968
rect 288 14936 328 14968
rect 360 14936 400 14968
rect 432 14936 472 14968
rect 504 14936 544 14968
rect 576 14936 616 14968
rect 648 14936 688 14968
rect 720 14936 760 14968
rect 792 14936 832 14968
rect 864 14936 904 14968
rect 936 14936 976 14968
rect 1008 14936 1048 14968
rect 1080 14936 1120 14968
rect 1152 14936 1192 14968
rect 1224 14936 1264 14968
rect 1296 14936 1336 14968
rect 1368 14936 1408 14968
rect 1440 14936 1480 14968
rect 1512 14936 1552 14968
rect 1584 14936 1624 14968
rect 1656 14936 1696 14968
rect 1728 14936 1768 14968
rect 1800 14936 1840 14968
rect 1872 14936 1912 14968
rect 1944 14936 1984 14968
rect 2016 14936 2056 14968
rect 2088 14936 2128 14968
rect 2160 14936 2200 14968
rect 2232 14936 2272 14968
rect 2304 14936 2344 14968
rect 2376 14936 2416 14968
rect 2448 14936 2488 14968
rect 2520 14936 2560 14968
rect 2592 14936 2632 14968
rect 2664 14936 2704 14968
rect 2736 14936 2776 14968
rect 2808 14936 2848 14968
rect 2880 14936 2920 14968
rect 2952 14936 2992 14968
rect 3024 14936 3064 14968
rect 3096 14936 3136 14968
rect 3168 14936 3208 14968
rect 3240 14936 3280 14968
rect 3312 14936 3352 14968
rect 3384 14936 3424 14968
rect 3456 14936 3496 14968
rect 3528 14936 3568 14968
rect 3600 14936 3640 14968
rect 3672 14936 3712 14968
rect 3744 14936 3784 14968
rect 3816 14936 3856 14968
rect 3888 14936 4000 14968
rect 0 14896 4000 14936
rect 0 14864 112 14896
rect 144 14864 184 14896
rect 216 14864 256 14896
rect 288 14864 328 14896
rect 360 14864 400 14896
rect 432 14864 472 14896
rect 504 14864 544 14896
rect 576 14864 616 14896
rect 648 14864 688 14896
rect 720 14864 760 14896
rect 792 14864 832 14896
rect 864 14864 904 14896
rect 936 14864 976 14896
rect 1008 14864 1048 14896
rect 1080 14864 1120 14896
rect 1152 14864 1192 14896
rect 1224 14864 1264 14896
rect 1296 14864 1336 14896
rect 1368 14864 1408 14896
rect 1440 14864 1480 14896
rect 1512 14864 1552 14896
rect 1584 14864 1624 14896
rect 1656 14864 1696 14896
rect 1728 14864 1768 14896
rect 1800 14864 1840 14896
rect 1872 14864 1912 14896
rect 1944 14864 1984 14896
rect 2016 14864 2056 14896
rect 2088 14864 2128 14896
rect 2160 14864 2200 14896
rect 2232 14864 2272 14896
rect 2304 14864 2344 14896
rect 2376 14864 2416 14896
rect 2448 14864 2488 14896
rect 2520 14864 2560 14896
rect 2592 14864 2632 14896
rect 2664 14864 2704 14896
rect 2736 14864 2776 14896
rect 2808 14864 2848 14896
rect 2880 14864 2920 14896
rect 2952 14864 2992 14896
rect 3024 14864 3064 14896
rect 3096 14864 3136 14896
rect 3168 14864 3208 14896
rect 3240 14864 3280 14896
rect 3312 14864 3352 14896
rect 3384 14864 3424 14896
rect 3456 14864 3496 14896
rect 3528 14864 3568 14896
rect 3600 14864 3640 14896
rect 3672 14864 3712 14896
rect 3744 14864 3784 14896
rect 3816 14864 3856 14896
rect 3888 14864 4000 14896
rect 0 14824 4000 14864
rect 0 14792 112 14824
rect 144 14792 184 14824
rect 216 14792 256 14824
rect 288 14792 328 14824
rect 360 14792 400 14824
rect 432 14792 472 14824
rect 504 14792 544 14824
rect 576 14792 616 14824
rect 648 14792 688 14824
rect 720 14792 760 14824
rect 792 14792 832 14824
rect 864 14792 904 14824
rect 936 14792 976 14824
rect 1008 14792 1048 14824
rect 1080 14792 1120 14824
rect 1152 14792 1192 14824
rect 1224 14792 1264 14824
rect 1296 14792 1336 14824
rect 1368 14792 1408 14824
rect 1440 14792 1480 14824
rect 1512 14792 1552 14824
rect 1584 14792 1624 14824
rect 1656 14792 1696 14824
rect 1728 14792 1768 14824
rect 1800 14792 1840 14824
rect 1872 14792 1912 14824
rect 1944 14792 1984 14824
rect 2016 14792 2056 14824
rect 2088 14792 2128 14824
rect 2160 14792 2200 14824
rect 2232 14792 2272 14824
rect 2304 14792 2344 14824
rect 2376 14792 2416 14824
rect 2448 14792 2488 14824
rect 2520 14792 2560 14824
rect 2592 14792 2632 14824
rect 2664 14792 2704 14824
rect 2736 14792 2776 14824
rect 2808 14792 2848 14824
rect 2880 14792 2920 14824
rect 2952 14792 2992 14824
rect 3024 14792 3064 14824
rect 3096 14792 3136 14824
rect 3168 14792 3208 14824
rect 3240 14792 3280 14824
rect 3312 14792 3352 14824
rect 3384 14792 3424 14824
rect 3456 14792 3496 14824
rect 3528 14792 3568 14824
rect 3600 14792 3640 14824
rect 3672 14792 3712 14824
rect 3744 14792 3784 14824
rect 3816 14792 3856 14824
rect 3888 14792 4000 14824
rect 0 14752 4000 14792
rect 0 14720 112 14752
rect 144 14720 184 14752
rect 216 14720 256 14752
rect 288 14720 328 14752
rect 360 14720 400 14752
rect 432 14720 472 14752
rect 504 14720 544 14752
rect 576 14720 616 14752
rect 648 14720 688 14752
rect 720 14720 760 14752
rect 792 14720 832 14752
rect 864 14720 904 14752
rect 936 14720 976 14752
rect 1008 14720 1048 14752
rect 1080 14720 1120 14752
rect 1152 14720 1192 14752
rect 1224 14720 1264 14752
rect 1296 14720 1336 14752
rect 1368 14720 1408 14752
rect 1440 14720 1480 14752
rect 1512 14720 1552 14752
rect 1584 14720 1624 14752
rect 1656 14720 1696 14752
rect 1728 14720 1768 14752
rect 1800 14720 1840 14752
rect 1872 14720 1912 14752
rect 1944 14720 1984 14752
rect 2016 14720 2056 14752
rect 2088 14720 2128 14752
rect 2160 14720 2200 14752
rect 2232 14720 2272 14752
rect 2304 14720 2344 14752
rect 2376 14720 2416 14752
rect 2448 14720 2488 14752
rect 2520 14720 2560 14752
rect 2592 14720 2632 14752
rect 2664 14720 2704 14752
rect 2736 14720 2776 14752
rect 2808 14720 2848 14752
rect 2880 14720 2920 14752
rect 2952 14720 2992 14752
rect 3024 14720 3064 14752
rect 3096 14720 3136 14752
rect 3168 14720 3208 14752
rect 3240 14720 3280 14752
rect 3312 14720 3352 14752
rect 3384 14720 3424 14752
rect 3456 14720 3496 14752
rect 3528 14720 3568 14752
rect 3600 14720 3640 14752
rect 3672 14720 3712 14752
rect 3744 14720 3784 14752
rect 3816 14720 3856 14752
rect 3888 14720 4000 14752
rect 0 14680 4000 14720
rect 0 14648 112 14680
rect 144 14648 184 14680
rect 216 14648 256 14680
rect 288 14648 328 14680
rect 360 14648 400 14680
rect 432 14648 472 14680
rect 504 14648 544 14680
rect 576 14648 616 14680
rect 648 14648 688 14680
rect 720 14648 760 14680
rect 792 14648 832 14680
rect 864 14648 904 14680
rect 936 14648 976 14680
rect 1008 14648 1048 14680
rect 1080 14648 1120 14680
rect 1152 14648 1192 14680
rect 1224 14648 1264 14680
rect 1296 14648 1336 14680
rect 1368 14648 1408 14680
rect 1440 14648 1480 14680
rect 1512 14648 1552 14680
rect 1584 14648 1624 14680
rect 1656 14648 1696 14680
rect 1728 14648 1768 14680
rect 1800 14648 1840 14680
rect 1872 14648 1912 14680
rect 1944 14648 1984 14680
rect 2016 14648 2056 14680
rect 2088 14648 2128 14680
rect 2160 14648 2200 14680
rect 2232 14648 2272 14680
rect 2304 14648 2344 14680
rect 2376 14648 2416 14680
rect 2448 14648 2488 14680
rect 2520 14648 2560 14680
rect 2592 14648 2632 14680
rect 2664 14648 2704 14680
rect 2736 14648 2776 14680
rect 2808 14648 2848 14680
rect 2880 14648 2920 14680
rect 2952 14648 2992 14680
rect 3024 14648 3064 14680
rect 3096 14648 3136 14680
rect 3168 14648 3208 14680
rect 3240 14648 3280 14680
rect 3312 14648 3352 14680
rect 3384 14648 3424 14680
rect 3456 14648 3496 14680
rect 3528 14648 3568 14680
rect 3600 14648 3640 14680
rect 3672 14648 3712 14680
rect 3744 14648 3784 14680
rect 3816 14648 3856 14680
rect 3888 14648 4000 14680
rect 0 14608 4000 14648
rect 0 14576 112 14608
rect 144 14576 184 14608
rect 216 14576 256 14608
rect 288 14576 328 14608
rect 360 14576 400 14608
rect 432 14576 472 14608
rect 504 14576 544 14608
rect 576 14576 616 14608
rect 648 14576 688 14608
rect 720 14576 760 14608
rect 792 14576 832 14608
rect 864 14576 904 14608
rect 936 14576 976 14608
rect 1008 14576 1048 14608
rect 1080 14576 1120 14608
rect 1152 14576 1192 14608
rect 1224 14576 1264 14608
rect 1296 14576 1336 14608
rect 1368 14576 1408 14608
rect 1440 14576 1480 14608
rect 1512 14576 1552 14608
rect 1584 14576 1624 14608
rect 1656 14576 1696 14608
rect 1728 14576 1768 14608
rect 1800 14576 1840 14608
rect 1872 14576 1912 14608
rect 1944 14576 1984 14608
rect 2016 14576 2056 14608
rect 2088 14576 2128 14608
rect 2160 14576 2200 14608
rect 2232 14576 2272 14608
rect 2304 14576 2344 14608
rect 2376 14576 2416 14608
rect 2448 14576 2488 14608
rect 2520 14576 2560 14608
rect 2592 14576 2632 14608
rect 2664 14576 2704 14608
rect 2736 14576 2776 14608
rect 2808 14576 2848 14608
rect 2880 14576 2920 14608
rect 2952 14576 2992 14608
rect 3024 14576 3064 14608
rect 3096 14576 3136 14608
rect 3168 14576 3208 14608
rect 3240 14576 3280 14608
rect 3312 14576 3352 14608
rect 3384 14576 3424 14608
rect 3456 14576 3496 14608
rect 3528 14576 3568 14608
rect 3600 14576 3640 14608
rect 3672 14576 3712 14608
rect 3744 14576 3784 14608
rect 3816 14576 3856 14608
rect 3888 14576 4000 14608
rect 0 14536 4000 14576
rect 0 14504 112 14536
rect 144 14504 184 14536
rect 216 14504 256 14536
rect 288 14504 328 14536
rect 360 14504 400 14536
rect 432 14504 472 14536
rect 504 14504 544 14536
rect 576 14504 616 14536
rect 648 14504 688 14536
rect 720 14504 760 14536
rect 792 14504 832 14536
rect 864 14504 904 14536
rect 936 14504 976 14536
rect 1008 14504 1048 14536
rect 1080 14504 1120 14536
rect 1152 14504 1192 14536
rect 1224 14504 1264 14536
rect 1296 14504 1336 14536
rect 1368 14504 1408 14536
rect 1440 14504 1480 14536
rect 1512 14504 1552 14536
rect 1584 14504 1624 14536
rect 1656 14504 1696 14536
rect 1728 14504 1768 14536
rect 1800 14504 1840 14536
rect 1872 14504 1912 14536
rect 1944 14504 1984 14536
rect 2016 14504 2056 14536
rect 2088 14504 2128 14536
rect 2160 14504 2200 14536
rect 2232 14504 2272 14536
rect 2304 14504 2344 14536
rect 2376 14504 2416 14536
rect 2448 14504 2488 14536
rect 2520 14504 2560 14536
rect 2592 14504 2632 14536
rect 2664 14504 2704 14536
rect 2736 14504 2776 14536
rect 2808 14504 2848 14536
rect 2880 14504 2920 14536
rect 2952 14504 2992 14536
rect 3024 14504 3064 14536
rect 3096 14504 3136 14536
rect 3168 14504 3208 14536
rect 3240 14504 3280 14536
rect 3312 14504 3352 14536
rect 3384 14504 3424 14536
rect 3456 14504 3496 14536
rect 3528 14504 3568 14536
rect 3600 14504 3640 14536
rect 3672 14504 3712 14536
rect 3744 14504 3784 14536
rect 3816 14504 3856 14536
rect 3888 14504 4000 14536
rect 0 14464 4000 14504
rect 0 14432 112 14464
rect 144 14432 184 14464
rect 216 14432 256 14464
rect 288 14432 328 14464
rect 360 14432 400 14464
rect 432 14432 472 14464
rect 504 14432 544 14464
rect 576 14432 616 14464
rect 648 14432 688 14464
rect 720 14432 760 14464
rect 792 14432 832 14464
rect 864 14432 904 14464
rect 936 14432 976 14464
rect 1008 14432 1048 14464
rect 1080 14432 1120 14464
rect 1152 14432 1192 14464
rect 1224 14432 1264 14464
rect 1296 14432 1336 14464
rect 1368 14432 1408 14464
rect 1440 14432 1480 14464
rect 1512 14432 1552 14464
rect 1584 14432 1624 14464
rect 1656 14432 1696 14464
rect 1728 14432 1768 14464
rect 1800 14432 1840 14464
rect 1872 14432 1912 14464
rect 1944 14432 1984 14464
rect 2016 14432 2056 14464
rect 2088 14432 2128 14464
rect 2160 14432 2200 14464
rect 2232 14432 2272 14464
rect 2304 14432 2344 14464
rect 2376 14432 2416 14464
rect 2448 14432 2488 14464
rect 2520 14432 2560 14464
rect 2592 14432 2632 14464
rect 2664 14432 2704 14464
rect 2736 14432 2776 14464
rect 2808 14432 2848 14464
rect 2880 14432 2920 14464
rect 2952 14432 2992 14464
rect 3024 14432 3064 14464
rect 3096 14432 3136 14464
rect 3168 14432 3208 14464
rect 3240 14432 3280 14464
rect 3312 14432 3352 14464
rect 3384 14432 3424 14464
rect 3456 14432 3496 14464
rect 3528 14432 3568 14464
rect 3600 14432 3640 14464
rect 3672 14432 3712 14464
rect 3744 14432 3784 14464
rect 3816 14432 3856 14464
rect 3888 14432 4000 14464
rect 0 14392 4000 14432
rect 0 14360 112 14392
rect 144 14360 184 14392
rect 216 14360 256 14392
rect 288 14360 328 14392
rect 360 14360 400 14392
rect 432 14360 472 14392
rect 504 14360 544 14392
rect 576 14360 616 14392
rect 648 14360 688 14392
rect 720 14360 760 14392
rect 792 14360 832 14392
rect 864 14360 904 14392
rect 936 14360 976 14392
rect 1008 14360 1048 14392
rect 1080 14360 1120 14392
rect 1152 14360 1192 14392
rect 1224 14360 1264 14392
rect 1296 14360 1336 14392
rect 1368 14360 1408 14392
rect 1440 14360 1480 14392
rect 1512 14360 1552 14392
rect 1584 14360 1624 14392
rect 1656 14360 1696 14392
rect 1728 14360 1768 14392
rect 1800 14360 1840 14392
rect 1872 14360 1912 14392
rect 1944 14360 1984 14392
rect 2016 14360 2056 14392
rect 2088 14360 2128 14392
rect 2160 14360 2200 14392
rect 2232 14360 2272 14392
rect 2304 14360 2344 14392
rect 2376 14360 2416 14392
rect 2448 14360 2488 14392
rect 2520 14360 2560 14392
rect 2592 14360 2632 14392
rect 2664 14360 2704 14392
rect 2736 14360 2776 14392
rect 2808 14360 2848 14392
rect 2880 14360 2920 14392
rect 2952 14360 2992 14392
rect 3024 14360 3064 14392
rect 3096 14360 3136 14392
rect 3168 14360 3208 14392
rect 3240 14360 3280 14392
rect 3312 14360 3352 14392
rect 3384 14360 3424 14392
rect 3456 14360 3496 14392
rect 3528 14360 3568 14392
rect 3600 14360 3640 14392
rect 3672 14360 3712 14392
rect 3744 14360 3784 14392
rect 3816 14360 3856 14392
rect 3888 14360 4000 14392
rect 0 14320 4000 14360
rect 0 14288 112 14320
rect 144 14288 184 14320
rect 216 14288 256 14320
rect 288 14288 328 14320
rect 360 14288 400 14320
rect 432 14288 472 14320
rect 504 14288 544 14320
rect 576 14288 616 14320
rect 648 14288 688 14320
rect 720 14288 760 14320
rect 792 14288 832 14320
rect 864 14288 904 14320
rect 936 14288 976 14320
rect 1008 14288 1048 14320
rect 1080 14288 1120 14320
rect 1152 14288 1192 14320
rect 1224 14288 1264 14320
rect 1296 14288 1336 14320
rect 1368 14288 1408 14320
rect 1440 14288 1480 14320
rect 1512 14288 1552 14320
rect 1584 14288 1624 14320
rect 1656 14288 1696 14320
rect 1728 14288 1768 14320
rect 1800 14288 1840 14320
rect 1872 14288 1912 14320
rect 1944 14288 1984 14320
rect 2016 14288 2056 14320
rect 2088 14288 2128 14320
rect 2160 14288 2200 14320
rect 2232 14288 2272 14320
rect 2304 14288 2344 14320
rect 2376 14288 2416 14320
rect 2448 14288 2488 14320
rect 2520 14288 2560 14320
rect 2592 14288 2632 14320
rect 2664 14288 2704 14320
rect 2736 14288 2776 14320
rect 2808 14288 2848 14320
rect 2880 14288 2920 14320
rect 2952 14288 2992 14320
rect 3024 14288 3064 14320
rect 3096 14288 3136 14320
rect 3168 14288 3208 14320
rect 3240 14288 3280 14320
rect 3312 14288 3352 14320
rect 3384 14288 3424 14320
rect 3456 14288 3496 14320
rect 3528 14288 3568 14320
rect 3600 14288 3640 14320
rect 3672 14288 3712 14320
rect 3744 14288 3784 14320
rect 3816 14288 3856 14320
rect 3888 14288 4000 14320
rect 0 14248 4000 14288
rect 0 14216 112 14248
rect 144 14216 184 14248
rect 216 14216 256 14248
rect 288 14216 328 14248
rect 360 14216 400 14248
rect 432 14216 472 14248
rect 504 14216 544 14248
rect 576 14216 616 14248
rect 648 14216 688 14248
rect 720 14216 760 14248
rect 792 14216 832 14248
rect 864 14216 904 14248
rect 936 14216 976 14248
rect 1008 14216 1048 14248
rect 1080 14216 1120 14248
rect 1152 14216 1192 14248
rect 1224 14216 1264 14248
rect 1296 14216 1336 14248
rect 1368 14216 1408 14248
rect 1440 14216 1480 14248
rect 1512 14216 1552 14248
rect 1584 14216 1624 14248
rect 1656 14216 1696 14248
rect 1728 14216 1768 14248
rect 1800 14216 1840 14248
rect 1872 14216 1912 14248
rect 1944 14216 1984 14248
rect 2016 14216 2056 14248
rect 2088 14216 2128 14248
rect 2160 14216 2200 14248
rect 2232 14216 2272 14248
rect 2304 14216 2344 14248
rect 2376 14216 2416 14248
rect 2448 14216 2488 14248
rect 2520 14216 2560 14248
rect 2592 14216 2632 14248
rect 2664 14216 2704 14248
rect 2736 14216 2776 14248
rect 2808 14216 2848 14248
rect 2880 14216 2920 14248
rect 2952 14216 2992 14248
rect 3024 14216 3064 14248
rect 3096 14216 3136 14248
rect 3168 14216 3208 14248
rect 3240 14216 3280 14248
rect 3312 14216 3352 14248
rect 3384 14216 3424 14248
rect 3456 14216 3496 14248
rect 3528 14216 3568 14248
rect 3600 14216 3640 14248
rect 3672 14216 3712 14248
rect 3744 14216 3784 14248
rect 3816 14216 3856 14248
rect 3888 14216 4000 14248
rect 0 14176 4000 14216
rect 0 14144 112 14176
rect 144 14144 184 14176
rect 216 14144 256 14176
rect 288 14144 328 14176
rect 360 14144 400 14176
rect 432 14144 472 14176
rect 504 14144 544 14176
rect 576 14144 616 14176
rect 648 14144 688 14176
rect 720 14144 760 14176
rect 792 14144 832 14176
rect 864 14144 904 14176
rect 936 14144 976 14176
rect 1008 14144 1048 14176
rect 1080 14144 1120 14176
rect 1152 14144 1192 14176
rect 1224 14144 1264 14176
rect 1296 14144 1336 14176
rect 1368 14144 1408 14176
rect 1440 14144 1480 14176
rect 1512 14144 1552 14176
rect 1584 14144 1624 14176
rect 1656 14144 1696 14176
rect 1728 14144 1768 14176
rect 1800 14144 1840 14176
rect 1872 14144 1912 14176
rect 1944 14144 1984 14176
rect 2016 14144 2056 14176
rect 2088 14144 2128 14176
rect 2160 14144 2200 14176
rect 2232 14144 2272 14176
rect 2304 14144 2344 14176
rect 2376 14144 2416 14176
rect 2448 14144 2488 14176
rect 2520 14144 2560 14176
rect 2592 14144 2632 14176
rect 2664 14144 2704 14176
rect 2736 14144 2776 14176
rect 2808 14144 2848 14176
rect 2880 14144 2920 14176
rect 2952 14144 2992 14176
rect 3024 14144 3064 14176
rect 3096 14144 3136 14176
rect 3168 14144 3208 14176
rect 3240 14144 3280 14176
rect 3312 14144 3352 14176
rect 3384 14144 3424 14176
rect 3456 14144 3496 14176
rect 3528 14144 3568 14176
rect 3600 14144 3640 14176
rect 3672 14144 3712 14176
rect 3744 14144 3784 14176
rect 3816 14144 3856 14176
rect 3888 14144 4000 14176
rect 0 14104 4000 14144
rect 0 14072 112 14104
rect 144 14072 184 14104
rect 216 14072 256 14104
rect 288 14072 328 14104
rect 360 14072 400 14104
rect 432 14072 472 14104
rect 504 14072 544 14104
rect 576 14072 616 14104
rect 648 14072 688 14104
rect 720 14072 760 14104
rect 792 14072 832 14104
rect 864 14072 904 14104
rect 936 14072 976 14104
rect 1008 14072 1048 14104
rect 1080 14072 1120 14104
rect 1152 14072 1192 14104
rect 1224 14072 1264 14104
rect 1296 14072 1336 14104
rect 1368 14072 1408 14104
rect 1440 14072 1480 14104
rect 1512 14072 1552 14104
rect 1584 14072 1624 14104
rect 1656 14072 1696 14104
rect 1728 14072 1768 14104
rect 1800 14072 1840 14104
rect 1872 14072 1912 14104
rect 1944 14072 1984 14104
rect 2016 14072 2056 14104
rect 2088 14072 2128 14104
rect 2160 14072 2200 14104
rect 2232 14072 2272 14104
rect 2304 14072 2344 14104
rect 2376 14072 2416 14104
rect 2448 14072 2488 14104
rect 2520 14072 2560 14104
rect 2592 14072 2632 14104
rect 2664 14072 2704 14104
rect 2736 14072 2776 14104
rect 2808 14072 2848 14104
rect 2880 14072 2920 14104
rect 2952 14072 2992 14104
rect 3024 14072 3064 14104
rect 3096 14072 3136 14104
rect 3168 14072 3208 14104
rect 3240 14072 3280 14104
rect 3312 14072 3352 14104
rect 3384 14072 3424 14104
rect 3456 14072 3496 14104
rect 3528 14072 3568 14104
rect 3600 14072 3640 14104
rect 3672 14072 3712 14104
rect 3744 14072 3784 14104
rect 3816 14072 3856 14104
rect 3888 14072 4000 14104
rect 0 14032 4000 14072
rect 0 14000 112 14032
rect 144 14000 184 14032
rect 216 14000 256 14032
rect 288 14000 328 14032
rect 360 14000 400 14032
rect 432 14000 472 14032
rect 504 14000 544 14032
rect 576 14000 616 14032
rect 648 14000 688 14032
rect 720 14000 760 14032
rect 792 14000 832 14032
rect 864 14000 904 14032
rect 936 14000 976 14032
rect 1008 14000 1048 14032
rect 1080 14000 1120 14032
rect 1152 14000 1192 14032
rect 1224 14000 1264 14032
rect 1296 14000 1336 14032
rect 1368 14000 1408 14032
rect 1440 14000 1480 14032
rect 1512 14000 1552 14032
rect 1584 14000 1624 14032
rect 1656 14000 1696 14032
rect 1728 14000 1768 14032
rect 1800 14000 1840 14032
rect 1872 14000 1912 14032
rect 1944 14000 1984 14032
rect 2016 14000 2056 14032
rect 2088 14000 2128 14032
rect 2160 14000 2200 14032
rect 2232 14000 2272 14032
rect 2304 14000 2344 14032
rect 2376 14000 2416 14032
rect 2448 14000 2488 14032
rect 2520 14000 2560 14032
rect 2592 14000 2632 14032
rect 2664 14000 2704 14032
rect 2736 14000 2776 14032
rect 2808 14000 2848 14032
rect 2880 14000 2920 14032
rect 2952 14000 2992 14032
rect 3024 14000 3064 14032
rect 3096 14000 3136 14032
rect 3168 14000 3208 14032
rect 3240 14000 3280 14032
rect 3312 14000 3352 14032
rect 3384 14000 3424 14032
rect 3456 14000 3496 14032
rect 3528 14000 3568 14032
rect 3600 14000 3640 14032
rect 3672 14000 3712 14032
rect 3744 14000 3784 14032
rect 3816 14000 3856 14032
rect 3888 14000 4000 14032
rect 0 13960 4000 14000
rect 0 13928 112 13960
rect 144 13928 184 13960
rect 216 13928 256 13960
rect 288 13928 328 13960
rect 360 13928 400 13960
rect 432 13928 472 13960
rect 504 13928 544 13960
rect 576 13928 616 13960
rect 648 13928 688 13960
rect 720 13928 760 13960
rect 792 13928 832 13960
rect 864 13928 904 13960
rect 936 13928 976 13960
rect 1008 13928 1048 13960
rect 1080 13928 1120 13960
rect 1152 13928 1192 13960
rect 1224 13928 1264 13960
rect 1296 13928 1336 13960
rect 1368 13928 1408 13960
rect 1440 13928 1480 13960
rect 1512 13928 1552 13960
rect 1584 13928 1624 13960
rect 1656 13928 1696 13960
rect 1728 13928 1768 13960
rect 1800 13928 1840 13960
rect 1872 13928 1912 13960
rect 1944 13928 1984 13960
rect 2016 13928 2056 13960
rect 2088 13928 2128 13960
rect 2160 13928 2200 13960
rect 2232 13928 2272 13960
rect 2304 13928 2344 13960
rect 2376 13928 2416 13960
rect 2448 13928 2488 13960
rect 2520 13928 2560 13960
rect 2592 13928 2632 13960
rect 2664 13928 2704 13960
rect 2736 13928 2776 13960
rect 2808 13928 2848 13960
rect 2880 13928 2920 13960
rect 2952 13928 2992 13960
rect 3024 13928 3064 13960
rect 3096 13928 3136 13960
rect 3168 13928 3208 13960
rect 3240 13928 3280 13960
rect 3312 13928 3352 13960
rect 3384 13928 3424 13960
rect 3456 13928 3496 13960
rect 3528 13928 3568 13960
rect 3600 13928 3640 13960
rect 3672 13928 3712 13960
rect 3744 13928 3784 13960
rect 3816 13928 3856 13960
rect 3888 13928 4000 13960
rect 0 13888 4000 13928
rect 0 13856 112 13888
rect 144 13856 184 13888
rect 216 13856 256 13888
rect 288 13856 328 13888
rect 360 13856 400 13888
rect 432 13856 472 13888
rect 504 13856 544 13888
rect 576 13856 616 13888
rect 648 13856 688 13888
rect 720 13856 760 13888
rect 792 13856 832 13888
rect 864 13856 904 13888
rect 936 13856 976 13888
rect 1008 13856 1048 13888
rect 1080 13856 1120 13888
rect 1152 13856 1192 13888
rect 1224 13856 1264 13888
rect 1296 13856 1336 13888
rect 1368 13856 1408 13888
rect 1440 13856 1480 13888
rect 1512 13856 1552 13888
rect 1584 13856 1624 13888
rect 1656 13856 1696 13888
rect 1728 13856 1768 13888
rect 1800 13856 1840 13888
rect 1872 13856 1912 13888
rect 1944 13856 1984 13888
rect 2016 13856 2056 13888
rect 2088 13856 2128 13888
rect 2160 13856 2200 13888
rect 2232 13856 2272 13888
rect 2304 13856 2344 13888
rect 2376 13856 2416 13888
rect 2448 13856 2488 13888
rect 2520 13856 2560 13888
rect 2592 13856 2632 13888
rect 2664 13856 2704 13888
rect 2736 13856 2776 13888
rect 2808 13856 2848 13888
rect 2880 13856 2920 13888
rect 2952 13856 2992 13888
rect 3024 13856 3064 13888
rect 3096 13856 3136 13888
rect 3168 13856 3208 13888
rect 3240 13856 3280 13888
rect 3312 13856 3352 13888
rect 3384 13856 3424 13888
rect 3456 13856 3496 13888
rect 3528 13856 3568 13888
rect 3600 13856 3640 13888
rect 3672 13856 3712 13888
rect 3744 13856 3784 13888
rect 3816 13856 3856 13888
rect 3888 13856 4000 13888
rect 0 13816 4000 13856
rect 0 13784 112 13816
rect 144 13784 184 13816
rect 216 13784 256 13816
rect 288 13784 328 13816
rect 360 13784 400 13816
rect 432 13784 472 13816
rect 504 13784 544 13816
rect 576 13784 616 13816
rect 648 13784 688 13816
rect 720 13784 760 13816
rect 792 13784 832 13816
rect 864 13784 904 13816
rect 936 13784 976 13816
rect 1008 13784 1048 13816
rect 1080 13784 1120 13816
rect 1152 13784 1192 13816
rect 1224 13784 1264 13816
rect 1296 13784 1336 13816
rect 1368 13784 1408 13816
rect 1440 13784 1480 13816
rect 1512 13784 1552 13816
rect 1584 13784 1624 13816
rect 1656 13784 1696 13816
rect 1728 13784 1768 13816
rect 1800 13784 1840 13816
rect 1872 13784 1912 13816
rect 1944 13784 1984 13816
rect 2016 13784 2056 13816
rect 2088 13784 2128 13816
rect 2160 13784 2200 13816
rect 2232 13784 2272 13816
rect 2304 13784 2344 13816
rect 2376 13784 2416 13816
rect 2448 13784 2488 13816
rect 2520 13784 2560 13816
rect 2592 13784 2632 13816
rect 2664 13784 2704 13816
rect 2736 13784 2776 13816
rect 2808 13784 2848 13816
rect 2880 13784 2920 13816
rect 2952 13784 2992 13816
rect 3024 13784 3064 13816
rect 3096 13784 3136 13816
rect 3168 13784 3208 13816
rect 3240 13784 3280 13816
rect 3312 13784 3352 13816
rect 3384 13784 3424 13816
rect 3456 13784 3496 13816
rect 3528 13784 3568 13816
rect 3600 13784 3640 13816
rect 3672 13784 3712 13816
rect 3744 13784 3784 13816
rect 3816 13784 3856 13816
rect 3888 13784 4000 13816
rect 0 13744 4000 13784
rect 0 13712 112 13744
rect 144 13712 184 13744
rect 216 13712 256 13744
rect 288 13712 328 13744
rect 360 13712 400 13744
rect 432 13712 472 13744
rect 504 13712 544 13744
rect 576 13712 616 13744
rect 648 13712 688 13744
rect 720 13712 760 13744
rect 792 13712 832 13744
rect 864 13712 904 13744
rect 936 13712 976 13744
rect 1008 13712 1048 13744
rect 1080 13712 1120 13744
rect 1152 13712 1192 13744
rect 1224 13712 1264 13744
rect 1296 13712 1336 13744
rect 1368 13712 1408 13744
rect 1440 13712 1480 13744
rect 1512 13712 1552 13744
rect 1584 13712 1624 13744
rect 1656 13712 1696 13744
rect 1728 13712 1768 13744
rect 1800 13712 1840 13744
rect 1872 13712 1912 13744
rect 1944 13712 1984 13744
rect 2016 13712 2056 13744
rect 2088 13712 2128 13744
rect 2160 13712 2200 13744
rect 2232 13712 2272 13744
rect 2304 13712 2344 13744
rect 2376 13712 2416 13744
rect 2448 13712 2488 13744
rect 2520 13712 2560 13744
rect 2592 13712 2632 13744
rect 2664 13712 2704 13744
rect 2736 13712 2776 13744
rect 2808 13712 2848 13744
rect 2880 13712 2920 13744
rect 2952 13712 2992 13744
rect 3024 13712 3064 13744
rect 3096 13712 3136 13744
rect 3168 13712 3208 13744
rect 3240 13712 3280 13744
rect 3312 13712 3352 13744
rect 3384 13712 3424 13744
rect 3456 13712 3496 13744
rect 3528 13712 3568 13744
rect 3600 13712 3640 13744
rect 3672 13712 3712 13744
rect 3744 13712 3784 13744
rect 3816 13712 3856 13744
rect 3888 13712 4000 13744
rect 0 13672 4000 13712
rect 0 13640 112 13672
rect 144 13640 184 13672
rect 216 13640 256 13672
rect 288 13640 328 13672
rect 360 13640 400 13672
rect 432 13640 472 13672
rect 504 13640 544 13672
rect 576 13640 616 13672
rect 648 13640 688 13672
rect 720 13640 760 13672
rect 792 13640 832 13672
rect 864 13640 904 13672
rect 936 13640 976 13672
rect 1008 13640 1048 13672
rect 1080 13640 1120 13672
rect 1152 13640 1192 13672
rect 1224 13640 1264 13672
rect 1296 13640 1336 13672
rect 1368 13640 1408 13672
rect 1440 13640 1480 13672
rect 1512 13640 1552 13672
rect 1584 13640 1624 13672
rect 1656 13640 1696 13672
rect 1728 13640 1768 13672
rect 1800 13640 1840 13672
rect 1872 13640 1912 13672
rect 1944 13640 1984 13672
rect 2016 13640 2056 13672
rect 2088 13640 2128 13672
rect 2160 13640 2200 13672
rect 2232 13640 2272 13672
rect 2304 13640 2344 13672
rect 2376 13640 2416 13672
rect 2448 13640 2488 13672
rect 2520 13640 2560 13672
rect 2592 13640 2632 13672
rect 2664 13640 2704 13672
rect 2736 13640 2776 13672
rect 2808 13640 2848 13672
rect 2880 13640 2920 13672
rect 2952 13640 2992 13672
rect 3024 13640 3064 13672
rect 3096 13640 3136 13672
rect 3168 13640 3208 13672
rect 3240 13640 3280 13672
rect 3312 13640 3352 13672
rect 3384 13640 3424 13672
rect 3456 13640 3496 13672
rect 3528 13640 3568 13672
rect 3600 13640 3640 13672
rect 3672 13640 3712 13672
rect 3744 13640 3784 13672
rect 3816 13640 3856 13672
rect 3888 13640 4000 13672
rect 0 13600 4000 13640
rect 0 13568 112 13600
rect 144 13568 184 13600
rect 216 13568 256 13600
rect 288 13568 328 13600
rect 360 13568 400 13600
rect 432 13568 472 13600
rect 504 13568 544 13600
rect 576 13568 616 13600
rect 648 13568 688 13600
rect 720 13568 760 13600
rect 792 13568 832 13600
rect 864 13568 904 13600
rect 936 13568 976 13600
rect 1008 13568 1048 13600
rect 1080 13568 1120 13600
rect 1152 13568 1192 13600
rect 1224 13568 1264 13600
rect 1296 13568 1336 13600
rect 1368 13568 1408 13600
rect 1440 13568 1480 13600
rect 1512 13568 1552 13600
rect 1584 13568 1624 13600
rect 1656 13568 1696 13600
rect 1728 13568 1768 13600
rect 1800 13568 1840 13600
rect 1872 13568 1912 13600
rect 1944 13568 1984 13600
rect 2016 13568 2056 13600
rect 2088 13568 2128 13600
rect 2160 13568 2200 13600
rect 2232 13568 2272 13600
rect 2304 13568 2344 13600
rect 2376 13568 2416 13600
rect 2448 13568 2488 13600
rect 2520 13568 2560 13600
rect 2592 13568 2632 13600
rect 2664 13568 2704 13600
rect 2736 13568 2776 13600
rect 2808 13568 2848 13600
rect 2880 13568 2920 13600
rect 2952 13568 2992 13600
rect 3024 13568 3064 13600
rect 3096 13568 3136 13600
rect 3168 13568 3208 13600
rect 3240 13568 3280 13600
rect 3312 13568 3352 13600
rect 3384 13568 3424 13600
rect 3456 13568 3496 13600
rect 3528 13568 3568 13600
rect 3600 13568 3640 13600
rect 3672 13568 3712 13600
rect 3744 13568 3784 13600
rect 3816 13568 3856 13600
rect 3888 13568 4000 13600
rect 0 13528 4000 13568
rect 0 13496 112 13528
rect 144 13496 184 13528
rect 216 13496 256 13528
rect 288 13496 328 13528
rect 360 13496 400 13528
rect 432 13496 472 13528
rect 504 13496 544 13528
rect 576 13496 616 13528
rect 648 13496 688 13528
rect 720 13496 760 13528
rect 792 13496 832 13528
rect 864 13496 904 13528
rect 936 13496 976 13528
rect 1008 13496 1048 13528
rect 1080 13496 1120 13528
rect 1152 13496 1192 13528
rect 1224 13496 1264 13528
rect 1296 13496 1336 13528
rect 1368 13496 1408 13528
rect 1440 13496 1480 13528
rect 1512 13496 1552 13528
rect 1584 13496 1624 13528
rect 1656 13496 1696 13528
rect 1728 13496 1768 13528
rect 1800 13496 1840 13528
rect 1872 13496 1912 13528
rect 1944 13496 1984 13528
rect 2016 13496 2056 13528
rect 2088 13496 2128 13528
rect 2160 13496 2200 13528
rect 2232 13496 2272 13528
rect 2304 13496 2344 13528
rect 2376 13496 2416 13528
rect 2448 13496 2488 13528
rect 2520 13496 2560 13528
rect 2592 13496 2632 13528
rect 2664 13496 2704 13528
rect 2736 13496 2776 13528
rect 2808 13496 2848 13528
rect 2880 13496 2920 13528
rect 2952 13496 2992 13528
rect 3024 13496 3064 13528
rect 3096 13496 3136 13528
rect 3168 13496 3208 13528
rect 3240 13496 3280 13528
rect 3312 13496 3352 13528
rect 3384 13496 3424 13528
rect 3456 13496 3496 13528
rect 3528 13496 3568 13528
rect 3600 13496 3640 13528
rect 3672 13496 3712 13528
rect 3744 13496 3784 13528
rect 3816 13496 3856 13528
rect 3888 13496 4000 13528
rect 0 13456 4000 13496
rect 0 13424 112 13456
rect 144 13424 184 13456
rect 216 13424 256 13456
rect 288 13424 328 13456
rect 360 13424 400 13456
rect 432 13424 472 13456
rect 504 13424 544 13456
rect 576 13424 616 13456
rect 648 13424 688 13456
rect 720 13424 760 13456
rect 792 13424 832 13456
rect 864 13424 904 13456
rect 936 13424 976 13456
rect 1008 13424 1048 13456
rect 1080 13424 1120 13456
rect 1152 13424 1192 13456
rect 1224 13424 1264 13456
rect 1296 13424 1336 13456
rect 1368 13424 1408 13456
rect 1440 13424 1480 13456
rect 1512 13424 1552 13456
rect 1584 13424 1624 13456
rect 1656 13424 1696 13456
rect 1728 13424 1768 13456
rect 1800 13424 1840 13456
rect 1872 13424 1912 13456
rect 1944 13424 1984 13456
rect 2016 13424 2056 13456
rect 2088 13424 2128 13456
rect 2160 13424 2200 13456
rect 2232 13424 2272 13456
rect 2304 13424 2344 13456
rect 2376 13424 2416 13456
rect 2448 13424 2488 13456
rect 2520 13424 2560 13456
rect 2592 13424 2632 13456
rect 2664 13424 2704 13456
rect 2736 13424 2776 13456
rect 2808 13424 2848 13456
rect 2880 13424 2920 13456
rect 2952 13424 2992 13456
rect 3024 13424 3064 13456
rect 3096 13424 3136 13456
rect 3168 13424 3208 13456
rect 3240 13424 3280 13456
rect 3312 13424 3352 13456
rect 3384 13424 3424 13456
rect 3456 13424 3496 13456
rect 3528 13424 3568 13456
rect 3600 13424 3640 13456
rect 3672 13424 3712 13456
rect 3744 13424 3784 13456
rect 3816 13424 3856 13456
rect 3888 13424 4000 13456
rect 0 13384 4000 13424
rect 0 13352 112 13384
rect 144 13352 184 13384
rect 216 13352 256 13384
rect 288 13352 328 13384
rect 360 13352 400 13384
rect 432 13352 472 13384
rect 504 13352 544 13384
rect 576 13352 616 13384
rect 648 13352 688 13384
rect 720 13352 760 13384
rect 792 13352 832 13384
rect 864 13352 904 13384
rect 936 13352 976 13384
rect 1008 13352 1048 13384
rect 1080 13352 1120 13384
rect 1152 13352 1192 13384
rect 1224 13352 1264 13384
rect 1296 13352 1336 13384
rect 1368 13352 1408 13384
rect 1440 13352 1480 13384
rect 1512 13352 1552 13384
rect 1584 13352 1624 13384
rect 1656 13352 1696 13384
rect 1728 13352 1768 13384
rect 1800 13352 1840 13384
rect 1872 13352 1912 13384
rect 1944 13352 1984 13384
rect 2016 13352 2056 13384
rect 2088 13352 2128 13384
rect 2160 13352 2200 13384
rect 2232 13352 2272 13384
rect 2304 13352 2344 13384
rect 2376 13352 2416 13384
rect 2448 13352 2488 13384
rect 2520 13352 2560 13384
rect 2592 13352 2632 13384
rect 2664 13352 2704 13384
rect 2736 13352 2776 13384
rect 2808 13352 2848 13384
rect 2880 13352 2920 13384
rect 2952 13352 2992 13384
rect 3024 13352 3064 13384
rect 3096 13352 3136 13384
rect 3168 13352 3208 13384
rect 3240 13352 3280 13384
rect 3312 13352 3352 13384
rect 3384 13352 3424 13384
rect 3456 13352 3496 13384
rect 3528 13352 3568 13384
rect 3600 13352 3640 13384
rect 3672 13352 3712 13384
rect 3744 13352 3784 13384
rect 3816 13352 3856 13384
rect 3888 13352 4000 13384
rect 0 13312 4000 13352
rect 0 13280 112 13312
rect 144 13280 184 13312
rect 216 13280 256 13312
rect 288 13280 328 13312
rect 360 13280 400 13312
rect 432 13280 472 13312
rect 504 13280 544 13312
rect 576 13280 616 13312
rect 648 13280 688 13312
rect 720 13280 760 13312
rect 792 13280 832 13312
rect 864 13280 904 13312
rect 936 13280 976 13312
rect 1008 13280 1048 13312
rect 1080 13280 1120 13312
rect 1152 13280 1192 13312
rect 1224 13280 1264 13312
rect 1296 13280 1336 13312
rect 1368 13280 1408 13312
rect 1440 13280 1480 13312
rect 1512 13280 1552 13312
rect 1584 13280 1624 13312
rect 1656 13280 1696 13312
rect 1728 13280 1768 13312
rect 1800 13280 1840 13312
rect 1872 13280 1912 13312
rect 1944 13280 1984 13312
rect 2016 13280 2056 13312
rect 2088 13280 2128 13312
rect 2160 13280 2200 13312
rect 2232 13280 2272 13312
rect 2304 13280 2344 13312
rect 2376 13280 2416 13312
rect 2448 13280 2488 13312
rect 2520 13280 2560 13312
rect 2592 13280 2632 13312
rect 2664 13280 2704 13312
rect 2736 13280 2776 13312
rect 2808 13280 2848 13312
rect 2880 13280 2920 13312
rect 2952 13280 2992 13312
rect 3024 13280 3064 13312
rect 3096 13280 3136 13312
rect 3168 13280 3208 13312
rect 3240 13280 3280 13312
rect 3312 13280 3352 13312
rect 3384 13280 3424 13312
rect 3456 13280 3496 13312
rect 3528 13280 3568 13312
rect 3600 13280 3640 13312
rect 3672 13280 3712 13312
rect 3744 13280 3784 13312
rect 3816 13280 3856 13312
rect 3888 13280 4000 13312
rect 0 13240 4000 13280
rect 0 13208 112 13240
rect 144 13208 184 13240
rect 216 13208 256 13240
rect 288 13208 328 13240
rect 360 13208 400 13240
rect 432 13208 472 13240
rect 504 13208 544 13240
rect 576 13208 616 13240
rect 648 13208 688 13240
rect 720 13208 760 13240
rect 792 13208 832 13240
rect 864 13208 904 13240
rect 936 13208 976 13240
rect 1008 13208 1048 13240
rect 1080 13208 1120 13240
rect 1152 13208 1192 13240
rect 1224 13208 1264 13240
rect 1296 13208 1336 13240
rect 1368 13208 1408 13240
rect 1440 13208 1480 13240
rect 1512 13208 1552 13240
rect 1584 13208 1624 13240
rect 1656 13208 1696 13240
rect 1728 13208 1768 13240
rect 1800 13208 1840 13240
rect 1872 13208 1912 13240
rect 1944 13208 1984 13240
rect 2016 13208 2056 13240
rect 2088 13208 2128 13240
rect 2160 13208 2200 13240
rect 2232 13208 2272 13240
rect 2304 13208 2344 13240
rect 2376 13208 2416 13240
rect 2448 13208 2488 13240
rect 2520 13208 2560 13240
rect 2592 13208 2632 13240
rect 2664 13208 2704 13240
rect 2736 13208 2776 13240
rect 2808 13208 2848 13240
rect 2880 13208 2920 13240
rect 2952 13208 2992 13240
rect 3024 13208 3064 13240
rect 3096 13208 3136 13240
rect 3168 13208 3208 13240
rect 3240 13208 3280 13240
rect 3312 13208 3352 13240
rect 3384 13208 3424 13240
rect 3456 13208 3496 13240
rect 3528 13208 3568 13240
rect 3600 13208 3640 13240
rect 3672 13208 3712 13240
rect 3744 13208 3784 13240
rect 3816 13208 3856 13240
rect 3888 13208 4000 13240
rect 0 13168 4000 13208
rect 0 13136 112 13168
rect 144 13136 184 13168
rect 216 13136 256 13168
rect 288 13136 328 13168
rect 360 13136 400 13168
rect 432 13136 472 13168
rect 504 13136 544 13168
rect 576 13136 616 13168
rect 648 13136 688 13168
rect 720 13136 760 13168
rect 792 13136 832 13168
rect 864 13136 904 13168
rect 936 13136 976 13168
rect 1008 13136 1048 13168
rect 1080 13136 1120 13168
rect 1152 13136 1192 13168
rect 1224 13136 1264 13168
rect 1296 13136 1336 13168
rect 1368 13136 1408 13168
rect 1440 13136 1480 13168
rect 1512 13136 1552 13168
rect 1584 13136 1624 13168
rect 1656 13136 1696 13168
rect 1728 13136 1768 13168
rect 1800 13136 1840 13168
rect 1872 13136 1912 13168
rect 1944 13136 1984 13168
rect 2016 13136 2056 13168
rect 2088 13136 2128 13168
rect 2160 13136 2200 13168
rect 2232 13136 2272 13168
rect 2304 13136 2344 13168
rect 2376 13136 2416 13168
rect 2448 13136 2488 13168
rect 2520 13136 2560 13168
rect 2592 13136 2632 13168
rect 2664 13136 2704 13168
rect 2736 13136 2776 13168
rect 2808 13136 2848 13168
rect 2880 13136 2920 13168
rect 2952 13136 2992 13168
rect 3024 13136 3064 13168
rect 3096 13136 3136 13168
rect 3168 13136 3208 13168
rect 3240 13136 3280 13168
rect 3312 13136 3352 13168
rect 3384 13136 3424 13168
rect 3456 13136 3496 13168
rect 3528 13136 3568 13168
rect 3600 13136 3640 13168
rect 3672 13136 3712 13168
rect 3744 13136 3784 13168
rect 3816 13136 3856 13168
rect 3888 13136 4000 13168
rect 0 13096 4000 13136
rect 0 13064 112 13096
rect 144 13064 184 13096
rect 216 13064 256 13096
rect 288 13064 328 13096
rect 360 13064 400 13096
rect 432 13064 472 13096
rect 504 13064 544 13096
rect 576 13064 616 13096
rect 648 13064 688 13096
rect 720 13064 760 13096
rect 792 13064 832 13096
rect 864 13064 904 13096
rect 936 13064 976 13096
rect 1008 13064 1048 13096
rect 1080 13064 1120 13096
rect 1152 13064 1192 13096
rect 1224 13064 1264 13096
rect 1296 13064 1336 13096
rect 1368 13064 1408 13096
rect 1440 13064 1480 13096
rect 1512 13064 1552 13096
rect 1584 13064 1624 13096
rect 1656 13064 1696 13096
rect 1728 13064 1768 13096
rect 1800 13064 1840 13096
rect 1872 13064 1912 13096
rect 1944 13064 1984 13096
rect 2016 13064 2056 13096
rect 2088 13064 2128 13096
rect 2160 13064 2200 13096
rect 2232 13064 2272 13096
rect 2304 13064 2344 13096
rect 2376 13064 2416 13096
rect 2448 13064 2488 13096
rect 2520 13064 2560 13096
rect 2592 13064 2632 13096
rect 2664 13064 2704 13096
rect 2736 13064 2776 13096
rect 2808 13064 2848 13096
rect 2880 13064 2920 13096
rect 2952 13064 2992 13096
rect 3024 13064 3064 13096
rect 3096 13064 3136 13096
rect 3168 13064 3208 13096
rect 3240 13064 3280 13096
rect 3312 13064 3352 13096
rect 3384 13064 3424 13096
rect 3456 13064 3496 13096
rect 3528 13064 3568 13096
rect 3600 13064 3640 13096
rect 3672 13064 3712 13096
rect 3744 13064 3784 13096
rect 3816 13064 3856 13096
rect 3888 13064 4000 13096
rect 0 13000 4000 13064
rect 0 12144 4000 12200
rect 0 12112 40 12144
rect 72 12112 112 12144
rect 144 12112 184 12144
rect 216 12112 256 12144
rect 288 12112 328 12144
rect 360 12112 400 12144
rect 432 12112 472 12144
rect 504 12112 544 12144
rect 576 12112 616 12144
rect 648 12112 688 12144
rect 720 12112 760 12144
rect 792 12112 832 12144
rect 864 12112 904 12144
rect 936 12112 976 12144
rect 1008 12112 1048 12144
rect 1080 12112 1120 12144
rect 1152 12112 1192 12144
rect 1224 12112 1264 12144
rect 1296 12112 1336 12144
rect 1368 12112 1408 12144
rect 1440 12112 1480 12144
rect 1512 12112 1552 12144
rect 1584 12112 1624 12144
rect 1656 12112 1696 12144
rect 1728 12112 1768 12144
rect 1800 12112 1840 12144
rect 1872 12112 1912 12144
rect 1944 12112 1984 12144
rect 2016 12112 2056 12144
rect 2088 12112 2128 12144
rect 2160 12112 2200 12144
rect 2232 12112 2272 12144
rect 2304 12112 2344 12144
rect 2376 12112 2416 12144
rect 2448 12112 2488 12144
rect 2520 12112 2560 12144
rect 2592 12112 2632 12144
rect 2664 12112 2704 12144
rect 2736 12112 2776 12144
rect 2808 12112 2848 12144
rect 2880 12112 2920 12144
rect 2952 12112 2992 12144
rect 3024 12112 3064 12144
rect 3096 12112 3136 12144
rect 3168 12112 3208 12144
rect 3240 12112 3280 12144
rect 3312 12112 3352 12144
rect 3384 12112 3424 12144
rect 3456 12112 3496 12144
rect 3528 12112 3568 12144
rect 3600 12112 3640 12144
rect 3672 12112 3712 12144
rect 3744 12112 3784 12144
rect 3816 12112 3856 12144
rect 3888 12112 3928 12144
rect 3960 12112 4000 12144
rect 0 12072 4000 12112
rect 0 12040 40 12072
rect 72 12040 112 12072
rect 144 12040 184 12072
rect 216 12040 256 12072
rect 288 12040 328 12072
rect 360 12040 400 12072
rect 432 12040 472 12072
rect 504 12040 544 12072
rect 576 12040 616 12072
rect 648 12040 688 12072
rect 720 12040 760 12072
rect 792 12040 832 12072
rect 864 12040 904 12072
rect 936 12040 976 12072
rect 1008 12040 1048 12072
rect 1080 12040 1120 12072
rect 1152 12040 1192 12072
rect 1224 12040 1264 12072
rect 1296 12040 1336 12072
rect 1368 12040 1408 12072
rect 1440 12040 1480 12072
rect 1512 12040 1552 12072
rect 1584 12040 1624 12072
rect 1656 12040 1696 12072
rect 1728 12040 1768 12072
rect 1800 12040 1840 12072
rect 1872 12040 1912 12072
rect 1944 12040 1984 12072
rect 2016 12040 2056 12072
rect 2088 12040 2128 12072
rect 2160 12040 2200 12072
rect 2232 12040 2272 12072
rect 2304 12040 2344 12072
rect 2376 12040 2416 12072
rect 2448 12040 2488 12072
rect 2520 12040 2560 12072
rect 2592 12040 2632 12072
rect 2664 12040 2704 12072
rect 2736 12040 2776 12072
rect 2808 12040 2848 12072
rect 2880 12040 2920 12072
rect 2952 12040 2992 12072
rect 3024 12040 3064 12072
rect 3096 12040 3136 12072
rect 3168 12040 3208 12072
rect 3240 12040 3280 12072
rect 3312 12040 3352 12072
rect 3384 12040 3424 12072
rect 3456 12040 3496 12072
rect 3528 12040 3568 12072
rect 3600 12040 3640 12072
rect 3672 12040 3712 12072
rect 3744 12040 3784 12072
rect 3816 12040 3856 12072
rect 3888 12040 3928 12072
rect 3960 12040 4000 12072
rect 0 12000 4000 12040
rect 0 11968 40 12000
rect 72 11968 112 12000
rect 144 11968 184 12000
rect 216 11968 256 12000
rect 288 11968 328 12000
rect 360 11968 400 12000
rect 432 11968 472 12000
rect 504 11968 544 12000
rect 576 11968 616 12000
rect 648 11968 688 12000
rect 720 11968 760 12000
rect 792 11968 832 12000
rect 864 11968 904 12000
rect 936 11968 976 12000
rect 1008 11968 1048 12000
rect 1080 11968 1120 12000
rect 1152 11968 1192 12000
rect 1224 11968 1264 12000
rect 1296 11968 1336 12000
rect 1368 11968 1408 12000
rect 1440 11968 1480 12000
rect 1512 11968 1552 12000
rect 1584 11968 1624 12000
rect 1656 11968 1696 12000
rect 1728 11968 1768 12000
rect 1800 11968 1840 12000
rect 1872 11968 1912 12000
rect 1944 11968 1984 12000
rect 2016 11968 2056 12000
rect 2088 11968 2128 12000
rect 2160 11968 2200 12000
rect 2232 11968 2272 12000
rect 2304 11968 2344 12000
rect 2376 11968 2416 12000
rect 2448 11968 2488 12000
rect 2520 11968 2560 12000
rect 2592 11968 2632 12000
rect 2664 11968 2704 12000
rect 2736 11968 2776 12000
rect 2808 11968 2848 12000
rect 2880 11968 2920 12000
rect 2952 11968 2992 12000
rect 3024 11968 3064 12000
rect 3096 11968 3136 12000
rect 3168 11968 3208 12000
rect 3240 11968 3280 12000
rect 3312 11968 3352 12000
rect 3384 11968 3424 12000
rect 3456 11968 3496 12000
rect 3528 11968 3568 12000
rect 3600 11968 3640 12000
rect 3672 11968 3712 12000
rect 3744 11968 3784 12000
rect 3816 11968 3856 12000
rect 3888 11968 3928 12000
rect 3960 11968 4000 12000
rect 0 11928 4000 11968
rect 0 11896 40 11928
rect 72 11896 112 11928
rect 144 11896 184 11928
rect 216 11896 256 11928
rect 288 11896 328 11928
rect 360 11896 400 11928
rect 432 11896 472 11928
rect 504 11896 544 11928
rect 576 11896 616 11928
rect 648 11896 688 11928
rect 720 11896 760 11928
rect 792 11896 832 11928
rect 864 11896 904 11928
rect 936 11896 976 11928
rect 1008 11896 1048 11928
rect 1080 11896 1120 11928
rect 1152 11896 1192 11928
rect 1224 11896 1264 11928
rect 1296 11896 1336 11928
rect 1368 11896 1408 11928
rect 1440 11896 1480 11928
rect 1512 11896 1552 11928
rect 1584 11896 1624 11928
rect 1656 11896 1696 11928
rect 1728 11896 1768 11928
rect 1800 11896 1840 11928
rect 1872 11896 1912 11928
rect 1944 11896 1984 11928
rect 2016 11896 2056 11928
rect 2088 11896 2128 11928
rect 2160 11896 2200 11928
rect 2232 11896 2272 11928
rect 2304 11896 2344 11928
rect 2376 11896 2416 11928
rect 2448 11896 2488 11928
rect 2520 11896 2560 11928
rect 2592 11896 2632 11928
rect 2664 11896 2704 11928
rect 2736 11896 2776 11928
rect 2808 11896 2848 11928
rect 2880 11896 2920 11928
rect 2952 11896 2992 11928
rect 3024 11896 3064 11928
rect 3096 11896 3136 11928
rect 3168 11896 3208 11928
rect 3240 11896 3280 11928
rect 3312 11896 3352 11928
rect 3384 11896 3424 11928
rect 3456 11896 3496 11928
rect 3528 11896 3568 11928
rect 3600 11896 3640 11928
rect 3672 11896 3712 11928
rect 3744 11896 3784 11928
rect 3816 11896 3856 11928
rect 3888 11896 3928 11928
rect 3960 11896 4000 11928
rect 0 11856 4000 11896
rect 0 11824 40 11856
rect 72 11824 112 11856
rect 144 11824 184 11856
rect 216 11824 256 11856
rect 288 11824 328 11856
rect 360 11824 400 11856
rect 432 11824 472 11856
rect 504 11824 544 11856
rect 576 11824 616 11856
rect 648 11824 688 11856
rect 720 11824 760 11856
rect 792 11824 832 11856
rect 864 11824 904 11856
rect 936 11824 976 11856
rect 1008 11824 1048 11856
rect 1080 11824 1120 11856
rect 1152 11824 1192 11856
rect 1224 11824 1264 11856
rect 1296 11824 1336 11856
rect 1368 11824 1408 11856
rect 1440 11824 1480 11856
rect 1512 11824 1552 11856
rect 1584 11824 1624 11856
rect 1656 11824 1696 11856
rect 1728 11824 1768 11856
rect 1800 11824 1840 11856
rect 1872 11824 1912 11856
rect 1944 11824 1984 11856
rect 2016 11824 2056 11856
rect 2088 11824 2128 11856
rect 2160 11824 2200 11856
rect 2232 11824 2272 11856
rect 2304 11824 2344 11856
rect 2376 11824 2416 11856
rect 2448 11824 2488 11856
rect 2520 11824 2560 11856
rect 2592 11824 2632 11856
rect 2664 11824 2704 11856
rect 2736 11824 2776 11856
rect 2808 11824 2848 11856
rect 2880 11824 2920 11856
rect 2952 11824 2992 11856
rect 3024 11824 3064 11856
rect 3096 11824 3136 11856
rect 3168 11824 3208 11856
rect 3240 11824 3280 11856
rect 3312 11824 3352 11856
rect 3384 11824 3424 11856
rect 3456 11824 3496 11856
rect 3528 11824 3568 11856
rect 3600 11824 3640 11856
rect 3672 11824 3712 11856
rect 3744 11824 3784 11856
rect 3816 11824 3856 11856
rect 3888 11824 3928 11856
rect 3960 11824 4000 11856
rect 0 11784 4000 11824
rect 0 11752 40 11784
rect 72 11752 112 11784
rect 144 11752 184 11784
rect 216 11752 256 11784
rect 288 11752 328 11784
rect 360 11752 400 11784
rect 432 11752 472 11784
rect 504 11752 544 11784
rect 576 11752 616 11784
rect 648 11752 688 11784
rect 720 11752 760 11784
rect 792 11752 832 11784
rect 864 11752 904 11784
rect 936 11752 976 11784
rect 1008 11752 1048 11784
rect 1080 11752 1120 11784
rect 1152 11752 1192 11784
rect 1224 11752 1264 11784
rect 1296 11752 1336 11784
rect 1368 11752 1408 11784
rect 1440 11752 1480 11784
rect 1512 11752 1552 11784
rect 1584 11752 1624 11784
rect 1656 11752 1696 11784
rect 1728 11752 1768 11784
rect 1800 11752 1840 11784
rect 1872 11752 1912 11784
rect 1944 11752 1984 11784
rect 2016 11752 2056 11784
rect 2088 11752 2128 11784
rect 2160 11752 2200 11784
rect 2232 11752 2272 11784
rect 2304 11752 2344 11784
rect 2376 11752 2416 11784
rect 2448 11752 2488 11784
rect 2520 11752 2560 11784
rect 2592 11752 2632 11784
rect 2664 11752 2704 11784
rect 2736 11752 2776 11784
rect 2808 11752 2848 11784
rect 2880 11752 2920 11784
rect 2952 11752 2992 11784
rect 3024 11752 3064 11784
rect 3096 11752 3136 11784
rect 3168 11752 3208 11784
rect 3240 11752 3280 11784
rect 3312 11752 3352 11784
rect 3384 11752 3424 11784
rect 3456 11752 3496 11784
rect 3528 11752 3568 11784
rect 3600 11752 3640 11784
rect 3672 11752 3712 11784
rect 3744 11752 3784 11784
rect 3816 11752 3856 11784
rect 3888 11752 3928 11784
rect 3960 11752 4000 11784
rect 0 11712 4000 11752
rect 0 11680 40 11712
rect 72 11680 112 11712
rect 144 11680 184 11712
rect 216 11680 256 11712
rect 288 11680 328 11712
rect 360 11680 400 11712
rect 432 11680 472 11712
rect 504 11680 544 11712
rect 576 11680 616 11712
rect 648 11680 688 11712
rect 720 11680 760 11712
rect 792 11680 832 11712
rect 864 11680 904 11712
rect 936 11680 976 11712
rect 1008 11680 1048 11712
rect 1080 11680 1120 11712
rect 1152 11680 1192 11712
rect 1224 11680 1264 11712
rect 1296 11680 1336 11712
rect 1368 11680 1408 11712
rect 1440 11680 1480 11712
rect 1512 11680 1552 11712
rect 1584 11680 1624 11712
rect 1656 11680 1696 11712
rect 1728 11680 1768 11712
rect 1800 11680 1840 11712
rect 1872 11680 1912 11712
rect 1944 11680 1984 11712
rect 2016 11680 2056 11712
rect 2088 11680 2128 11712
rect 2160 11680 2200 11712
rect 2232 11680 2272 11712
rect 2304 11680 2344 11712
rect 2376 11680 2416 11712
rect 2448 11680 2488 11712
rect 2520 11680 2560 11712
rect 2592 11680 2632 11712
rect 2664 11680 2704 11712
rect 2736 11680 2776 11712
rect 2808 11680 2848 11712
rect 2880 11680 2920 11712
rect 2952 11680 2992 11712
rect 3024 11680 3064 11712
rect 3096 11680 3136 11712
rect 3168 11680 3208 11712
rect 3240 11680 3280 11712
rect 3312 11680 3352 11712
rect 3384 11680 3424 11712
rect 3456 11680 3496 11712
rect 3528 11680 3568 11712
rect 3600 11680 3640 11712
rect 3672 11680 3712 11712
rect 3744 11680 3784 11712
rect 3816 11680 3856 11712
rect 3888 11680 3928 11712
rect 3960 11680 4000 11712
rect 0 11640 4000 11680
rect 0 11608 40 11640
rect 72 11608 112 11640
rect 144 11608 184 11640
rect 216 11608 256 11640
rect 288 11608 328 11640
rect 360 11608 400 11640
rect 432 11608 472 11640
rect 504 11608 544 11640
rect 576 11608 616 11640
rect 648 11608 688 11640
rect 720 11608 760 11640
rect 792 11608 832 11640
rect 864 11608 904 11640
rect 936 11608 976 11640
rect 1008 11608 1048 11640
rect 1080 11608 1120 11640
rect 1152 11608 1192 11640
rect 1224 11608 1264 11640
rect 1296 11608 1336 11640
rect 1368 11608 1408 11640
rect 1440 11608 1480 11640
rect 1512 11608 1552 11640
rect 1584 11608 1624 11640
rect 1656 11608 1696 11640
rect 1728 11608 1768 11640
rect 1800 11608 1840 11640
rect 1872 11608 1912 11640
rect 1944 11608 1984 11640
rect 2016 11608 2056 11640
rect 2088 11608 2128 11640
rect 2160 11608 2200 11640
rect 2232 11608 2272 11640
rect 2304 11608 2344 11640
rect 2376 11608 2416 11640
rect 2448 11608 2488 11640
rect 2520 11608 2560 11640
rect 2592 11608 2632 11640
rect 2664 11608 2704 11640
rect 2736 11608 2776 11640
rect 2808 11608 2848 11640
rect 2880 11608 2920 11640
rect 2952 11608 2992 11640
rect 3024 11608 3064 11640
rect 3096 11608 3136 11640
rect 3168 11608 3208 11640
rect 3240 11608 3280 11640
rect 3312 11608 3352 11640
rect 3384 11608 3424 11640
rect 3456 11608 3496 11640
rect 3528 11608 3568 11640
rect 3600 11608 3640 11640
rect 3672 11608 3712 11640
rect 3744 11608 3784 11640
rect 3816 11608 3856 11640
rect 3888 11608 3928 11640
rect 3960 11608 4000 11640
rect 0 11568 4000 11608
rect 0 11536 40 11568
rect 72 11536 112 11568
rect 144 11536 184 11568
rect 216 11536 256 11568
rect 288 11536 328 11568
rect 360 11536 400 11568
rect 432 11536 472 11568
rect 504 11536 544 11568
rect 576 11536 616 11568
rect 648 11536 688 11568
rect 720 11536 760 11568
rect 792 11536 832 11568
rect 864 11536 904 11568
rect 936 11536 976 11568
rect 1008 11536 1048 11568
rect 1080 11536 1120 11568
rect 1152 11536 1192 11568
rect 1224 11536 1264 11568
rect 1296 11536 1336 11568
rect 1368 11536 1408 11568
rect 1440 11536 1480 11568
rect 1512 11536 1552 11568
rect 1584 11536 1624 11568
rect 1656 11536 1696 11568
rect 1728 11536 1768 11568
rect 1800 11536 1840 11568
rect 1872 11536 1912 11568
rect 1944 11536 1984 11568
rect 2016 11536 2056 11568
rect 2088 11536 2128 11568
rect 2160 11536 2200 11568
rect 2232 11536 2272 11568
rect 2304 11536 2344 11568
rect 2376 11536 2416 11568
rect 2448 11536 2488 11568
rect 2520 11536 2560 11568
rect 2592 11536 2632 11568
rect 2664 11536 2704 11568
rect 2736 11536 2776 11568
rect 2808 11536 2848 11568
rect 2880 11536 2920 11568
rect 2952 11536 2992 11568
rect 3024 11536 3064 11568
rect 3096 11536 3136 11568
rect 3168 11536 3208 11568
rect 3240 11536 3280 11568
rect 3312 11536 3352 11568
rect 3384 11536 3424 11568
rect 3456 11536 3496 11568
rect 3528 11536 3568 11568
rect 3600 11536 3640 11568
rect 3672 11536 3712 11568
rect 3744 11536 3784 11568
rect 3816 11536 3856 11568
rect 3888 11536 3928 11568
rect 3960 11536 4000 11568
rect 0 11496 4000 11536
rect 0 11464 40 11496
rect 72 11464 112 11496
rect 144 11464 184 11496
rect 216 11464 256 11496
rect 288 11464 328 11496
rect 360 11464 400 11496
rect 432 11464 472 11496
rect 504 11464 544 11496
rect 576 11464 616 11496
rect 648 11464 688 11496
rect 720 11464 760 11496
rect 792 11464 832 11496
rect 864 11464 904 11496
rect 936 11464 976 11496
rect 1008 11464 1048 11496
rect 1080 11464 1120 11496
rect 1152 11464 1192 11496
rect 1224 11464 1264 11496
rect 1296 11464 1336 11496
rect 1368 11464 1408 11496
rect 1440 11464 1480 11496
rect 1512 11464 1552 11496
rect 1584 11464 1624 11496
rect 1656 11464 1696 11496
rect 1728 11464 1768 11496
rect 1800 11464 1840 11496
rect 1872 11464 1912 11496
rect 1944 11464 1984 11496
rect 2016 11464 2056 11496
rect 2088 11464 2128 11496
rect 2160 11464 2200 11496
rect 2232 11464 2272 11496
rect 2304 11464 2344 11496
rect 2376 11464 2416 11496
rect 2448 11464 2488 11496
rect 2520 11464 2560 11496
rect 2592 11464 2632 11496
rect 2664 11464 2704 11496
rect 2736 11464 2776 11496
rect 2808 11464 2848 11496
rect 2880 11464 2920 11496
rect 2952 11464 2992 11496
rect 3024 11464 3064 11496
rect 3096 11464 3136 11496
rect 3168 11464 3208 11496
rect 3240 11464 3280 11496
rect 3312 11464 3352 11496
rect 3384 11464 3424 11496
rect 3456 11464 3496 11496
rect 3528 11464 3568 11496
rect 3600 11464 3640 11496
rect 3672 11464 3712 11496
rect 3744 11464 3784 11496
rect 3816 11464 3856 11496
rect 3888 11464 3928 11496
rect 3960 11464 4000 11496
rect 0 11424 4000 11464
rect 0 11392 40 11424
rect 72 11392 112 11424
rect 144 11392 184 11424
rect 216 11392 256 11424
rect 288 11392 328 11424
rect 360 11392 400 11424
rect 432 11392 472 11424
rect 504 11392 544 11424
rect 576 11392 616 11424
rect 648 11392 688 11424
rect 720 11392 760 11424
rect 792 11392 832 11424
rect 864 11392 904 11424
rect 936 11392 976 11424
rect 1008 11392 1048 11424
rect 1080 11392 1120 11424
rect 1152 11392 1192 11424
rect 1224 11392 1264 11424
rect 1296 11392 1336 11424
rect 1368 11392 1408 11424
rect 1440 11392 1480 11424
rect 1512 11392 1552 11424
rect 1584 11392 1624 11424
rect 1656 11392 1696 11424
rect 1728 11392 1768 11424
rect 1800 11392 1840 11424
rect 1872 11392 1912 11424
rect 1944 11392 1984 11424
rect 2016 11392 2056 11424
rect 2088 11392 2128 11424
rect 2160 11392 2200 11424
rect 2232 11392 2272 11424
rect 2304 11392 2344 11424
rect 2376 11392 2416 11424
rect 2448 11392 2488 11424
rect 2520 11392 2560 11424
rect 2592 11392 2632 11424
rect 2664 11392 2704 11424
rect 2736 11392 2776 11424
rect 2808 11392 2848 11424
rect 2880 11392 2920 11424
rect 2952 11392 2992 11424
rect 3024 11392 3064 11424
rect 3096 11392 3136 11424
rect 3168 11392 3208 11424
rect 3240 11392 3280 11424
rect 3312 11392 3352 11424
rect 3384 11392 3424 11424
rect 3456 11392 3496 11424
rect 3528 11392 3568 11424
rect 3600 11392 3640 11424
rect 3672 11392 3712 11424
rect 3744 11392 3784 11424
rect 3816 11392 3856 11424
rect 3888 11392 3928 11424
rect 3960 11392 4000 11424
rect 0 11352 4000 11392
rect 0 11320 40 11352
rect 72 11320 112 11352
rect 144 11320 184 11352
rect 216 11320 256 11352
rect 288 11320 328 11352
rect 360 11320 400 11352
rect 432 11320 472 11352
rect 504 11320 544 11352
rect 576 11320 616 11352
rect 648 11320 688 11352
rect 720 11320 760 11352
rect 792 11320 832 11352
rect 864 11320 904 11352
rect 936 11320 976 11352
rect 1008 11320 1048 11352
rect 1080 11320 1120 11352
rect 1152 11320 1192 11352
rect 1224 11320 1264 11352
rect 1296 11320 1336 11352
rect 1368 11320 1408 11352
rect 1440 11320 1480 11352
rect 1512 11320 1552 11352
rect 1584 11320 1624 11352
rect 1656 11320 1696 11352
rect 1728 11320 1768 11352
rect 1800 11320 1840 11352
rect 1872 11320 1912 11352
rect 1944 11320 1984 11352
rect 2016 11320 2056 11352
rect 2088 11320 2128 11352
rect 2160 11320 2200 11352
rect 2232 11320 2272 11352
rect 2304 11320 2344 11352
rect 2376 11320 2416 11352
rect 2448 11320 2488 11352
rect 2520 11320 2560 11352
rect 2592 11320 2632 11352
rect 2664 11320 2704 11352
rect 2736 11320 2776 11352
rect 2808 11320 2848 11352
rect 2880 11320 2920 11352
rect 2952 11320 2992 11352
rect 3024 11320 3064 11352
rect 3096 11320 3136 11352
rect 3168 11320 3208 11352
rect 3240 11320 3280 11352
rect 3312 11320 3352 11352
rect 3384 11320 3424 11352
rect 3456 11320 3496 11352
rect 3528 11320 3568 11352
rect 3600 11320 3640 11352
rect 3672 11320 3712 11352
rect 3744 11320 3784 11352
rect 3816 11320 3856 11352
rect 3888 11320 3928 11352
rect 3960 11320 4000 11352
rect 0 11280 4000 11320
rect 0 11248 40 11280
rect 72 11248 112 11280
rect 144 11248 184 11280
rect 216 11248 256 11280
rect 288 11248 328 11280
rect 360 11248 400 11280
rect 432 11248 472 11280
rect 504 11248 544 11280
rect 576 11248 616 11280
rect 648 11248 688 11280
rect 720 11248 760 11280
rect 792 11248 832 11280
rect 864 11248 904 11280
rect 936 11248 976 11280
rect 1008 11248 1048 11280
rect 1080 11248 1120 11280
rect 1152 11248 1192 11280
rect 1224 11248 1264 11280
rect 1296 11248 1336 11280
rect 1368 11248 1408 11280
rect 1440 11248 1480 11280
rect 1512 11248 1552 11280
rect 1584 11248 1624 11280
rect 1656 11248 1696 11280
rect 1728 11248 1768 11280
rect 1800 11248 1840 11280
rect 1872 11248 1912 11280
rect 1944 11248 1984 11280
rect 2016 11248 2056 11280
rect 2088 11248 2128 11280
rect 2160 11248 2200 11280
rect 2232 11248 2272 11280
rect 2304 11248 2344 11280
rect 2376 11248 2416 11280
rect 2448 11248 2488 11280
rect 2520 11248 2560 11280
rect 2592 11248 2632 11280
rect 2664 11248 2704 11280
rect 2736 11248 2776 11280
rect 2808 11248 2848 11280
rect 2880 11248 2920 11280
rect 2952 11248 2992 11280
rect 3024 11248 3064 11280
rect 3096 11248 3136 11280
rect 3168 11248 3208 11280
rect 3240 11248 3280 11280
rect 3312 11248 3352 11280
rect 3384 11248 3424 11280
rect 3456 11248 3496 11280
rect 3528 11248 3568 11280
rect 3600 11248 3640 11280
rect 3672 11248 3712 11280
rect 3744 11248 3784 11280
rect 3816 11248 3856 11280
rect 3888 11248 3928 11280
rect 3960 11248 4000 11280
rect 0 11208 4000 11248
rect 0 11176 40 11208
rect 72 11176 112 11208
rect 144 11176 184 11208
rect 216 11176 256 11208
rect 288 11176 328 11208
rect 360 11176 400 11208
rect 432 11176 472 11208
rect 504 11176 544 11208
rect 576 11176 616 11208
rect 648 11176 688 11208
rect 720 11176 760 11208
rect 792 11176 832 11208
rect 864 11176 904 11208
rect 936 11176 976 11208
rect 1008 11176 1048 11208
rect 1080 11176 1120 11208
rect 1152 11176 1192 11208
rect 1224 11176 1264 11208
rect 1296 11176 1336 11208
rect 1368 11176 1408 11208
rect 1440 11176 1480 11208
rect 1512 11176 1552 11208
rect 1584 11176 1624 11208
rect 1656 11176 1696 11208
rect 1728 11176 1768 11208
rect 1800 11176 1840 11208
rect 1872 11176 1912 11208
rect 1944 11176 1984 11208
rect 2016 11176 2056 11208
rect 2088 11176 2128 11208
rect 2160 11176 2200 11208
rect 2232 11176 2272 11208
rect 2304 11176 2344 11208
rect 2376 11176 2416 11208
rect 2448 11176 2488 11208
rect 2520 11176 2560 11208
rect 2592 11176 2632 11208
rect 2664 11176 2704 11208
rect 2736 11176 2776 11208
rect 2808 11176 2848 11208
rect 2880 11176 2920 11208
rect 2952 11176 2992 11208
rect 3024 11176 3064 11208
rect 3096 11176 3136 11208
rect 3168 11176 3208 11208
rect 3240 11176 3280 11208
rect 3312 11176 3352 11208
rect 3384 11176 3424 11208
rect 3456 11176 3496 11208
rect 3528 11176 3568 11208
rect 3600 11176 3640 11208
rect 3672 11176 3712 11208
rect 3744 11176 3784 11208
rect 3816 11176 3856 11208
rect 3888 11176 3928 11208
rect 3960 11176 4000 11208
rect 0 11136 4000 11176
rect 0 11104 40 11136
rect 72 11104 112 11136
rect 144 11104 184 11136
rect 216 11104 256 11136
rect 288 11104 328 11136
rect 360 11104 400 11136
rect 432 11104 472 11136
rect 504 11104 544 11136
rect 576 11104 616 11136
rect 648 11104 688 11136
rect 720 11104 760 11136
rect 792 11104 832 11136
rect 864 11104 904 11136
rect 936 11104 976 11136
rect 1008 11104 1048 11136
rect 1080 11104 1120 11136
rect 1152 11104 1192 11136
rect 1224 11104 1264 11136
rect 1296 11104 1336 11136
rect 1368 11104 1408 11136
rect 1440 11104 1480 11136
rect 1512 11104 1552 11136
rect 1584 11104 1624 11136
rect 1656 11104 1696 11136
rect 1728 11104 1768 11136
rect 1800 11104 1840 11136
rect 1872 11104 1912 11136
rect 1944 11104 1984 11136
rect 2016 11104 2056 11136
rect 2088 11104 2128 11136
rect 2160 11104 2200 11136
rect 2232 11104 2272 11136
rect 2304 11104 2344 11136
rect 2376 11104 2416 11136
rect 2448 11104 2488 11136
rect 2520 11104 2560 11136
rect 2592 11104 2632 11136
rect 2664 11104 2704 11136
rect 2736 11104 2776 11136
rect 2808 11104 2848 11136
rect 2880 11104 2920 11136
rect 2952 11104 2992 11136
rect 3024 11104 3064 11136
rect 3096 11104 3136 11136
rect 3168 11104 3208 11136
rect 3240 11104 3280 11136
rect 3312 11104 3352 11136
rect 3384 11104 3424 11136
rect 3456 11104 3496 11136
rect 3528 11104 3568 11136
rect 3600 11104 3640 11136
rect 3672 11104 3712 11136
rect 3744 11104 3784 11136
rect 3816 11104 3856 11136
rect 3888 11104 3928 11136
rect 3960 11104 4000 11136
rect 0 11064 4000 11104
rect 0 11032 40 11064
rect 72 11032 112 11064
rect 144 11032 184 11064
rect 216 11032 256 11064
rect 288 11032 328 11064
rect 360 11032 400 11064
rect 432 11032 472 11064
rect 504 11032 544 11064
rect 576 11032 616 11064
rect 648 11032 688 11064
rect 720 11032 760 11064
rect 792 11032 832 11064
rect 864 11032 904 11064
rect 936 11032 976 11064
rect 1008 11032 1048 11064
rect 1080 11032 1120 11064
rect 1152 11032 1192 11064
rect 1224 11032 1264 11064
rect 1296 11032 1336 11064
rect 1368 11032 1408 11064
rect 1440 11032 1480 11064
rect 1512 11032 1552 11064
rect 1584 11032 1624 11064
rect 1656 11032 1696 11064
rect 1728 11032 1768 11064
rect 1800 11032 1840 11064
rect 1872 11032 1912 11064
rect 1944 11032 1984 11064
rect 2016 11032 2056 11064
rect 2088 11032 2128 11064
rect 2160 11032 2200 11064
rect 2232 11032 2272 11064
rect 2304 11032 2344 11064
rect 2376 11032 2416 11064
rect 2448 11032 2488 11064
rect 2520 11032 2560 11064
rect 2592 11032 2632 11064
rect 2664 11032 2704 11064
rect 2736 11032 2776 11064
rect 2808 11032 2848 11064
rect 2880 11032 2920 11064
rect 2952 11032 2992 11064
rect 3024 11032 3064 11064
rect 3096 11032 3136 11064
rect 3168 11032 3208 11064
rect 3240 11032 3280 11064
rect 3312 11032 3352 11064
rect 3384 11032 3424 11064
rect 3456 11032 3496 11064
rect 3528 11032 3568 11064
rect 3600 11032 3640 11064
rect 3672 11032 3712 11064
rect 3744 11032 3784 11064
rect 3816 11032 3856 11064
rect 3888 11032 3928 11064
rect 3960 11032 4000 11064
rect 0 10992 4000 11032
rect 0 10960 40 10992
rect 72 10960 112 10992
rect 144 10960 184 10992
rect 216 10960 256 10992
rect 288 10960 328 10992
rect 360 10960 400 10992
rect 432 10960 472 10992
rect 504 10960 544 10992
rect 576 10960 616 10992
rect 648 10960 688 10992
rect 720 10960 760 10992
rect 792 10960 832 10992
rect 864 10960 904 10992
rect 936 10960 976 10992
rect 1008 10960 1048 10992
rect 1080 10960 1120 10992
rect 1152 10960 1192 10992
rect 1224 10960 1264 10992
rect 1296 10960 1336 10992
rect 1368 10960 1408 10992
rect 1440 10960 1480 10992
rect 1512 10960 1552 10992
rect 1584 10960 1624 10992
rect 1656 10960 1696 10992
rect 1728 10960 1768 10992
rect 1800 10960 1840 10992
rect 1872 10960 1912 10992
rect 1944 10960 1984 10992
rect 2016 10960 2056 10992
rect 2088 10960 2128 10992
rect 2160 10960 2200 10992
rect 2232 10960 2272 10992
rect 2304 10960 2344 10992
rect 2376 10960 2416 10992
rect 2448 10960 2488 10992
rect 2520 10960 2560 10992
rect 2592 10960 2632 10992
rect 2664 10960 2704 10992
rect 2736 10960 2776 10992
rect 2808 10960 2848 10992
rect 2880 10960 2920 10992
rect 2952 10960 2992 10992
rect 3024 10960 3064 10992
rect 3096 10960 3136 10992
rect 3168 10960 3208 10992
rect 3240 10960 3280 10992
rect 3312 10960 3352 10992
rect 3384 10960 3424 10992
rect 3456 10960 3496 10992
rect 3528 10960 3568 10992
rect 3600 10960 3640 10992
rect 3672 10960 3712 10992
rect 3744 10960 3784 10992
rect 3816 10960 3856 10992
rect 3888 10960 3928 10992
rect 3960 10960 4000 10992
rect 0 10920 4000 10960
rect 0 10888 40 10920
rect 72 10888 112 10920
rect 144 10888 184 10920
rect 216 10888 256 10920
rect 288 10888 328 10920
rect 360 10888 400 10920
rect 432 10888 472 10920
rect 504 10888 544 10920
rect 576 10888 616 10920
rect 648 10888 688 10920
rect 720 10888 760 10920
rect 792 10888 832 10920
rect 864 10888 904 10920
rect 936 10888 976 10920
rect 1008 10888 1048 10920
rect 1080 10888 1120 10920
rect 1152 10888 1192 10920
rect 1224 10888 1264 10920
rect 1296 10888 1336 10920
rect 1368 10888 1408 10920
rect 1440 10888 1480 10920
rect 1512 10888 1552 10920
rect 1584 10888 1624 10920
rect 1656 10888 1696 10920
rect 1728 10888 1768 10920
rect 1800 10888 1840 10920
rect 1872 10888 1912 10920
rect 1944 10888 1984 10920
rect 2016 10888 2056 10920
rect 2088 10888 2128 10920
rect 2160 10888 2200 10920
rect 2232 10888 2272 10920
rect 2304 10888 2344 10920
rect 2376 10888 2416 10920
rect 2448 10888 2488 10920
rect 2520 10888 2560 10920
rect 2592 10888 2632 10920
rect 2664 10888 2704 10920
rect 2736 10888 2776 10920
rect 2808 10888 2848 10920
rect 2880 10888 2920 10920
rect 2952 10888 2992 10920
rect 3024 10888 3064 10920
rect 3096 10888 3136 10920
rect 3168 10888 3208 10920
rect 3240 10888 3280 10920
rect 3312 10888 3352 10920
rect 3384 10888 3424 10920
rect 3456 10888 3496 10920
rect 3528 10888 3568 10920
rect 3600 10888 3640 10920
rect 3672 10888 3712 10920
rect 3744 10888 3784 10920
rect 3816 10888 3856 10920
rect 3888 10888 3928 10920
rect 3960 10888 4000 10920
rect 0 10848 4000 10888
rect 0 10816 40 10848
rect 72 10816 112 10848
rect 144 10816 184 10848
rect 216 10816 256 10848
rect 288 10816 328 10848
rect 360 10816 400 10848
rect 432 10816 472 10848
rect 504 10816 544 10848
rect 576 10816 616 10848
rect 648 10816 688 10848
rect 720 10816 760 10848
rect 792 10816 832 10848
rect 864 10816 904 10848
rect 936 10816 976 10848
rect 1008 10816 1048 10848
rect 1080 10816 1120 10848
rect 1152 10816 1192 10848
rect 1224 10816 1264 10848
rect 1296 10816 1336 10848
rect 1368 10816 1408 10848
rect 1440 10816 1480 10848
rect 1512 10816 1552 10848
rect 1584 10816 1624 10848
rect 1656 10816 1696 10848
rect 1728 10816 1768 10848
rect 1800 10816 1840 10848
rect 1872 10816 1912 10848
rect 1944 10816 1984 10848
rect 2016 10816 2056 10848
rect 2088 10816 2128 10848
rect 2160 10816 2200 10848
rect 2232 10816 2272 10848
rect 2304 10816 2344 10848
rect 2376 10816 2416 10848
rect 2448 10816 2488 10848
rect 2520 10816 2560 10848
rect 2592 10816 2632 10848
rect 2664 10816 2704 10848
rect 2736 10816 2776 10848
rect 2808 10816 2848 10848
rect 2880 10816 2920 10848
rect 2952 10816 2992 10848
rect 3024 10816 3064 10848
rect 3096 10816 3136 10848
rect 3168 10816 3208 10848
rect 3240 10816 3280 10848
rect 3312 10816 3352 10848
rect 3384 10816 3424 10848
rect 3456 10816 3496 10848
rect 3528 10816 3568 10848
rect 3600 10816 3640 10848
rect 3672 10816 3712 10848
rect 3744 10816 3784 10848
rect 3816 10816 3856 10848
rect 3888 10816 3928 10848
rect 3960 10816 4000 10848
rect 0 10776 4000 10816
rect 0 10744 40 10776
rect 72 10744 112 10776
rect 144 10744 184 10776
rect 216 10744 256 10776
rect 288 10744 328 10776
rect 360 10744 400 10776
rect 432 10744 472 10776
rect 504 10744 544 10776
rect 576 10744 616 10776
rect 648 10744 688 10776
rect 720 10744 760 10776
rect 792 10744 832 10776
rect 864 10744 904 10776
rect 936 10744 976 10776
rect 1008 10744 1048 10776
rect 1080 10744 1120 10776
rect 1152 10744 1192 10776
rect 1224 10744 1264 10776
rect 1296 10744 1336 10776
rect 1368 10744 1408 10776
rect 1440 10744 1480 10776
rect 1512 10744 1552 10776
rect 1584 10744 1624 10776
rect 1656 10744 1696 10776
rect 1728 10744 1768 10776
rect 1800 10744 1840 10776
rect 1872 10744 1912 10776
rect 1944 10744 1984 10776
rect 2016 10744 2056 10776
rect 2088 10744 2128 10776
rect 2160 10744 2200 10776
rect 2232 10744 2272 10776
rect 2304 10744 2344 10776
rect 2376 10744 2416 10776
rect 2448 10744 2488 10776
rect 2520 10744 2560 10776
rect 2592 10744 2632 10776
rect 2664 10744 2704 10776
rect 2736 10744 2776 10776
rect 2808 10744 2848 10776
rect 2880 10744 2920 10776
rect 2952 10744 2992 10776
rect 3024 10744 3064 10776
rect 3096 10744 3136 10776
rect 3168 10744 3208 10776
rect 3240 10744 3280 10776
rect 3312 10744 3352 10776
rect 3384 10744 3424 10776
rect 3456 10744 3496 10776
rect 3528 10744 3568 10776
rect 3600 10744 3640 10776
rect 3672 10744 3712 10776
rect 3744 10744 3784 10776
rect 3816 10744 3856 10776
rect 3888 10744 3928 10776
rect 3960 10744 4000 10776
rect 0 10704 4000 10744
rect 0 10672 40 10704
rect 72 10672 112 10704
rect 144 10672 184 10704
rect 216 10672 256 10704
rect 288 10672 328 10704
rect 360 10672 400 10704
rect 432 10672 472 10704
rect 504 10672 544 10704
rect 576 10672 616 10704
rect 648 10672 688 10704
rect 720 10672 760 10704
rect 792 10672 832 10704
rect 864 10672 904 10704
rect 936 10672 976 10704
rect 1008 10672 1048 10704
rect 1080 10672 1120 10704
rect 1152 10672 1192 10704
rect 1224 10672 1264 10704
rect 1296 10672 1336 10704
rect 1368 10672 1408 10704
rect 1440 10672 1480 10704
rect 1512 10672 1552 10704
rect 1584 10672 1624 10704
rect 1656 10672 1696 10704
rect 1728 10672 1768 10704
rect 1800 10672 1840 10704
rect 1872 10672 1912 10704
rect 1944 10672 1984 10704
rect 2016 10672 2056 10704
rect 2088 10672 2128 10704
rect 2160 10672 2200 10704
rect 2232 10672 2272 10704
rect 2304 10672 2344 10704
rect 2376 10672 2416 10704
rect 2448 10672 2488 10704
rect 2520 10672 2560 10704
rect 2592 10672 2632 10704
rect 2664 10672 2704 10704
rect 2736 10672 2776 10704
rect 2808 10672 2848 10704
rect 2880 10672 2920 10704
rect 2952 10672 2992 10704
rect 3024 10672 3064 10704
rect 3096 10672 3136 10704
rect 3168 10672 3208 10704
rect 3240 10672 3280 10704
rect 3312 10672 3352 10704
rect 3384 10672 3424 10704
rect 3456 10672 3496 10704
rect 3528 10672 3568 10704
rect 3600 10672 3640 10704
rect 3672 10672 3712 10704
rect 3744 10672 3784 10704
rect 3816 10672 3856 10704
rect 3888 10672 3928 10704
rect 3960 10672 4000 10704
rect 0 10632 4000 10672
rect 0 10600 40 10632
rect 72 10600 112 10632
rect 144 10600 184 10632
rect 216 10600 256 10632
rect 288 10600 328 10632
rect 360 10600 400 10632
rect 432 10600 472 10632
rect 504 10600 544 10632
rect 576 10600 616 10632
rect 648 10600 688 10632
rect 720 10600 760 10632
rect 792 10600 832 10632
rect 864 10600 904 10632
rect 936 10600 976 10632
rect 1008 10600 1048 10632
rect 1080 10600 1120 10632
rect 1152 10600 1192 10632
rect 1224 10600 1264 10632
rect 1296 10600 1336 10632
rect 1368 10600 1408 10632
rect 1440 10600 1480 10632
rect 1512 10600 1552 10632
rect 1584 10600 1624 10632
rect 1656 10600 1696 10632
rect 1728 10600 1768 10632
rect 1800 10600 1840 10632
rect 1872 10600 1912 10632
rect 1944 10600 1984 10632
rect 2016 10600 2056 10632
rect 2088 10600 2128 10632
rect 2160 10600 2200 10632
rect 2232 10600 2272 10632
rect 2304 10600 2344 10632
rect 2376 10600 2416 10632
rect 2448 10600 2488 10632
rect 2520 10600 2560 10632
rect 2592 10600 2632 10632
rect 2664 10600 2704 10632
rect 2736 10600 2776 10632
rect 2808 10600 2848 10632
rect 2880 10600 2920 10632
rect 2952 10600 2992 10632
rect 3024 10600 3064 10632
rect 3096 10600 3136 10632
rect 3168 10600 3208 10632
rect 3240 10600 3280 10632
rect 3312 10600 3352 10632
rect 3384 10600 3424 10632
rect 3456 10600 3496 10632
rect 3528 10600 3568 10632
rect 3600 10600 3640 10632
rect 3672 10600 3712 10632
rect 3744 10600 3784 10632
rect 3816 10600 3856 10632
rect 3888 10600 3928 10632
rect 3960 10600 4000 10632
rect 0 10560 4000 10600
rect 0 10528 40 10560
rect 72 10528 112 10560
rect 144 10528 184 10560
rect 216 10528 256 10560
rect 288 10528 328 10560
rect 360 10528 400 10560
rect 432 10528 472 10560
rect 504 10528 544 10560
rect 576 10528 616 10560
rect 648 10528 688 10560
rect 720 10528 760 10560
rect 792 10528 832 10560
rect 864 10528 904 10560
rect 936 10528 976 10560
rect 1008 10528 1048 10560
rect 1080 10528 1120 10560
rect 1152 10528 1192 10560
rect 1224 10528 1264 10560
rect 1296 10528 1336 10560
rect 1368 10528 1408 10560
rect 1440 10528 1480 10560
rect 1512 10528 1552 10560
rect 1584 10528 1624 10560
rect 1656 10528 1696 10560
rect 1728 10528 1768 10560
rect 1800 10528 1840 10560
rect 1872 10528 1912 10560
rect 1944 10528 1984 10560
rect 2016 10528 2056 10560
rect 2088 10528 2128 10560
rect 2160 10528 2200 10560
rect 2232 10528 2272 10560
rect 2304 10528 2344 10560
rect 2376 10528 2416 10560
rect 2448 10528 2488 10560
rect 2520 10528 2560 10560
rect 2592 10528 2632 10560
rect 2664 10528 2704 10560
rect 2736 10528 2776 10560
rect 2808 10528 2848 10560
rect 2880 10528 2920 10560
rect 2952 10528 2992 10560
rect 3024 10528 3064 10560
rect 3096 10528 3136 10560
rect 3168 10528 3208 10560
rect 3240 10528 3280 10560
rect 3312 10528 3352 10560
rect 3384 10528 3424 10560
rect 3456 10528 3496 10560
rect 3528 10528 3568 10560
rect 3600 10528 3640 10560
rect 3672 10528 3712 10560
rect 3744 10528 3784 10560
rect 3816 10528 3856 10560
rect 3888 10528 3928 10560
rect 3960 10528 4000 10560
rect 0 10488 4000 10528
rect 0 10456 40 10488
rect 72 10456 112 10488
rect 144 10456 184 10488
rect 216 10456 256 10488
rect 288 10456 328 10488
rect 360 10456 400 10488
rect 432 10456 472 10488
rect 504 10456 544 10488
rect 576 10456 616 10488
rect 648 10456 688 10488
rect 720 10456 760 10488
rect 792 10456 832 10488
rect 864 10456 904 10488
rect 936 10456 976 10488
rect 1008 10456 1048 10488
rect 1080 10456 1120 10488
rect 1152 10456 1192 10488
rect 1224 10456 1264 10488
rect 1296 10456 1336 10488
rect 1368 10456 1408 10488
rect 1440 10456 1480 10488
rect 1512 10456 1552 10488
rect 1584 10456 1624 10488
rect 1656 10456 1696 10488
rect 1728 10456 1768 10488
rect 1800 10456 1840 10488
rect 1872 10456 1912 10488
rect 1944 10456 1984 10488
rect 2016 10456 2056 10488
rect 2088 10456 2128 10488
rect 2160 10456 2200 10488
rect 2232 10456 2272 10488
rect 2304 10456 2344 10488
rect 2376 10456 2416 10488
rect 2448 10456 2488 10488
rect 2520 10456 2560 10488
rect 2592 10456 2632 10488
rect 2664 10456 2704 10488
rect 2736 10456 2776 10488
rect 2808 10456 2848 10488
rect 2880 10456 2920 10488
rect 2952 10456 2992 10488
rect 3024 10456 3064 10488
rect 3096 10456 3136 10488
rect 3168 10456 3208 10488
rect 3240 10456 3280 10488
rect 3312 10456 3352 10488
rect 3384 10456 3424 10488
rect 3456 10456 3496 10488
rect 3528 10456 3568 10488
rect 3600 10456 3640 10488
rect 3672 10456 3712 10488
rect 3744 10456 3784 10488
rect 3816 10456 3856 10488
rect 3888 10456 3928 10488
rect 3960 10456 4000 10488
rect 0 10416 4000 10456
rect 0 10384 40 10416
rect 72 10384 112 10416
rect 144 10384 184 10416
rect 216 10384 256 10416
rect 288 10384 328 10416
rect 360 10384 400 10416
rect 432 10384 472 10416
rect 504 10384 544 10416
rect 576 10384 616 10416
rect 648 10384 688 10416
rect 720 10384 760 10416
rect 792 10384 832 10416
rect 864 10384 904 10416
rect 936 10384 976 10416
rect 1008 10384 1048 10416
rect 1080 10384 1120 10416
rect 1152 10384 1192 10416
rect 1224 10384 1264 10416
rect 1296 10384 1336 10416
rect 1368 10384 1408 10416
rect 1440 10384 1480 10416
rect 1512 10384 1552 10416
rect 1584 10384 1624 10416
rect 1656 10384 1696 10416
rect 1728 10384 1768 10416
rect 1800 10384 1840 10416
rect 1872 10384 1912 10416
rect 1944 10384 1984 10416
rect 2016 10384 2056 10416
rect 2088 10384 2128 10416
rect 2160 10384 2200 10416
rect 2232 10384 2272 10416
rect 2304 10384 2344 10416
rect 2376 10384 2416 10416
rect 2448 10384 2488 10416
rect 2520 10384 2560 10416
rect 2592 10384 2632 10416
rect 2664 10384 2704 10416
rect 2736 10384 2776 10416
rect 2808 10384 2848 10416
rect 2880 10384 2920 10416
rect 2952 10384 2992 10416
rect 3024 10384 3064 10416
rect 3096 10384 3136 10416
rect 3168 10384 3208 10416
rect 3240 10384 3280 10416
rect 3312 10384 3352 10416
rect 3384 10384 3424 10416
rect 3456 10384 3496 10416
rect 3528 10384 3568 10416
rect 3600 10384 3640 10416
rect 3672 10384 3712 10416
rect 3744 10384 3784 10416
rect 3816 10384 3856 10416
rect 3888 10384 3928 10416
rect 3960 10384 4000 10416
rect 0 10344 4000 10384
rect 0 10312 40 10344
rect 72 10312 112 10344
rect 144 10312 184 10344
rect 216 10312 256 10344
rect 288 10312 328 10344
rect 360 10312 400 10344
rect 432 10312 472 10344
rect 504 10312 544 10344
rect 576 10312 616 10344
rect 648 10312 688 10344
rect 720 10312 760 10344
rect 792 10312 832 10344
rect 864 10312 904 10344
rect 936 10312 976 10344
rect 1008 10312 1048 10344
rect 1080 10312 1120 10344
rect 1152 10312 1192 10344
rect 1224 10312 1264 10344
rect 1296 10312 1336 10344
rect 1368 10312 1408 10344
rect 1440 10312 1480 10344
rect 1512 10312 1552 10344
rect 1584 10312 1624 10344
rect 1656 10312 1696 10344
rect 1728 10312 1768 10344
rect 1800 10312 1840 10344
rect 1872 10312 1912 10344
rect 1944 10312 1984 10344
rect 2016 10312 2056 10344
rect 2088 10312 2128 10344
rect 2160 10312 2200 10344
rect 2232 10312 2272 10344
rect 2304 10312 2344 10344
rect 2376 10312 2416 10344
rect 2448 10312 2488 10344
rect 2520 10312 2560 10344
rect 2592 10312 2632 10344
rect 2664 10312 2704 10344
rect 2736 10312 2776 10344
rect 2808 10312 2848 10344
rect 2880 10312 2920 10344
rect 2952 10312 2992 10344
rect 3024 10312 3064 10344
rect 3096 10312 3136 10344
rect 3168 10312 3208 10344
rect 3240 10312 3280 10344
rect 3312 10312 3352 10344
rect 3384 10312 3424 10344
rect 3456 10312 3496 10344
rect 3528 10312 3568 10344
rect 3600 10312 3640 10344
rect 3672 10312 3712 10344
rect 3744 10312 3784 10344
rect 3816 10312 3856 10344
rect 3888 10312 3928 10344
rect 3960 10312 4000 10344
rect 0 10272 4000 10312
rect 0 10240 40 10272
rect 72 10240 112 10272
rect 144 10240 184 10272
rect 216 10240 256 10272
rect 288 10240 328 10272
rect 360 10240 400 10272
rect 432 10240 472 10272
rect 504 10240 544 10272
rect 576 10240 616 10272
rect 648 10240 688 10272
rect 720 10240 760 10272
rect 792 10240 832 10272
rect 864 10240 904 10272
rect 936 10240 976 10272
rect 1008 10240 1048 10272
rect 1080 10240 1120 10272
rect 1152 10240 1192 10272
rect 1224 10240 1264 10272
rect 1296 10240 1336 10272
rect 1368 10240 1408 10272
rect 1440 10240 1480 10272
rect 1512 10240 1552 10272
rect 1584 10240 1624 10272
rect 1656 10240 1696 10272
rect 1728 10240 1768 10272
rect 1800 10240 1840 10272
rect 1872 10240 1912 10272
rect 1944 10240 1984 10272
rect 2016 10240 2056 10272
rect 2088 10240 2128 10272
rect 2160 10240 2200 10272
rect 2232 10240 2272 10272
rect 2304 10240 2344 10272
rect 2376 10240 2416 10272
rect 2448 10240 2488 10272
rect 2520 10240 2560 10272
rect 2592 10240 2632 10272
rect 2664 10240 2704 10272
rect 2736 10240 2776 10272
rect 2808 10240 2848 10272
rect 2880 10240 2920 10272
rect 2952 10240 2992 10272
rect 3024 10240 3064 10272
rect 3096 10240 3136 10272
rect 3168 10240 3208 10272
rect 3240 10240 3280 10272
rect 3312 10240 3352 10272
rect 3384 10240 3424 10272
rect 3456 10240 3496 10272
rect 3528 10240 3568 10272
rect 3600 10240 3640 10272
rect 3672 10240 3712 10272
rect 3744 10240 3784 10272
rect 3816 10240 3856 10272
rect 3888 10240 3928 10272
rect 3960 10240 4000 10272
rect 0 10200 4000 10240
rect 0 10168 40 10200
rect 72 10168 112 10200
rect 144 10168 184 10200
rect 216 10168 256 10200
rect 288 10168 328 10200
rect 360 10168 400 10200
rect 432 10168 472 10200
rect 504 10168 544 10200
rect 576 10168 616 10200
rect 648 10168 688 10200
rect 720 10168 760 10200
rect 792 10168 832 10200
rect 864 10168 904 10200
rect 936 10168 976 10200
rect 1008 10168 1048 10200
rect 1080 10168 1120 10200
rect 1152 10168 1192 10200
rect 1224 10168 1264 10200
rect 1296 10168 1336 10200
rect 1368 10168 1408 10200
rect 1440 10168 1480 10200
rect 1512 10168 1552 10200
rect 1584 10168 1624 10200
rect 1656 10168 1696 10200
rect 1728 10168 1768 10200
rect 1800 10168 1840 10200
rect 1872 10168 1912 10200
rect 1944 10168 1984 10200
rect 2016 10168 2056 10200
rect 2088 10168 2128 10200
rect 2160 10168 2200 10200
rect 2232 10168 2272 10200
rect 2304 10168 2344 10200
rect 2376 10168 2416 10200
rect 2448 10168 2488 10200
rect 2520 10168 2560 10200
rect 2592 10168 2632 10200
rect 2664 10168 2704 10200
rect 2736 10168 2776 10200
rect 2808 10168 2848 10200
rect 2880 10168 2920 10200
rect 2952 10168 2992 10200
rect 3024 10168 3064 10200
rect 3096 10168 3136 10200
rect 3168 10168 3208 10200
rect 3240 10168 3280 10200
rect 3312 10168 3352 10200
rect 3384 10168 3424 10200
rect 3456 10168 3496 10200
rect 3528 10168 3568 10200
rect 3600 10168 3640 10200
rect 3672 10168 3712 10200
rect 3744 10168 3784 10200
rect 3816 10168 3856 10200
rect 3888 10168 3928 10200
rect 3960 10168 4000 10200
rect 0 10128 4000 10168
rect 0 10096 40 10128
rect 72 10096 112 10128
rect 144 10096 184 10128
rect 216 10096 256 10128
rect 288 10096 328 10128
rect 360 10096 400 10128
rect 432 10096 472 10128
rect 504 10096 544 10128
rect 576 10096 616 10128
rect 648 10096 688 10128
rect 720 10096 760 10128
rect 792 10096 832 10128
rect 864 10096 904 10128
rect 936 10096 976 10128
rect 1008 10096 1048 10128
rect 1080 10096 1120 10128
rect 1152 10096 1192 10128
rect 1224 10096 1264 10128
rect 1296 10096 1336 10128
rect 1368 10096 1408 10128
rect 1440 10096 1480 10128
rect 1512 10096 1552 10128
rect 1584 10096 1624 10128
rect 1656 10096 1696 10128
rect 1728 10096 1768 10128
rect 1800 10096 1840 10128
rect 1872 10096 1912 10128
rect 1944 10096 1984 10128
rect 2016 10096 2056 10128
rect 2088 10096 2128 10128
rect 2160 10096 2200 10128
rect 2232 10096 2272 10128
rect 2304 10096 2344 10128
rect 2376 10096 2416 10128
rect 2448 10096 2488 10128
rect 2520 10096 2560 10128
rect 2592 10096 2632 10128
rect 2664 10096 2704 10128
rect 2736 10096 2776 10128
rect 2808 10096 2848 10128
rect 2880 10096 2920 10128
rect 2952 10096 2992 10128
rect 3024 10096 3064 10128
rect 3096 10096 3136 10128
rect 3168 10096 3208 10128
rect 3240 10096 3280 10128
rect 3312 10096 3352 10128
rect 3384 10096 3424 10128
rect 3456 10096 3496 10128
rect 3528 10096 3568 10128
rect 3600 10096 3640 10128
rect 3672 10096 3712 10128
rect 3744 10096 3784 10128
rect 3816 10096 3856 10128
rect 3888 10096 3928 10128
rect 3960 10096 4000 10128
rect 0 10056 4000 10096
rect 0 10024 40 10056
rect 72 10024 112 10056
rect 144 10024 184 10056
rect 216 10024 256 10056
rect 288 10024 328 10056
rect 360 10024 400 10056
rect 432 10024 472 10056
rect 504 10024 544 10056
rect 576 10024 616 10056
rect 648 10024 688 10056
rect 720 10024 760 10056
rect 792 10024 832 10056
rect 864 10024 904 10056
rect 936 10024 976 10056
rect 1008 10024 1048 10056
rect 1080 10024 1120 10056
rect 1152 10024 1192 10056
rect 1224 10024 1264 10056
rect 1296 10024 1336 10056
rect 1368 10024 1408 10056
rect 1440 10024 1480 10056
rect 1512 10024 1552 10056
rect 1584 10024 1624 10056
rect 1656 10024 1696 10056
rect 1728 10024 1768 10056
rect 1800 10024 1840 10056
rect 1872 10024 1912 10056
rect 1944 10024 1984 10056
rect 2016 10024 2056 10056
rect 2088 10024 2128 10056
rect 2160 10024 2200 10056
rect 2232 10024 2272 10056
rect 2304 10024 2344 10056
rect 2376 10024 2416 10056
rect 2448 10024 2488 10056
rect 2520 10024 2560 10056
rect 2592 10024 2632 10056
rect 2664 10024 2704 10056
rect 2736 10024 2776 10056
rect 2808 10024 2848 10056
rect 2880 10024 2920 10056
rect 2952 10024 2992 10056
rect 3024 10024 3064 10056
rect 3096 10024 3136 10056
rect 3168 10024 3208 10056
rect 3240 10024 3280 10056
rect 3312 10024 3352 10056
rect 3384 10024 3424 10056
rect 3456 10024 3496 10056
rect 3528 10024 3568 10056
rect 3600 10024 3640 10056
rect 3672 10024 3712 10056
rect 3744 10024 3784 10056
rect 3816 10024 3856 10056
rect 3888 10024 3928 10056
rect 3960 10024 4000 10056
rect 0 9984 4000 10024
rect 0 9952 40 9984
rect 72 9952 112 9984
rect 144 9952 184 9984
rect 216 9952 256 9984
rect 288 9952 328 9984
rect 360 9952 400 9984
rect 432 9952 472 9984
rect 504 9952 544 9984
rect 576 9952 616 9984
rect 648 9952 688 9984
rect 720 9952 760 9984
rect 792 9952 832 9984
rect 864 9952 904 9984
rect 936 9952 976 9984
rect 1008 9952 1048 9984
rect 1080 9952 1120 9984
rect 1152 9952 1192 9984
rect 1224 9952 1264 9984
rect 1296 9952 1336 9984
rect 1368 9952 1408 9984
rect 1440 9952 1480 9984
rect 1512 9952 1552 9984
rect 1584 9952 1624 9984
rect 1656 9952 1696 9984
rect 1728 9952 1768 9984
rect 1800 9952 1840 9984
rect 1872 9952 1912 9984
rect 1944 9952 1984 9984
rect 2016 9952 2056 9984
rect 2088 9952 2128 9984
rect 2160 9952 2200 9984
rect 2232 9952 2272 9984
rect 2304 9952 2344 9984
rect 2376 9952 2416 9984
rect 2448 9952 2488 9984
rect 2520 9952 2560 9984
rect 2592 9952 2632 9984
rect 2664 9952 2704 9984
rect 2736 9952 2776 9984
rect 2808 9952 2848 9984
rect 2880 9952 2920 9984
rect 2952 9952 2992 9984
rect 3024 9952 3064 9984
rect 3096 9952 3136 9984
rect 3168 9952 3208 9984
rect 3240 9952 3280 9984
rect 3312 9952 3352 9984
rect 3384 9952 3424 9984
rect 3456 9952 3496 9984
rect 3528 9952 3568 9984
rect 3600 9952 3640 9984
rect 3672 9952 3712 9984
rect 3744 9952 3784 9984
rect 3816 9952 3856 9984
rect 3888 9952 3928 9984
rect 3960 9952 4000 9984
rect 0 9912 4000 9952
rect 0 9880 40 9912
rect 72 9880 112 9912
rect 144 9880 184 9912
rect 216 9880 256 9912
rect 288 9880 328 9912
rect 360 9880 400 9912
rect 432 9880 472 9912
rect 504 9880 544 9912
rect 576 9880 616 9912
rect 648 9880 688 9912
rect 720 9880 760 9912
rect 792 9880 832 9912
rect 864 9880 904 9912
rect 936 9880 976 9912
rect 1008 9880 1048 9912
rect 1080 9880 1120 9912
rect 1152 9880 1192 9912
rect 1224 9880 1264 9912
rect 1296 9880 1336 9912
rect 1368 9880 1408 9912
rect 1440 9880 1480 9912
rect 1512 9880 1552 9912
rect 1584 9880 1624 9912
rect 1656 9880 1696 9912
rect 1728 9880 1768 9912
rect 1800 9880 1840 9912
rect 1872 9880 1912 9912
rect 1944 9880 1984 9912
rect 2016 9880 2056 9912
rect 2088 9880 2128 9912
rect 2160 9880 2200 9912
rect 2232 9880 2272 9912
rect 2304 9880 2344 9912
rect 2376 9880 2416 9912
rect 2448 9880 2488 9912
rect 2520 9880 2560 9912
rect 2592 9880 2632 9912
rect 2664 9880 2704 9912
rect 2736 9880 2776 9912
rect 2808 9880 2848 9912
rect 2880 9880 2920 9912
rect 2952 9880 2992 9912
rect 3024 9880 3064 9912
rect 3096 9880 3136 9912
rect 3168 9880 3208 9912
rect 3240 9880 3280 9912
rect 3312 9880 3352 9912
rect 3384 9880 3424 9912
rect 3456 9880 3496 9912
rect 3528 9880 3568 9912
rect 3600 9880 3640 9912
rect 3672 9880 3712 9912
rect 3744 9880 3784 9912
rect 3816 9880 3856 9912
rect 3888 9880 3928 9912
rect 3960 9880 4000 9912
rect 0 9840 4000 9880
rect 0 9808 40 9840
rect 72 9808 112 9840
rect 144 9808 184 9840
rect 216 9808 256 9840
rect 288 9808 328 9840
rect 360 9808 400 9840
rect 432 9808 472 9840
rect 504 9808 544 9840
rect 576 9808 616 9840
rect 648 9808 688 9840
rect 720 9808 760 9840
rect 792 9808 832 9840
rect 864 9808 904 9840
rect 936 9808 976 9840
rect 1008 9808 1048 9840
rect 1080 9808 1120 9840
rect 1152 9808 1192 9840
rect 1224 9808 1264 9840
rect 1296 9808 1336 9840
rect 1368 9808 1408 9840
rect 1440 9808 1480 9840
rect 1512 9808 1552 9840
rect 1584 9808 1624 9840
rect 1656 9808 1696 9840
rect 1728 9808 1768 9840
rect 1800 9808 1840 9840
rect 1872 9808 1912 9840
rect 1944 9808 1984 9840
rect 2016 9808 2056 9840
rect 2088 9808 2128 9840
rect 2160 9808 2200 9840
rect 2232 9808 2272 9840
rect 2304 9808 2344 9840
rect 2376 9808 2416 9840
rect 2448 9808 2488 9840
rect 2520 9808 2560 9840
rect 2592 9808 2632 9840
rect 2664 9808 2704 9840
rect 2736 9808 2776 9840
rect 2808 9808 2848 9840
rect 2880 9808 2920 9840
rect 2952 9808 2992 9840
rect 3024 9808 3064 9840
rect 3096 9808 3136 9840
rect 3168 9808 3208 9840
rect 3240 9808 3280 9840
rect 3312 9808 3352 9840
rect 3384 9808 3424 9840
rect 3456 9808 3496 9840
rect 3528 9808 3568 9840
rect 3600 9808 3640 9840
rect 3672 9808 3712 9840
rect 3744 9808 3784 9840
rect 3816 9808 3856 9840
rect 3888 9808 3928 9840
rect 3960 9808 4000 9840
rect 0 9768 4000 9808
rect 0 9736 40 9768
rect 72 9736 112 9768
rect 144 9736 184 9768
rect 216 9736 256 9768
rect 288 9736 328 9768
rect 360 9736 400 9768
rect 432 9736 472 9768
rect 504 9736 544 9768
rect 576 9736 616 9768
rect 648 9736 688 9768
rect 720 9736 760 9768
rect 792 9736 832 9768
rect 864 9736 904 9768
rect 936 9736 976 9768
rect 1008 9736 1048 9768
rect 1080 9736 1120 9768
rect 1152 9736 1192 9768
rect 1224 9736 1264 9768
rect 1296 9736 1336 9768
rect 1368 9736 1408 9768
rect 1440 9736 1480 9768
rect 1512 9736 1552 9768
rect 1584 9736 1624 9768
rect 1656 9736 1696 9768
rect 1728 9736 1768 9768
rect 1800 9736 1840 9768
rect 1872 9736 1912 9768
rect 1944 9736 1984 9768
rect 2016 9736 2056 9768
rect 2088 9736 2128 9768
rect 2160 9736 2200 9768
rect 2232 9736 2272 9768
rect 2304 9736 2344 9768
rect 2376 9736 2416 9768
rect 2448 9736 2488 9768
rect 2520 9736 2560 9768
rect 2592 9736 2632 9768
rect 2664 9736 2704 9768
rect 2736 9736 2776 9768
rect 2808 9736 2848 9768
rect 2880 9736 2920 9768
rect 2952 9736 2992 9768
rect 3024 9736 3064 9768
rect 3096 9736 3136 9768
rect 3168 9736 3208 9768
rect 3240 9736 3280 9768
rect 3312 9736 3352 9768
rect 3384 9736 3424 9768
rect 3456 9736 3496 9768
rect 3528 9736 3568 9768
rect 3600 9736 3640 9768
rect 3672 9736 3712 9768
rect 3744 9736 3784 9768
rect 3816 9736 3856 9768
rect 3888 9736 3928 9768
rect 3960 9736 4000 9768
rect 0 9696 4000 9736
rect 0 9664 40 9696
rect 72 9664 112 9696
rect 144 9664 184 9696
rect 216 9664 256 9696
rect 288 9664 328 9696
rect 360 9664 400 9696
rect 432 9664 472 9696
rect 504 9664 544 9696
rect 576 9664 616 9696
rect 648 9664 688 9696
rect 720 9664 760 9696
rect 792 9664 832 9696
rect 864 9664 904 9696
rect 936 9664 976 9696
rect 1008 9664 1048 9696
rect 1080 9664 1120 9696
rect 1152 9664 1192 9696
rect 1224 9664 1264 9696
rect 1296 9664 1336 9696
rect 1368 9664 1408 9696
rect 1440 9664 1480 9696
rect 1512 9664 1552 9696
rect 1584 9664 1624 9696
rect 1656 9664 1696 9696
rect 1728 9664 1768 9696
rect 1800 9664 1840 9696
rect 1872 9664 1912 9696
rect 1944 9664 1984 9696
rect 2016 9664 2056 9696
rect 2088 9664 2128 9696
rect 2160 9664 2200 9696
rect 2232 9664 2272 9696
rect 2304 9664 2344 9696
rect 2376 9664 2416 9696
rect 2448 9664 2488 9696
rect 2520 9664 2560 9696
rect 2592 9664 2632 9696
rect 2664 9664 2704 9696
rect 2736 9664 2776 9696
rect 2808 9664 2848 9696
rect 2880 9664 2920 9696
rect 2952 9664 2992 9696
rect 3024 9664 3064 9696
rect 3096 9664 3136 9696
rect 3168 9664 3208 9696
rect 3240 9664 3280 9696
rect 3312 9664 3352 9696
rect 3384 9664 3424 9696
rect 3456 9664 3496 9696
rect 3528 9664 3568 9696
rect 3600 9664 3640 9696
rect 3672 9664 3712 9696
rect 3744 9664 3784 9696
rect 3816 9664 3856 9696
rect 3888 9664 3928 9696
rect 3960 9664 4000 9696
rect 0 9624 4000 9664
rect 0 9592 40 9624
rect 72 9592 112 9624
rect 144 9592 184 9624
rect 216 9592 256 9624
rect 288 9592 328 9624
rect 360 9592 400 9624
rect 432 9592 472 9624
rect 504 9592 544 9624
rect 576 9592 616 9624
rect 648 9592 688 9624
rect 720 9592 760 9624
rect 792 9592 832 9624
rect 864 9592 904 9624
rect 936 9592 976 9624
rect 1008 9592 1048 9624
rect 1080 9592 1120 9624
rect 1152 9592 1192 9624
rect 1224 9592 1264 9624
rect 1296 9592 1336 9624
rect 1368 9592 1408 9624
rect 1440 9592 1480 9624
rect 1512 9592 1552 9624
rect 1584 9592 1624 9624
rect 1656 9592 1696 9624
rect 1728 9592 1768 9624
rect 1800 9592 1840 9624
rect 1872 9592 1912 9624
rect 1944 9592 1984 9624
rect 2016 9592 2056 9624
rect 2088 9592 2128 9624
rect 2160 9592 2200 9624
rect 2232 9592 2272 9624
rect 2304 9592 2344 9624
rect 2376 9592 2416 9624
rect 2448 9592 2488 9624
rect 2520 9592 2560 9624
rect 2592 9592 2632 9624
rect 2664 9592 2704 9624
rect 2736 9592 2776 9624
rect 2808 9592 2848 9624
rect 2880 9592 2920 9624
rect 2952 9592 2992 9624
rect 3024 9592 3064 9624
rect 3096 9592 3136 9624
rect 3168 9592 3208 9624
rect 3240 9592 3280 9624
rect 3312 9592 3352 9624
rect 3384 9592 3424 9624
rect 3456 9592 3496 9624
rect 3528 9592 3568 9624
rect 3600 9592 3640 9624
rect 3672 9592 3712 9624
rect 3744 9592 3784 9624
rect 3816 9592 3856 9624
rect 3888 9592 3928 9624
rect 3960 9592 4000 9624
rect 0 9552 4000 9592
rect 0 9520 40 9552
rect 72 9520 112 9552
rect 144 9520 184 9552
rect 216 9520 256 9552
rect 288 9520 328 9552
rect 360 9520 400 9552
rect 432 9520 472 9552
rect 504 9520 544 9552
rect 576 9520 616 9552
rect 648 9520 688 9552
rect 720 9520 760 9552
rect 792 9520 832 9552
rect 864 9520 904 9552
rect 936 9520 976 9552
rect 1008 9520 1048 9552
rect 1080 9520 1120 9552
rect 1152 9520 1192 9552
rect 1224 9520 1264 9552
rect 1296 9520 1336 9552
rect 1368 9520 1408 9552
rect 1440 9520 1480 9552
rect 1512 9520 1552 9552
rect 1584 9520 1624 9552
rect 1656 9520 1696 9552
rect 1728 9520 1768 9552
rect 1800 9520 1840 9552
rect 1872 9520 1912 9552
rect 1944 9520 1984 9552
rect 2016 9520 2056 9552
rect 2088 9520 2128 9552
rect 2160 9520 2200 9552
rect 2232 9520 2272 9552
rect 2304 9520 2344 9552
rect 2376 9520 2416 9552
rect 2448 9520 2488 9552
rect 2520 9520 2560 9552
rect 2592 9520 2632 9552
rect 2664 9520 2704 9552
rect 2736 9520 2776 9552
rect 2808 9520 2848 9552
rect 2880 9520 2920 9552
rect 2952 9520 2992 9552
rect 3024 9520 3064 9552
rect 3096 9520 3136 9552
rect 3168 9520 3208 9552
rect 3240 9520 3280 9552
rect 3312 9520 3352 9552
rect 3384 9520 3424 9552
rect 3456 9520 3496 9552
rect 3528 9520 3568 9552
rect 3600 9520 3640 9552
rect 3672 9520 3712 9552
rect 3744 9520 3784 9552
rect 3816 9520 3856 9552
rect 3888 9520 3928 9552
rect 3960 9520 4000 9552
rect 0 9480 4000 9520
rect 0 9448 40 9480
rect 72 9448 112 9480
rect 144 9448 184 9480
rect 216 9448 256 9480
rect 288 9448 328 9480
rect 360 9448 400 9480
rect 432 9448 472 9480
rect 504 9448 544 9480
rect 576 9448 616 9480
rect 648 9448 688 9480
rect 720 9448 760 9480
rect 792 9448 832 9480
rect 864 9448 904 9480
rect 936 9448 976 9480
rect 1008 9448 1048 9480
rect 1080 9448 1120 9480
rect 1152 9448 1192 9480
rect 1224 9448 1264 9480
rect 1296 9448 1336 9480
rect 1368 9448 1408 9480
rect 1440 9448 1480 9480
rect 1512 9448 1552 9480
rect 1584 9448 1624 9480
rect 1656 9448 1696 9480
rect 1728 9448 1768 9480
rect 1800 9448 1840 9480
rect 1872 9448 1912 9480
rect 1944 9448 1984 9480
rect 2016 9448 2056 9480
rect 2088 9448 2128 9480
rect 2160 9448 2200 9480
rect 2232 9448 2272 9480
rect 2304 9448 2344 9480
rect 2376 9448 2416 9480
rect 2448 9448 2488 9480
rect 2520 9448 2560 9480
rect 2592 9448 2632 9480
rect 2664 9448 2704 9480
rect 2736 9448 2776 9480
rect 2808 9448 2848 9480
rect 2880 9448 2920 9480
rect 2952 9448 2992 9480
rect 3024 9448 3064 9480
rect 3096 9448 3136 9480
rect 3168 9448 3208 9480
rect 3240 9448 3280 9480
rect 3312 9448 3352 9480
rect 3384 9448 3424 9480
rect 3456 9448 3496 9480
rect 3528 9448 3568 9480
rect 3600 9448 3640 9480
rect 3672 9448 3712 9480
rect 3744 9448 3784 9480
rect 3816 9448 3856 9480
rect 3888 9448 3928 9480
rect 3960 9448 4000 9480
rect 0 9408 4000 9448
rect 0 9376 40 9408
rect 72 9376 112 9408
rect 144 9376 184 9408
rect 216 9376 256 9408
rect 288 9376 328 9408
rect 360 9376 400 9408
rect 432 9376 472 9408
rect 504 9376 544 9408
rect 576 9376 616 9408
rect 648 9376 688 9408
rect 720 9376 760 9408
rect 792 9376 832 9408
rect 864 9376 904 9408
rect 936 9376 976 9408
rect 1008 9376 1048 9408
rect 1080 9376 1120 9408
rect 1152 9376 1192 9408
rect 1224 9376 1264 9408
rect 1296 9376 1336 9408
rect 1368 9376 1408 9408
rect 1440 9376 1480 9408
rect 1512 9376 1552 9408
rect 1584 9376 1624 9408
rect 1656 9376 1696 9408
rect 1728 9376 1768 9408
rect 1800 9376 1840 9408
rect 1872 9376 1912 9408
rect 1944 9376 1984 9408
rect 2016 9376 2056 9408
rect 2088 9376 2128 9408
rect 2160 9376 2200 9408
rect 2232 9376 2272 9408
rect 2304 9376 2344 9408
rect 2376 9376 2416 9408
rect 2448 9376 2488 9408
rect 2520 9376 2560 9408
rect 2592 9376 2632 9408
rect 2664 9376 2704 9408
rect 2736 9376 2776 9408
rect 2808 9376 2848 9408
rect 2880 9376 2920 9408
rect 2952 9376 2992 9408
rect 3024 9376 3064 9408
rect 3096 9376 3136 9408
rect 3168 9376 3208 9408
rect 3240 9376 3280 9408
rect 3312 9376 3352 9408
rect 3384 9376 3424 9408
rect 3456 9376 3496 9408
rect 3528 9376 3568 9408
rect 3600 9376 3640 9408
rect 3672 9376 3712 9408
rect 3744 9376 3784 9408
rect 3816 9376 3856 9408
rect 3888 9376 3928 9408
rect 3960 9376 4000 9408
rect 0 9336 4000 9376
rect 0 9304 40 9336
rect 72 9304 112 9336
rect 144 9304 184 9336
rect 216 9304 256 9336
rect 288 9304 328 9336
rect 360 9304 400 9336
rect 432 9304 472 9336
rect 504 9304 544 9336
rect 576 9304 616 9336
rect 648 9304 688 9336
rect 720 9304 760 9336
rect 792 9304 832 9336
rect 864 9304 904 9336
rect 936 9304 976 9336
rect 1008 9304 1048 9336
rect 1080 9304 1120 9336
rect 1152 9304 1192 9336
rect 1224 9304 1264 9336
rect 1296 9304 1336 9336
rect 1368 9304 1408 9336
rect 1440 9304 1480 9336
rect 1512 9304 1552 9336
rect 1584 9304 1624 9336
rect 1656 9304 1696 9336
rect 1728 9304 1768 9336
rect 1800 9304 1840 9336
rect 1872 9304 1912 9336
rect 1944 9304 1984 9336
rect 2016 9304 2056 9336
rect 2088 9304 2128 9336
rect 2160 9304 2200 9336
rect 2232 9304 2272 9336
rect 2304 9304 2344 9336
rect 2376 9304 2416 9336
rect 2448 9304 2488 9336
rect 2520 9304 2560 9336
rect 2592 9304 2632 9336
rect 2664 9304 2704 9336
rect 2736 9304 2776 9336
rect 2808 9304 2848 9336
rect 2880 9304 2920 9336
rect 2952 9304 2992 9336
rect 3024 9304 3064 9336
rect 3096 9304 3136 9336
rect 3168 9304 3208 9336
rect 3240 9304 3280 9336
rect 3312 9304 3352 9336
rect 3384 9304 3424 9336
rect 3456 9304 3496 9336
rect 3528 9304 3568 9336
rect 3600 9304 3640 9336
rect 3672 9304 3712 9336
rect 3744 9304 3784 9336
rect 3816 9304 3856 9336
rect 3888 9304 3928 9336
rect 3960 9304 4000 9336
rect 0 9264 4000 9304
rect 0 9232 40 9264
rect 72 9232 112 9264
rect 144 9232 184 9264
rect 216 9232 256 9264
rect 288 9232 328 9264
rect 360 9232 400 9264
rect 432 9232 472 9264
rect 504 9232 544 9264
rect 576 9232 616 9264
rect 648 9232 688 9264
rect 720 9232 760 9264
rect 792 9232 832 9264
rect 864 9232 904 9264
rect 936 9232 976 9264
rect 1008 9232 1048 9264
rect 1080 9232 1120 9264
rect 1152 9232 1192 9264
rect 1224 9232 1264 9264
rect 1296 9232 1336 9264
rect 1368 9232 1408 9264
rect 1440 9232 1480 9264
rect 1512 9232 1552 9264
rect 1584 9232 1624 9264
rect 1656 9232 1696 9264
rect 1728 9232 1768 9264
rect 1800 9232 1840 9264
rect 1872 9232 1912 9264
rect 1944 9232 1984 9264
rect 2016 9232 2056 9264
rect 2088 9232 2128 9264
rect 2160 9232 2200 9264
rect 2232 9232 2272 9264
rect 2304 9232 2344 9264
rect 2376 9232 2416 9264
rect 2448 9232 2488 9264
rect 2520 9232 2560 9264
rect 2592 9232 2632 9264
rect 2664 9232 2704 9264
rect 2736 9232 2776 9264
rect 2808 9232 2848 9264
rect 2880 9232 2920 9264
rect 2952 9232 2992 9264
rect 3024 9232 3064 9264
rect 3096 9232 3136 9264
rect 3168 9232 3208 9264
rect 3240 9232 3280 9264
rect 3312 9232 3352 9264
rect 3384 9232 3424 9264
rect 3456 9232 3496 9264
rect 3528 9232 3568 9264
rect 3600 9232 3640 9264
rect 3672 9232 3712 9264
rect 3744 9232 3784 9264
rect 3816 9232 3856 9264
rect 3888 9232 3928 9264
rect 3960 9232 4000 9264
rect 0 9192 4000 9232
rect 0 9160 40 9192
rect 72 9160 112 9192
rect 144 9160 184 9192
rect 216 9160 256 9192
rect 288 9160 328 9192
rect 360 9160 400 9192
rect 432 9160 472 9192
rect 504 9160 544 9192
rect 576 9160 616 9192
rect 648 9160 688 9192
rect 720 9160 760 9192
rect 792 9160 832 9192
rect 864 9160 904 9192
rect 936 9160 976 9192
rect 1008 9160 1048 9192
rect 1080 9160 1120 9192
rect 1152 9160 1192 9192
rect 1224 9160 1264 9192
rect 1296 9160 1336 9192
rect 1368 9160 1408 9192
rect 1440 9160 1480 9192
rect 1512 9160 1552 9192
rect 1584 9160 1624 9192
rect 1656 9160 1696 9192
rect 1728 9160 1768 9192
rect 1800 9160 1840 9192
rect 1872 9160 1912 9192
rect 1944 9160 1984 9192
rect 2016 9160 2056 9192
rect 2088 9160 2128 9192
rect 2160 9160 2200 9192
rect 2232 9160 2272 9192
rect 2304 9160 2344 9192
rect 2376 9160 2416 9192
rect 2448 9160 2488 9192
rect 2520 9160 2560 9192
rect 2592 9160 2632 9192
rect 2664 9160 2704 9192
rect 2736 9160 2776 9192
rect 2808 9160 2848 9192
rect 2880 9160 2920 9192
rect 2952 9160 2992 9192
rect 3024 9160 3064 9192
rect 3096 9160 3136 9192
rect 3168 9160 3208 9192
rect 3240 9160 3280 9192
rect 3312 9160 3352 9192
rect 3384 9160 3424 9192
rect 3456 9160 3496 9192
rect 3528 9160 3568 9192
rect 3600 9160 3640 9192
rect 3672 9160 3712 9192
rect 3744 9160 3784 9192
rect 3816 9160 3856 9192
rect 3888 9160 3928 9192
rect 3960 9160 4000 9192
rect 0 9120 4000 9160
rect 0 9088 40 9120
rect 72 9088 112 9120
rect 144 9088 184 9120
rect 216 9088 256 9120
rect 288 9088 328 9120
rect 360 9088 400 9120
rect 432 9088 472 9120
rect 504 9088 544 9120
rect 576 9088 616 9120
rect 648 9088 688 9120
rect 720 9088 760 9120
rect 792 9088 832 9120
rect 864 9088 904 9120
rect 936 9088 976 9120
rect 1008 9088 1048 9120
rect 1080 9088 1120 9120
rect 1152 9088 1192 9120
rect 1224 9088 1264 9120
rect 1296 9088 1336 9120
rect 1368 9088 1408 9120
rect 1440 9088 1480 9120
rect 1512 9088 1552 9120
rect 1584 9088 1624 9120
rect 1656 9088 1696 9120
rect 1728 9088 1768 9120
rect 1800 9088 1840 9120
rect 1872 9088 1912 9120
rect 1944 9088 1984 9120
rect 2016 9088 2056 9120
rect 2088 9088 2128 9120
rect 2160 9088 2200 9120
rect 2232 9088 2272 9120
rect 2304 9088 2344 9120
rect 2376 9088 2416 9120
rect 2448 9088 2488 9120
rect 2520 9088 2560 9120
rect 2592 9088 2632 9120
rect 2664 9088 2704 9120
rect 2736 9088 2776 9120
rect 2808 9088 2848 9120
rect 2880 9088 2920 9120
rect 2952 9088 2992 9120
rect 3024 9088 3064 9120
rect 3096 9088 3136 9120
rect 3168 9088 3208 9120
rect 3240 9088 3280 9120
rect 3312 9088 3352 9120
rect 3384 9088 3424 9120
rect 3456 9088 3496 9120
rect 3528 9088 3568 9120
rect 3600 9088 3640 9120
rect 3672 9088 3712 9120
rect 3744 9088 3784 9120
rect 3816 9088 3856 9120
rect 3888 9088 3928 9120
rect 3960 9088 4000 9120
rect 0 9048 4000 9088
rect 0 9016 40 9048
rect 72 9016 112 9048
rect 144 9016 184 9048
rect 216 9016 256 9048
rect 288 9016 328 9048
rect 360 9016 400 9048
rect 432 9016 472 9048
rect 504 9016 544 9048
rect 576 9016 616 9048
rect 648 9016 688 9048
rect 720 9016 760 9048
rect 792 9016 832 9048
rect 864 9016 904 9048
rect 936 9016 976 9048
rect 1008 9016 1048 9048
rect 1080 9016 1120 9048
rect 1152 9016 1192 9048
rect 1224 9016 1264 9048
rect 1296 9016 1336 9048
rect 1368 9016 1408 9048
rect 1440 9016 1480 9048
rect 1512 9016 1552 9048
rect 1584 9016 1624 9048
rect 1656 9016 1696 9048
rect 1728 9016 1768 9048
rect 1800 9016 1840 9048
rect 1872 9016 1912 9048
rect 1944 9016 1984 9048
rect 2016 9016 2056 9048
rect 2088 9016 2128 9048
rect 2160 9016 2200 9048
rect 2232 9016 2272 9048
rect 2304 9016 2344 9048
rect 2376 9016 2416 9048
rect 2448 9016 2488 9048
rect 2520 9016 2560 9048
rect 2592 9016 2632 9048
rect 2664 9016 2704 9048
rect 2736 9016 2776 9048
rect 2808 9016 2848 9048
rect 2880 9016 2920 9048
rect 2952 9016 2992 9048
rect 3024 9016 3064 9048
rect 3096 9016 3136 9048
rect 3168 9016 3208 9048
rect 3240 9016 3280 9048
rect 3312 9016 3352 9048
rect 3384 9016 3424 9048
rect 3456 9016 3496 9048
rect 3528 9016 3568 9048
rect 3600 9016 3640 9048
rect 3672 9016 3712 9048
rect 3744 9016 3784 9048
rect 3816 9016 3856 9048
rect 3888 9016 3928 9048
rect 3960 9016 4000 9048
rect 0 8976 4000 9016
rect 0 8944 40 8976
rect 72 8944 112 8976
rect 144 8944 184 8976
rect 216 8944 256 8976
rect 288 8944 328 8976
rect 360 8944 400 8976
rect 432 8944 472 8976
rect 504 8944 544 8976
rect 576 8944 616 8976
rect 648 8944 688 8976
rect 720 8944 760 8976
rect 792 8944 832 8976
rect 864 8944 904 8976
rect 936 8944 976 8976
rect 1008 8944 1048 8976
rect 1080 8944 1120 8976
rect 1152 8944 1192 8976
rect 1224 8944 1264 8976
rect 1296 8944 1336 8976
rect 1368 8944 1408 8976
rect 1440 8944 1480 8976
rect 1512 8944 1552 8976
rect 1584 8944 1624 8976
rect 1656 8944 1696 8976
rect 1728 8944 1768 8976
rect 1800 8944 1840 8976
rect 1872 8944 1912 8976
rect 1944 8944 1984 8976
rect 2016 8944 2056 8976
rect 2088 8944 2128 8976
rect 2160 8944 2200 8976
rect 2232 8944 2272 8976
rect 2304 8944 2344 8976
rect 2376 8944 2416 8976
rect 2448 8944 2488 8976
rect 2520 8944 2560 8976
rect 2592 8944 2632 8976
rect 2664 8944 2704 8976
rect 2736 8944 2776 8976
rect 2808 8944 2848 8976
rect 2880 8944 2920 8976
rect 2952 8944 2992 8976
rect 3024 8944 3064 8976
rect 3096 8944 3136 8976
rect 3168 8944 3208 8976
rect 3240 8944 3280 8976
rect 3312 8944 3352 8976
rect 3384 8944 3424 8976
rect 3456 8944 3496 8976
rect 3528 8944 3568 8976
rect 3600 8944 3640 8976
rect 3672 8944 3712 8976
rect 3744 8944 3784 8976
rect 3816 8944 3856 8976
rect 3888 8944 3928 8976
rect 3960 8944 4000 8976
rect 0 8904 4000 8944
rect 0 8872 40 8904
rect 72 8872 112 8904
rect 144 8872 184 8904
rect 216 8872 256 8904
rect 288 8872 328 8904
rect 360 8872 400 8904
rect 432 8872 472 8904
rect 504 8872 544 8904
rect 576 8872 616 8904
rect 648 8872 688 8904
rect 720 8872 760 8904
rect 792 8872 832 8904
rect 864 8872 904 8904
rect 936 8872 976 8904
rect 1008 8872 1048 8904
rect 1080 8872 1120 8904
rect 1152 8872 1192 8904
rect 1224 8872 1264 8904
rect 1296 8872 1336 8904
rect 1368 8872 1408 8904
rect 1440 8872 1480 8904
rect 1512 8872 1552 8904
rect 1584 8872 1624 8904
rect 1656 8872 1696 8904
rect 1728 8872 1768 8904
rect 1800 8872 1840 8904
rect 1872 8872 1912 8904
rect 1944 8872 1984 8904
rect 2016 8872 2056 8904
rect 2088 8872 2128 8904
rect 2160 8872 2200 8904
rect 2232 8872 2272 8904
rect 2304 8872 2344 8904
rect 2376 8872 2416 8904
rect 2448 8872 2488 8904
rect 2520 8872 2560 8904
rect 2592 8872 2632 8904
rect 2664 8872 2704 8904
rect 2736 8872 2776 8904
rect 2808 8872 2848 8904
rect 2880 8872 2920 8904
rect 2952 8872 2992 8904
rect 3024 8872 3064 8904
rect 3096 8872 3136 8904
rect 3168 8872 3208 8904
rect 3240 8872 3280 8904
rect 3312 8872 3352 8904
rect 3384 8872 3424 8904
rect 3456 8872 3496 8904
rect 3528 8872 3568 8904
rect 3600 8872 3640 8904
rect 3672 8872 3712 8904
rect 3744 8872 3784 8904
rect 3816 8872 3856 8904
rect 3888 8872 3928 8904
rect 3960 8872 4000 8904
rect 0 8832 4000 8872
rect 0 8800 40 8832
rect 72 8800 112 8832
rect 144 8800 184 8832
rect 216 8800 256 8832
rect 288 8800 328 8832
rect 360 8800 400 8832
rect 432 8800 472 8832
rect 504 8800 544 8832
rect 576 8800 616 8832
rect 648 8800 688 8832
rect 720 8800 760 8832
rect 792 8800 832 8832
rect 864 8800 904 8832
rect 936 8800 976 8832
rect 1008 8800 1048 8832
rect 1080 8800 1120 8832
rect 1152 8800 1192 8832
rect 1224 8800 1264 8832
rect 1296 8800 1336 8832
rect 1368 8800 1408 8832
rect 1440 8800 1480 8832
rect 1512 8800 1552 8832
rect 1584 8800 1624 8832
rect 1656 8800 1696 8832
rect 1728 8800 1768 8832
rect 1800 8800 1840 8832
rect 1872 8800 1912 8832
rect 1944 8800 1984 8832
rect 2016 8800 2056 8832
rect 2088 8800 2128 8832
rect 2160 8800 2200 8832
rect 2232 8800 2272 8832
rect 2304 8800 2344 8832
rect 2376 8800 2416 8832
rect 2448 8800 2488 8832
rect 2520 8800 2560 8832
rect 2592 8800 2632 8832
rect 2664 8800 2704 8832
rect 2736 8800 2776 8832
rect 2808 8800 2848 8832
rect 2880 8800 2920 8832
rect 2952 8800 2992 8832
rect 3024 8800 3064 8832
rect 3096 8800 3136 8832
rect 3168 8800 3208 8832
rect 3240 8800 3280 8832
rect 3312 8800 3352 8832
rect 3384 8800 3424 8832
rect 3456 8800 3496 8832
rect 3528 8800 3568 8832
rect 3600 8800 3640 8832
rect 3672 8800 3712 8832
rect 3744 8800 3784 8832
rect 3816 8800 3856 8832
rect 3888 8800 3928 8832
rect 3960 8800 4000 8832
rect 0 8760 4000 8800
rect 0 8728 40 8760
rect 72 8728 112 8760
rect 144 8728 184 8760
rect 216 8728 256 8760
rect 288 8728 328 8760
rect 360 8728 400 8760
rect 432 8728 472 8760
rect 504 8728 544 8760
rect 576 8728 616 8760
rect 648 8728 688 8760
rect 720 8728 760 8760
rect 792 8728 832 8760
rect 864 8728 904 8760
rect 936 8728 976 8760
rect 1008 8728 1048 8760
rect 1080 8728 1120 8760
rect 1152 8728 1192 8760
rect 1224 8728 1264 8760
rect 1296 8728 1336 8760
rect 1368 8728 1408 8760
rect 1440 8728 1480 8760
rect 1512 8728 1552 8760
rect 1584 8728 1624 8760
rect 1656 8728 1696 8760
rect 1728 8728 1768 8760
rect 1800 8728 1840 8760
rect 1872 8728 1912 8760
rect 1944 8728 1984 8760
rect 2016 8728 2056 8760
rect 2088 8728 2128 8760
rect 2160 8728 2200 8760
rect 2232 8728 2272 8760
rect 2304 8728 2344 8760
rect 2376 8728 2416 8760
rect 2448 8728 2488 8760
rect 2520 8728 2560 8760
rect 2592 8728 2632 8760
rect 2664 8728 2704 8760
rect 2736 8728 2776 8760
rect 2808 8728 2848 8760
rect 2880 8728 2920 8760
rect 2952 8728 2992 8760
rect 3024 8728 3064 8760
rect 3096 8728 3136 8760
rect 3168 8728 3208 8760
rect 3240 8728 3280 8760
rect 3312 8728 3352 8760
rect 3384 8728 3424 8760
rect 3456 8728 3496 8760
rect 3528 8728 3568 8760
rect 3600 8728 3640 8760
rect 3672 8728 3712 8760
rect 3744 8728 3784 8760
rect 3816 8728 3856 8760
rect 3888 8728 3928 8760
rect 3960 8728 4000 8760
rect 0 8688 4000 8728
rect 0 8656 40 8688
rect 72 8656 112 8688
rect 144 8656 184 8688
rect 216 8656 256 8688
rect 288 8656 328 8688
rect 360 8656 400 8688
rect 432 8656 472 8688
rect 504 8656 544 8688
rect 576 8656 616 8688
rect 648 8656 688 8688
rect 720 8656 760 8688
rect 792 8656 832 8688
rect 864 8656 904 8688
rect 936 8656 976 8688
rect 1008 8656 1048 8688
rect 1080 8656 1120 8688
rect 1152 8656 1192 8688
rect 1224 8656 1264 8688
rect 1296 8656 1336 8688
rect 1368 8656 1408 8688
rect 1440 8656 1480 8688
rect 1512 8656 1552 8688
rect 1584 8656 1624 8688
rect 1656 8656 1696 8688
rect 1728 8656 1768 8688
rect 1800 8656 1840 8688
rect 1872 8656 1912 8688
rect 1944 8656 1984 8688
rect 2016 8656 2056 8688
rect 2088 8656 2128 8688
rect 2160 8656 2200 8688
rect 2232 8656 2272 8688
rect 2304 8656 2344 8688
rect 2376 8656 2416 8688
rect 2448 8656 2488 8688
rect 2520 8656 2560 8688
rect 2592 8656 2632 8688
rect 2664 8656 2704 8688
rect 2736 8656 2776 8688
rect 2808 8656 2848 8688
rect 2880 8656 2920 8688
rect 2952 8656 2992 8688
rect 3024 8656 3064 8688
rect 3096 8656 3136 8688
rect 3168 8656 3208 8688
rect 3240 8656 3280 8688
rect 3312 8656 3352 8688
rect 3384 8656 3424 8688
rect 3456 8656 3496 8688
rect 3528 8656 3568 8688
rect 3600 8656 3640 8688
rect 3672 8656 3712 8688
rect 3744 8656 3784 8688
rect 3816 8656 3856 8688
rect 3888 8656 3928 8688
rect 3960 8656 4000 8688
rect 0 8616 4000 8656
rect 0 8584 40 8616
rect 72 8584 112 8616
rect 144 8584 184 8616
rect 216 8584 256 8616
rect 288 8584 328 8616
rect 360 8584 400 8616
rect 432 8584 472 8616
rect 504 8584 544 8616
rect 576 8584 616 8616
rect 648 8584 688 8616
rect 720 8584 760 8616
rect 792 8584 832 8616
rect 864 8584 904 8616
rect 936 8584 976 8616
rect 1008 8584 1048 8616
rect 1080 8584 1120 8616
rect 1152 8584 1192 8616
rect 1224 8584 1264 8616
rect 1296 8584 1336 8616
rect 1368 8584 1408 8616
rect 1440 8584 1480 8616
rect 1512 8584 1552 8616
rect 1584 8584 1624 8616
rect 1656 8584 1696 8616
rect 1728 8584 1768 8616
rect 1800 8584 1840 8616
rect 1872 8584 1912 8616
rect 1944 8584 1984 8616
rect 2016 8584 2056 8616
rect 2088 8584 2128 8616
rect 2160 8584 2200 8616
rect 2232 8584 2272 8616
rect 2304 8584 2344 8616
rect 2376 8584 2416 8616
rect 2448 8584 2488 8616
rect 2520 8584 2560 8616
rect 2592 8584 2632 8616
rect 2664 8584 2704 8616
rect 2736 8584 2776 8616
rect 2808 8584 2848 8616
rect 2880 8584 2920 8616
rect 2952 8584 2992 8616
rect 3024 8584 3064 8616
rect 3096 8584 3136 8616
rect 3168 8584 3208 8616
rect 3240 8584 3280 8616
rect 3312 8584 3352 8616
rect 3384 8584 3424 8616
rect 3456 8584 3496 8616
rect 3528 8584 3568 8616
rect 3600 8584 3640 8616
rect 3672 8584 3712 8616
rect 3744 8584 3784 8616
rect 3816 8584 3856 8616
rect 3888 8584 3928 8616
rect 3960 8584 4000 8616
rect 0 8544 4000 8584
rect 0 8512 40 8544
rect 72 8512 112 8544
rect 144 8512 184 8544
rect 216 8512 256 8544
rect 288 8512 328 8544
rect 360 8512 400 8544
rect 432 8512 472 8544
rect 504 8512 544 8544
rect 576 8512 616 8544
rect 648 8512 688 8544
rect 720 8512 760 8544
rect 792 8512 832 8544
rect 864 8512 904 8544
rect 936 8512 976 8544
rect 1008 8512 1048 8544
rect 1080 8512 1120 8544
rect 1152 8512 1192 8544
rect 1224 8512 1264 8544
rect 1296 8512 1336 8544
rect 1368 8512 1408 8544
rect 1440 8512 1480 8544
rect 1512 8512 1552 8544
rect 1584 8512 1624 8544
rect 1656 8512 1696 8544
rect 1728 8512 1768 8544
rect 1800 8512 1840 8544
rect 1872 8512 1912 8544
rect 1944 8512 1984 8544
rect 2016 8512 2056 8544
rect 2088 8512 2128 8544
rect 2160 8512 2200 8544
rect 2232 8512 2272 8544
rect 2304 8512 2344 8544
rect 2376 8512 2416 8544
rect 2448 8512 2488 8544
rect 2520 8512 2560 8544
rect 2592 8512 2632 8544
rect 2664 8512 2704 8544
rect 2736 8512 2776 8544
rect 2808 8512 2848 8544
rect 2880 8512 2920 8544
rect 2952 8512 2992 8544
rect 3024 8512 3064 8544
rect 3096 8512 3136 8544
rect 3168 8512 3208 8544
rect 3240 8512 3280 8544
rect 3312 8512 3352 8544
rect 3384 8512 3424 8544
rect 3456 8512 3496 8544
rect 3528 8512 3568 8544
rect 3600 8512 3640 8544
rect 3672 8512 3712 8544
rect 3744 8512 3784 8544
rect 3816 8512 3856 8544
rect 3888 8512 3928 8544
rect 3960 8512 4000 8544
rect 0 8472 4000 8512
rect 0 8440 40 8472
rect 72 8440 112 8472
rect 144 8440 184 8472
rect 216 8440 256 8472
rect 288 8440 328 8472
rect 360 8440 400 8472
rect 432 8440 472 8472
rect 504 8440 544 8472
rect 576 8440 616 8472
rect 648 8440 688 8472
rect 720 8440 760 8472
rect 792 8440 832 8472
rect 864 8440 904 8472
rect 936 8440 976 8472
rect 1008 8440 1048 8472
rect 1080 8440 1120 8472
rect 1152 8440 1192 8472
rect 1224 8440 1264 8472
rect 1296 8440 1336 8472
rect 1368 8440 1408 8472
rect 1440 8440 1480 8472
rect 1512 8440 1552 8472
rect 1584 8440 1624 8472
rect 1656 8440 1696 8472
rect 1728 8440 1768 8472
rect 1800 8440 1840 8472
rect 1872 8440 1912 8472
rect 1944 8440 1984 8472
rect 2016 8440 2056 8472
rect 2088 8440 2128 8472
rect 2160 8440 2200 8472
rect 2232 8440 2272 8472
rect 2304 8440 2344 8472
rect 2376 8440 2416 8472
rect 2448 8440 2488 8472
rect 2520 8440 2560 8472
rect 2592 8440 2632 8472
rect 2664 8440 2704 8472
rect 2736 8440 2776 8472
rect 2808 8440 2848 8472
rect 2880 8440 2920 8472
rect 2952 8440 2992 8472
rect 3024 8440 3064 8472
rect 3096 8440 3136 8472
rect 3168 8440 3208 8472
rect 3240 8440 3280 8472
rect 3312 8440 3352 8472
rect 3384 8440 3424 8472
rect 3456 8440 3496 8472
rect 3528 8440 3568 8472
rect 3600 8440 3640 8472
rect 3672 8440 3712 8472
rect 3744 8440 3784 8472
rect 3816 8440 3856 8472
rect 3888 8440 3928 8472
rect 3960 8440 4000 8472
rect 0 8400 4000 8440
rect 0 8368 40 8400
rect 72 8368 112 8400
rect 144 8368 184 8400
rect 216 8368 256 8400
rect 288 8368 328 8400
rect 360 8368 400 8400
rect 432 8368 472 8400
rect 504 8368 544 8400
rect 576 8368 616 8400
rect 648 8368 688 8400
rect 720 8368 760 8400
rect 792 8368 832 8400
rect 864 8368 904 8400
rect 936 8368 976 8400
rect 1008 8368 1048 8400
rect 1080 8368 1120 8400
rect 1152 8368 1192 8400
rect 1224 8368 1264 8400
rect 1296 8368 1336 8400
rect 1368 8368 1408 8400
rect 1440 8368 1480 8400
rect 1512 8368 1552 8400
rect 1584 8368 1624 8400
rect 1656 8368 1696 8400
rect 1728 8368 1768 8400
rect 1800 8368 1840 8400
rect 1872 8368 1912 8400
rect 1944 8368 1984 8400
rect 2016 8368 2056 8400
rect 2088 8368 2128 8400
rect 2160 8368 2200 8400
rect 2232 8368 2272 8400
rect 2304 8368 2344 8400
rect 2376 8368 2416 8400
rect 2448 8368 2488 8400
rect 2520 8368 2560 8400
rect 2592 8368 2632 8400
rect 2664 8368 2704 8400
rect 2736 8368 2776 8400
rect 2808 8368 2848 8400
rect 2880 8368 2920 8400
rect 2952 8368 2992 8400
rect 3024 8368 3064 8400
rect 3096 8368 3136 8400
rect 3168 8368 3208 8400
rect 3240 8368 3280 8400
rect 3312 8368 3352 8400
rect 3384 8368 3424 8400
rect 3456 8368 3496 8400
rect 3528 8368 3568 8400
rect 3600 8368 3640 8400
rect 3672 8368 3712 8400
rect 3744 8368 3784 8400
rect 3816 8368 3856 8400
rect 3888 8368 3928 8400
rect 3960 8368 4000 8400
rect 0 8328 4000 8368
rect 0 8296 40 8328
rect 72 8296 112 8328
rect 144 8296 184 8328
rect 216 8296 256 8328
rect 288 8296 328 8328
rect 360 8296 400 8328
rect 432 8296 472 8328
rect 504 8296 544 8328
rect 576 8296 616 8328
rect 648 8296 688 8328
rect 720 8296 760 8328
rect 792 8296 832 8328
rect 864 8296 904 8328
rect 936 8296 976 8328
rect 1008 8296 1048 8328
rect 1080 8296 1120 8328
rect 1152 8296 1192 8328
rect 1224 8296 1264 8328
rect 1296 8296 1336 8328
rect 1368 8296 1408 8328
rect 1440 8296 1480 8328
rect 1512 8296 1552 8328
rect 1584 8296 1624 8328
rect 1656 8296 1696 8328
rect 1728 8296 1768 8328
rect 1800 8296 1840 8328
rect 1872 8296 1912 8328
rect 1944 8296 1984 8328
rect 2016 8296 2056 8328
rect 2088 8296 2128 8328
rect 2160 8296 2200 8328
rect 2232 8296 2272 8328
rect 2304 8296 2344 8328
rect 2376 8296 2416 8328
rect 2448 8296 2488 8328
rect 2520 8296 2560 8328
rect 2592 8296 2632 8328
rect 2664 8296 2704 8328
rect 2736 8296 2776 8328
rect 2808 8296 2848 8328
rect 2880 8296 2920 8328
rect 2952 8296 2992 8328
rect 3024 8296 3064 8328
rect 3096 8296 3136 8328
rect 3168 8296 3208 8328
rect 3240 8296 3280 8328
rect 3312 8296 3352 8328
rect 3384 8296 3424 8328
rect 3456 8296 3496 8328
rect 3528 8296 3568 8328
rect 3600 8296 3640 8328
rect 3672 8296 3712 8328
rect 3744 8296 3784 8328
rect 3816 8296 3856 8328
rect 3888 8296 3928 8328
rect 3960 8296 4000 8328
rect 0 8256 4000 8296
rect 0 8224 40 8256
rect 72 8224 112 8256
rect 144 8224 184 8256
rect 216 8224 256 8256
rect 288 8224 328 8256
rect 360 8224 400 8256
rect 432 8224 472 8256
rect 504 8224 544 8256
rect 576 8224 616 8256
rect 648 8224 688 8256
rect 720 8224 760 8256
rect 792 8224 832 8256
rect 864 8224 904 8256
rect 936 8224 976 8256
rect 1008 8224 1048 8256
rect 1080 8224 1120 8256
rect 1152 8224 1192 8256
rect 1224 8224 1264 8256
rect 1296 8224 1336 8256
rect 1368 8224 1408 8256
rect 1440 8224 1480 8256
rect 1512 8224 1552 8256
rect 1584 8224 1624 8256
rect 1656 8224 1696 8256
rect 1728 8224 1768 8256
rect 1800 8224 1840 8256
rect 1872 8224 1912 8256
rect 1944 8224 1984 8256
rect 2016 8224 2056 8256
rect 2088 8224 2128 8256
rect 2160 8224 2200 8256
rect 2232 8224 2272 8256
rect 2304 8224 2344 8256
rect 2376 8224 2416 8256
rect 2448 8224 2488 8256
rect 2520 8224 2560 8256
rect 2592 8224 2632 8256
rect 2664 8224 2704 8256
rect 2736 8224 2776 8256
rect 2808 8224 2848 8256
rect 2880 8224 2920 8256
rect 2952 8224 2992 8256
rect 3024 8224 3064 8256
rect 3096 8224 3136 8256
rect 3168 8224 3208 8256
rect 3240 8224 3280 8256
rect 3312 8224 3352 8256
rect 3384 8224 3424 8256
rect 3456 8224 3496 8256
rect 3528 8224 3568 8256
rect 3600 8224 3640 8256
rect 3672 8224 3712 8256
rect 3744 8224 3784 8256
rect 3816 8224 3856 8256
rect 3888 8224 3928 8256
rect 3960 8224 4000 8256
rect 0 8184 4000 8224
rect 0 8152 40 8184
rect 72 8152 112 8184
rect 144 8152 184 8184
rect 216 8152 256 8184
rect 288 8152 328 8184
rect 360 8152 400 8184
rect 432 8152 472 8184
rect 504 8152 544 8184
rect 576 8152 616 8184
rect 648 8152 688 8184
rect 720 8152 760 8184
rect 792 8152 832 8184
rect 864 8152 904 8184
rect 936 8152 976 8184
rect 1008 8152 1048 8184
rect 1080 8152 1120 8184
rect 1152 8152 1192 8184
rect 1224 8152 1264 8184
rect 1296 8152 1336 8184
rect 1368 8152 1408 8184
rect 1440 8152 1480 8184
rect 1512 8152 1552 8184
rect 1584 8152 1624 8184
rect 1656 8152 1696 8184
rect 1728 8152 1768 8184
rect 1800 8152 1840 8184
rect 1872 8152 1912 8184
rect 1944 8152 1984 8184
rect 2016 8152 2056 8184
rect 2088 8152 2128 8184
rect 2160 8152 2200 8184
rect 2232 8152 2272 8184
rect 2304 8152 2344 8184
rect 2376 8152 2416 8184
rect 2448 8152 2488 8184
rect 2520 8152 2560 8184
rect 2592 8152 2632 8184
rect 2664 8152 2704 8184
rect 2736 8152 2776 8184
rect 2808 8152 2848 8184
rect 2880 8152 2920 8184
rect 2952 8152 2992 8184
rect 3024 8152 3064 8184
rect 3096 8152 3136 8184
rect 3168 8152 3208 8184
rect 3240 8152 3280 8184
rect 3312 8152 3352 8184
rect 3384 8152 3424 8184
rect 3456 8152 3496 8184
rect 3528 8152 3568 8184
rect 3600 8152 3640 8184
rect 3672 8152 3712 8184
rect 3744 8152 3784 8184
rect 3816 8152 3856 8184
rect 3888 8152 3928 8184
rect 3960 8152 4000 8184
rect 0 8112 4000 8152
rect 0 8080 40 8112
rect 72 8080 112 8112
rect 144 8080 184 8112
rect 216 8080 256 8112
rect 288 8080 328 8112
rect 360 8080 400 8112
rect 432 8080 472 8112
rect 504 8080 544 8112
rect 576 8080 616 8112
rect 648 8080 688 8112
rect 720 8080 760 8112
rect 792 8080 832 8112
rect 864 8080 904 8112
rect 936 8080 976 8112
rect 1008 8080 1048 8112
rect 1080 8080 1120 8112
rect 1152 8080 1192 8112
rect 1224 8080 1264 8112
rect 1296 8080 1336 8112
rect 1368 8080 1408 8112
rect 1440 8080 1480 8112
rect 1512 8080 1552 8112
rect 1584 8080 1624 8112
rect 1656 8080 1696 8112
rect 1728 8080 1768 8112
rect 1800 8080 1840 8112
rect 1872 8080 1912 8112
rect 1944 8080 1984 8112
rect 2016 8080 2056 8112
rect 2088 8080 2128 8112
rect 2160 8080 2200 8112
rect 2232 8080 2272 8112
rect 2304 8080 2344 8112
rect 2376 8080 2416 8112
rect 2448 8080 2488 8112
rect 2520 8080 2560 8112
rect 2592 8080 2632 8112
rect 2664 8080 2704 8112
rect 2736 8080 2776 8112
rect 2808 8080 2848 8112
rect 2880 8080 2920 8112
rect 2952 8080 2992 8112
rect 3024 8080 3064 8112
rect 3096 8080 3136 8112
rect 3168 8080 3208 8112
rect 3240 8080 3280 8112
rect 3312 8080 3352 8112
rect 3384 8080 3424 8112
rect 3456 8080 3496 8112
rect 3528 8080 3568 8112
rect 3600 8080 3640 8112
rect 3672 8080 3712 8112
rect 3744 8080 3784 8112
rect 3816 8080 3856 8112
rect 3888 8080 3928 8112
rect 3960 8080 4000 8112
rect 0 8040 4000 8080
rect 0 8008 40 8040
rect 72 8008 112 8040
rect 144 8008 184 8040
rect 216 8008 256 8040
rect 288 8008 328 8040
rect 360 8008 400 8040
rect 432 8008 472 8040
rect 504 8008 544 8040
rect 576 8008 616 8040
rect 648 8008 688 8040
rect 720 8008 760 8040
rect 792 8008 832 8040
rect 864 8008 904 8040
rect 936 8008 976 8040
rect 1008 8008 1048 8040
rect 1080 8008 1120 8040
rect 1152 8008 1192 8040
rect 1224 8008 1264 8040
rect 1296 8008 1336 8040
rect 1368 8008 1408 8040
rect 1440 8008 1480 8040
rect 1512 8008 1552 8040
rect 1584 8008 1624 8040
rect 1656 8008 1696 8040
rect 1728 8008 1768 8040
rect 1800 8008 1840 8040
rect 1872 8008 1912 8040
rect 1944 8008 1984 8040
rect 2016 8008 2056 8040
rect 2088 8008 2128 8040
rect 2160 8008 2200 8040
rect 2232 8008 2272 8040
rect 2304 8008 2344 8040
rect 2376 8008 2416 8040
rect 2448 8008 2488 8040
rect 2520 8008 2560 8040
rect 2592 8008 2632 8040
rect 2664 8008 2704 8040
rect 2736 8008 2776 8040
rect 2808 8008 2848 8040
rect 2880 8008 2920 8040
rect 2952 8008 2992 8040
rect 3024 8008 3064 8040
rect 3096 8008 3136 8040
rect 3168 8008 3208 8040
rect 3240 8008 3280 8040
rect 3312 8008 3352 8040
rect 3384 8008 3424 8040
rect 3456 8008 3496 8040
rect 3528 8008 3568 8040
rect 3600 8008 3640 8040
rect 3672 8008 3712 8040
rect 3744 8008 3784 8040
rect 3816 8008 3856 8040
rect 3888 8008 3928 8040
rect 3960 8008 4000 8040
rect 0 7968 4000 8008
rect 0 7936 40 7968
rect 72 7936 112 7968
rect 144 7936 184 7968
rect 216 7936 256 7968
rect 288 7936 328 7968
rect 360 7936 400 7968
rect 432 7936 472 7968
rect 504 7936 544 7968
rect 576 7936 616 7968
rect 648 7936 688 7968
rect 720 7936 760 7968
rect 792 7936 832 7968
rect 864 7936 904 7968
rect 936 7936 976 7968
rect 1008 7936 1048 7968
rect 1080 7936 1120 7968
rect 1152 7936 1192 7968
rect 1224 7936 1264 7968
rect 1296 7936 1336 7968
rect 1368 7936 1408 7968
rect 1440 7936 1480 7968
rect 1512 7936 1552 7968
rect 1584 7936 1624 7968
rect 1656 7936 1696 7968
rect 1728 7936 1768 7968
rect 1800 7936 1840 7968
rect 1872 7936 1912 7968
rect 1944 7936 1984 7968
rect 2016 7936 2056 7968
rect 2088 7936 2128 7968
rect 2160 7936 2200 7968
rect 2232 7936 2272 7968
rect 2304 7936 2344 7968
rect 2376 7936 2416 7968
rect 2448 7936 2488 7968
rect 2520 7936 2560 7968
rect 2592 7936 2632 7968
rect 2664 7936 2704 7968
rect 2736 7936 2776 7968
rect 2808 7936 2848 7968
rect 2880 7936 2920 7968
rect 2952 7936 2992 7968
rect 3024 7936 3064 7968
rect 3096 7936 3136 7968
rect 3168 7936 3208 7968
rect 3240 7936 3280 7968
rect 3312 7936 3352 7968
rect 3384 7936 3424 7968
rect 3456 7936 3496 7968
rect 3528 7936 3568 7968
rect 3600 7936 3640 7968
rect 3672 7936 3712 7968
rect 3744 7936 3784 7968
rect 3816 7936 3856 7968
rect 3888 7936 3928 7968
rect 3960 7936 4000 7968
rect 0 7896 4000 7936
rect 0 7864 40 7896
rect 72 7864 112 7896
rect 144 7864 184 7896
rect 216 7864 256 7896
rect 288 7864 328 7896
rect 360 7864 400 7896
rect 432 7864 472 7896
rect 504 7864 544 7896
rect 576 7864 616 7896
rect 648 7864 688 7896
rect 720 7864 760 7896
rect 792 7864 832 7896
rect 864 7864 904 7896
rect 936 7864 976 7896
rect 1008 7864 1048 7896
rect 1080 7864 1120 7896
rect 1152 7864 1192 7896
rect 1224 7864 1264 7896
rect 1296 7864 1336 7896
rect 1368 7864 1408 7896
rect 1440 7864 1480 7896
rect 1512 7864 1552 7896
rect 1584 7864 1624 7896
rect 1656 7864 1696 7896
rect 1728 7864 1768 7896
rect 1800 7864 1840 7896
rect 1872 7864 1912 7896
rect 1944 7864 1984 7896
rect 2016 7864 2056 7896
rect 2088 7864 2128 7896
rect 2160 7864 2200 7896
rect 2232 7864 2272 7896
rect 2304 7864 2344 7896
rect 2376 7864 2416 7896
rect 2448 7864 2488 7896
rect 2520 7864 2560 7896
rect 2592 7864 2632 7896
rect 2664 7864 2704 7896
rect 2736 7864 2776 7896
rect 2808 7864 2848 7896
rect 2880 7864 2920 7896
rect 2952 7864 2992 7896
rect 3024 7864 3064 7896
rect 3096 7864 3136 7896
rect 3168 7864 3208 7896
rect 3240 7864 3280 7896
rect 3312 7864 3352 7896
rect 3384 7864 3424 7896
rect 3456 7864 3496 7896
rect 3528 7864 3568 7896
rect 3600 7864 3640 7896
rect 3672 7864 3712 7896
rect 3744 7864 3784 7896
rect 3816 7864 3856 7896
rect 3888 7864 3928 7896
rect 3960 7864 4000 7896
rect 0 7824 4000 7864
rect 0 7792 40 7824
rect 72 7792 112 7824
rect 144 7792 184 7824
rect 216 7792 256 7824
rect 288 7792 328 7824
rect 360 7792 400 7824
rect 432 7792 472 7824
rect 504 7792 544 7824
rect 576 7792 616 7824
rect 648 7792 688 7824
rect 720 7792 760 7824
rect 792 7792 832 7824
rect 864 7792 904 7824
rect 936 7792 976 7824
rect 1008 7792 1048 7824
rect 1080 7792 1120 7824
rect 1152 7792 1192 7824
rect 1224 7792 1264 7824
rect 1296 7792 1336 7824
rect 1368 7792 1408 7824
rect 1440 7792 1480 7824
rect 1512 7792 1552 7824
rect 1584 7792 1624 7824
rect 1656 7792 1696 7824
rect 1728 7792 1768 7824
rect 1800 7792 1840 7824
rect 1872 7792 1912 7824
rect 1944 7792 1984 7824
rect 2016 7792 2056 7824
rect 2088 7792 2128 7824
rect 2160 7792 2200 7824
rect 2232 7792 2272 7824
rect 2304 7792 2344 7824
rect 2376 7792 2416 7824
rect 2448 7792 2488 7824
rect 2520 7792 2560 7824
rect 2592 7792 2632 7824
rect 2664 7792 2704 7824
rect 2736 7792 2776 7824
rect 2808 7792 2848 7824
rect 2880 7792 2920 7824
rect 2952 7792 2992 7824
rect 3024 7792 3064 7824
rect 3096 7792 3136 7824
rect 3168 7792 3208 7824
rect 3240 7792 3280 7824
rect 3312 7792 3352 7824
rect 3384 7792 3424 7824
rect 3456 7792 3496 7824
rect 3528 7792 3568 7824
rect 3600 7792 3640 7824
rect 3672 7792 3712 7824
rect 3744 7792 3784 7824
rect 3816 7792 3856 7824
rect 3888 7792 3928 7824
rect 3960 7792 4000 7824
rect 0 7752 4000 7792
rect 0 7720 40 7752
rect 72 7720 112 7752
rect 144 7720 184 7752
rect 216 7720 256 7752
rect 288 7720 328 7752
rect 360 7720 400 7752
rect 432 7720 472 7752
rect 504 7720 544 7752
rect 576 7720 616 7752
rect 648 7720 688 7752
rect 720 7720 760 7752
rect 792 7720 832 7752
rect 864 7720 904 7752
rect 936 7720 976 7752
rect 1008 7720 1048 7752
rect 1080 7720 1120 7752
rect 1152 7720 1192 7752
rect 1224 7720 1264 7752
rect 1296 7720 1336 7752
rect 1368 7720 1408 7752
rect 1440 7720 1480 7752
rect 1512 7720 1552 7752
rect 1584 7720 1624 7752
rect 1656 7720 1696 7752
rect 1728 7720 1768 7752
rect 1800 7720 1840 7752
rect 1872 7720 1912 7752
rect 1944 7720 1984 7752
rect 2016 7720 2056 7752
rect 2088 7720 2128 7752
rect 2160 7720 2200 7752
rect 2232 7720 2272 7752
rect 2304 7720 2344 7752
rect 2376 7720 2416 7752
rect 2448 7720 2488 7752
rect 2520 7720 2560 7752
rect 2592 7720 2632 7752
rect 2664 7720 2704 7752
rect 2736 7720 2776 7752
rect 2808 7720 2848 7752
rect 2880 7720 2920 7752
rect 2952 7720 2992 7752
rect 3024 7720 3064 7752
rect 3096 7720 3136 7752
rect 3168 7720 3208 7752
rect 3240 7720 3280 7752
rect 3312 7720 3352 7752
rect 3384 7720 3424 7752
rect 3456 7720 3496 7752
rect 3528 7720 3568 7752
rect 3600 7720 3640 7752
rect 3672 7720 3712 7752
rect 3744 7720 3784 7752
rect 3816 7720 3856 7752
rect 3888 7720 3928 7752
rect 3960 7720 4000 7752
rect 0 7680 4000 7720
rect 0 7648 40 7680
rect 72 7648 112 7680
rect 144 7648 184 7680
rect 216 7648 256 7680
rect 288 7648 328 7680
rect 360 7648 400 7680
rect 432 7648 472 7680
rect 504 7648 544 7680
rect 576 7648 616 7680
rect 648 7648 688 7680
rect 720 7648 760 7680
rect 792 7648 832 7680
rect 864 7648 904 7680
rect 936 7648 976 7680
rect 1008 7648 1048 7680
rect 1080 7648 1120 7680
rect 1152 7648 1192 7680
rect 1224 7648 1264 7680
rect 1296 7648 1336 7680
rect 1368 7648 1408 7680
rect 1440 7648 1480 7680
rect 1512 7648 1552 7680
rect 1584 7648 1624 7680
rect 1656 7648 1696 7680
rect 1728 7648 1768 7680
rect 1800 7648 1840 7680
rect 1872 7648 1912 7680
rect 1944 7648 1984 7680
rect 2016 7648 2056 7680
rect 2088 7648 2128 7680
rect 2160 7648 2200 7680
rect 2232 7648 2272 7680
rect 2304 7648 2344 7680
rect 2376 7648 2416 7680
rect 2448 7648 2488 7680
rect 2520 7648 2560 7680
rect 2592 7648 2632 7680
rect 2664 7648 2704 7680
rect 2736 7648 2776 7680
rect 2808 7648 2848 7680
rect 2880 7648 2920 7680
rect 2952 7648 2992 7680
rect 3024 7648 3064 7680
rect 3096 7648 3136 7680
rect 3168 7648 3208 7680
rect 3240 7648 3280 7680
rect 3312 7648 3352 7680
rect 3384 7648 3424 7680
rect 3456 7648 3496 7680
rect 3528 7648 3568 7680
rect 3600 7648 3640 7680
rect 3672 7648 3712 7680
rect 3744 7648 3784 7680
rect 3816 7648 3856 7680
rect 3888 7648 3928 7680
rect 3960 7648 4000 7680
rect 0 7608 4000 7648
rect 0 7576 40 7608
rect 72 7576 112 7608
rect 144 7576 184 7608
rect 216 7576 256 7608
rect 288 7576 328 7608
rect 360 7576 400 7608
rect 432 7576 472 7608
rect 504 7576 544 7608
rect 576 7576 616 7608
rect 648 7576 688 7608
rect 720 7576 760 7608
rect 792 7576 832 7608
rect 864 7576 904 7608
rect 936 7576 976 7608
rect 1008 7576 1048 7608
rect 1080 7576 1120 7608
rect 1152 7576 1192 7608
rect 1224 7576 1264 7608
rect 1296 7576 1336 7608
rect 1368 7576 1408 7608
rect 1440 7576 1480 7608
rect 1512 7576 1552 7608
rect 1584 7576 1624 7608
rect 1656 7576 1696 7608
rect 1728 7576 1768 7608
rect 1800 7576 1840 7608
rect 1872 7576 1912 7608
rect 1944 7576 1984 7608
rect 2016 7576 2056 7608
rect 2088 7576 2128 7608
rect 2160 7576 2200 7608
rect 2232 7576 2272 7608
rect 2304 7576 2344 7608
rect 2376 7576 2416 7608
rect 2448 7576 2488 7608
rect 2520 7576 2560 7608
rect 2592 7576 2632 7608
rect 2664 7576 2704 7608
rect 2736 7576 2776 7608
rect 2808 7576 2848 7608
rect 2880 7576 2920 7608
rect 2952 7576 2992 7608
rect 3024 7576 3064 7608
rect 3096 7576 3136 7608
rect 3168 7576 3208 7608
rect 3240 7576 3280 7608
rect 3312 7576 3352 7608
rect 3384 7576 3424 7608
rect 3456 7576 3496 7608
rect 3528 7576 3568 7608
rect 3600 7576 3640 7608
rect 3672 7576 3712 7608
rect 3744 7576 3784 7608
rect 3816 7576 3856 7608
rect 3888 7576 3928 7608
rect 3960 7576 4000 7608
rect 0 7536 4000 7576
rect 0 7504 40 7536
rect 72 7504 112 7536
rect 144 7504 184 7536
rect 216 7504 256 7536
rect 288 7504 328 7536
rect 360 7504 400 7536
rect 432 7504 472 7536
rect 504 7504 544 7536
rect 576 7504 616 7536
rect 648 7504 688 7536
rect 720 7504 760 7536
rect 792 7504 832 7536
rect 864 7504 904 7536
rect 936 7504 976 7536
rect 1008 7504 1048 7536
rect 1080 7504 1120 7536
rect 1152 7504 1192 7536
rect 1224 7504 1264 7536
rect 1296 7504 1336 7536
rect 1368 7504 1408 7536
rect 1440 7504 1480 7536
rect 1512 7504 1552 7536
rect 1584 7504 1624 7536
rect 1656 7504 1696 7536
rect 1728 7504 1768 7536
rect 1800 7504 1840 7536
rect 1872 7504 1912 7536
rect 1944 7504 1984 7536
rect 2016 7504 2056 7536
rect 2088 7504 2128 7536
rect 2160 7504 2200 7536
rect 2232 7504 2272 7536
rect 2304 7504 2344 7536
rect 2376 7504 2416 7536
rect 2448 7504 2488 7536
rect 2520 7504 2560 7536
rect 2592 7504 2632 7536
rect 2664 7504 2704 7536
rect 2736 7504 2776 7536
rect 2808 7504 2848 7536
rect 2880 7504 2920 7536
rect 2952 7504 2992 7536
rect 3024 7504 3064 7536
rect 3096 7504 3136 7536
rect 3168 7504 3208 7536
rect 3240 7504 3280 7536
rect 3312 7504 3352 7536
rect 3384 7504 3424 7536
rect 3456 7504 3496 7536
rect 3528 7504 3568 7536
rect 3600 7504 3640 7536
rect 3672 7504 3712 7536
rect 3744 7504 3784 7536
rect 3816 7504 3856 7536
rect 3888 7504 3928 7536
rect 3960 7504 4000 7536
rect 0 7464 4000 7504
rect 0 7432 40 7464
rect 72 7432 112 7464
rect 144 7432 184 7464
rect 216 7432 256 7464
rect 288 7432 328 7464
rect 360 7432 400 7464
rect 432 7432 472 7464
rect 504 7432 544 7464
rect 576 7432 616 7464
rect 648 7432 688 7464
rect 720 7432 760 7464
rect 792 7432 832 7464
rect 864 7432 904 7464
rect 936 7432 976 7464
rect 1008 7432 1048 7464
rect 1080 7432 1120 7464
rect 1152 7432 1192 7464
rect 1224 7432 1264 7464
rect 1296 7432 1336 7464
rect 1368 7432 1408 7464
rect 1440 7432 1480 7464
rect 1512 7432 1552 7464
rect 1584 7432 1624 7464
rect 1656 7432 1696 7464
rect 1728 7432 1768 7464
rect 1800 7432 1840 7464
rect 1872 7432 1912 7464
rect 1944 7432 1984 7464
rect 2016 7432 2056 7464
rect 2088 7432 2128 7464
rect 2160 7432 2200 7464
rect 2232 7432 2272 7464
rect 2304 7432 2344 7464
rect 2376 7432 2416 7464
rect 2448 7432 2488 7464
rect 2520 7432 2560 7464
rect 2592 7432 2632 7464
rect 2664 7432 2704 7464
rect 2736 7432 2776 7464
rect 2808 7432 2848 7464
rect 2880 7432 2920 7464
rect 2952 7432 2992 7464
rect 3024 7432 3064 7464
rect 3096 7432 3136 7464
rect 3168 7432 3208 7464
rect 3240 7432 3280 7464
rect 3312 7432 3352 7464
rect 3384 7432 3424 7464
rect 3456 7432 3496 7464
rect 3528 7432 3568 7464
rect 3600 7432 3640 7464
rect 3672 7432 3712 7464
rect 3744 7432 3784 7464
rect 3816 7432 3856 7464
rect 3888 7432 3928 7464
rect 3960 7432 4000 7464
rect 0 7392 4000 7432
rect 0 7360 40 7392
rect 72 7360 112 7392
rect 144 7360 184 7392
rect 216 7360 256 7392
rect 288 7360 328 7392
rect 360 7360 400 7392
rect 432 7360 472 7392
rect 504 7360 544 7392
rect 576 7360 616 7392
rect 648 7360 688 7392
rect 720 7360 760 7392
rect 792 7360 832 7392
rect 864 7360 904 7392
rect 936 7360 976 7392
rect 1008 7360 1048 7392
rect 1080 7360 1120 7392
rect 1152 7360 1192 7392
rect 1224 7360 1264 7392
rect 1296 7360 1336 7392
rect 1368 7360 1408 7392
rect 1440 7360 1480 7392
rect 1512 7360 1552 7392
rect 1584 7360 1624 7392
rect 1656 7360 1696 7392
rect 1728 7360 1768 7392
rect 1800 7360 1840 7392
rect 1872 7360 1912 7392
rect 1944 7360 1984 7392
rect 2016 7360 2056 7392
rect 2088 7360 2128 7392
rect 2160 7360 2200 7392
rect 2232 7360 2272 7392
rect 2304 7360 2344 7392
rect 2376 7360 2416 7392
rect 2448 7360 2488 7392
rect 2520 7360 2560 7392
rect 2592 7360 2632 7392
rect 2664 7360 2704 7392
rect 2736 7360 2776 7392
rect 2808 7360 2848 7392
rect 2880 7360 2920 7392
rect 2952 7360 2992 7392
rect 3024 7360 3064 7392
rect 3096 7360 3136 7392
rect 3168 7360 3208 7392
rect 3240 7360 3280 7392
rect 3312 7360 3352 7392
rect 3384 7360 3424 7392
rect 3456 7360 3496 7392
rect 3528 7360 3568 7392
rect 3600 7360 3640 7392
rect 3672 7360 3712 7392
rect 3744 7360 3784 7392
rect 3816 7360 3856 7392
rect 3888 7360 3928 7392
rect 3960 7360 4000 7392
rect 0 7320 4000 7360
rect 0 7288 40 7320
rect 72 7288 112 7320
rect 144 7288 184 7320
rect 216 7288 256 7320
rect 288 7288 328 7320
rect 360 7288 400 7320
rect 432 7288 472 7320
rect 504 7288 544 7320
rect 576 7288 616 7320
rect 648 7288 688 7320
rect 720 7288 760 7320
rect 792 7288 832 7320
rect 864 7288 904 7320
rect 936 7288 976 7320
rect 1008 7288 1048 7320
rect 1080 7288 1120 7320
rect 1152 7288 1192 7320
rect 1224 7288 1264 7320
rect 1296 7288 1336 7320
rect 1368 7288 1408 7320
rect 1440 7288 1480 7320
rect 1512 7288 1552 7320
rect 1584 7288 1624 7320
rect 1656 7288 1696 7320
rect 1728 7288 1768 7320
rect 1800 7288 1840 7320
rect 1872 7288 1912 7320
rect 1944 7288 1984 7320
rect 2016 7288 2056 7320
rect 2088 7288 2128 7320
rect 2160 7288 2200 7320
rect 2232 7288 2272 7320
rect 2304 7288 2344 7320
rect 2376 7288 2416 7320
rect 2448 7288 2488 7320
rect 2520 7288 2560 7320
rect 2592 7288 2632 7320
rect 2664 7288 2704 7320
rect 2736 7288 2776 7320
rect 2808 7288 2848 7320
rect 2880 7288 2920 7320
rect 2952 7288 2992 7320
rect 3024 7288 3064 7320
rect 3096 7288 3136 7320
rect 3168 7288 3208 7320
rect 3240 7288 3280 7320
rect 3312 7288 3352 7320
rect 3384 7288 3424 7320
rect 3456 7288 3496 7320
rect 3528 7288 3568 7320
rect 3600 7288 3640 7320
rect 3672 7288 3712 7320
rect 3744 7288 3784 7320
rect 3816 7288 3856 7320
rect 3888 7288 3928 7320
rect 3960 7288 4000 7320
rect 0 7248 4000 7288
rect 0 7216 40 7248
rect 72 7216 112 7248
rect 144 7216 184 7248
rect 216 7216 256 7248
rect 288 7216 328 7248
rect 360 7216 400 7248
rect 432 7216 472 7248
rect 504 7216 544 7248
rect 576 7216 616 7248
rect 648 7216 688 7248
rect 720 7216 760 7248
rect 792 7216 832 7248
rect 864 7216 904 7248
rect 936 7216 976 7248
rect 1008 7216 1048 7248
rect 1080 7216 1120 7248
rect 1152 7216 1192 7248
rect 1224 7216 1264 7248
rect 1296 7216 1336 7248
rect 1368 7216 1408 7248
rect 1440 7216 1480 7248
rect 1512 7216 1552 7248
rect 1584 7216 1624 7248
rect 1656 7216 1696 7248
rect 1728 7216 1768 7248
rect 1800 7216 1840 7248
rect 1872 7216 1912 7248
rect 1944 7216 1984 7248
rect 2016 7216 2056 7248
rect 2088 7216 2128 7248
rect 2160 7216 2200 7248
rect 2232 7216 2272 7248
rect 2304 7216 2344 7248
rect 2376 7216 2416 7248
rect 2448 7216 2488 7248
rect 2520 7216 2560 7248
rect 2592 7216 2632 7248
rect 2664 7216 2704 7248
rect 2736 7216 2776 7248
rect 2808 7216 2848 7248
rect 2880 7216 2920 7248
rect 2952 7216 2992 7248
rect 3024 7216 3064 7248
rect 3096 7216 3136 7248
rect 3168 7216 3208 7248
rect 3240 7216 3280 7248
rect 3312 7216 3352 7248
rect 3384 7216 3424 7248
rect 3456 7216 3496 7248
rect 3528 7216 3568 7248
rect 3600 7216 3640 7248
rect 3672 7216 3712 7248
rect 3744 7216 3784 7248
rect 3816 7216 3856 7248
rect 3888 7216 3928 7248
rect 3960 7216 4000 7248
rect 0 7176 4000 7216
rect 0 7144 40 7176
rect 72 7144 112 7176
rect 144 7144 184 7176
rect 216 7144 256 7176
rect 288 7144 328 7176
rect 360 7144 400 7176
rect 432 7144 472 7176
rect 504 7144 544 7176
rect 576 7144 616 7176
rect 648 7144 688 7176
rect 720 7144 760 7176
rect 792 7144 832 7176
rect 864 7144 904 7176
rect 936 7144 976 7176
rect 1008 7144 1048 7176
rect 1080 7144 1120 7176
rect 1152 7144 1192 7176
rect 1224 7144 1264 7176
rect 1296 7144 1336 7176
rect 1368 7144 1408 7176
rect 1440 7144 1480 7176
rect 1512 7144 1552 7176
rect 1584 7144 1624 7176
rect 1656 7144 1696 7176
rect 1728 7144 1768 7176
rect 1800 7144 1840 7176
rect 1872 7144 1912 7176
rect 1944 7144 1984 7176
rect 2016 7144 2056 7176
rect 2088 7144 2128 7176
rect 2160 7144 2200 7176
rect 2232 7144 2272 7176
rect 2304 7144 2344 7176
rect 2376 7144 2416 7176
rect 2448 7144 2488 7176
rect 2520 7144 2560 7176
rect 2592 7144 2632 7176
rect 2664 7144 2704 7176
rect 2736 7144 2776 7176
rect 2808 7144 2848 7176
rect 2880 7144 2920 7176
rect 2952 7144 2992 7176
rect 3024 7144 3064 7176
rect 3096 7144 3136 7176
rect 3168 7144 3208 7176
rect 3240 7144 3280 7176
rect 3312 7144 3352 7176
rect 3384 7144 3424 7176
rect 3456 7144 3496 7176
rect 3528 7144 3568 7176
rect 3600 7144 3640 7176
rect 3672 7144 3712 7176
rect 3744 7144 3784 7176
rect 3816 7144 3856 7176
rect 3888 7144 3928 7176
rect 3960 7144 4000 7176
rect 0 7104 4000 7144
rect 0 7072 40 7104
rect 72 7072 112 7104
rect 144 7072 184 7104
rect 216 7072 256 7104
rect 288 7072 328 7104
rect 360 7072 400 7104
rect 432 7072 472 7104
rect 504 7072 544 7104
rect 576 7072 616 7104
rect 648 7072 688 7104
rect 720 7072 760 7104
rect 792 7072 832 7104
rect 864 7072 904 7104
rect 936 7072 976 7104
rect 1008 7072 1048 7104
rect 1080 7072 1120 7104
rect 1152 7072 1192 7104
rect 1224 7072 1264 7104
rect 1296 7072 1336 7104
rect 1368 7072 1408 7104
rect 1440 7072 1480 7104
rect 1512 7072 1552 7104
rect 1584 7072 1624 7104
rect 1656 7072 1696 7104
rect 1728 7072 1768 7104
rect 1800 7072 1840 7104
rect 1872 7072 1912 7104
rect 1944 7072 1984 7104
rect 2016 7072 2056 7104
rect 2088 7072 2128 7104
rect 2160 7072 2200 7104
rect 2232 7072 2272 7104
rect 2304 7072 2344 7104
rect 2376 7072 2416 7104
rect 2448 7072 2488 7104
rect 2520 7072 2560 7104
rect 2592 7072 2632 7104
rect 2664 7072 2704 7104
rect 2736 7072 2776 7104
rect 2808 7072 2848 7104
rect 2880 7072 2920 7104
rect 2952 7072 2992 7104
rect 3024 7072 3064 7104
rect 3096 7072 3136 7104
rect 3168 7072 3208 7104
rect 3240 7072 3280 7104
rect 3312 7072 3352 7104
rect 3384 7072 3424 7104
rect 3456 7072 3496 7104
rect 3528 7072 3568 7104
rect 3600 7072 3640 7104
rect 3672 7072 3712 7104
rect 3744 7072 3784 7104
rect 3816 7072 3856 7104
rect 3888 7072 3928 7104
rect 3960 7072 4000 7104
rect 0 7032 4000 7072
rect 0 7000 40 7032
rect 72 7000 112 7032
rect 144 7000 184 7032
rect 216 7000 256 7032
rect 288 7000 328 7032
rect 360 7000 400 7032
rect 432 7000 472 7032
rect 504 7000 544 7032
rect 576 7000 616 7032
rect 648 7000 688 7032
rect 720 7000 760 7032
rect 792 7000 832 7032
rect 864 7000 904 7032
rect 936 7000 976 7032
rect 1008 7000 1048 7032
rect 1080 7000 1120 7032
rect 1152 7000 1192 7032
rect 1224 7000 1264 7032
rect 1296 7000 1336 7032
rect 1368 7000 1408 7032
rect 1440 7000 1480 7032
rect 1512 7000 1552 7032
rect 1584 7000 1624 7032
rect 1656 7000 1696 7032
rect 1728 7000 1768 7032
rect 1800 7000 1840 7032
rect 1872 7000 1912 7032
rect 1944 7000 1984 7032
rect 2016 7000 2056 7032
rect 2088 7000 2128 7032
rect 2160 7000 2200 7032
rect 2232 7000 2272 7032
rect 2304 7000 2344 7032
rect 2376 7000 2416 7032
rect 2448 7000 2488 7032
rect 2520 7000 2560 7032
rect 2592 7000 2632 7032
rect 2664 7000 2704 7032
rect 2736 7000 2776 7032
rect 2808 7000 2848 7032
rect 2880 7000 2920 7032
rect 2952 7000 2992 7032
rect 3024 7000 3064 7032
rect 3096 7000 3136 7032
rect 3168 7000 3208 7032
rect 3240 7000 3280 7032
rect 3312 7000 3352 7032
rect 3384 7000 3424 7032
rect 3456 7000 3496 7032
rect 3528 7000 3568 7032
rect 3600 7000 3640 7032
rect 3672 7000 3712 7032
rect 3744 7000 3784 7032
rect 3816 7000 3856 7032
rect 3888 7000 3928 7032
rect 3960 7000 4000 7032
rect 0 6960 4000 7000
rect 0 6928 40 6960
rect 72 6928 112 6960
rect 144 6928 184 6960
rect 216 6928 256 6960
rect 288 6928 328 6960
rect 360 6928 400 6960
rect 432 6928 472 6960
rect 504 6928 544 6960
rect 576 6928 616 6960
rect 648 6928 688 6960
rect 720 6928 760 6960
rect 792 6928 832 6960
rect 864 6928 904 6960
rect 936 6928 976 6960
rect 1008 6928 1048 6960
rect 1080 6928 1120 6960
rect 1152 6928 1192 6960
rect 1224 6928 1264 6960
rect 1296 6928 1336 6960
rect 1368 6928 1408 6960
rect 1440 6928 1480 6960
rect 1512 6928 1552 6960
rect 1584 6928 1624 6960
rect 1656 6928 1696 6960
rect 1728 6928 1768 6960
rect 1800 6928 1840 6960
rect 1872 6928 1912 6960
rect 1944 6928 1984 6960
rect 2016 6928 2056 6960
rect 2088 6928 2128 6960
rect 2160 6928 2200 6960
rect 2232 6928 2272 6960
rect 2304 6928 2344 6960
rect 2376 6928 2416 6960
rect 2448 6928 2488 6960
rect 2520 6928 2560 6960
rect 2592 6928 2632 6960
rect 2664 6928 2704 6960
rect 2736 6928 2776 6960
rect 2808 6928 2848 6960
rect 2880 6928 2920 6960
rect 2952 6928 2992 6960
rect 3024 6928 3064 6960
rect 3096 6928 3136 6960
rect 3168 6928 3208 6960
rect 3240 6928 3280 6960
rect 3312 6928 3352 6960
rect 3384 6928 3424 6960
rect 3456 6928 3496 6960
rect 3528 6928 3568 6960
rect 3600 6928 3640 6960
rect 3672 6928 3712 6960
rect 3744 6928 3784 6960
rect 3816 6928 3856 6960
rect 3888 6928 3928 6960
rect 3960 6928 4000 6960
rect 0 6888 4000 6928
rect 0 6856 40 6888
rect 72 6856 112 6888
rect 144 6856 184 6888
rect 216 6856 256 6888
rect 288 6856 328 6888
rect 360 6856 400 6888
rect 432 6856 472 6888
rect 504 6856 544 6888
rect 576 6856 616 6888
rect 648 6856 688 6888
rect 720 6856 760 6888
rect 792 6856 832 6888
rect 864 6856 904 6888
rect 936 6856 976 6888
rect 1008 6856 1048 6888
rect 1080 6856 1120 6888
rect 1152 6856 1192 6888
rect 1224 6856 1264 6888
rect 1296 6856 1336 6888
rect 1368 6856 1408 6888
rect 1440 6856 1480 6888
rect 1512 6856 1552 6888
rect 1584 6856 1624 6888
rect 1656 6856 1696 6888
rect 1728 6856 1768 6888
rect 1800 6856 1840 6888
rect 1872 6856 1912 6888
rect 1944 6856 1984 6888
rect 2016 6856 2056 6888
rect 2088 6856 2128 6888
rect 2160 6856 2200 6888
rect 2232 6856 2272 6888
rect 2304 6856 2344 6888
rect 2376 6856 2416 6888
rect 2448 6856 2488 6888
rect 2520 6856 2560 6888
rect 2592 6856 2632 6888
rect 2664 6856 2704 6888
rect 2736 6856 2776 6888
rect 2808 6856 2848 6888
rect 2880 6856 2920 6888
rect 2952 6856 2992 6888
rect 3024 6856 3064 6888
rect 3096 6856 3136 6888
rect 3168 6856 3208 6888
rect 3240 6856 3280 6888
rect 3312 6856 3352 6888
rect 3384 6856 3424 6888
rect 3456 6856 3496 6888
rect 3528 6856 3568 6888
rect 3600 6856 3640 6888
rect 3672 6856 3712 6888
rect 3744 6856 3784 6888
rect 3816 6856 3856 6888
rect 3888 6856 3928 6888
rect 3960 6856 4000 6888
rect 0 6800 4000 6856
rect 0 6544 4000 6600
rect 0 6512 40 6544
rect 72 6512 112 6544
rect 144 6512 184 6544
rect 216 6512 256 6544
rect 288 6512 328 6544
rect 360 6512 400 6544
rect 432 6512 472 6544
rect 504 6512 544 6544
rect 576 6512 616 6544
rect 648 6512 688 6544
rect 720 6512 760 6544
rect 792 6512 832 6544
rect 864 6512 904 6544
rect 936 6512 976 6544
rect 1008 6512 1048 6544
rect 1080 6512 1120 6544
rect 1152 6512 1192 6544
rect 1224 6512 1264 6544
rect 1296 6512 1336 6544
rect 1368 6512 1408 6544
rect 1440 6512 1480 6544
rect 1512 6512 1552 6544
rect 1584 6512 1624 6544
rect 1656 6512 1696 6544
rect 1728 6512 1768 6544
rect 1800 6512 1840 6544
rect 1872 6512 1912 6544
rect 1944 6512 1984 6544
rect 2016 6512 2056 6544
rect 2088 6512 2128 6544
rect 2160 6512 2200 6544
rect 2232 6512 2272 6544
rect 2304 6512 2344 6544
rect 2376 6512 2416 6544
rect 2448 6512 2488 6544
rect 2520 6512 2560 6544
rect 2592 6512 2632 6544
rect 2664 6512 2704 6544
rect 2736 6512 2776 6544
rect 2808 6512 2848 6544
rect 2880 6512 2920 6544
rect 2952 6512 2992 6544
rect 3024 6512 3064 6544
rect 3096 6512 3136 6544
rect 3168 6512 3208 6544
rect 3240 6512 3280 6544
rect 3312 6512 3352 6544
rect 3384 6512 3424 6544
rect 3456 6512 3496 6544
rect 3528 6512 3568 6544
rect 3600 6512 3640 6544
rect 3672 6512 3712 6544
rect 3744 6512 3784 6544
rect 3816 6512 3856 6544
rect 3888 6512 3928 6544
rect 3960 6512 4000 6544
rect 0 6472 4000 6512
rect 0 6440 40 6472
rect 72 6440 112 6472
rect 144 6440 184 6472
rect 216 6440 256 6472
rect 288 6440 328 6472
rect 360 6440 400 6472
rect 432 6440 472 6472
rect 504 6440 544 6472
rect 576 6440 616 6472
rect 648 6440 688 6472
rect 720 6440 760 6472
rect 792 6440 832 6472
rect 864 6440 904 6472
rect 936 6440 976 6472
rect 1008 6440 1048 6472
rect 1080 6440 1120 6472
rect 1152 6440 1192 6472
rect 1224 6440 1264 6472
rect 1296 6440 1336 6472
rect 1368 6440 1408 6472
rect 1440 6440 1480 6472
rect 1512 6440 1552 6472
rect 1584 6440 1624 6472
rect 1656 6440 1696 6472
rect 1728 6440 1768 6472
rect 1800 6440 1840 6472
rect 1872 6440 1912 6472
rect 1944 6440 1984 6472
rect 2016 6440 2056 6472
rect 2088 6440 2128 6472
rect 2160 6440 2200 6472
rect 2232 6440 2272 6472
rect 2304 6440 2344 6472
rect 2376 6440 2416 6472
rect 2448 6440 2488 6472
rect 2520 6440 2560 6472
rect 2592 6440 2632 6472
rect 2664 6440 2704 6472
rect 2736 6440 2776 6472
rect 2808 6440 2848 6472
rect 2880 6440 2920 6472
rect 2952 6440 2992 6472
rect 3024 6440 3064 6472
rect 3096 6440 3136 6472
rect 3168 6440 3208 6472
rect 3240 6440 3280 6472
rect 3312 6440 3352 6472
rect 3384 6440 3424 6472
rect 3456 6440 3496 6472
rect 3528 6440 3568 6472
rect 3600 6440 3640 6472
rect 3672 6440 3712 6472
rect 3744 6440 3784 6472
rect 3816 6440 3856 6472
rect 3888 6440 3928 6472
rect 3960 6440 4000 6472
rect 0 6400 4000 6440
rect 0 6368 40 6400
rect 72 6368 112 6400
rect 144 6368 184 6400
rect 216 6368 256 6400
rect 288 6368 328 6400
rect 360 6368 400 6400
rect 432 6368 472 6400
rect 504 6368 544 6400
rect 576 6368 616 6400
rect 648 6368 688 6400
rect 720 6368 760 6400
rect 792 6368 832 6400
rect 864 6368 904 6400
rect 936 6368 976 6400
rect 1008 6368 1048 6400
rect 1080 6368 1120 6400
rect 1152 6368 1192 6400
rect 1224 6368 1264 6400
rect 1296 6368 1336 6400
rect 1368 6368 1408 6400
rect 1440 6368 1480 6400
rect 1512 6368 1552 6400
rect 1584 6368 1624 6400
rect 1656 6368 1696 6400
rect 1728 6368 1768 6400
rect 1800 6368 1840 6400
rect 1872 6368 1912 6400
rect 1944 6368 1984 6400
rect 2016 6368 2056 6400
rect 2088 6368 2128 6400
rect 2160 6368 2200 6400
rect 2232 6368 2272 6400
rect 2304 6368 2344 6400
rect 2376 6368 2416 6400
rect 2448 6368 2488 6400
rect 2520 6368 2560 6400
rect 2592 6368 2632 6400
rect 2664 6368 2704 6400
rect 2736 6368 2776 6400
rect 2808 6368 2848 6400
rect 2880 6368 2920 6400
rect 2952 6368 2992 6400
rect 3024 6368 3064 6400
rect 3096 6368 3136 6400
rect 3168 6368 3208 6400
rect 3240 6368 3280 6400
rect 3312 6368 3352 6400
rect 3384 6368 3424 6400
rect 3456 6368 3496 6400
rect 3528 6368 3568 6400
rect 3600 6368 3640 6400
rect 3672 6368 3712 6400
rect 3744 6368 3784 6400
rect 3816 6368 3856 6400
rect 3888 6368 3928 6400
rect 3960 6368 4000 6400
rect 0 6328 4000 6368
rect 0 6296 40 6328
rect 72 6296 112 6328
rect 144 6296 184 6328
rect 216 6296 256 6328
rect 288 6296 328 6328
rect 360 6296 400 6328
rect 432 6296 472 6328
rect 504 6296 544 6328
rect 576 6296 616 6328
rect 648 6296 688 6328
rect 720 6296 760 6328
rect 792 6296 832 6328
rect 864 6296 904 6328
rect 936 6296 976 6328
rect 1008 6296 1048 6328
rect 1080 6296 1120 6328
rect 1152 6296 1192 6328
rect 1224 6296 1264 6328
rect 1296 6296 1336 6328
rect 1368 6296 1408 6328
rect 1440 6296 1480 6328
rect 1512 6296 1552 6328
rect 1584 6296 1624 6328
rect 1656 6296 1696 6328
rect 1728 6296 1768 6328
rect 1800 6296 1840 6328
rect 1872 6296 1912 6328
rect 1944 6296 1984 6328
rect 2016 6296 2056 6328
rect 2088 6296 2128 6328
rect 2160 6296 2200 6328
rect 2232 6296 2272 6328
rect 2304 6296 2344 6328
rect 2376 6296 2416 6328
rect 2448 6296 2488 6328
rect 2520 6296 2560 6328
rect 2592 6296 2632 6328
rect 2664 6296 2704 6328
rect 2736 6296 2776 6328
rect 2808 6296 2848 6328
rect 2880 6296 2920 6328
rect 2952 6296 2992 6328
rect 3024 6296 3064 6328
rect 3096 6296 3136 6328
rect 3168 6296 3208 6328
rect 3240 6296 3280 6328
rect 3312 6296 3352 6328
rect 3384 6296 3424 6328
rect 3456 6296 3496 6328
rect 3528 6296 3568 6328
rect 3600 6296 3640 6328
rect 3672 6296 3712 6328
rect 3744 6296 3784 6328
rect 3816 6296 3856 6328
rect 3888 6296 3928 6328
rect 3960 6296 4000 6328
rect 0 6256 4000 6296
rect 0 6224 40 6256
rect 72 6224 112 6256
rect 144 6224 184 6256
rect 216 6224 256 6256
rect 288 6224 328 6256
rect 360 6224 400 6256
rect 432 6224 472 6256
rect 504 6224 544 6256
rect 576 6224 616 6256
rect 648 6224 688 6256
rect 720 6224 760 6256
rect 792 6224 832 6256
rect 864 6224 904 6256
rect 936 6224 976 6256
rect 1008 6224 1048 6256
rect 1080 6224 1120 6256
rect 1152 6224 1192 6256
rect 1224 6224 1264 6256
rect 1296 6224 1336 6256
rect 1368 6224 1408 6256
rect 1440 6224 1480 6256
rect 1512 6224 1552 6256
rect 1584 6224 1624 6256
rect 1656 6224 1696 6256
rect 1728 6224 1768 6256
rect 1800 6224 1840 6256
rect 1872 6224 1912 6256
rect 1944 6224 1984 6256
rect 2016 6224 2056 6256
rect 2088 6224 2128 6256
rect 2160 6224 2200 6256
rect 2232 6224 2272 6256
rect 2304 6224 2344 6256
rect 2376 6224 2416 6256
rect 2448 6224 2488 6256
rect 2520 6224 2560 6256
rect 2592 6224 2632 6256
rect 2664 6224 2704 6256
rect 2736 6224 2776 6256
rect 2808 6224 2848 6256
rect 2880 6224 2920 6256
rect 2952 6224 2992 6256
rect 3024 6224 3064 6256
rect 3096 6224 3136 6256
rect 3168 6224 3208 6256
rect 3240 6224 3280 6256
rect 3312 6224 3352 6256
rect 3384 6224 3424 6256
rect 3456 6224 3496 6256
rect 3528 6224 3568 6256
rect 3600 6224 3640 6256
rect 3672 6224 3712 6256
rect 3744 6224 3784 6256
rect 3816 6224 3856 6256
rect 3888 6224 3928 6256
rect 3960 6224 4000 6256
rect 0 6184 4000 6224
rect 0 6152 40 6184
rect 72 6152 112 6184
rect 144 6152 184 6184
rect 216 6152 256 6184
rect 288 6152 328 6184
rect 360 6152 400 6184
rect 432 6152 472 6184
rect 504 6152 544 6184
rect 576 6152 616 6184
rect 648 6152 688 6184
rect 720 6152 760 6184
rect 792 6152 832 6184
rect 864 6152 904 6184
rect 936 6152 976 6184
rect 1008 6152 1048 6184
rect 1080 6152 1120 6184
rect 1152 6152 1192 6184
rect 1224 6152 1264 6184
rect 1296 6152 1336 6184
rect 1368 6152 1408 6184
rect 1440 6152 1480 6184
rect 1512 6152 1552 6184
rect 1584 6152 1624 6184
rect 1656 6152 1696 6184
rect 1728 6152 1768 6184
rect 1800 6152 1840 6184
rect 1872 6152 1912 6184
rect 1944 6152 1984 6184
rect 2016 6152 2056 6184
rect 2088 6152 2128 6184
rect 2160 6152 2200 6184
rect 2232 6152 2272 6184
rect 2304 6152 2344 6184
rect 2376 6152 2416 6184
rect 2448 6152 2488 6184
rect 2520 6152 2560 6184
rect 2592 6152 2632 6184
rect 2664 6152 2704 6184
rect 2736 6152 2776 6184
rect 2808 6152 2848 6184
rect 2880 6152 2920 6184
rect 2952 6152 2992 6184
rect 3024 6152 3064 6184
rect 3096 6152 3136 6184
rect 3168 6152 3208 6184
rect 3240 6152 3280 6184
rect 3312 6152 3352 6184
rect 3384 6152 3424 6184
rect 3456 6152 3496 6184
rect 3528 6152 3568 6184
rect 3600 6152 3640 6184
rect 3672 6152 3712 6184
rect 3744 6152 3784 6184
rect 3816 6152 3856 6184
rect 3888 6152 3928 6184
rect 3960 6152 4000 6184
rect 0 6112 4000 6152
rect 0 6080 40 6112
rect 72 6080 112 6112
rect 144 6080 184 6112
rect 216 6080 256 6112
rect 288 6080 328 6112
rect 360 6080 400 6112
rect 432 6080 472 6112
rect 504 6080 544 6112
rect 576 6080 616 6112
rect 648 6080 688 6112
rect 720 6080 760 6112
rect 792 6080 832 6112
rect 864 6080 904 6112
rect 936 6080 976 6112
rect 1008 6080 1048 6112
rect 1080 6080 1120 6112
rect 1152 6080 1192 6112
rect 1224 6080 1264 6112
rect 1296 6080 1336 6112
rect 1368 6080 1408 6112
rect 1440 6080 1480 6112
rect 1512 6080 1552 6112
rect 1584 6080 1624 6112
rect 1656 6080 1696 6112
rect 1728 6080 1768 6112
rect 1800 6080 1840 6112
rect 1872 6080 1912 6112
rect 1944 6080 1984 6112
rect 2016 6080 2056 6112
rect 2088 6080 2128 6112
rect 2160 6080 2200 6112
rect 2232 6080 2272 6112
rect 2304 6080 2344 6112
rect 2376 6080 2416 6112
rect 2448 6080 2488 6112
rect 2520 6080 2560 6112
rect 2592 6080 2632 6112
rect 2664 6080 2704 6112
rect 2736 6080 2776 6112
rect 2808 6080 2848 6112
rect 2880 6080 2920 6112
rect 2952 6080 2992 6112
rect 3024 6080 3064 6112
rect 3096 6080 3136 6112
rect 3168 6080 3208 6112
rect 3240 6080 3280 6112
rect 3312 6080 3352 6112
rect 3384 6080 3424 6112
rect 3456 6080 3496 6112
rect 3528 6080 3568 6112
rect 3600 6080 3640 6112
rect 3672 6080 3712 6112
rect 3744 6080 3784 6112
rect 3816 6080 3856 6112
rect 3888 6080 3928 6112
rect 3960 6080 4000 6112
rect 0 6040 4000 6080
rect 0 6008 40 6040
rect 72 6008 112 6040
rect 144 6008 184 6040
rect 216 6008 256 6040
rect 288 6008 328 6040
rect 360 6008 400 6040
rect 432 6008 472 6040
rect 504 6008 544 6040
rect 576 6008 616 6040
rect 648 6008 688 6040
rect 720 6008 760 6040
rect 792 6008 832 6040
rect 864 6008 904 6040
rect 936 6008 976 6040
rect 1008 6008 1048 6040
rect 1080 6008 1120 6040
rect 1152 6008 1192 6040
rect 1224 6008 1264 6040
rect 1296 6008 1336 6040
rect 1368 6008 1408 6040
rect 1440 6008 1480 6040
rect 1512 6008 1552 6040
rect 1584 6008 1624 6040
rect 1656 6008 1696 6040
rect 1728 6008 1768 6040
rect 1800 6008 1840 6040
rect 1872 6008 1912 6040
rect 1944 6008 1984 6040
rect 2016 6008 2056 6040
rect 2088 6008 2128 6040
rect 2160 6008 2200 6040
rect 2232 6008 2272 6040
rect 2304 6008 2344 6040
rect 2376 6008 2416 6040
rect 2448 6008 2488 6040
rect 2520 6008 2560 6040
rect 2592 6008 2632 6040
rect 2664 6008 2704 6040
rect 2736 6008 2776 6040
rect 2808 6008 2848 6040
rect 2880 6008 2920 6040
rect 2952 6008 2992 6040
rect 3024 6008 3064 6040
rect 3096 6008 3136 6040
rect 3168 6008 3208 6040
rect 3240 6008 3280 6040
rect 3312 6008 3352 6040
rect 3384 6008 3424 6040
rect 3456 6008 3496 6040
rect 3528 6008 3568 6040
rect 3600 6008 3640 6040
rect 3672 6008 3712 6040
rect 3744 6008 3784 6040
rect 3816 6008 3856 6040
rect 3888 6008 3928 6040
rect 3960 6008 4000 6040
rect 0 5968 4000 6008
rect 0 5936 40 5968
rect 72 5936 112 5968
rect 144 5936 184 5968
rect 216 5936 256 5968
rect 288 5936 328 5968
rect 360 5936 400 5968
rect 432 5936 472 5968
rect 504 5936 544 5968
rect 576 5936 616 5968
rect 648 5936 688 5968
rect 720 5936 760 5968
rect 792 5936 832 5968
rect 864 5936 904 5968
rect 936 5936 976 5968
rect 1008 5936 1048 5968
rect 1080 5936 1120 5968
rect 1152 5936 1192 5968
rect 1224 5936 1264 5968
rect 1296 5936 1336 5968
rect 1368 5936 1408 5968
rect 1440 5936 1480 5968
rect 1512 5936 1552 5968
rect 1584 5936 1624 5968
rect 1656 5936 1696 5968
rect 1728 5936 1768 5968
rect 1800 5936 1840 5968
rect 1872 5936 1912 5968
rect 1944 5936 1984 5968
rect 2016 5936 2056 5968
rect 2088 5936 2128 5968
rect 2160 5936 2200 5968
rect 2232 5936 2272 5968
rect 2304 5936 2344 5968
rect 2376 5936 2416 5968
rect 2448 5936 2488 5968
rect 2520 5936 2560 5968
rect 2592 5936 2632 5968
rect 2664 5936 2704 5968
rect 2736 5936 2776 5968
rect 2808 5936 2848 5968
rect 2880 5936 2920 5968
rect 2952 5936 2992 5968
rect 3024 5936 3064 5968
rect 3096 5936 3136 5968
rect 3168 5936 3208 5968
rect 3240 5936 3280 5968
rect 3312 5936 3352 5968
rect 3384 5936 3424 5968
rect 3456 5936 3496 5968
rect 3528 5936 3568 5968
rect 3600 5936 3640 5968
rect 3672 5936 3712 5968
rect 3744 5936 3784 5968
rect 3816 5936 3856 5968
rect 3888 5936 3928 5968
rect 3960 5936 4000 5968
rect 0 5896 4000 5936
rect 0 5864 40 5896
rect 72 5864 112 5896
rect 144 5864 184 5896
rect 216 5864 256 5896
rect 288 5864 328 5896
rect 360 5864 400 5896
rect 432 5864 472 5896
rect 504 5864 544 5896
rect 576 5864 616 5896
rect 648 5864 688 5896
rect 720 5864 760 5896
rect 792 5864 832 5896
rect 864 5864 904 5896
rect 936 5864 976 5896
rect 1008 5864 1048 5896
rect 1080 5864 1120 5896
rect 1152 5864 1192 5896
rect 1224 5864 1264 5896
rect 1296 5864 1336 5896
rect 1368 5864 1408 5896
rect 1440 5864 1480 5896
rect 1512 5864 1552 5896
rect 1584 5864 1624 5896
rect 1656 5864 1696 5896
rect 1728 5864 1768 5896
rect 1800 5864 1840 5896
rect 1872 5864 1912 5896
rect 1944 5864 1984 5896
rect 2016 5864 2056 5896
rect 2088 5864 2128 5896
rect 2160 5864 2200 5896
rect 2232 5864 2272 5896
rect 2304 5864 2344 5896
rect 2376 5864 2416 5896
rect 2448 5864 2488 5896
rect 2520 5864 2560 5896
rect 2592 5864 2632 5896
rect 2664 5864 2704 5896
rect 2736 5864 2776 5896
rect 2808 5864 2848 5896
rect 2880 5864 2920 5896
rect 2952 5864 2992 5896
rect 3024 5864 3064 5896
rect 3096 5864 3136 5896
rect 3168 5864 3208 5896
rect 3240 5864 3280 5896
rect 3312 5864 3352 5896
rect 3384 5864 3424 5896
rect 3456 5864 3496 5896
rect 3528 5864 3568 5896
rect 3600 5864 3640 5896
rect 3672 5864 3712 5896
rect 3744 5864 3784 5896
rect 3816 5864 3856 5896
rect 3888 5864 3928 5896
rect 3960 5864 4000 5896
rect 0 5824 4000 5864
rect 0 5792 40 5824
rect 72 5792 112 5824
rect 144 5792 184 5824
rect 216 5792 256 5824
rect 288 5792 328 5824
rect 360 5792 400 5824
rect 432 5792 472 5824
rect 504 5792 544 5824
rect 576 5792 616 5824
rect 648 5792 688 5824
rect 720 5792 760 5824
rect 792 5792 832 5824
rect 864 5792 904 5824
rect 936 5792 976 5824
rect 1008 5792 1048 5824
rect 1080 5792 1120 5824
rect 1152 5792 1192 5824
rect 1224 5792 1264 5824
rect 1296 5792 1336 5824
rect 1368 5792 1408 5824
rect 1440 5792 1480 5824
rect 1512 5792 1552 5824
rect 1584 5792 1624 5824
rect 1656 5792 1696 5824
rect 1728 5792 1768 5824
rect 1800 5792 1840 5824
rect 1872 5792 1912 5824
rect 1944 5792 1984 5824
rect 2016 5792 2056 5824
rect 2088 5792 2128 5824
rect 2160 5792 2200 5824
rect 2232 5792 2272 5824
rect 2304 5792 2344 5824
rect 2376 5792 2416 5824
rect 2448 5792 2488 5824
rect 2520 5792 2560 5824
rect 2592 5792 2632 5824
rect 2664 5792 2704 5824
rect 2736 5792 2776 5824
rect 2808 5792 2848 5824
rect 2880 5792 2920 5824
rect 2952 5792 2992 5824
rect 3024 5792 3064 5824
rect 3096 5792 3136 5824
rect 3168 5792 3208 5824
rect 3240 5792 3280 5824
rect 3312 5792 3352 5824
rect 3384 5792 3424 5824
rect 3456 5792 3496 5824
rect 3528 5792 3568 5824
rect 3600 5792 3640 5824
rect 3672 5792 3712 5824
rect 3744 5792 3784 5824
rect 3816 5792 3856 5824
rect 3888 5792 3928 5824
rect 3960 5792 4000 5824
rect 0 5752 4000 5792
rect 0 5720 40 5752
rect 72 5720 112 5752
rect 144 5720 184 5752
rect 216 5720 256 5752
rect 288 5720 328 5752
rect 360 5720 400 5752
rect 432 5720 472 5752
rect 504 5720 544 5752
rect 576 5720 616 5752
rect 648 5720 688 5752
rect 720 5720 760 5752
rect 792 5720 832 5752
rect 864 5720 904 5752
rect 936 5720 976 5752
rect 1008 5720 1048 5752
rect 1080 5720 1120 5752
rect 1152 5720 1192 5752
rect 1224 5720 1264 5752
rect 1296 5720 1336 5752
rect 1368 5720 1408 5752
rect 1440 5720 1480 5752
rect 1512 5720 1552 5752
rect 1584 5720 1624 5752
rect 1656 5720 1696 5752
rect 1728 5720 1768 5752
rect 1800 5720 1840 5752
rect 1872 5720 1912 5752
rect 1944 5720 1984 5752
rect 2016 5720 2056 5752
rect 2088 5720 2128 5752
rect 2160 5720 2200 5752
rect 2232 5720 2272 5752
rect 2304 5720 2344 5752
rect 2376 5720 2416 5752
rect 2448 5720 2488 5752
rect 2520 5720 2560 5752
rect 2592 5720 2632 5752
rect 2664 5720 2704 5752
rect 2736 5720 2776 5752
rect 2808 5720 2848 5752
rect 2880 5720 2920 5752
rect 2952 5720 2992 5752
rect 3024 5720 3064 5752
rect 3096 5720 3136 5752
rect 3168 5720 3208 5752
rect 3240 5720 3280 5752
rect 3312 5720 3352 5752
rect 3384 5720 3424 5752
rect 3456 5720 3496 5752
rect 3528 5720 3568 5752
rect 3600 5720 3640 5752
rect 3672 5720 3712 5752
rect 3744 5720 3784 5752
rect 3816 5720 3856 5752
rect 3888 5720 3928 5752
rect 3960 5720 4000 5752
rect 0 5680 4000 5720
rect 0 5648 40 5680
rect 72 5648 112 5680
rect 144 5648 184 5680
rect 216 5648 256 5680
rect 288 5648 328 5680
rect 360 5648 400 5680
rect 432 5648 472 5680
rect 504 5648 544 5680
rect 576 5648 616 5680
rect 648 5648 688 5680
rect 720 5648 760 5680
rect 792 5648 832 5680
rect 864 5648 904 5680
rect 936 5648 976 5680
rect 1008 5648 1048 5680
rect 1080 5648 1120 5680
rect 1152 5648 1192 5680
rect 1224 5648 1264 5680
rect 1296 5648 1336 5680
rect 1368 5648 1408 5680
rect 1440 5648 1480 5680
rect 1512 5648 1552 5680
rect 1584 5648 1624 5680
rect 1656 5648 1696 5680
rect 1728 5648 1768 5680
rect 1800 5648 1840 5680
rect 1872 5648 1912 5680
rect 1944 5648 1984 5680
rect 2016 5648 2056 5680
rect 2088 5648 2128 5680
rect 2160 5648 2200 5680
rect 2232 5648 2272 5680
rect 2304 5648 2344 5680
rect 2376 5648 2416 5680
rect 2448 5648 2488 5680
rect 2520 5648 2560 5680
rect 2592 5648 2632 5680
rect 2664 5648 2704 5680
rect 2736 5648 2776 5680
rect 2808 5648 2848 5680
rect 2880 5648 2920 5680
rect 2952 5648 2992 5680
rect 3024 5648 3064 5680
rect 3096 5648 3136 5680
rect 3168 5648 3208 5680
rect 3240 5648 3280 5680
rect 3312 5648 3352 5680
rect 3384 5648 3424 5680
rect 3456 5648 3496 5680
rect 3528 5648 3568 5680
rect 3600 5648 3640 5680
rect 3672 5648 3712 5680
rect 3744 5648 3784 5680
rect 3816 5648 3856 5680
rect 3888 5648 3928 5680
rect 3960 5648 4000 5680
rect 0 5608 4000 5648
rect 0 5576 40 5608
rect 72 5576 112 5608
rect 144 5576 184 5608
rect 216 5576 256 5608
rect 288 5576 328 5608
rect 360 5576 400 5608
rect 432 5576 472 5608
rect 504 5576 544 5608
rect 576 5576 616 5608
rect 648 5576 688 5608
rect 720 5576 760 5608
rect 792 5576 832 5608
rect 864 5576 904 5608
rect 936 5576 976 5608
rect 1008 5576 1048 5608
rect 1080 5576 1120 5608
rect 1152 5576 1192 5608
rect 1224 5576 1264 5608
rect 1296 5576 1336 5608
rect 1368 5576 1408 5608
rect 1440 5576 1480 5608
rect 1512 5576 1552 5608
rect 1584 5576 1624 5608
rect 1656 5576 1696 5608
rect 1728 5576 1768 5608
rect 1800 5576 1840 5608
rect 1872 5576 1912 5608
rect 1944 5576 1984 5608
rect 2016 5576 2056 5608
rect 2088 5576 2128 5608
rect 2160 5576 2200 5608
rect 2232 5576 2272 5608
rect 2304 5576 2344 5608
rect 2376 5576 2416 5608
rect 2448 5576 2488 5608
rect 2520 5576 2560 5608
rect 2592 5576 2632 5608
rect 2664 5576 2704 5608
rect 2736 5576 2776 5608
rect 2808 5576 2848 5608
rect 2880 5576 2920 5608
rect 2952 5576 2992 5608
rect 3024 5576 3064 5608
rect 3096 5576 3136 5608
rect 3168 5576 3208 5608
rect 3240 5576 3280 5608
rect 3312 5576 3352 5608
rect 3384 5576 3424 5608
rect 3456 5576 3496 5608
rect 3528 5576 3568 5608
rect 3600 5576 3640 5608
rect 3672 5576 3712 5608
rect 3744 5576 3784 5608
rect 3816 5576 3856 5608
rect 3888 5576 3928 5608
rect 3960 5576 4000 5608
rect 0 5536 4000 5576
rect 0 5504 40 5536
rect 72 5504 112 5536
rect 144 5504 184 5536
rect 216 5504 256 5536
rect 288 5504 328 5536
rect 360 5504 400 5536
rect 432 5504 472 5536
rect 504 5504 544 5536
rect 576 5504 616 5536
rect 648 5504 688 5536
rect 720 5504 760 5536
rect 792 5504 832 5536
rect 864 5504 904 5536
rect 936 5504 976 5536
rect 1008 5504 1048 5536
rect 1080 5504 1120 5536
rect 1152 5504 1192 5536
rect 1224 5504 1264 5536
rect 1296 5504 1336 5536
rect 1368 5504 1408 5536
rect 1440 5504 1480 5536
rect 1512 5504 1552 5536
rect 1584 5504 1624 5536
rect 1656 5504 1696 5536
rect 1728 5504 1768 5536
rect 1800 5504 1840 5536
rect 1872 5504 1912 5536
rect 1944 5504 1984 5536
rect 2016 5504 2056 5536
rect 2088 5504 2128 5536
rect 2160 5504 2200 5536
rect 2232 5504 2272 5536
rect 2304 5504 2344 5536
rect 2376 5504 2416 5536
rect 2448 5504 2488 5536
rect 2520 5504 2560 5536
rect 2592 5504 2632 5536
rect 2664 5504 2704 5536
rect 2736 5504 2776 5536
rect 2808 5504 2848 5536
rect 2880 5504 2920 5536
rect 2952 5504 2992 5536
rect 3024 5504 3064 5536
rect 3096 5504 3136 5536
rect 3168 5504 3208 5536
rect 3240 5504 3280 5536
rect 3312 5504 3352 5536
rect 3384 5504 3424 5536
rect 3456 5504 3496 5536
rect 3528 5504 3568 5536
rect 3600 5504 3640 5536
rect 3672 5504 3712 5536
rect 3744 5504 3784 5536
rect 3816 5504 3856 5536
rect 3888 5504 3928 5536
rect 3960 5504 4000 5536
rect 0 5464 4000 5504
rect 0 5432 40 5464
rect 72 5432 112 5464
rect 144 5432 184 5464
rect 216 5432 256 5464
rect 288 5432 328 5464
rect 360 5432 400 5464
rect 432 5432 472 5464
rect 504 5432 544 5464
rect 576 5432 616 5464
rect 648 5432 688 5464
rect 720 5432 760 5464
rect 792 5432 832 5464
rect 864 5432 904 5464
rect 936 5432 976 5464
rect 1008 5432 1048 5464
rect 1080 5432 1120 5464
rect 1152 5432 1192 5464
rect 1224 5432 1264 5464
rect 1296 5432 1336 5464
rect 1368 5432 1408 5464
rect 1440 5432 1480 5464
rect 1512 5432 1552 5464
rect 1584 5432 1624 5464
rect 1656 5432 1696 5464
rect 1728 5432 1768 5464
rect 1800 5432 1840 5464
rect 1872 5432 1912 5464
rect 1944 5432 1984 5464
rect 2016 5432 2056 5464
rect 2088 5432 2128 5464
rect 2160 5432 2200 5464
rect 2232 5432 2272 5464
rect 2304 5432 2344 5464
rect 2376 5432 2416 5464
rect 2448 5432 2488 5464
rect 2520 5432 2560 5464
rect 2592 5432 2632 5464
rect 2664 5432 2704 5464
rect 2736 5432 2776 5464
rect 2808 5432 2848 5464
rect 2880 5432 2920 5464
rect 2952 5432 2992 5464
rect 3024 5432 3064 5464
rect 3096 5432 3136 5464
rect 3168 5432 3208 5464
rect 3240 5432 3280 5464
rect 3312 5432 3352 5464
rect 3384 5432 3424 5464
rect 3456 5432 3496 5464
rect 3528 5432 3568 5464
rect 3600 5432 3640 5464
rect 3672 5432 3712 5464
rect 3744 5432 3784 5464
rect 3816 5432 3856 5464
rect 3888 5432 3928 5464
rect 3960 5432 4000 5464
rect 0 5392 4000 5432
rect 0 5360 40 5392
rect 72 5360 112 5392
rect 144 5360 184 5392
rect 216 5360 256 5392
rect 288 5360 328 5392
rect 360 5360 400 5392
rect 432 5360 472 5392
rect 504 5360 544 5392
rect 576 5360 616 5392
rect 648 5360 688 5392
rect 720 5360 760 5392
rect 792 5360 832 5392
rect 864 5360 904 5392
rect 936 5360 976 5392
rect 1008 5360 1048 5392
rect 1080 5360 1120 5392
rect 1152 5360 1192 5392
rect 1224 5360 1264 5392
rect 1296 5360 1336 5392
rect 1368 5360 1408 5392
rect 1440 5360 1480 5392
rect 1512 5360 1552 5392
rect 1584 5360 1624 5392
rect 1656 5360 1696 5392
rect 1728 5360 1768 5392
rect 1800 5360 1840 5392
rect 1872 5360 1912 5392
rect 1944 5360 1984 5392
rect 2016 5360 2056 5392
rect 2088 5360 2128 5392
rect 2160 5360 2200 5392
rect 2232 5360 2272 5392
rect 2304 5360 2344 5392
rect 2376 5360 2416 5392
rect 2448 5360 2488 5392
rect 2520 5360 2560 5392
rect 2592 5360 2632 5392
rect 2664 5360 2704 5392
rect 2736 5360 2776 5392
rect 2808 5360 2848 5392
rect 2880 5360 2920 5392
rect 2952 5360 2992 5392
rect 3024 5360 3064 5392
rect 3096 5360 3136 5392
rect 3168 5360 3208 5392
rect 3240 5360 3280 5392
rect 3312 5360 3352 5392
rect 3384 5360 3424 5392
rect 3456 5360 3496 5392
rect 3528 5360 3568 5392
rect 3600 5360 3640 5392
rect 3672 5360 3712 5392
rect 3744 5360 3784 5392
rect 3816 5360 3856 5392
rect 3888 5360 3928 5392
rect 3960 5360 4000 5392
rect 0 5320 4000 5360
rect 0 5288 40 5320
rect 72 5288 112 5320
rect 144 5288 184 5320
rect 216 5288 256 5320
rect 288 5288 328 5320
rect 360 5288 400 5320
rect 432 5288 472 5320
rect 504 5288 544 5320
rect 576 5288 616 5320
rect 648 5288 688 5320
rect 720 5288 760 5320
rect 792 5288 832 5320
rect 864 5288 904 5320
rect 936 5288 976 5320
rect 1008 5288 1048 5320
rect 1080 5288 1120 5320
rect 1152 5288 1192 5320
rect 1224 5288 1264 5320
rect 1296 5288 1336 5320
rect 1368 5288 1408 5320
rect 1440 5288 1480 5320
rect 1512 5288 1552 5320
rect 1584 5288 1624 5320
rect 1656 5288 1696 5320
rect 1728 5288 1768 5320
rect 1800 5288 1840 5320
rect 1872 5288 1912 5320
rect 1944 5288 1984 5320
rect 2016 5288 2056 5320
rect 2088 5288 2128 5320
rect 2160 5288 2200 5320
rect 2232 5288 2272 5320
rect 2304 5288 2344 5320
rect 2376 5288 2416 5320
rect 2448 5288 2488 5320
rect 2520 5288 2560 5320
rect 2592 5288 2632 5320
rect 2664 5288 2704 5320
rect 2736 5288 2776 5320
rect 2808 5288 2848 5320
rect 2880 5288 2920 5320
rect 2952 5288 2992 5320
rect 3024 5288 3064 5320
rect 3096 5288 3136 5320
rect 3168 5288 3208 5320
rect 3240 5288 3280 5320
rect 3312 5288 3352 5320
rect 3384 5288 3424 5320
rect 3456 5288 3496 5320
rect 3528 5288 3568 5320
rect 3600 5288 3640 5320
rect 3672 5288 3712 5320
rect 3744 5288 3784 5320
rect 3816 5288 3856 5320
rect 3888 5288 3928 5320
rect 3960 5288 4000 5320
rect 0 5248 4000 5288
rect 0 5216 40 5248
rect 72 5216 112 5248
rect 144 5216 184 5248
rect 216 5216 256 5248
rect 288 5216 328 5248
rect 360 5216 400 5248
rect 432 5216 472 5248
rect 504 5216 544 5248
rect 576 5216 616 5248
rect 648 5216 688 5248
rect 720 5216 760 5248
rect 792 5216 832 5248
rect 864 5216 904 5248
rect 936 5216 976 5248
rect 1008 5216 1048 5248
rect 1080 5216 1120 5248
rect 1152 5216 1192 5248
rect 1224 5216 1264 5248
rect 1296 5216 1336 5248
rect 1368 5216 1408 5248
rect 1440 5216 1480 5248
rect 1512 5216 1552 5248
rect 1584 5216 1624 5248
rect 1656 5216 1696 5248
rect 1728 5216 1768 5248
rect 1800 5216 1840 5248
rect 1872 5216 1912 5248
rect 1944 5216 1984 5248
rect 2016 5216 2056 5248
rect 2088 5216 2128 5248
rect 2160 5216 2200 5248
rect 2232 5216 2272 5248
rect 2304 5216 2344 5248
rect 2376 5216 2416 5248
rect 2448 5216 2488 5248
rect 2520 5216 2560 5248
rect 2592 5216 2632 5248
rect 2664 5216 2704 5248
rect 2736 5216 2776 5248
rect 2808 5216 2848 5248
rect 2880 5216 2920 5248
rect 2952 5216 2992 5248
rect 3024 5216 3064 5248
rect 3096 5216 3136 5248
rect 3168 5216 3208 5248
rect 3240 5216 3280 5248
rect 3312 5216 3352 5248
rect 3384 5216 3424 5248
rect 3456 5216 3496 5248
rect 3528 5216 3568 5248
rect 3600 5216 3640 5248
rect 3672 5216 3712 5248
rect 3744 5216 3784 5248
rect 3816 5216 3856 5248
rect 3888 5216 3928 5248
rect 3960 5216 4000 5248
rect 0 5176 4000 5216
rect 0 5144 40 5176
rect 72 5144 112 5176
rect 144 5144 184 5176
rect 216 5144 256 5176
rect 288 5144 328 5176
rect 360 5144 400 5176
rect 432 5144 472 5176
rect 504 5144 544 5176
rect 576 5144 616 5176
rect 648 5144 688 5176
rect 720 5144 760 5176
rect 792 5144 832 5176
rect 864 5144 904 5176
rect 936 5144 976 5176
rect 1008 5144 1048 5176
rect 1080 5144 1120 5176
rect 1152 5144 1192 5176
rect 1224 5144 1264 5176
rect 1296 5144 1336 5176
rect 1368 5144 1408 5176
rect 1440 5144 1480 5176
rect 1512 5144 1552 5176
rect 1584 5144 1624 5176
rect 1656 5144 1696 5176
rect 1728 5144 1768 5176
rect 1800 5144 1840 5176
rect 1872 5144 1912 5176
rect 1944 5144 1984 5176
rect 2016 5144 2056 5176
rect 2088 5144 2128 5176
rect 2160 5144 2200 5176
rect 2232 5144 2272 5176
rect 2304 5144 2344 5176
rect 2376 5144 2416 5176
rect 2448 5144 2488 5176
rect 2520 5144 2560 5176
rect 2592 5144 2632 5176
rect 2664 5144 2704 5176
rect 2736 5144 2776 5176
rect 2808 5144 2848 5176
rect 2880 5144 2920 5176
rect 2952 5144 2992 5176
rect 3024 5144 3064 5176
rect 3096 5144 3136 5176
rect 3168 5144 3208 5176
rect 3240 5144 3280 5176
rect 3312 5144 3352 5176
rect 3384 5144 3424 5176
rect 3456 5144 3496 5176
rect 3528 5144 3568 5176
rect 3600 5144 3640 5176
rect 3672 5144 3712 5176
rect 3744 5144 3784 5176
rect 3816 5144 3856 5176
rect 3888 5144 3928 5176
rect 3960 5144 4000 5176
rect 0 5104 4000 5144
rect 0 5072 40 5104
rect 72 5072 112 5104
rect 144 5072 184 5104
rect 216 5072 256 5104
rect 288 5072 328 5104
rect 360 5072 400 5104
rect 432 5072 472 5104
rect 504 5072 544 5104
rect 576 5072 616 5104
rect 648 5072 688 5104
rect 720 5072 760 5104
rect 792 5072 832 5104
rect 864 5072 904 5104
rect 936 5072 976 5104
rect 1008 5072 1048 5104
rect 1080 5072 1120 5104
rect 1152 5072 1192 5104
rect 1224 5072 1264 5104
rect 1296 5072 1336 5104
rect 1368 5072 1408 5104
rect 1440 5072 1480 5104
rect 1512 5072 1552 5104
rect 1584 5072 1624 5104
rect 1656 5072 1696 5104
rect 1728 5072 1768 5104
rect 1800 5072 1840 5104
rect 1872 5072 1912 5104
rect 1944 5072 1984 5104
rect 2016 5072 2056 5104
rect 2088 5072 2128 5104
rect 2160 5072 2200 5104
rect 2232 5072 2272 5104
rect 2304 5072 2344 5104
rect 2376 5072 2416 5104
rect 2448 5072 2488 5104
rect 2520 5072 2560 5104
rect 2592 5072 2632 5104
rect 2664 5072 2704 5104
rect 2736 5072 2776 5104
rect 2808 5072 2848 5104
rect 2880 5072 2920 5104
rect 2952 5072 2992 5104
rect 3024 5072 3064 5104
rect 3096 5072 3136 5104
rect 3168 5072 3208 5104
rect 3240 5072 3280 5104
rect 3312 5072 3352 5104
rect 3384 5072 3424 5104
rect 3456 5072 3496 5104
rect 3528 5072 3568 5104
rect 3600 5072 3640 5104
rect 3672 5072 3712 5104
rect 3744 5072 3784 5104
rect 3816 5072 3856 5104
rect 3888 5072 3928 5104
rect 3960 5072 4000 5104
rect 0 5032 4000 5072
rect 0 5000 40 5032
rect 72 5000 112 5032
rect 144 5000 184 5032
rect 216 5000 256 5032
rect 288 5000 328 5032
rect 360 5000 400 5032
rect 432 5000 472 5032
rect 504 5000 544 5032
rect 576 5000 616 5032
rect 648 5000 688 5032
rect 720 5000 760 5032
rect 792 5000 832 5032
rect 864 5000 904 5032
rect 936 5000 976 5032
rect 1008 5000 1048 5032
rect 1080 5000 1120 5032
rect 1152 5000 1192 5032
rect 1224 5000 1264 5032
rect 1296 5000 1336 5032
rect 1368 5000 1408 5032
rect 1440 5000 1480 5032
rect 1512 5000 1552 5032
rect 1584 5000 1624 5032
rect 1656 5000 1696 5032
rect 1728 5000 1768 5032
rect 1800 5000 1840 5032
rect 1872 5000 1912 5032
rect 1944 5000 1984 5032
rect 2016 5000 2056 5032
rect 2088 5000 2128 5032
rect 2160 5000 2200 5032
rect 2232 5000 2272 5032
rect 2304 5000 2344 5032
rect 2376 5000 2416 5032
rect 2448 5000 2488 5032
rect 2520 5000 2560 5032
rect 2592 5000 2632 5032
rect 2664 5000 2704 5032
rect 2736 5000 2776 5032
rect 2808 5000 2848 5032
rect 2880 5000 2920 5032
rect 2952 5000 2992 5032
rect 3024 5000 3064 5032
rect 3096 5000 3136 5032
rect 3168 5000 3208 5032
rect 3240 5000 3280 5032
rect 3312 5000 3352 5032
rect 3384 5000 3424 5032
rect 3456 5000 3496 5032
rect 3528 5000 3568 5032
rect 3600 5000 3640 5032
rect 3672 5000 3712 5032
rect 3744 5000 3784 5032
rect 3816 5000 3856 5032
rect 3888 5000 3928 5032
rect 3960 5000 4000 5032
rect 0 4960 4000 5000
rect 0 4928 40 4960
rect 72 4928 112 4960
rect 144 4928 184 4960
rect 216 4928 256 4960
rect 288 4928 328 4960
rect 360 4928 400 4960
rect 432 4928 472 4960
rect 504 4928 544 4960
rect 576 4928 616 4960
rect 648 4928 688 4960
rect 720 4928 760 4960
rect 792 4928 832 4960
rect 864 4928 904 4960
rect 936 4928 976 4960
rect 1008 4928 1048 4960
rect 1080 4928 1120 4960
rect 1152 4928 1192 4960
rect 1224 4928 1264 4960
rect 1296 4928 1336 4960
rect 1368 4928 1408 4960
rect 1440 4928 1480 4960
rect 1512 4928 1552 4960
rect 1584 4928 1624 4960
rect 1656 4928 1696 4960
rect 1728 4928 1768 4960
rect 1800 4928 1840 4960
rect 1872 4928 1912 4960
rect 1944 4928 1984 4960
rect 2016 4928 2056 4960
rect 2088 4928 2128 4960
rect 2160 4928 2200 4960
rect 2232 4928 2272 4960
rect 2304 4928 2344 4960
rect 2376 4928 2416 4960
rect 2448 4928 2488 4960
rect 2520 4928 2560 4960
rect 2592 4928 2632 4960
rect 2664 4928 2704 4960
rect 2736 4928 2776 4960
rect 2808 4928 2848 4960
rect 2880 4928 2920 4960
rect 2952 4928 2992 4960
rect 3024 4928 3064 4960
rect 3096 4928 3136 4960
rect 3168 4928 3208 4960
rect 3240 4928 3280 4960
rect 3312 4928 3352 4960
rect 3384 4928 3424 4960
rect 3456 4928 3496 4960
rect 3528 4928 3568 4960
rect 3600 4928 3640 4960
rect 3672 4928 3712 4960
rect 3744 4928 3784 4960
rect 3816 4928 3856 4960
rect 3888 4928 3928 4960
rect 3960 4928 4000 4960
rect 0 4888 4000 4928
rect 0 4856 40 4888
rect 72 4856 112 4888
rect 144 4856 184 4888
rect 216 4856 256 4888
rect 288 4856 328 4888
rect 360 4856 400 4888
rect 432 4856 472 4888
rect 504 4856 544 4888
rect 576 4856 616 4888
rect 648 4856 688 4888
rect 720 4856 760 4888
rect 792 4856 832 4888
rect 864 4856 904 4888
rect 936 4856 976 4888
rect 1008 4856 1048 4888
rect 1080 4856 1120 4888
rect 1152 4856 1192 4888
rect 1224 4856 1264 4888
rect 1296 4856 1336 4888
rect 1368 4856 1408 4888
rect 1440 4856 1480 4888
rect 1512 4856 1552 4888
rect 1584 4856 1624 4888
rect 1656 4856 1696 4888
rect 1728 4856 1768 4888
rect 1800 4856 1840 4888
rect 1872 4856 1912 4888
rect 1944 4856 1984 4888
rect 2016 4856 2056 4888
rect 2088 4856 2128 4888
rect 2160 4856 2200 4888
rect 2232 4856 2272 4888
rect 2304 4856 2344 4888
rect 2376 4856 2416 4888
rect 2448 4856 2488 4888
rect 2520 4856 2560 4888
rect 2592 4856 2632 4888
rect 2664 4856 2704 4888
rect 2736 4856 2776 4888
rect 2808 4856 2848 4888
rect 2880 4856 2920 4888
rect 2952 4856 2992 4888
rect 3024 4856 3064 4888
rect 3096 4856 3136 4888
rect 3168 4856 3208 4888
rect 3240 4856 3280 4888
rect 3312 4856 3352 4888
rect 3384 4856 3424 4888
rect 3456 4856 3496 4888
rect 3528 4856 3568 4888
rect 3600 4856 3640 4888
rect 3672 4856 3712 4888
rect 3744 4856 3784 4888
rect 3816 4856 3856 4888
rect 3888 4856 3928 4888
rect 3960 4856 4000 4888
rect 0 4816 4000 4856
rect 0 4784 40 4816
rect 72 4784 112 4816
rect 144 4784 184 4816
rect 216 4784 256 4816
rect 288 4784 328 4816
rect 360 4784 400 4816
rect 432 4784 472 4816
rect 504 4784 544 4816
rect 576 4784 616 4816
rect 648 4784 688 4816
rect 720 4784 760 4816
rect 792 4784 832 4816
rect 864 4784 904 4816
rect 936 4784 976 4816
rect 1008 4784 1048 4816
rect 1080 4784 1120 4816
rect 1152 4784 1192 4816
rect 1224 4784 1264 4816
rect 1296 4784 1336 4816
rect 1368 4784 1408 4816
rect 1440 4784 1480 4816
rect 1512 4784 1552 4816
rect 1584 4784 1624 4816
rect 1656 4784 1696 4816
rect 1728 4784 1768 4816
rect 1800 4784 1840 4816
rect 1872 4784 1912 4816
rect 1944 4784 1984 4816
rect 2016 4784 2056 4816
rect 2088 4784 2128 4816
rect 2160 4784 2200 4816
rect 2232 4784 2272 4816
rect 2304 4784 2344 4816
rect 2376 4784 2416 4816
rect 2448 4784 2488 4816
rect 2520 4784 2560 4816
rect 2592 4784 2632 4816
rect 2664 4784 2704 4816
rect 2736 4784 2776 4816
rect 2808 4784 2848 4816
rect 2880 4784 2920 4816
rect 2952 4784 2992 4816
rect 3024 4784 3064 4816
rect 3096 4784 3136 4816
rect 3168 4784 3208 4816
rect 3240 4784 3280 4816
rect 3312 4784 3352 4816
rect 3384 4784 3424 4816
rect 3456 4784 3496 4816
rect 3528 4784 3568 4816
rect 3600 4784 3640 4816
rect 3672 4784 3712 4816
rect 3744 4784 3784 4816
rect 3816 4784 3856 4816
rect 3888 4784 3928 4816
rect 3960 4784 4000 4816
rect 0 4744 4000 4784
rect 0 4712 40 4744
rect 72 4712 112 4744
rect 144 4712 184 4744
rect 216 4712 256 4744
rect 288 4712 328 4744
rect 360 4712 400 4744
rect 432 4712 472 4744
rect 504 4712 544 4744
rect 576 4712 616 4744
rect 648 4712 688 4744
rect 720 4712 760 4744
rect 792 4712 832 4744
rect 864 4712 904 4744
rect 936 4712 976 4744
rect 1008 4712 1048 4744
rect 1080 4712 1120 4744
rect 1152 4712 1192 4744
rect 1224 4712 1264 4744
rect 1296 4712 1336 4744
rect 1368 4712 1408 4744
rect 1440 4712 1480 4744
rect 1512 4712 1552 4744
rect 1584 4712 1624 4744
rect 1656 4712 1696 4744
rect 1728 4712 1768 4744
rect 1800 4712 1840 4744
rect 1872 4712 1912 4744
rect 1944 4712 1984 4744
rect 2016 4712 2056 4744
rect 2088 4712 2128 4744
rect 2160 4712 2200 4744
rect 2232 4712 2272 4744
rect 2304 4712 2344 4744
rect 2376 4712 2416 4744
rect 2448 4712 2488 4744
rect 2520 4712 2560 4744
rect 2592 4712 2632 4744
rect 2664 4712 2704 4744
rect 2736 4712 2776 4744
rect 2808 4712 2848 4744
rect 2880 4712 2920 4744
rect 2952 4712 2992 4744
rect 3024 4712 3064 4744
rect 3096 4712 3136 4744
rect 3168 4712 3208 4744
rect 3240 4712 3280 4744
rect 3312 4712 3352 4744
rect 3384 4712 3424 4744
rect 3456 4712 3496 4744
rect 3528 4712 3568 4744
rect 3600 4712 3640 4744
rect 3672 4712 3712 4744
rect 3744 4712 3784 4744
rect 3816 4712 3856 4744
rect 3888 4712 3928 4744
rect 3960 4712 4000 4744
rect 0 4672 4000 4712
rect 0 4640 40 4672
rect 72 4640 112 4672
rect 144 4640 184 4672
rect 216 4640 256 4672
rect 288 4640 328 4672
rect 360 4640 400 4672
rect 432 4640 472 4672
rect 504 4640 544 4672
rect 576 4640 616 4672
rect 648 4640 688 4672
rect 720 4640 760 4672
rect 792 4640 832 4672
rect 864 4640 904 4672
rect 936 4640 976 4672
rect 1008 4640 1048 4672
rect 1080 4640 1120 4672
rect 1152 4640 1192 4672
rect 1224 4640 1264 4672
rect 1296 4640 1336 4672
rect 1368 4640 1408 4672
rect 1440 4640 1480 4672
rect 1512 4640 1552 4672
rect 1584 4640 1624 4672
rect 1656 4640 1696 4672
rect 1728 4640 1768 4672
rect 1800 4640 1840 4672
rect 1872 4640 1912 4672
rect 1944 4640 1984 4672
rect 2016 4640 2056 4672
rect 2088 4640 2128 4672
rect 2160 4640 2200 4672
rect 2232 4640 2272 4672
rect 2304 4640 2344 4672
rect 2376 4640 2416 4672
rect 2448 4640 2488 4672
rect 2520 4640 2560 4672
rect 2592 4640 2632 4672
rect 2664 4640 2704 4672
rect 2736 4640 2776 4672
rect 2808 4640 2848 4672
rect 2880 4640 2920 4672
rect 2952 4640 2992 4672
rect 3024 4640 3064 4672
rect 3096 4640 3136 4672
rect 3168 4640 3208 4672
rect 3240 4640 3280 4672
rect 3312 4640 3352 4672
rect 3384 4640 3424 4672
rect 3456 4640 3496 4672
rect 3528 4640 3568 4672
rect 3600 4640 3640 4672
rect 3672 4640 3712 4672
rect 3744 4640 3784 4672
rect 3816 4640 3856 4672
rect 3888 4640 3928 4672
rect 3960 4640 4000 4672
rect 0 4600 4000 4640
rect 0 4568 40 4600
rect 72 4568 112 4600
rect 144 4568 184 4600
rect 216 4568 256 4600
rect 288 4568 328 4600
rect 360 4568 400 4600
rect 432 4568 472 4600
rect 504 4568 544 4600
rect 576 4568 616 4600
rect 648 4568 688 4600
rect 720 4568 760 4600
rect 792 4568 832 4600
rect 864 4568 904 4600
rect 936 4568 976 4600
rect 1008 4568 1048 4600
rect 1080 4568 1120 4600
rect 1152 4568 1192 4600
rect 1224 4568 1264 4600
rect 1296 4568 1336 4600
rect 1368 4568 1408 4600
rect 1440 4568 1480 4600
rect 1512 4568 1552 4600
rect 1584 4568 1624 4600
rect 1656 4568 1696 4600
rect 1728 4568 1768 4600
rect 1800 4568 1840 4600
rect 1872 4568 1912 4600
rect 1944 4568 1984 4600
rect 2016 4568 2056 4600
rect 2088 4568 2128 4600
rect 2160 4568 2200 4600
rect 2232 4568 2272 4600
rect 2304 4568 2344 4600
rect 2376 4568 2416 4600
rect 2448 4568 2488 4600
rect 2520 4568 2560 4600
rect 2592 4568 2632 4600
rect 2664 4568 2704 4600
rect 2736 4568 2776 4600
rect 2808 4568 2848 4600
rect 2880 4568 2920 4600
rect 2952 4568 2992 4600
rect 3024 4568 3064 4600
rect 3096 4568 3136 4600
rect 3168 4568 3208 4600
rect 3240 4568 3280 4600
rect 3312 4568 3352 4600
rect 3384 4568 3424 4600
rect 3456 4568 3496 4600
rect 3528 4568 3568 4600
rect 3600 4568 3640 4600
rect 3672 4568 3712 4600
rect 3744 4568 3784 4600
rect 3816 4568 3856 4600
rect 3888 4568 3928 4600
rect 3960 4568 4000 4600
rect 0 4528 4000 4568
rect 0 4496 40 4528
rect 72 4496 112 4528
rect 144 4496 184 4528
rect 216 4496 256 4528
rect 288 4496 328 4528
rect 360 4496 400 4528
rect 432 4496 472 4528
rect 504 4496 544 4528
rect 576 4496 616 4528
rect 648 4496 688 4528
rect 720 4496 760 4528
rect 792 4496 832 4528
rect 864 4496 904 4528
rect 936 4496 976 4528
rect 1008 4496 1048 4528
rect 1080 4496 1120 4528
rect 1152 4496 1192 4528
rect 1224 4496 1264 4528
rect 1296 4496 1336 4528
rect 1368 4496 1408 4528
rect 1440 4496 1480 4528
rect 1512 4496 1552 4528
rect 1584 4496 1624 4528
rect 1656 4496 1696 4528
rect 1728 4496 1768 4528
rect 1800 4496 1840 4528
rect 1872 4496 1912 4528
rect 1944 4496 1984 4528
rect 2016 4496 2056 4528
rect 2088 4496 2128 4528
rect 2160 4496 2200 4528
rect 2232 4496 2272 4528
rect 2304 4496 2344 4528
rect 2376 4496 2416 4528
rect 2448 4496 2488 4528
rect 2520 4496 2560 4528
rect 2592 4496 2632 4528
rect 2664 4496 2704 4528
rect 2736 4496 2776 4528
rect 2808 4496 2848 4528
rect 2880 4496 2920 4528
rect 2952 4496 2992 4528
rect 3024 4496 3064 4528
rect 3096 4496 3136 4528
rect 3168 4496 3208 4528
rect 3240 4496 3280 4528
rect 3312 4496 3352 4528
rect 3384 4496 3424 4528
rect 3456 4496 3496 4528
rect 3528 4496 3568 4528
rect 3600 4496 3640 4528
rect 3672 4496 3712 4528
rect 3744 4496 3784 4528
rect 3816 4496 3856 4528
rect 3888 4496 3928 4528
rect 3960 4496 4000 4528
rect 0 4456 4000 4496
rect 0 4424 40 4456
rect 72 4424 112 4456
rect 144 4424 184 4456
rect 216 4424 256 4456
rect 288 4424 328 4456
rect 360 4424 400 4456
rect 432 4424 472 4456
rect 504 4424 544 4456
rect 576 4424 616 4456
rect 648 4424 688 4456
rect 720 4424 760 4456
rect 792 4424 832 4456
rect 864 4424 904 4456
rect 936 4424 976 4456
rect 1008 4424 1048 4456
rect 1080 4424 1120 4456
rect 1152 4424 1192 4456
rect 1224 4424 1264 4456
rect 1296 4424 1336 4456
rect 1368 4424 1408 4456
rect 1440 4424 1480 4456
rect 1512 4424 1552 4456
rect 1584 4424 1624 4456
rect 1656 4424 1696 4456
rect 1728 4424 1768 4456
rect 1800 4424 1840 4456
rect 1872 4424 1912 4456
rect 1944 4424 1984 4456
rect 2016 4424 2056 4456
rect 2088 4424 2128 4456
rect 2160 4424 2200 4456
rect 2232 4424 2272 4456
rect 2304 4424 2344 4456
rect 2376 4424 2416 4456
rect 2448 4424 2488 4456
rect 2520 4424 2560 4456
rect 2592 4424 2632 4456
rect 2664 4424 2704 4456
rect 2736 4424 2776 4456
rect 2808 4424 2848 4456
rect 2880 4424 2920 4456
rect 2952 4424 2992 4456
rect 3024 4424 3064 4456
rect 3096 4424 3136 4456
rect 3168 4424 3208 4456
rect 3240 4424 3280 4456
rect 3312 4424 3352 4456
rect 3384 4424 3424 4456
rect 3456 4424 3496 4456
rect 3528 4424 3568 4456
rect 3600 4424 3640 4456
rect 3672 4424 3712 4456
rect 3744 4424 3784 4456
rect 3816 4424 3856 4456
rect 3888 4424 3928 4456
rect 3960 4424 4000 4456
rect 0 4384 4000 4424
rect 0 4352 40 4384
rect 72 4352 112 4384
rect 144 4352 184 4384
rect 216 4352 256 4384
rect 288 4352 328 4384
rect 360 4352 400 4384
rect 432 4352 472 4384
rect 504 4352 544 4384
rect 576 4352 616 4384
rect 648 4352 688 4384
rect 720 4352 760 4384
rect 792 4352 832 4384
rect 864 4352 904 4384
rect 936 4352 976 4384
rect 1008 4352 1048 4384
rect 1080 4352 1120 4384
rect 1152 4352 1192 4384
rect 1224 4352 1264 4384
rect 1296 4352 1336 4384
rect 1368 4352 1408 4384
rect 1440 4352 1480 4384
rect 1512 4352 1552 4384
rect 1584 4352 1624 4384
rect 1656 4352 1696 4384
rect 1728 4352 1768 4384
rect 1800 4352 1840 4384
rect 1872 4352 1912 4384
rect 1944 4352 1984 4384
rect 2016 4352 2056 4384
rect 2088 4352 2128 4384
rect 2160 4352 2200 4384
rect 2232 4352 2272 4384
rect 2304 4352 2344 4384
rect 2376 4352 2416 4384
rect 2448 4352 2488 4384
rect 2520 4352 2560 4384
rect 2592 4352 2632 4384
rect 2664 4352 2704 4384
rect 2736 4352 2776 4384
rect 2808 4352 2848 4384
rect 2880 4352 2920 4384
rect 2952 4352 2992 4384
rect 3024 4352 3064 4384
rect 3096 4352 3136 4384
rect 3168 4352 3208 4384
rect 3240 4352 3280 4384
rect 3312 4352 3352 4384
rect 3384 4352 3424 4384
rect 3456 4352 3496 4384
rect 3528 4352 3568 4384
rect 3600 4352 3640 4384
rect 3672 4352 3712 4384
rect 3744 4352 3784 4384
rect 3816 4352 3856 4384
rect 3888 4352 3928 4384
rect 3960 4352 4000 4384
rect 0 4312 4000 4352
rect 0 4280 40 4312
rect 72 4280 112 4312
rect 144 4280 184 4312
rect 216 4280 256 4312
rect 288 4280 328 4312
rect 360 4280 400 4312
rect 432 4280 472 4312
rect 504 4280 544 4312
rect 576 4280 616 4312
rect 648 4280 688 4312
rect 720 4280 760 4312
rect 792 4280 832 4312
rect 864 4280 904 4312
rect 936 4280 976 4312
rect 1008 4280 1048 4312
rect 1080 4280 1120 4312
rect 1152 4280 1192 4312
rect 1224 4280 1264 4312
rect 1296 4280 1336 4312
rect 1368 4280 1408 4312
rect 1440 4280 1480 4312
rect 1512 4280 1552 4312
rect 1584 4280 1624 4312
rect 1656 4280 1696 4312
rect 1728 4280 1768 4312
rect 1800 4280 1840 4312
rect 1872 4280 1912 4312
rect 1944 4280 1984 4312
rect 2016 4280 2056 4312
rect 2088 4280 2128 4312
rect 2160 4280 2200 4312
rect 2232 4280 2272 4312
rect 2304 4280 2344 4312
rect 2376 4280 2416 4312
rect 2448 4280 2488 4312
rect 2520 4280 2560 4312
rect 2592 4280 2632 4312
rect 2664 4280 2704 4312
rect 2736 4280 2776 4312
rect 2808 4280 2848 4312
rect 2880 4280 2920 4312
rect 2952 4280 2992 4312
rect 3024 4280 3064 4312
rect 3096 4280 3136 4312
rect 3168 4280 3208 4312
rect 3240 4280 3280 4312
rect 3312 4280 3352 4312
rect 3384 4280 3424 4312
rect 3456 4280 3496 4312
rect 3528 4280 3568 4312
rect 3600 4280 3640 4312
rect 3672 4280 3712 4312
rect 3744 4280 3784 4312
rect 3816 4280 3856 4312
rect 3888 4280 3928 4312
rect 3960 4280 4000 4312
rect 0 4240 4000 4280
rect 0 4208 40 4240
rect 72 4208 112 4240
rect 144 4208 184 4240
rect 216 4208 256 4240
rect 288 4208 328 4240
rect 360 4208 400 4240
rect 432 4208 472 4240
rect 504 4208 544 4240
rect 576 4208 616 4240
rect 648 4208 688 4240
rect 720 4208 760 4240
rect 792 4208 832 4240
rect 864 4208 904 4240
rect 936 4208 976 4240
rect 1008 4208 1048 4240
rect 1080 4208 1120 4240
rect 1152 4208 1192 4240
rect 1224 4208 1264 4240
rect 1296 4208 1336 4240
rect 1368 4208 1408 4240
rect 1440 4208 1480 4240
rect 1512 4208 1552 4240
rect 1584 4208 1624 4240
rect 1656 4208 1696 4240
rect 1728 4208 1768 4240
rect 1800 4208 1840 4240
rect 1872 4208 1912 4240
rect 1944 4208 1984 4240
rect 2016 4208 2056 4240
rect 2088 4208 2128 4240
rect 2160 4208 2200 4240
rect 2232 4208 2272 4240
rect 2304 4208 2344 4240
rect 2376 4208 2416 4240
rect 2448 4208 2488 4240
rect 2520 4208 2560 4240
rect 2592 4208 2632 4240
rect 2664 4208 2704 4240
rect 2736 4208 2776 4240
rect 2808 4208 2848 4240
rect 2880 4208 2920 4240
rect 2952 4208 2992 4240
rect 3024 4208 3064 4240
rect 3096 4208 3136 4240
rect 3168 4208 3208 4240
rect 3240 4208 3280 4240
rect 3312 4208 3352 4240
rect 3384 4208 3424 4240
rect 3456 4208 3496 4240
rect 3528 4208 3568 4240
rect 3600 4208 3640 4240
rect 3672 4208 3712 4240
rect 3744 4208 3784 4240
rect 3816 4208 3856 4240
rect 3888 4208 3928 4240
rect 3960 4208 4000 4240
rect 0 4168 4000 4208
rect 0 4136 40 4168
rect 72 4136 112 4168
rect 144 4136 184 4168
rect 216 4136 256 4168
rect 288 4136 328 4168
rect 360 4136 400 4168
rect 432 4136 472 4168
rect 504 4136 544 4168
rect 576 4136 616 4168
rect 648 4136 688 4168
rect 720 4136 760 4168
rect 792 4136 832 4168
rect 864 4136 904 4168
rect 936 4136 976 4168
rect 1008 4136 1048 4168
rect 1080 4136 1120 4168
rect 1152 4136 1192 4168
rect 1224 4136 1264 4168
rect 1296 4136 1336 4168
rect 1368 4136 1408 4168
rect 1440 4136 1480 4168
rect 1512 4136 1552 4168
rect 1584 4136 1624 4168
rect 1656 4136 1696 4168
rect 1728 4136 1768 4168
rect 1800 4136 1840 4168
rect 1872 4136 1912 4168
rect 1944 4136 1984 4168
rect 2016 4136 2056 4168
rect 2088 4136 2128 4168
rect 2160 4136 2200 4168
rect 2232 4136 2272 4168
rect 2304 4136 2344 4168
rect 2376 4136 2416 4168
rect 2448 4136 2488 4168
rect 2520 4136 2560 4168
rect 2592 4136 2632 4168
rect 2664 4136 2704 4168
rect 2736 4136 2776 4168
rect 2808 4136 2848 4168
rect 2880 4136 2920 4168
rect 2952 4136 2992 4168
rect 3024 4136 3064 4168
rect 3096 4136 3136 4168
rect 3168 4136 3208 4168
rect 3240 4136 3280 4168
rect 3312 4136 3352 4168
rect 3384 4136 3424 4168
rect 3456 4136 3496 4168
rect 3528 4136 3568 4168
rect 3600 4136 3640 4168
rect 3672 4136 3712 4168
rect 3744 4136 3784 4168
rect 3816 4136 3856 4168
rect 3888 4136 3928 4168
rect 3960 4136 4000 4168
rect 0 4096 4000 4136
rect 0 4064 40 4096
rect 72 4064 112 4096
rect 144 4064 184 4096
rect 216 4064 256 4096
rect 288 4064 328 4096
rect 360 4064 400 4096
rect 432 4064 472 4096
rect 504 4064 544 4096
rect 576 4064 616 4096
rect 648 4064 688 4096
rect 720 4064 760 4096
rect 792 4064 832 4096
rect 864 4064 904 4096
rect 936 4064 976 4096
rect 1008 4064 1048 4096
rect 1080 4064 1120 4096
rect 1152 4064 1192 4096
rect 1224 4064 1264 4096
rect 1296 4064 1336 4096
rect 1368 4064 1408 4096
rect 1440 4064 1480 4096
rect 1512 4064 1552 4096
rect 1584 4064 1624 4096
rect 1656 4064 1696 4096
rect 1728 4064 1768 4096
rect 1800 4064 1840 4096
rect 1872 4064 1912 4096
rect 1944 4064 1984 4096
rect 2016 4064 2056 4096
rect 2088 4064 2128 4096
rect 2160 4064 2200 4096
rect 2232 4064 2272 4096
rect 2304 4064 2344 4096
rect 2376 4064 2416 4096
rect 2448 4064 2488 4096
rect 2520 4064 2560 4096
rect 2592 4064 2632 4096
rect 2664 4064 2704 4096
rect 2736 4064 2776 4096
rect 2808 4064 2848 4096
rect 2880 4064 2920 4096
rect 2952 4064 2992 4096
rect 3024 4064 3064 4096
rect 3096 4064 3136 4096
rect 3168 4064 3208 4096
rect 3240 4064 3280 4096
rect 3312 4064 3352 4096
rect 3384 4064 3424 4096
rect 3456 4064 3496 4096
rect 3528 4064 3568 4096
rect 3600 4064 3640 4096
rect 3672 4064 3712 4096
rect 3744 4064 3784 4096
rect 3816 4064 3856 4096
rect 3888 4064 3928 4096
rect 3960 4064 4000 4096
rect 0 4024 4000 4064
rect 0 3992 40 4024
rect 72 3992 112 4024
rect 144 3992 184 4024
rect 216 3992 256 4024
rect 288 3992 328 4024
rect 360 3992 400 4024
rect 432 3992 472 4024
rect 504 3992 544 4024
rect 576 3992 616 4024
rect 648 3992 688 4024
rect 720 3992 760 4024
rect 792 3992 832 4024
rect 864 3992 904 4024
rect 936 3992 976 4024
rect 1008 3992 1048 4024
rect 1080 3992 1120 4024
rect 1152 3992 1192 4024
rect 1224 3992 1264 4024
rect 1296 3992 1336 4024
rect 1368 3992 1408 4024
rect 1440 3992 1480 4024
rect 1512 3992 1552 4024
rect 1584 3992 1624 4024
rect 1656 3992 1696 4024
rect 1728 3992 1768 4024
rect 1800 3992 1840 4024
rect 1872 3992 1912 4024
rect 1944 3992 1984 4024
rect 2016 3992 2056 4024
rect 2088 3992 2128 4024
rect 2160 3992 2200 4024
rect 2232 3992 2272 4024
rect 2304 3992 2344 4024
rect 2376 3992 2416 4024
rect 2448 3992 2488 4024
rect 2520 3992 2560 4024
rect 2592 3992 2632 4024
rect 2664 3992 2704 4024
rect 2736 3992 2776 4024
rect 2808 3992 2848 4024
rect 2880 3992 2920 4024
rect 2952 3992 2992 4024
rect 3024 3992 3064 4024
rect 3096 3992 3136 4024
rect 3168 3992 3208 4024
rect 3240 3992 3280 4024
rect 3312 3992 3352 4024
rect 3384 3992 3424 4024
rect 3456 3992 3496 4024
rect 3528 3992 3568 4024
rect 3600 3992 3640 4024
rect 3672 3992 3712 4024
rect 3744 3992 3784 4024
rect 3816 3992 3856 4024
rect 3888 3992 3928 4024
rect 3960 3992 4000 4024
rect 0 3952 4000 3992
rect 0 3920 40 3952
rect 72 3920 112 3952
rect 144 3920 184 3952
rect 216 3920 256 3952
rect 288 3920 328 3952
rect 360 3920 400 3952
rect 432 3920 472 3952
rect 504 3920 544 3952
rect 576 3920 616 3952
rect 648 3920 688 3952
rect 720 3920 760 3952
rect 792 3920 832 3952
rect 864 3920 904 3952
rect 936 3920 976 3952
rect 1008 3920 1048 3952
rect 1080 3920 1120 3952
rect 1152 3920 1192 3952
rect 1224 3920 1264 3952
rect 1296 3920 1336 3952
rect 1368 3920 1408 3952
rect 1440 3920 1480 3952
rect 1512 3920 1552 3952
rect 1584 3920 1624 3952
rect 1656 3920 1696 3952
rect 1728 3920 1768 3952
rect 1800 3920 1840 3952
rect 1872 3920 1912 3952
rect 1944 3920 1984 3952
rect 2016 3920 2056 3952
rect 2088 3920 2128 3952
rect 2160 3920 2200 3952
rect 2232 3920 2272 3952
rect 2304 3920 2344 3952
rect 2376 3920 2416 3952
rect 2448 3920 2488 3952
rect 2520 3920 2560 3952
rect 2592 3920 2632 3952
rect 2664 3920 2704 3952
rect 2736 3920 2776 3952
rect 2808 3920 2848 3952
rect 2880 3920 2920 3952
rect 2952 3920 2992 3952
rect 3024 3920 3064 3952
rect 3096 3920 3136 3952
rect 3168 3920 3208 3952
rect 3240 3920 3280 3952
rect 3312 3920 3352 3952
rect 3384 3920 3424 3952
rect 3456 3920 3496 3952
rect 3528 3920 3568 3952
rect 3600 3920 3640 3952
rect 3672 3920 3712 3952
rect 3744 3920 3784 3952
rect 3816 3920 3856 3952
rect 3888 3920 3928 3952
rect 3960 3920 4000 3952
rect 0 3880 4000 3920
rect 0 3848 40 3880
rect 72 3848 112 3880
rect 144 3848 184 3880
rect 216 3848 256 3880
rect 288 3848 328 3880
rect 360 3848 400 3880
rect 432 3848 472 3880
rect 504 3848 544 3880
rect 576 3848 616 3880
rect 648 3848 688 3880
rect 720 3848 760 3880
rect 792 3848 832 3880
rect 864 3848 904 3880
rect 936 3848 976 3880
rect 1008 3848 1048 3880
rect 1080 3848 1120 3880
rect 1152 3848 1192 3880
rect 1224 3848 1264 3880
rect 1296 3848 1336 3880
rect 1368 3848 1408 3880
rect 1440 3848 1480 3880
rect 1512 3848 1552 3880
rect 1584 3848 1624 3880
rect 1656 3848 1696 3880
rect 1728 3848 1768 3880
rect 1800 3848 1840 3880
rect 1872 3848 1912 3880
rect 1944 3848 1984 3880
rect 2016 3848 2056 3880
rect 2088 3848 2128 3880
rect 2160 3848 2200 3880
rect 2232 3848 2272 3880
rect 2304 3848 2344 3880
rect 2376 3848 2416 3880
rect 2448 3848 2488 3880
rect 2520 3848 2560 3880
rect 2592 3848 2632 3880
rect 2664 3848 2704 3880
rect 2736 3848 2776 3880
rect 2808 3848 2848 3880
rect 2880 3848 2920 3880
rect 2952 3848 2992 3880
rect 3024 3848 3064 3880
rect 3096 3848 3136 3880
rect 3168 3848 3208 3880
rect 3240 3848 3280 3880
rect 3312 3848 3352 3880
rect 3384 3848 3424 3880
rect 3456 3848 3496 3880
rect 3528 3848 3568 3880
rect 3600 3848 3640 3880
rect 3672 3848 3712 3880
rect 3744 3848 3784 3880
rect 3816 3848 3856 3880
rect 3888 3848 3928 3880
rect 3960 3848 4000 3880
rect 0 3808 4000 3848
rect 0 3776 40 3808
rect 72 3776 112 3808
rect 144 3776 184 3808
rect 216 3776 256 3808
rect 288 3776 328 3808
rect 360 3776 400 3808
rect 432 3776 472 3808
rect 504 3776 544 3808
rect 576 3776 616 3808
rect 648 3776 688 3808
rect 720 3776 760 3808
rect 792 3776 832 3808
rect 864 3776 904 3808
rect 936 3776 976 3808
rect 1008 3776 1048 3808
rect 1080 3776 1120 3808
rect 1152 3776 1192 3808
rect 1224 3776 1264 3808
rect 1296 3776 1336 3808
rect 1368 3776 1408 3808
rect 1440 3776 1480 3808
rect 1512 3776 1552 3808
rect 1584 3776 1624 3808
rect 1656 3776 1696 3808
rect 1728 3776 1768 3808
rect 1800 3776 1840 3808
rect 1872 3776 1912 3808
rect 1944 3776 1984 3808
rect 2016 3776 2056 3808
rect 2088 3776 2128 3808
rect 2160 3776 2200 3808
rect 2232 3776 2272 3808
rect 2304 3776 2344 3808
rect 2376 3776 2416 3808
rect 2448 3776 2488 3808
rect 2520 3776 2560 3808
rect 2592 3776 2632 3808
rect 2664 3776 2704 3808
rect 2736 3776 2776 3808
rect 2808 3776 2848 3808
rect 2880 3776 2920 3808
rect 2952 3776 2992 3808
rect 3024 3776 3064 3808
rect 3096 3776 3136 3808
rect 3168 3776 3208 3808
rect 3240 3776 3280 3808
rect 3312 3776 3352 3808
rect 3384 3776 3424 3808
rect 3456 3776 3496 3808
rect 3528 3776 3568 3808
rect 3600 3776 3640 3808
rect 3672 3776 3712 3808
rect 3744 3776 3784 3808
rect 3816 3776 3856 3808
rect 3888 3776 3928 3808
rect 3960 3776 4000 3808
rect 0 3736 4000 3776
rect 0 3704 40 3736
rect 72 3704 112 3736
rect 144 3704 184 3736
rect 216 3704 256 3736
rect 288 3704 328 3736
rect 360 3704 400 3736
rect 432 3704 472 3736
rect 504 3704 544 3736
rect 576 3704 616 3736
rect 648 3704 688 3736
rect 720 3704 760 3736
rect 792 3704 832 3736
rect 864 3704 904 3736
rect 936 3704 976 3736
rect 1008 3704 1048 3736
rect 1080 3704 1120 3736
rect 1152 3704 1192 3736
rect 1224 3704 1264 3736
rect 1296 3704 1336 3736
rect 1368 3704 1408 3736
rect 1440 3704 1480 3736
rect 1512 3704 1552 3736
rect 1584 3704 1624 3736
rect 1656 3704 1696 3736
rect 1728 3704 1768 3736
rect 1800 3704 1840 3736
rect 1872 3704 1912 3736
rect 1944 3704 1984 3736
rect 2016 3704 2056 3736
rect 2088 3704 2128 3736
rect 2160 3704 2200 3736
rect 2232 3704 2272 3736
rect 2304 3704 2344 3736
rect 2376 3704 2416 3736
rect 2448 3704 2488 3736
rect 2520 3704 2560 3736
rect 2592 3704 2632 3736
rect 2664 3704 2704 3736
rect 2736 3704 2776 3736
rect 2808 3704 2848 3736
rect 2880 3704 2920 3736
rect 2952 3704 2992 3736
rect 3024 3704 3064 3736
rect 3096 3704 3136 3736
rect 3168 3704 3208 3736
rect 3240 3704 3280 3736
rect 3312 3704 3352 3736
rect 3384 3704 3424 3736
rect 3456 3704 3496 3736
rect 3528 3704 3568 3736
rect 3600 3704 3640 3736
rect 3672 3704 3712 3736
rect 3744 3704 3784 3736
rect 3816 3704 3856 3736
rect 3888 3704 3928 3736
rect 3960 3704 4000 3736
rect 0 3664 4000 3704
rect 0 3632 40 3664
rect 72 3632 112 3664
rect 144 3632 184 3664
rect 216 3632 256 3664
rect 288 3632 328 3664
rect 360 3632 400 3664
rect 432 3632 472 3664
rect 504 3632 544 3664
rect 576 3632 616 3664
rect 648 3632 688 3664
rect 720 3632 760 3664
rect 792 3632 832 3664
rect 864 3632 904 3664
rect 936 3632 976 3664
rect 1008 3632 1048 3664
rect 1080 3632 1120 3664
rect 1152 3632 1192 3664
rect 1224 3632 1264 3664
rect 1296 3632 1336 3664
rect 1368 3632 1408 3664
rect 1440 3632 1480 3664
rect 1512 3632 1552 3664
rect 1584 3632 1624 3664
rect 1656 3632 1696 3664
rect 1728 3632 1768 3664
rect 1800 3632 1840 3664
rect 1872 3632 1912 3664
rect 1944 3632 1984 3664
rect 2016 3632 2056 3664
rect 2088 3632 2128 3664
rect 2160 3632 2200 3664
rect 2232 3632 2272 3664
rect 2304 3632 2344 3664
rect 2376 3632 2416 3664
rect 2448 3632 2488 3664
rect 2520 3632 2560 3664
rect 2592 3632 2632 3664
rect 2664 3632 2704 3664
rect 2736 3632 2776 3664
rect 2808 3632 2848 3664
rect 2880 3632 2920 3664
rect 2952 3632 2992 3664
rect 3024 3632 3064 3664
rect 3096 3632 3136 3664
rect 3168 3632 3208 3664
rect 3240 3632 3280 3664
rect 3312 3632 3352 3664
rect 3384 3632 3424 3664
rect 3456 3632 3496 3664
rect 3528 3632 3568 3664
rect 3600 3632 3640 3664
rect 3672 3632 3712 3664
rect 3744 3632 3784 3664
rect 3816 3632 3856 3664
rect 3888 3632 3928 3664
rect 3960 3632 4000 3664
rect 0 3592 4000 3632
rect 0 3560 40 3592
rect 72 3560 112 3592
rect 144 3560 184 3592
rect 216 3560 256 3592
rect 288 3560 328 3592
rect 360 3560 400 3592
rect 432 3560 472 3592
rect 504 3560 544 3592
rect 576 3560 616 3592
rect 648 3560 688 3592
rect 720 3560 760 3592
rect 792 3560 832 3592
rect 864 3560 904 3592
rect 936 3560 976 3592
rect 1008 3560 1048 3592
rect 1080 3560 1120 3592
rect 1152 3560 1192 3592
rect 1224 3560 1264 3592
rect 1296 3560 1336 3592
rect 1368 3560 1408 3592
rect 1440 3560 1480 3592
rect 1512 3560 1552 3592
rect 1584 3560 1624 3592
rect 1656 3560 1696 3592
rect 1728 3560 1768 3592
rect 1800 3560 1840 3592
rect 1872 3560 1912 3592
rect 1944 3560 1984 3592
rect 2016 3560 2056 3592
rect 2088 3560 2128 3592
rect 2160 3560 2200 3592
rect 2232 3560 2272 3592
rect 2304 3560 2344 3592
rect 2376 3560 2416 3592
rect 2448 3560 2488 3592
rect 2520 3560 2560 3592
rect 2592 3560 2632 3592
rect 2664 3560 2704 3592
rect 2736 3560 2776 3592
rect 2808 3560 2848 3592
rect 2880 3560 2920 3592
rect 2952 3560 2992 3592
rect 3024 3560 3064 3592
rect 3096 3560 3136 3592
rect 3168 3560 3208 3592
rect 3240 3560 3280 3592
rect 3312 3560 3352 3592
rect 3384 3560 3424 3592
rect 3456 3560 3496 3592
rect 3528 3560 3568 3592
rect 3600 3560 3640 3592
rect 3672 3560 3712 3592
rect 3744 3560 3784 3592
rect 3816 3560 3856 3592
rect 3888 3560 3928 3592
rect 3960 3560 4000 3592
rect 0 3520 4000 3560
rect 0 3488 40 3520
rect 72 3488 112 3520
rect 144 3488 184 3520
rect 216 3488 256 3520
rect 288 3488 328 3520
rect 360 3488 400 3520
rect 432 3488 472 3520
rect 504 3488 544 3520
rect 576 3488 616 3520
rect 648 3488 688 3520
rect 720 3488 760 3520
rect 792 3488 832 3520
rect 864 3488 904 3520
rect 936 3488 976 3520
rect 1008 3488 1048 3520
rect 1080 3488 1120 3520
rect 1152 3488 1192 3520
rect 1224 3488 1264 3520
rect 1296 3488 1336 3520
rect 1368 3488 1408 3520
rect 1440 3488 1480 3520
rect 1512 3488 1552 3520
rect 1584 3488 1624 3520
rect 1656 3488 1696 3520
rect 1728 3488 1768 3520
rect 1800 3488 1840 3520
rect 1872 3488 1912 3520
rect 1944 3488 1984 3520
rect 2016 3488 2056 3520
rect 2088 3488 2128 3520
rect 2160 3488 2200 3520
rect 2232 3488 2272 3520
rect 2304 3488 2344 3520
rect 2376 3488 2416 3520
rect 2448 3488 2488 3520
rect 2520 3488 2560 3520
rect 2592 3488 2632 3520
rect 2664 3488 2704 3520
rect 2736 3488 2776 3520
rect 2808 3488 2848 3520
rect 2880 3488 2920 3520
rect 2952 3488 2992 3520
rect 3024 3488 3064 3520
rect 3096 3488 3136 3520
rect 3168 3488 3208 3520
rect 3240 3488 3280 3520
rect 3312 3488 3352 3520
rect 3384 3488 3424 3520
rect 3456 3488 3496 3520
rect 3528 3488 3568 3520
rect 3600 3488 3640 3520
rect 3672 3488 3712 3520
rect 3744 3488 3784 3520
rect 3816 3488 3856 3520
rect 3888 3488 3928 3520
rect 3960 3488 4000 3520
rect 0 3448 4000 3488
rect 0 3416 40 3448
rect 72 3416 112 3448
rect 144 3416 184 3448
rect 216 3416 256 3448
rect 288 3416 328 3448
rect 360 3416 400 3448
rect 432 3416 472 3448
rect 504 3416 544 3448
rect 576 3416 616 3448
rect 648 3416 688 3448
rect 720 3416 760 3448
rect 792 3416 832 3448
rect 864 3416 904 3448
rect 936 3416 976 3448
rect 1008 3416 1048 3448
rect 1080 3416 1120 3448
rect 1152 3416 1192 3448
rect 1224 3416 1264 3448
rect 1296 3416 1336 3448
rect 1368 3416 1408 3448
rect 1440 3416 1480 3448
rect 1512 3416 1552 3448
rect 1584 3416 1624 3448
rect 1656 3416 1696 3448
rect 1728 3416 1768 3448
rect 1800 3416 1840 3448
rect 1872 3416 1912 3448
rect 1944 3416 1984 3448
rect 2016 3416 2056 3448
rect 2088 3416 2128 3448
rect 2160 3416 2200 3448
rect 2232 3416 2272 3448
rect 2304 3416 2344 3448
rect 2376 3416 2416 3448
rect 2448 3416 2488 3448
rect 2520 3416 2560 3448
rect 2592 3416 2632 3448
rect 2664 3416 2704 3448
rect 2736 3416 2776 3448
rect 2808 3416 2848 3448
rect 2880 3416 2920 3448
rect 2952 3416 2992 3448
rect 3024 3416 3064 3448
rect 3096 3416 3136 3448
rect 3168 3416 3208 3448
rect 3240 3416 3280 3448
rect 3312 3416 3352 3448
rect 3384 3416 3424 3448
rect 3456 3416 3496 3448
rect 3528 3416 3568 3448
rect 3600 3416 3640 3448
rect 3672 3416 3712 3448
rect 3744 3416 3784 3448
rect 3816 3416 3856 3448
rect 3888 3416 3928 3448
rect 3960 3416 4000 3448
rect 0 3376 4000 3416
rect 0 3344 40 3376
rect 72 3344 112 3376
rect 144 3344 184 3376
rect 216 3344 256 3376
rect 288 3344 328 3376
rect 360 3344 400 3376
rect 432 3344 472 3376
rect 504 3344 544 3376
rect 576 3344 616 3376
rect 648 3344 688 3376
rect 720 3344 760 3376
rect 792 3344 832 3376
rect 864 3344 904 3376
rect 936 3344 976 3376
rect 1008 3344 1048 3376
rect 1080 3344 1120 3376
rect 1152 3344 1192 3376
rect 1224 3344 1264 3376
rect 1296 3344 1336 3376
rect 1368 3344 1408 3376
rect 1440 3344 1480 3376
rect 1512 3344 1552 3376
rect 1584 3344 1624 3376
rect 1656 3344 1696 3376
rect 1728 3344 1768 3376
rect 1800 3344 1840 3376
rect 1872 3344 1912 3376
rect 1944 3344 1984 3376
rect 2016 3344 2056 3376
rect 2088 3344 2128 3376
rect 2160 3344 2200 3376
rect 2232 3344 2272 3376
rect 2304 3344 2344 3376
rect 2376 3344 2416 3376
rect 2448 3344 2488 3376
rect 2520 3344 2560 3376
rect 2592 3344 2632 3376
rect 2664 3344 2704 3376
rect 2736 3344 2776 3376
rect 2808 3344 2848 3376
rect 2880 3344 2920 3376
rect 2952 3344 2992 3376
rect 3024 3344 3064 3376
rect 3096 3344 3136 3376
rect 3168 3344 3208 3376
rect 3240 3344 3280 3376
rect 3312 3344 3352 3376
rect 3384 3344 3424 3376
rect 3456 3344 3496 3376
rect 3528 3344 3568 3376
rect 3600 3344 3640 3376
rect 3672 3344 3712 3376
rect 3744 3344 3784 3376
rect 3816 3344 3856 3376
rect 3888 3344 3928 3376
rect 3960 3344 4000 3376
rect 0 3304 4000 3344
rect 0 3272 40 3304
rect 72 3272 112 3304
rect 144 3272 184 3304
rect 216 3272 256 3304
rect 288 3272 328 3304
rect 360 3272 400 3304
rect 432 3272 472 3304
rect 504 3272 544 3304
rect 576 3272 616 3304
rect 648 3272 688 3304
rect 720 3272 760 3304
rect 792 3272 832 3304
rect 864 3272 904 3304
rect 936 3272 976 3304
rect 1008 3272 1048 3304
rect 1080 3272 1120 3304
rect 1152 3272 1192 3304
rect 1224 3272 1264 3304
rect 1296 3272 1336 3304
rect 1368 3272 1408 3304
rect 1440 3272 1480 3304
rect 1512 3272 1552 3304
rect 1584 3272 1624 3304
rect 1656 3272 1696 3304
rect 1728 3272 1768 3304
rect 1800 3272 1840 3304
rect 1872 3272 1912 3304
rect 1944 3272 1984 3304
rect 2016 3272 2056 3304
rect 2088 3272 2128 3304
rect 2160 3272 2200 3304
rect 2232 3272 2272 3304
rect 2304 3272 2344 3304
rect 2376 3272 2416 3304
rect 2448 3272 2488 3304
rect 2520 3272 2560 3304
rect 2592 3272 2632 3304
rect 2664 3272 2704 3304
rect 2736 3272 2776 3304
rect 2808 3272 2848 3304
rect 2880 3272 2920 3304
rect 2952 3272 2992 3304
rect 3024 3272 3064 3304
rect 3096 3272 3136 3304
rect 3168 3272 3208 3304
rect 3240 3272 3280 3304
rect 3312 3272 3352 3304
rect 3384 3272 3424 3304
rect 3456 3272 3496 3304
rect 3528 3272 3568 3304
rect 3600 3272 3640 3304
rect 3672 3272 3712 3304
rect 3744 3272 3784 3304
rect 3816 3272 3856 3304
rect 3888 3272 3928 3304
rect 3960 3272 4000 3304
rect 0 3232 4000 3272
rect 0 3200 40 3232
rect 72 3200 112 3232
rect 144 3200 184 3232
rect 216 3200 256 3232
rect 288 3200 328 3232
rect 360 3200 400 3232
rect 432 3200 472 3232
rect 504 3200 544 3232
rect 576 3200 616 3232
rect 648 3200 688 3232
rect 720 3200 760 3232
rect 792 3200 832 3232
rect 864 3200 904 3232
rect 936 3200 976 3232
rect 1008 3200 1048 3232
rect 1080 3200 1120 3232
rect 1152 3200 1192 3232
rect 1224 3200 1264 3232
rect 1296 3200 1336 3232
rect 1368 3200 1408 3232
rect 1440 3200 1480 3232
rect 1512 3200 1552 3232
rect 1584 3200 1624 3232
rect 1656 3200 1696 3232
rect 1728 3200 1768 3232
rect 1800 3200 1840 3232
rect 1872 3200 1912 3232
rect 1944 3200 1984 3232
rect 2016 3200 2056 3232
rect 2088 3200 2128 3232
rect 2160 3200 2200 3232
rect 2232 3200 2272 3232
rect 2304 3200 2344 3232
rect 2376 3200 2416 3232
rect 2448 3200 2488 3232
rect 2520 3200 2560 3232
rect 2592 3200 2632 3232
rect 2664 3200 2704 3232
rect 2736 3200 2776 3232
rect 2808 3200 2848 3232
rect 2880 3200 2920 3232
rect 2952 3200 2992 3232
rect 3024 3200 3064 3232
rect 3096 3200 3136 3232
rect 3168 3200 3208 3232
rect 3240 3200 3280 3232
rect 3312 3200 3352 3232
rect 3384 3200 3424 3232
rect 3456 3200 3496 3232
rect 3528 3200 3568 3232
rect 3600 3200 3640 3232
rect 3672 3200 3712 3232
rect 3744 3200 3784 3232
rect 3816 3200 3856 3232
rect 3888 3200 3928 3232
rect 3960 3200 4000 3232
rect 0 3160 4000 3200
rect 0 3128 40 3160
rect 72 3128 112 3160
rect 144 3128 184 3160
rect 216 3128 256 3160
rect 288 3128 328 3160
rect 360 3128 400 3160
rect 432 3128 472 3160
rect 504 3128 544 3160
rect 576 3128 616 3160
rect 648 3128 688 3160
rect 720 3128 760 3160
rect 792 3128 832 3160
rect 864 3128 904 3160
rect 936 3128 976 3160
rect 1008 3128 1048 3160
rect 1080 3128 1120 3160
rect 1152 3128 1192 3160
rect 1224 3128 1264 3160
rect 1296 3128 1336 3160
rect 1368 3128 1408 3160
rect 1440 3128 1480 3160
rect 1512 3128 1552 3160
rect 1584 3128 1624 3160
rect 1656 3128 1696 3160
rect 1728 3128 1768 3160
rect 1800 3128 1840 3160
rect 1872 3128 1912 3160
rect 1944 3128 1984 3160
rect 2016 3128 2056 3160
rect 2088 3128 2128 3160
rect 2160 3128 2200 3160
rect 2232 3128 2272 3160
rect 2304 3128 2344 3160
rect 2376 3128 2416 3160
rect 2448 3128 2488 3160
rect 2520 3128 2560 3160
rect 2592 3128 2632 3160
rect 2664 3128 2704 3160
rect 2736 3128 2776 3160
rect 2808 3128 2848 3160
rect 2880 3128 2920 3160
rect 2952 3128 2992 3160
rect 3024 3128 3064 3160
rect 3096 3128 3136 3160
rect 3168 3128 3208 3160
rect 3240 3128 3280 3160
rect 3312 3128 3352 3160
rect 3384 3128 3424 3160
rect 3456 3128 3496 3160
rect 3528 3128 3568 3160
rect 3600 3128 3640 3160
rect 3672 3128 3712 3160
rect 3744 3128 3784 3160
rect 3816 3128 3856 3160
rect 3888 3128 3928 3160
rect 3960 3128 4000 3160
rect 0 3088 4000 3128
rect 0 3056 40 3088
rect 72 3056 112 3088
rect 144 3056 184 3088
rect 216 3056 256 3088
rect 288 3056 328 3088
rect 360 3056 400 3088
rect 432 3056 472 3088
rect 504 3056 544 3088
rect 576 3056 616 3088
rect 648 3056 688 3088
rect 720 3056 760 3088
rect 792 3056 832 3088
rect 864 3056 904 3088
rect 936 3056 976 3088
rect 1008 3056 1048 3088
rect 1080 3056 1120 3088
rect 1152 3056 1192 3088
rect 1224 3056 1264 3088
rect 1296 3056 1336 3088
rect 1368 3056 1408 3088
rect 1440 3056 1480 3088
rect 1512 3056 1552 3088
rect 1584 3056 1624 3088
rect 1656 3056 1696 3088
rect 1728 3056 1768 3088
rect 1800 3056 1840 3088
rect 1872 3056 1912 3088
rect 1944 3056 1984 3088
rect 2016 3056 2056 3088
rect 2088 3056 2128 3088
rect 2160 3056 2200 3088
rect 2232 3056 2272 3088
rect 2304 3056 2344 3088
rect 2376 3056 2416 3088
rect 2448 3056 2488 3088
rect 2520 3056 2560 3088
rect 2592 3056 2632 3088
rect 2664 3056 2704 3088
rect 2736 3056 2776 3088
rect 2808 3056 2848 3088
rect 2880 3056 2920 3088
rect 2952 3056 2992 3088
rect 3024 3056 3064 3088
rect 3096 3056 3136 3088
rect 3168 3056 3208 3088
rect 3240 3056 3280 3088
rect 3312 3056 3352 3088
rect 3384 3056 3424 3088
rect 3456 3056 3496 3088
rect 3528 3056 3568 3088
rect 3600 3056 3640 3088
rect 3672 3056 3712 3088
rect 3744 3056 3784 3088
rect 3816 3056 3856 3088
rect 3888 3056 3928 3088
rect 3960 3056 4000 3088
rect 0 3016 4000 3056
rect 0 2984 40 3016
rect 72 2984 112 3016
rect 144 2984 184 3016
rect 216 2984 256 3016
rect 288 2984 328 3016
rect 360 2984 400 3016
rect 432 2984 472 3016
rect 504 2984 544 3016
rect 576 2984 616 3016
rect 648 2984 688 3016
rect 720 2984 760 3016
rect 792 2984 832 3016
rect 864 2984 904 3016
rect 936 2984 976 3016
rect 1008 2984 1048 3016
rect 1080 2984 1120 3016
rect 1152 2984 1192 3016
rect 1224 2984 1264 3016
rect 1296 2984 1336 3016
rect 1368 2984 1408 3016
rect 1440 2984 1480 3016
rect 1512 2984 1552 3016
rect 1584 2984 1624 3016
rect 1656 2984 1696 3016
rect 1728 2984 1768 3016
rect 1800 2984 1840 3016
rect 1872 2984 1912 3016
rect 1944 2984 1984 3016
rect 2016 2984 2056 3016
rect 2088 2984 2128 3016
rect 2160 2984 2200 3016
rect 2232 2984 2272 3016
rect 2304 2984 2344 3016
rect 2376 2984 2416 3016
rect 2448 2984 2488 3016
rect 2520 2984 2560 3016
rect 2592 2984 2632 3016
rect 2664 2984 2704 3016
rect 2736 2984 2776 3016
rect 2808 2984 2848 3016
rect 2880 2984 2920 3016
rect 2952 2984 2992 3016
rect 3024 2984 3064 3016
rect 3096 2984 3136 3016
rect 3168 2984 3208 3016
rect 3240 2984 3280 3016
rect 3312 2984 3352 3016
rect 3384 2984 3424 3016
rect 3456 2984 3496 3016
rect 3528 2984 3568 3016
rect 3600 2984 3640 3016
rect 3672 2984 3712 3016
rect 3744 2984 3784 3016
rect 3816 2984 3856 3016
rect 3888 2984 3928 3016
rect 3960 2984 4000 3016
rect 0 2944 4000 2984
rect 0 2912 40 2944
rect 72 2912 112 2944
rect 144 2912 184 2944
rect 216 2912 256 2944
rect 288 2912 328 2944
rect 360 2912 400 2944
rect 432 2912 472 2944
rect 504 2912 544 2944
rect 576 2912 616 2944
rect 648 2912 688 2944
rect 720 2912 760 2944
rect 792 2912 832 2944
rect 864 2912 904 2944
rect 936 2912 976 2944
rect 1008 2912 1048 2944
rect 1080 2912 1120 2944
rect 1152 2912 1192 2944
rect 1224 2912 1264 2944
rect 1296 2912 1336 2944
rect 1368 2912 1408 2944
rect 1440 2912 1480 2944
rect 1512 2912 1552 2944
rect 1584 2912 1624 2944
rect 1656 2912 1696 2944
rect 1728 2912 1768 2944
rect 1800 2912 1840 2944
rect 1872 2912 1912 2944
rect 1944 2912 1984 2944
rect 2016 2912 2056 2944
rect 2088 2912 2128 2944
rect 2160 2912 2200 2944
rect 2232 2912 2272 2944
rect 2304 2912 2344 2944
rect 2376 2912 2416 2944
rect 2448 2912 2488 2944
rect 2520 2912 2560 2944
rect 2592 2912 2632 2944
rect 2664 2912 2704 2944
rect 2736 2912 2776 2944
rect 2808 2912 2848 2944
rect 2880 2912 2920 2944
rect 2952 2912 2992 2944
rect 3024 2912 3064 2944
rect 3096 2912 3136 2944
rect 3168 2912 3208 2944
rect 3240 2912 3280 2944
rect 3312 2912 3352 2944
rect 3384 2912 3424 2944
rect 3456 2912 3496 2944
rect 3528 2912 3568 2944
rect 3600 2912 3640 2944
rect 3672 2912 3712 2944
rect 3744 2912 3784 2944
rect 3816 2912 3856 2944
rect 3888 2912 3928 2944
rect 3960 2912 4000 2944
rect 0 2872 4000 2912
rect 0 2840 40 2872
rect 72 2840 112 2872
rect 144 2840 184 2872
rect 216 2840 256 2872
rect 288 2840 328 2872
rect 360 2840 400 2872
rect 432 2840 472 2872
rect 504 2840 544 2872
rect 576 2840 616 2872
rect 648 2840 688 2872
rect 720 2840 760 2872
rect 792 2840 832 2872
rect 864 2840 904 2872
rect 936 2840 976 2872
rect 1008 2840 1048 2872
rect 1080 2840 1120 2872
rect 1152 2840 1192 2872
rect 1224 2840 1264 2872
rect 1296 2840 1336 2872
rect 1368 2840 1408 2872
rect 1440 2840 1480 2872
rect 1512 2840 1552 2872
rect 1584 2840 1624 2872
rect 1656 2840 1696 2872
rect 1728 2840 1768 2872
rect 1800 2840 1840 2872
rect 1872 2840 1912 2872
rect 1944 2840 1984 2872
rect 2016 2840 2056 2872
rect 2088 2840 2128 2872
rect 2160 2840 2200 2872
rect 2232 2840 2272 2872
rect 2304 2840 2344 2872
rect 2376 2840 2416 2872
rect 2448 2840 2488 2872
rect 2520 2840 2560 2872
rect 2592 2840 2632 2872
rect 2664 2840 2704 2872
rect 2736 2840 2776 2872
rect 2808 2840 2848 2872
rect 2880 2840 2920 2872
rect 2952 2840 2992 2872
rect 3024 2840 3064 2872
rect 3096 2840 3136 2872
rect 3168 2840 3208 2872
rect 3240 2840 3280 2872
rect 3312 2840 3352 2872
rect 3384 2840 3424 2872
rect 3456 2840 3496 2872
rect 3528 2840 3568 2872
rect 3600 2840 3640 2872
rect 3672 2840 3712 2872
rect 3744 2840 3784 2872
rect 3816 2840 3856 2872
rect 3888 2840 3928 2872
rect 3960 2840 4000 2872
rect 0 2800 4000 2840
rect 0 2768 40 2800
rect 72 2768 112 2800
rect 144 2768 184 2800
rect 216 2768 256 2800
rect 288 2768 328 2800
rect 360 2768 400 2800
rect 432 2768 472 2800
rect 504 2768 544 2800
rect 576 2768 616 2800
rect 648 2768 688 2800
rect 720 2768 760 2800
rect 792 2768 832 2800
rect 864 2768 904 2800
rect 936 2768 976 2800
rect 1008 2768 1048 2800
rect 1080 2768 1120 2800
rect 1152 2768 1192 2800
rect 1224 2768 1264 2800
rect 1296 2768 1336 2800
rect 1368 2768 1408 2800
rect 1440 2768 1480 2800
rect 1512 2768 1552 2800
rect 1584 2768 1624 2800
rect 1656 2768 1696 2800
rect 1728 2768 1768 2800
rect 1800 2768 1840 2800
rect 1872 2768 1912 2800
rect 1944 2768 1984 2800
rect 2016 2768 2056 2800
rect 2088 2768 2128 2800
rect 2160 2768 2200 2800
rect 2232 2768 2272 2800
rect 2304 2768 2344 2800
rect 2376 2768 2416 2800
rect 2448 2768 2488 2800
rect 2520 2768 2560 2800
rect 2592 2768 2632 2800
rect 2664 2768 2704 2800
rect 2736 2768 2776 2800
rect 2808 2768 2848 2800
rect 2880 2768 2920 2800
rect 2952 2768 2992 2800
rect 3024 2768 3064 2800
rect 3096 2768 3136 2800
rect 3168 2768 3208 2800
rect 3240 2768 3280 2800
rect 3312 2768 3352 2800
rect 3384 2768 3424 2800
rect 3456 2768 3496 2800
rect 3528 2768 3568 2800
rect 3600 2768 3640 2800
rect 3672 2768 3712 2800
rect 3744 2768 3784 2800
rect 3816 2768 3856 2800
rect 3888 2768 3928 2800
rect 3960 2768 4000 2800
rect 0 2728 4000 2768
rect 0 2696 40 2728
rect 72 2696 112 2728
rect 144 2696 184 2728
rect 216 2696 256 2728
rect 288 2696 328 2728
rect 360 2696 400 2728
rect 432 2696 472 2728
rect 504 2696 544 2728
rect 576 2696 616 2728
rect 648 2696 688 2728
rect 720 2696 760 2728
rect 792 2696 832 2728
rect 864 2696 904 2728
rect 936 2696 976 2728
rect 1008 2696 1048 2728
rect 1080 2696 1120 2728
rect 1152 2696 1192 2728
rect 1224 2696 1264 2728
rect 1296 2696 1336 2728
rect 1368 2696 1408 2728
rect 1440 2696 1480 2728
rect 1512 2696 1552 2728
rect 1584 2696 1624 2728
rect 1656 2696 1696 2728
rect 1728 2696 1768 2728
rect 1800 2696 1840 2728
rect 1872 2696 1912 2728
rect 1944 2696 1984 2728
rect 2016 2696 2056 2728
rect 2088 2696 2128 2728
rect 2160 2696 2200 2728
rect 2232 2696 2272 2728
rect 2304 2696 2344 2728
rect 2376 2696 2416 2728
rect 2448 2696 2488 2728
rect 2520 2696 2560 2728
rect 2592 2696 2632 2728
rect 2664 2696 2704 2728
rect 2736 2696 2776 2728
rect 2808 2696 2848 2728
rect 2880 2696 2920 2728
rect 2952 2696 2992 2728
rect 3024 2696 3064 2728
rect 3096 2696 3136 2728
rect 3168 2696 3208 2728
rect 3240 2696 3280 2728
rect 3312 2696 3352 2728
rect 3384 2696 3424 2728
rect 3456 2696 3496 2728
rect 3528 2696 3568 2728
rect 3600 2696 3640 2728
rect 3672 2696 3712 2728
rect 3744 2696 3784 2728
rect 3816 2696 3856 2728
rect 3888 2696 3928 2728
rect 3960 2696 4000 2728
rect 0 2656 4000 2696
rect 0 2624 40 2656
rect 72 2624 112 2656
rect 144 2624 184 2656
rect 216 2624 256 2656
rect 288 2624 328 2656
rect 360 2624 400 2656
rect 432 2624 472 2656
rect 504 2624 544 2656
rect 576 2624 616 2656
rect 648 2624 688 2656
rect 720 2624 760 2656
rect 792 2624 832 2656
rect 864 2624 904 2656
rect 936 2624 976 2656
rect 1008 2624 1048 2656
rect 1080 2624 1120 2656
rect 1152 2624 1192 2656
rect 1224 2624 1264 2656
rect 1296 2624 1336 2656
rect 1368 2624 1408 2656
rect 1440 2624 1480 2656
rect 1512 2624 1552 2656
rect 1584 2624 1624 2656
rect 1656 2624 1696 2656
rect 1728 2624 1768 2656
rect 1800 2624 1840 2656
rect 1872 2624 1912 2656
rect 1944 2624 1984 2656
rect 2016 2624 2056 2656
rect 2088 2624 2128 2656
rect 2160 2624 2200 2656
rect 2232 2624 2272 2656
rect 2304 2624 2344 2656
rect 2376 2624 2416 2656
rect 2448 2624 2488 2656
rect 2520 2624 2560 2656
rect 2592 2624 2632 2656
rect 2664 2624 2704 2656
rect 2736 2624 2776 2656
rect 2808 2624 2848 2656
rect 2880 2624 2920 2656
rect 2952 2624 2992 2656
rect 3024 2624 3064 2656
rect 3096 2624 3136 2656
rect 3168 2624 3208 2656
rect 3240 2624 3280 2656
rect 3312 2624 3352 2656
rect 3384 2624 3424 2656
rect 3456 2624 3496 2656
rect 3528 2624 3568 2656
rect 3600 2624 3640 2656
rect 3672 2624 3712 2656
rect 3744 2624 3784 2656
rect 3816 2624 3856 2656
rect 3888 2624 3928 2656
rect 3960 2624 4000 2656
rect 0 2584 4000 2624
rect 0 2552 40 2584
rect 72 2552 112 2584
rect 144 2552 184 2584
rect 216 2552 256 2584
rect 288 2552 328 2584
rect 360 2552 400 2584
rect 432 2552 472 2584
rect 504 2552 544 2584
rect 576 2552 616 2584
rect 648 2552 688 2584
rect 720 2552 760 2584
rect 792 2552 832 2584
rect 864 2552 904 2584
rect 936 2552 976 2584
rect 1008 2552 1048 2584
rect 1080 2552 1120 2584
rect 1152 2552 1192 2584
rect 1224 2552 1264 2584
rect 1296 2552 1336 2584
rect 1368 2552 1408 2584
rect 1440 2552 1480 2584
rect 1512 2552 1552 2584
rect 1584 2552 1624 2584
rect 1656 2552 1696 2584
rect 1728 2552 1768 2584
rect 1800 2552 1840 2584
rect 1872 2552 1912 2584
rect 1944 2552 1984 2584
rect 2016 2552 2056 2584
rect 2088 2552 2128 2584
rect 2160 2552 2200 2584
rect 2232 2552 2272 2584
rect 2304 2552 2344 2584
rect 2376 2552 2416 2584
rect 2448 2552 2488 2584
rect 2520 2552 2560 2584
rect 2592 2552 2632 2584
rect 2664 2552 2704 2584
rect 2736 2552 2776 2584
rect 2808 2552 2848 2584
rect 2880 2552 2920 2584
rect 2952 2552 2992 2584
rect 3024 2552 3064 2584
rect 3096 2552 3136 2584
rect 3168 2552 3208 2584
rect 3240 2552 3280 2584
rect 3312 2552 3352 2584
rect 3384 2552 3424 2584
rect 3456 2552 3496 2584
rect 3528 2552 3568 2584
rect 3600 2552 3640 2584
rect 3672 2552 3712 2584
rect 3744 2552 3784 2584
rect 3816 2552 3856 2584
rect 3888 2552 3928 2584
rect 3960 2552 4000 2584
rect 0 2512 4000 2552
rect 0 2480 40 2512
rect 72 2480 112 2512
rect 144 2480 184 2512
rect 216 2480 256 2512
rect 288 2480 328 2512
rect 360 2480 400 2512
rect 432 2480 472 2512
rect 504 2480 544 2512
rect 576 2480 616 2512
rect 648 2480 688 2512
rect 720 2480 760 2512
rect 792 2480 832 2512
rect 864 2480 904 2512
rect 936 2480 976 2512
rect 1008 2480 1048 2512
rect 1080 2480 1120 2512
rect 1152 2480 1192 2512
rect 1224 2480 1264 2512
rect 1296 2480 1336 2512
rect 1368 2480 1408 2512
rect 1440 2480 1480 2512
rect 1512 2480 1552 2512
rect 1584 2480 1624 2512
rect 1656 2480 1696 2512
rect 1728 2480 1768 2512
rect 1800 2480 1840 2512
rect 1872 2480 1912 2512
rect 1944 2480 1984 2512
rect 2016 2480 2056 2512
rect 2088 2480 2128 2512
rect 2160 2480 2200 2512
rect 2232 2480 2272 2512
rect 2304 2480 2344 2512
rect 2376 2480 2416 2512
rect 2448 2480 2488 2512
rect 2520 2480 2560 2512
rect 2592 2480 2632 2512
rect 2664 2480 2704 2512
rect 2736 2480 2776 2512
rect 2808 2480 2848 2512
rect 2880 2480 2920 2512
rect 2952 2480 2992 2512
rect 3024 2480 3064 2512
rect 3096 2480 3136 2512
rect 3168 2480 3208 2512
rect 3240 2480 3280 2512
rect 3312 2480 3352 2512
rect 3384 2480 3424 2512
rect 3456 2480 3496 2512
rect 3528 2480 3568 2512
rect 3600 2480 3640 2512
rect 3672 2480 3712 2512
rect 3744 2480 3784 2512
rect 3816 2480 3856 2512
rect 3888 2480 3928 2512
rect 3960 2480 4000 2512
rect 0 2440 4000 2480
rect 0 2408 40 2440
rect 72 2408 112 2440
rect 144 2408 184 2440
rect 216 2408 256 2440
rect 288 2408 328 2440
rect 360 2408 400 2440
rect 432 2408 472 2440
rect 504 2408 544 2440
rect 576 2408 616 2440
rect 648 2408 688 2440
rect 720 2408 760 2440
rect 792 2408 832 2440
rect 864 2408 904 2440
rect 936 2408 976 2440
rect 1008 2408 1048 2440
rect 1080 2408 1120 2440
rect 1152 2408 1192 2440
rect 1224 2408 1264 2440
rect 1296 2408 1336 2440
rect 1368 2408 1408 2440
rect 1440 2408 1480 2440
rect 1512 2408 1552 2440
rect 1584 2408 1624 2440
rect 1656 2408 1696 2440
rect 1728 2408 1768 2440
rect 1800 2408 1840 2440
rect 1872 2408 1912 2440
rect 1944 2408 1984 2440
rect 2016 2408 2056 2440
rect 2088 2408 2128 2440
rect 2160 2408 2200 2440
rect 2232 2408 2272 2440
rect 2304 2408 2344 2440
rect 2376 2408 2416 2440
rect 2448 2408 2488 2440
rect 2520 2408 2560 2440
rect 2592 2408 2632 2440
rect 2664 2408 2704 2440
rect 2736 2408 2776 2440
rect 2808 2408 2848 2440
rect 2880 2408 2920 2440
rect 2952 2408 2992 2440
rect 3024 2408 3064 2440
rect 3096 2408 3136 2440
rect 3168 2408 3208 2440
rect 3240 2408 3280 2440
rect 3312 2408 3352 2440
rect 3384 2408 3424 2440
rect 3456 2408 3496 2440
rect 3528 2408 3568 2440
rect 3600 2408 3640 2440
rect 3672 2408 3712 2440
rect 3744 2408 3784 2440
rect 3816 2408 3856 2440
rect 3888 2408 3928 2440
rect 3960 2408 4000 2440
rect 0 2368 4000 2408
rect 0 2336 40 2368
rect 72 2336 112 2368
rect 144 2336 184 2368
rect 216 2336 256 2368
rect 288 2336 328 2368
rect 360 2336 400 2368
rect 432 2336 472 2368
rect 504 2336 544 2368
rect 576 2336 616 2368
rect 648 2336 688 2368
rect 720 2336 760 2368
rect 792 2336 832 2368
rect 864 2336 904 2368
rect 936 2336 976 2368
rect 1008 2336 1048 2368
rect 1080 2336 1120 2368
rect 1152 2336 1192 2368
rect 1224 2336 1264 2368
rect 1296 2336 1336 2368
rect 1368 2336 1408 2368
rect 1440 2336 1480 2368
rect 1512 2336 1552 2368
rect 1584 2336 1624 2368
rect 1656 2336 1696 2368
rect 1728 2336 1768 2368
rect 1800 2336 1840 2368
rect 1872 2336 1912 2368
rect 1944 2336 1984 2368
rect 2016 2336 2056 2368
rect 2088 2336 2128 2368
rect 2160 2336 2200 2368
rect 2232 2336 2272 2368
rect 2304 2336 2344 2368
rect 2376 2336 2416 2368
rect 2448 2336 2488 2368
rect 2520 2336 2560 2368
rect 2592 2336 2632 2368
rect 2664 2336 2704 2368
rect 2736 2336 2776 2368
rect 2808 2336 2848 2368
rect 2880 2336 2920 2368
rect 2952 2336 2992 2368
rect 3024 2336 3064 2368
rect 3096 2336 3136 2368
rect 3168 2336 3208 2368
rect 3240 2336 3280 2368
rect 3312 2336 3352 2368
rect 3384 2336 3424 2368
rect 3456 2336 3496 2368
rect 3528 2336 3568 2368
rect 3600 2336 3640 2368
rect 3672 2336 3712 2368
rect 3744 2336 3784 2368
rect 3816 2336 3856 2368
rect 3888 2336 3928 2368
rect 3960 2336 4000 2368
rect 0 2296 4000 2336
rect 0 2264 40 2296
rect 72 2264 112 2296
rect 144 2264 184 2296
rect 216 2264 256 2296
rect 288 2264 328 2296
rect 360 2264 400 2296
rect 432 2264 472 2296
rect 504 2264 544 2296
rect 576 2264 616 2296
rect 648 2264 688 2296
rect 720 2264 760 2296
rect 792 2264 832 2296
rect 864 2264 904 2296
rect 936 2264 976 2296
rect 1008 2264 1048 2296
rect 1080 2264 1120 2296
rect 1152 2264 1192 2296
rect 1224 2264 1264 2296
rect 1296 2264 1336 2296
rect 1368 2264 1408 2296
rect 1440 2264 1480 2296
rect 1512 2264 1552 2296
rect 1584 2264 1624 2296
rect 1656 2264 1696 2296
rect 1728 2264 1768 2296
rect 1800 2264 1840 2296
rect 1872 2264 1912 2296
rect 1944 2264 1984 2296
rect 2016 2264 2056 2296
rect 2088 2264 2128 2296
rect 2160 2264 2200 2296
rect 2232 2264 2272 2296
rect 2304 2264 2344 2296
rect 2376 2264 2416 2296
rect 2448 2264 2488 2296
rect 2520 2264 2560 2296
rect 2592 2264 2632 2296
rect 2664 2264 2704 2296
rect 2736 2264 2776 2296
rect 2808 2264 2848 2296
rect 2880 2264 2920 2296
rect 2952 2264 2992 2296
rect 3024 2264 3064 2296
rect 3096 2264 3136 2296
rect 3168 2264 3208 2296
rect 3240 2264 3280 2296
rect 3312 2264 3352 2296
rect 3384 2264 3424 2296
rect 3456 2264 3496 2296
rect 3528 2264 3568 2296
rect 3600 2264 3640 2296
rect 3672 2264 3712 2296
rect 3744 2264 3784 2296
rect 3816 2264 3856 2296
rect 3888 2264 3928 2296
rect 3960 2264 4000 2296
rect 0 2224 4000 2264
rect 0 2192 40 2224
rect 72 2192 112 2224
rect 144 2192 184 2224
rect 216 2192 256 2224
rect 288 2192 328 2224
rect 360 2192 400 2224
rect 432 2192 472 2224
rect 504 2192 544 2224
rect 576 2192 616 2224
rect 648 2192 688 2224
rect 720 2192 760 2224
rect 792 2192 832 2224
rect 864 2192 904 2224
rect 936 2192 976 2224
rect 1008 2192 1048 2224
rect 1080 2192 1120 2224
rect 1152 2192 1192 2224
rect 1224 2192 1264 2224
rect 1296 2192 1336 2224
rect 1368 2192 1408 2224
rect 1440 2192 1480 2224
rect 1512 2192 1552 2224
rect 1584 2192 1624 2224
rect 1656 2192 1696 2224
rect 1728 2192 1768 2224
rect 1800 2192 1840 2224
rect 1872 2192 1912 2224
rect 1944 2192 1984 2224
rect 2016 2192 2056 2224
rect 2088 2192 2128 2224
rect 2160 2192 2200 2224
rect 2232 2192 2272 2224
rect 2304 2192 2344 2224
rect 2376 2192 2416 2224
rect 2448 2192 2488 2224
rect 2520 2192 2560 2224
rect 2592 2192 2632 2224
rect 2664 2192 2704 2224
rect 2736 2192 2776 2224
rect 2808 2192 2848 2224
rect 2880 2192 2920 2224
rect 2952 2192 2992 2224
rect 3024 2192 3064 2224
rect 3096 2192 3136 2224
rect 3168 2192 3208 2224
rect 3240 2192 3280 2224
rect 3312 2192 3352 2224
rect 3384 2192 3424 2224
rect 3456 2192 3496 2224
rect 3528 2192 3568 2224
rect 3600 2192 3640 2224
rect 3672 2192 3712 2224
rect 3744 2192 3784 2224
rect 3816 2192 3856 2224
rect 3888 2192 3928 2224
rect 3960 2192 4000 2224
rect 0 2152 4000 2192
rect 0 2120 40 2152
rect 72 2120 112 2152
rect 144 2120 184 2152
rect 216 2120 256 2152
rect 288 2120 328 2152
rect 360 2120 400 2152
rect 432 2120 472 2152
rect 504 2120 544 2152
rect 576 2120 616 2152
rect 648 2120 688 2152
rect 720 2120 760 2152
rect 792 2120 832 2152
rect 864 2120 904 2152
rect 936 2120 976 2152
rect 1008 2120 1048 2152
rect 1080 2120 1120 2152
rect 1152 2120 1192 2152
rect 1224 2120 1264 2152
rect 1296 2120 1336 2152
rect 1368 2120 1408 2152
rect 1440 2120 1480 2152
rect 1512 2120 1552 2152
rect 1584 2120 1624 2152
rect 1656 2120 1696 2152
rect 1728 2120 1768 2152
rect 1800 2120 1840 2152
rect 1872 2120 1912 2152
rect 1944 2120 1984 2152
rect 2016 2120 2056 2152
rect 2088 2120 2128 2152
rect 2160 2120 2200 2152
rect 2232 2120 2272 2152
rect 2304 2120 2344 2152
rect 2376 2120 2416 2152
rect 2448 2120 2488 2152
rect 2520 2120 2560 2152
rect 2592 2120 2632 2152
rect 2664 2120 2704 2152
rect 2736 2120 2776 2152
rect 2808 2120 2848 2152
rect 2880 2120 2920 2152
rect 2952 2120 2992 2152
rect 3024 2120 3064 2152
rect 3096 2120 3136 2152
rect 3168 2120 3208 2152
rect 3240 2120 3280 2152
rect 3312 2120 3352 2152
rect 3384 2120 3424 2152
rect 3456 2120 3496 2152
rect 3528 2120 3568 2152
rect 3600 2120 3640 2152
rect 3672 2120 3712 2152
rect 3744 2120 3784 2152
rect 3816 2120 3856 2152
rect 3888 2120 3928 2152
rect 3960 2120 4000 2152
rect 0 2080 4000 2120
rect 0 2048 40 2080
rect 72 2048 112 2080
rect 144 2048 184 2080
rect 216 2048 256 2080
rect 288 2048 328 2080
rect 360 2048 400 2080
rect 432 2048 472 2080
rect 504 2048 544 2080
rect 576 2048 616 2080
rect 648 2048 688 2080
rect 720 2048 760 2080
rect 792 2048 832 2080
rect 864 2048 904 2080
rect 936 2048 976 2080
rect 1008 2048 1048 2080
rect 1080 2048 1120 2080
rect 1152 2048 1192 2080
rect 1224 2048 1264 2080
rect 1296 2048 1336 2080
rect 1368 2048 1408 2080
rect 1440 2048 1480 2080
rect 1512 2048 1552 2080
rect 1584 2048 1624 2080
rect 1656 2048 1696 2080
rect 1728 2048 1768 2080
rect 1800 2048 1840 2080
rect 1872 2048 1912 2080
rect 1944 2048 1984 2080
rect 2016 2048 2056 2080
rect 2088 2048 2128 2080
rect 2160 2048 2200 2080
rect 2232 2048 2272 2080
rect 2304 2048 2344 2080
rect 2376 2048 2416 2080
rect 2448 2048 2488 2080
rect 2520 2048 2560 2080
rect 2592 2048 2632 2080
rect 2664 2048 2704 2080
rect 2736 2048 2776 2080
rect 2808 2048 2848 2080
rect 2880 2048 2920 2080
rect 2952 2048 2992 2080
rect 3024 2048 3064 2080
rect 3096 2048 3136 2080
rect 3168 2048 3208 2080
rect 3240 2048 3280 2080
rect 3312 2048 3352 2080
rect 3384 2048 3424 2080
rect 3456 2048 3496 2080
rect 3528 2048 3568 2080
rect 3600 2048 3640 2080
rect 3672 2048 3712 2080
rect 3744 2048 3784 2080
rect 3816 2048 3856 2080
rect 3888 2048 3928 2080
rect 3960 2048 4000 2080
rect 0 2008 4000 2048
rect 0 1976 40 2008
rect 72 1976 112 2008
rect 144 1976 184 2008
rect 216 1976 256 2008
rect 288 1976 328 2008
rect 360 1976 400 2008
rect 432 1976 472 2008
rect 504 1976 544 2008
rect 576 1976 616 2008
rect 648 1976 688 2008
rect 720 1976 760 2008
rect 792 1976 832 2008
rect 864 1976 904 2008
rect 936 1976 976 2008
rect 1008 1976 1048 2008
rect 1080 1976 1120 2008
rect 1152 1976 1192 2008
rect 1224 1976 1264 2008
rect 1296 1976 1336 2008
rect 1368 1976 1408 2008
rect 1440 1976 1480 2008
rect 1512 1976 1552 2008
rect 1584 1976 1624 2008
rect 1656 1976 1696 2008
rect 1728 1976 1768 2008
rect 1800 1976 1840 2008
rect 1872 1976 1912 2008
rect 1944 1976 1984 2008
rect 2016 1976 2056 2008
rect 2088 1976 2128 2008
rect 2160 1976 2200 2008
rect 2232 1976 2272 2008
rect 2304 1976 2344 2008
rect 2376 1976 2416 2008
rect 2448 1976 2488 2008
rect 2520 1976 2560 2008
rect 2592 1976 2632 2008
rect 2664 1976 2704 2008
rect 2736 1976 2776 2008
rect 2808 1976 2848 2008
rect 2880 1976 2920 2008
rect 2952 1976 2992 2008
rect 3024 1976 3064 2008
rect 3096 1976 3136 2008
rect 3168 1976 3208 2008
rect 3240 1976 3280 2008
rect 3312 1976 3352 2008
rect 3384 1976 3424 2008
rect 3456 1976 3496 2008
rect 3528 1976 3568 2008
rect 3600 1976 3640 2008
rect 3672 1976 3712 2008
rect 3744 1976 3784 2008
rect 3816 1976 3856 2008
rect 3888 1976 3928 2008
rect 3960 1976 4000 2008
rect 0 1936 4000 1976
rect 0 1904 40 1936
rect 72 1904 112 1936
rect 144 1904 184 1936
rect 216 1904 256 1936
rect 288 1904 328 1936
rect 360 1904 400 1936
rect 432 1904 472 1936
rect 504 1904 544 1936
rect 576 1904 616 1936
rect 648 1904 688 1936
rect 720 1904 760 1936
rect 792 1904 832 1936
rect 864 1904 904 1936
rect 936 1904 976 1936
rect 1008 1904 1048 1936
rect 1080 1904 1120 1936
rect 1152 1904 1192 1936
rect 1224 1904 1264 1936
rect 1296 1904 1336 1936
rect 1368 1904 1408 1936
rect 1440 1904 1480 1936
rect 1512 1904 1552 1936
rect 1584 1904 1624 1936
rect 1656 1904 1696 1936
rect 1728 1904 1768 1936
rect 1800 1904 1840 1936
rect 1872 1904 1912 1936
rect 1944 1904 1984 1936
rect 2016 1904 2056 1936
rect 2088 1904 2128 1936
rect 2160 1904 2200 1936
rect 2232 1904 2272 1936
rect 2304 1904 2344 1936
rect 2376 1904 2416 1936
rect 2448 1904 2488 1936
rect 2520 1904 2560 1936
rect 2592 1904 2632 1936
rect 2664 1904 2704 1936
rect 2736 1904 2776 1936
rect 2808 1904 2848 1936
rect 2880 1904 2920 1936
rect 2952 1904 2992 1936
rect 3024 1904 3064 1936
rect 3096 1904 3136 1936
rect 3168 1904 3208 1936
rect 3240 1904 3280 1936
rect 3312 1904 3352 1936
rect 3384 1904 3424 1936
rect 3456 1904 3496 1936
rect 3528 1904 3568 1936
rect 3600 1904 3640 1936
rect 3672 1904 3712 1936
rect 3744 1904 3784 1936
rect 3816 1904 3856 1936
rect 3888 1904 3928 1936
rect 3960 1904 4000 1936
rect 0 1864 4000 1904
rect 0 1832 40 1864
rect 72 1832 112 1864
rect 144 1832 184 1864
rect 216 1832 256 1864
rect 288 1832 328 1864
rect 360 1832 400 1864
rect 432 1832 472 1864
rect 504 1832 544 1864
rect 576 1832 616 1864
rect 648 1832 688 1864
rect 720 1832 760 1864
rect 792 1832 832 1864
rect 864 1832 904 1864
rect 936 1832 976 1864
rect 1008 1832 1048 1864
rect 1080 1832 1120 1864
rect 1152 1832 1192 1864
rect 1224 1832 1264 1864
rect 1296 1832 1336 1864
rect 1368 1832 1408 1864
rect 1440 1832 1480 1864
rect 1512 1832 1552 1864
rect 1584 1832 1624 1864
rect 1656 1832 1696 1864
rect 1728 1832 1768 1864
rect 1800 1832 1840 1864
rect 1872 1832 1912 1864
rect 1944 1832 1984 1864
rect 2016 1832 2056 1864
rect 2088 1832 2128 1864
rect 2160 1832 2200 1864
rect 2232 1832 2272 1864
rect 2304 1832 2344 1864
rect 2376 1832 2416 1864
rect 2448 1832 2488 1864
rect 2520 1832 2560 1864
rect 2592 1832 2632 1864
rect 2664 1832 2704 1864
rect 2736 1832 2776 1864
rect 2808 1832 2848 1864
rect 2880 1832 2920 1864
rect 2952 1832 2992 1864
rect 3024 1832 3064 1864
rect 3096 1832 3136 1864
rect 3168 1832 3208 1864
rect 3240 1832 3280 1864
rect 3312 1832 3352 1864
rect 3384 1832 3424 1864
rect 3456 1832 3496 1864
rect 3528 1832 3568 1864
rect 3600 1832 3640 1864
rect 3672 1832 3712 1864
rect 3744 1832 3784 1864
rect 3816 1832 3856 1864
rect 3888 1832 3928 1864
rect 3960 1832 4000 1864
rect 0 1792 4000 1832
rect 0 1760 40 1792
rect 72 1760 112 1792
rect 144 1760 184 1792
rect 216 1760 256 1792
rect 288 1760 328 1792
rect 360 1760 400 1792
rect 432 1760 472 1792
rect 504 1760 544 1792
rect 576 1760 616 1792
rect 648 1760 688 1792
rect 720 1760 760 1792
rect 792 1760 832 1792
rect 864 1760 904 1792
rect 936 1760 976 1792
rect 1008 1760 1048 1792
rect 1080 1760 1120 1792
rect 1152 1760 1192 1792
rect 1224 1760 1264 1792
rect 1296 1760 1336 1792
rect 1368 1760 1408 1792
rect 1440 1760 1480 1792
rect 1512 1760 1552 1792
rect 1584 1760 1624 1792
rect 1656 1760 1696 1792
rect 1728 1760 1768 1792
rect 1800 1760 1840 1792
rect 1872 1760 1912 1792
rect 1944 1760 1984 1792
rect 2016 1760 2056 1792
rect 2088 1760 2128 1792
rect 2160 1760 2200 1792
rect 2232 1760 2272 1792
rect 2304 1760 2344 1792
rect 2376 1760 2416 1792
rect 2448 1760 2488 1792
rect 2520 1760 2560 1792
rect 2592 1760 2632 1792
rect 2664 1760 2704 1792
rect 2736 1760 2776 1792
rect 2808 1760 2848 1792
rect 2880 1760 2920 1792
rect 2952 1760 2992 1792
rect 3024 1760 3064 1792
rect 3096 1760 3136 1792
rect 3168 1760 3208 1792
rect 3240 1760 3280 1792
rect 3312 1760 3352 1792
rect 3384 1760 3424 1792
rect 3456 1760 3496 1792
rect 3528 1760 3568 1792
rect 3600 1760 3640 1792
rect 3672 1760 3712 1792
rect 3744 1760 3784 1792
rect 3816 1760 3856 1792
rect 3888 1760 3928 1792
rect 3960 1760 4000 1792
rect 0 1720 4000 1760
rect 0 1688 40 1720
rect 72 1688 112 1720
rect 144 1688 184 1720
rect 216 1688 256 1720
rect 288 1688 328 1720
rect 360 1688 400 1720
rect 432 1688 472 1720
rect 504 1688 544 1720
rect 576 1688 616 1720
rect 648 1688 688 1720
rect 720 1688 760 1720
rect 792 1688 832 1720
rect 864 1688 904 1720
rect 936 1688 976 1720
rect 1008 1688 1048 1720
rect 1080 1688 1120 1720
rect 1152 1688 1192 1720
rect 1224 1688 1264 1720
rect 1296 1688 1336 1720
rect 1368 1688 1408 1720
rect 1440 1688 1480 1720
rect 1512 1688 1552 1720
rect 1584 1688 1624 1720
rect 1656 1688 1696 1720
rect 1728 1688 1768 1720
rect 1800 1688 1840 1720
rect 1872 1688 1912 1720
rect 1944 1688 1984 1720
rect 2016 1688 2056 1720
rect 2088 1688 2128 1720
rect 2160 1688 2200 1720
rect 2232 1688 2272 1720
rect 2304 1688 2344 1720
rect 2376 1688 2416 1720
rect 2448 1688 2488 1720
rect 2520 1688 2560 1720
rect 2592 1688 2632 1720
rect 2664 1688 2704 1720
rect 2736 1688 2776 1720
rect 2808 1688 2848 1720
rect 2880 1688 2920 1720
rect 2952 1688 2992 1720
rect 3024 1688 3064 1720
rect 3096 1688 3136 1720
rect 3168 1688 3208 1720
rect 3240 1688 3280 1720
rect 3312 1688 3352 1720
rect 3384 1688 3424 1720
rect 3456 1688 3496 1720
rect 3528 1688 3568 1720
rect 3600 1688 3640 1720
rect 3672 1688 3712 1720
rect 3744 1688 3784 1720
rect 3816 1688 3856 1720
rect 3888 1688 3928 1720
rect 3960 1688 4000 1720
rect 0 1648 4000 1688
rect 0 1616 40 1648
rect 72 1616 112 1648
rect 144 1616 184 1648
rect 216 1616 256 1648
rect 288 1616 328 1648
rect 360 1616 400 1648
rect 432 1616 472 1648
rect 504 1616 544 1648
rect 576 1616 616 1648
rect 648 1616 688 1648
rect 720 1616 760 1648
rect 792 1616 832 1648
rect 864 1616 904 1648
rect 936 1616 976 1648
rect 1008 1616 1048 1648
rect 1080 1616 1120 1648
rect 1152 1616 1192 1648
rect 1224 1616 1264 1648
rect 1296 1616 1336 1648
rect 1368 1616 1408 1648
rect 1440 1616 1480 1648
rect 1512 1616 1552 1648
rect 1584 1616 1624 1648
rect 1656 1616 1696 1648
rect 1728 1616 1768 1648
rect 1800 1616 1840 1648
rect 1872 1616 1912 1648
rect 1944 1616 1984 1648
rect 2016 1616 2056 1648
rect 2088 1616 2128 1648
rect 2160 1616 2200 1648
rect 2232 1616 2272 1648
rect 2304 1616 2344 1648
rect 2376 1616 2416 1648
rect 2448 1616 2488 1648
rect 2520 1616 2560 1648
rect 2592 1616 2632 1648
rect 2664 1616 2704 1648
rect 2736 1616 2776 1648
rect 2808 1616 2848 1648
rect 2880 1616 2920 1648
rect 2952 1616 2992 1648
rect 3024 1616 3064 1648
rect 3096 1616 3136 1648
rect 3168 1616 3208 1648
rect 3240 1616 3280 1648
rect 3312 1616 3352 1648
rect 3384 1616 3424 1648
rect 3456 1616 3496 1648
rect 3528 1616 3568 1648
rect 3600 1616 3640 1648
rect 3672 1616 3712 1648
rect 3744 1616 3784 1648
rect 3816 1616 3856 1648
rect 3888 1616 3928 1648
rect 3960 1616 4000 1648
rect 0 1576 4000 1616
rect 0 1544 40 1576
rect 72 1544 112 1576
rect 144 1544 184 1576
rect 216 1544 256 1576
rect 288 1544 328 1576
rect 360 1544 400 1576
rect 432 1544 472 1576
rect 504 1544 544 1576
rect 576 1544 616 1576
rect 648 1544 688 1576
rect 720 1544 760 1576
rect 792 1544 832 1576
rect 864 1544 904 1576
rect 936 1544 976 1576
rect 1008 1544 1048 1576
rect 1080 1544 1120 1576
rect 1152 1544 1192 1576
rect 1224 1544 1264 1576
rect 1296 1544 1336 1576
rect 1368 1544 1408 1576
rect 1440 1544 1480 1576
rect 1512 1544 1552 1576
rect 1584 1544 1624 1576
rect 1656 1544 1696 1576
rect 1728 1544 1768 1576
rect 1800 1544 1840 1576
rect 1872 1544 1912 1576
rect 1944 1544 1984 1576
rect 2016 1544 2056 1576
rect 2088 1544 2128 1576
rect 2160 1544 2200 1576
rect 2232 1544 2272 1576
rect 2304 1544 2344 1576
rect 2376 1544 2416 1576
rect 2448 1544 2488 1576
rect 2520 1544 2560 1576
rect 2592 1544 2632 1576
rect 2664 1544 2704 1576
rect 2736 1544 2776 1576
rect 2808 1544 2848 1576
rect 2880 1544 2920 1576
rect 2952 1544 2992 1576
rect 3024 1544 3064 1576
rect 3096 1544 3136 1576
rect 3168 1544 3208 1576
rect 3240 1544 3280 1576
rect 3312 1544 3352 1576
rect 3384 1544 3424 1576
rect 3456 1544 3496 1576
rect 3528 1544 3568 1576
rect 3600 1544 3640 1576
rect 3672 1544 3712 1576
rect 3744 1544 3784 1576
rect 3816 1544 3856 1576
rect 3888 1544 3928 1576
rect 3960 1544 4000 1576
rect 0 1504 4000 1544
rect 0 1472 40 1504
rect 72 1472 112 1504
rect 144 1472 184 1504
rect 216 1472 256 1504
rect 288 1472 328 1504
rect 360 1472 400 1504
rect 432 1472 472 1504
rect 504 1472 544 1504
rect 576 1472 616 1504
rect 648 1472 688 1504
rect 720 1472 760 1504
rect 792 1472 832 1504
rect 864 1472 904 1504
rect 936 1472 976 1504
rect 1008 1472 1048 1504
rect 1080 1472 1120 1504
rect 1152 1472 1192 1504
rect 1224 1472 1264 1504
rect 1296 1472 1336 1504
rect 1368 1472 1408 1504
rect 1440 1472 1480 1504
rect 1512 1472 1552 1504
rect 1584 1472 1624 1504
rect 1656 1472 1696 1504
rect 1728 1472 1768 1504
rect 1800 1472 1840 1504
rect 1872 1472 1912 1504
rect 1944 1472 1984 1504
rect 2016 1472 2056 1504
rect 2088 1472 2128 1504
rect 2160 1472 2200 1504
rect 2232 1472 2272 1504
rect 2304 1472 2344 1504
rect 2376 1472 2416 1504
rect 2448 1472 2488 1504
rect 2520 1472 2560 1504
rect 2592 1472 2632 1504
rect 2664 1472 2704 1504
rect 2736 1472 2776 1504
rect 2808 1472 2848 1504
rect 2880 1472 2920 1504
rect 2952 1472 2992 1504
rect 3024 1472 3064 1504
rect 3096 1472 3136 1504
rect 3168 1472 3208 1504
rect 3240 1472 3280 1504
rect 3312 1472 3352 1504
rect 3384 1472 3424 1504
rect 3456 1472 3496 1504
rect 3528 1472 3568 1504
rect 3600 1472 3640 1504
rect 3672 1472 3712 1504
rect 3744 1472 3784 1504
rect 3816 1472 3856 1504
rect 3888 1472 3928 1504
rect 3960 1472 4000 1504
rect 0 1432 4000 1472
rect 0 1400 40 1432
rect 72 1400 112 1432
rect 144 1400 184 1432
rect 216 1400 256 1432
rect 288 1400 328 1432
rect 360 1400 400 1432
rect 432 1400 472 1432
rect 504 1400 544 1432
rect 576 1400 616 1432
rect 648 1400 688 1432
rect 720 1400 760 1432
rect 792 1400 832 1432
rect 864 1400 904 1432
rect 936 1400 976 1432
rect 1008 1400 1048 1432
rect 1080 1400 1120 1432
rect 1152 1400 1192 1432
rect 1224 1400 1264 1432
rect 1296 1400 1336 1432
rect 1368 1400 1408 1432
rect 1440 1400 1480 1432
rect 1512 1400 1552 1432
rect 1584 1400 1624 1432
rect 1656 1400 1696 1432
rect 1728 1400 1768 1432
rect 1800 1400 1840 1432
rect 1872 1400 1912 1432
rect 1944 1400 1984 1432
rect 2016 1400 2056 1432
rect 2088 1400 2128 1432
rect 2160 1400 2200 1432
rect 2232 1400 2272 1432
rect 2304 1400 2344 1432
rect 2376 1400 2416 1432
rect 2448 1400 2488 1432
rect 2520 1400 2560 1432
rect 2592 1400 2632 1432
rect 2664 1400 2704 1432
rect 2736 1400 2776 1432
rect 2808 1400 2848 1432
rect 2880 1400 2920 1432
rect 2952 1400 2992 1432
rect 3024 1400 3064 1432
rect 3096 1400 3136 1432
rect 3168 1400 3208 1432
rect 3240 1400 3280 1432
rect 3312 1400 3352 1432
rect 3384 1400 3424 1432
rect 3456 1400 3496 1432
rect 3528 1400 3568 1432
rect 3600 1400 3640 1432
rect 3672 1400 3712 1432
rect 3744 1400 3784 1432
rect 3816 1400 3856 1432
rect 3888 1400 3928 1432
rect 3960 1400 4000 1432
rect 0 1360 4000 1400
rect 0 1328 40 1360
rect 72 1328 112 1360
rect 144 1328 184 1360
rect 216 1328 256 1360
rect 288 1328 328 1360
rect 360 1328 400 1360
rect 432 1328 472 1360
rect 504 1328 544 1360
rect 576 1328 616 1360
rect 648 1328 688 1360
rect 720 1328 760 1360
rect 792 1328 832 1360
rect 864 1328 904 1360
rect 936 1328 976 1360
rect 1008 1328 1048 1360
rect 1080 1328 1120 1360
rect 1152 1328 1192 1360
rect 1224 1328 1264 1360
rect 1296 1328 1336 1360
rect 1368 1328 1408 1360
rect 1440 1328 1480 1360
rect 1512 1328 1552 1360
rect 1584 1328 1624 1360
rect 1656 1328 1696 1360
rect 1728 1328 1768 1360
rect 1800 1328 1840 1360
rect 1872 1328 1912 1360
rect 1944 1328 1984 1360
rect 2016 1328 2056 1360
rect 2088 1328 2128 1360
rect 2160 1328 2200 1360
rect 2232 1328 2272 1360
rect 2304 1328 2344 1360
rect 2376 1328 2416 1360
rect 2448 1328 2488 1360
rect 2520 1328 2560 1360
rect 2592 1328 2632 1360
rect 2664 1328 2704 1360
rect 2736 1328 2776 1360
rect 2808 1328 2848 1360
rect 2880 1328 2920 1360
rect 2952 1328 2992 1360
rect 3024 1328 3064 1360
rect 3096 1328 3136 1360
rect 3168 1328 3208 1360
rect 3240 1328 3280 1360
rect 3312 1328 3352 1360
rect 3384 1328 3424 1360
rect 3456 1328 3496 1360
rect 3528 1328 3568 1360
rect 3600 1328 3640 1360
rect 3672 1328 3712 1360
rect 3744 1328 3784 1360
rect 3816 1328 3856 1360
rect 3888 1328 3928 1360
rect 3960 1328 4000 1360
rect 0 1288 4000 1328
rect 0 1256 40 1288
rect 72 1256 112 1288
rect 144 1256 184 1288
rect 216 1256 256 1288
rect 288 1256 328 1288
rect 360 1256 400 1288
rect 432 1256 472 1288
rect 504 1256 544 1288
rect 576 1256 616 1288
rect 648 1256 688 1288
rect 720 1256 760 1288
rect 792 1256 832 1288
rect 864 1256 904 1288
rect 936 1256 976 1288
rect 1008 1256 1048 1288
rect 1080 1256 1120 1288
rect 1152 1256 1192 1288
rect 1224 1256 1264 1288
rect 1296 1256 1336 1288
rect 1368 1256 1408 1288
rect 1440 1256 1480 1288
rect 1512 1256 1552 1288
rect 1584 1256 1624 1288
rect 1656 1256 1696 1288
rect 1728 1256 1768 1288
rect 1800 1256 1840 1288
rect 1872 1256 1912 1288
rect 1944 1256 1984 1288
rect 2016 1256 2056 1288
rect 2088 1256 2128 1288
rect 2160 1256 2200 1288
rect 2232 1256 2272 1288
rect 2304 1256 2344 1288
rect 2376 1256 2416 1288
rect 2448 1256 2488 1288
rect 2520 1256 2560 1288
rect 2592 1256 2632 1288
rect 2664 1256 2704 1288
rect 2736 1256 2776 1288
rect 2808 1256 2848 1288
rect 2880 1256 2920 1288
rect 2952 1256 2992 1288
rect 3024 1256 3064 1288
rect 3096 1256 3136 1288
rect 3168 1256 3208 1288
rect 3240 1256 3280 1288
rect 3312 1256 3352 1288
rect 3384 1256 3424 1288
rect 3456 1256 3496 1288
rect 3528 1256 3568 1288
rect 3600 1256 3640 1288
rect 3672 1256 3712 1288
rect 3744 1256 3784 1288
rect 3816 1256 3856 1288
rect 3888 1256 3928 1288
rect 3960 1256 4000 1288
rect 0 1200 4000 1256
<< metal3 >>
rect 0 32000 4000 35600
rect 0 28000 4000 31600
rect 0 25200 4000 26800
rect 0 18700 4000 23800
rect 0 13200 4000 18300
rect 0 6900 4000 12000
rect 0 1400 4000 6500
<< metal4 >>
rect 0 32440 4000 35600
rect 0 28000 4000 31160
rect 0 25200 4000 26800
rect 0 18700 4000 23800
rect 0 13200 4000 18300
rect 0 6900 4000 12000
rect 0 1400 4000 6500
<< metal5 >>
rect 0 32000 4000 35600
rect 0 28000 4000 31600
rect 0 25200 4000 26800
rect 0 18700 4000 23800
rect 0 13200 4000 18300
rect 0 6900 4000 12000
rect 0 1400 4000 6500
<< metal6 >>
rect 0 32000 4000 35600
rect 0 28000 4000 31600
rect 0 25200 4000 26800
rect 0 18700 4000 23800
rect 0 13200 4000 18300
rect 0 6900 4000 12000
rect 0 1400 4000 6500
<< metal7 >>
rect 0 25500 4000 26500
rect 0 19000 4000 23500
rect 0 13500 4000 18000
rect 0 7200 4000 11700
rect 0 1700 4000 6200
<< labels >>
rlabel metal3 s 0 32000 4000 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 4000 31600 4 vss
port 1 nsew
rlabel metal3 s 0 18700 4000 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 13200 4000 18300 4 iovdd
port 4 nsew
rlabel metal3 s 0 25200 4000 26800 4 iovss
port 3 nsew
rlabel metal3 s 0 6900 4000 12000 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 4000 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 4000 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 4000 35600 4 vss
port 1 nsew
rlabel metal4 s 0 18700 4000 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 13200 4000 18300 4 iovdd
port 4 nsew
rlabel metal4 s 0 25200 4000 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 6900 4000 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 4000 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 4000 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 4000 35600 4 vss
port 1 nsew
rlabel metal5 s 0 18700 4000 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 13200 4000 18300 4 iovdd
port 4 nsew
rlabel metal5 s 0 25200 4000 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 6900 4000 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 4000 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 4000 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 4000 35600 4 vss
port 1 nsew
rlabel metal6 s 0 18700 4000 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 13200 4000 18300 4 iovdd
port 4 nsew
rlabel metal6 s 0 25200 4000 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 6900 4000 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 4000 6500 4 iovss
port 3 nsew
rlabel metal7 s 0 13500 4000 18000 4 iovdd
port 4 nsew
rlabel metal7 s 0 19000 4000 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 1700 4000 6200 4 iovss
port 3 nsew
rlabel metal7 s 0 7200 4000 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 25500 4000 26500 4 iovss
port 3 nsew
flabel comment s 441 13233 441 13233 0 FreeSans 1600 0 0 0 sub!
flabel comment s 434 18360 434 18360 0 FreeSans 1600 0 0 0 sub!
flabel comment s 441 23404 441 23404 0 FreeSans 1600 0 0 0 sub!
flabel comment s 571 31393 571 31393 0 FreeSans 1600 0 0 0 sub!
flabel metal1 s 655 8487 1204 9203 0 FreeSans 51 0 0 0 iovdd
port 4 nsew
flabel metal1 s 777 5239 1311 6017 0 FreeSans 51 0 0 0 iovdd
port 4 nsew
flabel metal1 s 224 31392 268 31409 0 FreeSans 51 0 0 0 vss
port 1 nsew
flabel metal1 s 500 16997 1242 17573 0 FreeSans 51 0 0 0 iovss
port 3 nsew
flabel metal1 s 500 21732 1242 22308 0 FreeSans 51 0 0 0 iovss
port 3 nsew
flabel metal1 s 500 26019 1242 26595 0 FreeSans 51 0 0 0 iovss
port 3 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 4000 36000
string GDS_END 5305084
string GDS_FILE sg13g2_io.gds
string GDS_START 4087280
<< end >>
