magic
tech ihp-sg13g2
magscale 1 2
timestamp 1749471858
<< metal1 >>
rect 3163 1428 15266 2104
rect 3163 -821 3336 1428
rect 3427 1289 3499 1428
rect 3535 1321 3907 1373
rect 3427 -683 3509 1289
rect 3671 393 3771 1321
rect 4063 1289 4135 1428
rect 4171 1321 4543 1373
rect 3671 213 3681 393
rect 3761 213 3771 393
rect 3671 -715 3771 213
rect 3933 -150 4015 1289
rect 3933 -330 3943 -150
rect 4005 -330 4015 -150
rect 3933 -683 4015 -330
rect 4063 -683 4145 1289
rect 4307 393 4407 1321
rect 4875 1289 4947 1428
rect 4983 1321 5355 1373
rect 4307 213 4317 393
rect 4397 213 4407 393
rect 4307 -715 4407 213
rect 4569 -150 4651 1289
rect 4569 -330 4579 -150
rect 4641 -330 4651 -150
rect 4569 -683 4651 -330
rect 4875 -683 4957 1289
rect 5119 393 5219 1321
rect 5511 1289 5583 1428
rect 5619 1321 5991 1373
rect 5119 213 5129 393
rect 5209 213 5219 393
rect 5119 -150 5219 213
rect 5119 -330 5129 -150
rect 5209 -330 5219 -150
rect 5119 -715 5219 -330
rect 5381 -150 5463 1289
rect 5381 -330 5391 -150
rect 5453 -330 5463 -150
rect 5381 -683 5463 -330
rect 5511 -683 5593 1289
rect 5755 393 5855 1321
rect 6323 1289 6395 1428
rect 6431 1321 6803 1373
rect 5755 213 5765 393
rect 5845 213 5855 393
rect 5755 -150 5855 213
rect 5755 -330 5765 -150
rect 5845 -330 5855 -150
rect 5755 -715 5855 -330
rect 6017 -150 6099 1289
rect 6017 -330 6027 -150
rect 6089 -330 6099 -150
rect 6017 -683 6099 -330
rect 6323 -683 6405 1289
rect 6567 393 6667 1321
rect 6959 1289 7031 1428
rect 7067 1321 7439 1373
rect 6567 213 6577 393
rect 6657 213 6667 393
rect 6567 -150 6667 213
rect 6567 -330 6577 -150
rect 6657 -330 6667 -150
rect 6567 -715 6667 -330
rect 6829 -150 6911 1289
rect 6829 -330 6839 -150
rect 6901 -330 6911 -150
rect 6829 -683 6911 -330
rect 6959 -683 7041 1289
rect 7203 393 7303 1321
rect 7771 1289 7843 1428
rect 7879 1321 8251 1373
rect 7203 213 7213 393
rect 7293 213 7303 393
rect 7203 -150 7303 213
rect 7203 -330 7213 -150
rect 7293 -330 7303 -150
rect 7203 -715 7303 -330
rect 7465 -150 7547 1289
rect 7465 -330 7475 -150
rect 7537 -330 7547 -150
rect 7465 -683 7547 -330
rect 7771 -683 7853 1289
rect 8015 393 8115 1321
rect 8407 1289 8479 1428
rect 8515 1321 8887 1373
rect 8015 213 8025 393
rect 8105 213 8115 393
rect 8015 -715 8115 213
rect 8277 -150 8359 1289
rect 8277 -330 8287 -150
rect 8349 -330 8359 -150
rect 8277 -683 8359 -330
rect 8407 -683 8489 1289
rect 8651 393 8751 1321
rect 9043 1289 9115 1428
rect 9151 1321 9523 1373
rect 8651 213 8661 393
rect 8741 213 8751 393
rect 8651 -715 8751 213
rect 8913 -150 8995 1289
rect 8913 -330 8923 -150
rect 8985 -330 8995 -150
rect 8913 -683 8995 -330
rect 9043 -683 9125 1289
rect 9287 393 9387 1321
rect 9679 1289 9751 1428
rect 9787 1321 10159 1373
rect 9287 213 9297 393
rect 9377 213 9387 393
rect 9287 -715 9387 213
rect 9549 -150 9631 1289
rect 9549 -330 9559 -150
rect 9621 -330 9631 -150
rect 9549 -683 9631 -330
rect 9679 -683 9761 1289
rect 9923 393 10023 1321
rect 10315 1289 10387 1428
rect 10423 1321 10795 1373
rect 9923 213 9933 393
rect 10013 213 10023 393
rect 9923 -715 10023 213
rect 10185 -150 10267 1289
rect 10185 -330 10195 -150
rect 10257 -330 10267 -150
rect 10185 -683 10267 -330
rect 10315 -683 10397 1289
rect 10559 393 10659 1321
rect 10951 1289 11023 1428
rect 11059 1321 11431 1373
rect 10559 213 10569 393
rect 10649 213 10659 393
rect 10559 -715 10659 213
rect 10821 -150 10903 1289
rect 10821 -330 10831 -150
rect 10893 -330 10903 -150
rect 10821 -683 10903 -330
rect 10951 -683 11033 1289
rect 11195 393 11295 1321
rect 11587 1289 11659 1428
rect 11695 1321 12067 1373
rect 11195 213 11205 393
rect 11285 213 11295 393
rect 11195 -715 11295 213
rect 11457 -150 11539 1289
rect 11457 -330 11467 -150
rect 11529 -330 11539 -150
rect 11457 -683 11539 -330
rect 11587 -683 11669 1289
rect 11831 393 11931 1321
rect 12223 1289 12295 1428
rect 12331 1321 12703 1373
rect 11831 213 11841 393
rect 11921 213 11931 393
rect 11831 -715 11931 213
rect 12093 -150 12175 1289
rect 12093 -330 12103 -150
rect 12165 -330 12175 -150
rect 12093 -683 12175 -330
rect 12223 -683 12305 1289
rect 12467 393 12567 1321
rect 12859 1289 12931 1428
rect 12967 1321 13339 1373
rect 12467 213 12477 393
rect 12557 213 12567 393
rect 12467 -715 12567 213
rect 12729 -150 12811 1289
rect 12729 -330 12739 -150
rect 12801 -330 12811 -150
rect 12729 -683 12811 -330
rect 12859 -683 12941 1289
rect 13103 393 13203 1321
rect 13495 1289 13567 1428
rect 13603 1321 13975 1373
rect 13103 213 13113 393
rect 13193 213 13203 393
rect 13103 -715 13203 213
rect 13365 -150 13447 1289
rect 13365 -330 13375 -150
rect 13437 -330 13447 -150
rect 13365 -683 13447 -330
rect 13495 -683 13577 1289
rect 13739 393 13839 1321
rect 13739 213 13749 393
rect 13829 213 13839 393
rect 13739 -715 13839 213
rect 14001 -150 14083 1289
rect 14001 -330 14011 -150
rect 14073 -330 14083 -150
rect 14001 -683 14083 -330
rect 3535 -767 3907 -715
rect 4171 -767 4543 -715
rect 4983 -767 5355 -715
rect 5619 -767 5991 -715
rect 6431 -767 6803 -715
rect 7067 -767 7439 -715
rect 7879 -767 8251 -715
rect 8515 -767 8887 -715
rect 9151 -767 9523 -715
rect 9787 -767 10159 -715
rect 10423 -767 10795 -715
rect 11059 -767 11431 -715
rect 11695 -767 12067 -715
rect 12331 -767 12703 -715
rect 12967 -767 13339 -715
rect 13603 -767 13975 -715
rect 14172 -821 15266 1428
rect 3163 -1242 15266 -821
rect 3163 -1259 10131 -1242
rect 3368 -1398 3668 -1388
rect 3368 -1673 3378 -1398
rect 3658 -1673 3668 -1398
rect 3368 -11669 3668 -1673
rect 3879 -1521 8983 -1388
rect 3879 -8762 4264 -1521
rect 4403 -1620 6375 -1610
rect 4403 -1684 5842 -1620
rect 6022 -1684 6375 -1620
rect 4403 -1694 6375 -1684
rect 6699 -1620 8671 -1610
rect 6699 -1684 7052 -1620
rect 7232 -1684 8671 -1620
rect 6699 -1694 8671 -1684
rect 4319 -1856 4371 -1720
rect 6407 -1856 6459 -1720
rect 4319 -1866 6459 -1856
rect 4319 -1946 4756 -1866
rect 4936 -1946 6459 -1866
rect 4319 -1956 6459 -1946
rect 4319 -2092 4371 -1956
rect 6407 -2092 6459 -1956
rect 6615 -1856 6667 -1720
rect 8703 -1856 8755 -1720
rect 6615 -1866 8755 -1856
rect 6615 -1946 8138 -1866
rect 8318 -1946 8755 -1866
rect 6615 -1956 8755 -1946
rect 6615 -2092 6667 -1956
rect 8703 -2092 8755 -1956
rect 4403 -2128 6375 -2118
rect 4403 -2192 5299 -2128
rect 5479 -2192 6375 -2128
rect 4403 -2202 6375 -2192
rect 6699 -2128 8671 -2118
rect 6699 -2192 7595 -2128
rect 7775 -2192 8671 -2128
rect 6699 -2202 8671 -2192
rect 4403 -2256 6375 -2246
rect 4403 -2320 5842 -2256
rect 6022 -2320 6375 -2256
rect 4403 -2330 6375 -2320
rect 6699 -2256 8671 -2246
rect 6699 -2320 7052 -2256
rect 7232 -2320 8671 -2256
rect 6699 -2330 8671 -2320
rect 4319 -2492 4371 -2356
rect 6407 -2492 6459 -2356
rect 4319 -2502 6459 -2492
rect 4319 -2582 4756 -2502
rect 4936 -2582 6459 -2502
rect 4319 -2592 6459 -2582
rect 4319 -2728 4371 -2592
rect 6407 -2728 6459 -2592
rect 6615 -2492 6667 -2356
rect 8703 -2492 8755 -2356
rect 6615 -2502 8755 -2492
rect 6615 -2582 8138 -2502
rect 8318 -2582 8755 -2502
rect 6615 -2592 8755 -2582
rect 6615 -2728 6667 -2592
rect 8703 -2728 8755 -2592
rect 4403 -2764 6375 -2754
rect 4403 -2828 5299 -2764
rect 5479 -2828 6375 -2764
rect 4403 -2838 6375 -2828
rect 6699 -2764 8671 -2754
rect 6699 -2828 7595 -2764
rect 7775 -2828 8671 -2764
rect 6699 -2838 8671 -2828
rect 4403 -2892 6375 -2882
rect 4403 -2956 5842 -2892
rect 6022 -2956 6375 -2892
rect 4403 -2966 6375 -2956
rect 6699 -2892 8671 -2882
rect 6699 -2956 7052 -2892
rect 7232 -2956 8671 -2892
rect 6699 -2966 8671 -2956
rect 4319 -3128 4371 -2992
rect 6407 -3128 6459 -2992
rect 4319 -3138 6459 -3128
rect 4319 -3218 4756 -3138
rect 4936 -3218 6459 -3138
rect 4319 -3228 6459 -3218
rect 4319 -3364 4371 -3228
rect 6407 -3364 6459 -3228
rect 6615 -3128 6667 -2992
rect 8703 -3128 8755 -2992
rect 6615 -3138 8755 -3128
rect 6615 -3218 8138 -3138
rect 8318 -3218 8755 -3138
rect 6615 -3228 8755 -3218
rect 6615 -3364 6667 -3228
rect 8703 -3364 8755 -3228
rect 4403 -3400 6375 -3390
rect 4403 -3464 5299 -3400
rect 5479 -3464 6375 -3400
rect 4403 -3474 6375 -3464
rect 6699 -3400 8671 -3390
rect 6699 -3464 7595 -3400
rect 7775 -3464 8671 -3400
rect 6699 -3474 8671 -3464
rect 4403 -3528 6375 -3518
rect 4403 -3592 5842 -3528
rect 6022 -3592 6375 -3528
rect 4403 -3602 6375 -3592
rect 6699 -3528 8671 -3518
rect 6699 -3592 7052 -3528
rect 7232 -3592 8671 -3528
rect 6699 -3602 8671 -3592
rect 4319 -3764 4371 -3628
rect 6407 -3764 6459 -3628
rect 4319 -3774 6459 -3764
rect 4319 -3854 4756 -3774
rect 4936 -3854 6459 -3774
rect 4319 -3864 6459 -3854
rect 4319 -4000 4371 -3864
rect 6407 -4000 6459 -3864
rect 6615 -3764 6667 -3628
rect 8703 -3764 8755 -3628
rect 6615 -3774 8755 -3764
rect 6615 -3854 8138 -3774
rect 8318 -3854 8755 -3774
rect 6615 -3864 8755 -3854
rect 6615 -4000 6667 -3864
rect 8703 -4000 8755 -3864
rect 4403 -4036 6375 -4026
rect 4403 -4100 5299 -4036
rect 5479 -4100 6375 -4036
rect 4403 -4110 6375 -4100
rect 6699 -4036 8671 -4026
rect 6699 -4100 7595 -4036
rect 7775 -4100 8671 -4036
rect 6699 -4110 8671 -4100
rect 4403 -4164 6375 -4154
rect 4403 -4228 5842 -4164
rect 6022 -4228 6375 -4164
rect 4403 -4238 6375 -4228
rect 6699 -4164 8671 -4154
rect 6699 -4228 7052 -4164
rect 7232 -4228 8671 -4164
rect 6699 -4238 8671 -4228
rect 4319 -4400 4371 -4264
rect 6407 -4400 6459 -4264
rect 4319 -4410 6459 -4400
rect 4319 -4490 4756 -4410
rect 4936 -4490 6459 -4410
rect 4319 -4500 6459 -4490
rect 4319 -4636 4371 -4500
rect 6407 -4636 6459 -4500
rect 6615 -4400 6667 -4264
rect 8703 -4400 8755 -4264
rect 6615 -4410 8755 -4400
rect 6615 -4490 8138 -4410
rect 8318 -4490 8755 -4410
rect 6615 -4500 8755 -4490
rect 6615 -4636 6667 -4500
rect 8703 -4636 8755 -4500
rect 4403 -4672 6375 -4662
rect 4403 -4736 5299 -4672
rect 5479 -4736 6375 -4672
rect 4403 -4746 6375 -4736
rect 6699 -4672 8671 -4662
rect 6699 -4736 7595 -4672
rect 7775 -4736 8671 -4672
rect 6699 -4746 8671 -4736
rect 4403 -4800 6375 -4790
rect 4403 -4864 5842 -4800
rect 6022 -4864 6375 -4800
rect 4403 -4874 6375 -4864
rect 6699 -4800 8671 -4790
rect 6699 -4864 7052 -4800
rect 7232 -4864 8671 -4800
rect 6699 -4874 8671 -4864
rect 4319 -5036 4371 -4900
rect 6407 -5036 6459 -4900
rect 4319 -5046 6459 -5036
rect 4319 -5126 4756 -5046
rect 4936 -5126 6459 -5046
rect 4319 -5136 6459 -5126
rect 4319 -5272 4371 -5136
rect 6407 -5272 6459 -5136
rect 6615 -5036 6667 -4900
rect 8703 -5036 8755 -4900
rect 6615 -5046 8755 -5036
rect 6615 -5126 8138 -5046
rect 8318 -5126 8755 -5046
rect 6615 -5136 8755 -5126
rect 6615 -5272 6667 -5136
rect 8703 -5272 8755 -5136
rect 4403 -5308 6375 -5298
rect 4403 -5372 5299 -5308
rect 5479 -5372 6375 -5308
rect 4403 -5382 6375 -5372
rect 6699 -5308 8671 -5298
rect 6699 -5372 7595 -5308
rect 7775 -5372 8671 -5308
rect 6699 -5382 8671 -5372
rect 4403 -5436 6375 -5426
rect 4403 -5500 5842 -5436
rect 6022 -5500 6375 -5436
rect 4403 -5510 6375 -5500
rect 6699 -5436 8671 -5426
rect 6699 -5500 7052 -5436
rect 7232 -5500 8671 -5436
rect 6699 -5510 8671 -5500
rect 4319 -5672 4371 -5536
rect 6407 -5672 6459 -5536
rect 4319 -5682 6459 -5672
rect 4319 -5762 4756 -5682
rect 4936 -5762 6459 -5682
rect 4319 -5772 6459 -5762
rect 4319 -5908 4371 -5772
rect 6407 -5908 6459 -5772
rect 6615 -5672 6667 -5536
rect 8703 -5672 8755 -5536
rect 6615 -5682 8755 -5672
rect 6615 -5762 8138 -5682
rect 8318 -5762 8755 -5682
rect 6615 -5772 8755 -5762
rect 6615 -5908 6667 -5772
rect 8703 -5908 8755 -5772
rect 4403 -5944 6375 -5934
rect 4403 -6008 5299 -5944
rect 5479 -6008 6375 -5944
rect 4403 -6018 6375 -6008
rect 6699 -5944 8671 -5934
rect 6699 -6008 7595 -5944
rect 7775 -6008 8671 -5944
rect 6699 -6018 8671 -6008
rect 4403 -6072 6375 -6062
rect 4403 -6136 5842 -6072
rect 6022 -6136 6375 -6072
rect 4403 -6146 6375 -6136
rect 6699 -6072 8671 -6062
rect 6699 -6136 7052 -6072
rect 7232 -6136 8671 -6072
rect 6699 -6146 8671 -6136
rect 4319 -6308 4371 -6172
rect 6407 -6308 6459 -6172
rect 4319 -6318 6459 -6308
rect 4319 -6398 4756 -6318
rect 4936 -6398 6459 -6318
rect 4319 -6408 6459 -6398
rect 4319 -6544 4371 -6408
rect 6407 -6544 6459 -6408
rect 6615 -6308 6667 -6172
rect 8703 -6308 8755 -6172
rect 6615 -6318 8755 -6308
rect 6615 -6398 8138 -6318
rect 8318 -6398 8755 -6318
rect 6615 -6408 8755 -6398
rect 6615 -6544 6667 -6408
rect 8703 -6544 8755 -6408
rect 4403 -6580 6375 -6570
rect 4403 -6644 5299 -6580
rect 5479 -6644 6375 -6580
rect 4403 -6654 6375 -6644
rect 6699 -6580 8671 -6570
rect 6699 -6644 7595 -6580
rect 7775 -6644 8671 -6580
rect 6699 -6654 8671 -6644
rect 4403 -6708 6375 -6698
rect 4403 -6772 5842 -6708
rect 6022 -6772 6375 -6708
rect 4403 -6782 6375 -6772
rect 6699 -6708 8671 -6698
rect 6699 -6772 7052 -6708
rect 7232 -6772 8671 -6708
rect 6699 -6782 8671 -6772
rect 4319 -6944 4371 -6808
rect 6407 -6944 6459 -6808
rect 4319 -6954 6459 -6944
rect 4319 -7034 4756 -6954
rect 4936 -7034 6459 -6954
rect 4319 -7044 6459 -7034
rect 4319 -7180 4371 -7044
rect 6407 -7180 6459 -7044
rect 6615 -6944 6667 -6808
rect 8703 -6944 8755 -6808
rect 6615 -6954 8755 -6944
rect 6615 -7034 8138 -6954
rect 8318 -7034 8755 -6954
rect 6615 -7044 8755 -7034
rect 6615 -7180 6667 -7044
rect 8703 -7180 8755 -7044
rect 4403 -7216 6375 -7206
rect 4403 -7280 5299 -7216
rect 5479 -7280 6375 -7216
rect 4403 -7290 6375 -7280
rect 6699 -7216 8671 -7206
rect 6699 -7280 7595 -7216
rect 7775 -7280 8671 -7216
rect 6699 -7290 8671 -7280
rect 4403 -7344 6375 -7334
rect 4403 -7408 5842 -7344
rect 6022 -7408 6375 -7344
rect 4403 -7418 6375 -7408
rect 6699 -7344 8671 -7334
rect 6699 -7408 7052 -7344
rect 7232 -7408 8671 -7344
rect 6699 -7418 8671 -7408
rect 4319 -7580 4371 -7444
rect 6407 -7580 6459 -7444
rect 4319 -7590 6459 -7580
rect 4319 -7670 4756 -7590
rect 4936 -7670 6459 -7590
rect 4319 -7680 6459 -7670
rect 4319 -7816 4371 -7680
rect 6407 -7816 6459 -7680
rect 6615 -7580 6667 -7444
rect 8703 -7580 8755 -7444
rect 6615 -7590 8755 -7580
rect 6615 -7670 8138 -7590
rect 8318 -7670 8755 -7590
rect 6615 -7680 8755 -7670
rect 6615 -7816 6667 -7680
rect 8703 -7816 8755 -7680
rect 4403 -7852 6375 -7842
rect 4403 -7916 5299 -7852
rect 5479 -7916 6375 -7852
rect 4403 -7926 6375 -7916
rect 6699 -7852 8671 -7842
rect 6699 -7916 7595 -7852
rect 7775 -7916 8671 -7852
rect 6699 -7926 8671 -7916
rect 6128 -8140 6328 -8130
rect 6128 -8236 6138 -8140
rect 6318 -8236 6328 -8140
rect 6128 -8585 6328 -8236
rect 6128 -8681 6138 -8585
rect 6318 -8681 6328 -8585
rect 6128 -8691 6328 -8681
rect 8813 -8762 8983 -1521
rect 9548 -1653 10131 -1259
rect 10711 -1653 13172 -1242
rect 13752 -1653 15266 -1242
rect 9548 -1663 15266 -1653
rect 9548 -8184 9725 -1663
rect 11894 -1761 11990 -1751
rect 9780 -1861 9822 -1761
rect 9864 -1771 11836 -1761
rect 9864 -1825 10988 -1771
rect 11568 -1825 11836 -1771
rect 9864 -1835 11836 -1825
rect 11894 -1861 11904 -1761
rect 9780 -1880 9832 -1861
rect 11868 -1880 11904 -1861
rect 9780 -1915 11904 -1880
rect 9780 -1933 9832 -1915
rect 11868 -1933 11904 -1915
rect 9780 -2177 9822 -1933
rect 9864 -1969 11836 -1959
rect 9864 -2023 10131 -1969
rect 10711 -2023 11836 -1969
rect 9864 -2033 11836 -2023
rect 9864 -2087 11836 -2077
rect 9864 -2141 10988 -2087
rect 11568 -2141 11836 -2087
rect 9864 -2151 11836 -2141
rect 11894 -2177 11904 -1933
rect 9780 -2196 9832 -2177
rect 11868 -2196 11904 -2177
rect 9780 -2231 11904 -2196
rect 9780 -2249 9832 -2231
rect 11868 -2249 11904 -2231
rect 9780 -2493 9822 -2249
rect 9864 -2285 11836 -2275
rect 9864 -2339 10131 -2285
rect 10711 -2339 11836 -2285
rect 9864 -2349 11836 -2339
rect 9864 -2403 11836 -2393
rect 9864 -2457 10988 -2403
rect 11568 -2457 11836 -2403
rect 9864 -2467 11836 -2457
rect 11894 -2493 11904 -2249
rect 9780 -2512 9832 -2493
rect 11868 -2512 11904 -2493
rect 9780 -2547 11904 -2512
rect 9780 -2565 9832 -2547
rect 11868 -2565 11904 -2547
rect 9780 -2809 9822 -2565
rect 9864 -2601 11836 -2591
rect 9864 -2655 10131 -2601
rect 10711 -2655 11836 -2601
rect 9864 -2665 11836 -2655
rect 9864 -2719 11836 -2709
rect 9864 -2773 10988 -2719
rect 11568 -2773 11836 -2719
rect 9864 -2783 11836 -2773
rect 11894 -2809 11904 -2565
rect 9780 -2828 9832 -2809
rect 11868 -2828 11904 -2809
rect 9780 -2863 11904 -2828
rect 9780 -2881 9832 -2863
rect 11868 -2881 11904 -2863
rect 9780 -3125 9822 -2881
rect 9864 -2917 11836 -2907
rect 9864 -2971 10131 -2917
rect 10711 -2971 11836 -2917
rect 9864 -2981 11836 -2971
rect 9864 -3035 11836 -3025
rect 9864 -3089 10988 -3035
rect 11568 -3089 11836 -3035
rect 9864 -3099 11836 -3089
rect 11894 -3125 11904 -2881
rect 9780 -3144 9832 -3125
rect 11868 -3144 11904 -3125
rect 9780 -3179 11904 -3144
rect 9780 -3197 9832 -3179
rect 11868 -3197 11904 -3179
rect 9780 -3441 9822 -3197
rect 9864 -3233 11836 -3223
rect 9864 -3287 10131 -3233
rect 10711 -3287 11836 -3233
rect 9864 -3297 11836 -3287
rect 9864 -3351 11836 -3341
rect 9864 -3405 10988 -3351
rect 11568 -3405 11836 -3351
rect 9864 -3415 11836 -3405
rect 11894 -3441 11904 -3197
rect 9780 -3460 9832 -3441
rect 11868 -3460 11904 -3441
rect 9780 -3495 11904 -3460
rect 9780 -3513 9832 -3495
rect 11868 -3513 11904 -3495
rect 9780 -3757 9822 -3513
rect 9864 -3549 11836 -3539
rect 9864 -3603 10131 -3549
rect 10711 -3603 11836 -3549
rect 9864 -3613 11836 -3603
rect 9864 -3667 11836 -3657
rect 9864 -3721 10988 -3667
rect 11568 -3721 11836 -3667
rect 9864 -3731 11836 -3721
rect 11894 -3757 11904 -3513
rect 9780 -3776 9832 -3757
rect 11868 -3776 11904 -3757
rect 9780 -3811 11904 -3776
rect 9780 -3829 9832 -3811
rect 11868 -3829 11904 -3811
rect 9780 -4073 9822 -3829
rect 9864 -3865 11836 -3855
rect 9864 -3919 10131 -3865
rect 10711 -3919 11836 -3865
rect 9864 -3929 11836 -3919
rect 9864 -3983 11836 -3973
rect 9864 -4037 10988 -3983
rect 11568 -4037 11836 -3983
rect 9864 -4047 11836 -4037
rect 11894 -4073 11904 -3829
rect 9780 -4092 9832 -4073
rect 11868 -4092 11904 -4073
rect 9780 -4127 11904 -4092
rect 9780 -4145 9832 -4127
rect 11868 -4145 11904 -4127
rect 9780 -4389 9822 -4145
rect 9864 -4181 11836 -4171
rect 9864 -4235 10131 -4181
rect 10711 -4235 11836 -4181
rect 9864 -4245 11836 -4235
rect 9864 -4299 11836 -4289
rect 9864 -4353 10988 -4299
rect 11568 -4353 11836 -4299
rect 9864 -4363 11836 -4353
rect 11894 -4389 11904 -4145
rect 9780 -4408 9832 -4389
rect 11868 -4408 11904 -4389
rect 9780 -4443 11904 -4408
rect 9780 -4461 9832 -4443
rect 11868 -4461 11904 -4443
rect 9780 -4705 9822 -4461
rect 9864 -4497 11836 -4487
rect 9864 -4551 10131 -4497
rect 10711 -4551 11836 -4497
rect 9864 -4561 11836 -4551
rect 9864 -4615 11836 -4605
rect 9864 -4669 10988 -4615
rect 11568 -4669 11836 -4615
rect 9864 -4679 11836 -4669
rect 11894 -4705 11904 -4461
rect 9780 -4724 9832 -4705
rect 11868 -4724 11904 -4705
rect 9780 -4759 11904 -4724
rect 9780 -4777 9832 -4759
rect 11868 -4777 11904 -4759
rect 9780 -5021 9822 -4777
rect 9864 -4813 11836 -4803
rect 9864 -4867 10131 -4813
rect 10711 -4867 11836 -4813
rect 9864 -4877 11836 -4867
rect 9864 -4931 11836 -4921
rect 9864 -4985 10988 -4931
rect 11568 -4985 11836 -4931
rect 9864 -4995 11836 -4985
rect 11894 -5021 11904 -4777
rect 9780 -5040 9832 -5021
rect 11868 -5040 11904 -5021
rect 9780 -5075 11904 -5040
rect 9780 -5093 9832 -5075
rect 11868 -5093 11904 -5075
rect 9780 -5337 9822 -5093
rect 9864 -5129 11836 -5119
rect 9864 -5183 10131 -5129
rect 10711 -5183 11836 -5129
rect 9864 -5193 11836 -5183
rect 9864 -5247 11836 -5237
rect 9864 -5301 10988 -5247
rect 11568 -5301 11836 -5247
rect 9864 -5311 11836 -5301
rect 11894 -5337 11904 -5093
rect 9780 -5356 9832 -5337
rect 11868 -5356 11904 -5337
rect 9780 -5391 11904 -5356
rect 9780 -5409 9832 -5391
rect 11868 -5409 11904 -5391
rect 9780 -5653 9822 -5409
rect 9864 -5445 11836 -5435
rect 9864 -5499 10131 -5445
rect 10711 -5499 11836 -5445
rect 9864 -5509 11836 -5499
rect 9864 -5563 11836 -5553
rect 9864 -5617 10988 -5563
rect 11568 -5617 11836 -5563
rect 9864 -5627 11836 -5617
rect 11894 -5653 11904 -5409
rect 9780 -5672 9832 -5653
rect 11868 -5672 11904 -5653
rect 9780 -5707 11904 -5672
rect 9780 -5725 9832 -5707
rect 11868 -5725 11904 -5707
rect 9780 -5969 9822 -5725
rect 9864 -5761 11836 -5751
rect 9864 -5815 10131 -5761
rect 10711 -5815 11836 -5761
rect 9864 -5825 11836 -5815
rect 9864 -5879 11836 -5869
rect 9864 -5933 10988 -5879
rect 11568 -5933 11836 -5879
rect 9864 -5943 11836 -5933
rect 11894 -5969 11904 -5725
rect 9780 -5988 9832 -5969
rect 11868 -5988 11904 -5969
rect 9780 -6023 11904 -5988
rect 9780 -6041 9832 -6023
rect 11868 -6041 11904 -6023
rect 9780 -6285 9822 -6041
rect 9864 -6077 11836 -6067
rect 9864 -6131 10131 -6077
rect 10711 -6131 11836 -6077
rect 9864 -6141 11836 -6131
rect 9864 -6195 11836 -6185
rect 9864 -6249 10988 -6195
rect 11568 -6249 11836 -6195
rect 9864 -6259 11836 -6249
rect 11894 -6285 11904 -6041
rect 9780 -6304 9832 -6285
rect 11868 -6304 11904 -6285
rect 9780 -6339 11904 -6304
rect 9780 -6357 9832 -6339
rect 11868 -6357 11904 -6339
rect 9780 -6601 9822 -6357
rect 9864 -6393 11836 -6383
rect 9864 -6447 10131 -6393
rect 10711 -6447 11836 -6393
rect 9864 -6457 11836 -6447
rect 9864 -6511 11836 -6501
rect 9864 -6565 10988 -6511
rect 11568 -6565 11836 -6511
rect 9864 -6575 11836 -6565
rect 11894 -6601 11904 -6357
rect 9780 -6620 9832 -6601
rect 11868 -6620 11904 -6601
rect 9780 -6655 11904 -6620
rect 9780 -6673 9832 -6655
rect 11868 -6673 11904 -6655
rect 9780 -6917 9822 -6673
rect 9864 -6709 11836 -6699
rect 9864 -6763 10131 -6709
rect 10711 -6763 11836 -6709
rect 9864 -6773 11836 -6763
rect 9864 -6827 11836 -6817
rect 9864 -6881 10988 -6827
rect 11568 -6881 11836 -6827
rect 9864 -6891 11836 -6881
rect 11894 -6917 11904 -6673
rect 9780 -6936 9832 -6917
rect 11868 -6936 11904 -6917
rect 9780 -6971 11904 -6936
rect 9780 -6989 9832 -6971
rect 11868 -6989 11904 -6971
rect 9780 -7233 9822 -6989
rect 9864 -7025 11836 -7015
rect 9864 -7079 10131 -7025
rect 10711 -7079 11836 -7025
rect 9864 -7089 11836 -7079
rect 9864 -7143 11836 -7133
rect 9864 -7197 10988 -7143
rect 11568 -7197 11836 -7143
rect 9864 -7207 11836 -7197
rect 11894 -7233 11904 -6989
rect 9780 -7252 9832 -7233
rect 11868 -7252 11904 -7233
rect 9780 -7287 11904 -7252
rect 9780 -7305 9832 -7287
rect 11868 -7305 11904 -7287
rect 9780 -7549 9822 -7305
rect 9864 -7341 11836 -7331
rect 9864 -7395 10131 -7341
rect 10711 -7395 11836 -7341
rect 9864 -7405 11836 -7395
rect 9864 -7459 11836 -7449
rect 9864 -7513 10988 -7459
rect 11568 -7513 11836 -7459
rect 9864 -7523 11836 -7513
rect 11894 -7549 11904 -7305
rect 9780 -7568 9832 -7549
rect 11868 -7568 11904 -7549
rect 9780 -7603 11904 -7568
rect 9780 -7621 9832 -7603
rect 11868 -7621 11904 -7603
rect 9780 -7865 9822 -7621
rect 9864 -7657 11836 -7647
rect 9864 -7711 10131 -7657
rect 10711 -7711 11836 -7657
rect 9864 -7721 11836 -7711
rect 9864 -7775 11836 -7765
rect 9864 -7829 10988 -7775
rect 11568 -7829 11836 -7775
rect 9864 -7839 11836 -7829
rect 11894 -7865 11904 -7621
rect 9780 -7884 9832 -7865
rect 11868 -7884 11904 -7865
rect 9780 -7919 11904 -7884
rect 9780 -7937 9832 -7919
rect 11868 -7937 11904 -7919
rect 9780 -8037 9822 -7937
rect 11894 -7952 11904 -7937
rect 11980 -1861 11990 -1761
rect 12048 -1771 14020 -1761
rect 12048 -1825 12315 -1771
rect 12895 -1825 14020 -1771
rect 12048 -1835 14020 -1825
rect 14062 -1861 14104 -1761
rect 11980 -1880 12016 -1861
rect 14052 -1880 14104 -1861
rect 11980 -1914 14104 -1880
rect 11980 -1933 12016 -1914
rect 14052 -1933 14104 -1914
rect 11980 -2177 11990 -1933
rect 12048 -1969 14020 -1959
rect 12048 -2023 13172 -1969
rect 13752 -2023 14020 -1969
rect 12048 -2033 14020 -2023
rect 12048 -2087 14020 -2077
rect 12048 -2141 12315 -2087
rect 12895 -2141 14020 -2087
rect 12048 -2151 14020 -2141
rect 14062 -2177 14104 -1933
rect 11980 -2196 12016 -2177
rect 14052 -2196 14104 -2177
rect 11980 -2230 14104 -2196
rect 11980 -2249 12016 -2230
rect 14052 -2249 14104 -2230
rect 11980 -2493 11990 -2249
rect 12048 -2285 14020 -2275
rect 12048 -2339 13172 -2285
rect 13752 -2339 14020 -2285
rect 12048 -2349 14020 -2339
rect 12048 -2403 14020 -2393
rect 12048 -2457 12315 -2403
rect 12895 -2457 14020 -2403
rect 12048 -2467 14020 -2457
rect 14062 -2493 14104 -2249
rect 11980 -2512 12016 -2493
rect 14052 -2512 14104 -2493
rect 11980 -2546 14104 -2512
rect 11980 -2565 12016 -2546
rect 14052 -2565 14104 -2546
rect 11980 -2809 11990 -2565
rect 12048 -2601 14020 -2591
rect 12048 -2655 13172 -2601
rect 13752 -2655 14020 -2601
rect 12048 -2665 14020 -2655
rect 12048 -2719 14020 -2709
rect 12048 -2773 12315 -2719
rect 12895 -2773 14020 -2719
rect 12048 -2783 14020 -2773
rect 14062 -2809 14104 -2565
rect 11980 -2828 12016 -2809
rect 14052 -2828 14104 -2809
rect 11980 -2862 14104 -2828
rect 11980 -2881 12016 -2862
rect 14052 -2881 14104 -2862
rect 11980 -3125 11990 -2881
rect 12048 -2917 14020 -2907
rect 12048 -2971 13172 -2917
rect 13752 -2971 14020 -2917
rect 12048 -2981 14020 -2971
rect 12048 -3035 14020 -3025
rect 12048 -3089 12315 -3035
rect 12895 -3089 14020 -3035
rect 12048 -3099 14020 -3089
rect 14062 -3125 14104 -2881
rect 11980 -3144 12016 -3125
rect 14052 -3144 14104 -3125
rect 11980 -3178 14104 -3144
rect 11980 -3197 12016 -3178
rect 14052 -3197 14104 -3178
rect 11980 -3441 11990 -3197
rect 12048 -3233 14020 -3223
rect 12048 -3287 13172 -3233
rect 13752 -3287 14020 -3233
rect 12048 -3297 14020 -3287
rect 12048 -3351 14020 -3341
rect 12048 -3405 12315 -3351
rect 12895 -3405 14020 -3351
rect 12048 -3415 14020 -3405
rect 14062 -3441 14104 -3197
rect 11980 -3460 12016 -3441
rect 14052 -3460 14104 -3441
rect 11980 -3494 14104 -3460
rect 11980 -3513 12016 -3494
rect 14052 -3513 14104 -3494
rect 11980 -3757 11990 -3513
rect 12048 -3549 14020 -3539
rect 12048 -3603 13172 -3549
rect 13752 -3603 14020 -3549
rect 12048 -3613 14020 -3603
rect 12048 -3667 14020 -3657
rect 12048 -3721 12315 -3667
rect 12895 -3721 14020 -3667
rect 12048 -3731 14020 -3721
rect 14062 -3757 14104 -3513
rect 11980 -3776 12016 -3757
rect 14052 -3776 14104 -3757
rect 11980 -3810 14104 -3776
rect 11980 -3829 12016 -3810
rect 14052 -3829 14104 -3810
rect 11980 -4073 11990 -3829
rect 12048 -3865 14020 -3855
rect 12048 -3919 13172 -3865
rect 13752 -3919 14020 -3865
rect 12048 -3929 14020 -3919
rect 12048 -3983 14020 -3973
rect 12048 -4037 12315 -3983
rect 12895 -4037 14020 -3983
rect 12048 -4047 14020 -4037
rect 14062 -4073 14104 -3829
rect 11980 -4092 12016 -4073
rect 14052 -4092 14104 -4073
rect 11980 -4126 14104 -4092
rect 11980 -4145 12016 -4126
rect 14052 -4145 14104 -4126
rect 11980 -4389 11990 -4145
rect 12048 -4181 14020 -4171
rect 12048 -4235 13172 -4181
rect 13752 -4235 14020 -4181
rect 12048 -4245 14020 -4235
rect 12048 -4299 14020 -4289
rect 12048 -4353 12315 -4299
rect 12895 -4353 14020 -4299
rect 12048 -4363 14020 -4353
rect 14062 -4389 14104 -4145
rect 11980 -4408 12016 -4389
rect 14052 -4408 14104 -4389
rect 11980 -4442 14104 -4408
rect 11980 -4461 12016 -4442
rect 14052 -4461 14104 -4442
rect 11980 -4705 11990 -4461
rect 12048 -4497 14020 -4487
rect 12048 -4551 13172 -4497
rect 13752 -4551 14020 -4497
rect 12048 -4561 14020 -4551
rect 12048 -4615 14020 -4605
rect 12048 -4669 12315 -4615
rect 12895 -4669 14020 -4615
rect 12048 -4679 14020 -4669
rect 14062 -4705 14104 -4461
rect 11980 -4724 12016 -4705
rect 14052 -4724 14104 -4705
rect 11980 -4758 14104 -4724
rect 11980 -4777 12016 -4758
rect 14052 -4777 14104 -4758
rect 11980 -5021 11990 -4777
rect 12048 -4813 14020 -4803
rect 12048 -4867 13172 -4813
rect 13752 -4867 14020 -4813
rect 12048 -4877 14020 -4867
rect 12048 -4931 14020 -4921
rect 12048 -4985 12315 -4931
rect 12895 -4985 14020 -4931
rect 12048 -4995 14020 -4985
rect 14062 -5021 14104 -4777
rect 11980 -5040 12016 -5021
rect 14052 -5040 14104 -5021
rect 11980 -5074 14104 -5040
rect 11980 -5093 12016 -5074
rect 14052 -5093 14104 -5074
rect 11980 -5337 11990 -5093
rect 12048 -5129 14020 -5119
rect 12048 -5183 13172 -5129
rect 13752 -5183 14020 -5129
rect 12048 -5193 14020 -5183
rect 12048 -5247 14020 -5237
rect 12048 -5301 12315 -5247
rect 12895 -5301 14020 -5247
rect 12048 -5311 14020 -5301
rect 14062 -5337 14104 -5093
rect 11980 -5356 12016 -5337
rect 14052 -5356 14104 -5337
rect 11980 -5390 14104 -5356
rect 11980 -5409 12016 -5390
rect 14052 -5409 14104 -5390
rect 11980 -5653 11990 -5409
rect 12048 -5445 14020 -5435
rect 12048 -5499 13172 -5445
rect 13752 -5499 14020 -5445
rect 12048 -5509 14020 -5499
rect 12048 -5563 14020 -5553
rect 12048 -5617 12315 -5563
rect 12895 -5617 14020 -5563
rect 12048 -5627 14020 -5617
rect 14062 -5653 14104 -5409
rect 11980 -5672 12016 -5653
rect 14052 -5672 14104 -5653
rect 11980 -5706 14104 -5672
rect 11980 -5725 12016 -5706
rect 14052 -5725 14104 -5706
rect 11980 -5969 11990 -5725
rect 12048 -5761 14020 -5751
rect 12048 -5815 13172 -5761
rect 13752 -5815 14020 -5761
rect 12048 -5825 14020 -5815
rect 12048 -5879 14020 -5869
rect 12048 -5933 12315 -5879
rect 12895 -5933 14020 -5879
rect 12048 -5943 14020 -5933
rect 14062 -5969 14104 -5725
rect 11980 -5988 12016 -5969
rect 14052 -5988 14104 -5969
rect 11980 -6022 14104 -5988
rect 11980 -6041 12016 -6022
rect 14052 -6041 14104 -6022
rect 11980 -6285 11990 -6041
rect 12048 -6077 14020 -6067
rect 12048 -6131 13172 -6077
rect 13752 -6131 14020 -6077
rect 12048 -6141 14020 -6131
rect 12048 -6195 14020 -6185
rect 12048 -6249 12315 -6195
rect 12895 -6249 14020 -6195
rect 12048 -6259 14020 -6249
rect 14062 -6285 14104 -6041
rect 11980 -6304 12016 -6285
rect 14052 -6304 14104 -6285
rect 11980 -6338 14104 -6304
rect 11980 -6357 12016 -6338
rect 14052 -6357 14104 -6338
rect 11980 -6601 11990 -6357
rect 12048 -6393 14020 -6383
rect 12048 -6447 13172 -6393
rect 13752 -6447 14020 -6393
rect 12048 -6457 14020 -6447
rect 12048 -6511 14020 -6501
rect 12048 -6565 12315 -6511
rect 12895 -6565 14020 -6511
rect 12048 -6575 14020 -6565
rect 14062 -6601 14104 -6357
rect 11980 -6620 12016 -6601
rect 14052 -6620 14104 -6601
rect 11980 -6654 14104 -6620
rect 11980 -6673 12016 -6654
rect 14052 -6673 14104 -6654
rect 11980 -6917 11990 -6673
rect 12048 -6709 14020 -6699
rect 12048 -6763 13172 -6709
rect 13752 -6763 14020 -6709
rect 12048 -6773 14020 -6763
rect 12048 -6827 14020 -6817
rect 12048 -6881 12315 -6827
rect 12895 -6881 14020 -6827
rect 12048 -6891 14020 -6881
rect 14062 -6917 14104 -6673
rect 11980 -6936 12016 -6917
rect 14052 -6936 14104 -6917
rect 11980 -6970 14104 -6936
rect 11980 -6989 12016 -6970
rect 14052 -6989 14104 -6970
rect 11980 -7233 11990 -6989
rect 12048 -7025 14020 -7015
rect 12048 -7079 13172 -7025
rect 13752 -7079 14020 -7025
rect 12048 -7089 14020 -7079
rect 12048 -7143 14020 -7133
rect 12048 -7197 12315 -7143
rect 12895 -7197 14020 -7143
rect 12048 -7207 14020 -7197
rect 14062 -7233 14104 -6989
rect 11980 -7252 12016 -7233
rect 14052 -7252 14104 -7233
rect 11980 -7286 14104 -7252
rect 11980 -7305 12016 -7286
rect 14052 -7305 14104 -7286
rect 11980 -7549 11990 -7305
rect 12048 -7341 14020 -7331
rect 12048 -7395 13172 -7341
rect 13752 -7395 14020 -7341
rect 12048 -7405 14020 -7395
rect 12048 -7459 14020 -7449
rect 12048 -7513 12315 -7459
rect 12895 -7513 14020 -7459
rect 12048 -7523 14020 -7513
rect 14062 -7549 14104 -7305
rect 11980 -7568 12016 -7549
rect 14052 -7568 14104 -7549
rect 11980 -7602 14104 -7568
rect 11980 -7621 12016 -7602
rect 14052 -7621 14104 -7602
rect 11980 -7865 11990 -7621
rect 12048 -7657 14020 -7647
rect 12048 -7711 13172 -7657
rect 13752 -7711 14020 -7657
rect 12048 -7721 14020 -7711
rect 12048 -7775 14020 -7765
rect 12048 -7829 12315 -7775
rect 12895 -7829 14020 -7775
rect 12048 -7839 14020 -7829
rect 14062 -7865 14104 -7621
rect 11980 -7884 12016 -7865
rect 14052 -7884 14104 -7865
rect 11980 -7918 14104 -7884
rect 11980 -7937 12016 -7918
rect 14052 -7937 14104 -7918
rect 11980 -7952 11990 -7937
rect 11894 -7963 11990 -7952
rect 9864 -7973 11836 -7963
rect 9864 -8027 10131 -7973
rect 10711 -8027 11836 -7973
rect 9864 -8037 11836 -8027
rect 12048 -7973 14020 -7963
rect 12048 -8027 13172 -7973
rect 13752 -8027 14020 -7973
rect 12048 -8037 14020 -8027
rect 14062 -8037 14104 -7937
rect 14160 -8182 15266 -1663
rect 9143 -8353 16281 -8343
rect 9143 -8526 9153 -8353
rect 9333 -8526 16281 -8353
rect 9143 -8536 16281 -8526
rect 3879 -9003 10849 -8762
rect 3879 -11344 4262 -9003
rect 4569 -9156 4941 -9104
rect 5205 -9156 5577 -9104
rect 6233 -9156 6605 -9104
rect 6869 -9156 7241 -9104
rect 4464 -11160 4543 -9188
rect 4705 -9722 4805 -9156
rect 4705 -9902 4715 -9722
rect 4795 -9902 4805 -9722
rect 4705 -10446 4805 -9902
rect 4705 -10625 4715 -10446
rect 4795 -10625 4805 -10446
rect 4464 -11344 4533 -11160
rect 4705 -11192 4805 -10625
rect 4967 -9722 5046 -9188
rect 4967 -9902 4977 -9722
rect 5036 -9902 5046 -9722
rect 4967 -11160 5046 -9902
rect 5100 -11160 5179 -9188
rect 5341 -9722 5441 -9156
rect 5341 -9902 5351 -9722
rect 5431 -9902 5441 -9722
rect 5341 -10446 5441 -9902
rect 5341 -10626 5351 -10446
rect 5431 -10626 5441 -10446
rect 4569 -11244 4941 -11192
rect 5100 -11344 5169 -11160
rect 5341 -11192 5441 -10626
rect 5603 -9722 5682 -9188
rect 5603 -9902 5613 -9722
rect 5672 -9902 5682 -9722
rect 5603 -11160 5682 -9902
rect 6128 -11160 6207 -9188
rect 6369 -10446 6469 -9156
rect 6369 -10626 6379 -10446
rect 6459 -10626 6469 -10446
rect 5205 -11244 5577 -11192
rect 6128 -11344 6197 -11160
rect 6369 -11192 6469 -10626
rect 6631 -9722 6710 -9188
rect 6631 -9902 6641 -9722
rect 6700 -9902 6710 -9722
rect 6631 -11160 6710 -9902
rect 6764 -11160 6843 -9188
rect 7005 -10446 7105 -9156
rect 7005 -10626 7015 -10446
rect 7095 -10626 7105 -10446
rect 6233 -11244 6605 -11192
rect 6764 -11344 6833 -11160
rect 7005 -11192 7105 -10626
rect 7267 -9722 7346 -9188
rect 7267 -9902 7277 -9722
rect 7336 -9902 7346 -9722
rect 7267 -11160 7346 -9902
rect 6869 -11244 7241 -11192
rect 7549 -11344 7824 -9003
rect 8054 -9091 8254 -9081
rect 8054 -9277 8064 -9091
rect 8244 -9277 8254 -9091
rect 8054 -11008 8254 -9277
rect 8054 -11194 8064 -11008
rect 8244 -11194 8254 -11008
rect 8054 -11204 8254 -11194
rect 8448 -11344 8723 -9003
rect 9028 -9156 9400 -9104
rect 9664 -9156 10036 -9104
rect 10300 -9156 10672 -9104
rect 10936 -9156 11308 -9104
rect 11572 -9156 11944 -9104
rect 12208 -9156 12580 -9104
rect 12844 -9156 13216 -9104
rect 13480 -9156 13852 -9104
rect 8923 -11160 9002 -9188
rect 9164 -10446 9264 -9156
rect 9164 -10626 9174 -10446
rect 9254 -10626 9264 -10446
rect 8923 -11344 8992 -11160
rect 9164 -11192 9264 -10626
rect 9426 -9722 9505 -9188
rect 9426 -9902 9436 -9722
rect 9495 -9902 9505 -9722
rect 9426 -11160 9505 -9902
rect 9559 -11160 9638 -9188
rect 9800 -10446 9900 -9156
rect 9800 -10626 9810 -10446
rect 9890 -10626 9900 -10446
rect 9028 -11244 9400 -11192
rect 9559 -11344 9628 -11160
rect 9800 -11192 9900 -10626
rect 10062 -9722 10141 -9188
rect 10062 -9902 10072 -9722
rect 10131 -9902 10141 -9722
rect 10062 -11160 10141 -9902
rect 10195 -11160 10274 -9188
rect 10436 -10446 10536 -9156
rect 10436 -10626 10446 -10446
rect 10526 -10626 10536 -10446
rect 9664 -11244 10036 -11192
rect 10195 -11344 10264 -11160
rect 10436 -11192 10536 -10626
rect 10698 -9722 10777 -9188
rect 10698 -9902 10708 -9722
rect 10767 -9902 10777 -9722
rect 10698 -11160 10777 -9902
rect 10831 -11160 10910 -9188
rect 11072 -10446 11172 -9156
rect 11072 -10626 11082 -10446
rect 11162 -10626 11172 -10446
rect 10300 -11244 10672 -11192
rect 10831 -11344 10900 -11160
rect 11072 -11192 11172 -10626
rect 11334 -9722 11413 -9188
rect 11334 -9902 11344 -9722
rect 11403 -9902 11413 -9722
rect 11334 -11160 11413 -9902
rect 11467 -11160 11546 -9188
rect 11708 -10446 11808 -9156
rect 11708 -10626 11718 -10446
rect 11798 -10626 11808 -10446
rect 10936 -11244 11308 -11192
rect 11467 -11344 11536 -11160
rect 11708 -11192 11808 -10626
rect 11970 -9722 12049 -9188
rect 11970 -9902 11980 -9722
rect 12039 -9902 12049 -9722
rect 11970 -11160 12049 -9902
rect 12103 -11160 12182 -9188
rect 12344 -10446 12444 -9156
rect 12344 -10626 12354 -10446
rect 12434 -10626 12444 -10446
rect 11572 -11244 11944 -11192
rect 12103 -11344 12172 -11160
rect 12344 -11192 12444 -10626
rect 12606 -9722 12685 -9188
rect 12606 -9902 12616 -9722
rect 12675 -9902 12685 -9722
rect 12606 -11160 12685 -9902
rect 12739 -11160 12818 -9188
rect 12980 -10446 13080 -9156
rect 12980 -10626 12990 -10446
rect 13070 -10626 13080 -10446
rect 12208 -11244 12580 -11192
rect 12739 -11344 12808 -11160
rect 12980 -11192 13080 -10626
rect 13242 -9722 13321 -9188
rect 13242 -9902 13252 -9722
rect 13311 -9902 13321 -9722
rect 13242 -11160 13321 -9902
rect 13375 -11160 13454 -9188
rect 13616 -10446 13716 -9156
rect 13616 -10626 13626 -10446
rect 13706 -10626 13716 -10446
rect 12844 -11244 13216 -11192
rect 13375 -11344 13444 -11160
rect 13616 -11192 13716 -10626
rect 13878 -9722 13957 -9188
rect 13878 -9902 13888 -9722
rect 13947 -9902 13957 -9722
rect 13878 -11160 13957 -9902
rect 13480 -11244 13852 -11192
rect 14159 -11344 14519 -9828
rect 14652 -9937 14844 -9927
rect 14652 -9994 14662 -9937
rect 14834 -9994 14844 -9937
rect 14652 -10060 14844 -9994
rect 3879 -11587 14519 -11344
rect 3368 -11679 4712 -11669
rect 3368 -11892 4398 -11679
rect 4702 -11892 4712 -11679
rect 3368 -11902 4712 -11892
rect 5563 -11696 14519 -11587
rect 5563 -14038 5785 -11696
rect 6092 -11851 6464 -11799
rect 6728 -11851 7100 -11799
rect 7756 -11851 8128 -11799
rect 8392 -11851 8764 -11799
rect 9028 -11851 9400 -11799
rect 9664 -11851 10036 -11799
rect 10300 -11851 10672 -11799
rect 10936 -11851 11308 -11799
rect 11572 -11851 11944 -11799
rect 12208 -11851 12580 -11799
rect 12844 -11851 13216 -11799
rect 13480 -11851 13852 -11799
rect 5987 -13855 6066 -11883
rect 6228 -12417 6328 -11851
rect 6228 -12597 6238 -12417
rect 6318 -12597 6328 -12417
rect 6228 -13140 6328 -12597
rect 6228 -13320 6238 -13140
rect 6318 -13320 6328 -13140
rect 5987 -14038 6056 -13855
rect 6228 -13887 6328 -13320
rect 6490 -12417 6569 -11883
rect 6490 -12597 6500 -12417
rect 6559 -12597 6569 -12417
rect 6490 -13855 6569 -12597
rect 6623 -13855 6702 -11883
rect 6864 -12417 6964 -11851
rect 6864 -12597 6874 -12417
rect 6954 -12597 6964 -12417
rect 6864 -13140 6964 -12597
rect 6864 -13320 6874 -13140
rect 6954 -13320 6964 -13140
rect 6092 -13939 6464 -13887
rect 6623 -14038 6692 -13855
rect 6864 -13887 6964 -13320
rect 7126 -12417 7205 -11883
rect 7126 -12597 7136 -12417
rect 7195 -12597 7205 -12417
rect 7126 -13855 7205 -12597
rect 7651 -13855 7730 -11883
rect 7892 -13140 7992 -11851
rect 7892 -13320 7902 -13140
rect 7982 -13320 7992 -13140
rect 6728 -13939 7100 -13887
rect 7651 -14037 7720 -13855
rect 7892 -13887 7992 -13320
rect 8154 -12416 8233 -11883
rect 8154 -12596 8164 -12416
rect 8223 -12596 8233 -12416
rect 8154 -13855 8233 -12596
rect 8287 -13855 8366 -11883
rect 8528 -13140 8628 -11851
rect 8528 -13320 8538 -13140
rect 8618 -13320 8628 -13140
rect 7756 -13939 8128 -13887
rect 8287 -14037 8356 -13855
rect 8528 -13887 8628 -13320
rect 8790 -12416 8869 -11883
rect 8790 -12596 8800 -12416
rect 8859 -12596 8869 -12416
rect 8790 -13855 8869 -12596
rect 8923 -13855 9002 -11883
rect 9164 -13140 9264 -11851
rect 9164 -13320 9174 -13140
rect 9254 -13320 9264 -13140
rect 8392 -13939 8764 -13887
rect 8923 -14037 8992 -13855
rect 9164 -13887 9264 -13320
rect 9426 -12416 9505 -11883
rect 9426 -12596 9436 -12416
rect 9495 -12596 9505 -12416
rect 9426 -13855 9505 -12596
rect 9559 -13855 9638 -11883
rect 9800 -13140 9900 -11851
rect 9800 -13320 9810 -13140
rect 9890 -13320 9900 -13140
rect 9028 -13939 9400 -13887
rect 9559 -14037 9628 -13855
rect 9800 -13887 9900 -13320
rect 10062 -12416 10141 -11883
rect 10062 -12596 10072 -12416
rect 10131 -12596 10141 -12416
rect 10062 -13855 10141 -12596
rect 10195 -13855 10274 -11883
rect 10436 -13140 10536 -11851
rect 10436 -13320 10446 -13140
rect 10526 -13320 10536 -13140
rect 9664 -13939 10036 -13887
rect 10195 -14037 10264 -13855
rect 10436 -13887 10536 -13320
rect 10698 -12416 10777 -11883
rect 10698 -12596 10708 -12416
rect 10767 -12596 10777 -12416
rect 10698 -13855 10777 -12596
rect 10831 -13855 10910 -11883
rect 11072 -13140 11172 -11851
rect 11072 -13320 11082 -13140
rect 11162 -13320 11172 -13140
rect 10300 -13939 10672 -13887
rect 10831 -14037 10900 -13855
rect 11072 -13887 11172 -13320
rect 11334 -12416 11413 -11883
rect 11334 -12596 11344 -12416
rect 11403 -12596 11413 -12416
rect 11334 -13855 11413 -12596
rect 11467 -13855 11546 -11883
rect 11708 -13140 11808 -11851
rect 11708 -13320 11718 -13140
rect 11798 -13320 11808 -13140
rect 10936 -13939 11308 -13887
rect 11467 -14037 11536 -13855
rect 11708 -13887 11808 -13320
rect 11970 -12416 12049 -11883
rect 11970 -12596 11980 -12416
rect 12039 -12596 12049 -12416
rect 11970 -13855 12049 -12596
rect 12103 -13855 12182 -11883
rect 12344 -13140 12444 -11851
rect 12344 -13320 12354 -13140
rect 12434 -13320 12444 -13140
rect 11572 -13939 11944 -13887
rect 12103 -14037 12172 -13855
rect 12344 -13887 12444 -13320
rect 12606 -12416 12685 -11883
rect 12606 -12596 12616 -12416
rect 12675 -12596 12685 -12416
rect 12606 -13855 12685 -12596
rect 12739 -13855 12818 -11883
rect 12980 -13140 13080 -11851
rect 12980 -13320 12990 -13140
rect 13070 -13320 13080 -13140
rect 12208 -13939 12580 -13887
rect 12739 -14037 12808 -13855
rect 12980 -13887 13080 -13320
rect 13242 -12416 13321 -11883
rect 13242 -12596 13252 -12416
rect 13311 -12596 13321 -12416
rect 13242 -13855 13321 -12596
rect 13375 -13855 13454 -11883
rect 13616 -13140 13716 -11851
rect 13616 -13320 13626 -13140
rect 13706 -13320 13716 -13140
rect 12844 -13939 13216 -13887
rect 13375 -14037 13444 -13855
rect 13616 -13887 13716 -13320
rect 13878 -12416 13957 -11883
rect 13878 -12596 13888 -12416
rect 13947 -12596 13957 -12416
rect 13878 -13855 13957 -12596
rect 14159 -12423 14519 -11696
rect 14652 -12306 14844 -12240
rect 14652 -12369 14662 -12306
rect 14834 -12369 14844 -12306
rect 14652 -12379 14844 -12369
rect 14978 -12423 15266 -9828
rect 16088 -10239 16281 -8536
rect 15621 -10319 16797 -10239
rect 15621 -11210 15701 -10319
rect 16717 -11210 16797 -10319
rect 15621 -11290 16797 -11210
rect 13480 -13939 13852 -13887
rect 14159 -14037 15266 -12423
rect 7528 -14038 15266 -14037
rect 5563 -14980 15266 -14038
<< via1 >>
rect 3681 213 3761 393
rect 3943 -330 4005 -150
rect 4317 213 4397 393
rect 4579 -330 4641 -150
rect 5129 213 5209 393
rect 5129 -330 5209 -150
rect 5391 -330 5453 -150
rect 5765 213 5845 393
rect 5765 -330 5845 -150
rect 6027 -330 6089 -150
rect 6577 213 6657 393
rect 6577 -330 6657 -150
rect 6839 -330 6901 -150
rect 7213 213 7293 393
rect 7213 -330 7293 -150
rect 7475 -330 7537 -150
rect 8025 213 8105 393
rect 8287 -330 8349 -150
rect 8661 213 8741 393
rect 8923 -330 8985 -150
rect 9297 213 9377 393
rect 9559 -330 9621 -150
rect 9933 213 10013 393
rect 10195 -330 10257 -150
rect 10569 213 10649 393
rect 10831 -330 10893 -150
rect 11205 213 11285 393
rect 11467 -330 11529 -150
rect 11841 213 11921 393
rect 12103 -330 12165 -150
rect 12477 213 12557 393
rect 12739 -330 12801 -150
rect 13113 213 13193 393
rect 13375 -330 13437 -150
rect 13749 213 13829 393
rect 14011 -330 14073 -150
rect 3378 -1673 3658 -1398
rect 5842 -1684 6022 -1620
rect 7052 -1684 7232 -1620
rect 4756 -1946 4936 -1866
rect 8138 -1946 8318 -1866
rect 5299 -2192 5479 -2128
rect 7595 -2192 7775 -2128
rect 5842 -2320 6022 -2256
rect 7052 -2320 7232 -2256
rect 4756 -2582 4936 -2502
rect 8138 -2582 8318 -2502
rect 5299 -2828 5479 -2764
rect 7595 -2828 7775 -2764
rect 5842 -2956 6022 -2892
rect 7052 -2956 7232 -2892
rect 4756 -3218 4936 -3138
rect 8138 -3218 8318 -3138
rect 5299 -3464 5479 -3400
rect 7595 -3464 7775 -3400
rect 5842 -3592 6022 -3528
rect 7052 -3592 7232 -3528
rect 4756 -3854 4936 -3774
rect 8138 -3854 8318 -3774
rect 5299 -4100 5479 -4036
rect 7595 -4100 7775 -4036
rect 5842 -4228 6022 -4164
rect 7052 -4228 7232 -4164
rect 4756 -4490 4936 -4410
rect 8138 -4490 8318 -4410
rect 5299 -4736 5479 -4672
rect 7595 -4736 7775 -4672
rect 5842 -4864 6022 -4800
rect 7052 -4864 7232 -4800
rect 4756 -5126 4936 -5046
rect 8138 -5126 8318 -5046
rect 5299 -5372 5479 -5308
rect 7595 -5372 7775 -5308
rect 5842 -5500 6022 -5436
rect 7052 -5500 7232 -5436
rect 4756 -5762 4936 -5682
rect 8138 -5762 8318 -5682
rect 5299 -6008 5479 -5944
rect 7595 -6008 7775 -5944
rect 5842 -6136 6022 -6072
rect 7052 -6136 7232 -6072
rect 4756 -6398 4936 -6318
rect 8138 -6398 8318 -6318
rect 5299 -6644 5479 -6580
rect 7595 -6644 7775 -6580
rect 5842 -6772 6022 -6708
rect 7052 -6772 7232 -6708
rect 4756 -7034 4936 -6954
rect 8138 -7034 8318 -6954
rect 5299 -7280 5479 -7216
rect 7595 -7280 7775 -7216
rect 5842 -7408 6022 -7344
rect 7052 -7408 7232 -7344
rect 4756 -7670 4936 -7590
rect 8138 -7670 8318 -7590
rect 5299 -7916 5479 -7852
rect 7595 -7916 7775 -7852
rect 6138 -8236 6318 -8140
rect 6138 -8681 6318 -8585
rect 10131 -1653 10711 -1242
rect 13172 -1653 13752 -1242
rect 10988 -1825 11568 -1771
rect 10131 -2023 10711 -1969
rect 10988 -2141 11568 -2087
rect 10131 -2339 10711 -2285
rect 10988 -2457 11568 -2403
rect 10131 -2655 10711 -2601
rect 10988 -2773 11568 -2719
rect 10131 -2971 10711 -2917
rect 10988 -3089 11568 -3035
rect 10131 -3287 10711 -3233
rect 10988 -3405 11568 -3351
rect 10131 -3603 10711 -3549
rect 10988 -3721 11568 -3667
rect 10131 -3919 10711 -3865
rect 10988 -4037 11568 -3983
rect 10131 -4235 10711 -4181
rect 10988 -4353 11568 -4299
rect 10131 -4551 10711 -4497
rect 10988 -4669 11568 -4615
rect 10131 -4867 10711 -4813
rect 10988 -4985 11568 -4931
rect 10131 -5183 10711 -5129
rect 10988 -5301 11568 -5247
rect 10131 -5499 10711 -5445
rect 10988 -5617 11568 -5563
rect 10131 -5815 10711 -5761
rect 10988 -5933 11568 -5879
rect 10131 -6131 10711 -6077
rect 10988 -6249 11568 -6195
rect 10131 -6447 10711 -6393
rect 10988 -6565 11568 -6511
rect 10131 -6763 10711 -6709
rect 10988 -6881 11568 -6827
rect 10131 -7079 10711 -7025
rect 10988 -7197 11568 -7143
rect 10131 -7395 10711 -7341
rect 10988 -7513 11568 -7459
rect 10131 -7711 10711 -7657
rect 10988 -7829 11568 -7775
rect 11904 -7952 11980 -1761
rect 12315 -1825 12895 -1771
rect 13172 -2023 13752 -1969
rect 12315 -2141 12895 -2087
rect 13172 -2339 13752 -2285
rect 12315 -2457 12895 -2403
rect 13172 -2655 13752 -2601
rect 12315 -2773 12895 -2719
rect 13172 -2971 13752 -2917
rect 12315 -3089 12895 -3035
rect 13172 -3287 13752 -3233
rect 12315 -3405 12895 -3351
rect 13172 -3603 13752 -3549
rect 12315 -3721 12895 -3667
rect 13172 -3919 13752 -3865
rect 12315 -4037 12895 -3983
rect 13172 -4235 13752 -4181
rect 12315 -4353 12895 -4299
rect 13172 -4551 13752 -4497
rect 12315 -4669 12895 -4615
rect 13172 -4867 13752 -4813
rect 12315 -4985 12895 -4931
rect 13172 -5183 13752 -5129
rect 12315 -5301 12895 -5247
rect 13172 -5499 13752 -5445
rect 12315 -5617 12895 -5563
rect 13172 -5815 13752 -5761
rect 12315 -5933 12895 -5879
rect 13172 -6131 13752 -6077
rect 12315 -6249 12895 -6195
rect 13172 -6447 13752 -6393
rect 12315 -6565 12895 -6511
rect 13172 -6763 13752 -6709
rect 12315 -6881 12895 -6827
rect 13172 -7079 13752 -7025
rect 12315 -7197 12895 -7143
rect 13172 -7395 13752 -7341
rect 12315 -7513 12895 -7459
rect 13172 -7711 13752 -7657
rect 12315 -7829 12895 -7775
rect 10131 -8027 10711 -7973
rect 13172 -8027 13752 -7973
rect 9153 -8526 9333 -8353
rect 4715 -9902 4795 -9722
rect 4715 -10625 4795 -10446
rect 4977 -9902 5036 -9722
rect 5351 -9902 5431 -9722
rect 5351 -10626 5431 -10446
rect 5613 -9902 5672 -9722
rect 6379 -10626 6459 -10446
rect 6641 -9902 6700 -9722
rect 7015 -10626 7095 -10446
rect 7277 -9902 7336 -9722
rect 8064 -9277 8244 -9091
rect 8064 -11194 8244 -11008
rect 9174 -10626 9254 -10446
rect 9436 -9902 9495 -9722
rect 9810 -10626 9890 -10446
rect 10072 -9902 10131 -9722
rect 10446 -10626 10526 -10446
rect 10708 -9902 10767 -9722
rect 11082 -10626 11162 -10446
rect 11344 -9902 11403 -9722
rect 11718 -10626 11798 -10446
rect 11980 -9902 12039 -9722
rect 12354 -10626 12434 -10446
rect 12616 -9902 12675 -9722
rect 12990 -10626 13070 -10446
rect 13252 -9902 13311 -9722
rect 13626 -10626 13706 -10446
rect 13888 -9902 13947 -9722
rect 14662 -9994 14834 -9937
rect 4398 -11892 4702 -11679
rect 6238 -12597 6318 -12417
rect 6238 -13320 6318 -13140
rect 6500 -12597 6559 -12417
rect 6874 -12597 6954 -12417
rect 6874 -13320 6954 -13140
rect 7136 -12597 7195 -12417
rect 7902 -13320 7982 -13140
rect 8164 -12596 8223 -12416
rect 8538 -13320 8618 -13140
rect 8800 -12596 8859 -12416
rect 9174 -13320 9254 -13140
rect 9436 -12596 9495 -12416
rect 9810 -13320 9890 -13140
rect 10072 -12596 10131 -12416
rect 10446 -13320 10526 -13140
rect 10708 -12596 10767 -12416
rect 11082 -13320 11162 -13140
rect 11344 -12596 11403 -12416
rect 11718 -13320 11798 -13140
rect 11980 -12596 12039 -12416
rect 12354 -13320 12434 -13140
rect 12616 -12596 12675 -12416
rect 12990 -13320 13070 -13140
rect 13252 -12596 13311 -12416
rect 13626 -13320 13706 -13140
rect 13888 -12596 13947 -12416
rect 14662 -12369 14834 -12306
rect 15701 -11210 16717 -10319
<< metal2 >>
rect 3427 393 6099 403
rect 3427 213 3681 393
rect 3761 213 4317 393
rect 4397 213 5129 393
rect 5209 213 5765 393
rect 5845 213 6099 393
rect 3427 203 6099 213
rect 6323 393 14083 403
rect 6323 213 6577 393
rect 6657 213 7213 393
rect 7293 213 8025 393
rect 8105 213 8661 393
rect 8741 213 9297 393
rect 9377 213 9933 393
rect 10013 213 10569 393
rect 10649 213 11205 393
rect 11285 213 11841 393
rect 11921 213 12477 393
rect 12557 213 13113 393
rect 13193 213 13749 393
rect 13829 213 14083 393
rect 6323 203 14083 213
rect 3427 -150 4651 -140
rect 3427 -330 3943 -150
rect 4005 -330 4579 -150
rect 4641 -330 4651 -150
rect 3427 -340 4651 -330
rect 4875 -150 6099 -140
rect 4875 -330 5129 -150
rect 5209 -330 5391 -150
rect 5453 -330 5765 -150
rect 5845 -330 6027 -150
rect 6089 -330 6099 -150
rect 4875 -340 6099 -330
rect 6323 -150 7547 -140
rect 6323 -330 6577 -150
rect 6657 -330 6839 -150
rect 6901 -330 7213 -150
rect 7293 -330 7475 -150
rect 7537 -330 7547 -150
rect 6323 -340 7547 -330
rect 7771 -150 14083 -140
rect 7771 -330 8287 -150
rect 8349 -330 8923 -150
rect 8985 -330 9559 -150
rect 9621 -330 10195 -150
rect 10257 -330 10831 -150
rect 10893 -330 11467 -150
rect 11529 -330 12103 -150
rect 12165 -330 12739 -150
rect 12801 -330 13375 -150
rect 13437 -330 14011 -150
rect 14073 -330 14083 -150
rect 7771 -340 14083 -330
rect 3989 -1053 4089 -340
rect 5437 -954 5537 -340
rect 3368 -1153 4089 -1053
rect 5289 -1051 5537 -954
rect 6885 -953 6985 -340
rect 6885 -1049 7785 -953
rect 3368 -1398 3668 -1153
rect 3368 -1673 3378 -1398
rect 3658 -1673 3668 -1398
rect 3368 -1683 3668 -1673
rect 4746 -1866 4946 -1610
rect 4746 -1946 4756 -1866
rect 4936 -1946 4946 -1866
rect 4746 -2502 4946 -1946
rect 4746 -2582 4756 -2502
rect 4936 -2582 4946 -2502
rect 4746 -3138 4946 -2582
rect 4746 -3218 4756 -3138
rect 4936 -3218 4946 -3138
rect 4746 -3774 4946 -3218
rect 4746 -3854 4756 -3774
rect 4936 -3854 4946 -3774
rect 4746 -4410 4946 -3854
rect 4746 -4490 4756 -4410
rect 4936 -4490 4946 -4410
rect 4746 -5046 4946 -4490
rect 4746 -5126 4756 -5046
rect 4936 -5126 4946 -5046
rect 4746 -5682 4946 -5126
rect 4746 -5762 4756 -5682
rect 4936 -5762 4946 -5682
rect 4746 -6318 4946 -5762
rect 4746 -6398 4756 -6318
rect 4936 -6398 4946 -6318
rect 4746 -6954 4946 -6398
rect 4746 -7034 4756 -6954
rect 4936 -7034 4946 -6954
rect 4746 -7590 4946 -7034
rect 4746 -7670 4756 -7590
rect 4936 -7670 4946 -7590
rect 3163 -8142 3587 -7832
rect 4746 -8142 4946 -7670
rect 5289 -2128 5489 -1051
rect 5289 -2192 5299 -2128
rect 5479 -2192 5489 -2128
rect 5289 -2764 5489 -2192
rect 5289 -2828 5299 -2764
rect 5479 -2828 5489 -2764
rect 5289 -3400 5489 -2828
rect 5289 -3464 5299 -3400
rect 5479 -3464 5489 -3400
rect 5289 -4036 5489 -3464
rect 5289 -4100 5299 -4036
rect 5479 -4100 5489 -4036
rect 5289 -4672 5489 -4100
rect 5289 -4736 5299 -4672
rect 5479 -4736 5489 -4672
rect 5289 -5308 5489 -4736
rect 5289 -5372 5299 -5308
rect 5479 -5372 5489 -5308
rect 5289 -5944 5489 -5372
rect 5289 -6008 5299 -5944
rect 5479 -6008 5489 -5944
rect 5289 -6580 5489 -6008
rect 5289 -6644 5299 -6580
rect 5479 -6644 5489 -6580
rect 5289 -7216 5489 -6644
rect 5289 -7280 5299 -7216
rect 5479 -7280 5489 -7216
rect 5289 -7852 5489 -7280
rect 5289 -7916 5299 -7852
rect 5479 -7916 5489 -7852
rect 5289 -7926 5489 -7916
rect 5832 -1620 6032 -1610
rect 5832 -1684 5842 -1620
rect 6022 -1684 6032 -1620
rect 5832 -2256 6032 -1684
rect 5832 -2320 5842 -2256
rect 6022 -2320 6032 -2256
rect 5832 -2892 6032 -2320
rect 5832 -2956 5842 -2892
rect 6022 -2956 6032 -2892
rect 5832 -3528 6032 -2956
rect 5832 -3592 5842 -3528
rect 6022 -3592 6032 -3528
rect 5832 -4164 6032 -3592
rect 5832 -4228 5842 -4164
rect 6022 -4228 6032 -4164
rect 5832 -4800 6032 -4228
rect 5832 -4864 5842 -4800
rect 6022 -4864 6032 -4800
rect 5832 -5436 6032 -4864
rect 5832 -5500 5842 -5436
rect 6022 -5500 6032 -5436
rect 5832 -6072 6032 -5500
rect 5832 -6136 5842 -6072
rect 6022 -6136 6032 -6072
rect 5832 -6708 6032 -6136
rect 5832 -6772 5842 -6708
rect 6022 -6772 6032 -6708
rect 5832 -7344 6032 -6772
rect 5832 -7408 5842 -7344
rect 6022 -7408 6032 -7344
rect 5832 -7852 6032 -7408
rect 7042 -1620 7242 -1610
rect 7042 -1684 7052 -1620
rect 7232 -1684 7242 -1620
rect 7042 -2256 7242 -1684
rect 7042 -2320 7052 -2256
rect 7232 -2320 7242 -2256
rect 7042 -2892 7242 -2320
rect 7042 -2956 7052 -2892
rect 7232 -2956 7242 -2892
rect 7042 -3528 7242 -2956
rect 7042 -3592 7052 -3528
rect 7232 -3592 7242 -3528
rect 7042 -4164 7242 -3592
rect 7042 -4228 7052 -4164
rect 7232 -4228 7242 -4164
rect 7042 -4800 7242 -4228
rect 7042 -4864 7052 -4800
rect 7232 -4864 7242 -4800
rect 7042 -5436 7242 -4864
rect 7042 -5500 7052 -5436
rect 7232 -5500 7242 -5436
rect 7042 -6072 7242 -5500
rect 7042 -6136 7052 -6072
rect 7232 -6136 7242 -6072
rect 7042 -6708 7242 -6136
rect 7042 -6772 7052 -6708
rect 7232 -6772 7242 -6708
rect 7042 -7344 7242 -6772
rect 7042 -7408 7052 -7344
rect 7232 -7408 7242 -7344
rect 7042 -7852 7242 -7408
rect 5832 -7975 7242 -7852
rect 7585 -2128 7785 -1049
rect 7585 -2192 7595 -2128
rect 7775 -2192 7785 -2128
rect 7585 -2764 7785 -2192
rect 7585 -2828 7595 -2764
rect 7775 -2828 7785 -2764
rect 7585 -3400 7785 -2828
rect 7585 -3464 7595 -3400
rect 7775 -3464 7785 -3400
rect 7585 -4036 7785 -3464
rect 7585 -4100 7595 -4036
rect 7775 -4100 7785 -4036
rect 7585 -4672 7785 -4100
rect 7585 -4736 7595 -4672
rect 7775 -4736 7785 -4672
rect 7585 -5308 7785 -4736
rect 7585 -5372 7595 -5308
rect 7775 -5372 7785 -5308
rect 7585 -5944 7785 -5372
rect 7585 -6008 7595 -5944
rect 7775 -6008 7785 -5944
rect 7585 -6580 7785 -6008
rect 7585 -6644 7595 -6580
rect 7775 -6644 7785 -6580
rect 7585 -7216 7785 -6644
rect 7585 -7280 7595 -7216
rect 7775 -7280 7785 -7216
rect 7585 -7852 7785 -7280
rect 7585 -7916 7595 -7852
rect 7775 -7916 7785 -7852
rect 7585 -7926 7785 -7916
rect 8128 -1866 8328 -1610
rect 8128 -1946 8138 -1866
rect 8318 -1946 8328 -1866
rect 8128 -2502 8328 -1946
rect 8128 -2582 8138 -2502
rect 8318 -2582 8328 -2502
rect 8128 -3138 8328 -2582
rect 8128 -3218 8138 -3138
rect 8318 -3218 8328 -3138
rect 8128 -3774 8328 -3218
rect 8128 -3854 8138 -3774
rect 8318 -3854 8328 -3774
rect 8128 -4410 8328 -3854
rect 8128 -4490 8138 -4410
rect 8318 -4490 8328 -4410
rect 8128 -5046 8328 -4490
rect 8128 -5126 8138 -5046
rect 8318 -5126 8328 -5046
rect 8128 -5682 8328 -5126
rect 8128 -5762 8138 -5682
rect 8318 -5762 8328 -5682
rect 8128 -6318 8328 -5762
rect 8128 -6398 8138 -6318
rect 8318 -6398 8328 -6318
rect 8128 -6954 8328 -6398
rect 8128 -7034 8138 -6954
rect 8318 -7034 8328 -6954
rect 8128 -7590 8328 -7034
rect 8128 -7670 8138 -7590
rect 8318 -7670 8328 -7590
rect 3163 -8260 4946 -8142
rect 6128 -8140 6328 -7975
rect 6128 -8236 6138 -8140
rect 6318 -8236 6328 -8140
rect 8128 -8142 8328 -7670
rect 6128 -8246 6328 -8236
rect 6873 -8260 8328 -8142
rect 6873 -8334 6991 -8260
rect 3163 -8452 6991 -8334
rect 9143 -8353 9343 -340
rect 10121 -1242 10721 -1232
rect 10121 -1653 10131 -1242
rect 10711 -1653 10721 -1242
rect 10121 -1969 10721 -1653
rect 11836 -1761 12048 -340
rect 13162 -1242 13762 -1232
rect 13162 -1653 13172 -1242
rect 13752 -1653 13762 -1242
rect 10121 -2023 10131 -1969
rect 10711 -2023 10721 -1969
rect 10121 -2285 10721 -2023
rect 10121 -2339 10131 -2285
rect 10711 -2339 10721 -2285
rect 10121 -2601 10721 -2339
rect 10121 -2655 10131 -2601
rect 10711 -2655 10721 -2601
rect 10121 -2917 10721 -2655
rect 10121 -2971 10131 -2917
rect 10711 -2971 10721 -2917
rect 10121 -3233 10721 -2971
rect 10121 -3287 10131 -3233
rect 10711 -3287 10721 -3233
rect 10121 -3549 10721 -3287
rect 10121 -3603 10131 -3549
rect 10711 -3603 10721 -3549
rect 10121 -3865 10721 -3603
rect 10121 -3919 10131 -3865
rect 10711 -3919 10721 -3865
rect 10121 -4181 10721 -3919
rect 10121 -4235 10131 -4181
rect 10711 -4235 10721 -4181
rect 10121 -4497 10721 -4235
rect 10121 -4551 10131 -4497
rect 10711 -4551 10721 -4497
rect 10121 -4813 10721 -4551
rect 10121 -4867 10131 -4813
rect 10711 -4867 10721 -4813
rect 10121 -5129 10721 -4867
rect 10121 -5183 10131 -5129
rect 10711 -5183 10721 -5129
rect 10121 -5445 10721 -5183
rect 10121 -5499 10131 -5445
rect 10711 -5499 10721 -5445
rect 10121 -5761 10721 -5499
rect 10121 -5815 10131 -5761
rect 10711 -5815 10721 -5761
rect 10121 -6077 10721 -5815
rect 10121 -6131 10131 -6077
rect 10711 -6131 10721 -6077
rect 10121 -6393 10721 -6131
rect 10121 -6447 10131 -6393
rect 10711 -6447 10721 -6393
rect 10121 -6709 10721 -6447
rect 10121 -6763 10131 -6709
rect 10711 -6763 10721 -6709
rect 10121 -7025 10721 -6763
rect 10121 -7079 10131 -7025
rect 10711 -7079 10721 -7025
rect 10121 -7341 10721 -7079
rect 10121 -7395 10131 -7341
rect 10711 -7395 10721 -7341
rect 10121 -7657 10721 -7395
rect 10121 -7711 10131 -7657
rect 10711 -7711 10721 -7657
rect 10121 -7973 10721 -7711
rect 10121 -8027 10131 -7973
rect 10711 -8027 10721 -7973
rect 10121 -8037 10721 -8027
rect 10978 -1771 11578 -1761
rect 10978 -1825 10988 -1771
rect 11568 -1825 11578 -1771
rect 10978 -2087 11578 -1825
rect 10978 -2141 10988 -2087
rect 11568 -2141 11578 -2087
rect 10978 -2403 11578 -2141
rect 10978 -2457 10988 -2403
rect 11568 -2457 11578 -2403
rect 10978 -2719 11578 -2457
rect 10978 -2773 10988 -2719
rect 11568 -2773 11578 -2719
rect 10978 -3035 11578 -2773
rect 10978 -3089 10988 -3035
rect 11568 -3089 11578 -3035
rect 10978 -3351 11578 -3089
rect 10978 -3405 10988 -3351
rect 11568 -3405 11578 -3351
rect 10978 -3667 11578 -3405
rect 10978 -3721 10988 -3667
rect 11568 -3721 11578 -3667
rect 10978 -3983 11578 -3721
rect 10978 -4037 10988 -3983
rect 11568 -4037 11578 -3983
rect 10978 -4299 11578 -4037
rect 10978 -4353 10988 -4299
rect 11568 -4353 11578 -4299
rect 10978 -4615 11578 -4353
rect 10978 -4669 10988 -4615
rect 11568 -4669 11578 -4615
rect 10978 -4931 11578 -4669
rect 10978 -4985 10988 -4931
rect 11568 -4985 11578 -4931
rect 10978 -5247 11578 -4985
rect 10978 -5301 10988 -5247
rect 11568 -5301 11578 -5247
rect 10978 -5563 11578 -5301
rect 10978 -5617 10988 -5563
rect 11568 -5617 11578 -5563
rect 10978 -5879 11578 -5617
rect 10978 -5933 10988 -5879
rect 11568 -5933 11578 -5879
rect 10978 -6195 11578 -5933
rect 10978 -6249 10988 -6195
rect 11568 -6249 11578 -6195
rect 10978 -6511 11578 -6249
rect 10978 -6565 10988 -6511
rect 11568 -6565 11578 -6511
rect 10978 -6827 11578 -6565
rect 10978 -6881 10988 -6827
rect 11568 -6881 11578 -6827
rect 10978 -7143 11578 -6881
rect 10978 -7197 10988 -7143
rect 11568 -7197 11578 -7143
rect 10978 -7459 11578 -7197
rect 10978 -7513 10988 -7459
rect 11568 -7513 11578 -7459
rect 10978 -7775 11578 -7513
rect 10978 -7829 10988 -7775
rect 11568 -7829 11578 -7775
rect 10978 -8037 11578 -7829
rect 11836 -7952 11904 -1761
rect 11980 -7952 12048 -1761
rect 11836 -7963 12048 -7952
rect 12305 -1771 12905 -1761
rect 12305 -1825 12315 -1771
rect 12895 -1825 12905 -1771
rect 12305 -2087 12905 -1825
rect 12305 -2141 12315 -2087
rect 12895 -2141 12905 -2087
rect 12305 -2403 12905 -2141
rect 12305 -2457 12315 -2403
rect 12895 -2457 12905 -2403
rect 12305 -2719 12905 -2457
rect 12305 -2773 12315 -2719
rect 12895 -2773 12905 -2719
rect 12305 -3035 12905 -2773
rect 12305 -3089 12315 -3035
rect 12895 -3089 12905 -3035
rect 12305 -3351 12905 -3089
rect 12305 -3405 12315 -3351
rect 12895 -3405 12905 -3351
rect 12305 -3667 12905 -3405
rect 12305 -3721 12315 -3667
rect 12895 -3721 12905 -3667
rect 12305 -3983 12905 -3721
rect 12305 -4037 12315 -3983
rect 12895 -4037 12905 -3983
rect 12305 -4299 12905 -4037
rect 12305 -4353 12315 -4299
rect 12895 -4353 12905 -4299
rect 12305 -4615 12905 -4353
rect 12305 -4669 12315 -4615
rect 12895 -4669 12905 -4615
rect 12305 -4931 12905 -4669
rect 12305 -4985 12315 -4931
rect 12895 -4985 12905 -4931
rect 12305 -5247 12905 -4985
rect 12305 -5301 12315 -5247
rect 12895 -5301 12905 -5247
rect 12305 -5563 12905 -5301
rect 12305 -5617 12315 -5563
rect 12895 -5617 12905 -5563
rect 12305 -5879 12905 -5617
rect 12305 -5933 12315 -5879
rect 12895 -5933 12905 -5879
rect 12305 -6195 12905 -5933
rect 12305 -6249 12315 -6195
rect 12895 -6249 12905 -6195
rect 12305 -6511 12905 -6249
rect 12305 -6565 12315 -6511
rect 12895 -6565 12905 -6511
rect 12305 -6827 12905 -6565
rect 12305 -6881 12315 -6827
rect 12895 -6881 12905 -6827
rect 12305 -7143 12905 -6881
rect 12305 -7197 12315 -7143
rect 12895 -7197 12905 -7143
rect 12305 -7459 12905 -7197
rect 12305 -7513 12315 -7459
rect 12895 -7513 12905 -7459
rect 12305 -7775 12905 -7513
rect 12305 -7829 12315 -7775
rect 12895 -7829 12905 -7775
rect 12305 -8037 12905 -7829
rect 13162 -1969 13762 -1653
rect 13162 -2023 13172 -1969
rect 13752 -2023 13762 -1969
rect 13162 -2285 13762 -2023
rect 13162 -2339 13172 -2285
rect 13752 -2339 13762 -2285
rect 13162 -2601 13762 -2339
rect 13162 -2655 13172 -2601
rect 13752 -2655 13762 -2601
rect 13162 -2917 13762 -2655
rect 13162 -2971 13172 -2917
rect 13752 -2971 13762 -2917
rect 13162 -3233 13762 -2971
rect 13162 -3287 13172 -3233
rect 13752 -3287 13762 -3233
rect 13162 -3549 13762 -3287
rect 13162 -3603 13172 -3549
rect 13752 -3603 13762 -3549
rect 13162 -3865 13762 -3603
rect 13162 -3919 13172 -3865
rect 13752 -3919 13762 -3865
rect 13162 -4181 13762 -3919
rect 13162 -4235 13172 -4181
rect 13752 -4235 13762 -4181
rect 13162 -4497 13762 -4235
rect 13162 -4551 13172 -4497
rect 13752 -4551 13762 -4497
rect 13162 -4813 13762 -4551
rect 13162 -4867 13172 -4813
rect 13752 -4867 13762 -4813
rect 13162 -5129 13762 -4867
rect 13162 -5183 13172 -5129
rect 13752 -5183 13762 -5129
rect 13162 -5445 13762 -5183
rect 13162 -5499 13172 -5445
rect 13752 -5499 13762 -5445
rect 13162 -5761 13762 -5499
rect 13162 -5815 13172 -5761
rect 13752 -5815 13762 -5761
rect 13162 -6077 13762 -5815
rect 13162 -6131 13172 -6077
rect 13752 -6131 13762 -6077
rect 13162 -6393 13762 -6131
rect 13162 -6447 13172 -6393
rect 13752 -6447 13762 -6393
rect 13162 -6709 13762 -6447
rect 13162 -6763 13172 -6709
rect 13752 -6763 13762 -6709
rect 13162 -7025 13762 -6763
rect 13162 -7079 13172 -7025
rect 13752 -7079 13762 -7025
rect 13162 -7341 13762 -7079
rect 13162 -7395 13172 -7341
rect 13752 -7395 13762 -7341
rect 13162 -7657 13762 -7395
rect 13162 -7711 13172 -7657
rect 13752 -7711 13762 -7657
rect 13162 -7973 13762 -7711
rect 13162 -8027 13172 -7973
rect 13752 -8027 13762 -7973
rect 13162 -8037 13762 -8027
rect 3163 -8761 3587 -8452
rect 9143 -8526 9153 -8353
rect 9333 -8526 9343 -8353
rect 9143 -8536 9343 -8526
rect 6128 -8585 6328 -8575
rect 6128 -8681 6138 -8585
rect 6318 -8681 6328 -8585
rect 3163 -9712 3589 -9530
rect 6128 -9712 6328 -8681
rect 8054 -8736 9343 -8536
rect 10978 -8304 12905 -8037
rect 15408 -8304 16698 2104
rect 8054 -9091 8254 -8736
rect 8054 -9277 8064 -9091
rect 8244 -9277 8254 -9091
rect 8054 -9287 8254 -9277
rect 10978 -9712 16698 -8304
rect 3163 -9722 5682 -9712
rect 3163 -9902 4715 -9722
rect 4795 -9902 4977 -9722
rect 5036 -9902 5351 -9722
rect 5431 -9902 5613 -9722
rect 5672 -9902 5682 -9722
rect 3163 -9912 5682 -9902
rect 6128 -9722 7346 -9712
rect 6128 -9902 6641 -9722
rect 6700 -9902 7277 -9722
rect 7336 -9902 7346 -9722
rect 6128 -9912 7346 -9902
rect 7856 -9722 13957 -9712
rect 7856 -9902 9436 -9722
rect 9495 -9902 10072 -9722
rect 10131 -9902 10708 -9722
rect 10767 -9902 11344 -9722
rect 11403 -9902 11980 -9722
rect 12039 -9902 12616 -9722
rect 12675 -9902 13252 -9722
rect 13311 -9902 13888 -9722
rect 13947 -9902 13957 -9722
rect 7856 -9912 13957 -9902
rect 7856 -10083 8056 -9912
rect 14652 -9937 14844 -9712
rect 14652 -9994 14662 -9937
rect 14834 -9994 14844 -9937
rect 14652 -10004 14844 -9994
rect 3718 -10283 8056 -10083
rect 3718 -11976 3918 -10283
rect 15621 -10319 16797 -10239
rect 4464 -10446 13957 -10436
rect 4464 -10625 4715 -10446
rect 4795 -10625 5351 -10446
rect 4464 -10626 5351 -10625
rect 5431 -10626 6379 -10446
rect 6459 -10626 7015 -10446
rect 7095 -10626 9174 -10446
rect 9254 -10626 9810 -10446
rect 9890 -10626 10446 -10446
rect 10526 -10626 11082 -10446
rect 11162 -10626 11718 -10446
rect 11798 -10626 12354 -10446
rect 12434 -10626 12990 -10446
rect 13070 -10626 13626 -10446
rect 13706 -10626 13957 -10446
rect 4464 -10636 13957 -10626
rect 8054 -11008 8254 -10998
rect 8054 -11194 8064 -11008
rect 8244 -11194 8254 -11008
rect 4388 -11679 5846 -11669
rect 4388 -11892 4398 -11679
rect 4702 -11892 5846 -11679
rect 4388 -11902 5846 -11892
rect 5613 -12407 5846 -11902
rect 8054 -12406 8254 -11194
rect 15621 -11210 15701 -10319
rect 16717 -11210 16797 -10319
rect 15621 -11290 16797 -11210
rect 15611 -12040 16787 -11960
rect 15611 -12296 15691 -12040
rect 14652 -12306 15691 -12296
rect 14652 -12369 14662 -12306
rect 14834 -12369 15691 -12306
rect 5613 -12417 7205 -12407
rect 5613 -12597 6238 -12417
rect 6318 -12597 6500 -12417
rect 6559 -12597 6874 -12417
rect 6954 -12597 7136 -12417
rect 7195 -12597 7205 -12417
rect 5613 -12607 7205 -12597
rect 7651 -12416 13957 -12406
rect 7651 -12596 8164 -12416
rect 8223 -12596 8800 -12416
rect 8859 -12596 9436 -12416
rect 9495 -12596 10072 -12416
rect 10131 -12596 10708 -12416
rect 10767 -12596 11344 -12416
rect 11403 -12596 11980 -12416
rect 12039 -12596 12616 -12416
rect 12675 -12596 13252 -12416
rect 13311 -12596 13888 -12416
rect 13947 -12596 13957 -12416
rect 14652 -12454 15691 -12369
rect 7651 -12606 13957 -12596
rect 15611 -12931 15691 -12454
rect 16707 -12931 16787 -12040
rect 15611 -13011 16787 -12931
rect 5987 -13140 13957 -13130
rect 5987 -13320 6238 -13140
rect 6318 -13320 6874 -13140
rect 6954 -13320 7902 -13140
rect 7982 -13320 8538 -13140
rect 8618 -13320 9174 -13140
rect 9254 -13320 9810 -13140
rect 9890 -13320 10446 -13140
rect 10526 -13320 11082 -13140
rect 11162 -13320 11718 -13140
rect 11798 -13320 12354 -13140
rect 12434 -13320 12990 -13140
rect 13070 -13320 13626 -13140
rect 13706 -13320 13957 -13140
rect 5987 -13330 13957 -13320
<< via2 >>
rect 15701 -11210 16717 -10319
rect 15691 -12931 16707 -12040
<< metal3 >>
rect 15621 -10319 16797 -10239
rect 15621 -11210 15701 -10319
rect 16717 -11210 16797 -10319
rect 15621 -11290 16797 -11210
rect 15611 -12040 16787 -11960
rect 15611 -12931 15691 -12040
rect 16707 -12931 16787 -12040
rect 15611 -13011 16787 -12931
<< via3 >>
rect 15701 -11210 16717 -10319
rect 15691 -12931 16707 -12040
<< metal4 >>
rect 17171 -1089 22211 911
rect 22611 -1089 27651 911
rect 28051 -1089 33091 911
rect 17171 -2129 33091 -1089
rect 17171 -4129 22211 -2129
rect 22611 -4129 27651 -2129
rect 28051 -4129 33091 -2129
rect 19171 -4529 20211 -4129
rect 24611 -4529 25651 -4129
rect 30051 -4529 31091 -4129
rect 17171 -6529 22211 -4529
rect 22611 -6529 27651 -4529
rect 28051 -6529 33091 -4529
rect 17171 -7569 33091 -6529
rect 17171 -9569 22211 -7569
rect 22611 -9569 27651 -7569
rect 28051 -9569 33091 -7569
rect 19171 -9969 20211 -9569
rect 24611 -9969 25651 -9569
rect 30051 -9969 31091 -9569
rect 17171 -10239 22211 -9969
rect 15621 -10319 22211 -10239
rect 15621 -11210 15701 -10319
rect 16717 -11210 22211 -10319
rect 15621 -11290 22211 -11210
rect 15611 -12040 16787 -11960
rect 15611 -12931 15691 -12040
rect 16707 -12931 16787 -12040
rect 15611 -13011 16787 -12931
rect 17171 -11969 22211 -11290
rect 22611 -11969 27651 -9969
rect 28051 -11969 33091 -9969
rect 17171 -13009 33091 -11969
rect 17171 -15009 22211 -13009
rect 22611 -15009 27651 -13009
rect 28051 -15009 33091 -13009
<< via4 >>
rect 15691 -12931 16707 -12040
<< metal5 >>
rect 15611 -12040 16787 -11960
rect 15611 -12931 15691 -12040
rect 16707 -12931 16787 -12040
rect 15611 -13011 16787 -12931
<< via5 >>
rect 15691 -12931 16707 -12040
<< metal6 >>
rect 17171 -1089 22211 911
rect 22611 -1089 27651 911
rect 28051 -1089 33091 911
rect 17171 -2129 33091 -1089
rect 17171 -4129 22211 -2129
rect 22611 -4129 27651 -2129
rect 28051 -4129 33091 -2129
rect 19171 -4529 20211 -4129
rect 24611 -4529 25651 -4129
rect 30051 -4529 31091 -4129
rect 17171 -6529 22211 -4529
rect 22611 -6529 27651 -4529
rect 28051 -6529 33091 -4529
rect 17171 -7569 33091 -6529
rect 17171 -9569 22211 -7569
rect 22611 -9569 27651 -7569
rect 28051 -9569 33091 -7569
rect 19171 -9969 20211 -9569
rect 24611 -9969 25651 -9569
rect 30051 -9969 31091 -9569
rect 17171 -11960 22211 -9969
rect 15611 -11969 22211 -11960
rect 22611 -11969 27651 -9969
rect 28051 -11969 33091 -9969
rect 15611 -12040 33091 -11969
rect 15611 -12931 15691 -12040
rect 16707 -12931 33091 -12040
rect 15611 -13009 33091 -12931
rect 15611 -13011 22211 -13009
rect 17171 -15009 22211 -13011
rect 22611 -15009 27651 -13009
rect 28051 -15009 33091 -13009
use cmim_KCDMMN  cmim_KCDMMN_0
timestamp 1749416725
transform 1 0 19691 0 1 -12489
box -2520 -2520 13400 13400
use hvnmos_2L3HPE  hvnmos_2L3HPE_0
timestamp 1749416725
transform 1 0 7942 0 1 -12869
box -544 -1222 6268 1222
use hvnmos_2L3PPE  hvnmos_2L3PPE_0
timestamp 1749416725
transform 0 1 5389 -1 0 -1906
box -436 -1178 6160 1178
use hvnmos_2L3PPE  hvnmos_2L3PPE_1
timestamp 1749416725
transform 0 1 7685 -1 0 -1906
box -436 -1178 6160 1178
use hvnmos_8GE7KN  hvnmos_8GE7KN_0
timestamp 1749416725
transform 1 0 6419 0 1 -10174
box -544 -1222 1180 1222
use hvnmos_8GE7KN  hvnmos_8GE7KN_1
timestamp 1749416725
transform 1 0 6278 0 1 -12869
box -544 -1222 1180 1222
use hvnmos_8GE7KN  hvnmos_8GE7KN_2
timestamp 1749416725
transform 1 0 4755 0 1 -10174
box -544 -1222 1180 1222
use hvnmos_84A7KN  hvnmos_84A7KN_0
timestamp 1749416725
transform 1 0 9214 0 1 -10174
box -544 -1222 4996 1222
use hvpmos_2L3PPE  hvpmos_2L3PPE_0
timestamp 1749416725
transform -1 0 13789 0 -1 303
box -560 -1302 6284 1302
use hvpmos_5SRWXM  hvpmos_5SRWXM_0
timestamp 1749416725
transform 0 -1 13034 1 0 -7901
box -410 -1302 6414 3486
use hvpmos_8GEZJN  hvpmos_8GEZJN_0
timestamp 1749416725
transform -1 0 4357 0 -1 303
box -560 -1302 1196 1302
use hvpmos_8GEZJN  hvpmos_8GEZJN_1
timestamp 1749416725
transform -1 0 5805 0 -1 303
box -560 -1302 1196 1302
use hvpmos_8GEZJN  hvpmos_8GEZJN_2
timestamp 1749416725
transform -1 0 7253 0 -1 303
box -560 -1302 1196 1302
use rppd_PAUPFW  rppd_PAUPFW_0
timestamp 1749416725
transform 1 0 14748 0 1 -11150
box -280 -1326 280 1326
<< labels >>
flabel metal2 15408 1498 16698 2104 0 FreeSans 800 0 0 0 VOUT
port 0 nsew
flabel metal1 3163 1605 4719 2104 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal2 3163 -9912 3589 -9530 0 FreeSans 800 0 0 0 IB
port 3 nsew
flabel metal2 3163 -8761 3587 -8334 0 FreeSans 800 0 0 0 INN
port 4 nsew
flabel metal2 3163 -8260 3587 -7832 0 FreeSans 800 0 0 0 INP
port 5 nsew
flabel metal1 5563 -14980 7119 -14481 0 FreeSans 800 0 0 0 VSS
port 2 nsew
<< end >>
