magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 35 56 453 314
rect -26 -56 506 56
<< nmos >>
rect 129 140 155 288
rect 231 140 257 288
rect 333 140 359 288
<< pmos >>
rect 129 412 155 636
rect 231 412 257 636
rect 333 412 359 636
<< ndiff >>
rect 61 186 129 288
rect 61 154 75 186
rect 107 154 129 186
rect 61 140 129 154
rect 155 254 231 288
rect 155 222 177 254
rect 209 222 231 254
rect 155 186 231 222
rect 155 154 177 186
rect 209 154 231 186
rect 155 140 231 154
rect 257 140 333 288
rect 359 254 427 288
rect 359 222 381 254
rect 413 222 427 254
rect 359 186 427 222
rect 359 154 381 186
rect 413 154 427 186
rect 359 140 427 154
<< pdiff >>
rect 61 622 129 636
rect 61 590 75 622
rect 107 590 129 622
rect 61 554 129 590
rect 61 522 75 554
rect 107 522 129 554
rect 61 486 129 522
rect 61 454 75 486
rect 107 454 129 486
rect 61 412 129 454
rect 155 622 231 636
rect 155 590 177 622
rect 209 590 231 622
rect 155 554 231 590
rect 155 522 177 554
rect 209 522 231 554
rect 155 412 231 522
rect 257 622 333 636
rect 257 590 279 622
rect 311 590 333 622
rect 257 412 333 590
rect 359 622 427 636
rect 359 590 381 622
rect 413 590 427 622
rect 359 554 427 590
rect 359 522 381 554
rect 413 522 427 554
rect 359 486 427 522
rect 359 454 381 486
rect 413 454 427 486
rect 359 412 427 454
<< ndiffc >>
rect 75 154 107 186
rect 177 222 209 254
rect 177 154 209 186
rect 381 222 413 254
rect 381 154 413 186
<< pdiffc >>
rect 75 590 107 622
rect 75 522 107 554
rect 75 454 107 486
rect 177 590 209 622
rect 177 522 209 554
rect 279 590 311 622
rect 381 590 413 622
rect 381 522 413 554
rect 381 454 413 486
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 416 740 448 772
<< poly >>
rect 129 636 155 672
rect 231 636 257 672
rect 333 636 359 672
rect 129 380 155 412
rect 61 366 155 380
rect 61 334 75 366
rect 107 334 155 366
rect 61 320 155 334
rect 129 288 155 320
rect 231 380 257 412
rect 333 380 359 412
rect 231 366 291 380
rect 231 334 245 366
rect 277 334 291 366
rect 231 320 291 334
rect 333 366 427 380
rect 333 334 381 366
rect 413 334 427 366
rect 333 320 427 334
rect 231 288 257 320
rect 333 288 359 320
rect 129 104 155 140
rect 231 104 257 140
rect 333 104 359 140
<< polycont >>
rect 75 334 107 366
rect 245 334 277 366
rect 381 334 413 366
<< metal1 >>
rect 0 772 480 800
rect 0 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 65 622 124 632
rect 65 590 75 622
rect 107 590 124 622
rect 65 554 124 590
rect 65 522 75 554
rect 107 522 124 554
rect 65 486 124 522
rect 167 622 219 632
rect 167 590 177 622
rect 209 590 219 622
rect 167 554 219 590
rect 269 622 321 712
rect 269 590 279 622
rect 311 590 321 622
rect 269 580 321 590
rect 371 622 423 632
rect 371 590 381 622
rect 413 590 423 622
rect 167 522 177 554
rect 209 543 219 554
rect 371 554 423 590
rect 371 543 381 554
rect 209 522 381 543
rect 413 522 423 554
rect 167 511 423 522
rect 65 454 75 486
rect 107 458 124 486
rect 371 486 423 511
rect 107 454 199 458
rect 65 416 199 454
rect 371 454 381 486
rect 413 454 423 486
rect 371 416 423 454
rect 65 366 120 376
rect 65 334 75 366
rect 107 334 120 366
rect 65 269 120 334
rect 167 264 199 416
rect 235 366 316 376
rect 235 334 245 366
rect 277 334 316 366
rect 235 324 316 334
rect 264 269 316 324
rect 354 366 423 376
rect 354 334 381 366
rect 413 334 423 366
rect 354 300 423 334
rect 167 254 219 264
rect 167 222 177 254
rect 209 222 219 254
rect 65 186 117 196
rect 65 154 75 186
rect 107 154 117 186
rect 65 44 117 154
rect 167 186 219 222
rect 167 154 177 186
rect 209 154 219 186
rect 167 144 219 154
rect 371 254 423 264
rect 371 222 381 254
rect 413 222 423 254
rect 371 186 423 222
rect 371 154 381 186
rect 413 154 423 186
rect 371 44 423 154
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 354 300 423 376 0 FreeSans 400 0 0 0 A2
port 4 nsew
flabel metal1 s 264 269 316 376 0 FreeSans 400 0 0 0 A1
port 5 nsew
flabel metal1 s 65 269 120 376 0 FreeSans 400 0 0 0 B1
port 6 nsew
flabel metal1 s 65 416 124 632 0 FreeSans 400 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 159078
string GDS_FILE 6_final.gds
string GDS_START 155362
<< end >>
