magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 27 56 343 292
rect -26 -56 410 56
<< nmos >>
rect 121 118 147 266
rect 223 118 249 266
<< pmos >>
rect 121 412 147 636
rect 223 412 249 636
<< ndiff >>
rect 53 232 121 266
rect 53 200 67 232
rect 99 200 121 232
rect 53 164 121 200
rect 53 132 67 164
rect 99 132 121 164
rect 53 118 121 132
rect 147 232 223 266
rect 147 200 169 232
rect 201 200 223 232
rect 147 164 223 200
rect 147 132 169 164
rect 201 132 223 164
rect 147 118 223 132
rect 249 232 317 266
rect 249 200 271 232
rect 303 200 317 232
rect 249 164 317 200
rect 249 132 271 164
rect 303 132 317 164
rect 249 118 317 132
<< pdiff >>
rect 53 622 121 636
rect 53 590 67 622
rect 99 590 121 622
rect 53 554 121 590
rect 53 522 67 554
rect 99 522 121 554
rect 53 486 121 522
rect 53 454 67 486
rect 99 454 121 486
rect 53 412 121 454
rect 147 622 223 636
rect 147 590 169 622
rect 201 590 223 622
rect 147 554 223 590
rect 147 522 169 554
rect 201 522 223 554
rect 147 486 223 522
rect 147 454 169 486
rect 201 454 223 486
rect 147 412 223 454
rect 249 622 318 636
rect 249 590 272 622
rect 304 590 318 622
rect 249 554 318 590
rect 249 522 272 554
rect 304 522 318 554
rect 249 486 318 522
rect 249 454 272 486
rect 304 454 318 486
rect 249 412 318 454
<< ndiffc >>
rect 67 200 99 232
rect 67 132 99 164
rect 169 200 201 232
rect 169 132 201 164
rect 271 200 303 232
rect 271 132 303 164
<< pdiffc >>
rect 67 590 99 622
rect 67 522 99 554
rect 67 454 99 486
rect 169 590 201 622
rect 169 522 201 554
rect 169 454 201 486
rect 272 590 304 622
rect 272 522 304 554
rect 272 454 304 486
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 121 636 147 672
rect 223 636 249 672
rect 121 370 147 412
rect 61 353 147 370
rect 61 321 78 353
rect 110 334 147 353
rect 223 334 249 412
rect 110 321 249 334
rect 61 304 249 321
rect 121 266 147 304
rect 223 266 249 304
rect 121 82 147 118
rect 223 82 249 118
<< polycont >>
rect 78 321 110 353
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 57 622 109 712
rect 57 590 67 622
rect 99 590 109 622
rect 57 554 109 590
rect 57 522 67 554
rect 99 522 109 554
rect 57 486 109 522
rect 57 454 67 486
rect 99 454 109 486
rect 57 444 109 454
rect 159 622 211 636
rect 159 590 169 622
rect 201 590 211 622
rect 159 554 211 590
rect 159 522 169 554
rect 201 522 211 554
rect 159 486 211 522
rect 159 454 169 486
rect 201 454 211 486
rect 159 444 211 454
rect 262 622 314 712
rect 262 590 272 622
rect 304 590 314 622
rect 262 554 314 590
rect 262 522 272 554
rect 304 522 314 554
rect 262 486 314 522
rect 262 454 272 486
rect 304 454 314 486
rect 262 444 314 454
rect 174 370 211 444
rect 51 353 127 370
rect 51 321 78 353
rect 110 321 127 353
rect 51 304 127 321
rect 174 304 318 370
rect 174 242 211 304
rect 57 232 109 242
rect 57 200 67 232
rect 99 200 109 232
rect 57 164 109 200
rect 57 132 67 164
rect 99 132 109 164
rect 57 44 109 132
rect 159 232 211 242
rect 159 200 169 232
rect 201 200 211 232
rect 159 164 211 200
rect 159 132 169 164
rect 201 132 211 164
rect 159 122 211 132
rect 261 232 313 242
rect 261 200 271 232
rect 303 200 313 232
rect 261 164 313 200
rect 261 132 271 164
rect 303 132 313 164
rect 261 44 313 132
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 174 304 318 370 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 51 304 127 370 0 FreeSans 400 0 0 0 A
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 228462
string GDS_FILE 6_final.gds
string GDS_START 224758
<< end >>
