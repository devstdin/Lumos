magic
tech ihp-sg13g2
timestamp 1748514843
<< error_p >>
rect -43 1664 -38 1669
rect 38 1664 43 1669
rect 185 1664 190 1669
rect 266 1664 271 1669
rect 413 1664 418 1669
rect 494 1664 499 1669
rect 641 1664 646 1669
rect 722 1664 727 1669
rect 869 1664 874 1669
rect 950 1664 955 1669
rect 1097 1664 1102 1669
rect 1178 1664 1183 1669
rect 1325 1664 1330 1669
rect 1406 1664 1411 1669
rect 1553 1664 1558 1669
rect 1634 1664 1639 1669
rect 1781 1664 1786 1669
rect 1862 1664 1867 1669
rect 2009 1664 2014 1669
rect 2090 1664 2095 1669
rect 2237 1664 2242 1669
rect 2318 1664 2323 1669
rect 2465 1664 2470 1669
rect 2546 1664 2551 1669
rect 2693 1664 2698 1669
rect 2774 1664 2779 1669
rect 2921 1664 2926 1669
rect 3002 1664 3007 1669
rect 3149 1664 3154 1669
rect 3230 1664 3235 1669
rect 3377 1664 3382 1669
rect 3458 1664 3463 1669
rect -48 1659 -43 1664
rect 43 1659 48 1664
rect 180 1659 185 1664
rect 271 1659 276 1664
rect 408 1659 413 1664
rect 499 1659 504 1664
rect 636 1659 641 1664
rect 727 1659 732 1664
rect 864 1659 869 1664
rect 955 1659 960 1664
rect 1092 1659 1097 1664
rect 1183 1659 1188 1664
rect 1320 1659 1325 1664
rect 1411 1659 1416 1664
rect 1548 1659 1553 1664
rect 1639 1659 1644 1664
rect 1776 1659 1781 1664
rect 1867 1659 1872 1664
rect 2004 1659 2009 1664
rect 2095 1659 2100 1664
rect 2232 1659 2237 1664
rect 2323 1659 2328 1664
rect 2460 1659 2465 1664
rect 2551 1659 2556 1664
rect 2688 1659 2693 1664
rect 2779 1659 2784 1664
rect 2916 1659 2921 1664
rect 3007 1659 3012 1664
rect 3144 1659 3149 1664
rect 3235 1659 3240 1664
rect 3372 1659 3377 1664
rect 3463 1659 3468 1664
rect -48 1648 -43 1653
rect 43 1648 48 1653
rect 180 1648 185 1653
rect 271 1648 276 1653
rect 408 1648 413 1653
rect 499 1648 504 1653
rect 636 1648 641 1653
rect 727 1648 732 1653
rect 864 1648 869 1653
rect 955 1648 960 1653
rect 1092 1648 1097 1653
rect 1183 1648 1188 1653
rect 1320 1648 1325 1653
rect 1411 1648 1416 1653
rect 1548 1648 1553 1653
rect 1639 1648 1644 1653
rect 1776 1648 1781 1653
rect 1867 1648 1872 1653
rect 2004 1648 2009 1653
rect 2095 1648 2100 1653
rect 2232 1648 2237 1653
rect 2323 1648 2328 1653
rect 2460 1648 2465 1653
rect 2551 1648 2556 1653
rect 2688 1648 2693 1653
rect 2779 1648 2784 1653
rect 2916 1648 2921 1653
rect 3007 1648 3012 1653
rect 3144 1648 3149 1653
rect 3235 1648 3240 1653
rect 3372 1648 3377 1653
rect 3463 1648 3468 1653
rect -43 1643 -38 1648
rect 38 1643 43 1648
rect 185 1643 190 1648
rect 266 1643 271 1648
rect 413 1643 418 1648
rect 494 1643 499 1648
rect 641 1643 646 1648
rect 722 1643 727 1648
rect 869 1643 874 1648
rect 950 1643 955 1648
rect 1097 1643 1102 1648
rect 1178 1643 1183 1648
rect 1325 1643 1330 1648
rect 1406 1643 1411 1648
rect 1553 1643 1558 1648
rect 1634 1643 1639 1648
rect 1781 1643 1786 1648
rect 1862 1643 1867 1648
rect 2009 1643 2014 1648
rect 2090 1643 2095 1648
rect 2237 1643 2242 1648
rect 2318 1643 2323 1648
rect 2465 1643 2470 1648
rect 2546 1643 2551 1648
rect 2693 1643 2698 1648
rect 2774 1643 2779 1648
rect 2921 1643 2926 1648
rect 3002 1643 3007 1648
rect 3149 1643 3154 1648
rect 3230 1643 3235 1648
rect 3377 1643 3382 1648
rect 3458 1643 3463 1648
rect -77 1627 -72 1632
rect -66 1627 -61 1632
rect 61 1627 66 1632
rect 72 1627 77 1632
rect 151 1627 156 1632
rect 162 1627 167 1632
rect 289 1627 294 1632
rect 300 1627 305 1632
rect 379 1627 384 1632
rect 390 1627 395 1632
rect 517 1627 522 1632
rect 528 1627 533 1632
rect 607 1627 612 1632
rect 618 1627 623 1632
rect 745 1627 750 1632
rect 756 1627 761 1632
rect 835 1627 840 1632
rect 846 1627 851 1632
rect 973 1627 978 1632
rect 984 1627 989 1632
rect 1063 1627 1068 1632
rect 1074 1627 1079 1632
rect 1201 1627 1206 1632
rect 1212 1627 1217 1632
rect 1291 1627 1296 1632
rect 1302 1627 1307 1632
rect 1429 1627 1434 1632
rect 1440 1627 1445 1632
rect 1519 1627 1524 1632
rect 1530 1627 1535 1632
rect 1657 1627 1662 1632
rect 1668 1627 1673 1632
rect 1747 1627 1752 1632
rect 1758 1627 1763 1632
rect 1885 1627 1890 1632
rect 1896 1627 1901 1632
rect 1975 1627 1980 1632
rect 1986 1627 1991 1632
rect 2113 1627 2118 1632
rect 2124 1627 2129 1632
rect 2203 1627 2208 1632
rect 2214 1627 2219 1632
rect 2341 1627 2346 1632
rect 2352 1627 2357 1632
rect 2431 1627 2436 1632
rect 2442 1627 2447 1632
rect 2569 1627 2574 1632
rect 2580 1627 2585 1632
rect 2659 1627 2664 1632
rect 2670 1627 2675 1632
rect 2797 1627 2802 1632
rect 2808 1627 2813 1632
rect 2887 1627 2892 1632
rect 2898 1627 2903 1632
rect 3025 1627 3030 1632
rect 3036 1627 3041 1632
rect 3115 1627 3120 1632
rect 3126 1627 3131 1632
rect 3253 1627 3258 1632
rect 3264 1627 3269 1632
rect 3343 1627 3348 1632
rect 3354 1627 3359 1632
rect 3481 1627 3486 1632
rect 3492 1627 3497 1632
rect -82 1622 -77 1627
rect -61 1622 -56 1627
rect 56 1622 61 1627
rect 77 1622 82 1627
rect 146 1622 151 1627
rect 167 1622 172 1627
rect 284 1622 289 1627
rect 305 1622 310 1627
rect 374 1622 379 1627
rect 395 1622 400 1627
rect 512 1622 517 1627
rect 533 1622 538 1627
rect 602 1622 607 1627
rect 623 1622 628 1627
rect 740 1622 745 1627
rect 761 1622 766 1627
rect 830 1622 835 1627
rect 851 1622 856 1627
rect 968 1622 973 1627
rect 989 1622 994 1627
rect 1058 1622 1063 1627
rect 1079 1622 1084 1627
rect 1196 1622 1201 1627
rect 1217 1622 1222 1627
rect 1286 1622 1291 1627
rect 1307 1622 1312 1627
rect 1424 1622 1429 1627
rect 1445 1622 1450 1627
rect 1514 1622 1519 1627
rect 1535 1622 1540 1627
rect 1652 1622 1657 1627
rect 1673 1622 1678 1627
rect 1742 1622 1747 1627
rect 1763 1622 1768 1627
rect 1880 1622 1885 1627
rect 1901 1622 1906 1627
rect 1970 1622 1975 1627
rect 1991 1622 1996 1627
rect 2108 1622 2113 1627
rect 2129 1622 2134 1627
rect 2198 1622 2203 1627
rect 2219 1622 2224 1627
rect 2336 1622 2341 1627
rect 2357 1622 2362 1627
rect 2426 1622 2431 1627
rect 2447 1622 2452 1627
rect 2564 1622 2569 1627
rect 2585 1622 2590 1627
rect 2654 1622 2659 1627
rect 2675 1622 2680 1627
rect 2792 1622 2797 1627
rect 2813 1622 2818 1627
rect 2882 1622 2887 1627
rect 2903 1622 2908 1627
rect 3020 1622 3025 1627
rect 3041 1622 3046 1627
rect 3110 1622 3115 1627
rect 3131 1622 3136 1627
rect 3248 1622 3253 1627
rect 3269 1622 3274 1627
rect 3338 1622 3343 1627
rect 3359 1622 3364 1627
rect 3476 1622 3481 1627
rect 3497 1622 3502 1627
rect -82 641 -77 646
rect -61 641 -56 646
rect 56 641 61 646
rect 77 641 82 646
rect 146 641 151 646
rect 167 641 172 646
rect 284 641 289 646
rect 305 641 310 646
rect 374 641 379 646
rect 395 641 400 646
rect 512 641 517 646
rect 533 641 538 646
rect 602 641 607 646
rect 623 641 628 646
rect 740 641 745 646
rect 761 641 766 646
rect 830 641 835 646
rect 851 641 856 646
rect 968 641 973 646
rect 989 641 994 646
rect 1058 641 1063 646
rect 1079 641 1084 646
rect 1196 641 1201 646
rect 1217 641 1222 646
rect 1286 641 1291 646
rect 1307 641 1312 646
rect 1424 641 1429 646
rect 1445 641 1450 646
rect 1514 641 1519 646
rect 1535 641 1540 646
rect 1652 641 1657 646
rect 1673 641 1678 646
rect 1742 641 1747 646
rect 1763 641 1768 646
rect 1880 641 1885 646
rect 1901 641 1906 646
rect 1970 641 1975 646
rect 1991 641 1996 646
rect 2108 641 2113 646
rect 2129 641 2134 646
rect 2198 641 2203 646
rect 2219 641 2224 646
rect 2336 641 2341 646
rect 2357 641 2362 646
rect 2426 641 2431 646
rect 2447 641 2452 646
rect 2564 641 2569 646
rect 2585 641 2590 646
rect 2654 641 2659 646
rect 2675 641 2680 646
rect 2792 641 2797 646
rect 2813 641 2818 646
rect 2882 641 2887 646
rect 2903 641 2908 646
rect 3020 641 3025 646
rect 3041 641 3046 646
rect 3110 641 3115 646
rect 3131 641 3136 646
rect 3248 641 3253 646
rect 3269 641 3274 646
rect 3338 641 3343 646
rect 3359 641 3364 646
rect 3476 641 3481 646
rect 3497 641 3502 646
rect -77 636 -72 641
rect -66 636 -61 641
rect 61 636 66 641
rect 72 636 77 641
rect 151 636 156 641
rect 162 636 167 641
rect 289 636 294 641
rect 300 636 305 641
rect 379 636 384 641
rect 390 636 395 641
rect 517 636 522 641
rect 528 636 533 641
rect 607 636 612 641
rect 618 636 623 641
rect 745 636 750 641
rect 756 636 761 641
rect 835 636 840 641
rect 846 636 851 641
rect 973 636 978 641
rect 984 636 989 641
rect 1063 636 1068 641
rect 1074 636 1079 641
rect 1201 636 1206 641
rect 1212 636 1217 641
rect 1291 636 1296 641
rect 1302 636 1307 641
rect 1429 636 1434 641
rect 1440 636 1445 641
rect 1519 636 1524 641
rect 1530 636 1535 641
rect 1657 636 1662 641
rect 1668 636 1673 641
rect 1747 636 1752 641
rect 1758 636 1763 641
rect 1885 636 1890 641
rect 1896 636 1901 641
rect 1975 636 1980 641
rect 1986 636 1991 641
rect 2113 636 2118 641
rect 2124 636 2129 641
rect 2203 636 2208 641
rect 2214 636 2219 641
rect 2341 636 2346 641
rect 2352 636 2357 641
rect 2431 636 2436 641
rect 2442 636 2447 641
rect 2569 636 2574 641
rect 2580 636 2585 641
rect 2659 636 2664 641
rect 2670 636 2675 641
rect 2797 636 2802 641
rect 2808 636 2813 641
rect 2887 636 2892 641
rect 2898 636 2903 641
rect 3025 636 3030 641
rect 3036 636 3041 641
rect 3115 636 3120 641
rect 3126 636 3131 641
rect 3253 636 3258 641
rect 3264 636 3269 641
rect 3343 636 3348 641
rect 3354 636 3359 641
rect 3481 636 3486 641
rect 3492 636 3497 641
rect -43 620 -38 625
rect 38 620 43 625
rect 185 620 190 625
rect 266 620 271 625
rect 413 620 418 625
rect 494 620 499 625
rect 641 620 646 625
rect 722 620 727 625
rect 869 620 874 625
rect 950 620 955 625
rect 1097 620 1102 625
rect 1178 620 1183 625
rect 1325 620 1330 625
rect 1406 620 1411 625
rect 1553 620 1558 625
rect 1634 620 1639 625
rect 1781 620 1786 625
rect 1862 620 1867 625
rect 2009 620 2014 625
rect 2090 620 2095 625
rect 2237 620 2242 625
rect 2318 620 2323 625
rect 2465 620 2470 625
rect 2546 620 2551 625
rect 2693 620 2698 625
rect 2774 620 2779 625
rect 2921 620 2926 625
rect 3002 620 3007 625
rect 3149 620 3154 625
rect 3230 620 3235 625
rect 3377 620 3382 625
rect 3458 620 3463 625
rect -48 615 -43 620
rect 43 615 48 620
rect 180 615 185 620
rect 271 615 276 620
rect 408 615 413 620
rect 499 615 504 620
rect 636 615 641 620
rect 727 615 732 620
rect 864 615 869 620
rect 955 615 960 620
rect 1092 615 1097 620
rect 1183 615 1188 620
rect 1320 615 1325 620
rect 1411 615 1416 620
rect 1548 615 1553 620
rect 1639 615 1644 620
rect 1776 615 1781 620
rect 1867 615 1872 620
rect 2004 615 2009 620
rect 2095 615 2100 620
rect 2232 615 2237 620
rect 2323 615 2328 620
rect 2460 615 2465 620
rect 2551 615 2556 620
rect 2688 615 2693 620
rect 2779 615 2784 620
rect 2916 615 2921 620
rect 3007 615 3012 620
rect 3144 615 3149 620
rect 3235 615 3240 620
rect 3372 615 3377 620
rect 3463 615 3468 620
rect -48 604 -43 609
rect 43 604 48 609
rect 180 604 185 609
rect 271 604 276 609
rect 408 604 413 609
rect 499 604 504 609
rect 636 604 641 609
rect 727 604 732 609
rect 864 604 869 609
rect 955 604 960 609
rect 1092 604 1097 609
rect 1183 604 1188 609
rect 1320 604 1325 609
rect 1411 604 1416 609
rect 1548 604 1553 609
rect 1639 604 1644 609
rect 1776 604 1781 609
rect 1867 604 1872 609
rect 2004 604 2009 609
rect 2095 604 2100 609
rect 2232 604 2237 609
rect 2323 604 2328 609
rect 2460 604 2465 609
rect 2551 604 2556 609
rect 2688 604 2693 609
rect 2779 604 2784 609
rect 2916 604 2921 609
rect 3007 604 3012 609
rect 3144 604 3149 609
rect 3235 604 3240 609
rect 3372 604 3377 609
rect 3463 604 3468 609
rect -43 599 -38 604
rect 38 599 43 604
rect 185 599 190 604
rect 266 599 271 604
rect 413 599 418 604
rect 494 599 499 604
rect 641 599 646 604
rect 722 599 727 604
rect 869 599 874 604
rect 950 599 955 604
rect 1097 599 1102 604
rect 1178 599 1183 604
rect 1325 599 1330 604
rect 1406 599 1411 604
rect 1553 599 1558 604
rect 1634 599 1639 604
rect 1781 599 1786 604
rect 1862 599 1867 604
rect 2009 599 2014 604
rect 2090 599 2095 604
rect 2237 599 2242 604
rect 2318 599 2323 604
rect 2465 599 2470 604
rect 2546 599 2551 604
rect 2693 599 2698 604
rect 2774 599 2779 604
rect 2921 599 2926 604
rect 3002 599 3007 604
rect 3149 599 3154 604
rect 3230 599 3235 604
rect 3377 599 3382 604
rect 3458 599 3463 604
rect -43 530 -38 535
rect 38 530 43 535
rect 185 530 190 535
rect 266 530 271 535
rect 413 530 418 535
rect 494 530 499 535
rect 641 530 646 535
rect 722 530 727 535
rect 869 530 874 535
rect 950 530 955 535
rect 1097 530 1102 535
rect 1178 530 1183 535
rect 1325 530 1330 535
rect 1406 530 1411 535
rect 1553 530 1558 535
rect 1634 530 1639 535
rect 1781 530 1786 535
rect 1862 530 1867 535
rect 2009 530 2014 535
rect 2090 530 2095 535
rect 2237 530 2242 535
rect 2318 530 2323 535
rect 2465 530 2470 535
rect 2546 530 2551 535
rect 2693 530 2698 535
rect 2774 530 2779 535
rect 2921 530 2926 535
rect 3002 530 3007 535
rect 3149 530 3154 535
rect 3230 530 3235 535
rect 3377 530 3382 535
rect 3458 530 3463 535
rect -48 525 -43 530
rect 43 525 48 530
rect 180 525 185 530
rect 271 525 276 530
rect 408 525 413 530
rect 499 525 504 530
rect 636 525 641 530
rect 727 525 732 530
rect 864 525 869 530
rect 955 525 960 530
rect 1092 525 1097 530
rect 1183 525 1188 530
rect 1320 525 1325 530
rect 1411 525 1416 530
rect 1548 525 1553 530
rect 1639 525 1644 530
rect 1776 525 1781 530
rect 1867 525 1872 530
rect 2004 525 2009 530
rect 2095 525 2100 530
rect 2232 525 2237 530
rect 2323 525 2328 530
rect 2460 525 2465 530
rect 2551 525 2556 530
rect 2688 525 2693 530
rect 2779 525 2784 530
rect 2916 525 2921 530
rect 3007 525 3012 530
rect 3144 525 3149 530
rect 3235 525 3240 530
rect 3372 525 3377 530
rect 3463 525 3468 530
rect -48 514 -43 519
rect 43 514 48 519
rect 180 514 185 519
rect 271 514 276 519
rect 408 514 413 519
rect 499 514 504 519
rect 636 514 641 519
rect 727 514 732 519
rect 864 514 869 519
rect 955 514 960 519
rect 1092 514 1097 519
rect 1183 514 1188 519
rect 1320 514 1325 519
rect 1411 514 1416 519
rect 1548 514 1553 519
rect 1639 514 1644 519
rect 1776 514 1781 519
rect 1867 514 1872 519
rect 2004 514 2009 519
rect 2095 514 2100 519
rect 2232 514 2237 519
rect 2323 514 2328 519
rect 2460 514 2465 519
rect 2551 514 2556 519
rect 2688 514 2693 519
rect 2779 514 2784 519
rect 2916 514 2921 519
rect 3007 514 3012 519
rect 3144 514 3149 519
rect 3235 514 3240 519
rect 3372 514 3377 519
rect 3463 514 3468 519
rect -43 509 -38 514
rect 38 509 43 514
rect 185 509 190 514
rect 266 509 271 514
rect 413 509 418 514
rect 494 509 499 514
rect 641 509 646 514
rect 722 509 727 514
rect 869 509 874 514
rect 950 509 955 514
rect 1097 509 1102 514
rect 1178 509 1183 514
rect 1325 509 1330 514
rect 1406 509 1411 514
rect 1553 509 1558 514
rect 1634 509 1639 514
rect 1781 509 1786 514
rect 1862 509 1867 514
rect 2009 509 2014 514
rect 2090 509 2095 514
rect 2237 509 2242 514
rect 2318 509 2323 514
rect 2465 509 2470 514
rect 2546 509 2551 514
rect 2693 509 2698 514
rect 2774 509 2779 514
rect 2921 509 2926 514
rect 3002 509 3007 514
rect 3149 509 3154 514
rect 3230 509 3235 514
rect 3377 509 3382 514
rect 3458 509 3463 514
rect -77 493 -72 498
rect -66 493 -61 498
rect 61 493 66 498
rect 72 493 77 498
rect 151 493 156 498
rect 162 493 167 498
rect 289 493 294 498
rect 300 493 305 498
rect 379 493 384 498
rect 390 493 395 498
rect 517 493 522 498
rect 528 493 533 498
rect 607 493 612 498
rect 618 493 623 498
rect 745 493 750 498
rect 756 493 761 498
rect 835 493 840 498
rect 846 493 851 498
rect 973 493 978 498
rect 984 493 989 498
rect 1063 493 1068 498
rect 1074 493 1079 498
rect 1201 493 1206 498
rect 1212 493 1217 498
rect 1291 493 1296 498
rect 1302 493 1307 498
rect 1429 493 1434 498
rect 1440 493 1445 498
rect 1519 493 1524 498
rect 1530 493 1535 498
rect 1657 493 1662 498
rect 1668 493 1673 498
rect 1747 493 1752 498
rect 1758 493 1763 498
rect 1885 493 1890 498
rect 1896 493 1901 498
rect 1975 493 1980 498
rect 1986 493 1991 498
rect 2113 493 2118 498
rect 2124 493 2129 498
rect 2203 493 2208 498
rect 2214 493 2219 498
rect 2341 493 2346 498
rect 2352 493 2357 498
rect 2431 493 2436 498
rect 2442 493 2447 498
rect 2569 493 2574 498
rect 2580 493 2585 498
rect 2659 493 2664 498
rect 2670 493 2675 498
rect 2797 493 2802 498
rect 2808 493 2813 498
rect 2887 493 2892 498
rect 2898 493 2903 498
rect 3025 493 3030 498
rect 3036 493 3041 498
rect 3115 493 3120 498
rect 3126 493 3131 498
rect 3253 493 3258 498
rect 3264 493 3269 498
rect 3343 493 3348 498
rect 3354 493 3359 498
rect 3481 493 3486 498
rect 3492 493 3497 498
rect -82 488 -77 493
rect -61 488 -56 493
rect 56 488 61 493
rect 77 488 82 493
rect 146 488 151 493
rect 167 488 172 493
rect 284 488 289 493
rect 305 488 310 493
rect 374 488 379 493
rect 395 488 400 493
rect 512 488 517 493
rect 533 488 538 493
rect 602 488 607 493
rect 623 488 628 493
rect 740 488 745 493
rect 761 488 766 493
rect 830 488 835 493
rect 851 488 856 493
rect 968 488 973 493
rect 989 488 994 493
rect 1058 488 1063 493
rect 1079 488 1084 493
rect 1196 488 1201 493
rect 1217 488 1222 493
rect 1286 488 1291 493
rect 1307 488 1312 493
rect 1424 488 1429 493
rect 1445 488 1450 493
rect 1514 488 1519 493
rect 1535 488 1540 493
rect 1652 488 1657 493
rect 1673 488 1678 493
rect 1742 488 1747 493
rect 1763 488 1768 493
rect 1880 488 1885 493
rect 1901 488 1906 493
rect 1970 488 1975 493
rect 1991 488 1996 493
rect 2108 488 2113 493
rect 2129 488 2134 493
rect 2198 488 2203 493
rect 2219 488 2224 493
rect 2336 488 2341 493
rect 2357 488 2362 493
rect 2426 488 2431 493
rect 2447 488 2452 493
rect 2564 488 2569 493
rect 2585 488 2590 493
rect 2654 488 2659 493
rect 2675 488 2680 493
rect 2792 488 2797 493
rect 2813 488 2818 493
rect 2882 488 2887 493
rect 2903 488 2908 493
rect 3020 488 3025 493
rect 3041 488 3046 493
rect 3110 488 3115 493
rect 3131 488 3136 493
rect 3248 488 3253 493
rect 3269 488 3274 493
rect 3338 488 3343 493
rect 3359 488 3364 493
rect 3476 488 3481 493
rect 3497 488 3502 493
rect -82 -493 -77 -488
rect -61 -493 -56 -488
rect 56 -493 61 -488
rect 77 -493 82 -488
rect 146 -493 151 -488
rect 167 -493 172 -488
rect 284 -493 289 -488
rect 305 -493 310 -488
rect 374 -493 379 -488
rect 395 -493 400 -488
rect 512 -493 517 -488
rect 533 -493 538 -488
rect 602 -493 607 -488
rect 623 -493 628 -488
rect 740 -493 745 -488
rect 761 -493 766 -488
rect 830 -493 835 -488
rect 851 -493 856 -488
rect 968 -493 973 -488
rect 989 -493 994 -488
rect 1058 -493 1063 -488
rect 1079 -493 1084 -488
rect 1196 -493 1201 -488
rect 1217 -493 1222 -488
rect 1286 -493 1291 -488
rect 1307 -493 1312 -488
rect 1424 -493 1429 -488
rect 1445 -493 1450 -488
rect 1514 -493 1519 -488
rect 1535 -493 1540 -488
rect 1652 -493 1657 -488
rect 1673 -493 1678 -488
rect 1742 -493 1747 -488
rect 1763 -493 1768 -488
rect 1880 -493 1885 -488
rect 1901 -493 1906 -488
rect 1970 -493 1975 -488
rect 1991 -493 1996 -488
rect 2108 -493 2113 -488
rect 2129 -493 2134 -488
rect 2198 -493 2203 -488
rect 2219 -493 2224 -488
rect 2336 -493 2341 -488
rect 2357 -493 2362 -488
rect 2426 -493 2431 -488
rect 2447 -493 2452 -488
rect 2564 -493 2569 -488
rect 2585 -493 2590 -488
rect 2654 -493 2659 -488
rect 2675 -493 2680 -488
rect 2792 -493 2797 -488
rect 2813 -493 2818 -488
rect 2882 -493 2887 -488
rect 2903 -493 2908 -488
rect 3020 -493 3025 -488
rect 3041 -493 3046 -488
rect 3110 -493 3115 -488
rect 3131 -493 3136 -488
rect 3248 -493 3253 -488
rect 3269 -493 3274 -488
rect 3338 -493 3343 -488
rect 3359 -493 3364 -488
rect 3476 -493 3481 -488
rect 3497 -493 3502 -488
rect -77 -498 -72 -493
rect -66 -498 -61 -493
rect 61 -498 66 -493
rect 72 -498 77 -493
rect 151 -498 156 -493
rect 162 -498 167 -493
rect 289 -498 294 -493
rect 300 -498 305 -493
rect 379 -498 384 -493
rect 390 -498 395 -493
rect 517 -498 522 -493
rect 528 -498 533 -493
rect 607 -498 612 -493
rect 618 -498 623 -493
rect 745 -498 750 -493
rect 756 -498 761 -493
rect 835 -498 840 -493
rect 846 -498 851 -493
rect 973 -498 978 -493
rect 984 -498 989 -493
rect 1063 -498 1068 -493
rect 1074 -498 1079 -493
rect 1201 -498 1206 -493
rect 1212 -498 1217 -493
rect 1291 -498 1296 -493
rect 1302 -498 1307 -493
rect 1429 -498 1434 -493
rect 1440 -498 1445 -493
rect 1519 -498 1524 -493
rect 1530 -498 1535 -493
rect 1657 -498 1662 -493
rect 1668 -498 1673 -493
rect 1747 -498 1752 -493
rect 1758 -498 1763 -493
rect 1885 -498 1890 -493
rect 1896 -498 1901 -493
rect 1975 -498 1980 -493
rect 1986 -498 1991 -493
rect 2113 -498 2118 -493
rect 2124 -498 2129 -493
rect 2203 -498 2208 -493
rect 2214 -498 2219 -493
rect 2341 -498 2346 -493
rect 2352 -498 2357 -493
rect 2431 -498 2436 -493
rect 2442 -498 2447 -493
rect 2569 -498 2574 -493
rect 2580 -498 2585 -493
rect 2659 -498 2664 -493
rect 2670 -498 2675 -493
rect 2797 -498 2802 -493
rect 2808 -498 2813 -493
rect 2887 -498 2892 -493
rect 2898 -498 2903 -493
rect 3025 -498 3030 -493
rect 3036 -498 3041 -493
rect 3115 -498 3120 -493
rect 3126 -498 3131 -493
rect 3253 -498 3258 -493
rect 3264 -498 3269 -493
rect 3343 -498 3348 -493
rect 3354 -498 3359 -493
rect 3481 -498 3486 -493
rect 3492 -498 3497 -493
rect -43 -514 -38 -509
rect 38 -514 43 -509
rect 185 -514 190 -509
rect 266 -514 271 -509
rect 413 -514 418 -509
rect 494 -514 499 -509
rect 641 -514 646 -509
rect 722 -514 727 -509
rect 869 -514 874 -509
rect 950 -514 955 -509
rect 1097 -514 1102 -509
rect 1178 -514 1183 -509
rect 1325 -514 1330 -509
rect 1406 -514 1411 -509
rect 1553 -514 1558 -509
rect 1634 -514 1639 -509
rect 1781 -514 1786 -509
rect 1862 -514 1867 -509
rect 2009 -514 2014 -509
rect 2090 -514 2095 -509
rect 2237 -514 2242 -509
rect 2318 -514 2323 -509
rect 2465 -514 2470 -509
rect 2546 -514 2551 -509
rect 2693 -514 2698 -509
rect 2774 -514 2779 -509
rect 2921 -514 2926 -509
rect 3002 -514 3007 -509
rect 3149 -514 3154 -509
rect 3230 -514 3235 -509
rect 3377 -514 3382 -509
rect 3458 -514 3463 -509
rect -48 -519 -43 -514
rect 43 -519 48 -514
rect 180 -519 185 -514
rect 271 -519 276 -514
rect 408 -519 413 -514
rect 499 -519 504 -514
rect 636 -519 641 -514
rect 727 -519 732 -514
rect 864 -519 869 -514
rect 955 -519 960 -514
rect 1092 -519 1097 -514
rect 1183 -519 1188 -514
rect 1320 -519 1325 -514
rect 1411 -519 1416 -514
rect 1548 -519 1553 -514
rect 1639 -519 1644 -514
rect 1776 -519 1781 -514
rect 1867 -519 1872 -514
rect 2004 -519 2009 -514
rect 2095 -519 2100 -514
rect 2232 -519 2237 -514
rect 2323 -519 2328 -514
rect 2460 -519 2465 -514
rect 2551 -519 2556 -514
rect 2688 -519 2693 -514
rect 2779 -519 2784 -514
rect 2916 -519 2921 -514
rect 3007 -519 3012 -514
rect 3144 -519 3149 -514
rect 3235 -519 3240 -514
rect 3372 -519 3377 -514
rect 3463 -519 3468 -514
rect -48 -530 -43 -525
rect 43 -530 48 -525
rect 180 -530 185 -525
rect 271 -530 276 -525
rect 408 -530 413 -525
rect 499 -530 504 -525
rect 636 -530 641 -525
rect 727 -530 732 -525
rect 864 -530 869 -525
rect 955 -530 960 -525
rect 1092 -530 1097 -525
rect 1183 -530 1188 -525
rect 1320 -530 1325 -525
rect 1411 -530 1416 -525
rect 1548 -530 1553 -525
rect 1639 -530 1644 -525
rect 1776 -530 1781 -525
rect 1867 -530 1872 -525
rect 2004 -530 2009 -525
rect 2095 -530 2100 -525
rect 2232 -530 2237 -525
rect 2323 -530 2328 -525
rect 2460 -530 2465 -525
rect 2551 -530 2556 -525
rect 2688 -530 2693 -525
rect 2779 -530 2784 -525
rect 2916 -530 2921 -525
rect 3007 -530 3012 -525
rect 3144 -530 3149 -525
rect 3235 -530 3240 -525
rect 3372 -530 3377 -525
rect 3463 -530 3468 -525
rect -43 -535 -38 -530
rect 38 -535 43 -530
rect 185 -535 190 -530
rect 266 -535 271 -530
rect 413 -535 418 -530
rect 494 -535 499 -530
rect 641 -535 646 -530
rect 722 -535 727 -530
rect 869 -535 874 -530
rect 950 -535 955 -530
rect 1097 -535 1102 -530
rect 1178 -535 1183 -530
rect 1325 -535 1330 -530
rect 1406 -535 1411 -530
rect 1553 -535 1558 -530
rect 1634 -535 1639 -530
rect 1781 -535 1786 -530
rect 1862 -535 1867 -530
rect 2009 -535 2014 -530
rect 2090 -535 2095 -530
rect 2237 -535 2242 -530
rect 2318 -535 2323 -530
rect 2465 -535 2470 -530
rect 2546 -535 2551 -530
rect 2693 -535 2698 -530
rect 2774 -535 2779 -530
rect 2921 -535 2926 -530
rect 3002 -535 3007 -530
rect 3149 -535 3154 -530
rect 3230 -535 3235 -530
rect 3377 -535 3382 -530
rect 3458 -535 3463 -530
<< nwell >>
rect -230 -651 3650 1785
<< hvpmos >>
rect -50 634 50 1634
rect 178 634 278 1634
rect 406 634 506 1634
rect 634 634 734 1634
rect 862 634 962 1634
rect 1090 634 1190 1634
rect 1318 634 1418 1634
rect 1546 634 1646 1634
rect 1774 634 1874 1634
rect 2002 634 2102 1634
rect 2230 634 2330 1634
rect 2458 634 2558 1634
rect 2686 634 2786 1634
rect 2914 634 3014 1634
rect 3142 634 3242 1634
rect 3370 634 3470 1634
rect -50 -500 50 500
rect 178 -500 278 500
rect 406 -500 506 500
rect 634 -500 734 500
rect 862 -500 962 500
rect 1090 -500 1190 500
rect 1318 -500 1418 500
rect 1546 -500 1646 500
rect 1774 -500 1874 500
rect 2002 -500 2102 500
rect 2230 -500 2330 500
rect 2458 -500 2558 500
rect 2686 -500 2786 500
rect 2914 -500 3014 500
rect 3142 -500 3242 500
rect 3370 -500 3470 500
<< hvpdiff >>
rect -84 1627 -50 1634
rect -84 641 -77 1627
rect -61 641 -50 1627
rect -84 634 -50 641
rect 50 1627 84 1634
rect 50 641 61 1627
rect 77 641 84 1627
rect 50 634 84 641
rect 144 1627 178 1634
rect 144 641 151 1627
rect 167 641 178 1627
rect 144 634 178 641
rect 278 1627 312 1634
rect 278 641 289 1627
rect 305 641 312 1627
rect 278 634 312 641
rect 372 1627 406 1634
rect 372 641 379 1627
rect 395 641 406 1627
rect 372 634 406 641
rect 506 1627 540 1634
rect 506 641 517 1627
rect 533 641 540 1627
rect 506 634 540 641
rect 600 1627 634 1634
rect 600 641 607 1627
rect 623 641 634 1627
rect 600 634 634 641
rect 734 1627 768 1634
rect 734 641 745 1627
rect 761 641 768 1627
rect 734 634 768 641
rect 828 1627 862 1634
rect 828 641 835 1627
rect 851 641 862 1627
rect 828 634 862 641
rect 962 1627 996 1634
rect 962 641 973 1627
rect 989 641 996 1627
rect 962 634 996 641
rect 1056 1627 1090 1634
rect 1056 641 1063 1627
rect 1079 641 1090 1627
rect 1056 634 1090 641
rect 1190 1627 1224 1634
rect 1190 641 1201 1627
rect 1217 641 1224 1627
rect 1190 634 1224 641
rect 1284 1627 1318 1634
rect 1284 641 1291 1627
rect 1307 641 1318 1627
rect 1284 634 1318 641
rect 1418 1627 1452 1634
rect 1418 641 1429 1627
rect 1445 641 1452 1627
rect 1418 634 1452 641
rect 1512 1627 1546 1634
rect 1512 641 1519 1627
rect 1535 641 1546 1627
rect 1512 634 1546 641
rect 1646 1627 1680 1634
rect 1646 641 1657 1627
rect 1673 641 1680 1627
rect 1646 634 1680 641
rect 1740 1627 1774 1634
rect 1740 641 1747 1627
rect 1763 641 1774 1627
rect 1740 634 1774 641
rect 1874 1627 1908 1634
rect 1874 641 1885 1627
rect 1901 641 1908 1627
rect 1874 634 1908 641
rect 1968 1627 2002 1634
rect 1968 641 1975 1627
rect 1991 641 2002 1627
rect 1968 634 2002 641
rect 2102 1627 2136 1634
rect 2102 641 2113 1627
rect 2129 641 2136 1627
rect 2102 634 2136 641
rect 2196 1627 2230 1634
rect 2196 641 2203 1627
rect 2219 641 2230 1627
rect 2196 634 2230 641
rect 2330 1627 2364 1634
rect 2330 641 2341 1627
rect 2357 641 2364 1627
rect 2330 634 2364 641
rect 2424 1627 2458 1634
rect 2424 641 2431 1627
rect 2447 641 2458 1627
rect 2424 634 2458 641
rect 2558 1627 2592 1634
rect 2558 641 2569 1627
rect 2585 641 2592 1627
rect 2558 634 2592 641
rect 2652 1627 2686 1634
rect 2652 641 2659 1627
rect 2675 641 2686 1627
rect 2652 634 2686 641
rect 2786 1627 2820 1634
rect 2786 641 2797 1627
rect 2813 641 2820 1627
rect 2786 634 2820 641
rect 2880 1627 2914 1634
rect 2880 641 2887 1627
rect 2903 641 2914 1627
rect 2880 634 2914 641
rect 3014 1627 3048 1634
rect 3014 641 3025 1627
rect 3041 641 3048 1627
rect 3014 634 3048 641
rect 3108 1627 3142 1634
rect 3108 641 3115 1627
rect 3131 641 3142 1627
rect 3108 634 3142 641
rect 3242 1627 3276 1634
rect 3242 641 3253 1627
rect 3269 641 3276 1627
rect 3242 634 3276 641
rect 3336 1627 3370 1634
rect 3336 641 3343 1627
rect 3359 641 3370 1627
rect 3336 634 3370 641
rect 3470 1627 3504 1634
rect 3470 641 3481 1627
rect 3497 641 3504 1627
rect 3470 634 3504 641
rect -84 493 -50 500
rect -84 -493 -77 493
rect -61 -493 -50 493
rect -84 -500 -50 -493
rect 50 493 84 500
rect 50 -493 61 493
rect 77 -493 84 493
rect 50 -500 84 -493
rect 144 493 178 500
rect 144 -493 151 493
rect 167 -493 178 493
rect 144 -500 178 -493
rect 278 493 312 500
rect 278 -493 289 493
rect 305 -493 312 493
rect 278 -500 312 -493
rect 372 493 406 500
rect 372 -493 379 493
rect 395 -493 406 493
rect 372 -500 406 -493
rect 506 493 540 500
rect 506 -493 517 493
rect 533 -493 540 493
rect 506 -500 540 -493
rect 600 493 634 500
rect 600 -493 607 493
rect 623 -493 634 493
rect 600 -500 634 -493
rect 734 493 768 500
rect 734 -493 745 493
rect 761 -493 768 493
rect 734 -500 768 -493
rect 828 493 862 500
rect 828 -493 835 493
rect 851 -493 862 493
rect 828 -500 862 -493
rect 962 493 996 500
rect 962 -493 973 493
rect 989 -493 996 493
rect 962 -500 996 -493
rect 1056 493 1090 500
rect 1056 -493 1063 493
rect 1079 -493 1090 493
rect 1056 -500 1090 -493
rect 1190 493 1224 500
rect 1190 -493 1201 493
rect 1217 -493 1224 493
rect 1190 -500 1224 -493
rect 1284 493 1318 500
rect 1284 -493 1291 493
rect 1307 -493 1318 493
rect 1284 -500 1318 -493
rect 1418 493 1452 500
rect 1418 -493 1429 493
rect 1445 -493 1452 493
rect 1418 -500 1452 -493
rect 1512 493 1546 500
rect 1512 -493 1519 493
rect 1535 -493 1546 493
rect 1512 -500 1546 -493
rect 1646 493 1680 500
rect 1646 -493 1657 493
rect 1673 -493 1680 493
rect 1646 -500 1680 -493
rect 1740 493 1774 500
rect 1740 -493 1747 493
rect 1763 -493 1774 493
rect 1740 -500 1774 -493
rect 1874 493 1908 500
rect 1874 -493 1885 493
rect 1901 -493 1908 493
rect 1874 -500 1908 -493
rect 1968 493 2002 500
rect 1968 -493 1975 493
rect 1991 -493 2002 493
rect 1968 -500 2002 -493
rect 2102 493 2136 500
rect 2102 -493 2113 493
rect 2129 -493 2136 493
rect 2102 -500 2136 -493
rect 2196 493 2230 500
rect 2196 -493 2203 493
rect 2219 -493 2230 493
rect 2196 -500 2230 -493
rect 2330 493 2364 500
rect 2330 -493 2341 493
rect 2357 -493 2364 493
rect 2330 -500 2364 -493
rect 2424 493 2458 500
rect 2424 -493 2431 493
rect 2447 -493 2458 493
rect 2424 -500 2458 -493
rect 2558 493 2592 500
rect 2558 -493 2569 493
rect 2585 -493 2592 493
rect 2558 -500 2592 -493
rect 2652 493 2686 500
rect 2652 -493 2659 493
rect 2675 -493 2686 493
rect 2652 -500 2686 -493
rect 2786 493 2820 500
rect 2786 -493 2797 493
rect 2813 -493 2820 493
rect 2786 -500 2820 -493
rect 2880 493 2914 500
rect 2880 -493 2887 493
rect 2903 -493 2914 493
rect 2880 -500 2914 -493
rect 3014 493 3048 500
rect 3014 -493 3025 493
rect 3041 -493 3048 493
rect 3014 -500 3048 -493
rect 3108 493 3142 500
rect 3108 -493 3115 493
rect 3131 -493 3142 493
rect 3108 -500 3142 -493
rect 3242 493 3276 500
rect 3242 -493 3253 493
rect 3269 -493 3276 493
rect 3242 -500 3276 -493
rect 3336 493 3370 500
rect 3336 -493 3343 493
rect 3359 -493 3370 493
rect 3336 -500 3370 -493
rect 3470 493 3504 500
rect 3470 -493 3481 493
rect 3497 -493 3504 493
rect 3470 -500 3504 -493
<< hvpdiffc >>
rect -77 641 -61 1627
rect 61 641 77 1627
rect 151 641 167 1627
rect 289 641 305 1627
rect 379 641 395 1627
rect 517 641 533 1627
rect 607 641 623 1627
rect 745 641 761 1627
rect 835 641 851 1627
rect 973 641 989 1627
rect 1063 641 1079 1627
rect 1201 641 1217 1627
rect 1291 641 1307 1627
rect 1429 641 1445 1627
rect 1519 641 1535 1627
rect 1657 641 1673 1627
rect 1747 641 1763 1627
rect 1885 641 1901 1627
rect 1975 641 1991 1627
rect 2113 641 2129 1627
rect 2203 641 2219 1627
rect 2341 641 2357 1627
rect 2431 641 2447 1627
rect 2569 641 2585 1627
rect 2659 641 2675 1627
rect 2797 641 2813 1627
rect 2887 641 2903 1627
rect 3025 641 3041 1627
rect 3115 641 3131 1627
rect 3253 641 3269 1627
rect 3343 641 3359 1627
rect 3481 641 3497 1627
rect -77 -493 -61 493
rect 61 -493 77 493
rect 151 -493 167 493
rect 289 -493 305 493
rect 379 -493 395 493
rect 517 -493 533 493
rect 607 -493 623 493
rect 745 -493 761 493
rect 835 -493 851 493
rect 973 -493 989 493
rect 1063 -493 1079 493
rect 1201 -493 1217 493
rect 1291 -493 1307 493
rect 1429 -493 1445 493
rect 1519 -493 1535 493
rect 1657 -493 1673 493
rect 1747 -493 1763 493
rect 1885 -493 1901 493
rect 1975 -493 1991 493
rect 2113 -493 2129 493
rect 2203 -493 2219 493
rect 2341 -493 2357 493
rect 2431 -493 2447 493
rect 2569 -493 2585 493
rect 2659 -493 2675 493
rect 2797 -493 2813 493
rect 2887 -493 2903 493
rect 3025 -493 3041 493
rect 3115 -493 3131 493
rect 3253 -493 3269 493
rect 3343 -493 3359 493
rect 3481 -493 3497 493
<< nsubdiff >>
rect -168 1716 3588 1723
rect -168 1700 -131 1716
rect 3551 1700 3588 1716
rect -168 1693 3588 1700
rect -168 1686 -138 1693
rect -168 -552 -161 1686
rect -145 -552 -138 1686
rect 3558 1686 3588 1693
rect -168 -559 -138 -552
rect 3558 -552 3565 1686
rect 3581 -552 3588 1686
rect 3558 -559 3588 -552
rect -168 -566 3588 -559
rect -168 -582 -131 -566
rect 3551 -582 3588 -566
rect -168 -589 3588 -582
<< nsubdiffcont >>
rect -131 1700 3551 1716
rect -161 -552 -145 1686
rect 3565 -552 3581 1686
rect -131 -582 3551 -566
<< poly >>
rect -50 1664 50 1671
rect -50 1648 -43 1664
rect 43 1648 50 1664
rect -50 1634 50 1648
rect 178 1664 278 1671
rect 178 1648 185 1664
rect 271 1648 278 1664
rect 178 1634 278 1648
rect 406 1664 506 1671
rect 406 1648 413 1664
rect 499 1648 506 1664
rect 406 1634 506 1648
rect 634 1664 734 1671
rect 634 1648 641 1664
rect 727 1648 734 1664
rect 634 1634 734 1648
rect 862 1664 962 1671
rect 862 1648 869 1664
rect 955 1648 962 1664
rect 862 1634 962 1648
rect 1090 1664 1190 1671
rect 1090 1648 1097 1664
rect 1183 1648 1190 1664
rect 1090 1634 1190 1648
rect 1318 1664 1418 1671
rect 1318 1648 1325 1664
rect 1411 1648 1418 1664
rect 1318 1634 1418 1648
rect 1546 1664 1646 1671
rect 1546 1648 1553 1664
rect 1639 1648 1646 1664
rect 1546 1634 1646 1648
rect 1774 1664 1874 1671
rect 1774 1648 1781 1664
rect 1867 1648 1874 1664
rect 1774 1634 1874 1648
rect 2002 1664 2102 1671
rect 2002 1648 2009 1664
rect 2095 1648 2102 1664
rect 2002 1634 2102 1648
rect 2230 1664 2330 1671
rect 2230 1648 2237 1664
rect 2323 1648 2330 1664
rect 2230 1634 2330 1648
rect 2458 1664 2558 1671
rect 2458 1648 2465 1664
rect 2551 1648 2558 1664
rect 2458 1634 2558 1648
rect 2686 1664 2786 1671
rect 2686 1648 2693 1664
rect 2779 1648 2786 1664
rect 2686 1634 2786 1648
rect 2914 1664 3014 1671
rect 2914 1648 2921 1664
rect 3007 1648 3014 1664
rect 2914 1634 3014 1648
rect 3142 1664 3242 1671
rect 3142 1648 3149 1664
rect 3235 1648 3242 1664
rect 3142 1634 3242 1648
rect 3370 1664 3470 1671
rect 3370 1648 3377 1664
rect 3463 1648 3470 1664
rect 3370 1634 3470 1648
rect -50 620 50 634
rect -50 604 -43 620
rect 43 604 50 620
rect -50 597 50 604
rect 178 620 278 634
rect 178 604 185 620
rect 271 604 278 620
rect 178 597 278 604
rect 406 620 506 634
rect 406 604 413 620
rect 499 604 506 620
rect 406 597 506 604
rect 634 620 734 634
rect 634 604 641 620
rect 727 604 734 620
rect 634 597 734 604
rect 862 620 962 634
rect 862 604 869 620
rect 955 604 962 620
rect 862 597 962 604
rect 1090 620 1190 634
rect 1090 604 1097 620
rect 1183 604 1190 620
rect 1090 597 1190 604
rect 1318 620 1418 634
rect 1318 604 1325 620
rect 1411 604 1418 620
rect 1318 597 1418 604
rect 1546 620 1646 634
rect 1546 604 1553 620
rect 1639 604 1646 620
rect 1546 597 1646 604
rect 1774 620 1874 634
rect 1774 604 1781 620
rect 1867 604 1874 620
rect 1774 597 1874 604
rect 2002 620 2102 634
rect 2002 604 2009 620
rect 2095 604 2102 620
rect 2002 597 2102 604
rect 2230 620 2330 634
rect 2230 604 2237 620
rect 2323 604 2330 620
rect 2230 597 2330 604
rect 2458 620 2558 634
rect 2458 604 2465 620
rect 2551 604 2558 620
rect 2458 597 2558 604
rect 2686 620 2786 634
rect 2686 604 2693 620
rect 2779 604 2786 620
rect 2686 597 2786 604
rect 2914 620 3014 634
rect 2914 604 2921 620
rect 3007 604 3014 620
rect 2914 597 3014 604
rect 3142 620 3242 634
rect 3142 604 3149 620
rect 3235 604 3242 620
rect 3142 597 3242 604
rect 3370 620 3470 634
rect 3370 604 3377 620
rect 3463 604 3470 620
rect 3370 597 3470 604
rect -50 530 50 537
rect -50 514 -43 530
rect 43 514 50 530
rect -50 500 50 514
rect 178 530 278 537
rect 178 514 185 530
rect 271 514 278 530
rect 178 500 278 514
rect 406 530 506 537
rect 406 514 413 530
rect 499 514 506 530
rect 406 500 506 514
rect 634 530 734 537
rect 634 514 641 530
rect 727 514 734 530
rect 634 500 734 514
rect 862 530 962 537
rect 862 514 869 530
rect 955 514 962 530
rect 862 500 962 514
rect 1090 530 1190 537
rect 1090 514 1097 530
rect 1183 514 1190 530
rect 1090 500 1190 514
rect 1318 530 1418 537
rect 1318 514 1325 530
rect 1411 514 1418 530
rect 1318 500 1418 514
rect 1546 530 1646 537
rect 1546 514 1553 530
rect 1639 514 1646 530
rect 1546 500 1646 514
rect 1774 530 1874 537
rect 1774 514 1781 530
rect 1867 514 1874 530
rect 1774 500 1874 514
rect 2002 530 2102 537
rect 2002 514 2009 530
rect 2095 514 2102 530
rect 2002 500 2102 514
rect 2230 530 2330 537
rect 2230 514 2237 530
rect 2323 514 2330 530
rect 2230 500 2330 514
rect 2458 530 2558 537
rect 2458 514 2465 530
rect 2551 514 2558 530
rect 2458 500 2558 514
rect 2686 530 2786 537
rect 2686 514 2693 530
rect 2779 514 2786 530
rect 2686 500 2786 514
rect 2914 530 3014 537
rect 2914 514 2921 530
rect 3007 514 3014 530
rect 2914 500 3014 514
rect 3142 530 3242 537
rect 3142 514 3149 530
rect 3235 514 3242 530
rect 3142 500 3242 514
rect 3370 530 3470 537
rect 3370 514 3377 530
rect 3463 514 3470 530
rect 3370 500 3470 514
rect -50 -514 50 -500
rect -50 -530 -43 -514
rect 43 -530 50 -514
rect -50 -537 50 -530
rect 178 -514 278 -500
rect 178 -530 185 -514
rect 271 -530 278 -514
rect 178 -537 278 -530
rect 406 -514 506 -500
rect 406 -530 413 -514
rect 499 -530 506 -514
rect 406 -537 506 -530
rect 634 -514 734 -500
rect 634 -530 641 -514
rect 727 -530 734 -514
rect 634 -537 734 -530
rect 862 -514 962 -500
rect 862 -530 869 -514
rect 955 -530 962 -514
rect 862 -537 962 -530
rect 1090 -514 1190 -500
rect 1090 -530 1097 -514
rect 1183 -530 1190 -514
rect 1090 -537 1190 -530
rect 1318 -514 1418 -500
rect 1318 -530 1325 -514
rect 1411 -530 1418 -514
rect 1318 -537 1418 -530
rect 1546 -514 1646 -500
rect 1546 -530 1553 -514
rect 1639 -530 1646 -514
rect 1546 -537 1646 -530
rect 1774 -514 1874 -500
rect 1774 -530 1781 -514
rect 1867 -530 1874 -514
rect 1774 -537 1874 -530
rect 2002 -514 2102 -500
rect 2002 -530 2009 -514
rect 2095 -530 2102 -514
rect 2002 -537 2102 -530
rect 2230 -514 2330 -500
rect 2230 -530 2237 -514
rect 2323 -530 2330 -514
rect 2230 -537 2330 -530
rect 2458 -514 2558 -500
rect 2458 -530 2465 -514
rect 2551 -530 2558 -514
rect 2458 -537 2558 -530
rect 2686 -514 2786 -500
rect 2686 -530 2693 -514
rect 2779 -530 2786 -514
rect 2686 -537 2786 -530
rect 2914 -514 3014 -500
rect 2914 -530 2921 -514
rect 3007 -530 3014 -514
rect 2914 -537 3014 -530
rect 3142 -514 3242 -500
rect 3142 -530 3149 -514
rect 3235 -530 3242 -514
rect 3142 -537 3242 -530
rect 3370 -514 3470 -500
rect 3370 -530 3377 -514
rect 3463 -530 3470 -514
rect 3370 -537 3470 -530
<< polycont >>
rect -43 1648 43 1664
rect 185 1648 271 1664
rect 413 1648 499 1664
rect 641 1648 727 1664
rect 869 1648 955 1664
rect 1097 1648 1183 1664
rect 1325 1648 1411 1664
rect 1553 1648 1639 1664
rect 1781 1648 1867 1664
rect 2009 1648 2095 1664
rect 2237 1648 2323 1664
rect 2465 1648 2551 1664
rect 2693 1648 2779 1664
rect 2921 1648 3007 1664
rect 3149 1648 3235 1664
rect 3377 1648 3463 1664
rect -43 604 43 620
rect 185 604 271 620
rect 413 604 499 620
rect 641 604 727 620
rect 869 604 955 620
rect 1097 604 1183 620
rect 1325 604 1411 620
rect 1553 604 1639 620
rect 1781 604 1867 620
rect 2009 604 2095 620
rect 2237 604 2323 620
rect 2465 604 2551 620
rect 2693 604 2779 620
rect 2921 604 3007 620
rect 3149 604 3235 620
rect 3377 604 3463 620
rect -43 514 43 530
rect 185 514 271 530
rect 413 514 499 530
rect 641 514 727 530
rect 869 514 955 530
rect 1097 514 1183 530
rect 1325 514 1411 530
rect 1553 514 1639 530
rect 1781 514 1867 530
rect 2009 514 2095 530
rect 2237 514 2323 530
rect 2465 514 2551 530
rect 2693 514 2779 530
rect 2921 514 3007 530
rect 3149 514 3235 530
rect 3377 514 3463 530
rect -43 -530 43 -514
rect 185 -530 271 -514
rect 413 -530 499 -514
rect 641 -530 727 -514
rect 869 -530 955 -514
rect 1097 -530 1183 -514
rect 1325 -530 1411 -514
rect 1553 -530 1639 -514
rect 1781 -530 1867 -514
rect 2009 -530 2095 -514
rect 2237 -530 2323 -514
rect 2465 -530 2551 -514
rect 2693 -530 2779 -514
rect 2921 -530 3007 -514
rect 3149 -530 3235 -514
rect 3377 -530 3463 -514
<< metal1 >>
rect -166 1716 3586 1721
rect -166 1700 -131 1716
rect 3551 1700 3586 1716
rect -166 1695 3586 1700
rect -166 1686 -140 1695
rect -166 -552 -161 1686
rect -145 -552 -140 1686
rect 3560 1686 3586 1695
rect -166 -561 -140 -552
rect 3560 -552 3565 1686
rect 3581 -552 3586 1686
rect 3560 -561 3586 -552
rect -166 -566 3586 -561
rect -166 -582 -131 -566
rect 3551 -582 3586 -566
rect -166 -587 3586 -582
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 10 l 1 nf 1 nx 16 dx 0.6 ny 2 dy 0.6 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
