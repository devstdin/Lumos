magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -924 4124 37600
<< isosubstrate >>
rect 50 23124 1950 28034
rect 50 18112 1950 22924
rect 50 13000 1950 17912
<< nwell >>
rect -124 33246 2124 33554
rect -124 29546 2124 29854
rect -124 1076 2124 12324
<< pwell >>
rect 24 31344 1976 31456
rect 24 12974 1976 28060
<< psubdiff >>
rect 768 31384 800 31416
rect 838 31384 870 31416
rect 907 31384 939 31416
rect 978 31384 1010 31416
rect 1048 31384 1080 31416
rect 1116 31384 1148 31416
rect 1186 31384 1218 31416
rect 192 27939 224 27971
rect 264 27939 296 27971
rect 336 27939 368 27971
rect 408 27939 440 27971
rect 480 27939 512 27971
rect 552 27939 584 27971
rect 624 27939 656 27971
rect 696 27939 728 27971
rect 768 27939 800 27971
rect 840 27939 872 27971
rect 912 27939 944 27971
rect 984 27939 1016 27971
rect 1056 27939 1088 27971
rect 1128 27939 1160 27971
rect 1200 27939 1232 27971
rect 1272 27939 1304 27971
rect 1344 27939 1376 27971
rect 1416 27939 1448 27971
rect 1488 27939 1520 27971
rect 1560 27939 1592 27971
rect 1632 27939 1664 27971
rect 1704 27939 1736 27971
rect 1776 27939 1808 27971
rect 1848 27939 1880 27971
rect 120 27867 152 27899
rect 192 27867 224 27899
rect 264 27867 296 27899
rect 336 27867 368 27899
rect 408 27867 440 27899
rect 480 27867 512 27899
rect 552 27867 584 27899
rect 624 27867 656 27899
rect 696 27867 728 27899
rect 768 27867 800 27899
rect 840 27867 872 27899
rect 912 27867 944 27899
rect 984 27867 1016 27899
rect 1056 27867 1088 27899
rect 1128 27867 1160 27899
rect 1200 27867 1232 27899
rect 1272 27867 1304 27899
rect 1344 27867 1376 27899
rect 1416 27867 1448 27899
rect 1488 27867 1520 27899
rect 1560 27867 1592 27899
rect 1632 27867 1664 27899
rect 1704 27867 1736 27899
rect 1776 27867 1808 27899
rect 1848 27867 1880 27899
rect 120 27795 152 27827
rect 192 27795 224 27827
rect 264 27795 296 27827
rect 336 27795 368 27827
rect 408 27795 440 27827
rect 480 27795 512 27827
rect 552 27795 584 27827
rect 624 27795 656 27827
rect 696 27795 728 27827
rect 768 27795 800 27827
rect 840 27795 872 27827
rect 912 27795 944 27827
rect 984 27795 1016 27827
rect 1056 27795 1088 27827
rect 1128 27795 1160 27827
rect 1200 27795 1232 27827
rect 1272 27795 1304 27827
rect 1344 27795 1376 27827
rect 1416 27795 1448 27827
rect 1488 27795 1520 27827
rect 1560 27795 1592 27827
rect 1632 27795 1664 27827
rect 1704 27795 1736 27827
rect 1776 27795 1808 27827
rect 1848 27795 1880 27827
rect 120 27723 152 27755
rect 192 27723 224 27755
rect 264 27723 296 27755
rect 336 27723 368 27755
rect 408 27723 440 27755
rect 480 27723 512 27755
rect 552 27723 584 27755
rect 624 27723 656 27755
rect 696 27723 728 27755
rect 768 27723 800 27755
rect 840 27723 872 27755
rect 912 27723 944 27755
rect 984 27723 1016 27755
rect 1056 27723 1088 27755
rect 1128 27723 1160 27755
rect 1200 27723 1232 27755
rect 1272 27723 1304 27755
rect 1344 27723 1376 27755
rect 1416 27723 1448 27755
rect 1488 27723 1520 27755
rect 1560 27723 1592 27755
rect 1632 27723 1664 27755
rect 1704 27723 1736 27755
rect 1776 27723 1808 27755
rect 1848 27723 1880 27755
rect 120 27651 152 27683
rect 192 27651 224 27683
rect 264 27651 296 27683
rect 336 27651 368 27683
rect 408 27651 440 27683
rect 480 27651 512 27683
rect 552 27651 584 27683
rect 624 27651 656 27683
rect 696 27651 728 27683
rect 768 27651 800 27683
rect 840 27651 872 27683
rect 912 27651 944 27683
rect 984 27651 1016 27683
rect 1056 27651 1088 27683
rect 1128 27651 1160 27683
rect 1200 27651 1232 27683
rect 1272 27651 1304 27683
rect 1344 27651 1376 27683
rect 1416 27651 1448 27683
rect 1488 27651 1520 27683
rect 1560 27651 1592 27683
rect 1632 27651 1664 27683
rect 1704 27651 1736 27683
rect 1776 27651 1808 27683
rect 1848 27651 1880 27683
rect 120 27579 152 27611
rect 192 27579 224 27611
rect 264 27579 296 27611
rect 336 27579 368 27611
rect 408 27579 440 27611
rect 480 27579 512 27611
rect 552 27579 584 27611
rect 624 27579 656 27611
rect 696 27579 728 27611
rect 768 27579 800 27611
rect 840 27579 872 27611
rect 912 27579 944 27611
rect 984 27579 1016 27611
rect 1056 27579 1088 27611
rect 1128 27579 1160 27611
rect 1200 27579 1232 27611
rect 1272 27579 1304 27611
rect 1344 27579 1376 27611
rect 1416 27579 1448 27611
rect 1488 27579 1520 27611
rect 1560 27579 1592 27611
rect 1632 27579 1664 27611
rect 1704 27579 1736 27611
rect 1776 27579 1808 27611
rect 1848 27579 1880 27611
rect 120 27507 152 27539
rect 192 27507 224 27539
rect 264 27507 296 27539
rect 336 27507 368 27539
rect 408 27507 440 27539
rect 480 27507 512 27539
rect 552 27507 584 27539
rect 624 27507 656 27539
rect 696 27507 728 27539
rect 768 27507 800 27539
rect 840 27507 872 27539
rect 912 27507 944 27539
rect 984 27507 1016 27539
rect 1056 27507 1088 27539
rect 1128 27507 1160 27539
rect 1200 27507 1232 27539
rect 1272 27507 1304 27539
rect 1344 27507 1376 27539
rect 1416 27507 1448 27539
rect 1488 27507 1520 27539
rect 1560 27507 1592 27539
rect 1632 27507 1664 27539
rect 1704 27507 1736 27539
rect 1776 27507 1808 27539
rect 1848 27507 1880 27539
rect 120 27435 152 27467
rect 192 27435 224 27467
rect 264 27435 296 27467
rect 336 27435 368 27467
rect 408 27435 440 27467
rect 480 27435 512 27467
rect 552 27435 584 27467
rect 624 27435 656 27467
rect 696 27435 728 27467
rect 768 27435 800 27467
rect 840 27435 872 27467
rect 912 27435 944 27467
rect 984 27435 1016 27467
rect 1056 27435 1088 27467
rect 1128 27435 1160 27467
rect 1200 27435 1232 27467
rect 1272 27435 1304 27467
rect 1344 27435 1376 27467
rect 1416 27435 1448 27467
rect 1488 27435 1520 27467
rect 1560 27435 1592 27467
rect 1632 27435 1664 27467
rect 1704 27435 1736 27467
rect 1776 27435 1808 27467
rect 1848 27435 1880 27467
rect 120 27363 152 27395
rect 192 27363 224 27395
rect 264 27363 296 27395
rect 336 27363 368 27395
rect 408 27363 440 27395
rect 480 27363 512 27395
rect 552 27363 584 27395
rect 624 27363 656 27395
rect 696 27363 728 27395
rect 768 27363 800 27395
rect 840 27363 872 27395
rect 912 27363 944 27395
rect 984 27363 1016 27395
rect 1056 27363 1088 27395
rect 1128 27363 1160 27395
rect 1200 27363 1232 27395
rect 1272 27363 1304 27395
rect 1344 27363 1376 27395
rect 1416 27363 1448 27395
rect 1488 27363 1520 27395
rect 1560 27363 1592 27395
rect 1632 27363 1664 27395
rect 1704 27363 1736 27395
rect 1776 27363 1808 27395
rect 1848 27363 1880 27395
rect 120 27291 152 27323
rect 192 27291 224 27323
rect 264 27291 296 27323
rect 336 27291 368 27323
rect 408 27291 440 27323
rect 480 27291 512 27323
rect 552 27291 584 27323
rect 624 27291 656 27323
rect 696 27291 728 27323
rect 768 27291 800 27323
rect 840 27291 872 27323
rect 912 27291 944 27323
rect 984 27291 1016 27323
rect 1056 27291 1088 27323
rect 1128 27291 1160 27323
rect 1200 27291 1232 27323
rect 1272 27291 1304 27323
rect 1344 27291 1376 27323
rect 1416 27291 1448 27323
rect 1488 27291 1520 27323
rect 1560 27291 1592 27323
rect 1632 27291 1664 27323
rect 1704 27291 1736 27323
rect 1776 27291 1808 27323
rect 1848 27291 1880 27323
rect 120 27219 152 27251
rect 192 27219 224 27251
rect 264 27219 296 27251
rect 336 27219 368 27251
rect 408 27219 440 27251
rect 480 27219 512 27251
rect 552 27219 584 27251
rect 624 27219 656 27251
rect 696 27219 728 27251
rect 768 27219 800 27251
rect 840 27219 872 27251
rect 912 27219 944 27251
rect 984 27219 1016 27251
rect 1056 27219 1088 27251
rect 1128 27219 1160 27251
rect 1200 27219 1232 27251
rect 1272 27219 1304 27251
rect 1344 27219 1376 27251
rect 1416 27219 1448 27251
rect 1488 27219 1520 27251
rect 1560 27219 1592 27251
rect 1632 27219 1664 27251
rect 1704 27219 1736 27251
rect 1776 27219 1808 27251
rect 1848 27219 1880 27251
rect 120 27147 152 27179
rect 192 27147 224 27179
rect 264 27147 296 27179
rect 336 27147 368 27179
rect 408 27147 440 27179
rect 480 27147 512 27179
rect 552 27147 584 27179
rect 624 27147 656 27179
rect 696 27147 728 27179
rect 768 27147 800 27179
rect 840 27147 872 27179
rect 912 27147 944 27179
rect 984 27147 1016 27179
rect 1056 27147 1088 27179
rect 1128 27147 1160 27179
rect 1200 27147 1232 27179
rect 1272 27147 1304 27179
rect 1344 27147 1376 27179
rect 1416 27147 1448 27179
rect 1488 27147 1520 27179
rect 1560 27147 1592 27179
rect 1632 27147 1664 27179
rect 1704 27147 1736 27179
rect 1776 27147 1808 27179
rect 1848 27147 1880 27179
rect 120 27075 152 27107
rect 192 27075 224 27107
rect 264 27075 296 27107
rect 336 27075 368 27107
rect 408 27075 440 27107
rect 480 27075 512 27107
rect 552 27075 584 27107
rect 624 27075 656 27107
rect 696 27075 728 27107
rect 768 27075 800 27107
rect 840 27075 872 27107
rect 912 27075 944 27107
rect 984 27075 1016 27107
rect 1056 27075 1088 27107
rect 1128 27075 1160 27107
rect 1200 27075 1232 27107
rect 1272 27075 1304 27107
rect 1344 27075 1376 27107
rect 1416 27075 1448 27107
rect 1488 27075 1520 27107
rect 1560 27075 1592 27107
rect 1632 27075 1664 27107
rect 1704 27075 1736 27107
rect 1776 27075 1808 27107
rect 1848 27075 1880 27107
rect 120 27003 152 27035
rect 192 27003 224 27035
rect 264 27003 296 27035
rect 336 27003 368 27035
rect 408 27003 440 27035
rect 480 27003 512 27035
rect 552 27003 584 27035
rect 624 27003 656 27035
rect 696 27003 728 27035
rect 768 27003 800 27035
rect 840 27003 872 27035
rect 912 27003 944 27035
rect 984 27003 1016 27035
rect 1056 27003 1088 27035
rect 1128 27003 1160 27035
rect 1200 27003 1232 27035
rect 1272 27003 1304 27035
rect 1344 27003 1376 27035
rect 1416 27003 1448 27035
rect 1488 27003 1520 27035
rect 1560 27003 1592 27035
rect 1632 27003 1664 27035
rect 1704 27003 1736 27035
rect 1776 27003 1808 27035
rect 1848 27003 1880 27035
rect 120 26931 152 26963
rect 192 26931 224 26963
rect 264 26931 296 26963
rect 336 26931 368 26963
rect 408 26931 440 26963
rect 480 26931 512 26963
rect 552 26931 584 26963
rect 624 26931 656 26963
rect 696 26931 728 26963
rect 768 26931 800 26963
rect 840 26931 872 26963
rect 912 26931 944 26963
rect 984 26931 1016 26963
rect 1056 26931 1088 26963
rect 1128 26931 1160 26963
rect 1200 26931 1232 26963
rect 1272 26931 1304 26963
rect 1344 26931 1376 26963
rect 1416 26931 1448 26963
rect 1488 26931 1520 26963
rect 1560 26931 1592 26963
rect 1632 26931 1664 26963
rect 1704 26931 1736 26963
rect 1776 26931 1808 26963
rect 1848 26931 1880 26963
rect 120 26859 152 26891
rect 192 26859 224 26891
rect 264 26859 296 26891
rect 336 26859 368 26891
rect 408 26859 440 26891
rect 480 26859 512 26891
rect 552 26859 584 26891
rect 624 26859 656 26891
rect 696 26859 728 26891
rect 768 26859 800 26891
rect 840 26859 872 26891
rect 912 26859 944 26891
rect 984 26859 1016 26891
rect 1056 26859 1088 26891
rect 1128 26859 1160 26891
rect 1200 26859 1232 26891
rect 1272 26859 1304 26891
rect 1344 26859 1376 26891
rect 1416 26859 1448 26891
rect 1488 26859 1520 26891
rect 1560 26859 1592 26891
rect 1632 26859 1664 26891
rect 1704 26859 1736 26891
rect 1776 26859 1808 26891
rect 1848 26859 1880 26891
rect 120 26787 152 26819
rect 192 26787 224 26819
rect 264 26787 296 26819
rect 336 26787 368 26819
rect 408 26787 440 26819
rect 480 26787 512 26819
rect 552 26787 584 26819
rect 624 26787 656 26819
rect 696 26787 728 26819
rect 768 26787 800 26819
rect 840 26787 872 26819
rect 912 26787 944 26819
rect 984 26787 1016 26819
rect 1056 26787 1088 26819
rect 1128 26787 1160 26819
rect 1200 26787 1232 26819
rect 1272 26787 1304 26819
rect 1344 26787 1376 26819
rect 1416 26787 1448 26819
rect 1488 26787 1520 26819
rect 1560 26787 1592 26819
rect 1632 26787 1664 26819
rect 1704 26787 1736 26819
rect 1776 26787 1808 26819
rect 1848 26787 1880 26819
rect 120 26715 152 26747
rect 192 26715 224 26747
rect 264 26715 296 26747
rect 336 26715 368 26747
rect 408 26715 440 26747
rect 480 26715 512 26747
rect 552 26715 584 26747
rect 624 26715 656 26747
rect 696 26715 728 26747
rect 768 26715 800 26747
rect 840 26715 872 26747
rect 912 26715 944 26747
rect 984 26715 1016 26747
rect 1056 26715 1088 26747
rect 1128 26715 1160 26747
rect 1200 26715 1232 26747
rect 1272 26715 1304 26747
rect 1344 26715 1376 26747
rect 1416 26715 1448 26747
rect 1488 26715 1520 26747
rect 1560 26715 1592 26747
rect 1632 26715 1664 26747
rect 1704 26715 1736 26747
rect 1776 26715 1808 26747
rect 1848 26715 1880 26747
rect 120 26643 152 26675
rect 192 26643 224 26675
rect 264 26643 296 26675
rect 336 26643 368 26675
rect 408 26643 440 26675
rect 480 26643 512 26675
rect 552 26643 584 26675
rect 624 26643 656 26675
rect 696 26643 728 26675
rect 768 26643 800 26675
rect 840 26643 872 26675
rect 912 26643 944 26675
rect 984 26643 1016 26675
rect 1056 26643 1088 26675
rect 1128 26643 1160 26675
rect 1200 26643 1232 26675
rect 1272 26643 1304 26675
rect 1344 26643 1376 26675
rect 1416 26643 1448 26675
rect 1488 26643 1520 26675
rect 1560 26643 1592 26675
rect 1632 26643 1664 26675
rect 1704 26643 1736 26675
rect 1776 26643 1808 26675
rect 1848 26643 1880 26675
rect 120 26571 152 26603
rect 192 26571 224 26603
rect 264 26571 296 26603
rect 336 26571 368 26603
rect 408 26571 440 26603
rect 480 26571 512 26603
rect 552 26571 584 26603
rect 624 26571 656 26603
rect 696 26571 728 26603
rect 768 26571 800 26603
rect 840 26571 872 26603
rect 912 26571 944 26603
rect 984 26571 1016 26603
rect 1056 26571 1088 26603
rect 1128 26571 1160 26603
rect 1200 26571 1232 26603
rect 1272 26571 1304 26603
rect 1344 26571 1376 26603
rect 1416 26571 1448 26603
rect 1488 26571 1520 26603
rect 1560 26571 1592 26603
rect 1632 26571 1664 26603
rect 1704 26571 1736 26603
rect 1776 26571 1808 26603
rect 1848 26571 1880 26603
rect 120 26499 152 26531
rect 192 26499 224 26531
rect 264 26499 296 26531
rect 336 26499 368 26531
rect 408 26499 440 26531
rect 480 26499 512 26531
rect 552 26499 584 26531
rect 624 26499 656 26531
rect 696 26499 728 26531
rect 768 26499 800 26531
rect 840 26499 872 26531
rect 912 26499 944 26531
rect 984 26499 1016 26531
rect 1056 26499 1088 26531
rect 1128 26499 1160 26531
rect 1200 26499 1232 26531
rect 1272 26499 1304 26531
rect 1344 26499 1376 26531
rect 1416 26499 1448 26531
rect 1488 26499 1520 26531
rect 1560 26499 1592 26531
rect 1632 26499 1664 26531
rect 1704 26499 1736 26531
rect 1776 26499 1808 26531
rect 1848 26499 1880 26531
rect 120 26427 152 26459
rect 192 26427 224 26459
rect 264 26427 296 26459
rect 336 26427 368 26459
rect 408 26427 440 26459
rect 480 26427 512 26459
rect 552 26427 584 26459
rect 624 26427 656 26459
rect 696 26427 728 26459
rect 768 26427 800 26459
rect 840 26427 872 26459
rect 912 26427 944 26459
rect 984 26427 1016 26459
rect 1056 26427 1088 26459
rect 1128 26427 1160 26459
rect 1200 26427 1232 26459
rect 1272 26427 1304 26459
rect 1344 26427 1376 26459
rect 1416 26427 1448 26459
rect 1488 26427 1520 26459
rect 1560 26427 1592 26459
rect 1632 26427 1664 26459
rect 1704 26427 1736 26459
rect 1776 26427 1808 26459
rect 1848 26427 1880 26459
rect 120 26355 152 26387
rect 192 26355 224 26387
rect 264 26355 296 26387
rect 336 26355 368 26387
rect 408 26355 440 26387
rect 480 26355 512 26387
rect 552 26355 584 26387
rect 624 26355 656 26387
rect 696 26355 728 26387
rect 768 26355 800 26387
rect 840 26355 872 26387
rect 912 26355 944 26387
rect 984 26355 1016 26387
rect 1056 26355 1088 26387
rect 1128 26355 1160 26387
rect 1200 26355 1232 26387
rect 1272 26355 1304 26387
rect 1344 26355 1376 26387
rect 1416 26355 1448 26387
rect 1488 26355 1520 26387
rect 1560 26355 1592 26387
rect 1632 26355 1664 26387
rect 1704 26355 1736 26387
rect 1776 26355 1808 26387
rect 1848 26355 1880 26387
rect 120 26283 152 26315
rect 192 26283 224 26315
rect 264 26283 296 26315
rect 336 26283 368 26315
rect 408 26283 440 26315
rect 480 26283 512 26315
rect 552 26283 584 26315
rect 624 26283 656 26315
rect 696 26283 728 26315
rect 768 26283 800 26315
rect 840 26283 872 26315
rect 912 26283 944 26315
rect 984 26283 1016 26315
rect 1056 26283 1088 26315
rect 1128 26283 1160 26315
rect 1200 26283 1232 26315
rect 1272 26283 1304 26315
rect 1344 26283 1376 26315
rect 1416 26283 1448 26315
rect 1488 26283 1520 26315
rect 1560 26283 1592 26315
rect 1632 26283 1664 26315
rect 1704 26283 1736 26315
rect 1776 26283 1808 26315
rect 1848 26283 1880 26315
rect 120 26211 152 26243
rect 192 26211 224 26243
rect 264 26211 296 26243
rect 336 26211 368 26243
rect 408 26211 440 26243
rect 480 26211 512 26243
rect 552 26211 584 26243
rect 624 26211 656 26243
rect 696 26211 728 26243
rect 768 26211 800 26243
rect 840 26211 872 26243
rect 912 26211 944 26243
rect 984 26211 1016 26243
rect 1056 26211 1088 26243
rect 1128 26211 1160 26243
rect 1200 26211 1232 26243
rect 1272 26211 1304 26243
rect 1344 26211 1376 26243
rect 1416 26211 1448 26243
rect 1488 26211 1520 26243
rect 1560 26211 1592 26243
rect 1632 26211 1664 26243
rect 1704 26211 1736 26243
rect 1776 26211 1808 26243
rect 1848 26211 1880 26243
rect 120 26139 152 26171
rect 192 26139 224 26171
rect 264 26139 296 26171
rect 336 26139 368 26171
rect 408 26139 440 26171
rect 480 26139 512 26171
rect 552 26139 584 26171
rect 624 26139 656 26171
rect 696 26139 728 26171
rect 768 26139 800 26171
rect 840 26139 872 26171
rect 912 26139 944 26171
rect 984 26139 1016 26171
rect 1056 26139 1088 26171
rect 1128 26139 1160 26171
rect 1200 26139 1232 26171
rect 1272 26139 1304 26171
rect 1344 26139 1376 26171
rect 1416 26139 1448 26171
rect 1488 26139 1520 26171
rect 1560 26139 1592 26171
rect 1632 26139 1664 26171
rect 1704 26139 1736 26171
rect 1776 26139 1808 26171
rect 1848 26139 1880 26171
rect 120 26067 152 26099
rect 192 26067 224 26099
rect 264 26067 296 26099
rect 336 26067 368 26099
rect 408 26067 440 26099
rect 480 26067 512 26099
rect 552 26067 584 26099
rect 624 26067 656 26099
rect 696 26067 728 26099
rect 768 26067 800 26099
rect 840 26067 872 26099
rect 912 26067 944 26099
rect 984 26067 1016 26099
rect 1056 26067 1088 26099
rect 1128 26067 1160 26099
rect 1200 26067 1232 26099
rect 1272 26067 1304 26099
rect 1344 26067 1376 26099
rect 1416 26067 1448 26099
rect 1488 26067 1520 26099
rect 1560 26067 1592 26099
rect 1632 26067 1664 26099
rect 1704 26067 1736 26099
rect 1776 26067 1808 26099
rect 1848 26067 1880 26099
rect 120 25995 152 26027
rect 192 25995 224 26027
rect 264 25995 296 26027
rect 336 25995 368 26027
rect 408 25995 440 26027
rect 480 25995 512 26027
rect 552 25995 584 26027
rect 624 25995 656 26027
rect 696 25995 728 26027
rect 768 25995 800 26027
rect 840 25995 872 26027
rect 912 25995 944 26027
rect 984 25995 1016 26027
rect 1056 25995 1088 26027
rect 1128 25995 1160 26027
rect 1200 25995 1232 26027
rect 1272 25995 1304 26027
rect 1344 25995 1376 26027
rect 1416 25995 1448 26027
rect 1488 25995 1520 26027
rect 1560 25995 1592 26027
rect 1632 25995 1664 26027
rect 1704 25995 1736 26027
rect 1776 25995 1808 26027
rect 1848 25995 1880 26027
rect 120 25923 152 25955
rect 192 25923 224 25955
rect 264 25923 296 25955
rect 336 25923 368 25955
rect 408 25923 440 25955
rect 480 25923 512 25955
rect 552 25923 584 25955
rect 624 25923 656 25955
rect 696 25923 728 25955
rect 768 25923 800 25955
rect 840 25923 872 25955
rect 912 25923 944 25955
rect 984 25923 1016 25955
rect 1056 25923 1088 25955
rect 1128 25923 1160 25955
rect 1200 25923 1232 25955
rect 1272 25923 1304 25955
rect 1344 25923 1376 25955
rect 1416 25923 1448 25955
rect 1488 25923 1520 25955
rect 1560 25923 1592 25955
rect 1632 25923 1664 25955
rect 1704 25923 1736 25955
rect 1776 25923 1808 25955
rect 1848 25923 1880 25955
rect 120 25851 152 25883
rect 192 25851 224 25883
rect 264 25851 296 25883
rect 336 25851 368 25883
rect 408 25851 440 25883
rect 480 25851 512 25883
rect 552 25851 584 25883
rect 624 25851 656 25883
rect 696 25851 728 25883
rect 768 25851 800 25883
rect 840 25851 872 25883
rect 912 25851 944 25883
rect 984 25851 1016 25883
rect 1056 25851 1088 25883
rect 1128 25851 1160 25883
rect 1200 25851 1232 25883
rect 1272 25851 1304 25883
rect 1344 25851 1376 25883
rect 1416 25851 1448 25883
rect 1488 25851 1520 25883
rect 1560 25851 1592 25883
rect 1632 25851 1664 25883
rect 1704 25851 1736 25883
rect 1776 25851 1808 25883
rect 1848 25851 1880 25883
rect 120 25779 152 25811
rect 192 25779 224 25811
rect 264 25779 296 25811
rect 336 25779 368 25811
rect 408 25779 440 25811
rect 480 25779 512 25811
rect 552 25779 584 25811
rect 624 25779 656 25811
rect 696 25779 728 25811
rect 768 25779 800 25811
rect 840 25779 872 25811
rect 912 25779 944 25811
rect 984 25779 1016 25811
rect 1056 25779 1088 25811
rect 1128 25779 1160 25811
rect 1200 25779 1232 25811
rect 1272 25779 1304 25811
rect 1344 25779 1376 25811
rect 1416 25779 1448 25811
rect 1488 25779 1520 25811
rect 1560 25779 1592 25811
rect 1632 25779 1664 25811
rect 1704 25779 1736 25811
rect 1776 25779 1808 25811
rect 1848 25779 1880 25811
rect 120 25707 152 25739
rect 192 25707 224 25739
rect 264 25707 296 25739
rect 336 25707 368 25739
rect 408 25707 440 25739
rect 480 25707 512 25739
rect 552 25707 584 25739
rect 624 25707 656 25739
rect 696 25707 728 25739
rect 768 25707 800 25739
rect 840 25707 872 25739
rect 912 25707 944 25739
rect 984 25707 1016 25739
rect 1056 25707 1088 25739
rect 1128 25707 1160 25739
rect 1200 25707 1232 25739
rect 1272 25707 1304 25739
rect 1344 25707 1376 25739
rect 1416 25707 1448 25739
rect 1488 25707 1520 25739
rect 1560 25707 1592 25739
rect 1632 25707 1664 25739
rect 1704 25707 1736 25739
rect 1776 25707 1808 25739
rect 1848 25707 1880 25739
rect 120 25635 152 25667
rect 192 25635 224 25667
rect 264 25635 296 25667
rect 336 25635 368 25667
rect 408 25635 440 25667
rect 480 25635 512 25667
rect 552 25635 584 25667
rect 624 25635 656 25667
rect 696 25635 728 25667
rect 768 25635 800 25667
rect 840 25635 872 25667
rect 912 25635 944 25667
rect 984 25635 1016 25667
rect 1056 25635 1088 25667
rect 1128 25635 1160 25667
rect 1200 25635 1232 25667
rect 1272 25635 1304 25667
rect 1344 25635 1376 25667
rect 1416 25635 1448 25667
rect 1488 25635 1520 25667
rect 1560 25635 1592 25667
rect 1632 25635 1664 25667
rect 1704 25635 1736 25667
rect 1776 25635 1808 25667
rect 1848 25635 1880 25667
rect 120 25563 152 25595
rect 192 25563 224 25595
rect 264 25563 296 25595
rect 336 25563 368 25595
rect 408 25563 440 25595
rect 480 25563 512 25595
rect 552 25563 584 25595
rect 624 25563 656 25595
rect 696 25563 728 25595
rect 768 25563 800 25595
rect 840 25563 872 25595
rect 912 25563 944 25595
rect 984 25563 1016 25595
rect 1056 25563 1088 25595
rect 1128 25563 1160 25595
rect 1200 25563 1232 25595
rect 1272 25563 1304 25595
rect 1344 25563 1376 25595
rect 1416 25563 1448 25595
rect 1488 25563 1520 25595
rect 1560 25563 1592 25595
rect 1632 25563 1664 25595
rect 1704 25563 1736 25595
rect 1776 25563 1808 25595
rect 1848 25563 1880 25595
rect 120 25491 152 25523
rect 192 25491 224 25523
rect 264 25491 296 25523
rect 336 25491 368 25523
rect 408 25491 440 25523
rect 480 25491 512 25523
rect 552 25491 584 25523
rect 624 25491 656 25523
rect 696 25491 728 25523
rect 768 25491 800 25523
rect 840 25491 872 25523
rect 912 25491 944 25523
rect 984 25491 1016 25523
rect 1056 25491 1088 25523
rect 1128 25491 1160 25523
rect 1200 25491 1232 25523
rect 1272 25491 1304 25523
rect 1344 25491 1376 25523
rect 1416 25491 1448 25523
rect 1488 25491 1520 25523
rect 1560 25491 1592 25523
rect 1632 25491 1664 25523
rect 1704 25491 1736 25523
rect 1776 25491 1808 25523
rect 1848 25491 1880 25523
rect 120 25419 152 25451
rect 192 25419 224 25451
rect 264 25419 296 25451
rect 336 25419 368 25451
rect 408 25419 440 25451
rect 480 25419 512 25451
rect 552 25419 584 25451
rect 624 25419 656 25451
rect 696 25419 728 25451
rect 768 25419 800 25451
rect 840 25419 872 25451
rect 912 25419 944 25451
rect 984 25419 1016 25451
rect 1056 25419 1088 25451
rect 1128 25419 1160 25451
rect 1200 25419 1232 25451
rect 1272 25419 1304 25451
rect 1344 25419 1376 25451
rect 1416 25419 1448 25451
rect 1488 25419 1520 25451
rect 1560 25419 1592 25451
rect 1632 25419 1664 25451
rect 1704 25419 1736 25451
rect 1776 25419 1808 25451
rect 1848 25419 1880 25451
rect 120 25347 152 25379
rect 192 25347 224 25379
rect 264 25347 296 25379
rect 336 25347 368 25379
rect 408 25347 440 25379
rect 480 25347 512 25379
rect 552 25347 584 25379
rect 624 25347 656 25379
rect 696 25347 728 25379
rect 768 25347 800 25379
rect 840 25347 872 25379
rect 912 25347 944 25379
rect 984 25347 1016 25379
rect 1056 25347 1088 25379
rect 1128 25347 1160 25379
rect 1200 25347 1232 25379
rect 1272 25347 1304 25379
rect 1344 25347 1376 25379
rect 1416 25347 1448 25379
rect 1488 25347 1520 25379
rect 1560 25347 1592 25379
rect 1632 25347 1664 25379
rect 1704 25347 1736 25379
rect 1776 25347 1808 25379
rect 1848 25347 1880 25379
rect 120 25275 152 25307
rect 192 25275 224 25307
rect 264 25275 296 25307
rect 336 25275 368 25307
rect 408 25275 440 25307
rect 480 25275 512 25307
rect 552 25275 584 25307
rect 624 25275 656 25307
rect 696 25275 728 25307
rect 768 25275 800 25307
rect 840 25275 872 25307
rect 912 25275 944 25307
rect 984 25275 1016 25307
rect 1056 25275 1088 25307
rect 1128 25275 1160 25307
rect 1200 25275 1232 25307
rect 1272 25275 1304 25307
rect 1344 25275 1376 25307
rect 1416 25275 1448 25307
rect 1488 25275 1520 25307
rect 1560 25275 1592 25307
rect 1632 25275 1664 25307
rect 1704 25275 1736 25307
rect 1776 25275 1808 25307
rect 1848 25275 1880 25307
rect 120 25203 152 25235
rect 192 25203 224 25235
rect 264 25203 296 25235
rect 336 25203 368 25235
rect 408 25203 440 25235
rect 480 25203 512 25235
rect 552 25203 584 25235
rect 624 25203 656 25235
rect 696 25203 728 25235
rect 768 25203 800 25235
rect 840 25203 872 25235
rect 912 25203 944 25235
rect 984 25203 1016 25235
rect 1056 25203 1088 25235
rect 1128 25203 1160 25235
rect 1200 25203 1232 25235
rect 1272 25203 1304 25235
rect 1344 25203 1376 25235
rect 1416 25203 1448 25235
rect 1488 25203 1520 25235
rect 1560 25203 1592 25235
rect 1632 25203 1664 25235
rect 1704 25203 1736 25235
rect 1776 25203 1808 25235
rect 1848 25203 1880 25235
rect 120 25131 152 25163
rect 192 25131 224 25163
rect 264 25131 296 25163
rect 336 25131 368 25163
rect 408 25131 440 25163
rect 480 25131 512 25163
rect 552 25131 584 25163
rect 624 25131 656 25163
rect 696 25131 728 25163
rect 768 25131 800 25163
rect 840 25131 872 25163
rect 912 25131 944 25163
rect 984 25131 1016 25163
rect 1056 25131 1088 25163
rect 1128 25131 1160 25163
rect 1200 25131 1232 25163
rect 1272 25131 1304 25163
rect 1344 25131 1376 25163
rect 1416 25131 1448 25163
rect 1488 25131 1520 25163
rect 1560 25131 1592 25163
rect 1632 25131 1664 25163
rect 1704 25131 1736 25163
rect 1776 25131 1808 25163
rect 1848 25131 1880 25163
rect 120 25059 152 25091
rect 192 25059 224 25091
rect 264 25059 296 25091
rect 336 25059 368 25091
rect 408 25059 440 25091
rect 480 25059 512 25091
rect 552 25059 584 25091
rect 624 25059 656 25091
rect 696 25059 728 25091
rect 768 25059 800 25091
rect 840 25059 872 25091
rect 912 25059 944 25091
rect 984 25059 1016 25091
rect 1056 25059 1088 25091
rect 1128 25059 1160 25091
rect 1200 25059 1232 25091
rect 1272 25059 1304 25091
rect 1344 25059 1376 25091
rect 1416 25059 1448 25091
rect 1488 25059 1520 25091
rect 1560 25059 1592 25091
rect 1632 25059 1664 25091
rect 1704 25059 1736 25091
rect 1776 25059 1808 25091
rect 1848 25059 1880 25091
rect 120 24987 152 25019
rect 192 24987 224 25019
rect 264 24987 296 25019
rect 336 24987 368 25019
rect 408 24987 440 25019
rect 480 24987 512 25019
rect 552 24987 584 25019
rect 624 24987 656 25019
rect 696 24987 728 25019
rect 768 24987 800 25019
rect 840 24987 872 25019
rect 912 24987 944 25019
rect 984 24987 1016 25019
rect 1056 24987 1088 25019
rect 1128 24987 1160 25019
rect 1200 24987 1232 25019
rect 1272 24987 1304 25019
rect 1344 24987 1376 25019
rect 1416 24987 1448 25019
rect 1488 24987 1520 25019
rect 1560 24987 1592 25019
rect 1632 24987 1664 25019
rect 1704 24987 1736 25019
rect 1776 24987 1808 25019
rect 1848 24987 1880 25019
rect 120 24915 152 24947
rect 192 24915 224 24947
rect 264 24915 296 24947
rect 336 24915 368 24947
rect 408 24915 440 24947
rect 480 24915 512 24947
rect 552 24915 584 24947
rect 624 24915 656 24947
rect 696 24915 728 24947
rect 768 24915 800 24947
rect 840 24915 872 24947
rect 912 24915 944 24947
rect 984 24915 1016 24947
rect 1056 24915 1088 24947
rect 1128 24915 1160 24947
rect 1200 24915 1232 24947
rect 1272 24915 1304 24947
rect 1344 24915 1376 24947
rect 1416 24915 1448 24947
rect 1488 24915 1520 24947
rect 1560 24915 1592 24947
rect 1632 24915 1664 24947
rect 1704 24915 1736 24947
rect 1776 24915 1808 24947
rect 1848 24915 1880 24947
rect 120 24843 152 24875
rect 192 24843 224 24875
rect 264 24843 296 24875
rect 336 24843 368 24875
rect 408 24843 440 24875
rect 480 24843 512 24875
rect 552 24843 584 24875
rect 624 24843 656 24875
rect 696 24843 728 24875
rect 768 24843 800 24875
rect 840 24843 872 24875
rect 912 24843 944 24875
rect 984 24843 1016 24875
rect 1056 24843 1088 24875
rect 1128 24843 1160 24875
rect 1200 24843 1232 24875
rect 1272 24843 1304 24875
rect 1344 24843 1376 24875
rect 1416 24843 1448 24875
rect 1488 24843 1520 24875
rect 1560 24843 1592 24875
rect 1632 24843 1664 24875
rect 1704 24843 1736 24875
rect 1776 24843 1808 24875
rect 1848 24843 1880 24875
rect 120 24771 152 24803
rect 192 24771 224 24803
rect 264 24771 296 24803
rect 336 24771 368 24803
rect 408 24771 440 24803
rect 480 24771 512 24803
rect 552 24771 584 24803
rect 624 24771 656 24803
rect 696 24771 728 24803
rect 768 24771 800 24803
rect 840 24771 872 24803
rect 912 24771 944 24803
rect 984 24771 1016 24803
rect 1056 24771 1088 24803
rect 1128 24771 1160 24803
rect 1200 24771 1232 24803
rect 1272 24771 1304 24803
rect 1344 24771 1376 24803
rect 1416 24771 1448 24803
rect 1488 24771 1520 24803
rect 1560 24771 1592 24803
rect 1632 24771 1664 24803
rect 1704 24771 1736 24803
rect 1776 24771 1808 24803
rect 1848 24771 1880 24803
rect 120 24699 152 24731
rect 192 24699 224 24731
rect 264 24699 296 24731
rect 336 24699 368 24731
rect 408 24699 440 24731
rect 480 24699 512 24731
rect 552 24699 584 24731
rect 624 24699 656 24731
rect 696 24699 728 24731
rect 768 24699 800 24731
rect 840 24699 872 24731
rect 912 24699 944 24731
rect 984 24699 1016 24731
rect 1056 24699 1088 24731
rect 1128 24699 1160 24731
rect 1200 24699 1232 24731
rect 1272 24699 1304 24731
rect 1344 24699 1376 24731
rect 1416 24699 1448 24731
rect 1488 24699 1520 24731
rect 1560 24699 1592 24731
rect 1632 24699 1664 24731
rect 1704 24699 1736 24731
rect 1776 24699 1808 24731
rect 1848 24699 1880 24731
rect 120 24627 152 24659
rect 192 24627 224 24659
rect 264 24627 296 24659
rect 336 24627 368 24659
rect 408 24627 440 24659
rect 480 24627 512 24659
rect 552 24627 584 24659
rect 624 24627 656 24659
rect 696 24627 728 24659
rect 768 24627 800 24659
rect 840 24627 872 24659
rect 912 24627 944 24659
rect 984 24627 1016 24659
rect 1056 24627 1088 24659
rect 1128 24627 1160 24659
rect 1200 24627 1232 24659
rect 1272 24627 1304 24659
rect 1344 24627 1376 24659
rect 1416 24627 1448 24659
rect 1488 24627 1520 24659
rect 1560 24627 1592 24659
rect 1632 24627 1664 24659
rect 1704 24627 1736 24659
rect 1776 24627 1808 24659
rect 1848 24627 1880 24659
rect 120 24555 152 24587
rect 192 24555 224 24587
rect 264 24555 296 24587
rect 336 24555 368 24587
rect 408 24555 440 24587
rect 480 24555 512 24587
rect 552 24555 584 24587
rect 624 24555 656 24587
rect 696 24555 728 24587
rect 768 24555 800 24587
rect 840 24555 872 24587
rect 912 24555 944 24587
rect 984 24555 1016 24587
rect 1056 24555 1088 24587
rect 1128 24555 1160 24587
rect 1200 24555 1232 24587
rect 1272 24555 1304 24587
rect 1344 24555 1376 24587
rect 1416 24555 1448 24587
rect 1488 24555 1520 24587
rect 1560 24555 1592 24587
rect 1632 24555 1664 24587
rect 1704 24555 1736 24587
rect 1776 24555 1808 24587
rect 1848 24555 1880 24587
rect 120 24483 152 24515
rect 192 24483 224 24515
rect 264 24483 296 24515
rect 336 24483 368 24515
rect 408 24483 440 24515
rect 480 24483 512 24515
rect 552 24483 584 24515
rect 624 24483 656 24515
rect 696 24483 728 24515
rect 768 24483 800 24515
rect 840 24483 872 24515
rect 912 24483 944 24515
rect 984 24483 1016 24515
rect 1056 24483 1088 24515
rect 1128 24483 1160 24515
rect 1200 24483 1232 24515
rect 1272 24483 1304 24515
rect 1344 24483 1376 24515
rect 1416 24483 1448 24515
rect 1488 24483 1520 24515
rect 1560 24483 1592 24515
rect 1632 24483 1664 24515
rect 1704 24483 1736 24515
rect 1776 24483 1808 24515
rect 1848 24483 1880 24515
rect 120 24411 152 24443
rect 192 24411 224 24443
rect 264 24411 296 24443
rect 336 24411 368 24443
rect 408 24411 440 24443
rect 480 24411 512 24443
rect 552 24411 584 24443
rect 624 24411 656 24443
rect 696 24411 728 24443
rect 768 24411 800 24443
rect 840 24411 872 24443
rect 912 24411 944 24443
rect 984 24411 1016 24443
rect 1056 24411 1088 24443
rect 1128 24411 1160 24443
rect 1200 24411 1232 24443
rect 1272 24411 1304 24443
rect 1344 24411 1376 24443
rect 1416 24411 1448 24443
rect 1488 24411 1520 24443
rect 1560 24411 1592 24443
rect 1632 24411 1664 24443
rect 1704 24411 1736 24443
rect 1776 24411 1808 24443
rect 1848 24411 1880 24443
rect 120 24339 152 24371
rect 192 24339 224 24371
rect 264 24339 296 24371
rect 336 24339 368 24371
rect 408 24339 440 24371
rect 480 24339 512 24371
rect 552 24339 584 24371
rect 624 24339 656 24371
rect 696 24339 728 24371
rect 768 24339 800 24371
rect 840 24339 872 24371
rect 912 24339 944 24371
rect 984 24339 1016 24371
rect 1056 24339 1088 24371
rect 1128 24339 1160 24371
rect 1200 24339 1232 24371
rect 1272 24339 1304 24371
rect 1344 24339 1376 24371
rect 1416 24339 1448 24371
rect 1488 24339 1520 24371
rect 1560 24339 1592 24371
rect 1632 24339 1664 24371
rect 1704 24339 1736 24371
rect 1776 24339 1808 24371
rect 1848 24339 1880 24371
rect 120 24267 152 24299
rect 192 24267 224 24299
rect 264 24267 296 24299
rect 336 24267 368 24299
rect 408 24267 440 24299
rect 480 24267 512 24299
rect 552 24267 584 24299
rect 624 24267 656 24299
rect 696 24267 728 24299
rect 768 24267 800 24299
rect 840 24267 872 24299
rect 912 24267 944 24299
rect 984 24267 1016 24299
rect 1056 24267 1088 24299
rect 1128 24267 1160 24299
rect 1200 24267 1232 24299
rect 1272 24267 1304 24299
rect 1344 24267 1376 24299
rect 1416 24267 1448 24299
rect 1488 24267 1520 24299
rect 1560 24267 1592 24299
rect 1632 24267 1664 24299
rect 1704 24267 1736 24299
rect 1776 24267 1808 24299
rect 1848 24267 1880 24299
rect 120 24195 152 24227
rect 192 24195 224 24227
rect 264 24195 296 24227
rect 336 24195 368 24227
rect 408 24195 440 24227
rect 480 24195 512 24227
rect 552 24195 584 24227
rect 624 24195 656 24227
rect 696 24195 728 24227
rect 768 24195 800 24227
rect 840 24195 872 24227
rect 912 24195 944 24227
rect 984 24195 1016 24227
rect 1056 24195 1088 24227
rect 1128 24195 1160 24227
rect 1200 24195 1232 24227
rect 1272 24195 1304 24227
rect 1344 24195 1376 24227
rect 1416 24195 1448 24227
rect 1488 24195 1520 24227
rect 1560 24195 1592 24227
rect 1632 24195 1664 24227
rect 1704 24195 1736 24227
rect 1776 24195 1808 24227
rect 1848 24195 1880 24227
rect 120 24123 152 24155
rect 192 24123 224 24155
rect 264 24123 296 24155
rect 336 24123 368 24155
rect 408 24123 440 24155
rect 480 24123 512 24155
rect 552 24123 584 24155
rect 624 24123 656 24155
rect 696 24123 728 24155
rect 768 24123 800 24155
rect 840 24123 872 24155
rect 912 24123 944 24155
rect 984 24123 1016 24155
rect 1056 24123 1088 24155
rect 1128 24123 1160 24155
rect 1200 24123 1232 24155
rect 1272 24123 1304 24155
rect 1344 24123 1376 24155
rect 1416 24123 1448 24155
rect 1488 24123 1520 24155
rect 1560 24123 1592 24155
rect 1632 24123 1664 24155
rect 1704 24123 1736 24155
rect 1776 24123 1808 24155
rect 1848 24123 1880 24155
rect 120 24051 152 24083
rect 192 24051 224 24083
rect 264 24051 296 24083
rect 336 24051 368 24083
rect 408 24051 440 24083
rect 480 24051 512 24083
rect 552 24051 584 24083
rect 624 24051 656 24083
rect 696 24051 728 24083
rect 768 24051 800 24083
rect 840 24051 872 24083
rect 912 24051 944 24083
rect 984 24051 1016 24083
rect 1056 24051 1088 24083
rect 1128 24051 1160 24083
rect 1200 24051 1232 24083
rect 1272 24051 1304 24083
rect 1344 24051 1376 24083
rect 1416 24051 1448 24083
rect 1488 24051 1520 24083
rect 1560 24051 1592 24083
rect 1632 24051 1664 24083
rect 1704 24051 1736 24083
rect 1776 24051 1808 24083
rect 1848 24051 1880 24083
rect 120 23979 152 24011
rect 192 23979 224 24011
rect 264 23979 296 24011
rect 336 23979 368 24011
rect 408 23979 440 24011
rect 480 23979 512 24011
rect 552 23979 584 24011
rect 624 23979 656 24011
rect 696 23979 728 24011
rect 768 23979 800 24011
rect 840 23979 872 24011
rect 912 23979 944 24011
rect 984 23979 1016 24011
rect 1056 23979 1088 24011
rect 1128 23979 1160 24011
rect 1200 23979 1232 24011
rect 1272 23979 1304 24011
rect 1344 23979 1376 24011
rect 1416 23979 1448 24011
rect 1488 23979 1520 24011
rect 1560 23979 1592 24011
rect 1632 23979 1664 24011
rect 1704 23979 1736 24011
rect 1776 23979 1808 24011
rect 1848 23979 1880 24011
rect 120 23907 152 23939
rect 192 23907 224 23939
rect 264 23907 296 23939
rect 336 23907 368 23939
rect 408 23907 440 23939
rect 480 23907 512 23939
rect 552 23907 584 23939
rect 624 23907 656 23939
rect 696 23907 728 23939
rect 768 23907 800 23939
rect 840 23907 872 23939
rect 912 23907 944 23939
rect 984 23907 1016 23939
rect 1056 23907 1088 23939
rect 1128 23907 1160 23939
rect 1200 23907 1232 23939
rect 1272 23907 1304 23939
rect 1344 23907 1376 23939
rect 1416 23907 1448 23939
rect 1488 23907 1520 23939
rect 1560 23907 1592 23939
rect 1632 23907 1664 23939
rect 1704 23907 1736 23939
rect 1776 23907 1808 23939
rect 1848 23907 1880 23939
rect 120 23835 152 23867
rect 192 23835 224 23867
rect 264 23835 296 23867
rect 336 23835 368 23867
rect 408 23835 440 23867
rect 480 23835 512 23867
rect 552 23835 584 23867
rect 624 23835 656 23867
rect 696 23835 728 23867
rect 768 23835 800 23867
rect 840 23835 872 23867
rect 912 23835 944 23867
rect 984 23835 1016 23867
rect 1056 23835 1088 23867
rect 1128 23835 1160 23867
rect 1200 23835 1232 23867
rect 1272 23835 1304 23867
rect 1344 23835 1376 23867
rect 1416 23835 1448 23867
rect 1488 23835 1520 23867
rect 1560 23835 1592 23867
rect 1632 23835 1664 23867
rect 1704 23835 1736 23867
rect 1776 23835 1808 23867
rect 1848 23835 1880 23867
rect 120 23763 152 23795
rect 192 23763 224 23795
rect 264 23763 296 23795
rect 336 23763 368 23795
rect 408 23763 440 23795
rect 480 23763 512 23795
rect 552 23763 584 23795
rect 624 23763 656 23795
rect 696 23763 728 23795
rect 768 23763 800 23795
rect 840 23763 872 23795
rect 912 23763 944 23795
rect 984 23763 1016 23795
rect 1056 23763 1088 23795
rect 1128 23763 1160 23795
rect 1200 23763 1232 23795
rect 1272 23763 1304 23795
rect 1344 23763 1376 23795
rect 1416 23763 1448 23795
rect 1488 23763 1520 23795
rect 1560 23763 1592 23795
rect 1632 23763 1664 23795
rect 1704 23763 1736 23795
rect 1776 23763 1808 23795
rect 1848 23763 1880 23795
rect 120 23691 152 23723
rect 192 23691 224 23723
rect 264 23691 296 23723
rect 336 23691 368 23723
rect 408 23691 440 23723
rect 480 23691 512 23723
rect 552 23691 584 23723
rect 624 23691 656 23723
rect 696 23691 728 23723
rect 768 23691 800 23723
rect 840 23691 872 23723
rect 912 23691 944 23723
rect 984 23691 1016 23723
rect 1056 23691 1088 23723
rect 1128 23691 1160 23723
rect 1200 23691 1232 23723
rect 1272 23691 1304 23723
rect 1344 23691 1376 23723
rect 1416 23691 1448 23723
rect 1488 23691 1520 23723
rect 1560 23691 1592 23723
rect 1632 23691 1664 23723
rect 1704 23691 1736 23723
rect 1776 23691 1808 23723
rect 1848 23691 1880 23723
rect 120 23619 152 23651
rect 192 23619 224 23651
rect 264 23619 296 23651
rect 336 23619 368 23651
rect 408 23619 440 23651
rect 480 23619 512 23651
rect 552 23619 584 23651
rect 624 23619 656 23651
rect 696 23619 728 23651
rect 768 23619 800 23651
rect 840 23619 872 23651
rect 912 23619 944 23651
rect 984 23619 1016 23651
rect 1056 23619 1088 23651
rect 1128 23619 1160 23651
rect 1200 23619 1232 23651
rect 1272 23619 1304 23651
rect 1344 23619 1376 23651
rect 1416 23619 1448 23651
rect 1488 23619 1520 23651
rect 1560 23619 1592 23651
rect 1632 23619 1664 23651
rect 1704 23619 1736 23651
rect 1776 23619 1808 23651
rect 1848 23619 1880 23651
rect 120 23547 152 23579
rect 192 23547 224 23579
rect 264 23547 296 23579
rect 336 23547 368 23579
rect 408 23547 440 23579
rect 480 23547 512 23579
rect 552 23547 584 23579
rect 624 23547 656 23579
rect 696 23547 728 23579
rect 768 23547 800 23579
rect 840 23547 872 23579
rect 912 23547 944 23579
rect 984 23547 1016 23579
rect 1056 23547 1088 23579
rect 1128 23547 1160 23579
rect 1200 23547 1232 23579
rect 1272 23547 1304 23579
rect 1344 23547 1376 23579
rect 1416 23547 1448 23579
rect 1488 23547 1520 23579
rect 1560 23547 1592 23579
rect 1632 23547 1664 23579
rect 1704 23547 1736 23579
rect 1776 23547 1808 23579
rect 1848 23547 1880 23579
rect 120 23475 152 23507
rect 192 23475 224 23507
rect 264 23475 296 23507
rect 336 23475 368 23507
rect 408 23475 440 23507
rect 480 23475 512 23507
rect 552 23475 584 23507
rect 624 23475 656 23507
rect 696 23475 728 23507
rect 768 23475 800 23507
rect 840 23475 872 23507
rect 912 23475 944 23507
rect 984 23475 1016 23507
rect 1056 23475 1088 23507
rect 1128 23475 1160 23507
rect 1200 23475 1232 23507
rect 1272 23475 1304 23507
rect 1344 23475 1376 23507
rect 1416 23475 1448 23507
rect 1488 23475 1520 23507
rect 1560 23475 1592 23507
rect 1632 23475 1664 23507
rect 1704 23475 1736 23507
rect 1776 23475 1808 23507
rect 1848 23475 1880 23507
rect 120 23403 152 23435
rect 192 23403 224 23435
rect 264 23403 296 23435
rect 336 23403 368 23435
rect 408 23403 440 23435
rect 480 23403 512 23435
rect 552 23403 584 23435
rect 624 23403 656 23435
rect 696 23403 728 23435
rect 768 23403 800 23435
rect 840 23403 872 23435
rect 912 23403 944 23435
rect 984 23403 1016 23435
rect 1056 23403 1088 23435
rect 1128 23403 1160 23435
rect 1200 23403 1232 23435
rect 1272 23403 1304 23435
rect 1344 23403 1376 23435
rect 1416 23403 1448 23435
rect 1488 23403 1520 23435
rect 1560 23403 1592 23435
rect 1632 23403 1664 23435
rect 1704 23403 1736 23435
rect 1776 23403 1808 23435
rect 1848 23403 1880 23435
rect 120 23331 152 23363
rect 192 23331 224 23363
rect 264 23331 296 23363
rect 336 23331 368 23363
rect 408 23331 440 23363
rect 480 23331 512 23363
rect 552 23331 584 23363
rect 624 23331 656 23363
rect 696 23331 728 23363
rect 768 23331 800 23363
rect 840 23331 872 23363
rect 912 23331 944 23363
rect 984 23331 1016 23363
rect 1056 23331 1088 23363
rect 1128 23331 1160 23363
rect 1200 23331 1232 23363
rect 1272 23331 1304 23363
rect 1344 23331 1376 23363
rect 1416 23331 1448 23363
rect 1488 23331 1520 23363
rect 1560 23331 1592 23363
rect 1632 23331 1664 23363
rect 1704 23331 1736 23363
rect 1776 23331 1808 23363
rect 1848 23331 1880 23363
rect 120 23259 152 23291
rect 192 23259 224 23291
rect 264 23259 296 23291
rect 336 23259 368 23291
rect 408 23259 440 23291
rect 480 23259 512 23291
rect 552 23259 584 23291
rect 624 23259 656 23291
rect 696 23259 728 23291
rect 768 23259 800 23291
rect 840 23259 872 23291
rect 912 23259 944 23291
rect 984 23259 1016 23291
rect 1056 23259 1088 23291
rect 1128 23259 1160 23291
rect 1200 23259 1232 23291
rect 1272 23259 1304 23291
rect 1344 23259 1376 23291
rect 1416 23259 1448 23291
rect 1488 23259 1520 23291
rect 1560 23259 1592 23291
rect 1632 23259 1664 23291
rect 1704 23259 1736 23291
rect 1776 23259 1808 23291
rect 1848 23259 1880 23291
rect 120 23187 152 23219
rect 192 23187 224 23219
rect 264 23187 296 23219
rect 336 23187 368 23219
rect 408 23187 440 23219
rect 480 23187 512 23219
rect 552 23187 584 23219
rect 624 23187 656 23219
rect 696 23187 728 23219
rect 768 23187 800 23219
rect 840 23187 872 23219
rect 912 23187 944 23219
rect 984 23187 1016 23219
rect 1056 23187 1088 23219
rect 1128 23187 1160 23219
rect 1200 23187 1232 23219
rect 1272 23187 1304 23219
rect 1344 23187 1376 23219
rect 1416 23187 1448 23219
rect 1488 23187 1520 23219
rect 1560 23187 1592 23219
rect 1632 23187 1664 23219
rect 1704 23187 1736 23219
rect 1776 23187 1808 23219
rect 1848 23187 1880 23219
rect 192 22842 224 22874
rect 264 22842 296 22874
rect 336 22842 368 22874
rect 408 22842 440 22874
rect 480 22842 512 22874
rect 552 22842 584 22874
rect 624 22842 656 22874
rect 696 22842 728 22874
rect 768 22842 800 22874
rect 840 22842 872 22874
rect 912 22842 944 22874
rect 984 22842 1016 22874
rect 1056 22842 1088 22874
rect 1128 22842 1160 22874
rect 1200 22842 1232 22874
rect 1272 22842 1304 22874
rect 1344 22842 1376 22874
rect 1416 22842 1448 22874
rect 1488 22842 1520 22874
rect 1560 22842 1592 22874
rect 1632 22842 1664 22874
rect 1704 22842 1736 22874
rect 1776 22842 1808 22874
rect 1848 22842 1880 22874
rect 120 22770 152 22802
rect 192 22770 224 22802
rect 264 22770 296 22802
rect 336 22770 368 22802
rect 408 22770 440 22802
rect 480 22770 512 22802
rect 552 22770 584 22802
rect 624 22770 656 22802
rect 696 22770 728 22802
rect 768 22770 800 22802
rect 840 22770 872 22802
rect 912 22770 944 22802
rect 984 22770 1016 22802
rect 1056 22770 1088 22802
rect 1128 22770 1160 22802
rect 1200 22770 1232 22802
rect 1272 22770 1304 22802
rect 1344 22770 1376 22802
rect 1416 22770 1448 22802
rect 1488 22770 1520 22802
rect 1560 22770 1592 22802
rect 1632 22770 1664 22802
rect 1704 22770 1736 22802
rect 1776 22770 1808 22802
rect 1848 22770 1880 22802
rect 120 22698 152 22730
rect 192 22698 224 22730
rect 264 22698 296 22730
rect 336 22698 368 22730
rect 408 22698 440 22730
rect 480 22698 512 22730
rect 552 22698 584 22730
rect 624 22698 656 22730
rect 696 22698 728 22730
rect 768 22698 800 22730
rect 840 22698 872 22730
rect 912 22698 944 22730
rect 984 22698 1016 22730
rect 1056 22698 1088 22730
rect 1128 22698 1160 22730
rect 1200 22698 1232 22730
rect 1272 22698 1304 22730
rect 1344 22698 1376 22730
rect 1416 22698 1448 22730
rect 1488 22698 1520 22730
rect 1560 22698 1592 22730
rect 1632 22698 1664 22730
rect 1704 22698 1736 22730
rect 1776 22698 1808 22730
rect 1848 22698 1880 22730
rect 120 22626 152 22658
rect 192 22626 224 22658
rect 264 22626 296 22658
rect 336 22626 368 22658
rect 408 22626 440 22658
rect 480 22626 512 22658
rect 552 22626 584 22658
rect 624 22626 656 22658
rect 696 22626 728 22658
rect 768 22626 800 22658
rect 840 22626 872 22658
rect 912 22626 944 22658
rect 984 22626 1016 22658
rect 1056 22626 1088 22658
rect 1128 22626 1160 22658
rect 1200 22626 1232 22658
rect 1272 22626 1304 22658
rect 1344 22626 1376 22658
rect 1416 22626 1448 22658
rect 1488 22626 1520 22658
rect 1560 22626 1592 22658
rect 1632 22626 1664 22658
rect 1704 22626 1736 22658
rect 1776 22626 1808 22658
rect 1848 22626 1880 22658
rect 120 22554 152 22586
rect 192 22554 224 22586
rect 264 22554 296 22586
rect 336 22554 368 22586
rect 408 22554 440 22586
rect 480 22554 512 22586
rect 552 22554 584 22586
rect 624 22554 656 22586
rect 696 22554 728 22586
rect 768 22554 800 22586
rect 840 22554 872 22586
rect 912 22554 944 22586
rect 984 22554 1016 22586
rect 1056 22554 1088 22586
rect 1128 22554 1160 22586
rect 1200 22554 1232 22586
rect 1272 22554 1304 22586
rect 1344 22554 1376 22586
rect 1416 22554 1448 22586
rect 1488 22554 1520 22586
rect 1560 22554 1592 22586
rect 1632 22554 1664 22586
rect 1704 22554 1736 22586
rect 1776 22554 1808 22586
rect 1848 22554 1880 22586
rect 120 22482 152 22514
rect 192 22482 224 22514
rect 264 22482 296 22514
rect 336 22482 368 22514
rect 408 22482 440 22514
rect 480 22482 512 22514
rect 552 22482 584 22514
rect 624 22482 656 22514
rect 696 22482 728 22514
rect 768 22482 800 22514
rect 840 22482 872 22514
rect 912 22482 944 22514
rect 984 22482 1016 22514
rect 1056 22482 1088 22514
rect 1128 22482 1160 22514
rect 1200 22482 1232 22514
rect 1272 22482 1304 22514
rect 1344 22482 1376 22514
rect 1416 22482 1448 22514
rect 1488 22482 1520 22514
rect 1560 22482 1592 22514
rect 1632 22482 1664 22514
rect 1704 22482 1736 22514
rect 1776 22482 1808 22514
rect 1848 22482 1880 22514
rect 120 22410 152 22442
rect 192 22410 224 22442
rect 264 22410 296 22442
rect 336 22410 368 22442
rect 408 22410 440 22442
rect 480 22410 512 22442
rect 552 22410 584 22442
rect 624 22410 656 22442
rect 696 22410 728 22442
rect 768 22410 800 22442
rect 840 22410 872 22442
rect 912 22410 944 22442
rect 984 22410 1016 22442
rect 1056 22410 1088 22442
rect 1128 22410 1160 22442
rect 1200 22410 1232 22442
rect 1272 22410 1304 22442
rect 1344 22410 1376 22442
rect 1416 22410 1448 22442
rect 1488 22410 1520 22442
rect 1560 22410 1592 22442
rect 1632 22410 1664 22442
rect 1704 22410 1736 22442
rect 1776 22410 1808 22442
rect 1848 22410 1880 22442
rect 120 22338 152 22370
rect 192 22338 224 22370
rect 264 22338 296 22370
rect 336 22338 368 22370
rect 408 22338 440 22370
rect 480 22338 512 22370
rect 552 22338 584 22370
rect 624 22338 656 22370
rect 696 22338 728 22370
rect 768 22338 800 22370
rect 840 22338 872 22370
rect 912 22338 944 22370
rect 984 22338 1016 22370
rect 1056 22338 1088 22370
rect 1128 22338 1160 22370
rect 1200 22338 1232 22370
rect 1272 22338 1304 22370
rect 1344 22338 1376 22370
rect 1416 22338 1448 22370
rect 1488 22338 1520 22370
rect 1560 22338 1592 22370
rect 1632 22338 1664 22370
rect 1704 22338 1736 22370
rect 1776 22338 1808 22370
rect 1848 22338 1880 22370
rect 120 22266 152 22298
rect 192 22266 224 22298
rect 264 22266 296 22298
rect 336 22266 368 22298
rect 408 22266 440 22298
rect 480 22266 512 22298
rect 552 22266 584 22298
rect 624 22266 656 22298
rect 696 22266 728 22298
rect 768 22266 800 22298
rect 840 22266 872 22298
rect 912 22266 944 22298
rect 984 22266 1016 22298
rect 1056 22266 1088 22298
rect 1128 22266 1160 22298
rect 1200 22266 1232 22298
rect 1272 22266 1304 22298
rect 1344 22266 1376 22298
rect 1416 22266 1448 22298
rect 1488 22266 1520 22298
rect 1560 22266 1592 22298
rect 1632 22266 1664 22298
rect 1704 22266 1736 22298
rect 1776 22266 1808 22298
rect 1848 22266 1880 22298
rect 120 22194 152 22226
rect 192 22194 224 22226
rect 264 22194 296 22226
rect 336 22194 368 22226
rect 408 22194 440 22226
rect 480 22194 512 22226
rect 552 22194 584 22226
rect 624 22194 656 22226
rect 696 22194 728 22226
rect 768 22194 800 22226
rect 840 22194 872 22226
rect 912 22194 944 22226
rect 984 22194 1016 22226
rect 1056 22194 1088 22226
rect 1128 22194 1160 22226
rect 1200 22194 1232 22226
rect 1272 22194 1304 22226
rect 1344 22194 1376 22226
rect 1416 22194 1448 22226
rect 1488 22194 1520 22226
rect 1560 22194 1592 22226
rect 1632 22194 1664 22226
rect 1704 22194 1736 22226
rect 1776 22194 1808 22226
rect 1848 22194 1880 22226
rect 120 22122 152 22154
rect 192 22122 224 22154
rect 264 22122 296 22154
rect 336 22122 368 22154
rect 408 22122 440 22154
rect 480 22122 512 22154
rect 552 22122 584 22154
rect 624 22122 656 22154
rect 696 22122 728 22154
rect 768 22122 800 22154
rect 840 22122 872 22154
rect 912 22122 944 22154
rect 984 22122 1016 22154
rect 1056 22122 1088 22154
rect 1128 22122 1160 22154
rect 1200 22122 1232 22154
rect 1272 22122 1304 22154
rect 1344 22122 1376 22154
rect 1416 22122 1448 22154
rect 1488 22122 1520 22154
rect 1560 22122 1592 22154
rect 1632 22122 1664 22154
rect 1704 22122 1736 22154
rect 1776 22122 1808 22154
rect 1848 22122 1880 22154
rect 120 22050 152 22082
rect 192 22050 224 22082
rect 264 22050 296 22082
rect 336 22050 368 22082
rect 408 22050 440 22082
rect 480 22050 512 22082
rect 552 22050 584 22082
rect 624 22050 656 22082
rect 696 22050 728 22082
rect 768 22050 800 22082
rect 840 22050 872 22082
rect 912 22050 944 22082
rect 984 22050 1016 22082
rect 1056 22050 1088 22082
rect 1128 22050 1160 22082
rect 1200 22050 1232 22082
rect 1272 22050 1304 22082
rect 1344 22050 1376 22082
rect 1416 22050 1448 22082
rect 1488 22050 1520 22082
rect 1560 22050 1592 22082
rect 1632 22050 1664 22082
rect 1704 22050 1736 22082
rect 1776 22050 1808 22082
rect 1848 22050 1880 22082
rect 120 21978 152 22010
rect 192 21978 224 22010
rect 264 21978 296 22010
rect 336 21978 368 22010
rect 408 21978 440 22010
rect 480 21978 512 22010
rect 552 21978 584 22010
rect 624 21978 656 22010
rect 696 21978 728 22010
rect 768 21978 800 22010
rect 840 21978 872 22010
rect 912 21978 944 22010
rect 984 21978 1016 22010
rect 1056 21978 1088 22010
rect 1128 21978 1160 22010
rect 1200 21978 1232 22010
rect 1272 21978 1304 22010
rect 1344 21978 1376 22010
rect 1416 21978 1448 22010
rect 1488 21978 1520 22010
rect 1560 21978 1592 22010
rect 1632 21978 1664 22010
rect 1704 21978 1736 22010
rect 1776 21978 1808 22010
rect 1848 21978 1880 22010
rect 120 21906 152 21938
rect 192 21906 224 21938
rect 264 21906 296 21938
rect 336 21906 368 21938
rect 408 21906 440 21938
rect 480 21906 512 21938
rect 552 21906 584 21938
rect 624 21906 656 21938
rect 696 21906 728 21938
rect 768 21906 800 21938
rect 840 21906 872 21938
rect 912 21906 944 21938
rect 984 21906 1016 21938
rect 1056 21906 1088 21938
rect 1128 21906 1160 21938
rect 1200 21906 1232 21938
rect 1272 21906 1304 21938
rect 1344 21906 1376 21938
rect 1416 21906 1448 21938
rect 1488 21906 1520 21938
rect 1560 21906 1592 21938
rect 1632 21906 1664 21938
rect 1704 21906 1736 21938
rect 1776 21906 1808 21938
rect 1848 21906 1880 21938
rect 120 21834 152 21866
rect 192 21834 224 21866
rect 264 21834 296 21866
rect 336 21834 368 21866
rect 408 21834 440 21866
rect 480 21834 512 21866
rect 552 21834 584 21866
rect 624 21834 656 21866
rect 696 21834 728 21866
rect 768 21834 800 21866
rect 840 21834 872 21866
rect 912 21834 944 21866
rect 984 21834 1016 21866
rect 1056 21834 1088 21866
rect 1128 21834 1160 21866
rect 1200 21834 1232 21866
rect 1272 21834 1304 21866
rect 1344 21834 1376 21866
rect 1416 21834 1448 21866
rect 1488 21834 1520 21866
rect 1560 21834 1592 21866
rect 1632 21834 1664 21866
rect 1704 21834 1736 21866
rect 1776 21834 1808 21866
rect 1848 21834 1880 21866
rect 120 21762 152 21794
rect 192 21762 224 21794
rect 264 21762 296 21794
rect 336 21762 368 21794
rect 408 21762 440 21794
rect 480 21762 512 21794
rect 552 21762 584 21794
rect 624 21762 656 21794
rect 696 21762 728 21794
rect 768 21762 800 21794
rect 840 21762 872 21794
rect 912 21762 944 21794
rect 984 21762 1016 21794
rect 1056 21762 1088 21794
rect 1128 21762 1160 21794
rect 1200 21762 1232 21794
rect 1272 21762 1304 21794
rect 1344 21762 1376 21794
rect 1416 21762 1448 21794
rect 1488 21762 1520 21794
rect 1560 21762 1592 21794
rect 1632 21762 1664 21794
rect 1704 21762 1736 21794
rect 1776 21762 1808 21794
rect 1848 21762 1880 21794
rect 120 21690 152 21722
rect 192 21690 224 21722
rect 264 21690 296 21722
rect 336 21690 368 21722
rect 408 21690 440 21722
rect 480 21690 512 21722
rect 552 21690 584 21722
rect 624 21690 656 21722
rect 696 21690 728 21722
rect 768 21690 800 21722
rect 840 21690 872 21722
rect 912 21690 944 21722
rect 984 21690 1016 21722
rect 1056 21690 1088 21722
rect 1128 21690 1160 21722
rect 1200 21690 1232 21722
rect 1272 21690 1304 21722
rect 1344 21690 1376 21722
rect 1416 21690 1448 21722
rect 1488 21690 1520 21722
rect 1560 21690 1592 21722
rect 1632 21690 1664 21722
rect 1704 21690 1736 21722
rect 1776 21690 1808 21722
rect 1848 21690 1880 21722
rect 120 21618 152 21650
rect 192 21618 224 21650
rect 264 21618 296 21650
rect 336 21618 368 21650
rect 408 21618 440 21650
rect 480 21618 512 21650
rect 552 21618 584 21650
rect 624 21618 656 21650
rect 696 21618 728 21650
rect 768 21618 800 21650
rect 840 21618 872 21650
rect 912 21618 944 21650
rect 984 21618 1016 21650
rect 1056 21618 1088 21650
rect 1128 21618 1160 21650
rect 1200 21618 1232 21650
rect 1272 21618 1304 21650
rect 1344 21618 1376 21650
rect 1416 21618 1448 21650
rect 1488 21618 1520 21650
rect 1560 21618 1592 21650
rect 1632 21618 1664 21650
rect 1704 21618 1736 21650
rect 1776 21618 1808 21650
rect 1848 21618 1880 21650
rect 120 21546 152 21578
rect 192 21546 224 21578
rect 264 21546 296 21578
rect 336 21546 368 21578
rect 408 21546 440 21578
rect 480 21546 512 21578
rect 552 21546 584 21578
rect 624 21546 656 21578
rect 696 21546 728 21578
rect 768 21546 800 21578
rect 840 21546 872 21578
rect 912 21546 944 21578
rect 984 21546 1016 21578
rect 1056 21546 1088 21578
rect 1128 21546 1160 21578
rect 1200 21546 1232 21578
rect 1272 21546 1304 21578
rect 1344 21546 1376 21578
rect 1416 21546 1448 21578
rect 1488 21546 1520 21578
rect 1560 21546 1592 21578
rect 1632 21546 1664 21578
rect 1704 21546 1736 21578
rect 1776 21546 1808 21578
rect 1848 21546 1880 21578
rect 120 21474 152 21506
rect 192 21474 224 21506
rect 264 21474 296 21506
rect 336 21474 368 21506
rect 408 21474 440 21506
rect 480 21474 512 21506
rect 552 21474 584 21506
rect 624 21474 656 21506
rect 696 21474 728 21506
rect 768 21474 800 21506
rect 840 21474 872 21506
rect 912 21474 944 21506
rect 984 21474 1016 21506
rect 1056 21474 1088 21506
rect 1128 21474 1160 21506
rect 1200 21474 1232 21506
rect 1272 21474 1304 21506
rect 1344 21474 1376 21506
rect 1416 21474 1448 21506
rect 1488 21474 1520 21506
rect 1560 21474 1592 21506
rect 1632 21474 1664 21506
rect 1704 21474 1736 21506
rect 1776 21474 1808 21506
rect 1848 21474 1880 21506
rect 120 21402 152 21434
rect 192 21402 224 21434
rect 264 21402 296 21434
rect 336 21402 368 21434
rect 408 21402 440 21434
rect 480 21402 512 21434
rect 552 21402 584 21434
rect 624 21402 656 21434
rect 696 21402 728 21434
rect 768 21402 800 21434
rect 840 21402 872 21434
rect 912 21402 944 21434
rect 984 21402 1016 21434
rect 1056 21402 1088 21434
rect 1128 21402 1160 21434
rect 1200 21402 1232 21434
rect 1272 21402 1304 21434
rect 1344 21402 1376 21434
rect 1416 21402 1448 21434
rect 1488 21402 1520 21434
rect 1560 21402 1592 21434
rect 1632 21402 1664 21434
rect 1704 21402 1736 21434
rect 1776 21402 1808 21434
rect 1848 21402 1880 21434
rect 120 21330 152 21362
rect 192 21330 224 21362
rect 264 21330 296 21362
rect 336 21330 368 21362
rect 408 21330 440 21362
rect 480 21330 512 21362
rect 552 21330 584 21362
rect 624 21330 656 21362
rect 696 21330 728 21362
rect 768 21330 800 21362
rect 840 21330 872 21362
rect 912 21330 944 21362
rect 984 21330 1016 21362
rect 1056 21330 1088 21362
rect 1128 21330 1160 21362
rect 1200 21330 1232 21362
rect 1272 21330 1304 21362
rect 1344 21330 1376 21362
rect 1416 21330 1448 21362
rect 1488 21330 1520 21362
rect 1560 21330 1592 21362
rect 1632 21330 1664 21362
rect 1704 21330 1736 21362
rect 1776 21330 1808 21362
rect 1848 21330 1880 21362
rect 120 21258 152 21290
rect 192 21258 224 21290
rect 264 21258 296 21290
rect 336 21258 368 21290
rect 408 21258 440 21290
rect 480 21258 512 21290
rect 552 21258 584 21290
rect 624 21258 656 21290
rect 696 21258 728 21290
rect 768 21258 800 21290
rect 840 21258 872 21290
rect 912 21258 944 21290
rect 984 21258 1016 21290
rect 1056 21258 1088 21290
rect 1128 21258 1160 21290
rect 1200 21258 1232 21290
rect 1272 21258 1304 21290
rect 1344 21258 1376 21290
rect 1416 21258 1448 21290
rect 1488 21258 1520 21290
rect 1560 21258 1592 21290
rect 1632 21258 1664 21290
rect 1704 21258 1736 21290
rect 1776 21258 1808 21290
rect 1848 21258 1880 21290
rect 120 21186 152 21218
rect 192 21186 224 21218
rect 264 21186 296 21218
rect 336 21186 368 21218
rect 408 21186 440 21218
rect 480 21186 512 21218
rect 552 21186 584 21218
rect 624 21186 656 21218
rect 696 21186 728 21218
rect 768 21186 800 21218
rect 840 21186 872 21218
rect 912 21186 944 21218
rect 984 21186 1016 21218
rect 1056 21186 1088 21218
rect 1128 21186 1160 21218
rect 1200 21186 1232 21218
rect 1272 21186 1304 21218
rect 1344 21186 1376 21218
rect 1416 21186 1448 21218
rect 1488 21186 1520 21218
rect 1560 21186 1592 21218
rect 1632 21186 1664 21218
rect 1704 21186 1736 21218
rect 1776 21186 1808 21218
rect 1848 21186 1880 21218
rect 120 21114 152 21146
rect 192 21114 224 21146
rect 264 21114 296 21146
rect 336 21114 368 21146
rect 408 21114 440 21146
rect 480 21114 512 21146
rect 552 21114 584 21146
rect 624 21114 656 21146
rect 696 21114 728 21146
rect 768 21114 800 21146
rect 840 21114 872 21146
rect 912 21114 944 21146
rect 984 21114 1016 21146
rect 1056 21114 1088 21146
rect 1128 21114 1160 21146
rect 1200 21114 1232 21146
rect 1272 21114 1304 21146
rect 1344 21114 1376 21146
rect 1416 21114 1448 21146
rect 1488 21114 1520 21146
rect 1560 21114 1592 21146
rect 1632 21114 1664 21146
rect 1704 21114 1736 21146
rect 1776 21114 1808 21146
rect 1848 21114 1880 21146
rect 120 21042 152 21074
rect 192 21042 224 21074
rect 264 21042 296 21074
rect 336 21042 368 21074
rect 408 21042 440 21074
rect 480 21042 512 21074
rect 552 21042 584 21074
rect 624 21042 656 21074
rect 696 21042 728 21074
rect 768 21042 800 21074
rect 840 21042 872 21074
rect 912 21042 944 21074
rect 984 21042 1016 21074
rect 1056 21042 1088 21074
rect 1128 21042 1160 21074
rect 1200 21042 1232 21074
rect 1272 21042 1304 21074
rect 1344 21042 1376 21074
rect 1416 21042 1448 21074
rect 1488 21042 1520 21074
rect 1560 21042 1592 21074
rect 1632 21042 1664 21074
rect 1704 21042 1736 21074
rect 1776 21042 1808 21074
rect 1848 21042 1880 21074
rect 120 20970 152 21002
rect 192 20970 224 21002
rect 264 20970 296 21002
rect 336 20970 368 21002
rect 408 20970 440 21002
rect 480 20970 512 21002
rect 552 20970 584 21002
rect 624 20970 656 21002
rect 696 20970 728 21002
rect 768 20970 800 21002
rect 840 20970 872 21002
rect 912 20970 944 21002
rect 984 20970 1016 21002
rect 1056 20970 1088 21002
rect 1128 20970 1160 21002
rect 1200 20970 1232 21002
rect 1272 20970 1304 21002
rect 1344 20970 1376 21002
rect 1416 20970 1448 21002
rect 1488 20970 1520 21002
rect 1560 20970 1592 21002
rect 1632 20970 1664 21002
rect 1704 20970 1736 21002
rect 1776 20970 1808 21002
rect 1848 20970 1880 21002
rect 120 20898 152 20930
rect 192 20898 224 20930
rect 264 20898 296 20930
rect 336 20898 368 20930
rect 408 20898 440 20930
rect 480 20898 512 20930
rect 552 20898 584 20930
rect 624 20898 656 20930
rect 696 20898 728 20930
rect 768 20898 800 20930
rect 840 20898 872 20930
rect 912 20898 944 20930
rect 984 20898 1016 20930
rect 1056 20898 1088 20930
rect 1128 20898 1160 20930
rect 1200 20898 1232 20930
rect 1272 20898 1304 20930
rect 1344 20898 1376 20930
rect 1416 20898 1448 20930
rect 1488 20898 1520 20930
rect 1560 20898 1592 20930
rect 1632 20898 1664 20930
rect 1704 20898 1736 20930
rect 1776 20898 1808 20930
rect 1848 20898 1880 20930
rect 120 20826 152 20858
rect 192 20826 224 20858
rect 264 20826 296 20858
rect 336 20826 368 20858
rect 408 20826 440 20858
rect 480 20826 512 20858
rect 552 20826 584 20858
rect 624 20826 656 20858
rect 696 20826 728 20858
rect 768 20826 800 20858
rect 840 20826 872 20858
rect 912 20826 944 20858
rect 984 20826 1016 20858
rect 1056 20826 1088 20858
rect 1128 20826 1160 20858
rect 1200 20826 1232 20858
rect 1272 20826 1304 20858
rect 1344 20826 1376 20858
rect 1416 20826 1448 20858
rect 1488 20826 1520 20858
rect 1560 20826 1592 20858
rect 1632 20826 1664 20858
rect 1704 20826 1736 20858
rect 1776 20826 1808 20858
rect 1848 20826 1880 20858
rect 120 20754 152 20786
rect 192 20754 224 20786
rect 264 20754 296 20786
rect 336 20754 368 20786
rect 408 20754 440 20786
rect 480 20754 512 20786
rect 552 20754 584 20786
rect 624 20754 656 20786
rect 696 20754 728 20786
rect 768 20754 800 20786
rect 840 20754 872 20786
rect 912 20754 944 20786
rect 984 20754 1016 20786
rect 1056 20754 1088 20786
rect 1128 20754 1160 20786
rect 1200 20754 1232 20786
rect 1272 20754 1304 20786
rect 1344 20754 1376 20786
rect 1416 20754 1448 20786
rect 1488 20754 1520 20786
rect 1560 20754 1592 20786
rect 1632 20754 1664 20786
rect 1704 20754 1736 20786
rect 1776 20754 1808 20786
rect 1848 20754 1880 20786
rect 120 20682 152 20714
rect 192 20682 224 20714
rect 264 20682 296 20714
rect 336 20682 368 20714
rect 408 20682 440 20714
rect 480 20682 512 20714
rect 552 20682 584 20714
rect 624 20682 656 20714
rect 696 20682 728 20714
rect 768 20682 800 20714
rect 840 20682 872 20714
rect 912 20682 944 20714
rect 984 20682 1016 20714
rect 1056 20682 1088 20714
rect 1128 20682 1160 20714
rect 1200 20682 1232 20714
rect 1272 20682 1304 20714
rect 1344 20682 1376 20714
rect 1416 20682 1448 20714
rect 1488 20682 1520 20714
rect 1560 20682 1592 20714
rect 1632 20682 1664 20714
rect 1704 20682 1736 20714
rect 1776 20682 1808 20714
rect 1848 20682 1880 20714
rect 120 20610 152 20642
rect 192 20610 224 20642
rect 264 20610 296 20642
rect 336 20610 368 20642
rect 408 20610 440 20642
rect 480 20610 512 20642
rect 552 20610 584 20642
rect 624 20610 656 20642
rect 696 20610 728 20642
rect 768 20610 800 20642
rect 840 20610 872 20642
rect 912 20610 944 20642
rect 984 20610 1016 20642
rect 1056 20610 1088 20642
rect 1128 20610 1160 20642
rect 1200 20610 1232 20642
rect 1272 20610 1304 20642
rect 1344 20610 1376 20642
rect 1416 20610 1448 20642
rect 1488 20610 1520 20642
rect 1560 20610 1592 20642
rect 1632 20610 1664 20642
rect 1704 20610 1736 20642
rect 1776 20610 1808 20642
rect 1848 20610 1880 20642
rect 120 20538 152 20570
rect 192 20538 224 20570
rect 264 20538 296 20570
rect 336 20538 368 20570
rect 408 20538 440 20570
rect 480 20538 512 20570
rect 552 20538 584 20570
rect 624 20538 656 20570
rect 696 20538 728 20570
rect 768 20538 800 20570
rect 840 20538 872 20570
rect 912 20538 944 20570
rect 984 20538 1016 20570
rect 1056 20538 1088 20570
rect 1128 20538 1160 20570
rect 1200 20538 1232 20570
rect 1272 20538 1304 20570
rect 1344 20538 1376 20570
rect 1416 20538 1448 20570
rect 1488 20538 1520 20570
rect 1560 20538 1592 20570
rect 1632 20538 1664 20570
rect 1704 20538 1736 20570
rect 1776 20538 1808 20570
rect 1848 20538 1880 20570
rect 120 20466 152 20498
rect 192 20466 224 20498
rect 264 20466 296 20498
rect 336 20466 368 20498
rect 408 20466 440 20498
rect 480 20466 512 20498
rect 552 20466 584 20498
rect 624 20466 656 20498
rect 696 20466 728 20498
rect 768 20466 800 20498
rect 840 20466 872 20498
rect 912 20466 944 20498
rect 984 20466 1016 20498
rect 1056 20466 1088 20498
rect 1128 20466 1160 20498
rect 1200 20466 1232 20498
rect 1272 20466 1304 20498
rect 1344 20466 1376 20498
rect 1416 20466 1448 20498
rect 1488 20466 1520 20498
rect 1560 20466 1592 20498
rect 1632 20466 1664 20498
rect 1704 20466 1736 20498
rect 1776 20466 1808 20498
rect 1848 20466 1880 20498
rect 120 20394 152 20426
rect 192 20394 224 20426
rect 264 20394 296 20426
rect 336 20394 368 20426
rect 408 20394 440 20426
rect 480 20394 512 20426
rect 552 20394 584 20426
rect 624 20394 656 20426
rect 696 20394 728 20426
rect 768 20394 800 20426
rect 840 20394 872 20426
rect 912 20394 944 20426
rect 984 20394 1016 20426
rect 1056 20394 1088 20426
rect 1128 20394 1160 20426
rect 1200 20394 1232 20426
rect 1272 20394 1304 20426
rect 1344 20394 1376 20426
rect 1416 20394 1448 20426
rect 1488 20394 1520 20426
rect 1560 20394 1592 20426
rect 1632 20394 1664 20426
rect 1704 20394 1736 20426
rect 1776 20394 1808 20426
rect 1848 20394 1880 20426
rect 120 20322 152 20354
rect 192 20322 224 20354
rect 264 20322 296 20354
rect 336 20322 368 20354
rect 408 20322 440 20354
rect 480 20322 512 20354
rect 552 20322 584 20354
rect 624 20322 656 20354
rect 696 20322 728 20354
rect 768 20322 800 20354
rect 840 20322 872 20354
rect 912 20322 944 20354
rect 984 20322 1016 20354
rect 1056 20322 1088 20354
rect 1128 20322 1160 20354
rect 1200 20322 1232 20354
rect 1272 20322 1304 20354
rect 1344 20322 1376 20354
rect 1416 20322 1448 20354
rect 1488 20322 1520 20354
rect 1560 20322 1592 20354
rect 1632 20322 1664 20354
rect 1704 20322 1736 20354
rect 1776 20322 1808 20354
rect 1848 20322 1880 20354
rect 120 20250 152 20282
rect 192 20250 224 20282
rect 264 20250 296 20282
rect 336 20250 368 20282
rect 408 20250 440 20282
rect 480 20250 512 20282
rect 552 20250 584 20282
rect 624 20250 656 20282
rect 696 20250 728 20282
rect 768 20250 800 20282
rect 840 20250 872 20282
rect 912 20250 944 20282
rect 984 20250 1016 20282
rect 1056 20250 1088 20282
rect 1128 20250 1160 20282
rect 1200 20250 1232 20282
rect 1272 20250 1304 20282
rect 1344 20250 1376 20282
rect 1416 20250 1448 20282
rect 1488 20250 1520 20282
rect 1560 20250 1592 20282
rect 1632 20250 1664 20282
rect 1704 20250 1736 20282
rect 1776 20250 1808 20282
rect 1848 20250 1880 20282
rect 120 20178 152 20210
rect 192 20178 224 20210
rect 264 20178 296 20210
rect 336 20178 368 20210
rect 408 20178 440 20210
rect 480 20178 512 20210
rect 552 20178 584 20210
rect 624 20178 656 20210
rect 696 20178 728 20210
rect 768 20178 800 20210
rect 840 20178 872 20210
rect 912 20178 944 20210
rect 984 20178 1016 20210
rect 1056 20178 1088 20210
rect 1128 20178 1160 20210
rect 1200 20178 1232 20210
rect 1272 20178 1304 20210
rect 1344 20178 1376 20210
rect 1416 20178 1448 20210
rect 1488 20178 1520 20210
rect 1560 20178 1592 20210
rect 1632 20178 1664 20210
rect 1704 20178 1736 20210
rect 1776 20178 1808 20210
rect 1848 20178 1880 20210
rect 120 20106 152 20138
rect 192 20106 224 20138
rect 264 20106 296 20138
rect 336 20106 368 20138
rect 408 20106 440 20138
rect 480 20106 512 20138
rect 552 20106 584 20138
rect 624 20106 656 20138
rect 696 20106 728 20138
rect 768 20106 800 20138
rect 840 20106 872 20138
rect 912 20106 944 20138
rect 984 20106 1016 20138
rect 1056 20106 1088 20138
rect 1128 20106 1160 20138
rect 1200 20106 1232 20138
rect 1272 20106 1304 20138
rect 1344 20106 1376 20138
rect 1416 20106 1448 20138
rect 1488 20106 1520 20138
rect 1560 20106 1592 20138
rect 1632 20106 1664 20138
rect 1704 20106 1736 20138
rect 1776 20106 1808 20138
rect 1848 20106 1880 20138
rect 120 20034 152 20066
rect 192 20034 224 20066
rect 264 20034 296 20066
rect 336 20034 368 20066
rect 408 20034 440 20066
rect 480 20034 512 20066
rect 552 20034 584 20066
rect 624 20034 656 20066
rect 696 20034 728 20066
rect 768 20034 800 20066
rect 840 20034 872 20066
rect 912 20034 944 20066
rect 984 20034 1016 20066
rect 1056 20034 1088 20066
rect 1128 20034 1160 20066
rect 1200 20034 1232 20066
rect 1272 20034 1304 20066
rect 1344 20034 1376 20066
rect 1416 20034 1448 20066
rect 1488 20034 1520 20066
rect 1560 20034 1592 20066
rect 1632 20034 1664 20066
rect 1704 20034 1736 20066
rect 1776 20034 1808 20066
rect 1848 20034 1880 20066
rect 120 19962 152 19994
rect 192 19962 224 19994
rect 264 19962 296 19994
rect 336 19962 368 19994
rect 408 19962 440 19994
rect 480 19962 512 19994
rect 552 19962 584 19994
rect 624 19962 656 19994
rect 696 19962 728 19994
rect 768 19962 800 19994
rect 840 19962 872 19994
rect 912 19962 944 19994
rect 984 19962 1016 19994
rect 1056 19962 1088 19994
rect 1128 19962 1160 19994
rect 1200 19962 1232 19994
rect 1272 19962 1304 19994
rect 1344 19962 1376 19994
rect 1416 19962 1448 19994
rect 1488 19962 1520 19994
rect 1560 19962 1592 19994
rect 1632 19962 1664 19994
rect 1704 19962 1736 19994
rect 1776 19962 1808 19994
rect 1848 19962 1880 19994
rect 120 19890 152 19922
rect 192 19890 224 19922
rect 264 19890 296 19922
rect 336 19890 368 19922
rect 408 19890 440 19922
rect 480 19890 512 19922
rect 552 19890 584 19922
rect 624 19890 656 19922
rect 696 19890 728 19922
rect 768 19890 800 19922
rect 840 19890 872 19922
rect 912 19890 944 19922
rect 984 19890 1016 19922
rect 1056 19890 1088 19922
rect 1128 19890 1160 19922
rect 1200 19890 1232 19922
rect 1272 19890 1304 19922
rect 1344 19890 1376 19922
rect 1416 19890 1448 19922
rect 1488 19890 1520 19922
rect 1560 19890 1592 19922
rect 1632 19890 1664 19922
rect 1704 19890 1736 19922
rect 1776 19890 1808 19922
rect 1848 19890 1880 19922
rect 120 19818 152 19850
rect 192 19818 224 19850
rect 264 19818 296 19850
rect 336 19818 368 19850
rect 408 19818 440 19850
rect 480 19818 512 19850
rect 552 19818 584 19850
rect 624 19818 656 19850
rect 696 19818 728 19850
rect 768 19818 800 19850
rect 840 19818 872 19850
rect 912 19818 944 19850
rect 984 19818 1016 19850
rect 1056 19818 1088 19850
rect 1128 19818 1160 19850
rect 1200 19818 1232 19850
rect 1272 19818 1304 19850
rect 1344 19818 1376 19850
rect 1416 19818 1448 19850
rect 1488 19818 1520 19850
rect 1560 19818 1592 19850
rect 1632 19818 1664 19850
rect 1704 19818 1736 19850
rect 1776 19818 1808 19850
rect 1848 19818 1880 19850
rect 120 19746 152 19778
rect 192 19746 224 19778
rect 264 19746 296 19778
rect 336 19746 368 19778
rect 408 19746 440 19778
rect 480 19746 512 19778
rect 552 19746 584 19778
rect 624 19746 656 19778
rect 696 19746 728 19778
rect 768 19746 800 19778
rect 840 19746 872 19778
rect 912 19746 944 19778
rect 984 19746 1016 19778
rect 1056 19746 1088 19778
rect 1128 19746 1160 19778
rect 1200 19746 1232 19778
rect 1272 19746 1304 19778
rect 1344 19746 1376 19778
rect 1416 19746 1448 19778
rect 1488 19746 1520 19778
rect 1560 19746 1592 19778
rect 1632 19746 1664 19778
rect 1704 19746 1736 19778
rect 1776 19746 1808 19778
rect 1848 19746 1880 19778
rect 120 19674 152 19706
rect 192 19674 224 19706
rect 264 19674 296 19706
rect 336 19674 368 19706
rect 408 19674 440 19706
rect 480 19674 512 19706
rect 552 19674 584 19706
rect 624 19674 656 19706
rect 696 19674 728 19706
rect 768 19674 800 19706
rect 840 19674 872 19706
rect 912 19674 944 19706
rect 984 19674 1016 19706
rect 1056 19674 1088 19706
rect 1128 19674 1160 19706
rect 1200 19674 1232 19706
rect 1272 19674 1304 19706
rect 1344 19674 1376 19706
rect 1416 19674 1448 19706
rect 1488 19674 1520 19706
rect 1560 19674 1592 19706
rect 1632 19674 1664 19706
rect 1704 19674 1736 19706
rect 1776 19674 1808 19706
rect 1848 19674 1880 19706
rect 120 19602 152 19634
rect 192 19602 224 19634
rect 264 19602 296 19634
rect 336 19602 368 19634
rect 408 19602 440 19634
rect 480 19602 512 19634
rect 552 19602 584 19634
rect 624 19602 656 19634
rect 696 19602 728 19634
rect 768 19602 800 19634
rect 840 19602 872 19634
rect 912 19602 944 19634
rect 984 19602 1016 19634
rect 1056 19602 1088 19634
rect 1128 19602 1160 19634
rect 1200 19602 1232 19634
rect 1272 19602 1304 19634
rect 1344 19602 1376 19634
rect 1416 19602 1448 19634
rect 1488 19602 1520 19634
rect 1560 19602 1592 19634
rect 1632 19602 1664 19634
rect 1704 19602 1736 19634
rect 1776 19602 1808 19634
rect 1848 19602 1880 19634
rect 120 19530 152 19562
rect 192 19530 224 19562
rect 264 19530 296 19562
rect 336 19530 368 19562
rect 408 19530 440 19562
rect 480 19530 512 19562
rect 552 19530 584 19562
rect 624 19530 656 19562
rect 696 19530 728 19562
rect 768 19530 800 19562
rect 840 19530 872 19562
rect 912 19530 944 19562
rect 984 19530 1016 19562
rect 1056 19530 1088 19562
rect 1128 19530 1160 19562
rect 1200 19530 1232 19562
rect 1272 19530 1304 19562
rect 1344 19530 1376 19562
rect 1416 19530 1448 19562
rect 1488 19530 1520 19562
rect 1560 19530 1592 19562
rect 1632 19530 1664 19562
rect 1704 19530 1736 19562
rect 1776 19530 1808 19562
rect 1848 19530 1880 19562
rect 120 19458 152 19490
rect 192 19458 224 19490
rect 264 19458 296 19490
rect 336 19458 368 19490
rect 408 19458 440 19490
rect 480 19458 512 19490
rect 552 19458 584 19490
rect 624 19458 656 19490
rect 696 19458 728 19490
rect 768 19458 800 19490
rect 840 19458 872 19490
rect 912 19458 944 19490
rect 984 19458 1016 19490
rect 1056 19458 1088 19490
rect 1128 19458 1160 19490
rect 1200 19458 1232 19490
rect 1272 19458 1304 19490
rect 1344 19458 1376 19490
rect 1416 19458 1448 19490
rect 1488 19458 1520 19490
rect 1560 19458 1592 19490
rect 1632 19458 1664 19490
rect 1704 19458 1736 19490
rect 1776 19458 1808 19490
rect 1848 19458 1880 19490
rect 120 19386 152 19418
rect 192 19386 224 19418
rect 264 19386 296 19418
rect 336 19386 368 19418
rect 408 19386 440 19418
rect 480 19386 512 19418
rect 552 19386 584 19418
rect 624 19386 656 19418
rect 696 19386 728 19418
rect 768 19386 800 19418
rect 840 19386 872 19418
rect 912 19386 944 19418
rect 984 19386 1016 19418
rect 1056 19386 1088 19418
rect 1128 19386 1160 19418
rect 1200 19386 1232 19418
rect 1272 19386 1304 19418
rect 1344 19386 1376 19418
rect 1416 19386 1448 19418
rect 1488 19386 1520 19418
rect 1560 19386 1592 19418
rect 1632 19386 1664 19418
rect 1704 19386 1736 19418
rect 1776 19386 1808 19418
rect 1848 19386 1880 19418
rect 120 19314 152 19346
rect 192 19314 224 19346
rect 264 19314 296 19346
rect 336 19314 368 19346
rect 408 19314 440 19346
rect 480 19314 512 19346
rect 552 19314 584 19346
rect 624 19314 656 19346
rect 696 19314 728 19346
rect 768 19314 800 19346
rect 840 19314 872 19346
rect 912 19314 944 19346
rect 984 19314 1016 19346
rect 1056 19314 1088 19346
rect 1128 19314 1160 19346
rect 1200 19314 1232 19346
rect 1272 19314 1304 19346
rect 1344 19314 1376 19346
rect 1416 19314 1448 19346
rect 1488 19314 1520 19346
rect 1560 19314 1592 19346
rect 1632 19314 1664 19346
rect 1704 19314 1736 19346
rect 1776 19314 1808 19346
rect 1848 19314 1880 19346
rect 120 19242 152 19274
rect 192 19242 224 19274
rect 264 19242 296 19274
rect 336 19242 368 19274
rect 408 19242 440 19274
rect 480 19242 512 19274
rect 552 19242 584 19274
rect 624 19242 656 19274
rect 696 19242 728 19274
rect 768 19242 800 19274
rect 840 19242 872 19274
rect 912 19242 944 19274
rect 984 19242 1016 19274
rect 1056 19242 1088 19274
rect 1128 19242 1160 19274
rect 1200 19242 1232 19274
rect 1272 19242 1304 19274
rect 1344 19242 1376 19274
rect 1416 19242 1448 19274
rect 1488 19242 1520 19274
rect 1560 19242 1592 19274
rect 1632 19242 1664 19274
rect 1704 19242 1736 19274
rect 1776 19242 1808 19274
rect 1848 19242 1880 19274
rect 120 19170 152 19202
rect 192 19170 224 19202
rect 264 19170 296 19202
rect 336 19170 368 19202
rect 408 19170 440 19202
rect 480 19170 512 19202
rect 552 19170 584 19202
rect 624 19170 656 19202
rect 696 19170 728 19202
rect 768 19170 800 19202
rect 840 19170 872 19202
rect 912 19170 944 19202
rect 984 19170 1016 19202
rect 1056 19170 1088 19202
rect 1128 19170 1160 19202
rect 1200 19170 1232 19202
rect 1272 19170 1304 19202
rect 1344 19170 1376 19202
rect 1416 19170 1448 19202
rect 1488 19170 1520 19202
rect 1560 19170 1592 19202
rect 1632 19170 1664 19202
rect 1704 19170 1736 19202
rect 1776 19170 1808 19202
rect 1848 19170 1880 19202
rect 120 19098 152 19130
rect 192 19098 224 19130
rect 264 19098 296 19130
rect 336 19098 368 19130
rect 408 19098 440 19130
rect 480 19098 512 19130
rect 552 19098 584 19130
rect 624 19098 656 19130
rect 696 19098 728 19130
rect 768 19098 800 19130
rect 840 19098 872 19130
rect 912 19098 944 19130
rect 984 19098 1016 19130
rect 1056 19098 1088 19130
rect 1128 19098 1160 19130
rect 1200 19098 1232 19130
rect 1272 19098 1304 19130
rect 1344 19098 1376 19130
rect 1416 19098 1448 19130
rect 1488 19098 1520 19130
rect 1560 19098 1592 19130
rect 1632 19098 1664 19130
rect 1704 19098 1736 19130
rect 1776 19098 1808 19130
rect 1848 19098 1880 19130
rect 120 19026 152 19058
rect 192 19026 224 19058
rect 264 19026 296 19058
rect 336 19026 368 19058
rect 408 19026 440 19058
rect 480 19026 512 19058
rect 552 19026 584 19058
rect 624 19026 656 19058
rect 696 19026 728 19058
rect 768 19026 800 19058
rect 840 19026 872 19058
rect 912 19026 944 19058
rect 984 19026 1016 19058
rect 1056 19026 1088 19058
rect 1128 19026 1160 19058
rect 1200 19026 1232 19058
rect 1272 19026 1304 19058
rect 1344 19026 1376 19058
rect 1416 19026 1448 19058
rect 1488 19026 1520 19058
rect 1560 19026 1592 19058
rect 1632 19026 1664 19058
rect 1704 19026 1736 19058
rect 1776 19026 1808 19058
rect 1848 19026 1880 19058
rect 120 18954 152 18986
rect 192 18954 224 18986
rect 264 18954 296 18986
rect 336 18954 368 18986
rect 408 18954 440 18986
rect 480 18954 512 18986
rect 552 18954 584 18986
rect 624 18954 656 18986
rect 696 18954 728 18986
rect 768 18954 800 18986
rect 840 18954 872 18986
rect 912 18954 944 18986
rect 984 18954 1016 18986
rect 1056 18954 1088 18986
rect 1128 18954 1160 18986
rect 1200 18954 1232 18986
rect 1272 18954 1304 18986
rect 1344 18954 1376 18986
rect 1416 18954 1448 18986
rect 1488 18954 1520 18986
rect 1560 18954 1592 18986
rect 1632 18954 1664 18986
rect 1704 18954 1736 18986
rect 1776 18954 1808 18986
rect 1848 18954 1880 18986
rect 120 18882 152 18914
rect 192 18882 224 18914
rect 264 18882 296 18914
rect 336 18882 368 18914
rect 408 18882 440 18914
rect 480 18882 512 18914
rect 552 18882 584 18914
rect 624 18882 656 18914
rect 696 18882 728 18914
rect 768 18882 800 18914
rect 840 18882 872 18914
rect 912 18882 944 18914
rect 984 18882 1016 18914
rect 1056 18882 1088 18914
rect 1128 18882 1160 18914
rect 1200 18882 1232 18914
rect 1272 18882 1304 18914
rect 1344 18882 1376 18914
rect 1416 18882 1448 18914
rect 1488 18882 1520 18914
rect 1560 18882 1592 18914
rect 1632 18882 1664 18914
rect 1704 18882 1736 18914
rect 1776 18882 1808 18914
rect 1848 18882 1880 18914
rect 120 18810 152 18842
rect 192 18810 224 18842
rect 264 18810 296 18842
rect 336 18810 368 18842
rect 408 18810 440 18842
rect 480 18810 512 18842
rect 552 18810 584 18842
rect 624 18810 656 18842
rect 696 18810 728 18842
rect 768 18810 800 18842
rect 840 18810 872 18842
rect 912 18810 944 18842
rect 984 18810 1016 18842
rect 1056 18810 1088 18842
rect 1128 18810 1160 18842
rect 1200 18810 1232 18842
rect 1272 18810 1304 18842
rect 1344 18810 1376 18842
rect 1416 18810 1448 18842
rect 1488 18810 1520 18842
rect 1560 18810 1592 18842
rect 1632 18810 1664 18842
rect 1704 18810 1736 18842
rect 1776 18810 1808 18842
rect 1848 18810 1880 18842
rect 120 18738 152 18770
rect 192 18738 224 18770
rect 264 18738 296 18770
rect 336 18738 368 18770
rect 408 18738 440 18770
rect 480 18738 512 18770
rect 552 18738 584 18770
rect 624 18738 656 18770
rect 696 18738 728 18770
rect 768 18738 800 18770
rect 840 18738 872 18770
rect 912 18738 944 18770
rect 984 18738 1016 18770
rect 1056 18738 1088 18770
rect 1128 18738 1160 18770
rect 1200 18738 1232 18770
rect 1272 18738 1304 18770
rect 1344 18738 1376 18770
rect 1416 18738 1448 18770
rect 1488 18738 1520 18770
rect 1560 18738 1592 18770
rect 1632 18738 1664 18770
rect 1704 18738 1736 18770
rect 1776 18738 1808 18770
rect 1848 18738 1880 18770
rect 120 18666 152 18698
rect 192 18666 224 18698
rect 264 18666 296 18698
rect 336 18666 368 18698
rect 408 18666 440 18698
rect 480 18666 512 18698
rect 552 18666 584 18698
rect 624 18666 656 18698
rect 696 18666 728 18698
rect 768 18666 800 18698
rect 840 18666 872 18698
rect 912 18666 944 18698
rect 984 18666 1016 18698
rect 1056 18666 1088 18698
rect 1128 18666 1160 18698
rect 1200 18666 1232 18698
rect 1272 18666 1304 18698
rect 1344 18666 1376 18698
rect 1416 18666 1448 18698
rect 1488 18666 1520 18698
rect 1560 18666 1592 18698
rect 1632 18666 1664 18698
rect 1704 18666 1736 18698
rect 1776 18666 1808 18698
rect 1848 18666 1880 18698
rect 120 18594 152 18626
rect 192 18594 224 18626
rect 264 18594 296 18626
rect 336 18594 368 18626
rect 408 18594 440 18626
rect 480 18594 512 18626
rect 552 18594 584 18626
rect 624 18594 656 18626
rect 696 18594 728 18626
rect 768 18594 800 18626
rect 840 18594 872 18626
rect 912 18594 944 18626
rect 984 18594 1016 18626
rect 1056 18594 1088 18626
rect 1128 18594 1160 18626
rect 1200 18594 1232 18626
rect 1272 18594 1304 18626
rect 1344 18594 1376 18626
rect 1416 18594 1448 18626
rect 1488 18594 1520 18626
rect 1560 18594 1592 18626
rect 1632 18594 1664 18626
rect 1704 18594 1736 18626
rect 1776 18594 1808 18626
rect 1848 18594 1880 18626
rect 120 18522 152 18554
rect 192 18522 224 18554
rect 264 18522 296 18554
rect 336 18522 368 18554
rect 408 18522 440 18554
rect 480 18522 512 18554
rect 552 18522 584 18554
rect 624 18522 656 18554
rect 696 18522 728 18554
rect 768 18522 800 18554
rect 840 18522 872 18554
rect 912 18522 944 18554
rect 984 18522 1016 18554
rect 1056 18522 1088 18554
rect 1128 18522 1160 18554
rect 1200 18522 1232 18554
rect 1272 18522 1304 18554
rect 1344 18522 1376 18554
rect 1416 18522 1448 18554
rect 1488 18522 1520 18554
rect 1560 18522 1592 18554
rect 1632 18522 1664 18554
rect 1704 18522 1736 18554
rect 1776 18522 1808 18554
rect 1848 18522 1880 18554
rect 120 18450 152 18482
rect 192 18450 224 18482
rect 264 18450 296 18482
rect 336 18450 368 18482
rect 408 18450 440 18482
rect 480 18450 512 18482
rect 552 18450 584 18482
rect 624 18450 656 18482
rect 696 18450 728 18482
rect 768 18450 800 18482
rect 840 18450 872 18482
rect 912 18450 944 18482
rect 984 18450 1016 18482
rect 1056 18450 1088 18482
rect 1128 18450 1160 18482
rect 1200 18450 1232 18482
rect 1272 18450 1304 18482
rect 1344 18450 1376 18482
rect 1416 18450 1448 18482
rect 1488 18450 1520 18482
rect 1560 18450 1592 18482
rect 1632 18450 1664 18482
rect 1704 18450 1736 18482
rect 1776 18450 1808 18482
rect 1848 18450 1880 18482
rect 120 18378 152 18410
rect 192 18378 224 18410
rect 264 18378 296 18410
rect 336 18378 368 18410
rect 408 18378 440 18410
rect 480 18378 512 18410
rect 552 18378 584 18410
rect 624 18378 656 18410
rect 696 18378 728 18410
rect 768 18378 800 18410
rect 840 18378 872 18410
rect 912 18378 944 18410
rect 984 18378 1016 18410
rect 1056 18378 1088 18410
rect 1128 18378 1160 18410
rect 1200 18378 1232 18410
rect 1272 18378 1304 18410
rect 1344 18378 1376 18410
rect 1416 18378 1448 18410
rect 1488 18378 1520 18410
rect 1560 18378 1592 18410
rect 1632 18378 1664 18410
rect 1704 18378 1736 18410
rect 1776 18378 1808 18410
rect 1848 18378 1880 18410
rect 120 18306 152 18338
rect 192 18306 224 18338
rect 264 18306 296 18338
rect 336 18306 368 18338
rect 408 18306 440 18338
rect 480 18306 512 18338
rect 552 18306 584 18338
rect 624 18306 656 18338
rect 696 18306 728 18338
rect 768 18306 800 18338
rect 840 18306 872 18338
rect 912 18306 944 18338
rect 984 18306 1016 18338
rect 1056 18306 1088 18338
rect 1128 18306 1160 18338
rect 1200 18306 1232 18338
rect 1272 18306 1304 18338
rect 1344 18306 1376 18338
rect 1416 18306 1448 18338
rect 1488 18306 1520 18338
rect 1560 18306 1592 18338
rect 1632 18306 1664 18338
rect 1704 18306 1736 18338
rect 1776 18306 1808 18338
rect 1848 18306 1880 18338
rect 120 18234 152 18266
rect 192 18234 224 18266
rect 264 18234 296 18266
rect 336 18234 368 18266
rect 408 18234 440 18266
rect 480 18234 512 18266
rect 552 18234 584 18266
rect 624 18234 656 18266
rect 696 18234 728 18266
rect 768 18234 800 18266
rect 840 18234 872 18266
rect 912 18234 944 18266
rect 984 18234 1016 18266
rect 1056 18234 1088 18266
rect 1128 18234 1160 18266
rect 1200 18234 1232 18266
rect 1272 18234 1304 18266
rect 1344 18234 1376 18266
rect 1416 18234 1448 18266
rect 1488 18234 1520 18266
rect 1560 18234 1592 18266
rect 1632 18234 1664 18266
rect 1704 18234 1736 18266
rect 1776 18234 1808 18266
rect 1848 18234 1880 18266
rect 120 18162 152 18194
rect 192 18162 224 18194
rect 264 18162 296 18194
rect 336 18162 368 18194
rect 408 18162 440 18194
rect 480 18162 512 18194
rect 552 18162 584 18194
rect 624 18162 656 18194
rect 696 18162 728 18194
rect 768 18162 800 18194
rect 840 18162 872 18194
rect 912 18162 944 18194
rect 984 18162 1016 18194
rect 1056 18162 1088 18194
rect 1128 18162 1160 18194
rect 1200 18162 1232 18194
rect 1272 18162 1304 18194
rect 1344 18162 1376 18194
rect 1416 18162 1448 18194
rect 1488 18162 1520 18194
rect 1560 18162 1592 18194
rect 1632 18162 1664 18194
rect 1704 18162 1736 18194
rect 1776 18162 1808 18194
rect 1848 18162 1880 18194
rect 192 17816 224 17848
rect 264 17816 296 17848
rect 336 17816 368 17848
rect 408 17816 440 17848
rect 480 17816 512 17848
rect 552 17816 584 17848
rect 624 17816 656 17848
rect 696 17816 728 17848
rect 768 17816 800 17848
rect 840 17816 872 17848
rect 912 17816 944 17848
rect 984 17816 1016 17848
rect 1056 17816 1088 17848
rect 1128 17816 1160 17848
rect 1200 17816 1232 17848
rect 1272 17816 1304 17848
rect 1344 17816 1376 17848
rect 1416 17816 1448 17848
rect 1488 17816 1520 17848
rect 1560 17816 1592 17848
rect 1632 17816 1664 17848
rect 1704 17816 1736 17848
rect 1776 17816 1808 17848
rect 1848 17816 1880 17848
rect 120 17744 152 17776
rect 192 17744 224 17776
rect 264 17744 296 17776
rect 336 17744 368 17776
rect 408 17744 440 17776
rect 480 17744 512 17776
rect 552 17744 584 17776
rect 624 17744 656 17776
rect 696 17744 728 17776
rect 768 17744 800 17776
rect 840 17744 872 17776
rect 912 17744 944 17776
rect 984 17744 1016 17776
rect 1056 17744 1088 17776
rect 1128 17744 1160 17776
rect 1200 17744 1232 17776
rect 1272 17744 1304 17776
rect 1344 17744 1376 17776
rect 1416 17744 1448 17776
rect 1488 17744 1520 17776
rect 1560 17744 1592 17776
rect 1632 17744 1664 17776
rect 1704 17744 1736 17776
rect 1776 17744 1808 17776
rect 1848 17744 1880 17776
rect 120 17672 152 17704
rect 192 17672 224 17704
rect 264 17672 296 17704
rect 336 17672 368 17704
rect 408 17672 440 17704
rect 480 17672 512 17704
rect 552 17672 584 17704
rect 624 17672 656 17704
rect 696 17672 728 17704
rect 768 17672 800 17704
rect 840 17672 872 17704
rect 912 17672 944 17704
rect 984 17672 1016 17704
rect 1056 17672 1088 17704
rect 1128 17672 1160 17704
rect 1200 17672 1232 17704
rect 1272 17672 1304 17704
rect 1344 17672 1376 17704
rect 1416 17672 1448 17704
rect 1488 17672 1520 17704
rect 1560 17672 1592 17704
rect 1632 17672 1664 17704
rect 1704 17672 1736 17704
rect 1776 17672 1808 17704
rect 1848 17672 1880 17704
rect 120 17600 152 17632
rect 192 17600 224 17632
rect 264 17600 296 17632
rect 336 17600 368 17632
rect 408 17600 440 17632
rect 480 17600 512 17632
rect 552 17600 584 17632
rect 624 17600 656 17632
rect 696 17600 728 17632
rect 768 17600 800 17632
rect 840 17600 872 17632
rect 912 17600 944 17632
rect 984 17600 1016 17632
rect 1056 17600 1088 17632
rect 1128 17600 1160 17632
rect 1200 17600 1232 17632
rect 1272 17600 1304 17632
rect 1344 17600 1376 17632
rect 1416 17600 1448 17632
rect 1488 17600 1520 17632
rect 1560 17600 1592 17632
rect 1632 17600 1664 17632
rect 1704 17600 1736 17632
rect 1776 17600 1808 17632
rect 1848 17600 1880 17632
rect 120 17528 152 17560
rect 192 17528 224 17560
rect 264 17528 296 17560
rect 336 17528 368 17560
rect 408 17528 440 17560
rect 480 17528 512 17560
rect 552 17528 584 17560
rect 624 17528 656 17560
rect 696 17528 728 17560
rect 768 17528 800 17560
rect 840 17528 872 17560
rect 912 17528 944 17560
rect 984 17528 1016 17560
rect 1056 17528 1088 17560
rect 1128 17528 1160 17560
rect 1200 17528 1232 17560
rect 1272 17528 1304 17560
rect 1344 17528 1376 17560
rect 1416 17528 1448 17560
rect 1488 17528 1520 17560
rect 1560 17528 1592 17560
rect 1632 17528 1664 17560
rect 1704 17528 1736 17560
rect 1776 17528 1808 17560
rect 1848 17528 1880 17560
rect 120 17456 152 17488
rect 192 17456 224 17488
rect 264 17456 296 17488
rect 336 17456 368 17488
rect 408 17456 440 17488
rect 480 17456 512 17488
rect 552 17456 584 17488
rect 624 17456 656 17488
rect 696 17456 728 17488
rect 768 17456 800 17488
rect 840 17456 872 17488
rect 912 17456 944 17488
rect 984 17456 1016 17488
rect 1056 17456 1088 17488
rect 1128 17456 1160 17488
rect 1200 17456 1232 17488
rect 1272 17456 1304 17488
rect 1344 17456 1376 17488
rect 1416 17456 1448 17488
rect 1488 17456 1520 17488
rect 1560 17456 1592 17488
rect 1632 17456 1664 17488
rect 1704 17456 1736 17488
rect 1776 17456 1808 17488
rect 1848 17456 1880 17488
rect 120 17384 152 17416
rect 192 17384 224 17416
rect 264 17384 296 17416
rect 336 17384 368 17416
rect 408 17384 440 17416
rect 480 17384 512 17416
rect 552 17384 584 17416
rect 624 17384 656 17416
rect 696 17384 728 17416
rect 768 17384 800 17416
rect 840 17384 872 17416
rect 912 17384 944 17416
rect 984 17384 1016 17416
rect 1056 17384 1088 17416
rect 1128 17384 1160 17416
rect 1200 17384 1232 17416
rect 1272 17384 1304 17416
rect 1344 17384 1376 17416
rect 1416 17384 1448 17416
rect 1488 17384 1520 17416
rect 1560 17384 1592 17416
rect 1632 17384 1664 17416
rect 1704 17384 1736 17416
rect 1776 17384 1808 17416
rect 1848 17384 1880 17416
rect 120 17312 152 17344
rect 192 17312 224 17344
rect 264 17312 296 17344
rect 336 17312 368 17344
rect 408 17312 440 17344
rect 480 17312 512 17344
rect 552 17312 584 17344
rect 624 17312 656 17344
rect 696 17312 728 17344
rect 768 17312 800 17344
rect 840 17312 872 17344
rect 912 17312 944 17344
rect 984 17312 1016 17344
rect 1056 17312 1088 17344
rect 1128 17312 1160 17344
rect 1200 17312 1232 17344
rect 1272 17312 1304 17344
rect 1344 17312 1376 17344
rect 1416 17312 1448 17344
rect 1488 17312 1520 17344
rect 1560 17312 1592 17344
rect 1632 17312 1664 17344
rect 1704 17312 1736 17344
rect 1776 17312 1808 17344
rect 1848 17312 1880 17344
rect 120 17240 152 17272
rect 192 17240 224 17272
rect 264 17240 296 17272
rect 336 17240 368 17272
rect 408 17240 440 17272
rect 480 17240 512 17272
rect 552 17240 584 17272
rect 624 17240 656 17272
rect 696 17240 728 17272
rect 768 17240 800 17272
rect 840 17240 872 17272
rect 912 17240 944 17272
rect 984 17240 1016 17272
rect 1056 17240 1088 17272
rect 1128 17240 1160 17272
rect 1200 17240 1232 17272
rect 1272 17240 1304 17272
rect 1344 17240 1376 17272
rect 1416 17240 1448 17272
rect 1488 17240 1520 17272
rect 1560 17240 1592 17272
rect 1632 17240 1664 17272
rect 1704 17240 1736 17272
rect 1776 17240 1808 17272
rect 1848 17240 1880 17272
rect 120 17168 152 17200
rect 192 17168 224 17200
rect 264 17168 296 17200
rect 336 17168 368 17200
rect 408 17168 440 17200
rect 480 17168 512 17200
rect 552 17168 584 17200
rect 624 17168 656 17200
rect 696 17168 728 17200
rect 768 17168 800 17200
rect 840 17168 872 17200
rect 912 17168 944 17200
rect 984 17168 1016 17200
rect 1056 17168 1088 17200
rect 1128 17168 1160 17200
rect 1200 17168 1232 17200
rect 1272 17168 1304 17200
rect 1344 17168 1376 17200
rect 1416 17168 1448 17200
rect 1488 17168 1520 17200
rect 1560 17168 1592 17200
rect 1632 17168 1664 17200
rect 1704 17168 1736 17200
rect 1776 17168 1808 17200
rect 1848 17168 1880 17200
rect 120 17096 152 17128
rect 192 17096 224 17128
rect 264 17096 296 17128
rect 336 17096 368 17128
rect 408 17096 440 17128
rect 480 17096 512 17128
rect 552 17096 584 17128
rect 624 17096 656 17128
rect 696 17096 728 17128
rect 768 17096 800 17128
rect 840 17096 872 17128
rect 912 17096 944 17128
rect 984 17096 1016 17128
rect 1056 17096 1088 17128
rect 1128 17096 1160 17128
rect 1200 17096 1232 17128
rect 1272 17096 1304 17128
rect 1344 17096 1376 17128
rect 1416 17096 1448 17128
rect 1488 17096 1520 17128
rect 1560 17096 1592 17128
rect 1632 17096 1664 17128
rect 1704 17096 1736 17128
rect 1776 17096 1808 17128
rect 1848 17096 1880 17128
rect 120 17024 152 17056
rect 192 17024 224 17056
rect 264 17024 296 17056
rect 336 17024 368 17056
rect 408 17024 440 17056
rect 480 17024 512 17056
rect 552 17024 584 17056
rect 624 17024 656 17056
rect 696 17024 728 17056
rect 768 17024 800 17056
rect 840 17024 872 17056
rect 912 17024 944 17056
rect 984 17024 1016 17056
rect 1056 17024 1088 17056
rect 1128 17024 1160 17056
rect 1200 17024 1232 17056
rect 1272 17024 1304 17056
rect 1344 17024 1376 17056
rect 1416 17024 1448 17056
rect 1488 17024 1520 17056
rect 1560 17024 1592 17056
rect 1632 17024 1664 17056
rect 1704 17024 1736 17056
rect 1776 17024 1808 17056
rect 1848 17024 1880 17056
rect 120 16952 152 16984
rect 192 16952 224 16984
rect 264 16952 296 16984
rect 336 16952 368 16984
rect 408 16952 440 16984
rect 480 16952 512 16984
rect 552 16952 584 16984
rect 624 16952 656 16984
rect 696 16952 728 16984
rect 768 16952 800 16984
rect 840 16952 872 16984
rect 912 16952 944 16984
rect 984 16952 1016 16984
rect 1056 16952 1088 16984
rect 1128 16952 1160 16984
rect 1200 16952 1232 16984
rect 1272 16952 1304 16984
rect 1344 16952 1376 16984
rect 1416 16952 1448 16984
rect 1488 16952 1520 16984
rect 1560 16952 1592 16984
rect 1632 16952 1664 16984
rect 1704 16952 1736 16984
rect 1776 16952 1808 16984
rect 1848 16952 1880 16984
rect 120 16880 152 16912
rect 192 16880 224 16912
rect 264 16880 296 16912
rect 336 16880 368 16912
rect 408 16880 440 16912
rect 480 16880 512 16912
rect 552 16880 584 16912
rect 624 16880 656 16912
rect 696 16880 728 16912
rect 768 16880 800 16912
rect 840 16880 872 16912
rect 912 16880 944 16912
rect 984 16880 1016 16912
rect 1056 16880 1088 16912
rect 1128 16880 1160 16912
rect 1200 16880 1232 16912
rect 1272 16880 1304 16912
rect 1344 16880 1376 16912
rect 1416 16880 1448 16912
rect 1488 16880 1520 16912
rect 1560 16880 1592 16912
rect 1632 16880 1664 16912
rect 1704 16880 1736 16912
rect 1776 16880 1808 16912
rect 1848 16880 1880 16912
rect 120 16808 152 16840
rect 192 16808 224 16840
rect 264 16808 296 16840
rect 336 16808 368 16840
rect 408 16808 440 16840
rect 480 16808 512 16840
rect 552 16808 584 16840
rect 624 16808 656 16840
rect 696 16808 728 16840
rect 768 16808 800 16840
rect 840 16808 872 16840
rect 912 16808 944 16840
rect 984 16808 1016 16840
rect 1056 16808 1088 16840
rect 1128 16808 1160 16840
rect 1200 16808 1232 16840
rect 1272 16808 1304 16840
rect 1344 16808 1376 16840
rect 1416 16808 1448 16840
rect 1488 16808 1520 16840
rect 1560 16808 1592 16840
rect 1632 16808 1664 16840
rect 1704 16808 1736 16840
rect 1776 16808 1808 16840
rect 1848 16808 1880 16840
rect 120 16736 152 16768
rect 192 16736 224 16768
rect 264 16736 296 16768
rect 336 16736 368 16768
rect 408 16736 440 16768
rect 480 16736 512 16768
rect 552 16736 584 16768
rect 624 16736 656 16768
rect 696 16736 728 16768
rect 768 16736 800 16768
rect 840 16736 872 16768
rect 912 16736 944 16768
rect 984 16736 1016 16768
rect 1056 16736 1088 16768
rect 1128 16736 1160 16768
rect 1200 16736 1232 16768
rect 1272 16736 1304 16768
rect 1344 16736 1376 16768
rect 1416 16736 1448 16768
rect 1488 16736 1520 16768
rect 1560 16736 1592 16768
rect 1632 16736 1664 16768
rect 1704 16736 1736 16768
rect 1776 16736 1808 16768
rect 1848 16736 1880 16768
rect 120 16664 152 16696
rect 192 16664 224 16696
rect 264 16664 296 16696
rect 336 16664 368 16696
rect 408 16664 440 16696
rect 480 16664 512 16696
rect 552 16664 584 16696
rect 624 16664 656 16696
rect 696 16664 728 16696
rect 768 16664 800 16696
rect 840 16664 872 16696
rect 912 16664 944 16696
rect 984 16664 1016 16696
rect 1056 16664 1088 16696
rect 1128 16664 1160 16696
rect 1200 16664 1232 16696
rect 1272 16664 1304 16696
rect 1344 16664 1376 16696
rect 1416 16664 1448 16696
rect 1488 16664 1520 16696
rect 1560 16664 1592 16696
rect 1632 16664 1664 16696
rect 1704 16664 1736 16696
rect 1776 16664 1808 16696
rect 1848 16664 1880 16696
rect 120 16592 152 16624
rect 192 16592 224 16624
rect 264 16592 296 16624
rect 336 16592 368 16624
rect 408 16592 440 16624
rect 480 16592 512 16624
rect 552 16592 584 16624
rect 624 16592 656 16624
rect 696 16592 728 16624
rect 768 16592 800 16624
rect 840 16592 872 16624
rect 912 16592 944 16624
rect 984 16592 1016 16624
rect 1056 16592 1088 16624
rect 1128 16592 1160 16624
rect 1200 16592 1232 16624
rect 1272 16592 1304 16624
rect 1344 16592 1376 16624
rect 1416 16592 1448 16624
rect 1488 16592 1520 16624
rect 1560 16592 1592 16624
rect 1632 16592 1664 16624
rect 1704 16592 1736 16624
rect 1776 16592 1808 16624
rect 1848 16592 1880 16624
rect 120 16520 152 16552
rect 192 16520 224 16552
rect 264 16520 296 16552
rect 336 16520 368 16552
rect 408 16520 440 16552
rect 480 16520 512 16552
rect 552 16520 584 16552
rect 624 16520 656 16552
rect 696 16520 728 16552
rect 768 16520 800 16552
rect 840 16520 872 16552
rect 912 16520 944 16552
rect 984 16520 1016 16552
rect 1056 16520 1088 16552
rect 1128 16520 1160 16552
rect 1200 16520 1232 16552
rect 1272 16520 1304 16552
rect 1344 16520 1376 16552
rect 1416 16520 1448 16552
rect 1488 16520 1520 16552
rect 1560 16520 1592 16552
rect 1632 16520 1664 16552
rect 1704 16520 1736 16552
rect 1776 16520 1808 16552
rect 1848 16520 1880 16552
rect 120 16448 152 16480
rect 192 16448 224 16480
rect 264 16448 296 16480
rect 336 16448 368 16480
rect 408 16448 440 16480
rect 480 16448 512 16480
rect 552 16448 584 16480
rect 624 16448 656 16480
rect 696 16448 728 16480
rect 768 16448 800 16480
rect 840 16448 872 16480
rect 912 16448 944 16480
rect 984 16448 1016 16480
rect 1056 16448 1088 16480
rect 1128 16448 1160 16480
rect 1200 16448 1232 16480
rect 1272 16448 1304 16480
rect 1344 16448 1376 16480
rect 1416 16448 1448 16480
rect 1488 16448 1520 16480
rect 1560 16448 1592 16480
rect 1632 16448 1664 16480
rect 1704 16448 1736 16480
rect 1776 16448 1808 16480
rect 1848 16448 1880 16480
rect 120 16376 152 16408
rect 192 16376 224 16408
rect 264 16376 296 16408
rect 336 16376 368 16408
rect 408 16376 440 16408
rect 480 16376 512 16408
rect 552 16376 584 16408
rect 624 16376 656 16408
rect 696 16376 728 16408
rect 768 16376 800 16408
rect 840 16376 872 16408
rect 912 16376 944 16408
rect 984 16376 1016 16408
rect 1056 16376 1088 16408
rect 1128 16376 1160 16408
rect 1200 16376 1232 16408
rect 1272 16376 1304 16408
rect 1344 16376 1376 16408
rect 1416 16376 1448 16408
rect 1488 16376 1520 16408
rect 1560 16376 1592 16408
rect 1632 16376 1664 16408
rect 1704 16376 1736 16408
rect 1776 16376 1808 16408
rect 1848 16376 1880 16408
rect 120 16304 152 16336
rect 192 16304 224 16336
rect 264 16304 296 16336
rect 336 16304 368 16336
rect 408 16304 440 16336
rect 480 16304 512 16336
rect 552 16304 584 16336
rect 624 16304 656 16336
rect 696 16304 728 16336
rect 768 16304 800 16336
rect 840 16304 872 16336
rect 912 16304 944 16336
rect 984 16304 1016 16336
rect 1056 16304 1088 16336
rect 1128 16304 1160 16336
rect 1200 16304 1232 16336
rect 1272 16304 1304 16336
rect 1344 16304 1376 16336
rect 1416 16304 1448 16336
rect 1488 16304 1520 16336
rect 1560 16304 1592 16336
rect 1632 16304 1664 16336
rect 1704 16304 1736 16336
rect 1776 16304 1808 16336
rect 1848 16304 1880 16336
rect 120 16232 152 16264
rect 192 16232 224 16264
rect 264 16232 296 16264
rect 336 16232 368 16264
rect 408 16232 440 16264
rect 480 16232 512 16264
rect 552 16232 584 16264
rect 624 16232 656 16264
rect 696 16232 728 16264
rect 768 16232 800 16264
rect 840 16232 872 16264
rect 912 16232 944 16264
rect 984 16232 1016 16264
rect 1056 16232 1088 16264
rect 1128 16232 1160 16264
rect 1200 16232 1232 16264
rect 1272 16232 1304 16264
rect 1344 16232 1376 16264
rect 1416 16232 1448 16264
rect 1488 16232 1520 16264
rect 1560 16232 1592 16264
rect 1632 16232 1664 16264
rect 1704 16232 1736 16264
rect 1776 16232 1808 16264
rect 1848 16232 1880 16264
rect 120 16160 152 16192
rect 192 16160 224 16192
rect 264 16160 296 16192
rect 336 16160 368 16192
rect 408 16160 440 16192
rect 480 16160 512 16192
rect 552 16160 584 16192
rect 624 16160 656 16192
rect 696 16160 728 16192
rect 768 16160 800 16192
rect 840 16160 872 16192
rect 912 16160 944 16192
rect 984 16160 1016 16192
rect 1056 16160 1088 16192
rect 1128 16160 1160 16192
rect 1200 16160 1232 16192
rect 1272 16160 1304 16192
rect 1344 16160 1376 16192
rect 1416 16160 1448 16192
rect 1488 16160 1520 16192
rect 1560 16160 1592 16192
rect 1632 16160 1664 16192
rect 1704 16160 1736 16192
rect 1776 16160 1808 16192
rect 1848 16160 1880 16192
rect 120 16088 152 16120
rect 192 16088 224 16120
rect 264 16088 296 16120
rect 336 16088 368 16120
rect 408 16088 440 16120
rect 480 16088 512 16120
rect 552 16088 584 16120
rect 624 16088 656 16120
rect 696 16088 728 16120
rect 768 16088 800 16120
rect 840 16088 872 16120
rect 912 16088 944 16120
rect 984 16088 1016 16120
rect 1056 16088 1088 16120
rect 1128 16088 1160 16120
rect 1200 16088 1232 16120
rect 1272 16088 1304 16120
rect 1344 16088 1376 16120
rect 1416 16088 1448 16120
rect 1488 16088 1520 16120
rect 1560 16088 1592 16120
rect 1632 16088 1664 16120
rect 1704 16088 1736 16120
rect 1776 16088 1808 16120
rect 1848 16088 1880 16120
rect 120 16016 152 16048
rect 192 16016 224 16048
rect 264 16016 296 16048
rect 336 16016 368 16048
rect 408 16016 440 16048
rect 480 16016 512 16048
rect 552 16016 584 16048
rect 624 16016 656 16048
rect 696 16016 728 16048
rect 768 16016 800 16048
rect 840 16016 872 16048
rect 912 16016 944 16048
rect 984 16016 1016 16048
rect 1056 16016 1088 16048
rect 1128 16016 1160 16048
rect 1200 16016 1232 16048
rect 1272 16016 1304 16048
rect 1344 16016 1376 16048
rect 1416 16016 1448 16048
rect 1488 16016 1520 16048
rect 1560 16016 1592 16048
rect 1632 16016 1664 16048
rect 1704 16016 1736 16048
rect 1776 16016 1808 16048
rect 1848 16016 1880 16048
rect 120 15944 152 15976
rect 192 15944 224 15976
rect 264 15944 296 15976
rect 336 15944 368 15976
rect 408 15944 440 15976
rect 480 15944 512 15976
rect 552 15944 584 15976
rect 624 15944 656 15976
rect 696 15944 728 15976
rect 768 15944 800 15976
rect 840 15944 872 15976
rect 912 15944 944 15976
rect 984 15944 1016 15976
rect 1056 15944 1088 15976
rect 1128 15944 1160 15976
rect 1200 15944 1232 15976
rect 1272 15944 1304 15976
rect 1344 15944 1376 15976
rect 1416 15944 1448 15976
rect 1488 15944 1520 15976
rect 1560 15944 1592 15976
rect 1632 15944 1664 15976
rect 1704 15944 1736 15976
rect 1776 15944 1808 15976
rect 1848 15944 1880 15976
rect 120 15872 152 15904
rect 192 15872 224 15904
rect 264 15872 296 15904
rect 336 15872 368 15904
rect 408 15872 440 15904
rect 480 15872 512 15904
rect 552 15872 584 15904
rect 624 15872 656 15904
rect 696 15872 728 15904
rect 768 15872 800 15904
rect 840 15872 872 15904
rect 912 15872 944 15904
rect 984 15872 1016 15904
rect 1056 15872 1088 15904
rect 1128 15872 1160 15904
rect 1200 15872 1232 15904
rect 1272 15872 1304 15904
rect 1344 15872 1376 15904
rect 1416 15872 1448 15904
rect 1488 15872 1520 15904
rect 1560 15872 1592 15904
rect 1632 15872 1664 15904
rect 1704 15872 1736 15904
rect 1776 15872 1808 15904
rect 1848 15872 1880 15904
rect 120 15800 152 15832
rect 192 15800 224 15832
rect 264 15800 296 15832
rect 336 15800 368 15832
rect 408 15800 440 15832
rect 480 15800 512 15832
rect 552 15800 584 15832
rect 624 15800 656 15832
rect 696 15800 728 15832
rect 768 15800 800 15832
rect 840 15800 872 15832
rect 912 15800 944 15832
rect 984 15800 1016 15832
rect 1056 15800 1088 15832
rect 1128 15800 1160 15832
rect 1200 15800 1232 15832
rect 1272 15800 1304 15832
rect 1344 15800 1376 15832
rect 1416 15800 1448 15832
rect 1488 15800 1520 15832
rect 1560 15800 1592 15832
rect 1632 15800 1664 15832
rect 1704 15800 1736 15832
rect 1776 15800 1808 15832
rect 1848 15800 1880 15832
rect 120 15728 152 15760
rect 192 15728 224 15760
rect 264 15728 296 15760
rect 336 15728 368 15760
rect 408 15728 440 15760
rect 480 15728 512 15760
rect 552 15728 584 15760
rect 624 15728 656 15760
rect 696 15728 728 15760
rect 768 15728 800 15760
rect 840 15728 872 15760
rect 912 15728 944 15760
rect 984 15728 1016 15760
rect 1056 15728 1088 15760
rect 1128 15728 1160 15760
rect 1200 15728 1232 15760
rect 1272 15728 1304 15760
rect 1344 15728 1376 15760
rect 1416 15728 1448 15760
rect 1488 15728 1520 15760
rect 1560 15728 1592 15760
rect 1632 15728 1664 15760
rect 1704 15728 1736 15760
rect 1776 15728 1808 15760
rect 1848 15728 1880 15760
rect 120 15656 152 15688
rect 192 15656 224 15688
rect 264 15656 296 15688
rect 336 15656 368 15688
rect 408 15656 440 15688
rect 480 15656 512 15688
rect 552 15656 584 15688
rect 624 15656 656 15688
rect 696 15656 728 15688
rect 768 15656 800 15688
rect 840 15656 872 15688
rect 912 15656 944 15688
rect 984 15656 1016 15688
rect 1056 15656 1088 15688
rect 1128 15656 1160 15688
rect 1200 15656 1232 15688
rect 1272 15656 1304 15688
rect 1344 15656 1376 15688
rect 1416 15656 1448 15688
rect 1488 15656 1520 15688
rect 1560 15656 1592 15688
rect 1632 15656 1664 15688
rect 1704 15656 1736 15688
rect 1776 15656 1808 15688
rect 1848 15656 1880 15688
rect 120 15584 152 15616
rect 192 15584 224 15616
rect 264 15584 296 15616
rect 336 15584 368 15616
rect 408 15584 440 15616
rect 480 15584 512 15616
rect 552 15584 584 15616
rect 624 15584 656 15616
rect 696 15584 728 15616
rect 768 15584 800 15616
rect 840 15584 872 15616
rect 912 15584 944 15616
rect 984 15584 1016 15616
rect 1056 15584 1088 15616
rect 1128 15584 1160 15616
rect 1200 15584 1232 15616
rect 1272 15584 1304 15616
rect 1344 15584 1376 15616
rect 1416 15584 1448 15616
rect 1488 15584 1520 15616
rect 1560 15584 1592 15616
rect 1632 15584 1664 15616
rect 1704 15584 1736 15616
rect 1776 15584 1808 15616
rect 1848 15584 1880 15616
rect 120 15512 152 15544
rect 192 15512 224 15544
rect 264 15512 296 15544
rect 336 15512 368 15544
rect 408 15512 440 15544
rect 480 15512 512 15544
rect 552 15512 584 15544
rect 624 15512 656 15544
rect 696 15512 728 15544
rect 768 15512 800 15544
rect 840 15512 872 15544
rect 912 15512 944 15544
rect 984 15512 1016 15544
rect 1056 15512 1088 15544
rect 1128 15512 1160 15544
rect 1200 15512 1232 15544
rect 1272 15512 1304 15544
rect 1344 15512 1376 15544
rect 1416 15512 1448 15544
rect 1488 15512 1520 15544
rect 1560 15512 1592 15544
rect 1632 15512 1664 15544
rect 1704 15512 1736 15544
rect 1776 15512 1808 15544
rect 1848 15512 1880 15544
rect 120 15440 152 15472
rect 192 15440 224 15472
rect 264 15440 296 15472
rect 336 15440 368 15472
rect 408 15440 440 15472
rect 480 15440 512 15472
rect 552 15440 584 15472
rect 624 15440 656 15472
rect 696 15440 728 15472
rect 768 15440 800 15472
rect 840 15440 872 15472
rect 912 15440 944 15472
rect 984 15440 1016 15472
rect 1056 15440 1088 15472
rect 1128 15440 1160 15472
rect 1200 15440 1232 15472
rect 1272 15440 1304 15472
rect 1344 15440 1376 15472
rect 1416 15440 1448 15472
rect 1488 15440 1520 15472
rect 1560 15440 1592 15472
rect 1632 15440 1664 15472
rect 1704 15440 1736 15472
rect 1776 15440 1808 15472
rect 1848 15440 1880 15472
rect 120 15368 152 15400
rect 192 15368 224 15400
rect 264 15368 296 15400
rect 336 15368 368 15400
rect 408 15368 440 15400
rect 480 15368 512 15400
rect 552 15368 584 15400
rect 624 15368 656 15400
rect 696 15368 728 15400
rect 768 15368 800 15400
rect 840 15368 872 15400
rect 912 15368 944 15400
rect 984 15368 1016 15400
rect 1056 15368 1088 15400
rect 1128 15368 1160 15400
rect 1200 15368 1232 15400
rect 1272 15368 1304 15400
rect 1344 15368 1376 15400
rect 1416 15368 1448 15400
rect 1488 15368 1520 15400
rect 1560 15368 1592 15400
rect 1632 15368 1664 15400
rect 1704 15368 1736 15400
rect 1776 15368 1808 15400
rect 1848 15368 1880 15400
rect 120 15296 152 15328
rect 192 15296 224 15328
rect 264 15296 296 15328
rect 336 15296 368 15328
rect 408 15296 440 15328
rect 480 15296 512 15328
rect 552 15296 584 15328
rect 624 15296 656 15328
rect 696 15296 728 15328
rect 768 15296 800 15328
rect 840 15296 872 15328
rect 912 15296 944 15328
rect 984 15296 1016 15328
rect 1056 15296 1088 15328
rect 1128 15296 1160 15328
rect 1200 15296 1232 15328
rect 1272 15296 1304 15328
rect 1344 15296 1376 15328
rect 1416 15296 1448 15328
rect 1488 15296 1520 15328
rect 1560 15296 1592 15328
rect 1632 15296 1664 15328
rect 1704 15296 1736 15328
rect 1776 15296 1808 15328
rect 1848 15296 1880 15328
rect 120 15224 152 15256
rect 192 15224 224 15256
rect 264 15224 296 15256
rect 336 15224 368 15256
rect 408 15224 440 15256
rect 480 15224 512 15256
rect 552 15224 584 15256
rect 624 15224 656 15256
rect 696 15224 728 15256
rect 768 15224 800 15256
rect 840 15224 872 15256
rect 912 15224 944 15256
rect 984 15224 1016 15256
rect 1056 15224 1088 15256
rect 1128 15224 1160 15256
rect 1200 15224 1232 15256
rect 1272 15224 1304 15256
rect 1344 15224 1376 15256
rect 1416 15224 1448 15256
rect 1488 15224 1520 15256
rect 1560 15224 1592 15256
rect 1632 15224 1664 15256
rect 1704 15224 1736 15256
rect 1776 15224 1808 15256
rect 1848 15224 1880 15256
rect 120 15152 152 15184
rect 192 15152 224 15184
rect 264 15152 296 15184
rect 336 15152 368 15184
rect 408 15152 440 15184
rect 480 15152 512 15184
rect 552 15152 584 15184
rect 624 15152 656 15184
rect 696 15152 728 15184
rect 768 15152 800 15184
rect 840 15152 872 15184
rect 912 15152 944 15184
rect 984 15152 1016 15184
rect 1056 15152 1088 15184
rect 1128 15152 1160 15184
rect 1200 15152 1232 15184
rect 1272 15152 1304 15184
rect 1344 15152 1376 15184
rect 1416 15152 1448 15184
rect 1488 15152 1520 15184
rect 1560 15152 1592 15184
rect 1632 15152 1664 15184
rect 1704 15152 1736 15184
rect 1776 15152 1808 15184
rect 1848 15152 1880 15184
rect 120 15080 152 15112
rect 192 15080 224 15112
rect 264 15080 296 15112
rect 336 15080 368 15112
rect 408 15080 440 15112
rect 480 15080 512 15112
rect 552 15080 584 15112
rect 624 15080 656 15112
rect 696 15080 728 15112
rect 768 15080 800 15112
rect 840 15080 872 15112
rect 912 15080 944 15112
rect 984 15080 1016 15112
rect 1056 15080 1088 15112
rect 1128 15080 1160 15112
rect 1200 15080 1232 15112
rect 1272 15080 1304 15112
rect 1344 15080 1376 15112
rect 1416 15080 1448 15112
rect 1488 15080 1520 15112
rect 1560 15080 1592 15112
rect 1632 15080 1664 15112
rect 1704 15080 1736 15112
rect 1776 15080 1808 15112
rect 1848 15080 1880 15112
rect 120 15008 152 15040
rect 192 15008 224 15040
rect 264 15008 296 15040
rect 336 15008 368 15040
rect 408 15008 440 15040
rect 480 15008 512 15040
rect 552 15008 584 15040
rect 624 15008 656 15040
rect 696 15008 728 15040
rect 768 15008 800 15040
rect 840 15008 872 15040
rect 912 15008 944 15040
rect 984 15008 1016 15040
rect 1056 15008 1088 15040
rect 1128 15008 1160 15040
rect 1200 15008 1232 15040
rect 1272 15008 1304 15040
rect 1344 15008 1376 15040
rect 1416 15008 1448 15040
rect 1488 15008 1520 15040
rect 1560 15008 1592 15040
rect 1632 15008 1664 15040
rect 1704 15008 1736 15040
rect 1776 15008 1808 15040
rect 1848 15008 1880 15040
rect 120 14936 152 14968
rect 192 14936 224 14968
rect 264 14936 296 14968
rect 336 14936 368 14968
rect 408 14936 440 14968
rect 480 14936 512 14968
rect 552 14936 584 14968
rect 624 14936 656 14968
rect 696 14936 728 14968
rect 768 14936 800 14968
rect 840 14936 872 14968
rect 912 14936 944 14968
rect 984 14936 1016 14968
rect 1056 14936 1088 14968
rect 1128 14936 1160 14968
rect 1200 14936 1232 14968
rect 1272 14936 1304 14968
rect 1344 14936 1376 14968
rect 1416 14936 1448 14968
rect 1488 14936 1520 14968
rect 1560 14936 1592 14968
rect 1632 14936 1664 14968
rect 1704 14936 1736 14968
rect 1776 14936 1808 14968
rect 1848 14936 1880 14968
rect 120 14864 152 14896
rect 192 14864 224 14896
rect 264 14864 296 14896
rect 336 14864 368 14896
rect 408 14864 440 14896
rect 480 14864 512 14896
rect 552 14864 584 14896
rect 624 14864 656 14896
rect 696 14864 728 14896
rect 768 14864 800 14896
rect 840 14864 872 14896
rect 912 14864 944 14896
rect 984 14864 1016 14896
rect 1056 14864 1088 14896
rect 1128 14864 1160 14896
rect 1200 14864 1232 14896
rect 1272 14864 1304 14896
rect 1344 14864 1376 14896
rect 1416 14864 1448 14896
rect 1488 14864 1520 14896
rect 1560 14864 1592 14896
rect 1632 14864 1664 14896
rect 1704 14864 1736 14896
rect 1776 14864 1808 14896
rect 1848 14864 1880 14896
rect 120 14792 152 14824
rect 192 14792 224 14824
rect 264 14792 296 14824
rect 336 14792 368 14824
rect 408 14792 440 14824
rect 480 14792 512 14824
rect 552 14792 584 14824
rect 624 14792 656 14824
rect 696 14792 728 14824
rect 768 14792 800 14824
rect 840 14792 872 14824
rect 912 14792 944 14824
rect 984 14792 1016 14824
rect 1056 14792 1088 14824
rect 1128 14792 1160 14824
rect 1200 14792 1232 14824
rect 1272 14792 1304 14824
rect 1344 14792 1376 14824
rect 1416 14792 1448 14824
rect 1488 14792 1520 14824
rect 1560 14792 1592 14824
rect 1632 14792 1664 14824
rect 1704 14792 1736 14824
rect 1776 14792 1808 14824
rect 1848 14792 1880 14824
rect 120 14720 152 14752
rect 192 14720 224 14752
rect 264 14720 296 14752
rect 336 14720 368 14752
rect 408 14720 440 14752
rect 480 14720 512 14752
rect 552 14720 584 14752
rect 624 14720 656 14752
rect 696 14720 728 14752
rect 768 14720 800 14752
rect 840 14720 872 14752
rect 912 14720 944 14752
rect 984 14720 1016 14752
rect 1056 14720 1088 14752
rect 1128 14720 1160 14752
rect 1200 14720 1232 14752
rect 1272 14720 1304 14752
rect 1344 14720 1376 14752
rect 1416 14720 1448 14752
rect 1488 14720 1520 14752
rect 1560 14720 1592 14752
rect 1632 14720 1664 14752
rect 1704 14720 1736 14752
rect 1776 14720 1808 14752
rect 1848 14720 1880 14752
rect 120 14648 152 14680
rect 192 14648 224 14680
rect 264 14648 296 14680
rect 336 14648 368 14680
rect 408 14648 440 14680
rect 480 14648 512 14680
rect 552 14648 584 14680
rect 624 14648 656 14680
rect 696 14648 728 14680
rect 768 14648 800 14680
rect 840 14648 872 14680
rect 912 14648 944 14680
rect 984 14648 1016 14680
rect 1056 14648 1088 14680
rect 1128 14648 1160 14680
rect 1200 14648 1232 14680
rect 1272 14648 1304 14680
rect 1344 14648 1376 14680
rect 1416 14648 1448 14680
rect 1488 14648 1520 14680
rect 1560 14648 1592 14680
rect 1632 14648 1664 14680
rect 1704 14648 1736 14680
rect 1776 14648 1808 14680
rect 1848 14648 1880 14680
rect 120 14576 152 14608
rect 192 14576 224 14608
rect 264 14576 296 14608
rect 336 14576 368 14608
rect 408 14576 440 14608
rect 480 14576 512 14608
rect 552 14576 584 14608
rect 624 14576 656 14608
rect 696 14576 728 14608
rect 768 14576 800 14608
rect 840 14576 872 14608
rect 912 14576 944 14608
rect 984 14576 1016 14608
rect 1056 14576 1088 14608
rect 1128 14576 1160 14608
rect 1200 14576 1232 14608
rect 1272 14576 1304 14608
rect 1344 14576 1376 14608
rect 1416 14576 1448 14608
rect 1488 14576 1520 14608
rect 1560 14576 1592 14608
rect 1632 14576 1664 14608
rect 1704 14576 1736 14608
rect 1776 14576 1808 14608
rect 1848 14576 1880 14608
rect 120 14504 152 14536
rect 192 14504 224 14536
rect 264 14504 296 14536
rect 336 14504 368 14536
rect 408 14504 440 14536
rect 480 14504 512 14536
rect 552 14504 584 14536
rect 624 14504 656 14536
rect 696 14504 728 14536
rect 768 14504 800 14536
rect 840 14504 872 14536
rect 912 14504 944 14536
rect 984 14504 1016 14536
rect 1056 14504 1088 14536
rect 1128 14504 1160 14536
rect 1200 14504 1232 14536
rect 1272 14504 1304 14536
rect 1344 14504 1376 14536
rect 1416 14504 1448 14536
rect 1488 14504 1520 14536
rect 1560 14504 1592 14536
rect 1632 14504 1664 14536
rect 1704 14504 1736 14536
rect 1776 14504 1808 14536
rect 1848 14504 1880 14536
rect 120 14432 152 14464
rect 192 14432 224 14464
rect 264 14432 296 14464
rect 336 14432 368 14464
rect 408 14432 440 14464
rect 480 14432 512 14464
rect 552 14432 584 14464
rect 624 14432 656 14464
rect 696 14432 728 14464
rect 768 14432 800 14464
rect 840 14432 872 14464
rect 912 14432 944 14464
rect 984 14432 1016 14464
rect 1056 14432 1088 14464
rect 1128 14432 1160 14464
rect 1200 14432 1232 14464
rect 1272 14432 1304 14464
rect 1344 14432 1376 14464
rect 1416 14432 1448 14464
rect 1488 14432 1520 14464
rect 1560 14432 1592 14464
rect 1632 14432 1664 14464
rect 1704 14432 1736 14464
rect 1776 14432 1808 14464
rect 1848 14432 1880 14464
rect 120 14360 152 14392
rect 192 14360 224 14392
rect 264 14360 296 14392
rect 336 14360 368 14392
rect 408 14360 440 14392
rect 480 14360 512 14392
rect 552 14360 584 14392
rect 624 14360 656 14392
rect 696 14360 728 14392
rect 768 14360 800 14392
rect 840 14360 872 14392
rect 912 14360 944 14392
rect 984 14360 1016 14392
rect 1056 14360 1088 14392
rect 1128 14360 1160 14392
rect 1200 14360 1232 14392
rect 1272 14360 1304 14392
rect 1344 14360 1376 14392
rect 1416 14360 1448 14392
rect 1488 14360 1520 14392
rect 1560 14360 1592 14392
rect 1632 14360 1664 14392
rect 1704 14360 1736 14392
rect 1776 14360 1808 14392
rect 1848 14360 1880 14392
rect 120 14288 152 14320
rect 192 14288 224 14320
rect 264 14288 296 14320
rect 336 14288 368 14320
rect 408 14288 440 14320
rect 480 14288 512 14320
rect 552 14288 584 14320
rect 624 14288 656 14320
rect 696 14288 728 14320
rect 768 14288 800 14320
rect 840 14288 872 14320
rect 912 14288 944 14320
rect 984 14288 1016 14320
rect 1056 14288 1088 14320
rect 1128 14288 1160 14320
rect 1200 14288 1232 14320
rect 1272 14288 1304 14320
rect 1344 14288 1376 14320
rect 1416 14288 1448 14320
rect 1488 14288 1520 14320
rect 1560 14288 1592 14320
rect 1632 14288 1664 14320
rect 1704 14288 1736 14320
rect 1776 14288 1808 14320
rect 1848 14288 1880 14320
rect 120 14216 152 14248
rect 192 14216 224 14248
rect 264 14216 296 14248
rect 336 14216 368 14248
rect 408 14216 440 14248
rect 480 14216 512 14248
rect 552 14216 584 14248
rect 624 14216 656 14248
rect 696 14216 728 14248
rect 768 14216 800 14248
rect 840 14216 872 14248
rect 912 14216 944 14248
rect 984 14216 1016 14248
rect 1056 14216 1088 14248
rect 1128 14216 1160 14248
rect 1200 14216 1232 14248
rect 1272 14216 1304 14248
rect 1344 14216 1376 14248
rect 1416 14216 1448 14248
rect 1488 14216 1520 14248
rect 1560 14216 1592 14248
rect 1632 14216 1664 14248
rect 1704 14216 1736 14248
rect 1776 14216 1808 14248
rect 1848 14216 1880 14248
rect 120 14144 152 14176
rect 192 14144 224 14176
rect 264 14144 296 14176
rect 336 14144 368 14176
rect 408 14144 440 14176
rect 480 14144 512 14176
rect 552 14144 584 14176
rect 624 14144 656 14176
rect 696 14144 728 14176
rect 768 14144 800 14176
rect 840 14144 872 14176
rect 912 14144 944 14176
rect 984 14144 1016 14176
rect 1056 14144 1088 14176
rect 1128 14144 1160 14176
rect 1200 14144 1232 14176
rect 1272 14144 1304 14176
rect 1344 14144 1376 14176
rect 1416 14144 1448 14176
rect 1488 14144 1520 14176
rect 1560 14144 1592 14176
rect 1632 14144 1664 14176
rect 1704 14144 1736 14176
rect 1776 14144 1808 14176
rect 1848 14144 1880 14176
rect 120 14072 152 14104
rect 192 14072 224 14104
rect 264 14072 296 14104
rect 336 14072 368 14104
rect 408 14072 440 14104
rect 480 14072 512 14104
rect 552 14072 584 14104
rect 624 14072 656 14104
rect 696 14072 728 14104
rect 768 14072 800 14104
rect 840 14072 872 14104
rect 912 14072 944 14104
rect 984 14072 1016 14104
rect 1056 14072 1088 14104
rect 1128 14072 1160 14104
rect 1200 14072 1232 14104
rect 1272 14072 1304 14104
rect 1344 14072 1376 14104
rect 1416 14072 1448 14104
rect 1488 14072 1520 14104
rect 1560 14072 1592 14104
rect 1632 14072 1664 14104
rect 1704 14072 1736 14104
rect 1776 14072 1808 14104
rect 1848 14072 1880 14104
rect 120 14000 152 14032
rect 192 14000 224 14032
rect 264 14000 296 14032
rect 336 14000 368 14032
rect 408 14000 440 14032
rect 480 14000 512 14032
rect 552 14000 584 14032
rect 624 14000 656 14032
rect 696 14000 728 14032
rect 768 14000 800 14032
rect 840 14000 872 14032
rect 912 14000 944 14032
rect 984 14000 1016 14032
rect 1056 14000 1088 14032
rect 1128 14000 1160 14032
rect 1200 14000 1232 14032
rect 1272 14000 1304 14032
rect 1344 14000 1376 14032
rect 1416 14000 1448 14032
rect 1488 14000 1520 14032
rect 1560 14000 1592 14032
rect 1632 14000 1664 14032
rect 1704 14000 1736 14032
rect 1776 14000 1808 14032
rect 1848 14000 1880 14032
rect 120 13928 152 13960
rect 192 13928 224 13960
rect 264 13928 296 13960
rect 336 13928 368 13960
rect 408 13928 440 13960
rect 480 13928 512 13960
rect 552 13928 584 13960
rect 624 13928 656 13960
rect 696 13928 728 13960
rect 768 13928 800 13960
rect 840 13928 872 13960
rect 912 13928 944 13960
rect 984 13928 1016 13960
rect 1056 13928 1088 13960
rect 1128 13928 1160 13960
rect 1200 13928 1232 13960
rect 1272 13928 1304 13960
rect 1344 13928 1376 13960
rect 1416 13928 1448 13960
rect 1488 13928 1520 13960
rect 1560 13928 1592 13960
rect 1632 13928 1664 13960
rect 1704 13928 1736 13960
rect 1776 13928 1808 13960
rect 1848 13928 1880 13960
rect 120 13856 152 13888
rect 192 13856 224 13888
rect 264 13856 296 13888
rect 336 13856 368 13888
rect 408 13856 440 13888
rect 480 13856 512 13888
rect 552 13856 584 13888
rect 624 13856 656 13888
rect 696 13856 728 13888
rect 768 13856 800 13888
rect 840 13856 872 13888
rect 912 13856 944 13888
rect 984 13856 1016 13888
rect 1056 13856 1088 13888
rect 1128 13856 1160 13888
rect 1200 13856 1232 13888
rect 1272 13856 1304 13888
rect 1344 13856 1376 13888
rect 1416 13856 1448 13888
rect 1488 13856 1520 13888
rect 1560 13856 1592 13888
rect 1632 13856 1664 13888
rect 1704 13856 1736 13888
rect 1776 13856 1808 13888
rect 1848 13856 1880 13888
rect 120 13784 152 13816
rect 192 13784 224 13816
rect 264 13784 296 13816
rect 336 13784 368 13816
rect 408 13784 440 13816
rect 480 13784 512 13816
rect 552 13784 584 13816
rect 624 13784 656 13816
rect 696 13784 728 13816
rect 768 13784 800 13816
rect 840 13784 872 13816
rect 912 13784 944 13816
rect 984 13784 1016 13816
rect 1056 13784 1088 13816
rect 1128 13784 1160 13816
rect 1200 13784 1232 13816
rect 1272 13784 1304 13816
rect 1344 13784 1376 13816
rect 1416 13784 1448 13816
rect 1488 13784 1520 13816
rect 1560 13784 1592 13816
rect 1632 13784 1664 13816
rect 1704 13784 1736 13816
rect 1776 13784 1808 13816
rect 1848 13784 1880 13816
rect 120 13712 152 13744
rect 192 13712 224 13744
rect 264 13712 296 13744
rect 336 13712 368 13744
rect 408 13712 440 13744
rect 480 13712 512 13744
rect 552 13712 584 13744
rect 624 13712 656 13744
rect 696 13712 728 13744
rect 768 13712 800 13744
rect 840 13712 872 13744
rect 912 13712 944 13744
rect 984 13712 1016 13744
rect 1056 13712 1088 13744
rect 1128 13712 1160 13744
rect 1200 13712 1232 13744
rect 1272 13712 1304 13744
rect 1344 13712 1376 13744
rect 1416 13712 1448 13744
rect 1488 13712 1520 13744
rect 1560 13712 1592 13744
rect 1632 13712 1664 13744
rect 1704 13712 1736 13744
rect 1776 13712 1808 13744
rect 1848 13712 1880 13744
rect 120 13640 152 13672
rect 192 13640 224 13672
rect 264 13640 296 13672
rect 336 13640 368 13672
rect 408 13640 440 13672
rect 480 13640 512 13672
rect 552 13640 584 13672
rect 624 13640 656 13672
rect 696 13640 728 13672
rect 768 13640 800 13672
rect 840 13640 872 13672
rect 912 13640 944 13672
rect 984 13640 1016 13672
rect 1056 13640 1088 13672
rect 1128 13640 1160 13672
rect 1200 13640 1232 13672
rect 1272 13640 1304 13672
rect 1344 13640 1376 13672
rect 1416 13640 1448 13672
rect 1488 13640 1520 13672
rect 1560 13640 1592 13672
rect 1632 13640 1664 13672
rect 1704 13640 1736 13672
rect 1776 13640 1808 13672
rect 1848 13640 1880 13672
rect 120 13568 152 13600
rect 192 13568 224 13600
rect 264 13568 296 13600
rect 336 13568 368 13600
rect 408 13568 440 13600
rect 480 13568 512 13600
rect 552 13568 584 13600
rect 624 13568 656 13600
rect 696 13568 728 13600
rect 768 13568 800 13600
rect 840 13568 872 13600
rect 912 13568 944 13600
rect 984 13568 1016 13600
rect 1056 13568 1088 13600
rect 1128 13568 1160 13600
rect 1200 13568 1232 13600
rect 1272 13568 1304 13600
rect 1344 13568 1376 13600
rect 1416 13568 1448 13600
rect 1488 13568 1520 13600
rect 1560 13568 1592 13600
rect 1632 13568 1664 13600
rect 1704 13568 1736 13600
rect 1776 13568 1808 13600
rect 1848 13568 1880 13600
rect 120 13496 152 13528
rect 192 13496 224 13528
rect 264 13496 296 13528
rect 336 13496 368 13528
rect 408 13496 440 13528
rect 480 13496 512 13528
rect 552 13496 584 13528
rect 624 13496 656 13528
rect 696 13496 728 13528
rect 768 13496 800 13528
rect 840 13496 872 13528
rect 912 13496 944 13528
rect 984 13496 1016 13528
rect 1056 13496 1088 13528
rect 1128 13496 1160 13528
rect 1200 13496 1232 13528
rect 1272 13496 1304 13528
rect 1344 13496 1376 13528
rect 1416 13496 1448 13528
rect 1488 13496 1520 13528
rect 1560 13496 1592 13528
rect 1632 13496 1664 13528
rect 1704 13496 1736 13528
rect 1776 13496 1808 13528
rect 1848 13496 1880 13528
rect 120 13424 152 13456
rect 192 13424 224 13456
rect 264 13424 296 13456
rect 336 13424 368 13456
rect 408 13424 440 13456
rect 480 13424 512 13456
rect 552 13424 584 13456
rect 624 13424 656 13456
rect 696 13424 728 13456
rect 768 13424 800 13456
rect 840 13424 872 13456
rect 912 13424 944 13456
rect 984 13424 1016 13456
rect 1056 13424 1088 13456
rect 1128 13424 1160 13456
rect 1200 13424 1232 13456
rect 1272 13424 1304 13456
rect 1344 13424 1376 13456
rect 1416 13424 1448 13456
rect 1488 13424 1520 13456
rect 1560 13424 1592 13456
rect 1632 13424 1664 13456
rect 1704 13424 1736 13456
rect 1776 13424 1808 13456
rect 1848 13424 1880 13456
rect 120 13352 152 13384
rect 192 13352 224 13384
rect 264 13352 296 13384
rect 336 13352 368 13384
rect 408 13352 440 13384
rect 480 13352 512 13384
rect 552 13352 584 13384
rect 624 13352 656 13384
rect 696 13352 728 13384
rect 768 13352 800 13384
rect 840 13352 872 13384
rect 912 13352 944 13384
rect 984 13352 1016 13384
rect 1056 13352 1088 13384
rect 1128 13352 1160 13384
rect 1200 13352 1232 13384
rect 1272 13352 1304 13384
rect 1344 13352 1376 13384
rect 1416 13352 1448 13384
rect 1488 13352 1520 13384
rect 1560 13352 1592 13384
rect 1632 13352 1664 13384
rect 1704 13352 1736 13384
rect 1776 13352 1808 13384
rect 1848 13352 1880 13384
rect 120 13280 152 13312
rect 192 13280 224 13312
rect 264 13280 296 13312
rect 336 13280 368 13312
rect 408 13280 440 13312
rect 480 13280 512 13312
rect 552 13280 584 13312
rect 624 13280 656 13312
rect 696 13280 728 13312
rect 768 13280 800 13312
rect 840 13280 872 13312
rect 912 13280 944 13312
rect 984 13280 1016 13312
rect 1056 13280 1088 13312
rect 1128 13280 1160 13312
rect 1200 13280 1232 13312
rect 1272 13280 1304 13312
rect 1344 13280 1376 13312
rect 1416 13280 1448 13312
rect 1488 13280 1520 13312
rect 1560 13280 1592 13312
rect 1632 13280 1664 13312
rect 1704 13280 1736 13312
rect 1776 13280 1808 13312
rect 1848 13280 1880 13312
rect 120 13208 152 13240
rect 192 13208 224 13240
rect 264 13208 296 13240
rect 336 13208 368 13240
rect 408 13208 440 13240
rect 480 13208 512 13240
rect 552 13208 584 13240
rect 624 13208 656 13240
rect 696 13208 728 13240
rect 768 13208 800 13240
rect 840 13208 872 13240
rect 912 13208 944 13240
rect 984 13208 1016 13240
rect 1056 13208 1088 13240
rect 1128 13208 1160 13240
rect 1200 13208 1232 13240
rect 1272 13208 1304 13240
rect 1344 13208 1376 13240
rect 1416 13208 1448 13240
rect 1488 13208 1520 13240
rect 1560 13208 1592 13240
rect 1632 13208 1664 13240
rect 1704 13208 1736 13240
rect 1776 13208 1808 13240
rect 1848 13208 1880 13240
rect 120 13136 152 13168
rect 192 13136 224 13168
rect 264 13136 296 13168
rect 336 13136 368 13168
rect 408 13136 440 13168
rect 480 13136 512 13168
rect 552 13136 584 13168
rect 624 13136 656 13168
rect 696 13136 728 13168
rect 768 13136 800 13168
rect 840 13136 872 13168
rect 912 13136 944 13168
rect 984 13136 1016 13168
rect 1056 13136 1088 13168
rect 1128 13136 1160 13168
rect 1200 13136 1232 13168
rect 1272 13136 1304 13168
rect 1344 13136 1376 13168
rect 1416 13136 1448 13168
rect 1488 13136 1520 13168
rect 1560 13136 1592 13168
rect 1632 13136 1664 13168
rect 1704 13136 1736 13168
rect 1776 13136 1808 13168
rect 1848 13136 1880 13168
rect 120 13064 152 13096
rect 192 13064 224 13096
rect 264 13064 296 13096
rect 336 13064 368 13096
rect 408 13064 440 13096
rect 480 13064 512 13096
rect 552 13064 584 13096
rect 624 13064 656 13096
rect 696 13064 728 13096
rect 768 13064 800 13096
rect 840 13064 872 13096
rect 912 13064 944 13096
rect 984 13064 1016 13096
rect 1056 13064 1088 13096
rect 1128 13064 1160 13096
rect 1200 13064 1232 13096
rect 1272 13064 1304 13096
rect 1344 13064 1376 13096
rect 1416 13064 1448 13096
rect 1488 13064 1520 13096
rect 1560 13064 1592 13096
rect 1632 13064 1664 13096
rect 1704 13064 1736 13096
rect 1776 13064 1808 13096
rect 1848 13064 1880 13096
rect 50 31416 1950 31430
rect 50 31384 699 31416
rect 731 31384 768 31416
rect 800 31384 838 31416
rect 870 31384 907 31416
rect 939 31384 978 31416
rect 1010 31384 1048 31416
rect 1080 31384 1116 31416
rect 1148 31384 1186 31416
rect 1218 31384 1950 31416
rect 50 31370 1950 31384
rect 50 27971 1950 28034
rect 50 27939 120 27971
rect 152 27939 192 27971
rect 224 27939 264 27971
rect 296 27939 336 27971
rect 368 27939 408 27971
rect 440 27939 480 27971
rect 512 27939 552 27971
rect 584 27939 624 27971
rect 656 27939 696 27971
rect 728 27939 768 27971
rect 800 27939 840 27971
rect 872 27939 912 27971
rect 944 27939 984 27971
rect 1016 27939 1056 27971
rect 1088 27939 1128 27971
rect 1160 27939 1200 27971
rect 1232 27939 1272 27971
rect 1304 27939 1344 27971
rect 1376 27939 1416 27971
rect 1448 27939 1488 27971
rect 1520 27939 1560 27971
rect 1592 27939 1632 27971
rect 1664 27939 1704 27971
rect 1736 27939 1776 27971
rect 1808 27939 1848 27971
rect 1880 27939 1950 27971
rect 50 27899 1950 27939
rect 50 27867 120 27899
rect 152 27867 192 27899
rect 224 27867 264 27899
rect 296 27867 336 27899
rect 368 27867 408 27899
rect 440 27867 480 27899
rect 512 27867 552 27899
rect 584 27867 624 27899
rect 656 27867 696 27899
rect 728 27867 768 27899
rect 800 27867 840 27899
rect 872 27867 912 27899
rect 944 27867 984 27899
rect 1016 27867 1056 27899
rect 1088 27867 1128 27899
rect 1160 27867 1200 27899
rect 1232 27867 1272 27899
rect 1304 27867 1344 27899
rect 1376 27867 1416 27899
rect 1448 27867 1488 27899
rect 1520 27867 1560 27899
rect 1592 27867 1632 27899
rect 1664 27867 1704 27899
rect 1736 27867 1776 27899
rect 1808 27867 1848 27899
rect 1880 27867 1950 27899
rect 50 27827 1950 27867
rect 50 27795 120 27827
rect 152 27795 192 27827
rect 224 27795 264 27827
rect 296 27795 336 27827
rect 368 27795 408 27827
rect 440 27795 480 27827
rect 512 27795 552 27827
rect 584 27795 624 27827
rect 656 27795 696 27827
rect 728 27795 768 27827
rect 800 27795 840 27827
rect 872 27795 912 27827
rect 944 27795 984 27827
rect 1016 27795 1056 27827
rect 1088 27795 1128 27827
rect 1160 27795 1200 27827
rect 1232 27795 1272 27827
rect 1304 27795 1344 27827
rect 1376 27795 1416 27827
rect 1448 27795 1488 27827
rect 1520 27795 1560 27827
rect 1592 27795 1632 27827
rect 1664 27795 1704 27827
rect 1736 27795 1776 27827
rect 1808 27795 1848 27827
rect 1880 27795 1950 27827
rect 50 27755 1950 27795
rect 50 27723 120 27755
rect 152 27723 192 27755
rect 224 27723 264 27755
rect 296 27723 336 27755
rect 368 27723 408 27755
rect 440 27723 480 27755
rect 512 27723 552 27755
rect 584 27723 624 27755
rect 656 27723 696 27755
rect 728 27723 768 27755
rect 800 27723 840 27755
rect 872 27723 912 27755
rect 944 27723 984 27755
rect 1016 27723 1056 27755
rect 1088 27723 1128 27755
rect 1160 27723 1200 27755
rect 1232 27723 1272 27755
rect 1304 27723 1344 27755
rect 1376 27723 1416 27755
rect 1448 27723 1488 27755
rect 1520 27723 1560 27755
rect 1592 27723 1632 27755
rect 1664 27723 1704 27755
rect 1736 27723 1776 27755
rect 1808 27723 1848 27755
rect 1880 27723 1950 27755
rect 50 27683 1950 27723
rect 50 27651 120 27683
rect 152 27651 192 27683
rect 224 27651 264 27683
rect 296 27651 336 27683
rect 368 27651 408 27683
rect 440 27651 480 27683
rect 512 27651 552 27683
rect 584 27651 624 27683
rect 656 27651 696 27683
rect 728 27651 768 27683
rect 800 27651 840 27683
rect 872 27651 912 27683
rect 944 27651 984 27683
rect 1016 27651 1056 27683
rect 1088 27651 1128 27683
rect 1160 27651 1200 27683
rect 1232 27651 1272 27683
rect 1304 27651 1344 27683
rect 1376 27651 1416 27683
rect 1448 27651 1488 27683
rect 1520 27651 1560 27683
rect 1592 27651 1632 27683
rect 1664 27651 1704 27683
rect 1736 27651 1776 27683
rect 1808 27651 1848 27683
rect 1880 27651 1950 27683
rect 50 27611 1950 27651
rect 50 27579 120 27611
rect 152 27579 192 27611
rect 224 27579 264 27611
rect 296 27579 336 27611
rect 368 27579 408 27611
rect 440 27579 480 27611
rect 512 27579 552 27611
rect 584 27579 624 27611
rect 656 27579 696 27611
rect 728 27579 768 27611
rect 800 27579 840 27611
rect 872 27579 912 27611
rect 944 27579 984 27611
rect 1016 27579 1056 27611
rect 1088 27579 1128 27611
rect 1160 27579 1200 27611
rect 1232 27579 1272 27611
rect 1304 27579 1344 27611
rect 1376 27579 1416 27611
rect 1448 27579 1488 27611
rect 1520 27579 1560 27611
rect 1592 27579 1632 27611
rect 1664 27579 1704 27611
rect 1736 27579 1776 27611
rect 1808 27579 1848 27611
rect 1880 27579 1950 27611
rect 50 27539 1950 27579
rect 50 27507 120 27539
rect 152 27507 192 27539
rect 224 27507 264 27539
rect 296 27507 336 27539
rect 368 27507 408 27539
rect 440 27507 480 27539
rect 512 27507 552 27539
rect 584 27507 624 27539
rect 656 27507 696 27539
rect 728 27507 768 27539
rect 800 27507 840 27539
rect 872 27507 912 27539
rect 944 27507 984 27539
rect 1016 27507 1056 27539
rect 1088 27507 1128 27539
rect 1160 27507 1200 27539
rect 1232 27507 1272 27539
rect 1304 27507 1344 27539
rect 1376 27507 1416 27539
rect 1448 27507 1488 27539
rect 1520 27507 1560 27539
rect 1592 27507 1632 27539
rect 1664 27507 1704 27539
rect 1736 27507 1776 27539
rect 1808 27507 1848 27539
rect 1880 27507 1950 27539
rect 50 27467 1950 27507
rect 50 27435 120 27467
rect 152 27435 192 27467
rect 224 27435 264 27467
rect 296 27435 336 27467
rect 368 27435 408 27467
rect 440 27435 480 27467
rect 512 27435 552 27467
rect 584 27435 624 27467
rect 656 27435 696 27467
rect 728 27435 768 27467
rect 800 27435 840 27467
rect 872 27435 912 27467
rect 944 27435 984 27467
rect 1016 27435 1056 27467
rect 1088 27435 1128 27467
rect 1160 27435 1200 27467
rect 1232 27435 1272 27467
rect 1304 27435 1344 27467
rect 1376 27435 1416 27467
rect 1448 27435 1488 27467
rect 1520 27435 1560 27467
rect 1592 27435 1632 27467
rect 1664 27435 1704 27467
rect 1736 27435 1776 27467
rect 1808 27435 1848 27467
rect 1880 27435 1950 27467
rect 50 27395 1950 27435
rect 50 27363 120 27395
rect 152 27363 192 27395
rect 224 27363 264 27395
rect 296 27363 336 27395
rect 368 27363 408 27395
rect 440 27363 480 27395
rect 512 27363 552 27395
rect 584 27363 624 27395
rect 656 27363 696 27395
rect 728 27363 768 27395
rect 800 27363 840 27395
rect 872 27363 912 27395
rect 944 27363 984 27395
rect 1016 27363 1056 27395
rect 1088 27363 1128 27395
rect 1160 27363 1200 27395
rect 1232 27363 1272 27395
rect 1304 27363 1344 27395
rect 1376 27363 1416 27395
rect 1448 27363 1488 27395
rect 1520 27363 1560 27395
rect 1592 27363 1632 27395
rect 1664 27363 1704 27395
rect 1736 27363 1776 27395
rect 1808 27363 1848 27395
rect 1880 27363 1950 27395
rect 50 27323 1950 27363
rect 50 27291 120 27323
rect 152 27291 192 27323
rect 224 27291 264 27323
rect 296 27291 336 27323
rect 368 27291 408 27323
rect 440 27291 480 27323
rect 512 27291 552 27323
rect 584 27291 624 27323
rect 656 27291 696 27323
rect 728 27291 768 27323
rect 800 27291 840 27323
rect 872 27291 912 27323
rect 944 27291 984 27323
rect 1016 27291 1056 27323
rect 1088 27291 1128 27323
rect 1160 27291 1200 27323
rect 1232 27291 1272 27323
rect 1304 27291 1344 27323
rect 1376 27291 1416 27323
rect 1448 27291 1488 27323
rect 1520 27291 1560 27323
rect 1592 27291 1632 27323
rect 1664 27291 1704 27323
rect 1736 27291 1776 27323
rect 1808 27291 1848 27323
rect 1880 27291 1950 27323
rect 50 27251 1950 27291
rect 50 27219 120 27251
rect 152 27219 192 27251
rect 224 27219 264 27251
rect 296 27219 336 27251
rect 368 27219 408 27251
rect 440 27219 480 27251
rect 512 27219 552 27251
rect 584 27219 624 27251
rect 656 27219 696 27251
rect 728 27219 768 27251
rect 800 27219 840 27251
rect 872 27219 912 27251
rect 944 27219 984 27251
rect 1016 27219 1056 27251
rect 1088 27219 1128 27251
rect 1160 27219 1200 27251
rect 1232 27219 1272 27251
rect 1304 27219 1344 27251
rect 1376 27219 1416 27251
rect 1448 27219 1488 27251
rect 1520 27219 1560 27251
rect 1592 27219 1632 27251
rect 1664 27219 1704 27251
rect 1736 27219 1776 27251
rect 1808 27219 1848 27251
rect 1880 27219 1950 27251
rect 50 27179 1950 27219
rect 50 27147 120 27179
rect 152 27147 192 27179
rect 224 27147 264 27179
rect 296 27147 336 27179
rect 368 27147 408 27179
rect 440 27147 480 27179
rect 512 27147 552 27179
rect 584 27147 624 27179
rect 656 27147 696 27179
rect 728 27147 768 27179
rect 800 27147 840 27179
rect 872 27147 912 27179
rect 944 27147 984 27179
rect 1016 27147 1056 27179
rect 1088 27147 1128 27179
rect 1160 27147 1200 27179
rect 1232 27147 1272 27179
rect 1304 27147 1344 27179
rect 1376 27147 1416 27179
rect 1448 27147 1488 27179
rect 1520 27147 1560 27179
rect 1592 27147 1632 27179
rect 1664 27147 1704 27179
rect 1736 27147 1776 27179
rect 1808 27147 1848 27179
rect 1880 27147 1950 27179
rect 50 27107 1950 27147
rect 50 27075 120 27107
rect 152 27075 192 27107
rect 224 27075 264 27107
rect 296 27075 336 27107
rect 368 27075 408 27107
rect 440 27075 480 27107
rect 512 27075 552 27107
rect 584 27075 624 27107
rect 656 27075 696 27107
rect 728 27075 768 27107
rect 800 27075 840 27107
rect 872 27075 912 27107
rect 944 27075 984 27107
rect 1016 27075 1056 27107
rect 1088 27075 1128 27107
rect 1160 27075 1200 27107
rect 1232 27075 1272 27107
rect 1304 27075 1344 27107
rect 1376 27075 1416 27107
rect 1448 27075 1488 27107
rect 1520 27075 1560 27107
rect 1592 27075 1632 27107
rect 1664 27075 1704 27107
rect 1736 27075 1776 27107
rect 1808 27075 1848 27107
rect 1880 27075 1950 27107
rect 50 27035 1950 27075
rect 50 27003 120 27035
rect 152 27003 192 27035
rect 224 27003 264 27035
rect 296 27003 336 27035
rect 368 27003 408 27035
rect 440 27003 480 27035
rect 512 27003 552 27035
rect 584 27003 624 27035
rect 656 27003 696 27035
rect 728 27003 768 27035
rect 800 27003 840 27035
rect 872 27003 912 27035
rect 944 27003 984 27035
rect 1016 27003 1056 27035
rect 1088 27003 1128 27035
rect 1160 27003 1200 27035
rect 1232 27003 1272 27035
rect 1304 27003 1344 27035
rect 1376 27003 1416 27035
rect 1448 27003 1488 27035
rect 1520 27003 1560 27035
rect 1592 27003 1632 27035
rect 1664 27003 1704 27035
rect 1736 27003 1776 27035
rect 1808 27003 1848 27035
rect 1880 27003 1950 27035
rect 50 26963 1950 27003
rect 50 26931 120 26963
rect 152 26931 192 26963
rect 224 26931 264 26963
rect 296 26931 336 26963
rect 368 26931 408 26963
rect 440 26931 480 26963
rect 512 26931 552 26963
rect 584 26931 624 26963
rect 656 26931 696 26963
rect 728 26931 768 26963
rect 800 26931 840 26963
rect 872 26931 912 26963
rect 944 26931 984 26963
rect 1016 26931 1056 26963
rect 1088 26931 1128 26963
rect 1160 26931 1200 26963
rect 1232 26931 1272 26963
rect 1304 26931 1344 26963
rect 1376 26931 1416 26963
rect 1448 26931 1488 26963
rect 1520 26931 1560 26963
rect 1592 26931 1632 26963
rect 1664 26931 1704 26963
rect 1736 26931 1776 26963
rect 1808 26931 1848 26963
rect 1880 26931 1950 26963
rect 50 26891 1950 26931
rect 50 26859 120 26891
rect 152 26859 192 26891
rect 224 26859 264 26891
rect 296 26859 336 26891
rect 368 26859 408 26891
rect 440 26859 480 26891
rect 512 26859 552 26891
rect 584 26859 624 26891
rect 656 26859 696 26891
rect 728 26859 768 26891
rect 800 26859 840 26891
rect 872 26859 912 26891
rect 944 26859 984 26891
rect 1016 26859 1056 26891
rect 1088 26859 1128 26891
rect 1160 26859 1200 26891
rect 1232 26859 1272 26891
rect 1304 26859 1344 26891
rect 1376 26859 1416 26891
rect 1448 26859 1488 26891
rect 1520 26859 1560 26891
rect 1592 26859 1632 26891
rect 1664 26859 1704 26891
rect 1736 26859 1776 26891
rect 1808 26859 1848 26891
rect 1880 26859 1950 26891
rect 50 26819 1950 26859
rect 50 26787 120 26819
rect 152 26787 192 26819
rect 224 26787 264 26819
rect 296 26787 336 26819
rect 368 26787 408 26819
rect 440 26787 480 26819
rect 512 26787 552 26819
rect 584 26787 624 26819
rect 656 26787 696 26819
rect 728 26787 768 26819
rect 800 26787 840 26819
rect 872 26787 912 26819
rect 944 26787 984 26819
rect 1016 26787 1056 26819
rect 1088 26787 1128 26819
rect 1160 26787 1200 26819
rect 1232 26787 1272 26819
rect 1304 26787 1344 26819
rect 1376 26787 1416 26819
rect 1448 26787 1488 26819
rect 1520 26787 1560 26819
rect 1592 26787 1632 26819
rect 1664 26787 1704 26819
rect 1736 26787 1776 26819
rect 1808 26787 1848 26819
rect 1880 26787 1950 26819
rect 50 26747 1950 26787
rect 50 26715 120 26747
rect 152 26715 192 26747
rect 224 26715 264 26747
rect 296 26715 336 26747
rect 368 26715 408 26747
rect 440 26715 480 26747
rect 512 26715 552 26747
rect 584 26715 624 26747
rect 656 26715 696 26747
rect 728 26715 768 26747
rect 800 26715 840 26747
rect 872 26715 912 26747
rect 944 26715 984 26747
rect 1016 26715 1056 26747
rect 1088 26715 1128 26747
rect 1160 26715 1200 26747
rect 1232 26715 1272 26747
rect 1304 26715 1344 26747
rect 1376 26715 1416 26747
rect 1448 26715 1488 26747
rect 1520 26715 1560 26747
rect 1592 26715 1632 26747
rect 1664 26715 1704 26747
rect 1736 26715 1776 26747
rect 1808 26715 1848 26747
rect 1880 26715 1950 26747
rect 50 26675 1950 26715
rect 50 26643 120 26675
rect 152 26643 192 26675
rect 224 26643 264 26675
rect 296 26643 336 26675
rect 368 26643 408 26675
rect 440 26643 480 26675
rect 512 26643 552 26675
rect 584 26643 624 26675
rect 656 26643 696 26675
rect 728 26643 768 26675
rect 800 26643 840 26675
rect 872 26643 912 26675
rect 944 26643 984 26675
rect 1016 26643 1056 26675
rect 1088 26643 1128 26675
rect 1160 26643 1200 26675
rect 1232 26643 1272 26675
rect 1304 26643 1344 26675
rect 1376 26643 1416 26675
rect 1448 26643 1488 26675
rect 1520 26643 1560 26675
rect 1592 26643 1632 26675
rect 1664 26643 1704 26675
rect 1736 26643 1776 26675
rect 1808 26643 1848 26675
rect 1880 26643 1950 26675
rect 50 26603 1950 26643
rect 50 26571 120 26603
rect 152 26571 192 26603
rect 224 26571 264 26603
rect 296 26571 336 26603
rect 368 26571 408 26603
rect 440 26571 480 26603
rect 512 26571 552 26603
rect 584 26571 624 26603
rect 656 26571 696 26603
rect 728 26571 768 26603
rect 800 26571 840 26603
rect 872 26571 912 26603
rect 944 26571 984 26603
rect 1016 26571 1056 26603
rect 1088 26571 1128 26603
rect 1160 26571 1200 26603
rect 1232 26571 1272 26603
rect 1304 26571 1344 26603
rect 1376 26571 1416 26603
rect 1448 26571 1488 26603
rect 1520 26571 1560 26603
rect 1592 26571 1632 26603
rect 1664 26571 1704 26603
rect 1736 26571 1776 26603
rect 1808 26571 1848 26603
rect 1880 26571 1950 26603
rect 50 26531 1950 26571
rect 50 26499 120 26531
rect 152 26499 192 26531
rect 224 26499 264 26531
rect 296 26499 336 26531
rect 368 26499 408 26531
rect 440 26499 480 26531
rect 512 26499 552 26531
rect 584 26499 624 26531
rect 656 26499 696 26531
rect 728 26499 768 26531
rect 800 26499 840 26531
rect 872 26499 912 26531
rect 944 26499 984 26531
rect 1016 26499 1056 26531
rect 1088 26499 1128 26531
rect 1160 26499 1200 26531
rect 1232 26499 1272 26531
rect 1304 26499 1344 26531
rect 1376 26499 1416 26531
rect 1448 26499 1488 26531
rect 1520 26499 1560 26531
rect 1592 26499 1632 26531
rect 1664 26499 1704 26531
rect 1736 26499 1776 26531
rect 1808 26499 1848 26531
rect 1880 26499 1950 26531
rect 50 26459 1950 26499
rect 50 26427 120 26459
rect 152 26427 192 26459
rect 224 26427 264 26459
rect 296 26427 336 26459
rect 368 26427 408 26459
rect 440 26427 480 26459
rect 512 26427 552 26459
rect 584 26427 624 26459
rect 656 26427 696 26459
rect 728 26427 768 26459
rect 800 26427 840 26459
rect 872 26427 912 26459
rect 944 26427 984 26459
rect 1016 26427 1056 26459
rect 1088 26427 1128 26459
rect 1160 26427 1200 26459
rect 1232 26427 1272 26459
rect 1304 26427 1344 26459
rect 1376 26427 1416 26459
rect 1448 26427 1488 26459
rect 1520 26427 1560 26459
rect 1592 26427 1632 26459
rect 1664 26427 1704 26459
rect 1736 26427 1776 26459
rect 1808 26427 1848 26459
rect 1880 26427 1950 26459
rect 50 26387 1950 26427
rect 50 26355 120 26387
rect 152 26355 192 26387
rect 224 26355 264 26387
rect 296 26355 336 26387
rect 368 26355 408 26387
rect 440 26355 480 26387
rect 512 26355 552 26387
rect 584 26355 624 26387
rect 656 26355 696 26387
rect 728 26355 768 26387
rect 800 26355 840 26387
rect 872 26355 912 26387
rect 944 26355 984 26387
rect 1016 26355 1056 26387
rect 1088 26355 1128 26387
rect 1160 26355 1200 26387
rect 1232 26355 1272 26387
rect 1304 26355 1344 26387
rect 1376 26355 1416 26387
rect 1448 26355 1488 26387
rect 1520 26355 1560 26387
rect 1592 26355 1632 26387
rect 1664 26355 1704 26387
rect 1736 26355 1776 26387
rect 1808 26355 1848 26387
rect 1880 26355 1950 26387
rect 50 26315 1950 26355
rect 50 26283 120 26315
rect 152 26283 192 26315
rect 224 26283 264 26315
rect 296 26283 336 26315
rect 368 26283 408 26315
rect 440 26283 480 26315
rect 512 26283 552 26315
rect 584 26283 624 26315
rect 656 26283 696 26315
rect 728 26283 768 26315
rect 800 26283 840 26315
rect 872 26283 912 26315
rect 944 26283 984 26315
rect 1016 26283 1056 26315
rect 1088 26283 1128 26315
rect 1160 26283 1200 26315
rect 1232 26283 1272 26315
rect 1304 26283 1344 26315
rect 1376 26283 1416 26315
rect 1448 26283 1488 26315
rect 1520 26283 1560 26315
rect 1592 26283 1632 26315
rect 1664 26283 1704 26315
rect 1736 26283 1776 26315
rect 1808 26283 1848 26315
rect 1880 26283 1950 26315
rect 50 26243 1950 26283
rect 50 26211 120 26243
rect 152 26211 192 26243
rect 224 26211 264 26243
rect 296 26211 336 26243
rect 368 26211 408 26243
rect 440 26211 480 26243
rect 512 26211 552 26243
rect 584 26211 624 26243
rect 656 26211 696 26243
rect 728 26211 768 26243
rect 800 26211 840 26243
rect 872 26211 912 26243
rect 944 26211 984 26243
rect 1016 26211 1056 26243
rect 1088 26211 1128 26243
rect 1160 26211 1200 26243
rect 1232 26211 1272 26243
rect 1304 26211 1344 26243
rect 1376 26211 1416 26243
rect 1448 26211 1488 26243
rect 1520 26211 1560 26243
rect 1592 26211 1632 26243
rect 1664 26211 1704 26243
rect 1736 26211 1776 26243
rect 1808 26211 1848 26243
rect 1880 26211 1950 26243
rect 50 26171 1950 26211
rect 50 26139 120 26171
rect 152 26139 192 26171
rect 224 26139 264 26171
rect 296 26139 336 26171
rect 368 26139 408 26171
rect 440 26139 480 26171
rect 512 26139 552 26171
rect 584 26139 624 26171
rect 656 26139 696 26171
rect 728 26139 768 26171
rect 800 26139 840 26171
rect 872 26139 912 26171
rect 944 26139 984 26171
rect 1016 26139 1056 26171
rect 1088 26139 1128 26171
rect 1160 26139 1200 26171
rect 1232 26139 1272 26171
rect 1304 26139 1344 26171
rect 1376 26139 1416 26171
rect 1448 26139 1488 26171
rect 1520 26139 1560 26171
rect 1592 26139 1632 26171
rect 1664 26139 1704 26171
rect 1736 26139 1776 26171
rect 1808 26139 1848 26171
rect 1880 26139 1950 26171
rect 50 26099 1950 26139
rect 50 26067 120 26099
rect 152 26067 192 26099
rect 224 26067 264 26099
rect 296 26067 336 26099
rect 368 26067 408 26099
rect 440 26067 480 26099
rect 512 26067 552 26099
rect 584 26067 624 26099
rect 656 26067 696 26099
rect 728 26067 768 26099
rect 800 26067 840 26099
rect 872 26067 912 26099
rect 944 26067 984 26099
rect 1016 26067 1056 26099
rect 1088 26067 1128 26099
rect 1160 26067 1200 26099
rect 1232 26067 1272 26099
rect 1304 26067 1344 26099
rect 1376 26067 1416 26099
rect 1448 26067 1488 26099
rect 1520 26067 1560 26099
rect 1592 26067 1632 26099
rect 1664 26067 1704 26099
rect 1736 26067 1776 26099
rect 1808 26067 1848 26099
rect 1880 26067 1950 26099
rect 50 26027 1950 26067
rect 50 25995 120 26027
rect 152 25995 192 26027
rect 224 25995 264 26027
rect 296 25995 336 26027
rect 368 25995 408 26027
rect 440 25995 480 26027
rect 512 25995 552 26027
rect 584 25995 624 26027
rect 656 25995 696 26027
rect 728 25995 768 26027
rect 800 25995 840 26027
rect 872 25995 912 26027
rect 944 25995 984 26027
rect 1016 25995 1056 26027
rect 1088 25995 1128 26027
rect 1160 25995 1200 26027
rect 1232 25995 1272 26027
rect 1304 25995 1344 26027
rect 1376 25995 1416 26027
rect 1448 25995 1488 26027
rect 1520 25995 1560 26027
rect 1592 25995 1632 26027
rect 1664 25995 1704 26027
rect 1736 25995 1776 26027
rect 1808 25995 1848 26027
rect 1880 25995 1950 26027
rect 50 25955 1950 25995
rect 50 25923 120 25955
rect 152 25923 192 25955
rect 224 25923 264 25955
rect 296 25923 336 25955
rect 368 25923 408 25955
rect 440 25923 480 25955
rect 512 25923 552 25955
rect 584 25923 624 25955
rect 656 25923 696 25955
rect 728 25923 768 25955
rect 800 25923 840 25955
rect 872 25923 912 25955
rect 944 25923 984 25955
rect 1016 25923 1056 25955
rect 1088 25923 1128 25955
rect 1160 25923 1200 25955
rect 1232 25923 1272 25955
rect 1304 25923 1344 25955
rect 1376 25923 1416 25955
rect 1448 25923 1488 25955
rect 1520 25923 1560 25955
rect 1592 25923 1632 25955
rect 1664 25923 1704 25955
rect 1736 25923 1776 25955
rect 1808 25923 1848 25955
rect 1880 25923 1950 25955
rect 50 25883 1950 25923
rect 50 25851 120 25883
rect 152 25851 192 25883
rect 224 25851 264 25883
rect 296 25851 336 25883
rect 368 25851 408 25883
rect 440 25851 480 25883
rect 512 25851 552 25883
rect 584 25851 624 25883
rect 656 25851 696 25883
rect 728 25851 768 25883
rect 800 25851 840 25883
rect 872 25851 912 25883
rect 944 25851 984 25883
rect 1016 25851 1056 25883
rect 1088 25851 1128 25883
rect 1160 25851 1200 25883
rect 1232 25851 1272 25883
rect 1304 25851 1344 25883
rect 1376 25851 1416 25883
rect 1448 25851 1488 25883
rect 1520 25851 1560 25883
rect 1592 25851 1632 25883
rect 1664 25851 1704 25883
rect 1736 25851 1776 25883
rect 1808 25851 1848 25883
rect 1880 25851 1950 25883
rect 50 25811 1950 25851
rect 50 25779 120 25811
rect 152 25779 192 25811
rect 224 25779 264 25811
rect 296 25779 336 25811
rect 368 25779 408 25811
rect 440 25779 480 25811
rect 512 25779 552 25811
rect 584 25779 624 25811
rect 656 25779 696 25811
rect 728 25779 768 25811
rect 800 25779 840 25811
rect 872 25779 912 25811
rect 944 25779 984 25811
rect 1016 25779 1056 25811
rect 1088 25779 1128 25811
rect 1160 25779 1200 25811
rect 1232 25779 1272 25811
rect 1304 25779 1344 25811
rect 1376 25779 1416 25811
rect 1448 25779 1488 25811
rect 1520 25779 1560 25811
rect 1592 25779 1632 25811
rect 1664 25779 1704 25811
rect 1736 25779 1776 25811
rect 1808 25779 1848 25811
rect 1880 25779 1950 25811
rect 50 25739 1950 25779
rect 50 25707 120 25739
rect 152 25707 192 25739
rect 224 25707 264 25739
rect 296 25707 336 25739
rect 368 25707 408 25739
rect 440 25707 480 25739
rect 512 25707 552 25739
rect 584 25707 624 25739
rect 656 25707 696 25739
rect 728 25707 768 25739
rect 800 25707 840 25739
rect 872 25707 912 25739
rect 944 25707 984 25739
rect 1016 25707 1056 25739
rect 1088 25707 1128 25739
rect 1160 25707 1200 25739
rect 1232 25707 1272 25739
rect 1304 25707 1344 25739
rect 1376 25707 1416 25739
rect 1448 25707 1488 25739
rect 1520 25707 1560 25739
rect 1592 25707 1632 25739
rect 1664 25707 1704 25739
rect 1736 25707 1776 25739
rect 1808 25707 1848 25739
rect 1880 25707 1950 25739
rect 50 25667 1950 25707
rect 50 25635 120 25667
rect 152 25635 192 25667
rect 224 25635 264 25667
rect 296 25635 336 25667
rect 368 25635 408 25667
rect 440 25635 480 25667
rect 512 25635 552 25667
rect 584 25635 624 25667
rect 656 25635 696 25667
rect 728 25635 768 25667
rect 800 25635 840 25667
rect 872 25635 912 25667
rect 944 25635 984 25667
rect 1016 25635 1056 25667
rect 1088 25635 1128 25667
rect 1160 25635 1200 25667
rect 1232 25635 1272 25667
rect 1304 25635 1344 25667
rect 1376 25635 1416 25667
rect 1448 25635 1488 25667
rect 1520 25635 1560 25667
rect 1592 25635 1632 25667
rect 1664 25635 1704 25667
rect 1736 25635 1776 25667
rect 1808 25635 1848 25667
rect 1880 25635 1950 25667
rect 50 25595 1950 25635
rect 50 25563 120 25595
rect 152 25563 192 25595
rect 224 25563 264 25595
rect 296 25563 336 25595
rect 368 25563 408 25595
rect 440 25563 480 25595
rect 512 25563 552 25595
rect 584 25563 624 25595
rect 656 25563 696 25595
rect 728 25563 768 25595
rect 800 25563 840 25595
rect 872 25563 912 25595
rect 944 25563 984 25595
rect 1016 25563 1056 25595
rect 1088 25563 1128 25595
rect 1160 25563 1200 25595
rect 1232 25563 1272 25595
rect 1304 25563 1344 25595
rect 1376 25563 1416 25595
rect 1448 25563 1488 25595
rect 1520 25563 1560 25595
rect 1592 25563 1632 25595
rect 1664 25563 1704 25595
rect 1736 25563 1776 25595
rect 1808 25563 1848 25595
rect 1880 25563 1950 25595
rect 50 25523 1950 25563
rect 50 25491 120 25523
rect 152 25491 192 25523
rect 224 25491 264 25523
rect 296 25491 336 25523
rect 368 25491 408 25523
rect 440 25491 480 25523
rect 512 25491 552 25523
rect 584 25491 624 25523
rect 656 25491 696 25523
rect 728 25491 768 25523
rect 800 25491 840 25523
rect 872 25491 912 25523
rect 944 25491 984 25523
rect 1016 25491 1056 25523
rect 1088 25491 1128 25523
rect 1160 25491 1200 25523
rect 1232 25491 1272 25523
rect 1304 25491 1344 25523
rect 1376 25491 1416 25523
rect 1448 25491 1488 25523
rect 1520 25491 1560 25523
rect 1592 25491 1632 25523
rect 1664 25491 1704 25523
rect 1736 25491 1776 25523
rect 1808 25491 1848 25523
rect 1880 25491 1950 25523
rect 50 25451 1950 25491
rect 50 25419 120 25451
rect 152 25419 192 25451
rect 224 25419 264 25451
rect 296 25419 336 25451
rect 368 25419 408 25451
rect 440 25419 480 25451
rect 512 25419 552 25451
rect 584 25419 624 25451
rect 656 25419 696 25451
rect 728 25419 768 25451
rect 800 25419 840 25451
rect 872 25419 912 25451
rect 944 25419 984 25451
rect 1016 25419 1056 25451
rect 1088 25419 1128 25451
rect 1160 25419 1200 25451
rect 1232 25419 1272 25451
rect 1304 25419 1344 25451
rect 1376 25419 1416 25451
rect 1448 25419 1488 25451
rect 1520 25419 1560 25451
rect 1592 25419 1632 25451
rect 1664 25419 1704 25451
rect 1736 25419 1776 25451
rect 1808 25419 1848 25451
rect 1880 25419 1950 25451
rect 50 25379 1950 25419
rect 50 25347 120 25379
rect 152 25347 192 25379
rect 224 25347 264 25379
rect 296 25347 336 25379
rect 368 25347 408 25379
rect 440 25347 480 25379
rect 512 25347 552 25379
rect 584 25347 624 25379
rect 656 25347 696 25379
rect 728 25347 768 25379
rect 800 25347 840 25379
rect 872 25347 912 25379
rect 944 25347 984 25379
rect 1016 25347 1056 25379
rect 1088 25347 1128 25379
rect 1160 25347 1200 25379
rect 1232 25347 1272 25379
rect 1304 25347 1344 25379
rect 1376 25347 1416 25379
rect 1448 25347 1488 25379
rect 1520 25347 1560 25379
rect 1592 25347 1632 25379
rect 1664 25347 1704 25379
rect 1736 25347 1776 25379
rect 1808 25347 1848 25379
rect 1880 25347 1950 25379
rect 50 25307 1950 25347
rect 50 25275 120 25307
rect 152 25275 192 25307
rect 224 25275 264 25307
rect 296 25275 336 25307
rect 368 25275 408 25307
rect 440 25275 480 25307
rect 512 25275 552 25307
rect 584 25275 624 25307
rect 656 25275 696 25307
rect 728 25275 768 25307
rect 800 25275 840 25307
rect 872 25275 912 25307
rect 944 25275 984 25307
rect 1016 25275 1056 25307
rect 1088 25275 1128 25307
rect 1160 25275 1200 25307
rect 1232 25275 1272 25307
rect 1304 25275 1344 25307
rect 1376 25275 1416 25307
rect 1448 25275 1488 25307
rect 1520 25275 1560 25307
rect 1592 25275 1632 25307
rect 1664 25275 1704 25307
rect 1736 25275 1776 25307
rect 1808 25275 1848 25307
rect 1880 25275 1950 25307
rect 50 25235 1950 25275
rect 50 25203 120 25235
rect 152 25203 192 25235
rect 224 25203 264 25235
rect 296 25203 336 25235
rect 368 25203 408 25235
rect 440 25203 480 25235
rect 512 25203 552 25235
rect 584 25203 624 25235
rect 656 25203 696 25235
rect 728 25203 768 25235
rect 800 25203 840 25235
rect 872 25203 912 25235
rect 944 25203 984 25235
rect 1016 25203 1056 25235
rect 1088 25203 1128 25235
rect 1160 25203 1200 25235
rect 1232 25203 1272 25235
rect 1304 25203 1344 25235
rect 1376 25203 1416 25235
rect 1448 25203 1488 25235
rect 1520 25203 1560 25235
rect 1592 25203 1632 25235
rect 1664 25203 1704 25235
rect 1736 25203 1776 25235
rect 1808 25203 1848 25235
rect 1880 25203 1950 25235
rect 50 25163 1950 25203
rect 50 25131 120 25163
rect 152 25131 192 25163
rect 224 25131 264 25163
rect 296 25131 336 25163
rect 368 25131 408 25163
rect 440 25131 480 25163
rect 512 25131 552 25163
rect 584 25131 624 25163
rect 656 25131 696 25163
rect 728 25131 768 25163
rect 800 25131 840 25163
rect 872 25131 912 25163
rect 944 25131 984 25163
rect 1016 25131 1056 25163
rect 1088 25131 1128 25163
rect 1160 25131 1200 25163
rect 1232 25131 1272 25163
rect 1304 25131 1344 25163
rect 1376 25131 1416 25163
rect 1448 25131 1488 25163
rect 1520 25131 1560 25163
rect 1592 25131 1632 25163
rect 1664 25131 1704 25163
rect 1736 25131 1776 25163
rect 1808 25131 1848 25163
rect 1880 25131 1950 25163
rect 50 25091 1950 25131
rect 50 25059 120 25091
rect 152 25059 192 25091
rect 224 25059 264 25091
rect 296 25059 336 25091
rect 368 25059 408 25091
rect 440 25059 480 25091
rect 512 25059 552 25091
rect 584 25059 624 25091
rect 656 25059 696 25091
rect 728 25059 768 25091
rect 800 25059 840 25091
rect 872 25059 912 25091
rect 944 25059 984 25091
rect 1016 25059 1056 25091
rect 1088 25059 1128 25091
rect 1160 25059 1200 25091
rect 1232 25059 1272 25091
rect 1304 25059 1344 25091
rect 1376 25059 1416 25091
rect 1448 25059 1488 25091
rect 1520 25059 1560 25091
rect 1592 25059 1632 25091
rect 1664 25059 1704 25091
rect 1736 25059 1776 25091
rect 1808 25059 1848 25091
rect 1880 25059 1950 25091
rect 50 25019 1950 25059
rect 50 24987 120 25019
rect 152 24987 192 25019
rect 224 24987 264 25019
rect 296 24987 336 25019
rect 368 24987 408 25019
rect 440 24987 480 25019
rect 512 24987 552 25019
rect 584 24987 624 25019
rect 656 24987 696 25019
rect 728 24987 768 25019
rect 800 24987 840 25019
rect 872 24987 912 25019
rect 944 24987 984 25019
rect 1016 24987 1056 25019
rect 1088 24987 1128 25019
rect 1160 24987 1200 25019
rect 1232 24987 1272 25019
rect 1304 24987 1344 25019
rect 1376 24987 1416 25019
rect 1448 24987 1488 25019
rect 1520 24987 1560 25019
rect 1592 24987 1632 25019
rect 1664 24987 1704 25019
rect 1736 24987 1776 25019
rect 1808 24987 1848 25019
rect 1880 24987 1950 25019
rect 50 24947 1950 24987
rect 50 24915 120 24947
rect 152 24915 192 24947
rect 224 24915 264 24947
rect 296 24915 336 24947
rect 368 24915 408 24947
rect 440 24915 480 24947
rect 512 24915 552 24947
rect 584 24915 624 24947
rect 656 24915 696 24947
rect 728 24915 768 24947
rect 800 24915 840 24947
rect 872 24915 912 24947
rect 944 24915 984 24947
rect 1016 24915 1056 24947
rect 1088 24915 1128 24947
rect 1160 24915 1200 24947
rect 1232 24915 1272 24947
rect 1304 24915 1344 24947
rect 1376 24915 1416 24947
rect 1448 24915 1488 24947
rect 1520 24915 1560 24947
rect 1592 24915 1632 24947
rect 1664 24915 1704 24947
rect 1736 24915 1776 24947
rect 1808 24915 1848 24947
rect 1880 24915 1950 24947
rect 50 24875 1950 24915
rect 50 24843 120 24875
rect 152 24843 192 24875
rect 224 24843 264 24875
rect 296 24843 336 24875
rect 368 24843 408 24875
rect 440 24843 480 24875
rect 512 24843 552 24875
rect 584 24843 624 24875
rect 656 24843 696 24875
rect 728 24843 768 24875
rect 800 24843 840 24875
rect 872 24843 912 24875
rect 944 24843 984 24875
rect 1016 24843 1056 24875
rect 1088 24843 1128 24875
rect 1160 24843 1200 24875
rect 1232 24843 1272 24875
rect 1304 24843 1344 24875
rect 1376 24843 1416 24875
rect 1448 24843 1488 24875
rect 1520 24843 1560 24875
rect 1592 24843 1632 24875
rect 1664 24843 1704 24875
rect 1736 24843 1776 24875
rect 1808 24843 1848 24875
rect 1880 24843 1950 24875
rect 50 24803 1950 24843
rect 50 24771 120 24803
rect 152 24771 192 24803
rect 224 24771 264 24803
rect 296 24771 336 24803
rect 368 24771 408 24803
rect 440 24771 480 24803
rect 512 24771 552 24803
rect 584 24771 624 24803
rect 656 24771 696 24803
rect 728 24771 768 24803
rect 800 24771 840 24803
rect 872 24771 912 24803
rect 944 24771 984 24803
rect 1016 24771 1056 24803
rect 1088 24771 1128 24803
rect 1160 24771 1200 24803
rect 1232 24771 1272 24803
rect 1304 24771 1344 24803
rect 1376 24771 1416 24803
rect 1448 24771 1488 24803
rect 1520 24771 1560 24803
rect 1592 24771 1632 24803
rect 1664 24771 1704 24803
rect 1736 24771 1776 24803
rect 1808 24771 1848 24803
rect 1880 24771 1950 24803
rect 50 24731 1950 24771
rect 50 24699 120 24731
rect 152 24699 192 24731
rect 224 24699 264 24731
rect 296 24699 336 24731
rect 368 24699 408 24731
rect 440 24699 480 24731
rect 512 24699 552 24731
rect 584 24699 624 24731
rect 656 24699 696 24731
rect 728 24699 768 24731
rect 800 24699 840 24731
rect 872 24699 912 24731
rect 944 24699 984 24731
rect 1016 24699 1056 24731
rect 1088 24699 1128 24731
rect 1160 24699 1200 24731
rect 1232 24699 1272 24731
rect 1304 24699 1344 24731
rect 1376 24699 1416 24731
rect 1448 24699 1488 24731
rect 1520 24699 1560 24731
rect 1592 24699 1632 24731
rect 1664 24699 1704 24731
rect 1736 24699 1776 24731
rect 1808 24699 1848 24731
rect 1880 24699 1950 24731
rect 50 24659 1950 24699
rect 50 24627 120 24659
rect 152 24627 192 24659
rect 224 24627 264 24659
rect 296 24627 336 24659
rect 368 24627 408 24659
rect 440 24627 480 24659
rect 512 24627 552 24659
rect 584 24627 624 24659
rect 656 24627 696 24659
rect 728 24627 768 24659
rect 800 24627 840 24659
rect 872 24627 912 24659
rect 944 24627 984 24659
rect 1016 24627 1056 24659
rect 1088 24627 1128 24659
rect 1160 24627 1200 24659
rect 1232 24627 1272 24659
rect 1304 24627 1344 24659
rect 1376 24627 1416 24659
rect 1448 24627 1488 24659
rect 1520 24627 1560 24659
rect 1592 24627 1632 24659
rect 1664 24627 1704 24659
rect 1736 24627 1776 24659
rect 1808 24627 1848 24659
rect 1880 24627 1950 24659
rect 50 24587 1950 24627
rect 50 24555 120 24587
rect 152 24555 192 24587
rect 224 24555 264 24587
rect 296 24555 336 24587
rect 368 24555 408 24587
rect 440 24555 480 24587
rect 512 24555 552 24587
rect 584 24555 624 24587
rect 656 24555 696 24587
rect 728 24555 768 24587
rect 800 24555 840 24587
rect 872 24555 912 24587
rect 944 24555 984 24587
rect 1016 24555 1056 24587
rect 1088 24555 1128 24587
rect 1160 24555 1200 24587
rect 1232 24555 1272 24587
rect 1304 24555 1344 24587
rect 1376 24555 1416 24587
rect 1448 24555 1488 24587
rect 1520 24555 1560 24587
rect 1592 24555 1632 24587
rect 1664 24555 1704 24587
rect 1736 24555 1776 24587
rect 1808 24555 1848 24587
rect 1880 24555 1950 24587
rect 50 24515 1950 24555
rect 50 24483 120 24515
rect 152 24483 192 24515
rect 224 24483 264 24515
rect 296 24483 336 24515
rect 368 24483 408 24515
rect 440 24483 480 24515
rect 512 24483 552 24515
rect 584 24483 624 24515
rect 656 24483 696 24515
rect 728 24483 768 24515
rect 800 24483 840 24515
rect 872 24483 912 24515
rect 944 24483 984 24515
rect 1016 24483 1056 24515
rect 1088 24483 1128 24515
rect 1160 24483 1200 24515
rect 1232 24483 1272 24515
rect 1304 24483 1344 24515
rect 1376 24483 1416 24515
rect 1448 24483 1488 24515
rect 1520 24483 1560 24515
rect 1592 24483 1632 24515
rect 1664 24483 1704 24515
rect 1736 24483 1776 24515
rect 1808 24483 1848 24515
rect 1880 24483 1950 24515
rect 50 24443 1950 24483
rect 50 24411 120 24443
rect 152 24411 192 24443
rect 224 24411 264 24443
rect 296 24411 336 24443
rect 368 24411 408 24443
rect 440 24411 480 24443
rect 512 24411 552 24443
rect 584 24411 624 24443
rect 656 24411 696 24443
rect 728 24411 768 24443
rect 800 24411 840 24443
rect 872 24411 912 24443
rect 944 24411 984 24443
rect 1016 24411 1056 24443
rect 1088 24411 1128 24443
rect 1160 24411 1200 24443
rect 1232 24411 1272 24443
rect 1304 24411 1344 24443
rect 1376 24411 1416 24443
rect 1448 24411 1488 24443
rect 1520 24411 1560 24443
rect 1592 24411 1632 24443
rect 1664 24411 1704 24443
rect 1736 24411 1776 24443
rect 1808 24411 1848 24443
rect 1880 24411 1950 24443
rect 50 24371 1950 24411
rect 50 24339 120 24371
rect 152 24339 192 24371
rect 224 24339 264 24371
rect 296 24339 336 24371
rect 368 24339 408 24371
rect 440 24339 480 24371
rect 512 24339 552 24371
rect 584 24339 624 24371
rect 656 24339 696 24371
rect 728 24339 768 24371
rect 800 24339 840 24371
rect 872 24339 912 24371
rect 944 24339 984 24371
rect 1016 24339 1056 24371
rect 1088 24339 1128 24371
rect 1160 24339 1200 24371
rect 1232 24339 1272 24371
rect 1304 24339 1344 24371
rect 1376 24339 1416 24371
rect 1448 24339 1488 24371
rect 1520 24339 1560 24371
rect 1592 24339 1632 24371
rect 1664 24339 1704 24371
rect 1736 24339 1776 24371
rect 1808 24339 1848 24371
rect 1880 24339 1950 24371
rect 50 24299 1950 24339
rect 50 24267 120 24299
rect 152 24267 192 24299
rect 224 24267 264 24299
rect 296 24267 336 24299
rect 368 24267 408 24299
rect 440 24267 480 24299
rect 512 24267 552 24299
rect 584 24267 624 24299
rect 656 24267 696 24299
rect 728 24267 768 24299
rect 800 24267 840 24299
rect 872 24267 912 24299
rect 944 24267 984 24299
rect 1016 24267 1056 24299
rect 1088 24267 1128 24299
rect 1160 24267 1200 24299
rect 1232 24267 1272 24299
rect 1304 24267 1344 24299
rect 1376 24267 1416 24299
rect 1448 24267 1488 24299
rect 1520 24267 1560 24299
rect 1592 24267 1632 24299
rect 1664 24267 1704 24299
rect 1736 24267 1776 24299
rect 1808 24267 1848 24299
rect 1880 24267 1950 24299
rect 50 24227 1950 24267
rect 50 24195 120 24227
rect 152 24195 192 24227
rect 224 24195 264 24227
rect 296 24195 336 24227
rect 368 24195 408 24227
rect 440 24195 480 24227
rect 512 24195 552 24227
rect 584 24195 624 24227
rect 656 24195 696 24227
rect 728 24195 768 24227
rect 800 24195 840 24227
rect 872 24195 912 24227
rect 944 24195 984 24227
rect 1016 24195 1056 24227
rect 1088 24195 1128 24227
rect 1160 24195 1200 24227
rect 1232 24195 1272 24227
rect 1304 24195 1344 24227
rect 1376 24195 1416 24227
rect 1448 24195 1488 24227
rect 1520 24195 1560 24227
rect 1592 24195 1632 24227
rect 1664 24195 1704 24227
rect 1736 24195 1776 24227
rect 1808 24195 1848 24227
rect 1880 24195 1950 24227
rect 50 24155 1950 24195
rect 50 24123 120 24155
rect 152 24123 192 24155
rect 224 24123 264 24155
rect 296 24123 336 24155
rect 368 24123 408 24155
rect 440 24123 480 24155
rect 512 24123 552 24155
rect 584 24123 624 24155
rect 656 24123 696 24155
rect 728 24123 768 24155
rect 800 24123 840 24155
rect 872 24123 912 24155
rect 944 24123 984 24155
rect 1016 24123 1056 24155
rect 1088 24123 1128 24155
rect 1160 24123 1200 24155
rect 1232 24123 1272 24155
rect 1304 24123 1344 24155
rect 1376 24123 1416 24155
rect 1448 24123 1488 24155
rect 1520 24123 1560 24155
rect 1592 24123 1632 24155
rect 1664 24123 1704 24155
rect 1736 24123 1776 24155
rect 1808 24123 1848 24155
rect 1880 24123 1950 24155
rect 50 24083 1950 24123
rect 50 24051 120 24083
rect 152 24051 192 24083
rect 224 24051 264 24083
rect 296 24051 336 24083
rect 368 24051 408 24083
rect 440 24051 480 24083
rect 512 24051 552 24083
rect 584 24051 624 24083
rect 656 24051 696 24083
rect 728 24051 768 24083
rect 800 24051 840 24083
rect 872 24051 912 24083
rect 944 24051 984 24083
rect 1016 24051 1056 24083
rect 1088 24051 1128 24083
rect 1160 24051 1200 24083
rect 1232 24051 1272 24083
rect 1304 24051 1344 24083
rect 1376 24051 1416 24083
rect 1448 24051 1488 24083
rect 1520 24051 1560 24083
rect 1592 24051 1632 24083
rect 1664 24051 1704 24083
rect 1736 24051 1776 24083
rect 1808 24051 1848 24083
rect 1880 24051 1950 24083
rect 50 24011 1950 24051
rect 50 23979 120 24011
rect 152 23979 192 24011
rect 224 23979 264 24011
rect 296 23979 336 24011
rect 368 23979 408 24011
rect 440 23979 480 24011
rect 512 23979 552 24011
rect 584 23979 624 24011
rect 656 23979 696 24011
rect 728 23979 768 24011
rect 800 23979 840 24011
rect 872 23979 912 24011
rect 944 23979 984 24011
rect 1016 23979 1056 24011
rect 1088 23979 1128 24011
rect 1160 23979 1200 24011
rect 1232 23979 1272 24011
rect 1304 23979 1344 24011
rect 1376 23979 1416 24011
rect 1448 23979 1488 24011
rect 1520 23979 1560 24011
rect 1592 23979 1632 24011
rect 1664 23979 1704 24011
rect 1736 23979 1776 24011
rect 1808 23979 1848 24011
rect 1880 23979 1950 24011
rect 50 23939 1950 23979
rect 50 23907 120 23939
rect 152 23907 192 23939
rect 224 23907 264 23939
rect 296 23907 336 23939
rect 368 23907 408 23939
rect 440 23907 480 23939
rect 512 23907 552 23939
rect 584 23907 624 23939
rect 656 23907 696 23939
rect 728 23907 768 23939
rect 800 23907 840 23939
rect 872 23907 912 23939
rect 944 23907 984 23939
rect 1016 23907 1056 23939
rect 1088 23907 1128 23939
rect 1160 23907 1200 23939
rect 1232 23907 1272 23939
rect 1304 23907 1344 23939
rect 1376 23907 1416 23939
rect 1448 23907 1488 23939
rect 1520 23907 1560 23939
rect 1592 23907 1632 23939
rect 1664 23907 1704 23939
rect 1736 23907 1776 23939
rect 1808 23907 1848 23939
rect 1880 23907 1950 23939
rect 50 23867 1950 23907
rect 50 23835 120 23867
rect 152 23835 192 23867
rect 224 23835 264 23867
rect 296 23835 336 23867
rect 368 23835 408 23867
rect 440 23835 480 23867
rect 512 23835 552 23867
rect 584 23835 624 23867
rect 656 23835 696 23867
rect 728 23835 768 23867
rect 800 23835 840 23867
rect 872 23835 912 23867
rect 944 23835 984 23867
rect 1016 23835 1056 23867
rect 1088 23835 1128 23867
rect 1160 23835 1200 23867
rect 1232 23835 1272 23867
rect 1304 23835 1344 23867
rect 1376 23835 1416 23867
rect 1448 23835 1488 23867
rect 1520 23835 1560 23867
rect 1592 23835 1632 23867
rect 1664 23835 1704 23867
rect 1736 23835 1776 23867
rect 1808 23835 1848 23867
rect 1880 23835 1950 23867
rect 50 23795 1950 23835
rect 50 23763 120 23795
rect 152 23763 192 23795
rect 224 23763 264 23795
rect 296 23763 336 23795
rect 368 23763 408 23795
rect 440 23763 480 23795
rect 512 23763 552 23795
rect 584 23763 624 23795
rect 656 23763 696 23795
rect 728 23763 768 23795
rect 800 23763 840 23795
rect 872 23763 912 23795
rect 944 23763 984 23795
rect 1016 23763 1056 23795
rect 1088 23763 1128 23795
rect 1160 23763 1200 23795
rect 1232 23763 1272 23795
rect 1304 23763 1344 23795
rect 1376 23763 1416 23795
rect 1448 23763 1488 23795
rect 1520 23763 1560 23795
rect 1592 23763 1632 23795
rect 1664 23763 1704 23795
rect 1736 23763 1776 23795
rect 1808 23763 1848 23795
rect 1880 23763 1950 23795
rect 50 23723 1950 23763
rect 50 23691 120 23723
rect 152 23691 192 23723
rect 224 23691 264 23723
rect 296 23691 336 23723
rect 368 23691 408 23723
rect 440 23691 480 23723
rect 512 23691 552 23723
rect 584 23691 624 23723
rect 656 23691 696 23723
rect 728 23691 768 23723
rect 800 23691 840 23723
rect 872 23691 912 23723
rect 944 23691 984 23723
rect 1016 23691 1056 23723
rect 1088 23691 1128 23723
rect 1160 23691 1200 23723
rect 1232 23691 1272 23723
rect 1304 23691 1344 23723
rect 1376 23691 1416 23723
rect 1448 23691 1488 23723
rect 1520 23691 1560 23723
rect 1592 23691 1632 23723
rect 1664 23691 1704 23723
rect 1736 23691 1776 23723
rect 1808 23691 1848 23723
rect 1880 23691 1950 23723
rect 50 23651 1950 23691
rect 50 23619 120 23651
rect 152 23619 192 23651
rect 224 23619 264 23651
rect 296 23619 336 23651
rect 368 23619 408 23651
rect 440 23619 480 23651
rect 512 23619 552 23651
rect 584 23619 624 23651
rect 656 23619 696 23651
rect 728 23619 768 23651
rect 800 23619 840 23651
rect 872 23619 912 23651
rect 944 23619 984 23651
rect 1016 23619 1056 23651
rect 1088 23619 1128 23651
rect 1160 23619 1200 23651
rect 1232 23619 1272 23651
rect 1304 23619 1344 23651
rect 1376 23619 1416 23651
rect 1448 23619 1488 23651
rect 1520 23619 1560 23651
rect 1592 23619 1632 23651
rect 1664 23619 1704 23651
rect 1736 23619 1776 23651
rect 1808 23619 1848 23651
rect 1880 23619 1950 23651
rect 50 23579 1950 23619
rect 50 23547 120 23579
rect 152 23547 192 23579
rect 224 23547 264 23579
rect 296 23547 336 23579
rect 368 23547 408 23579
rect 440 23547 480 23579
rect 512 23547 552 23579
rect 584 23547 624 23579
rect 656 23547 696 23579
rect 728 23547 768 23579
rect 800 23547 840 23579
rect 872 23547 912 23579
rect 944 23547 984 23579
rect 1016 23547 1056 23579
rect 1088 23547 1128 23579
rect 1160 23547 1200 23579
rect 1232 23547 1272 23579
rect 1304 23547 1344 23579
rect 1376 23547 1416 23579
rect 1448 23547 1488 23579
rect 1520 23547 1560 23579
rect 1592 23547 1632 23579
rect 1664 23547 1704 23579
rect 1736 23547 1776 23579
rect 1808 23547 1848 23579
rect 1880 23547 1950 23579
rect 50 23507 1950 23547
rect 50 23475 120 23507
rect 152 23475 192 23507
rect 224 23475 264 23507
rect 296 23475 336 23507
rect 368 23475 408 23507
rect 440 23475 480 23507
rect 512 23475 552 23507
rect 584 23475 624 23507
rect 656 23475 696 23507
rect 728 23475 768 23507
rect 800 23475 840 23507
rect 872 23475 912 23507
rect 944 23475 984 23507
rect 1016 23475 1056 23507
rect 1088 23475 1128 23507
rect 1160 23475 1200 23507
rect 1232 23475 1272 23507
rect 1304 23475 1344 23507
rect 1376 23475 1416 23507
rect 1448 23475 1488 23507
rect 1520 23475 1560 23507
rect 1592 23475 1632 23507
rect 1664 23475 1704 23507
rect 1736 23475 1776 23507
rect 1808 23475 1848 23507
rect 1880 23475 1950 23507
rect 50 23435 1950 23475
rect 50 23403 120 23435
rect 152 23403 192 23435
rect 224 23403 264 23435
rect 296 23403 336 23435
rect 368 23403 408 23435
rect 440 23403 480 23435
rect 512 23403 552 23435
rect 584 23403 624 23435
rect 656 23403 696 23435
rect 728 23403 768 23435
rect 800 23403 840 23435
rect 872 23403 912 23435
rect 944 23403 984 23435
rect 1016 23403 1056 23435
rect 1088 23403 1128 23435
rect 1160 23403 1200 23435
rect 1232 23403 1272 23435
rect 1304 23403 1344 23435
rect 1376 23403 1416 23435
rect 1448 23403 1488 23435
rect 1520 23403 1560 23435
rect 1592 23403 1632 23435
rect 1664 23403 1704 23435
rect 1736 23403 1776 23435
rect 1808 23403 1848 23435
rect 1880 23403 1950 23435
rect 50 23363 1950 23403
rect 50 23331 120 23363
rect 152 23331 192 23363
rect 224 23331 264 23363
rect 296 23331 336 23363
rect 368 23331 408 23363
rect 440 23331 480 23363
rect 512 23331 552 23363
rect 584 23331 624 23363
rect 656 23331 696 23363
rect 728 23331 768 23363
rect 800 23331 840 23363
rect 872 23331 912 23363
rect 944 23331 984 23363
rect 1016 23331 1056 23363
rect 1088 23331 1128 23363
rect 1160 23331 1200 23363
rect 1232 23331 1272 23363
rect 1304 23331 1344 23363
rect 1376 23331 1416 23363
rect 1448 23331 1488 23363
rect 1520 23331 1560 23363
rect 1592 23331 1632 23363
rect 1664 23331 1704 23363
rect 1736 23331 1776 23363
rect 1808 23331 1848 23363
rect 1880 23331 1950 23363
rect 50 23291 1950 23331
rect 50 23259 120 23291
rect 152 23259 192 23291
rect 224 23259 264 23291
rect 296 23259 336 23291
rect 368 23259 408 23291
rect 440 23259 480 23291
rect 512 23259 552 23291
rect 584 23259 624 23291
rect 656 23259 696 23291
rect 728 23259 768 23291
rect 800 23259 840 23291
rect 872 23259 912 23291
rect 944 23259 984 23291
rect 1016 23259 1056 23291
rect 1088 23259 1128 23291
rect 1160 23259 1200 23291
rect 1232 23259 1272 23291
rect 1304 23259 1344 23291
rect 1376 23259 1416 23291
rect 1448 23259 1488 23291
rect 1520 23259 1560 23291
rect 1592 23259 1632 23291
rect 1664 23259 1704 23291
rect 1736 23259 1776 23291
rect 1808 23259 1848 23291
rect 1880 23259 1950 23291
rect 50 23219 1950 23259
rect 50 23187 120 23219
rect 152 23187 192 23219
rect 224 23187 264 23219
rect 296 23187 336 23219
rect 368 23187 408 23219
rect 440 23187 480 23219
rect 512 23187 552 23219
rect 584 23187 624 23219
rect 656 23187 696 23219
rect 728 23187 768 23219
rect 800 23187 840 23219
rect 872 23187 912 23219
rect 944 23187 984 23219
rect 1016 23187 1056 23219
rect 1088 23187 1128 23219
rect 1160 23187 1200 23219
rect 1232 23187 1272 23219
rect 1304 23187 1344 23219
rect 1376 23187 1416 23219
rect 1448 23187 1488 23219
rect 1520 23187 1560 23219
rect 1592 23187 1632 23219
rect 1664 23187 1704 23219
rect 1736 23187 1776 23219
rect 1808 23187 1848 23219
rect 1880 23187 1950 23219
rect 50 23124 1950 23187
rect 50 22874 1950 22924
rect 50 22842 120 22874
rect 152 22842 192 22874
rect 224 22842 264 22874
rect 296 22842 336 22874
rect 368 22842 408 22874
rect 440 22842 480 22874
rect 512 22842 552 22874
rect 584 22842 624 22874
rect 656 22842 696 22874
rect 728 22842 768 22874
rect 800 22842 840 22874
rect 872 22842 912 22874
rect 944 22842 984 22874
rect 1016 22842 1056 22874
rect 1088 22842 1128 22874
rect 1160 22842 1200 22874
rect 1232 22842 1272 22874
rect 1304 22842 1344 22874
rect 1376 22842 1416 22874
rect 1448 22842 1488 22874
rect 1520 22842 1560 22874
rect 1592 22842 1632 22874
rect 1664 22842 1704 22874
rect 1736 22842 1776 22874
rect 1808 22842 1848 22874
rect 1880 22842 1950 22874
rect 50 22802 1950 22842
rect 50 22770 120 22802
rect 152 22770 192 22802
rect 224 22770 264 22802
rect 296 22770 336 22802
rect 368 22770 408 22802
rect 440 22770 480 22802
rect 512 22770 552 22802
rect 584 22770 624 22802
rect 656 22770 696 22802
rect 728 22770 768 22802
rect 800 22770 840 22802
rect 872 22770 912 22802
rect 944 22770 984 22802
rect 1016 22770 1056 22802
rect 1088 22770 1128 22802
rect 1160 22770 1200 22802
rect 1232 22770 1272 22802
rect 1304 22770 1344 22802
rect 1376 22770 1416 22802
rect 1448 22770 1488 22802
rect 1520 22770 1560 22802
rect 1592 22770 1632 22802
rect 1664 22770 1704 22802
rect 1736 22770 1776 22802
rect 1808 22770 1848 22802
rect 1880 22770 1950 22802
rect 50 22730 1950 22770
rect 50 22698 120 22730
rect 152 22698 192 22730
rect 224 22698 264 22730
rect 296 22698 336 22730
rect 368 22698 408 22730
rect 440 22698 480 22730
rect 512 22698 552 22730
rect 584 22698 624 22730
rect 656 22698 696 22730
rect 728 22698 768 22730
rect 800 22698 840 22730
rect 872 22698 912 22730
rect 944 22698 984 22730
rect 1016 22698 1056 22730
rect 1088 22698 1128 22730
rect 1160 22698 1200 22730
rect 1232 22698 1272 22730
rect 1304 22698 1344 22730
rect 1376 22698 1416 22730
rect 1448 22698 1488 22730
rect 1520 22698 1560 22730
rect 1592 22698 1632 22730
rect 1664 22698 1704 22730
rect 1736 22698 1776 22730
rect 1808 22698 1848 22730
rect 1880 22698 1950 22730
rect 50 22658 1950 22698
rect 50 22626 120 22658
rect 152 22626 192 22658
rect 224 22626 264 22658
rect 296 22626 336 22658
rect 368 22626 408 22658
rect 440 22626 480 22658
rect 512 22626 552 22658
rect 584 22626 624 22658
rect 656 22626 696 22658
rect 728 22626 768 22658
rect 800 22626 840 22658
rect 872 22626 912 22658
rect 944 22626 984 22658
rect 1016 22626 1056 22658
rect 1088 22626 1128 22658
rect 1160 22626 1200 22658
rect 1232 22626 1272 22658
rect 1304 22626 1344 22658
rect 1376 22626 1416 22658
rect 1448 22626 1488 22658
rect 1520 22626 1560 22658
rect 1592 22626 1632 22658
rect 1664 22626 1704 22658
rect 1736 22626 1776 22658
rect 1808 22626 1848 22658
rect 1880 22626 1950 22658
rect 50 22586 1950 22626
rect 50 22554 120 22586
rect 152 22554 192 22586
rect 224 22554 264 22586
rect 296 22554 336 22586
rect 368 22554 408 22586
rect 440 22554 480 22586
rect 512 22554 552 22586
rect 584 22554 624 22586
rect 656 22554 696 22586
rect 728 22554 768 22586
rect 800 22554 840 22586
rect 872 22554 912 22586
rect 944 22554 984 22586
rect 1016 22554 1056 22586
rect 1088 22554 1128 22586
rect 1160 22554 1200 22586
rect 1232 22554 1272 22586
rect 1304 22554 1344 22586
rect 1376 22554 1416 22586
rect 1448 22554 1488 22586
rect 1520 22554 1560 22586
rect 1592 22554 1632 22586
rect 1664 22554 1704 22586
rect 1736 22554 1776 22586
rect 1808 22554 1848 22586
rect 1880 22554 1950 22586
rect 50 22514 1950 22554
rect 50 22482 120 22514
rect 152 22482 192 22514
rect 224 22482 264 22514
rect 296 22482 336 22514
rect 368 22482 408 22514
rect 440 22482 480 22514
rect 512 22482 552 22514
rect 584 22482 624 22514
rect 656 22482 696 22514
rect 728 22482 768 22514
rect 800 22482 840 22514
rect 872 22482 912 22514
rect 944 22482 984 22514
rect 1016 22482 1056 22514
rect 1088 22482 1128 22514
rect 1160 22482 1200 22514
rect 1232 22482 1272 22514
rect 1304 22482 1344 22514
rect 1376 22482 1416 22514
rect 1448 22482 1488 22514
rect 1520 22482 1560 22514
rect 1592 22482 1632 22514
rect 1664 22482 1704 22514
rect 1736 22482 1776 22514
rect 1808 22482 1848 22514
rect 1880 22482 1950 22514
rect 50 22442 1950 22482
rect 50 22410 120 22442
rect 152 22410 192 22442
rect 224 22410 264 22442
rect 296 22410 336 22442
rect 368 22410 408 22442
rect 440 22410 480 22442
rect 512 22410 552 22442
rect 584 22410 624 22442
rect 656 22410 696 22442
rect 728 22410 768 22442
rect 800 22410 840 22442
rect 872 22410 912 22442
rect 944 22410 984 22442
rect 1016 22410 1056 22442
rect 1088 22410 1128 22442
rect 1160 22410 1200 22442
rect 1232 22410 1272 22442
rect 1304 22410 1344 22442
rect 1376 22410 1416 22442
rect 1448 22410 1488 22442
rect 1520 22410 1560 22442
rect 1592 22410 1632 22442
rect 1664 22410 1704 22442
rect 1736 22410 1776 22442
rect 1808 22410 1848 22442
rect 1880 22410 1950 22442
rect 50 22370 1950 22410
rect 50 22338 120 22370
rect 152 22338 192 22370
rect 224 22338 264 22370
rect 296 22338 336 22370
rect 368 22338 408 22370
rect 440 22338 480 22370
rect 512 22338 552 22370
rect 584 22338 624 22370
rect 656 22338 696 22370
rect 728 22338 768 22370
rect 800 22338 840 22370
rect 872 22338 912 22370
rect 944 22338 984 22370
rect 1016 22338 1056 22370
rect 1088 22338 1128 22370
rect 1160 22338 1200 22370
rect 1232 22338 1272 22370
rect 1304 22338 1344 22370
rect 1376 22338 1416 22370
rect 1448 22338 1488 22370
rect 1520 22338 1560 22370
rect 1592 22338 1632 22370
rect 1664 22338 1704 22370
rect 1736 22338 1776 22370
rect 1808 22338 1848 22370
rect 1880 22338 1950 22370
rect 50 22298 1950 22338
rect 50 22266 120 22298
rect 152 22266 192 22298
rect 224 22266 264 22298
rect 296 22266 336 22298
rect 368 22266 408 22298
rect 440 22266 480 22298
rect 512 22266 552 22298
rect 584 22266 624 22298
rect 656 22266 696 22298
rect 728 22266 768 22298
rect 800 22266 840 22298
rect 872 22266 912 22298
rect 944 22266 984 22298
rect 1016 22266 1056 22298
rect 1088 22266 1128 22298
rect 1160 22266 1200 22298
rect 1232 22266 1272 22298
rect 1304 22266 1344 22298
rect 1376 22266 1416 22298
rect 1448 22266 1488 22298
rect 1520 22266 1560 22298
rect 1592 22266 1632 22298
rect 1664 22266 1704 22298
rect 1736 22266 1776 22298
rect 1808 22266 1848 22298
rect 1880 22266 1950 22298
rect 50 22226 1950 22266
rect 50 22194 120 22226
rect 152 22194 192 22226
rect 224 22194 264 22226
rect 296 22194 336 22226
rect 368 22194 408 22226
rect 440 22194 480 22226
rect 512 22194 552 22226
rect 584 22194 624 22226
rect 656 22194 696 22226
rect 728 22194 768 22226
rect 800 22194 840 22226
rect 872 22194 912 22226
rect 944 22194 984 22226
rect 1016 22194 1056 22226
rect 1088 22194 1128 22226
rect 1160 22194 1200 22226
rect 1232 22194 1272 22226
rect 1304 22194 1344 22226
rect 1376 22194 1416 22226
rect 1448 22194 1488 22226
rect 1520 22194 1560 22226
rect 1592 22194 1632 22226
rect 1664 22194 1704 22226
rect 1736 22194 1776 22226
rect 1808 22194 1848 22226
rect 1880 22194 1950 22226
rect 50 22154 1950 22194
rect 50 22122 120 22154
rect 152 22122 192 22154
rect 224 22122 264 22154
rect 296 22122 336 22154
rect 368 22122 408 22154
rect 440 22122 480 22154
rect 512 22122 552 22154
rect 584 22122 624 22154
rect 656 22122 696 22154
rect 728 22122 768 22154
rect 800 22122 840 22154
rect 872 22122 912 22154
rect 944 22122 984 22154
rect 1016 22122 1056 22154
rect 1088 22122 1128 22154
rect 1160 22122 1200 22154
rect 1232 22122 1272 22154
rect 1304 22122 1344 22154
rect 1376 22122 1416 22154
rect 1448 22122 1488 22154
rect 1520 22122 1560 22154
rect 1592 22122 1632 22154
rect 1664 22122 1704 22154
rect 1736 22122 1776 22154
rect 1808 22122 1848 22154
rect 1880 22122 1950 22154
rect 50 22082 1950 22122
rect 50 22050 120 22082
rect 152 22050 192 22082
rect 224 22050 264 22082
rect 296 22050 336 22082
rect 368 22050 408 22082
rect 440 22050 480 22082
rect 512 22050 552 22082
rect 584 22050 624 22082
rect 656 22050 696 22082
rect 728 22050 768 22082
rect 800 22050 840 22082
rect 872 22050 912 22082
rect 944 22050 984 22082
rect 1016 22050 1056 22082
rect 1088 22050 1128 22082
rect 1160 22050 1200 22082
rect 1232 22050 1272 22082
rect 1304 22050 1344 22082
rect 1376 22050 1416 22082
rect 1448 22050 1488 22082
rect 1520 22050 1560 22082
rect 1592 22050 1632 22082
rect 1664 22050 1704 22082
rect 1736 22050 1776 22082
rect 1808 22050 1848 22082
rect 1880 22050 1950 22082
rect 50 22010 1950 22050
rect 50 21978 120 22010
rect 152 21978 192 22010
rect 224 21978 264 22010
rect 296 21978 336 22010
rect 368 21978 408 22010
rect 440 21978 480 22010
rect 512 21978 552 22010
rect 584 21978 624 22010
rect 656 21978 696 22010
rect 728 21978 768 22010
rect 800 21978 840 22010
rect 872 21978 912 22010
rect 944 21978 984 22010
rect 1016 21978 1056 22010
rect 1088 21978 1128 22010
rect 1160 21978 1200 22010
rect 1232 21978 1272 22010
rect 1304 21978 1344 22010
rect 1376 21978 1416 22010
rect 1448 21978 1488 22010
rect 1520 21978 1560 22010
rect 1592 21978 1632 22010
rect 1664 21978 1704 22010
rect 1736 21978 1776 22010
rect 1808 21978 1848 22010
rect 1880 21978 1950 22010
rect 50 21938 1950 21978
rect 50 21906 120 21938
rect 152 21906 192 21938
rect 224 21906 264 21938
rect 296 21906 336 21938
rect 368 21906 408 21938
rect 440 21906 480 21938
rect 512 21906 552 21938
rect 584 21906 624 21938
rect 656 21906 696 21938
rect 728 21906 768 21938
rect 800 21906 840 21938
rect 872 21906 912 21938
rect 944 21906 984 21938
rect 1016 21906 1056 21938
rect 1088 21906 1128 21938
rect 1160 21906 1200 21938
rect 1232 21906 1272 21938
rect 1304 21906 1344 21938
rect 1376 21906 1416 21938
rect 1448 21906 1488 21938
rect 1520 21906 1560 21938
rect 1592 21906 1632 21938
rect 1664 21906 1704 21938
rect 1736 21906 1776 21938
rect 1808 21906 1848 21938
rect 1880 21906 1950 21938
rect 50 21866 1950 21906
rect 50 21834 120 21866
rect 152 21834 192 21866
rect 224 21834 264 21866
rect 296 21834 336 21866
rect 368 21834 408 21866
rect 440 21834 480 21866
rect 512 21834 552 21866
rect 584 21834 624 21866
rect 656 21834 696 21866
rect 728 21834 768 21866
rect 800 21834 840 21866
rect 872 21834 912 21866
rect 944 21834 984 21866
rect 1016 21834 1056 21866
rect 1088 21834 1128 21866
rect 1160 21834 1200 21866
rect 1232 21834 1272 21866
rect 1304 21834 1344 21866
rect 1376 21834 1416 21866
rect 1448 21834 1488 21866
rect 1520 21834 1560 21866
rect 1592 21834 1632 21866
rect 1664 21834 1704 21866
rect 1736 21834 1776 21866
rect 1808 21834 1848 21866
rect 1880 21834 1950 21866
rect 50 21794 1950 21834
rect 50 21762 120 21794
rect 152 21762 192 21794
rect 224 21762 264 21794
rect 296 21762 336 21794
rect 368 21762 408 21794
rect 440 21762 480 21794
rect 512 21762 552 21794
rect 584 21762 624 21794
rect 656 21762 696 21794
rect 728 21762 768 21794
rect 800 21762 840 21794
rect 872 21762 912 21794
rect 944 21762 984 21794
rect 1016 21762 1056 21794
rect 1088 21762 1128 21794
rect 1160 21762 1200 21794
rect 1232 21762 1272 21794
rect 1304 21762 1344 21794
rect 1376 21762 1416 21794
rect 1448 21762 1488 21794
rect 1520 21762 1560 21794
rect 1592 21762 1632 21794
rect 1664 21762 1704 21794
rect 1736 21762 1776 21794
rect 1808 21762 1848 21794
rect 1880 21762 1950 21794
rect 50 21722 1950 21762
rect 50 21690 120 21722
rect 152 21690 192 21722
rect 224 21690 264 21722
rect 296 21690 336 21722
rect 368 21690 408 21722
rect 440 21690 480 21722
rect 512 21690 552 21722
rect 584 21690 624 21722
rect 656 21690 696 21722
rect 728 21690 768 21722
rect 800 21690 840 21722
rect 872 21690 912 21722
rect 944 21690 984 21722
rect 1016 21690 1056 21722
rect 1088 21690 1128 21722
rect 1160 21690 1200 21722
rect 1232 21690 1272 21722
rect 1304 21690 1344 21722
rect 1376 21690 1416 21722
rect 1448 21690 1488 21722
rect 1520 21690 1560 21722
rect 1592 21690 1632 21722
rect 1664 21690 1704 21722
rect 1736 21690 1776 21722
rect 1808 21690 1848 21722
rect 1880 21690 1950 21722
rect 50 21650 1950 21690
rect 50 21618 120 21650
rect 152 21618 192 21650
rect 224 21618 264 21650
rect 296 21618 336 21650
rect 368 21618 408 21650
rect 440 21618 480 21650
rect 512 21618 552 21650
rect 584 21618 624 21650
rect 656 21618 696 21650
rect 728 21618 768 21650
rect 800 21618 840 21650
rect 872 21618 912 21650
rect 944 21618 984 21650
rect 1016 21618 1056 21650
rect 1088 21618 1128 21650
rect 1160 21618 1200 21650
rect 1232 21618 1272 21650
rect 1304 21618 1344 21650
rect 1376 21618 1416 21650
rect 1448 21618 1488 21650
rect 1520 21618 1560 21650
rect 1592 21618 1632 21650
rect 1664 21618 1704 21650
rect 1736 21618 1776 21650
rect 1808 21618 1848 21650
rect 1880 21618 1950 21650
rect 50 21578 1950 21618
rect 50 21546 120 21578
rect 152 21546 192 21578
rect 224 21546 264 21578
rect 296 21546 336 21578
rect 368 21546 408 21578
rect 440 21546 480 21578
rect 512 21546 552 21578
rect 584 21546 624 21578
rect 656 21546 696 21578
rect 728 21546 768 21578
rect 800 21546 840 21578
rect 872 21546 912 21578
rect 944 21546 984 21578
rect 1016 21546 1056 21578
rect 1088 21546 1128 21578
rect 1160 21546 1200 21578
rect 1232 21546 1272 21578
rect 1304 21546 1344 21578
rect 1376 21546 1416 21578
rect 1448 21546 1488 21578
rect 1520 21546 1560 21578
rect 1592 21546 1632 21578
rect 1664 21546 1704 21578
rect 1736 21546 1776 21578
rect 1808 21546 1848 21578
rect 1880 21546 1950 21578
rect 50 21506 1950 21546
rect 50 21474 120 21506
rect 152 21474 192 21506
rect 224 21474 264 21506
rect 296 21474 336 21506
rect 368 21474 408 21506
rect 440 21474 480 21506
rect 512 21474 552 21506
rect 584 21474 624 21506
rect 656 21474 696 21506
rect 728 21474 768 21506
rect 800 21474 840 21506
rect 872 21474 912 21506
rect 944 21474 984 21506
rect 1016 21474 1056 21506
rect 1088 21474 1128 21506
rect 1160 21474 1200 21506
rect 1232 21474 1272 21506
rect 1304 21474 1344 21506
rect 1376 21474 1416 21506
rect 1448 21474 1488 21506
rect 1520 21474 1560 21506
rect 1592 21474 1632 21506
rect 1664 21474 1704 21506
rect 1736 21474 1776 21506
rect 1808 21474 1848 21506
rect 1880 21474 1950 21506
rect 50 21434 1950 21474
rect 50 21402 120 21434
rect 152 21402 192 21434
rect 224 21402 264 21434
rect 296 21402 336 21434
rect 368 21402 408 21434
rect 440 21402 480 21434
rect 512 21402 552 21434
rect 584 21402 624 21434
rect 656 21402 696 21434
rect 728 21402 768 21434
rect 800 21402 840 21434
rect 872 21402 912 21434
rect 944 21402 984 21434
rect 1016 21402 1056 21434
rect 1088 21402 1128 21434
rect 1160 21402 1200 21434
rect 1232 21402 1272 21434
rect 1304 21402 1344 21434
rect 1376 21402 1416 21434
rect 1448 21402 1488 21434
rect 1520 21402 1560 21434
rect 1592 21402 1632 21434
rect 1664 21402 1704 21434
rect 1736 21402 1776 21434
rect 1808 21402 1848 21434
rect 1880 21402 1950 21434
rect 50 21362 1950 21402
rect 50 21330 120 21362
rect 152 21330 192 21362
rect 224 21330 264 21362
rect 296 21330 336 21362
rect 368 21330 408 21362
rect 440 21330 480 21362
rect 512 21330 552 21362
rect 584 21330 624 21362
rect 656 21330 696 21362
rect 728 21330 768 21362
rect 800 21330 840 21362
rect 872 21330 912 21362
rect 944 21330 984 21362
rect 1016 21330 1056 21362
rect 1088 21330 1128 21362
rect 1160 21330 1200 21362
rect 1232 21330 1272 21362
rect 1304 21330 1344 21362
rect 1376 21330 1416 21362
rect 1448 21330 1488 21362
rect 1520 21330 1560 21362
rect 1592 21330 1632 21362
rect 1664 21330 1704 21362
rect 1736 21330 1776 21362
rect 1808 21330 1848 21362
rect 1880 21330 1950 21362
rect 50 21290 1950 21330
rect 50 21258 120 21290
rect 152 21258 192 21290
rect 224 21258 264 21290
rect 296 21258 336 21290
rect 368 21258 408 21290
rect 440 21258 480 21290
rect 512 21258 552 21290
rect 584 21258 624 21290
rect 656 21258 696 21290
rect 728 21258 768 21290
rect 800 21258 840 21290
rect 872 21258 912 21290
rect 944 21258 984 21290
rect 1016 21258 1056 21290
rect 1088 21258 1128 21290
rect 1160 21258 1200 21290
rect 1232 21258 1272 21290
rect 1304 21258 1344 21290
rect 1376 21258 1416 21290
rect 1448 21258 1488 21290
rect 1520 21258 1560 21290
rect 1592 21258 1632 21290
rect 1664 21258 1704 21290
rect 1736 21258 1776 21290
rect 1808 21258 1848 21290
rect 1880 21258 1950 21290
rect 50 21218 1950 21258
rect 50 21186 120 21218
rect 152 21186 192 21218
rect 224 21186 264 21218
rect 296 21186 336 21218
rect 368 21186 408 21218
rect 440 21186 480 21218
rect 512 21186 552 21218
rect 584 21186 624 21218
rect 656 21186 696 21218
rect 728 21186 768 21218
rect 800 21186 840 21218
rect 872 21186 912 21218
rect 944 21186 984 21218
rect 1016 21186 1056 21218
rect 1088 21186 1128 21218
rect 1160 21186 1200 21218
rect 1232 21186 1272 21218
rect 1304 21186 1344 21218
rect 1376 21186 1416 21218
rect 1448 21186 1488 21218
rect 1520 21186 1560 21218
rect 1592 21186 1632 21218
rect 1664 21186 1704 21218
rect 1736 21186 1776 21218
rect 1808 21186 1848 21218
rect 1880 21186 1950 21218
rect 50 21146 1950 21186
rect 50 21114 120 21146
rect 152 21114 192 21146
rect 224 21114 264 21146
rect 296 21114 336 21146
rect 368 21114 408 21146
rect 440 21114 480 21146
rect 512 21114 552 21146
rect 584 21114 624 21146
rect 656 21114 696 21146
rect 728 21114 768 21146
rect 800 21114 840 21146
rect 872 21114 912 21146
rect 944 21114 984 21146
rect 1016 21114 1056 21146
rect 1088 21114 1128 21146
rect 1160 21114 1200 21146
rect 1232 21114 1272 21146
rect 1304 21114 1344 21146
rect 1376 21114 1416 21146
rect 1448 21114 1488 21146
rect 1520 21114 1560 21146
rect 1592 21114 1632 21146
rect 1664 21114 1704 21146
rect 1736 21114 1776 21146
rect 1808 21114 1848 21146
rect 1880 21114 1950 21146
rect 50 21074 1950 21114
rect 50 21042 120 21074
rect 152 21042 192 21074
rect 224 21042 264 21074
rect 296 21042 336 21074
rect 368 21042 408 21074
rect 440 21042 480 21074
rect 512 21042 552 21074
rect 584 21042 624 21074
rect 656 21042 696 21074
rect 728 21042 768 21074
rect 800 21042 840 21074
rect 872 21042 912 21074
rect 944 21042 984 21074
rect 1016 21042 1056 21074
rect 1088 21042 1128 21074
rect 1160 21042 1200 21074
rect 1232 21042 1272 21074
rect 1304 21042 1344 21074
rect 1376 21042 1416 21074
rect 1448 21042 1488 21074
rect 1520 21042 1560 21074
rect 1592 21042 1632 21074
rect 1664 21042 1704 21074
rect 1736 21042 1776 21074
rect 1808 21042 1848 21074
rect 1880 21042 1950 21074
rect 50 21002 1950 21042
rect 50 20970 120 21002
rect 152 20970 192 21002
rect 224 20970 264 21002
rect 296 20970 336 21002
rect 368 20970 408 21002
rect 440 20970 480 21002
rect 512 20970 552 21002
rect 584 20970 624 21002
rect 656 20970 696 21002
rect 728 20970 768 21002
rect 800 20970 840 21002
rect 872 20970 912 21002
rect 944 20970 984 21002
rect 1016 20970 1056 21002
rect 1088 20970 1128 21002
rect 1160 20970 1200 21002
rect 1232 20970 1272 21002
rect 1304 20970 1344 21002
rect 1376 20970 1416 21002
rect 1448 20970 1488 21002
rect 1520 20970 1560 21002
rect 1592 20970 1632 21002
rect 1664 20970 1704 21002
rect 1736 20970 1776 21002
rect 1808 20970 1848 21002
rect 1880 20970 1950 21002
rect 50 20930 1950 20970
rect 50 20898 120 20930
rect 152 20898 192 20930
rect 224 20898 264 20930
rect 296 20898 336 20930
rect 368 20898 408 20930
rect 440 20898 480 20930
rect 512 20898 552 20930
rect 584 20898 624 20930
rect 656 20898 696 20930
rect 728 20898 768 20930
rect 800 20898 840 20930
rect 872 20898 912 20930
rect 944 20898 984 20930
rect 1016 20898 1056 20930
rect 1088 20898 1128 20930
rect 1160 20898 1200 20930
rect 1232 20898 1272 20930
rect 1304 20898 1344 20930
rect 1376 20898 1416 20930
rect 1448 20898 1488 20930
rect 1520 20898 1560 20930
rect 1592 20898 1632 20930
rect 1664 20898 1704 20930
rect 1736 20898 1776 20930
rect 1808 20898 1848 20930
rect 1880 20898 1950 20930
rect 50 20858 1950 20898
rect 50 20826 120 20858
rect 152 20826 192 20858
rect 224 20826 264 20858
rect 296 20826 336 20858
rect 368 20826 408 20858
rect 440 20826 480 20858
rect 512 20826 552 20858
rect 584 20826 624 20858
rect 656 20826 696 20858
rect 728 20826 768 20858
rect 800 20826 840 20858
rect 872 20826 912 20858
rect 944 20826 984 20858
rect 1016 20826 1056 20858
rect 1088 20826 1128 20858
rect 1160 20826 1200 20858
rect 1232 20826 1272 20858
rect 1304 20826 1344 20858
rect 1376 20826 1416 20858
rect 1448 20826 1488 20858
rect 1520 20826 1560 20858
rect 1592 20826 1632 20858
rect 1664 20826 1704 20858
rect 1736 20826 1776 20858
rect 1808 20826 1848 20858
rect 1880 20826 1950 20858
rect 50 20786 1950 20826
rect 50 20754 120 20786
rect 152 20754 192 20786
rect 224 20754 264 20786
rect 296 20754 336 20786
rect 368 20754 408 20786
rect 440 20754 480 20786
rect 512 20754 552 20786
rect 584 20754 624 20786
rect 656 20754 696 20786
rect 728 20754 768 20786
rect 800 20754 840 20786
rect 872 20754 912 20786
rect 944 20754 984 20786
rect 1016 20754 1056 20786
rect 1088 20754 1128 20786
rect 1160 20754 1200 20786
rect 1232 20754 1272 20786
rect 1304 20754 1344 20786
rect 1376 20754 1416 20786
rect 1448 20754 1488 20786
rect 1520 20754 1560 20786
rect 1592 20754 1632 20786
rect 1664 20754 1704 20786
rect 1736 20754 1776 20786
rect 1808 20754 1848 20786
rect 1880 20754 1950 20786
rect 50 20714 1950 20754
rect 50 20682 120 20714
rect 152 20682 192 20714
rect 224 20682 264 20714
rect 296 20682 336 20714
rect 368 20682 408 20714
rect 440 20682 480 20714
rect 512 20682 552 20714
rect 584 20682 624 20714
rect 656 20682 696 20714
rect 728 20682 768 20714
rect 800 20682 840 20714
rect 872 20682 912 20714
rect 944 20682 984 20714
rect 1016 20682 1056 20714
rect 1088 20682 1128 20714
rect 1160 20682 1200 20714
rect 1232 20682 1272 20714
rect 1304 20682 1344 20714
rect 1376 20682 1416 20714
rect 1448 20682 1488 20714
rect 1520 20682 1560 20714
rect 1592 20682 1632 20714
rect 1664 20682 1704 20714
rect 1736 20682 1776 20714
rect 1808 20682 1848 20714
rect 1880 20682 1950 20714
rect 50 20642 1950 20682
rect 50 20610 120 20642
rect 152 20610 192 20642
rect 224 20610 264 20642
rect 296 20610 336 20642
rect 368 20610 408 20642
rect 440 20610 480 20642
rect 512 20610 552 20642
rect 584 20610 624 20642
rect 656 20610 696 20642
rect 728 20610 768 20642
rect 800 20610 840 20642
rect 872 20610 912 20642
rect 944 20610 984 20642
rect 1016 20610 1056 20642
rect 1088 20610 1128 20642
rect 1160 20610 1200 20642
rect 1232 20610 1272 20642
rect 1304 20610 1344 20642
rect 1376 20610 1416 20642
rect 1448 20610 1488 20642
rect 1520 20610 1560 20642
rect 1592 20610 1632 20642
rect 1664 20610 1704 20642
rect 1736 20610 1776 20642
rect 1808 20610 1848 20642
rect 1880 20610 1950 20642
rect 50 20570 1950 20610
rect 50 20538 120 20570
rect 152 20538 192 20570
rect 224 20538 264 20570
rect 296 20538 336 20570
rect 368 20538 408 20570
rect 440 20538 480 20570
rect 512 20538 552 20570
rect 584 20538 624 20570
rect 656 20538 696 20570
rect 728 20538 768 20570
rect 800 20538 840 20570
rect 872 20538 912 20570
rect 944 20538 984 20570
rect 1016 20538 1056 20570
rect 1088 20538 1128 20570
rect 1160 20538 1200 20570
rect 1232 20538 1272 20570
rect 1304 20538 1344 20570
rect 1376 20538 1416 20570
rect 1448 20538 1488 20570
rect 1520 20538 1560 20570
rect 1592 20538 1632 20570
rect 1664 20538 1704 20570
rect 1736 20538 1776 20570
rect 1808 20538 1848 20570
rect 1880 20538 1950 20570
rect 50 20498 1950 20538
rect 50 20466 120 20498
rect 152 20466 192 20498
rect 224 20466 264 20498
rect 296 20466 336 20498
rect 368 20466 408 20498
rect 440 20466 480 20498
rect 512 20466 552 20498
rect 584 20466 624 20498
rect 656 20466 696 20498
rect 728 20466 768 20498
rect 800 20466 840 20498
rect 872 20466 912 20498
rect 944 20466 984 20498
rect 1016 20466 1056 20498
rect 1088 20466 1128 20498
rect 1160 20466 1200 20498
rect 1232 20466 1272 20498
rect 1304 20466 1344 20498
rect 1376 20466 1416 20498
rect 1448 20466 1488 20498
rect 1520 20466 1560 20498
rect 1592 20466 1632 20498
rect 1664 20466 1704 20498
rect 1736 20466 1776 20498
rect 1808 20466 1848 20498
rect 1880 20466 1950 20498
rect 50 20426 1950 20466
rect 50 20394 120 20426
rect 152 20394 192 20426
rect 224 20394 264 20426
rect 296 20394 336 20426
rect 368 20394 408 20426
rect 440 20394 480 20426
rect 512 20394 552 20426
rect 584 20394 624 20426
rect 656 20394 696 20426
rect 728 20394 768 20426
rect 800 20394 840 20426
rect 872 20394 912 20426
rect 944 20394 984 20426
rect 1016 20394 1056 20426
rect 1088 20394 1128 20426
rect 1160 20394 1200 20426
rect 1232 20394 1272 20426
rect 1304 20394 1344 20426
rect 1376 20394 1416 20426
rect 1448 20394 1488 20426
rect 1520 20394 1560 20426
rect 1592 20394 1632 20426
rect 1664 20394 1704 20426
rect 1736 20394 1776 20426
rect 1808 20394 1848 20426
rect 1880 20394 1950 20426
rect 50 20354 1950 20394
rect 50 20322 120 20354
rect 152 20322 192 20354
rect 224 20322 264 20354
rect 296 20322 336 20354
rect 368 20322 408 20354
rect 440 20322 480 20354
rect 512 20322 552 20354
rect 584 20322 624 20354
rect 656 20322 696 20354
rect 728 20322 768 20354
rect 800 20322 840 20354
rect 872 20322 912 20354
rect 944 20322 984 20354
rect 1016 20322 1056 20354
rect 1088 20322 1128 20354
rect 1160 20322 1200 20354
rect 1232 20322 1272 20354
rect 1304 20322 1344 20354
rect 1376 20322 1416 20354
rect 1448 20322 1488 20354
rect 1520 20322 1560 20354
rect 1592 20322 1632 20354
rect 1664 20322 1704 20354
rect 1736 20322 1776 20354
rect 1808 20322 1848 20354
rect 1880 20322 1950 20354
rect 50 20282 1950 20322
rect 50 20250 120 20282
rect 152 20250 192 20282
rect 224 20250 264 20282
rect 296 20250 336 20282
rect 368 20250 408 20282
rect 440 20250 480 20282
rect 512 20250 552 20282
rect 584 20250 624 20282
rect 656 20250 696 20282
rect 728 20250 768 20282
rect 800 20250 840 20282
rect 872 20250 912 20282
rect 944 20250 984 20282
rect 1016 20250 1056 20282
rect 1088 20250 1128 20282
rect 1160 20250 1200 20282
rect 1232 20250 1272 20282
rect 1304 20250 1344 20282
rect 1376 20250 1416 20282
rect 1448 20250 1488 20282
rect 1520 20250 1560 20282
rect 1592 20250 1632 20282
rect 1664 20250 1704 20282
rect 1736 20250 1776 20282
rect 1808 20250 1848 20282
rect 1880 20250 1950 20282
rect 50 20210 1950 20250
rect 50 20178 120 20210
rect 152 20178 192 20210
rect 224 20178 264 20210
rect 296 20178 336 20210
rect 368 20178 408 20210
rect 440 20178 480 20210
rect 512 20178 552 20210
rect 584 20178 624 20210
rect 656 20178 696 20210
rect 728 20178 768 20210
rect 800 20178 840 20210
rect 872 20178 912 20210
rect 944 20178 984 20210
rect 1016 20178 1056 20210
rect 1088 20178 1128 20210
rect 1160 20178 1200 20210
rect 1232 20178 1272 20210
rect 1304 20178 1344 20210
rect 1376 20178 1416 20210
rect 1448 20178 1488 20210
rect 1520 20178 1560 20210
rect 1592 20178 1632 20210
rect 1664 20178 1704 20210
rect 1736 20178 1776 20210
rect 1808 20178 1848 20210
rect 1880 20178 1950 20210
rect 50 20138 1950 20178
rect 50 20106 120 20138
rect 152 20106 192 20138
rect 224 20106 264 20138
rect 296 20106 336 20138
rect 368 20106 408 20138
rect 440 20106 480 20138
rect 512 20106 552 20138
rect 584 20106 624 20138
rect 656 20106 696 20138
rect 728 20106 768 20138
rect 800 20106 840 20138
rect 872 20106 912 20138
rect 944 20106 984 20138
rect 1016 20106 1056 20138
rect 1088 20106 1128 20138
rect 1160 20106 1200 20138
rect 1232 20106 1272 20138
rect 1304 20106 1344 20138
rect 1376 20106 1416 20138
rect 1448 20106 1488 20138
rect 1520 20106 1560 20138
rect 1592 20106 1632 20138
rect 1664 20106 1704 20138
rect 1736 20106 1776 20138
rect 1808 20106 1848 20138
rect 1880 20106 1950 20138
rect 50 20066 1950 20106
rect 50 20034 120 20066
rect 152 20034 192 20066
rect 224 20034 264 20066
rect 296 20034 336 20066
rect 368 20034 408 20066
rect 440 20034 480 20066
rect 512 20034 552 20066
rect 584 20034 624 20066
rect 656 20034 696 20066
rect 728 20034 768 20066
rect 800 20034 840 20066
rect 872 20034 912 20066
rect 944 20034 984 20066
rect 1016 20034 1056 20066
rect 1088 20034 1128 20066
rect 1160 20034 1200 20066
rect 1232 20034 1272 20066
rect 1304 20034 1344 20066
rect 1376 20034 1416 20066
rect 1448 20034 1488 20066
rect 1520 20034 1560 20066
rect 1592 20034 1632 20066
rect 1664 20034 1704 20066
rect 1736 20034 1776 20066
rect 1808 20034 1848 20066
rect 1880 20034 1950 20066
rect 50 19994 1950 20034
rect 50 19962 120 19994
rect 152 19962 192 19994
rect 224 19962 264 19994
rect 296 19962 336 19994
rect 368 19962 408 19994
rect 440 19962 480 19994
rect 512 19962 552 19994
rect 584 19962 624 19994
rect 656 19962 696 19994
rect 728 19962 768 19994
rect 800 19962 840 19994
rect 872 19962 912 19994
rect 944 19962 984 19994
rect 1016 19962 1056 19994
rect 1088 19962 1128 19994
rect 1160 19962 1200 19994
rect 1232 19962 1272 19994
rect 1304 19962 1344 19994
rect 1376 19962 1416 19994
rect 1448 19962 1488 19994
rect 1520 19962 1560 19994
rect 1592 19962 1632 19994
rect 1664 19962 1704 19994
rect 1736 19962 1776 19994
rect 1808 19962 1848 19994
rect 1880 19962 1950 19994
rect 50 19922 1950 19962
rect 50 19890 120 19922
rect 152 19890 192 19922
rect 224 19890 264 19922
rect 296 19890 336 19922
rect 368 19890 408 19922
rect 440 19890 480 19922
rect 512 19890 552 19922
rect 584 19890 624 19922
rect 656 19890 696 19922
rect 728 19890 768 19922
rect 800 19890 840 19922
rect 872 19890 912 19922
rect 944 19890 984 19922
rect 1016 19890 1056 19922
rect 1088 19890 1128 19922
rect 1160 19890 1200 19922
rect 1232 19890 1272 19922
rect 1304 19890 1344 19922
rect 1376 19890 1416 19922
rect 1448 19890 1488 19922
rect 1520 19890 1560 19922
rect 1592 19890 1632 19922
rect 1664 19890 1704 19922
rect 1736 19890 1776 19922
rect 1808 19890 1848 19922
rect 1880 19890 1950 19922
rect 50 19850 1950 19890
rect 50 19818 120 19850
rect 152 19818 192 19850
rect 224 19818 264 19850
rect 296 19818 336 19850
rect 368 19818 408 19850
rect 440 19818 480 19850
rect 512 19818 552 19850
rect 584 19818 624 19850
rect 656 19818 696 19850
rect 728 19818 768 19850
rect 800 19818 840 19850
rect 872 19818 912 19850
rect 944 19818 984 19850
rect 1016 19818 1056 19850
rect 1088 19818 1128 19850
rect 1160 19818 1200 19850
rect 1232 19818 1272 19850
rect 1304 19818 1344 19850
rect 1376 19818 1416 19850
rect 1448 19818 1488 19850
rect 1520 19818 1560 19850
rect 1592 19818 1632 19850
rect 1664 19818 1704 19850
rect 1736 19818 1776 19850
rect 1808 19818 1848 19850
rect 1880 19818 1950 19850
rect 50 19778 1950 19818
rect 50 19746 120 19778
rect 152 19746 192 19778
rect 224 19746 264 19778
rect 296 19746 336 19778
rect 368 19746 408 19778
rect 440 19746 480 19778
rect 512 19746 552 19778
rect 584 19746 624 19778
rect 656 19746 696 19778
rect 728 19746 768 19778
rect 800 19746 840 19778
rect 872 19746 912 19778
rect 944 19746 984 19778
rect 1016 19746 1056 19778
rect 1088 19746 1128 19778
rect 1160 19746 1200 19778
rect 1232 19746 1272 19778
rect 1304 19746 1344 19778
rect 1376 19746 1416 19778
rect 1448 19746 1488 19778
rect 1520 19746 1560 19778
rect 1592 19746 1632 19778
rect 1664 19746 1704 19778
rect 1736 19746 1776 19778
rect 1808 19746 1848 19778
rect 1880 19746 1950 19778
rect 50 19706 1950 19746
rect 50 19674 120 19706
rect 152 19674 192 19706
rect 224 19674 264 19706
rect 296 19674 336 19706
rect 368 19674 408 19706
rect 440 19674 480 19706
rect 512 19674 552 19706
rect 584 19674 624 19706
rect 656 19674 696 19706
rect 728 19674 768 19706
rect 800 19674 840 19706
rect 872 19674 912 19706
rect 944 19674 984 19706
rect 1016 19674 1056 19706
rect 1088 19674 1128 19706
rect 1160 19674 1200 19706
rect 1232 19674 1272 19706
rect 1304 19674 1344 19706
rect 1376 19674 1416 19706
rect 1448 19674 1488 19706
rect 1520 19674 1560 19706
rect 1592 19674 1632 19706
rect 1664 19674 1704 19706
rect 1736 19674 1776 19706
rect 1808 19674 1848 19706
rect 1880 19674 1950 19706
rect 50 19634 1950 19674
rect 50 19602 120 19634
rect 152 19602 192 19634
rect 224 19602 264 19634
rect 296 19602 336 19634
rect 368 19602 408 19634
rect 440 19602 480 19634
rect 512 19602 552 19634
rect 584 19602 624 19634
rect 656 19602 696 19634
rect 728 19602 768 19634
rect 800 19602 840 19634
rect 872 19602 912 19634
rect 944 19602 984 19634
rect 1016 19602 1056 19634
rect 1088 19602 1128 19634
rect 1160 19602 1200 19634
rect 1232 19602 1272 19634
rect 1304 19602 1344 19634
rect 1376 19602 1416 19634
rect 1448 19602 1488 19634
rect 1520 19602 1560 19634
rect 1592 19602 1632 19634
rect 1664 19602 1704 19634
rect 1736 19602 1776 19634
rect 1808 19602 1848 19634
rect 1880 19602 1950 19634
rect 50 19562 1950 19602
rect 50 19530 120 19562
rect 152 19530 192 19562
rect 224 19530 264 19562
rect 296 19530 336 19562
rect 368 19530 408 19562
rect 440 19530 480 19562
rect 512 19530 552 19562
rect 584 19530 624 19562
rect 656 19530 696 19562
rect 728 19530 768 19562
rect 800 19530 840 19562
rect 872 19530 912 19562
rect 944 19530 984 19562
rect 1016 19530 1056 19562
rect 1088 19530 1128 19562
rect 1160 19530 1200 19562
rect 1232 19530 1272 19562
rect 1304 19530 1344 19562
rect 1376 19530 1416 19562
rect 1448 19530 1488 19562
rect 1520 19530 1560 19562
rect 1592 19530 1632 19562
rect 1664 19530 1704 19562
rect 1736 19530 1776 19562
rect 1808 19530 1848 19562
rect 1880 19530 1950 19562
rect 50 19490 1950 19530
rect 50 19458 120 19490
rect 152 19458 192 19490
rect 224 19458 264 19490
rect 296 19458 336 19490
rect 368 19458 408 19490
rect 440 19458 480 19490
rect 512 19458 552 19490
rect 584 19458 624 19490
rect 656 19458 696 19490
rect 728 19458 768 19490
rect 800 19458 840 19490
rect 872 19458 912 19490
rect 944 19458 984 19490
rect 1016 19458 1056 19490
rect 1088 19458 1128 19490
rect 1160 19458 1200 19490
rect 1232 19458 1272 19490
rect 1304 19458 1344 19490
rect 1376 19458 1416 19490
rect 1448 19458 1488 19490
rect 1520 19458 1560 19490
rect 1592 19458 1632 19490
rect 1664 19458 1704 19490
rect 1736 19458 1776 19490
rect 1808 19458 1848 19490
rect 1880 19458 1950 19490
rect 50 19418 1950 19458
rect 50 19386 120 19418
rect 152 19386 192 19418
rect 224 19386 264 19418
rect 296 19386 336 19418
rect 368 19386 408 19418
rect 440 19386 480 19418
rect 512 19386 552 19418
rect 584 19386 624 19418
rect 656 19386 696 19418
rect 728 19386 768 19418
rect 800 19386 840 19418
rect 872 19386 912 19418
rect 944 19386 984 19418
rect 1016 19386 1056 19418
rect 1088 19386 1128 19418
rect 1160 19386 1200 19418
rect 1232 19386 1272 19418
rect 1304 19386 1344 19418
rect 1376 19386 1416 19418
rect 1448 19386 1488 19418
rect 1520 19386 1560 19418
rect 1592 19386 1632 19418
rect 1664 19386 1704 19418
rect 1736 19386 1776 19418
rect 1808 19386 1848 19418
rect 1880 19386 1950 19418
rect 50 19346 1950 19386
rect 50 19314 120 19346
rect 152 19314 192 19346
rect 224 19314 264 19346
rect 296 19314 336 19346
rect 368 19314 408 19346
rect 440 19314 480 19346
rect 512 19314 552 19346
rect 584 19314 624 19346
rect 656 19314 696 19346
rect 728 19314 768 19346
rect 800 19314 840 19346
rect 872 19314 912 19346
rect 944 19314 984 19346
rect 1016 19314 1056 19346
rect 1088 19314 1128 19346
rect 1160 19314 1200 19346
rect 1232 19314 1272 19346
rect 1304 19314 1344 19346
rect 1376 19314 1416 19346
rect 1448 19314 1488 19346
rect 1520 19314 1560 19346
rect 1592 19314 1632 19346
rect 1664 19314 1704 19346
rect 1736 19314 1776 19346
rect 1808 19314 1848 19346
rect 1880 19314 1950 19346
rect 50 19274 1950 19314
rect 50 19242 120 19274
rect 152 19242 192 19274
rect 224 19242 264 19274
rect 296 19242 336 19274
rect 368 19242 408 19274
rect 440 19242 480 19274
rect 512 19242 552 19274
rect 584 19242 624 19274
rect 656 19242 696 19274
rect 728 19242 768 19274
rect 800 19242 840 19274
rect 872 19242 912 19274
rect 944 19242 984 19274
rect 1016 19242 1056 19274
rect 1088 19242 1128 19274
rect 1160 19242 1200 19274
rect 1232 19242 1272 19274
rect 1304 19242 1344 19274
rect 1376 19242 1416 19274
rect 1448 19242 1488 19274
rect 1520 19242 1560 19274
rect 1592 19242 1632 19274
rect 1664 19242 1704 19274
rect 1736 19242 1776 19274
rect 1808 19242 1848 19274
rect 1880 19242 1950 19274
rect 50 19202 1950 19242
rect 50 19170 120 19202
rect 152 19170 192 19202
rect 224 19170 264 19202
rect 296 19170 336 19202
rect 368 19170 408 19202
rect 440 19170 480 19202
rect 512 19170 552 19202
rect 584 19170 624 19202
rect 656 19170 696 19202
rect 728 19170 768 19202
rect 800 19170 840 19202
rect 872 19170 912 19202
rect 944 19170 984 19202
rect 1016 19170 1056 19202
rect 1088 19170 1128 19202
rect 1160 19170 1200 19202
rect 1232 19170 1272 19202
rect 1304 19170 1344 19202
rect 1376 19170 1416 19202
rect 1448 19170 1488 19202
rect 1520 19170 1560 19202
rect 1592 19170 1632 19202
rect 1664 19170 1704 19202
rect 1736 19170 1776 19202
rect 1808 19170 1848 19202
rect 1880 19170 1950 19202
rect 50 19130 1950 19170
rect 50 19098 120 19130
rect 152 19098 192 19130
rect 224 19098 264 19130
rect 296 19098 336 19130
rect 368 19098 408 19130
rect 440 19098 480 19130
rect 512 19098 552 19130
rect 584 19098 624 19130
rect 656 19098 696 19130
rect 728 19098 768 19130
rect 800 19098 840 19130
rect 872 19098 912 19130
rect 944 19098 984 19130
rect 1016 19098 1056 19130
rect 1088 19098 1128 19130
rect 1160 19098 1200 19130
rect 1232 19098 1272 19130
rect 1304 19098 1344 19130
rect 1376 19098 1416 19130
rect 1448 19098 1488 19130
rect 1520 19098 1560 19130
rect 1592 19098 1632 19130
rect 1664 19098 1704 19130
rect 1736 19098 1776 19130
rect 1808 19098 1848 19130
rect 1880 19098 1950 19130
rect 50 19058 1950 19098
rect 50 19026 120 19058
rect 152 19026 192 19058
rect 224 19026 264 19058
rect 296 19026 336 19058
rect 368 19026 408 19058
rect 440 19026 480 19058
rect 512 19026 552 19058
rect 584 19026 624 19058
rect 656 19026 696 19058
rect 728 19026 768 19058
rect 800 19026 840 19058
rect 872 19026 912 19058
rect 944 19026 984 19058
rect 1016 19026 1056 19058
rect 1088 19026 1128 19058
rect 1160 19026 1200 19058
rect 1232 19026 1272 19058
rect 1304 19026 1344 19058
rect 1376 19026 1416 19058
rect 1448 19026 1488 19058
rect 1520 19026 1560 19058
rect 1592 19026 1632 19058
rect 1664 19026 1704 19058
rect 1736 19026 1776 19058
rect 1808 19026 1848 19058
rect 1880 19026 1950 19058
rect 50 18986 1950 19026
rect 50 18954 120 18986
rect 152 18954 192 18986
rect 224 18954 264 18986
rect 296 18954 336 18986
rect 368 18954 408 18986
rect 440 18954 480 18986
rect 512 18954 552 18986
rect 584 18954 624 18986
rect 656 18954 696 18986
rect 728 18954 768 18986
rect 800 18954 840 18986
rect 872 18954 912 18986
rect 944 18954 984 18986
rect 1016 18954 1056 18986
rect 1088 18954 1128 18986
rect 1160 18954 1200 18986
rect 1232 18954 1272 18986
rect 1304 18954 1344 18986
rect 1376 18954 1416 18986
rect 1448 18954 1488 18986
rect 1520 18954 1560 18986
rect 1592 18954 1632 18986
rect 1664 18954 1704 18986
rect 1736 18954 1776 18986
rect 1808 18954 1848 18986
rect 1880 18954 1950 18986
rect 50 18914 1950 18954
rect 50 18882 120 18914
rect 152 18882 192 18914
rect 224 18882 264 18914
rect 296 18882 336 18914
rect 368 18882 408 18914
rect 440 18882 480 18914
rect 512 18882 552 18914
rect 584 18882 624 18914
rect 656 18882 696 18914
rect 728 18882 768 18914
rect 800 18882 840 18914
rect 872 18882 912 18914
rect 944 18882 984 18914
rect 1016 18882 1056 18914
rect 1088 18882 1128 18914
rect 1160 18882 1200 18914
rect 1232 18882 1272 18914
rect 1304 18882 1344 18914
rect 1376 18882 1416 18914
rect 1448 18882 1488 18914
rect 1520 18882 1560 18914
rect 1592 18882 1632 18914
rect 1664 18882 1704 18914
rect 1736 18882 1776 18914
rect 1808 18882 1848 18914
rect 1880 18882 1950 18914
rect 50 18842 1950 18882
rect 50 18810 120 18842
rect 152 18810 192 18842
rect 224 18810 264 18842
rect 296 18810 336 18842
rect 368 18810 408 18842
rect 440 18810 480 18842
rect 512 18810 552 18842
rect 584 18810 624 18842
rect 656 18810 696 18842
rect 728 18810 768 18842
rect 800 18810 840 18842
rect 872 18810 912 18842
rect 944 18810 984 18842
rect 1016 18810 1056 18842
rect 1088 18810 1128 18842
rect 1160 18810 1200 18842
rect 1232 18810 1272 18842
rect 1304 18810 1344 18842
rect 1376 18810 1416 18842
rect 1448 18810 1488 18842
rect 1520 18810 1560 18842
rect 1592 18810 1632 18842
rect 1664 18810 1704 18842
rect 1736 18810 1776 18842
rect 1808 18810 1848 18842
rect 1880 18810 1950 18842
rect 50 18770 1950 18810
rect 50 18738 120 18770
rect 152 18738 192 18770
rect 224 18738 264 18770
rect 296 18738 336 18770
rect 368 18738 408 18770
rect 440 18738 480 18770
rect 512 18738 552 18770
rect 584 18738 624 18770
rect 656 18738 696 18770
rect 728 18738 768 18770
rect 800 18738 840 18770
rect 872 18738 912 18770
rect 944 18738 984 18770
rect 1016 18738 1056 18770
rect 1088 18738 1128 18770
rect 1160 18738 1200 18770
rect 1232 18738 1272 18770
rect 1304 18738 1344 18770
rect 1376 18738 1416 18770
rect 1448 18738 1488 18770
rect 1520 18738 1560 18770
rect 1592 18738 1632 18770
rect 1664 18738 1704 18770
rect 1736 18738 1776 18770
rect 1808 18738 1848 18770
rect 1880 18738 1950 18770
rect 50 18698 1950 18738
rect 50 18666 120 18698
rect 152 18666 192 18698
rect 224 18666 264 18698
rect 296 18666 336 18698
rect 368 18666 408 18698
rect 440 18666 480 18698
rect 512 18666 552 18698
rect 584 18666 624 18698
rect 656 18666 696 18698
rect 728 18666 768 18698
rect 800 18666 840 18698
rect 872 18666 912 18698
rect 944 18666 984 18698
rect 1016 18666 1056 18698
rect 1088 18666 1128 18698
rect 1160 18666 1200 18698
rect 1232 18666 1272 18698
rect 1304 18666 1344 18698
rect 1376 18666 1416 18698
rect 1448 18666 1488 18698
rect 1520 18666 1560 18698
rect 1592 18666 1632 18698
rect 1664 18666 1704 18698
rect 1736 18666 1776 18698
rect 1808 18666 1848 18698
rect 1880 18666 1950 18698
rect 50 18626 1950 18666
rect 50 18594 120 18626
rect 152 18594 192 18626
rect 224 18594 264 18626
rect 296 18594 336 18626
rect 368 18594 408 18626
rect 440 18594 480 18626
rect 512 18594 552 18626
rect 584 18594 624 18626
rect 656 18594 696 18626
rect 728 18594 768 18626
rect 800 18594 840 18626
rect 872 18594 912 18626
rect 944 18594 984 18626
rect 1016 18594 1056 18626
rect 1088 18594 1128 18626
rect 1160 18594 1200 18626
rect 1232 18594 1272 18626
rect 1304 18594 1344 18626
rect 1376 18594 1416 18626
rect 1448 18594 1488 18626
rect 1520 18594 1560 18626
rect 1592 18594 1632 18626
rect 1664 18594 1704 18626
rect 1736 18594 1776 18626
rect 1808 18594 1848 18626
rect 1880 18594 1950 18626
rect 50 18554 1950 18594
rect 50 18522 120 18554
rect 152 18522 192 18554
rect 224 18522 264 18554
rect 296 18522 336 18554
rect 368 18522 408 18554
rect 440 18522 480 18554
rect 512 18522 552 18554
rect 584 18522 624 18554
rect 656 18522 696 18554
rect 728 18522 768 18554
rect 800 18522 840 18554
rect 872 18522 912 18554
rect 944 18522 984 18554
rect 1016 18522 1056 18554
rect 1088 18522 1128 18554
rect 1160 18522 1200 18554
rect 1232 18522 1272 18554
rect 1304 18522 1344 18554
rect 1376 18522 1416 18554
rect 1448 18522 1488 18554
rect 1520 18522 1560 18554
rect 1592 18522 1632 18554
rect 1664 18522 1704 18554
rect 1736 18522 1776 18554
rect 1808 18522 1848 18554
rect 1880 18522 1950 18554
rect 50 18482 1950 18522
rect 50 18450 120 18482
rect 152 18450 192 18482
rect 224 18450 264 18482
rect 296 18450 336 18482
rect 368 18450 408 18482
rect 440 18450 480 18482
rect 512 18450 552 18482
rect 584 18450 624 18482
rect 656 18450 696 18482
rect 728 18450 768 18482
rect 800 18450 840 18482
rect 872 18450 912 18482
rect 944 18450 984 18482
rect 1016 18450 1056 18482
rect 1088 18450 1128 18482
rect 1160 18450 1200 18482
rect 1232 18450 1272 18482
rect 1304 18450 1344 18482
rect 1376 18450 1416 18482
rect 1448 18450 1488 18482
rect 1520 18450 1560 18482
rect 1592 18450 1632 18482
rect 1664 18450 1704 18482
rect 1736 18450 1776 18482
rect 1808 18450 1848 18482
rect 1880 18450 1950 18482
rect 50 18410 1950 18450
rect 50 18378 120 18410
rect 152 18378 192 18410
rect 224 18378 264 18410
rect 296 18378 336 18410
rect 368 18378 408 18410
rect 440 18378 480 18410
rect 512 18378 552 18410
rect 584 18378 624 18410
rect 656 18378 696 18410
rect 728 18378 768 18410
rect 800 18378 840 18410
rect 872 18378 912 18410
rect 944 18378 984 18410
rect 1016 18378 1056 18410
rect 1088 18378 1128 18410
rect 1160 18378 1200 18410
rect 1232 18378 1272 18410
rect 1304 18378 1344 18410
rect 1376 18378 1416 18410
rect 1448 18378 1488 18410
rect 1520 18378 1560 18410
rect 1592 18378 1632 18410
rect 1664 18378 1704 18410
rect 1736 18378 1776 18410
rect 1808 18378 1848 18410
rect 1880 18378 1950 18410
rect 50 18338 1950 18378
rect 50 18306 120 18338
rect 152 18306 192 18338
rect 224 18306 264 18338
rect 296 18306 336 18338
rect 368 18306 408 18338
rect 440 18306 480 18338
rect 512 18306 552 18338
rect 584 18306 624 18338
rect 656 18306 696 18338
rect 728 18306 768 18338
rect 800 18306 840 18338
rect 872 18306 912 18338
rect 944 18306 984 18338
rect 1016 18306 1056 18338
rect 1088 18306 1128 18338
rect 1160 18306 1200 18338
rect 1232 18306 1272 18338
rect 1304 18306 1344 18338
rect 1376 18306 1416 18338
rect 1448 18306 1488 18338
rect 1520 18306 1560 18338
rect 1592 18306 1632 18338
rect 1664 18306 1704 18338
rect 1736 18306 1776 18338
rect 1808 18306 1848 18338
rect 1880 18306 1950 18338
rect 50 18266 1950 18306
rect 50 18234 120 18266
rect 152 18234 192 18266
rect 224 18234 264 18266
rect 296 18234 336 18266
rect 368 18234 408 18266
rect 440 18234 480 18266
rect 512 18234 552 18266
rect 584 18234 624 18266
rect 656 18234 696 18266
rect 728 18234 768 18266
rect 800 18234 840 18266
rect 872 18234 912 18266
rect 944 18234 984 18266
rect 1016 18234 1056 18266
rect 1088 18234 1128 18266
rect 1160 18234 1200 18266
rect 1232 18234 1272 18266
rect 1304 18234 1344 18266
rect 1376 18234 1416 18266
rect 1448 18234 1488 18266
rect 1520 18234 1560 18266
rect 1592 18234 1632 18266
rect 1664 18234 1704 18266
rect 1736 18234 1776 18266
rect 1808 18234 1848 18266
rect 1880 18234 1950 18266
rect 50 18194 1950 18234
rect 50 18162 120 18194
rect 152 18162 192 18194
rect 224 18162 264 18194
rect 296 18162 336 18194
rect 368 18162 408 18194
rect 440 18162 480 18194
rect 512 18162 552 18194
rect 584 18162 624 18194
rect 656 18162 696 18194
rect 728 18162 768 18194
rect 800 18162 840 18194
rect 872 18162 912 18194
rect 944 18162 984 18194
rect 1016 18162 1056 18194
rect 1088 18162 1128 18194
rect 1160 18162 1200 18194
rect 1232 18162 1272 18194
rect 1304 18162 1344 18194
rect 1376 18162 1416 18194
rect 1448 18162 1488 18194
rect 1520 18162 1560 18194
rect 1592 18162 1632 18194
rect 1664 18162 1704 18194
rect 1736 18162 1776 18194
rect 1808 18162 1848 18194
rect 1880 18162 1950 18194
rect 50 18112 1950 18162
rect 50 17848 1950 17912
rect 50 17816 120 17848
rect 152 17816 192 17848
rect 224 17816 264 17848
rect 296 17816 336 17848
rect 368 17816 408 17848
rect 440 17816 480 17848
rect 512 17816 552 17848
rect 584 17816 624 17848
rect 656 17816 696 17848
rect 728 17816 768 17848
rect 800 17816 840 17848
rect 872 17816 912 17848
rect 944 17816 984 17848
rect 1016 17816 1056 17848
rect 1088 17816 1128 17848
rect 1160 17816 1200 17848
rect 1232 17816 1272 17848
rect 1304 17816 1344 17848
rect 1376 17816 1416 17848
rect 1448 17816 1488 17848
rect 1520 17816 1560 17848
rect 1592 17816 1632 17848
rect 1664 17816 1704 17848
rect 1736 17816 1776 17848
rect 1808 17816 1848 17848
rect 1880 17816 1950 17848
rect 50 17776 1950 17816
rect 50 17744 120 17776
rect 152 17744 192 17776
rect 224 17744 264 17776
rect 296 17744 336 17776
rect 368 17744 408 17776
rect 440 17744 480 17776
rect 512 17744 552 17776
rect 584 17744 624 17776
rect 656 17744 696 17776
rect 728 17744 768 17776
rect 800 17744 840 17776
rect 872 17744 912 17776
rect 944 17744 984 17776
rect 1016 17744 1056 17776
rect 1088 17744 1128 17776
rect 1160 17744 1200 17776
rect 1232 17744 1272 17776
rect 1304 17744 1344 17776
rect 1376 17744 1416 17776
rect 1448 17744 1488 17776
rect 1520 17744 1560 17776
rect 1592 17744 1632 17776
rect 1664 17744 1704 17776
rect 1736 17744 1776 17776
rect 1808 17744 1848 17776
rect 1880 17744 1950 17776
rect 50 17704 1950 17744
rect 50 17672 120 17704
rect 152 17672 192 17704
rect 224 17672 264 17704
rect 296 17672 336 17704
rect 368 17672 408 17704
rect 440 17672 480 17704
rect 512 17672 552 17704
rect 584 17672 624 17704
rect 656 17672 696 17704
rect 728 17672 768 17704
rect 800 17672 840 17704
rect 872 17672 912 17704
rect 944 17672 984 17704
rect 1016 17672 1056 17704
rect 1088 17672 1128 17704
rect 1160 17672 1200 17704
rect 1232 17672 1272 17704
rect 1304 17672 1344 17704
rect 1376 17672 1416 17704
rect 1448 17672 1488 17704
rect 1520 17672 1560 17704
rect 1592 17672 1632 17704
rect 1664 17672 1704 17704
rect 1736 17672 1776 17704
rect 1808 17672 1848 17704
rect 1880 17672 1950 17704
rect 50 17632 1950 17672
rect 50 17600 120 17632
rect 152 17600 192 17632
rect 224 17600 264 17632
rect 296 17600 336 17632
rect 368 17600 408 17632
rect 440 17600 480 17632
rect 512 17600 552 17632
rect 584 17600 624 17632
rect 656 17600 696 17632
rect 728 17600 768 17632
rect 800 17600 840 17632
rect 872 17600 912 17632
rect 944 17600 984 17632
rect 1016 17600 1056 17632
rect 1088 17600 1128 17632
rect 1160 17600 1200 17632
rect 1232 17600 1272 17632
rect 1304 17600 1344 17632
rect 1376 17600 1416 17632
rect 1448 17600 1488 17632
rect 1520 17600 1560 17632
rect 1592 17600 1632 17632
rect 1664 17600 1704 17632
rect 1736 17600 1776 17632
rect 1808 17600 1848 17632
rect 1880 17600 1950 17632
rect 50 17560 1950 17600
rect 50 17528 120 17560
rect 152 17528 192 17560
rect 224 17528 264 17560
rect 296 17528 336 17560
rect 368 17528 408 17560
rect 440 17528 480 17560
rect 512 17528 552 17560
rect 584 17528 624 17560
rect 656 17528 696 17560
rect 728 17528 768 17560
rect 800 17528 840 17560
rect 872 17528 912 17560
rect 944 17528 984 17560
rect 1016 17528 1056 17560
rect 1088 17528 1128 17560
rect 1160 17528 1200 17560
rect 1232 17528 1272 17560
rect 1304 17528 1344 17560
rect 1376 17528 1416 17560
rect 1448 17528 1488 17560
rect 1520 17528 1560 17560
rect 1592 17528 1632 17560
rect 1664 17528 1704 17560
rect 1736 17528 1776 17560
rect 1808 17528 1848 17560
rect 1880 17528 1950 17560
rect 50 17488 1950 17528
rect 50 17456 120 17488
rect 152 17456 192 17488
rect 224 17456 264 17488
rect 296 17456 336 17488
rect 368 17456 408 17488
rect 440 17456 480 17488
rect 512 17456 552 17488
rect 584 17456 624 17488
rect 656 17456 696 17488
rect 728 17456 768 17488
rect 800 17456 840 17488
rect 872 17456 912 17488
rect 944 17456 984 17488
rect 1016 17456 1056 17488
rect 1088 17456 1128 17488
rect 1160 17456 1200 17488
rect 1232 17456 1272 17488
rect 1304 17456 1344 17488
rect 1376 17456 1416 17488
rect 1448 17456 1488 17488
rect 1520 17456 1560 17488
rect 1592 17456 1632 17488
rect 1664 17456 1704 17488
rect 1736 17456 1776 17488
rect 1808 17456 1848 17488
rect 1880 17456 1950 17488
rect 50 17416 1950 17456
rect 50 17384 120 17416
rect 152 17384 192 17416
rect 224 17384 264 17416
rect 296 17384 336 17416
rect 368 17384 408 17416
rect 440 17384 480 17416
rect 512 17384 552 17416
rect 584 17384 624 17416
rect 656 17384 696 17416
rect 728 17384 768 17416
rect 800 17384 840 17416
rect 872 17384 912 17416
rect 944 17384 984 17416
rect 1016 17384 1056 17416
rect 1088 17384 1128 17416
rect 1160 17384 1200 17416
rect 1232 17384 1272 17416
rect 1304 17384 1344 17416
rect 1376 17384 1416 17416
rect 1448 17384 1488 17416
rect 1520 17384 1560 17416
rect 1592 17384 1632 17416
rect 1664 17384 1704 17416
rect 1736 17384 1776 17416
rect 1808 17384 1848 17416
rect 1880 17384 1950 17416
rect 50 17344 1950 17384
rect 50 17312 120 17344
rect 152 17312 192 17344
rect 224 17312 264 17344
rect 296 17312 336 17344
rect 368 17312 408 17344
rect 440 17312 480 17344
rect 512 17312 552 17344
rect 584 17312 624 17344
rect 656 17312 696 17344
rect 728 17312 768 17344
rect 800 17312 840 17344
rect 872 17312 912 17344
rect 944 17312 984 17344
rect 1016 17312 1056 17344
rect 1088 17312 1128 17344
rect 1160 17312 1200 17344
rect 1232 17312 1272 17344
rect 1304 17312 1344 17344
rect 1376 17312 1416 17344
rect 1448 17312 1488 17344
rect 1520 17312 1560 17344
rect 1592 17312 1632 17344
rect 1664 17312 1704 17344
rect 1736 17312 1776 17344
rect 1808 17312 1848 17344
rect 1880 17312 1950 17344
rect 50 17272 1950 17312
rect 50 17240 120 17272
rect 152 17240 192 17272
rect 224 17240 264 17272
rect 296 17240 336 17272
rect 368 17240 408 17272
rect 440 17240 480 17272
rect 512 17240 552 17272
rect 584 17240 624 17272
rect 656 17240 696 17272
rect 728 17240 768 17272
rect 800 17240 840 17272
rect 872 17240 912 17272
rect 944 17240 984 17272
rect 1016 17240 1056 17272
rect 1088 17240 1128 17272
rect 1160 17240 1200 17272
rect 1232 17240 1272 17272
rect 1304 17240 1344 17272
rect 1376 17240 1416 17272
rect 1448 17240 1488 17272
rect 1520 17240 1560 17272
rect 1592 17240 1632 17272
rect 1664 17240 1704 17272
rect 1736 17240 1776 17272
rect 1808 17240 1848 17272
rect 1880 17240 1950 17272
rect 50 17200 1950 17240
rect 50 17168 120 17200
rect 152 17168 192 17200
rect 224 17168 264 17200
rect 296 17168 336 17200
rect 368 17168 408 17200
rect 440 17168 480 17200
rect 512 17168 552 17200
rect 584 17168 624 17200
rect 656 17168 696 17200
rect 728 17168 768 17200
rect 800 17168 840 17200
rect 872 17168 912 17200
rect 944 17168 984 17200
rect 1016 17168 1056 17200
rect 1088 17168 1128 17200
rect 1160 17168 1200 17200
rect 1232 17168 1272 17200
rect 1304 17168 1344 17200
rect 1376 17168 1416 17200
rect 1448 17168 1488 17200
rect 1520 17168 1560 17200
rect 1592 17168 1632 17200
rect 1664 17168 1704 17200
rect 1736 17168 1776 17200
rect 1808 17168 1848 17200
rect 1880 17168 1950 17200
rect 50 17128 1950 17168
rect 50 17096 120 17128
rect 152 17096 192 17128
rect 224 17096 264 17128
rect 296 17096 336 17128
rect 368 17096 408 17128
rect 440 17096 480 17128
rect 512 17096 552 17128
rect 584 17096 624 17128
rect 656 17096 696 17128
rect 728 17096 768 17128
rect 800 17096 840 17128
rect 872 17096 912 17128
rect 944 17096 984 17128
rect 1016 17096 1056 17128
rect 1088 17096 1128 17128
rect 1160 17096 1200 17128
rect 1232 17096 1272 17128
rect 1304 17096 1344 17128
rect 1376 17096 1416 17128
rect 1448 17096 1488 17128
rect 1520 17096 1560 17128
rect 1592 17096 1632 17128
rect 1664 17096 1704 17128
rect 1736 17096 1776 17128
rect 1808 17096 1848 17128
rect 1880 17096 1950 17128
rect 50 17056 1950 17096
rect 50 17024 120 17056
rect 152 17024 192 17056
rect 224 17024 264 17056
rect 296 17024 336 17056
rect 368 17024 408 17056
rect 440 17024 480 17056
rect 512 17024 552 17056
rect 584 17024 624 17056
rect 656 17024 696 17056
rect 728 17024 768 17056
rect 800 17024 840 17056
rect 872 17024 912 17056
rect 944 17024 984 17056
rect 1016 17024 1056 17056
rect 1088 17024 1128 17056
rect 1160 17024 1200 17056
rect 1232 17024 1272 17056
rect 1304 17024 1344 17056
rect 1376 17024 1416 17056
rect 1448 17024 1488 17056
rect 1520 17024 1560 17056
rect 1592 17024 1632 17056
rect 1664 17024 1704 17056
rect 1736 17024 1776 17056
rect 1808 17024 1848 17056
rect 1880 17024 1950 17056
rect 50 16984 1950 17024
rect 50 16952 120 16984
rect 152 16952 192 16984
rect 224 16952 264 16984
rect 296 16952 336 16984
rect 368 16952 408 16984
rect 440 16952 480 16984
rect 512 16952 552 16984
rect 584 16952 624 16984
rect 656 16952 696 16984
rect 728 16952 768 16984
rect 800 16952 840 16984
rect 872 16952 912 16984
rect 944 16952 984 16984
rect 1016 16952 1056 16984
rect 1088 16952 1128 16984
rect 1160 16952 1200 16984
rect 1232 16952 1272 16984
rect 1304 16952 1344 16984
rect 1376 16952 1416 16984
rect 1448 16952 1488 16984
rect 1520 16952 1560 16984
rect 1592 16952 1632 16984
rect 1664 16952 1704 16984
rect 1736 16952 1776 16984
rect 1808 16952 1848 16984
rect 1880 16952 1950 16984
rect 50 16912 1950 16952
rect 50 16880 120 16912
rect 152 16880 192 16912
rect 224 16880 264 16912
rect 296 16880 336 16912
rect 368 16880 408 16912
rect 440 16880 480 16912
rect 512 16880 552 16912
rect 584 16880 624 16912
rect 656 16880 696 16912
rect 728 16880 768 16912
rect 800 16880 840 16912
rect 872 16880 912 16912
rect 944 16880 984 16912
rect 1016 16880 1056 16912
rect 1088 16880 1128 16912
rect 1160 16880 1200 16912
rect 1232 16880 1272 16912
rect 1304 16880 1344 16912
rect 1376 16880 1416 16912
rect 1448 16880 1488 16912
rect 1520 16880 1560 16912
rect 1592 16880 1632 16912
rect 1664 16880 1704 16912
rect 1736 16880 1776 16912
rect 1808 16880 1848 16912
rect 1880 16880 1950 16912
rect 50 16840 1950 16880
rect 50 16808 120 16840
rect 152 16808 192 16840
rect 224 16808 264 16840
rect 296 16808 336 16840
rect 368 16808 408 16840
rect 440 16808 480 16840
rect 512 16808 552 16840
rect 584 16808 624 16840
rect 656 16808 696 16840
rect 728 16808 768 16840
rect 800 16808 840 16840
rect 872 16808 912 16840
rect 944 16808 984 16840
rect 1016 16808 1056 16840
rect 1088 16808 1128 16840
rect 1160 16808 1200 16840
rect 1232 16808 1272 16840
rect 1304 16808 1344 16840
rect 1376 16808 1416 16840
rect 1448 16808 1488 16840
rect 1520 16808 1560 16840
rect 1592 16808 1632 16840
rect 1664 16808 1704 16840
rect 1736 16808 1776 16840
rect 1808 16808 1848 16840
rect 1880 16808 1950 16840
rect 50 16768 1950 16808
rect 50 16736 120 16768
rect 152 16736 192 16768
rect 224 16736 264 16768
rect 296 16736 336 16768
rect 368 16736 408 16768
rect 440 16736 480 16768
rect 512 16736 552 16768
rect 584 16736 624 16768
rect 656 16736 696 16768
rect 728 16736 768 16768
rect 800 16736 840 16768
rect 872 16736 912 16768
rect 944 16736 984 16768
rect 1016 16736 1056 16768
rect 1088 16736 1128 16768
rect 1160 16736 1200 16768
rect 1232 16736 1272 16768
rect 1304 16736 1344 16768
rect 1376 16736 1416 16768
rect 1448 16736 1488 16768
rect 1520 16736 1560 16768
rect 1592 16736 1632 16768
rect 1664 16736 1704 16768
rect 1736 16736 1776 16768
rect 1808 16736 1848 16768
rect 1880 16736 1950 16768
rect 50 16696 1950 16736
rect 50 16664 120 16696
rect 152 16664 192 16696
rect 224 16664 264 16696
rect 296 16664 336 16696
rect 368 16664 408 16696
rect 440 16664 480 16696
rect 512 16664 552 16696
rect 584 16664 624 16696
rect 656 16664 696 16696
rect 728 16664 768 16696
rect 800 16664 840 16696
rect 872 16664 912 16696
rect 944 16664 984 16696
rect 1016 16664 1056 16696
rect 1088 16664 1128 16696
rect 1160 16664 1200 16696
rect 1232 16664 1272 16696
rect 1304 16664 1344 16696
rect 1376 16664 1416 16696
rect 1448 16664 1488 16696
rect 1520 16664 1560 16696
rect 1592 16664 1632 16696
rect 1664 16664 1704 16696
rect 1736 16664 1776 16696
rect 1808 16664 1848 16696
rect 1880 16664 1950 16696
rect 50 16624 1950 16664
rect 50 16592 120 16624
rect 152 16592 192 16624
rect 224 16592 264 16624
rect 296 16592 336 16624
rect 368 16592 408 16624
rect 440 16592 480 16624
rect 512 16592 552 16624
rect 584 16592 624 16624
rect 656 16592 696 16624
rect 728 16592 768 16624
rect 800 16592 840 16624
rect 872 16592 912 16624
rect 944 16592 984 16624
rect 1016 16592 1056 16624
rect 1088 16592 1128 16624
rect 1160 16592 1200 16624
rect 1232 16592 1272 16624
rect 1304 16592 1344 16624
rect 1376 16592 1416 16624
rect 1448 16592 1488 16624
rect 1520 16592 1560 16624
rect 1592 16592 1632 16624
rect 1664 16592 1704 16624
rect 1736 16592 1776 16624
rect 1808 16592 1848 16624
rect 1880 16592 1950 16624
rect 50 16552 1950 16592
rect 50 16520 120 16552
rect 152 16520 192 16552
rect 224 16520 264 16552
rect 296 16520 336 16552
rect 368 16520 408 16552
rect 440 16520 480 16552
rect 512 16520 552 16552
rect 584 16520 624 16552
rect 656 16520 696 16552
rect 728 16520 768 16552
rect 800 16520 840 16552
rect 872 16520 912 16552
rect 944 16520 984 16552
rect 1016 16520 1056 16552
rect 1088 16520 1128 16552
rect 1160 16520 1200 16552
rect 1232 16520 1272 16552
rect 1304 16520 1344 16552
rect 1376 16520 1416 16552
rect 1448 16520 1488 16552
rect 1520 16520 1560 16552
rect 1592 16520 1632 16552
rect 1664 16520 1704 16552
rect 1736 16520 1776 16552
rect 1808 16520 1848 16552
rect 1880 16520 1950 16552
rect 50 16480 1950 16520
rect 50 16448 120 16480
rect 152 16448 192 16480
rect 224 16448 264 16480
rect 296 16448 336 16480
rect 368 16448 408 16480
rect 440 16448 480 16480
rect 512 16448 552 16480
rect 584 16448 624 16480
rect 656 16448 696 16480
rect 728 16448 768 16480
rect 800 16448 840 16480
rect 872 16448 912 16480
rect 944 16448 984 16480
rect 1016 16448 1056 16480
rect 1088 16448 1128 16480
rect 1160 16448 1200 16480
rect 1232 16448 1272 16480
rect 1304 16448 1344 16480
rect 1376 16448 1416 16480
rect 1448 16448 1488 16480
rect 1520 16448 1560 16480
rect 1592 16448 1632 16480
rect 1664 16448 1704 16480
rect 1736 16448 1776 16480
rect 1808 16448 1848 16480
rect 1880 16448 1950 16480
rect 50 16408 1950 16448
rect 50 16376 120 16408
rect 152 16376 192 16408
rect 224 16376 264 16408
rect 296 16376 336 16408
rect 368 16376 408 16408
rect 440 16376 480 16408
rect 512 16376 552 16408
rect 584 16376 624 16408
rect 656 16376 696 16408
rect 728 16376 768 16408
rect 800 16376 840 16408
rect 872 16376 912 16408
rect 944 16376 984 16408
rect 1016 16376 1056 16408
rect 1088 16376 1128 16408
rect 1160 16376 1200 16408
rect 1232 16376 1272 16408
rect 1304 16376 1344 16408
rect 1376 16376 1416 16408
rect 1448 16376 1488 16408
rect 1520 16376 1560 16408
rect 1592 16376 1632 16408
rect 1664 16376 1704 16408
rect 1736 16376 1776 16408
rect 1808 16376 1848 16408
rect 1880 16376 1950 16408
rect 50 16336 1950 16376
rect 50 16304 120 16336
rect 152 16304 192 16336
rect 224 16304 264 16336
rect 296 16304 336 16336
rect 368 16304 408 16336
rect 440 16304 480 16336
rect 512 16304 552 16336
rect 584 16304 624 16336
rect 656 16304 696 16336
rect 728 16304 768 16336
rect 800 16304 840 16336
rect 872 16304 912 16336
rect 944 16304 984 16336
rect 1016 16304 1056 16336
rect 1088 16304 1128 16336
rect 1160 16304 1200 16336
rect 1232 16304 1272 16336
rect 1304 16304 1344 16336
rect 1376 16304 1416 16336
rect 1448 16304 1488 16336
rect 1520 16304 1560 16336
rect 1592 16304 1632 16336
rect 1664 16304 1704 16336
rect 1736 16304 1776 16336
rect 1808 16304 1848 16336
rect 1880 16304 1950 16336
rect 50 16264 1950 16304
rect 50 16232 120 16264
rect 152 16232 192 16264
rect 224 16232 264 16264
rect 296 16232 336 16264
rect 368 16232 408 16264
rect 440 16232 480 16264
rect 512 16232 552 16264
rect 584 16232 624 16264
rect 656 16232 696 16264
rect 728 16232 768 16264
rect 800 16232 840 16264
rect 872 16232 912 16264
rect 944 16232 984 16264
rect 1016 16232 1056 16264
rect 1088 16232 1128 16264
rect 1160 16232 1200 16264
rect 1232 16232 1272 16264
rect 1304 16232 1344 16264
rect 1376 16232 1416 16264
rect 1448 16232 1488 16264
rect 1520 16232 1560 16264
rect 1592 16232 1632 16264
rect 1664 16232 1704 16264
rect 1736 16232 1776 16264
rect 1808 16232 1848 16264
rect 1880 16232 1950 16264
rect 50 16192 1950 16232
rect 50 16160 120 16192
rect 152 16160 192 16192
rect 224 16160 264 16192
rect 296 16160 336 16192
rect 368 16160 408 16192
rect 440 16160 480 16192
rect 512 16160 552 16192
rect 584 16160 624 16192
rect 656 16160 696 16192
rect 728 16160 768 16192
rect 800 16160 840 16192
rect 872 16160 912 16192
rect 944 16160 984 16192
rect 1016 16160 1056 16192
rect 1088 16160 1128 16192
rect 1160 16160 1200 16192
rect 1232 16160 1272 16192
rect 1304 16160 1344 16192
rect 1376 16160 1416 16192
rect 1448 16160 1488 16192
rect 1520 16160 1560 16192
rect 1592 16160 1632 16192
rect 1664 16160 1704 16192
rect 1736 16160 1776 16192
rect 1808 16160 1848 16192
rect 1880 16160 1950 16192
rect 50 16120 1950 16160
rect 50 16088 120 16120
rect 152 16088 192 16120
rect 224 16088 264 16120
rect 296 16088 336 16120
rect 368 16088 408 16120
rect 440 16088 480 16120
rect 512 16088 552 16120
rect 584 16088 624 16120
rect 656 16088 696 16120
rect 728 16088 768 16120
rect 800 16088 840 16120
rect 872 16088 912 16120
rect 944 16088 984 16120
rect 1016 16088 1056 16120
rect 1088 16088 1128 16120
rect 1160 16088 1200 16120
rect 1232 16088 1272 16120
rect 1304 16088 1344 16120
rect 1376 16088 1416 16120
rect 1448 16088 1488 16120
rect 1520 16088 1560 16120
rect 1592 16088 1632 16120
rect 1664 16088 1704 16120
rect 1736 16088 1776 16120
rect 1808 16088 1848 16120
rect 1880 16088 1950 16120
rect 50 16048 1950 16088
rect 50 16016 120 16048
rect 152 16016 192 16048
rect 224 16016 264 16048
rect 296 16016 336 16048
rect 368 16016 408 16048
rect 440 16016 480 16048
rect 512 16016 552 16048
rect 584 16016 624 16048
rect 656 16016 696 16048
rect 728 16016 768 16048
rect 800 16016 840 16048
rect 872 16016 912 16048
rect 944 16016 984 16048
rect 1016 16016 1056 16048
rect 1088 16016 1128 16048
rect 1160 16016 1200 16048
rect 1232 16016 1272 16048
rect 1304 16016 1344 16048
rect 1376 16016 1416 16048
rect 1448 16016 1488 16048
rect 1520 16016 1560 16048
rect 1592 16016 1632 16048
rect 1664 16016 1704 16048
rect 1736 16016 1776 16048
rect 1808 16016 1848 16048
rect 1880 16016 1950 16048
rect 50 15976 1950 16016
rect 50 15944 120 15976
rect 152 15944 192 15976
rect 224 15944 264 15976
rect 296 15944 336 15976
rect 368 15944 408 15976
rect 440 15944 480 15976
rect 512 15944 552 15976
rect 584 15944 624 15976
rect 656 15944 696 15976
rect 728 15944 768 15976
rect 800 15944 840 15976
rect 872 15944 912 15976
rect 944 15944 984 15976
rect 1016 15944 1056 15976
rect 1088 15944 1128 15976
rect 1160 15944 1200 15976
rect 1232 15944 1272 15976
rect 1304 15944 1344 15976
rect 1376 15944 1416 15976
rect 1448 15944 1488 15976
rect 1520 15944 1560 15976
rect 1592 15944 1632 15976
rect 1664 15944 1704 15976
rect 1736 15944 1776 15976
rect 1808 15944 1848 15976
rect 1880 15944 1950 15976
rect 50 15904 1950 15944
rect 50 15872 120 15904
rect 152 15872 192 15904
rect 224 15872 264 15904
rect 296 15872 336 15904
rect 368 15872 408 15904
rect 440 15872 480 15904
rect 512 15872 552 15904
rect 584 15872 624 15904
rect 656 15872 696 15904
rect 728 15872 768 15904
rect 800 15872 840 15904
rect 872 15872 912 15904
rect 944 15872 984 15904
rect 1016 15872 1056 15904
rect 1088 15872 1128 15904
rect 1160 15872 1200 15904
rect 1232 15872 1272 15904
rect 1304 15872 1344 15904
rect 1376 15872 1416 15904
rect 1448 15872 1488 15904
rect 1520 15872 1560 15904
rect 1592 15872 1632 15904
rect 1664 15872 1704 15904
rect 1736 15872 1776 15904
rect 1808 15872 1848 15904
rect 1880 15872 1950 15904
rect 50 15832 1950 15872
rect 50 15800 120 15832
rect 152 15800 192 15832
rect 224 15800 264 15832
rect 296 15800 336 15832
rect 368 15800 408 15832
rect 440 15800 480 15832
rect 512 15800 552 15832
rect 584 15800 624 15832
rect 656 15800 696 15832
rect 728 15800 768 15832
rect 800 15800 840 15832
rect 872 15800 912 15832
rect 944 15800 984 15832
rect 1016 15800 1056 15832
rect 1088 15800 1128 15832
rect 1160 15800 1200 15832
rect 1232 15800 1272 15832
rect 1304 15800 1344 15832
rect 1376 15800 1416 15832
rect 1448 15800 1488 15832
rect 1520 15800 1560 15832
rect 1592 15800 1632 15832
rect 1664 15800 1704 15832
rect 1736 15800 1776 15832
rect 1808 15800 1848 15832
rect 1880 15800 1950 15832
rect 50 15760 1950 15800
rect 50 15728 120 15760
rect 152 15728 192 15760
rect 224 15728 264 15760
rect 296 15728 336 15760
rect 368 15728 408 15760
rect 440 15728 480 15760
rect 512 15728 552 15760
rect 584 15728 624 15760
rect 656 15728 696 15760
rect 728 15728 768 15760
rect 800 15728 840 15760
rect 872 15728 912 15760
rect 944 15728 984 15760
rect 1016 15728 1056 15760
rect 1088 15728 1128 15760
rect 1160 15728 1200 15760
rect 1232 15728 1272 15760
rect 1304 15728 1344 15760
rect 1376 15728 1416 15760
rect 1448 15728 1488 15760
rect 1520 15728 1560 15760
rect 1592 15728 1632 15760
rect 1664 15728 1704 15760
rect 1736 15728 1776 15760
rect 1808 15728 1848 15760
rect 1880 15728 1950 15760
rect 50 15688 1950 15728
rect 50 15656 120 15688
rect 152 15656 192 15688
rect 224 15656 264 15688
rect 296 15656 336 15688
rect 368 15656 408 15688
rect 440 15656 480 15688
rect 512 15656 552 15688
rect 584 15656 624 15688
rect 656 15656 696 15688
rect 728 15656 768 15688
rect 800 15656 840 15688
rect 872 15656 912 15688
rect 944 15656 984 15688
rect 1016 15656 1056 15688
rect 1088 15656 1128 15688
rect 1160 15656 1200 15688
rect 1232 15656 1272 15688
rect 1304 15656 1344 15688
rect 1376 15656 1416 15688
rect 1448 15656 1488 15688
rect 1520 15656 1560 15688
rect 1592 15656 1632 15688
rect 1664 15656 1704 15688
rect 1736 15656 1776 15688
rect 1808 15656 1848 15688
rect 1880 15656 1950 15688
rect 50 15616 1950 15656
rect 50 15584 120 15616
rect 152 15584 192 15616
rect 224 15584 264 15616
rect 296 15584 336 15616
rect 368 15584 408 15616
rect 440 15584 480 15616
rect 512 15584 552 15616
rect 584 15584 624 15616
rect 656 15584 696 15616
rect 728 15584 768 15616
rect 800 15584 840 15616
rect 872 15584 912 15616
rect 944 15584 984 15616
rect 1016 15584 1056 15616
rect 1088 15584 1128 15616
rect 1160 15584 1200 15616
rect 1232 15584 1272 15616
rect 1304 15584 1344 15616
rect 1376 15584 1416 15616
rect 1448 15584 1488 15616
rect 1520 15584 1560 15616
rect 1592 15584 1632 15616
rect 1664 15584 1704 15616
rect 1736 15584 1776 15616
rect 1808 15584 1848 15616
rect 1880 15584 1950 15616
rect 50 15544 1950 15584
rect 50 15512 120 15544
rect 152 15512 192 15544
rect 224 15512 264 15544
rect 296 15512 336 15544
rect 368 15512 408 15544
rect 440 15512 480 15544
rect 512 15512 552 15544
rect 584 15512 624 15544
rect 656 15512 696 15544
rect 728 15512 768 15544
rect 800 15512 840 15544
rect 872 15512 912 15544
rect 944 15512 984 15544
rect 1016 15512 1056 15544
rect 1088 15512 1128 15544
rect 1160 15512 1200 15544
rect 1232 15512 1272 15544
rect 1304 15512 1344 15544
rect 1376 15512 1416 15544
rect 1448 15512 1488 15544
rect 1520 15512 1560 15544
rect 1592 15512 1632 15544
rect 1664 15512 1704 15544
rect 1736 15512 1776 15544
rect 1808 15512 1848 15544
rect 1880 15512 1950 15544
rect 50 15472 1950 15512
rect 50 15440 120 15472
rect 152 15440 192 15472
rect 224 15440 264 15472
rect 296 15440 336 15472
rect 368 15440 408 15472
rect 440 15440 480 15472
rect 512 15440 552 15472
rect 584 15440 624 15472
rect 656 15440 696 15472
rect 728 15440 768 15472
rect 800 15440 840 15472
rect 872 15440 912 15472
rect 944 15440 984 15472
rect 1016 15440 1056 15472
rect 1088 15440 1128 15472
rect 1160 15440 1200 15472
rect 1232 15440 1272 15472
rect 1304 15440 1344 15472
rect 1376 15440 1416 15472
rect 1448 15440 1488 15472
rect 1520 15440 1560 15472
rect 1592 15440 1632 15472
rect 1664 15440 1704 15472
rect 1736 15440 1776 15472
rect 1808 15440 1848 15472
rect 1880 15440 1950 15472
rect 50 15400 1950 15440
rect 50 15368 120 15400
rect 152 15368 192 15400
rect 224 15368 264 15400
rect 296 15368 336 15400
rect 368 15368 408 15400
rect 440 15368 480 15400
rect 512 15368 552 15400
rect 584 15368 624 15400
rect 656 15368 696 15400
rect 728 15368 768 15400
rect 800 15368 840 15400
rect 872 15368 912 15400
rect 944 15368 984 15400
rect 1016 15368 1056 15400
rect 1088 15368 1128 15400
rect 1160 15368 1200 15400
rect 1232 15368 1272 15400
rect 1304 15368 1344 15400
rect 1376 15368 1416 15400
rect 1448 15368 1488 15400
rect 1520 15368 1560 15400
rect 1592 15368 1632 15400
rect 1664 15368 1704 15400
rect 1736 15368 1776 15400
rect 1808 15368 1848 15400
rect 1880 15368 1950 15400
rect 50 15328 1950 15368
rect 50 15296 120 15328
rect 152 15296 192 15328
rect 224 15296 264 15328
rect 296 15296 336 15328
rect 368 15296 408 15328
rect 440 15296 480 15328
rect 512 15296 552 15328
rect 584 15296 624 15328
rect 656 15296 696 15328
rect 728 15296 768 15328
rect 800 15296 840 15328
rect 872 15296 912 15328
rect 944 15296 984 15328
rect 1016 15296 1056 15328
rect 1088 15296 1128 15328
rect 1160 15296 1200 15328
rect 1232 15296 1272 15328
rect 1304 15296 1344 15328
rect 1376 15296 1416 15328
rect 1448 15296 1488 15328
rect 1520 15296 1560 15328
rect 1592 15296 1632 15328
rect 1664 15296 1704 15328
rect 1736 15296 1776 15328
rect 1808 15296 1848 15328
rect 1880 15296 1950 15328
rect 50 15256 1950 15296
rect 50 15224 120 15256
rect 152 15224 192 15256
rect 224 15224 264 15256
rect 296 15224 336 15256
rect 368 15224 408 15256
rect 440 15224 480 15256
rect 512 15224 552 15256
rect 584 15224 624 15256
rect 656 15224 696 15256
rect 728 15224 768 15256
rect 800 15224 840 15256
rect 872 15224 912 15256
rect 944 15224 984 15256
rect 1016 15224 1056 15256
rect 1088 15224 1128 15256
rect 1160 15224 1200 15256
rect 1232 15224 1272 15256
rect 1304 15224 1344 15256
rect 1376 15224 1416 15256
rect 1448 15224 1488 15256
rect 1520 15224 1560 15256
rect 1592 15224 1632 15256
rect 1664 15224 1704 15256
rect 1736 15224 1776 15256
rect 1808 15224 1848 15256
rect 1880 15224 1950 15256
rect 50 15184 1950 15224
rect 50 15152 120 15184
rect 152 15152 192 15184
rect 224 15152 264 15184
rect 296 15152 336 15184
rect 368 15152 408 15184
rect 440 15152 480 15184
rect 512 15152 552 15184
rect 584 15152 624 15184
rect 656 15152 696 15184
rect 728 15152 768 15184
rect 800 15152 840 15184
rect 872 15152 912 15184
rect 944 15152 984 15184
rect 1016 15152 1056 15184
rect 1088 15152 1128 15184
rect 1160 15152 1200 15184
rect 1232 15152 1272 15184
rect 1304 15152 1344 15184
rect 1376 15152 1416 15184
rect 1448 15152 1488 15184
rect 1520 15152 1560 15184
rect 1592 15152 1632 15184
rect 1664 15152 1704 15184
rect 1736 15152 1776 15184
rect 1808 15152 1848 15184
rect 1880 15152 1950 15184
rect 50 15112 1950 15152
rect 50 15080 120 15112
rect 152 15080 192 15112
rect 224 15080 264 15112
rect 296 15080 336 15112
rect 368 15080 408 15112
rect 440 15080 480 15112
rect 512 15080 552 15112
rect 584 15080 624 15112
rect 656 15080 696 15112
rect 728 15080 768 15112
rect 800 15080 840 15112
rect 872 15080 912 15112
rect 944 15080 984 15112
rect 1016 15080 1056 15112
rect 1088 15080 1128 15112
rect 1160 15080 1200 15112
rect 1232 15080 1272 15112
rect 1304 15080 1344 15112
rect 1376 15080 1416 15112
rect 1448 15080 1488 15112
rect 1520 15080 1560 15112
rect 1592 15080 1632 15112
rect 1664 15080 1704 15112
rect 1736 15080 1776 15112
rect 1808 15080 1848 15112
rect 1880 15080 1950 15112
rect 50 15040 1950 15080
rect 50 15008 120 15040
rect 152 15008 192 15040
rect 224 15008 264 15040
rect 296 15008 336 15040
rect 368 15008 408 15040
rect 440 15008 480 15040
rect 512 15008 552 15040
rect 584 15008 624 15040
rect 656 15008 696 15040
rect 728 15008 768 15040
rect 800 15008 840 15040
rect 872 15008 912 15040
rect 944 15008 984 15040
rect 1016 15008 1056 15040
rect 1088 15008 1128 15040
rect 1160 15008 1200 15040
rect 1232 15008 1272 15040
rect 1304 15008 1344 15040
rect 1376 15008 1416 15040
rect 1448 15008 1488 15040
rect 1520 15008 1560 15040
rect 1592 15008 1632 15040
rect 1664 15008 1704 15040
rect 1736 15008 1776 15040
rect 1808 15008 1848 15040
rect 1880 15008 1950 15040
rect 50 14968 1950 15008
rect 50 14936 120 14968
rect 152 14936 192 14968
rect 224 14936 264 14968
rect 296 14936 336 14968
rect 368 14936 408 14968
rect 440 14936 480 14968
rect 512 14936 552 14968
rect 584 14936 624 14968
rect 656 14936 696 14968
rect 728 14936 768 14968
rect 800 14936 840 14968
rect 872 14936 912 14968
rect 944 14936 984 14968
rect 1016 14936 1056 14968
rect 1088 14936 1128 14968
rect 1160 14936 1200 14968
rect 1232 14936 1272 14968
rect 1304 14936 1344 14968
rect 1376 14936 1416 14968
rect 1448 14936 1488 14968
rect 1520 14936 1560 14968
rect 1592 14936 1632 14968
rect 1664 14936 1704 14968
rect 1736 14936 1776 14968
rect 1808 14936 1848 14968
rect 1880 14936 1950 14968
rect 50 14896 1950 14936
rect 50 14864 120 14896
rect 152 14864 192 14896
rect 224 14864 264 14896
rect 296 14864 336 14896
rect 368 14864 408 14896
rect 440 14864 480 14896
rect 512 14864 552 14896
rect 584 14864 624 14896
rect 656 14864 696 14896
rect 728 14864 768 14896
rect 800 14864 840 14896
rect 872 14864 912 14896
rect 944 14864 984 14896
rect 1016 14864 1056 14896
rect 1088 14864 1128 14896
rect 1160 14864 1200 14896
rect 1232 14864 1272 14896
rect 1304 14864 1344 14896
rect 1376 14864 1416 14896
rect 1448 14864 1488 14896
rect 1520 14864 1560 14896
rect 1592 14864 1632 14896
rect 1664 14864 1704 14896
rect 1736 14864 1776 14896
rect 1808 14864 1848 14896
rect 1880 14864 1950 14896
rect 50 14824 1950 14864
rect 50 14792 120 14824
rect 152 14792 192 14824
rect 224 14792 264 14824
rect 296 14792 336 14824
rect 368 14792 408 14824
rect 440 14792 480 14824
rect 512 14792 552 14824
rect 584 14792 624 14824
rect 656 14792 696 14824
rect 728 14792 768 14824
rect 800 14792 840 14824
rect 872 14792 912 14824
rect 944 14792 984 14824
rect 1016 14792 1056 14824
rect 1088 14792 1128 14824
rect 1160 14792 1200 14824
rect 1232 14792 1272 14824
rect 1304 14792 1344 14824
rect 1376 14792 1416 14824
rect 1448 14792 1488 14824
rect 1520 14792 1560 14824
rect 1592 14792 1632 14824
rect 1664 14792 1704 14824
rect 1736 14792 1776 14824
rect 1808 14792 1848 14824
rect 1880 14792 1950 14824
rect 50 14752 1950 14792
rect 50 14720 120 14752
rect 152 14720 192 14752
rect 224 14720 264 14752
rect 296 14720 336 14752
rect 368 14720 408 14752
rect 440 14720 480 14752
rect 512 14720 552 14752
rect 584 14720 624 14752
rect 656 14720 696 14752
rect 728 14720 768 14752
rect 800 14720 840 14752
rect 872 14720 912 14752
rect 944 14720 984 14752
rect 1016 14720 1056 14752
rect 1088 14720 1128 14752
rect 1160 14720 1200 14752
rect 1232 14720 1272 14752
rect 1304 14720 1344 14752
rect 1376 14720 1416 14752
rect 1448 14720 1488 14752
rect 1520 14720 1560 14752
rect 1592 14720 1632 14752
rect 1664 14720 1704 14752
rect 1736 14720 1776 14752
rect 1808 14720 1848 14752
rect 1880 14720 1950 14752
rect 50 14680 1950 14720
rect 50 14648 120 14680
rect 152 14648 192 14680
rect 224 14648 264 14680
rect 296 14648 336 14680
rect 368 14648 408 14680
rect 440 14648 480 14680
rect 512 14648 552 14680
rect 584 14648 624 14680
rect 656 14648 696 14680
rect 728 14648 768 14680
rect 800 14648 840 14680
rect 872 14648 912 14680
rect 944 14648 984 14680
rect 1016 14648 1056 14680
rect 1088 14648 1128 14680
rect 1160 14648 1200 14680
rect 1232 14648 1272 14680
rect 1304 14648 1344 14680
rect 1376 14648 1416 14680
rect 1448 14648 1488 14680
rect 1520 14648 1560 14680
rect 1592 14648 1632 14680
rect 1664 14648 1704 14680
rect 1736 14648 1776 14680
rect 1808 14648 1848 14680
rect 1880 14648 1950 14680
rect 50 14608 1950 14648
rect 50 14576 120 14608
rect 152 14576 192 14608
rect 224 14576 264 14608
rect 296 14576 336 14608
rect 368 14576 408 14608
rect 440 14576 480 14608
rect 512 14576 552 14608
rect 584 14576 624 14608
rect 656 14576 696 14608
rect 728 14576 768 14608
rect 800 14576 840 14608
rect 872 14576 912 14608
rect 944 14576 984 14608
rect 1016 14576 1056 14608
rect 1088 14576 1128 14608
rect 1160 14576 1200 14608
rect 1232 14576 1272 14608
rect 1304 14576 1344 14608
rect 1376 14576 1416 14608
rect 1448 14576 1488 14608
rect 1520 14576 1560 14608
rect 1592 14576 1632 14608
rect 1664 14576 1704 14608
rect 1736 14576 1776 14608
rect 1808 14576 1848 14608
rect 1880 14576 1950 14608
rect 50 14536 1950 14576
rect 50 14504 120 14536
rect 152 14504 192 14536
rect 224 14504 264 14536
rect 296 14504 336 14536
rect 368 14504 408 14536
rect 440 14504 480 14536
rect 512 14504 552 14536
rect 584 14504 624 14536
rect 656 14504 696 14536
rect 728 14504 768 14536
rect 800 14504 840 14536
rect 872 14504 912 14536
rect 944 14504 984 14536
rect 1016 14504 1056 14536
rect 1088 14504 1128 14536
rect 1160 14504 1200 14536
rect 1232 14504 1272 14536
rect 1304 14504 1344 14536
rect 1376 14504 1416 14536
rect 1448 14504 1488 14536
rect 1520 14504 1560 14536
rect 1592 14504 1632 14536
rect 1664 14504 1704 14536
rect 1736 14504 1776 14536
rect 1808 14504 1848 14536
rect 1880 14504 1950 14536
rect 50 14464 1950 14504
rect 50 14432 120 14464
rect 152 14432 192 14464
rect 224 14432 264 14464
rect 296 14432 336 14464
rect 368 14432 408 14464
rect 440 14432 480 14464
rect 512 14432 552 14464
rect 584 14432 624 14464
rect 656 14432 696 14464
rect 728 14432 768 14464
rect 800 14432 840 14464
rect 872 14432 912 14464
rect 944 14432 984 14464
rect 1016 14432 1056 14464
rect 1088 14432 1128 14464
rect 1160 14432 1200 14464
rect 1232 14432 1272 14464
rect 1304 14432 1344 14464
rect 1376 14432 1416 14464
rect 1448 14432 1488 14464
rect 1520 14432 1560 14464
rect 1592 14432 1632 14464
rect 1664 14432 1704 14464
rect 1736 14432 1776 14464
rect 1808 14432 1848 14464
rect 1880 14432 1950 14464
rect 50 14392 1950 14432
rect 50 14360 120 14392
rect 152 14360 192 14392
rect 224 14360 264 14392
rect 296 14360 336 14392
rect 368 14360 408 14392
rect 440 14360 480 14392
rect 512 14360 552 14392
rect 584 14360 624 14392
rect 656 14360 696 14392
rect 728 14360 768 14392
rect 800 14360 840 14392
rect 872 14360 912 14392
rect 944 14360 984 14392
rect 1016 14360 1056 14392
rect 1088 14360 1128 14392
rect 1160 14360 1200 14392
rect 1232 14360 1272 14392
rect 1304 14360 1344 14392
rect 1376 14360 1416 14392
rect 1448 14360 1488 14392
rect 1520 14360 1560 14392
rect 1592 14360 1632 14392
rect 1664 14360 1704 14392
rect 1736 14360 1776 14392
rect 1808 14360 1848 14392
rect 1880 14360 1950 14392
rect 50 14320 1950 14360
rect 50 14288 120 14320
rect 152 14288 192 14320
rect 224 14288 264 14320
rect 296 14288 336 14320
rect 368 14288 408 14320
rect 440 14288 480 14320
rect 512 14288 552 14320
rect 584 14288 624 14320
rect 656 14288 696 14320
rect 728 14288 768 14320
rect 800 14288 840 14320
rect 872 14288 912 14320
rect 944 14288 984 14320
rect 1016 14288 1056 14320
rect 1088 14288 1128 14320
rect 1160 14288 1200 14320
rect 1232 14288 1272 14320
rect 1304 14288 1344 14320
rect 1376 14288 1416 14320
rect 1448 14288 1488 14320
rect 1520 14288 1560 14320
rect 1592 14288 1632 14320
rect 1664 14288 1704 14320
rect 1736 14288 1776 14320
rect 1808 14288 1848 14320
rect 1880 14288 1950 14320
rect 50 14248 1950 14288
rect 50 14216 120 14248
rect 152 14216 192 14248
rect 224 14216 264 14248
rect 296 14216 336 14248
rect 368 14216 408 14248
rect 440 14216 480 14248
rect 512 14216 552 14248
rect 584 14216 624 14248
rect 656 14216 696 14248
rect 728 14216 768 14248
rect 800 14216 840 14248
rect 872 14216 912 14248
rect 944 14216 984 14248
rect 1016 14216 1056 14248
rect 1088 14216 1128 14248
rect 1160 14216 1200 14248
rect 1232 14216 1272 14248
rect 1304 14216 1344 14248
rect 1376 14216 1416 14248
rect 1448 14216 1488 14248
rect 1520 14216 1560 14248
rect 1592 14216 1632 14248
rect 1664 14216 1704 14248
rect 1736 14216 1776 14248
rect 1808 14216 1848 14248
rect 1880 14216 1950 14248
rect 50 14176 1950 14216
rect 50 14144 120 14176
rect 152 14144 192 14176
rect 224 14144 264 14176
rect 296 14144 336 14176
rect 368 14144 408 14176
rect 440 14144 480 14176
rect 512 14144 552 14176
rect 584 14144 624 14176
rect 656 14144 696 14176
rect 728 14144 768 14176
rect 800 14144 840 14176
rect 872 14144 912 14176
rect 944 14144 984 14176
rect 1016 14144 1056 14176
rect 1088 14144 1128 14176
rect 1160 14144 1200 14176
rect 1232 14144 1272 14176
rect 1304 14144 1344 14176
rect 1376 14144 1416 14176
rect 1448 14144 1488 14176
rect 1520 14144 1560 14176
rect 1592 14144 1632 14176
rect 1664 14144 1704 14176
rect 1736 14144 1776 14176
rect 1808 14144 1848 14176
rect 1880 14144 1950 14176
rect 50 14104 1950 14144
rect 50 14072 120 14104
rect 152 14072 192 14104
rect 224 14072 264 14104
rect 296 14072 336 14104
rect 368 14072 408 14104
rect 440 14072 480 14104
rect 512 14072 552 14104
rect 584 14072 624 14104
rect 656 14072 696 14104
rect 728 14072 768 14104
rect 800 14072 840 14104
rect 872 14072 912 14104
rect 944 14072 984 14104
rect 1016 14072 1056 14104
rect 1088 14072 1128 14104
rect 1160 14072 1200 14104
rect 1232 14072 1272 14104
rect 1304 14072 1344 14104
rect 1376 14072 1416 14104
rect 1448 14072 1488 14104
rect 1520 14072 1560 14104
rect 1592 14072 1632 14104
rect 1664 14072 1704 14104
rect 1736 14072 1776 14104
rect 1808 14072 1848 14104
rect 1880 14072 1950 14104
rect 50 14032 1950 14072
rect 50 14000 120 14032
rect 152 14000 192 14032
rect 224 14000 264 14032
rect 296 14000 336 14032
rect 368 14000 408 14032
rect 440 14000 480 14032
rect 512 14000 552 14032
rect 584 14000 624 14032
rect 656 14000 696 14032
rect 728 14000 768 14032
rect 800 14000 840 14032
rect 872 14000 912 14032
rect 944 14000 984 14032
rect 1016 14000 1056 14032
rect 1088 14000 1128 14032
rect 1160 14000 1200 14032
rect 1232 14000 1272 14032
rect 1304 14000 1344 14032
rect 1376 14000 1416 14032
rect 1448 14000 1488 14032
rect 1520 14000 1560 14032
rect 1592 14000 1632 14032
rect 1664 14000 1704 14032
rect 1736 14000 1776 14032
rect 1808 14000 1848 14032
rect 1880 14000 1950 14032
rect 50 13960 1950 14000
rect 50 13928 120 13960
rect 152 13928 192 13960
rect 224 13928 264 13960
rect 296 13928 336 13960
rect 368 13928 408 13960
rect 440 13928 480 13960
rect 512 13928 552 13960
rect 584 13928 624 13960
rect 656 13928 696 13960
rect 728 13928 768 13960
rect 800 13928 840 13960
rect 872 13928 912 13960
rect 944 13928 984 13960
rect 1016 13928 1056 13960
rect 1088 13928 1128 13960
rect 1160 13928 1200 13960
rect 1232 13928 1272 13960
rect 1304 13928 1344 13960
rect 1376 13928 1416 13960
rect 1448 13928 1488 13960
rect 1520 13928 1560 13960
rect 1592 13928 1632 13960
rect 1664 13928 1704 13960
rect 1736 13928 1776 13960
rect 1808 13928 1848 13960
rect 1880 13928 1950 13960
rect 50 13888 1950 13928
rect 50 13856 120 13888
rect 152 13856 192 13888
rect 224 13856 264 13888
rect 296 13856 336 13888
rect 368 13856 408 13888
rect 440 13856 480 13888
rect 512 13856 552 13888
rect 584 13856 624 13888
rect 656 13856 696 13888
rect 728 13856 768 13888
rect 800 13856 840 13888
rect 872 13856 912 13888
rect 944 13856 984 13888
rect 1016 13856 1056 13888
rect 1088 13856 1128 13888
rect 1160 13856 1200 13888
rect 1232 13856 1272 13888
rect 1304 13856 1344 13888
rect 1376 13856 1416 13888
rect 1448 13856 1488 13888
rect 1520 13856 1560 13888
rect 1592 13856 1632 13888
rect 1664 13856 1704 13888
rect 1736 13856 1776 13888
rect 1808 13856 1848 13888
rect 1880 13856 1950 13888
rect 50 13816 1950 13856
rect 50 13784 120 13816
rect 152 13784 192 13816
rect 224 13784 264 13816
rect 296 13784 336 13816
rect 368 13784 408 13816
rect 440 13784 480 13816
rect 512 13784 552 13816
rect 584 13784 624 13816
rect 656 13784 696 13816
rect 728 13784 768 13816
rect 800 13784 840 13816
rect 872 13784 912 13816
rect 944 13784 984 13816
rect 1016 13784 1056 13816
rect 1088 13784 1128 13816
rect 1160 13784 1200 13816
rect 1232 13784 1272 13816
rect 1304 13784 1344 13816
rect 1376 13784 1416 13816
rect 1448 13784 1488 13816
rect 1520 13784 1560 13816
rect 1592 13784 1632 13816
rect 1664 13784 1704 13816
rect 1736 13784 1776 13816
rect 1808 13784 1848 13816
rect 1880 13784 1950 13816
rect 50 13744 1950 13784
rect 50 13712 120 13744
rect 152 13712 192 13744
rect 224 13712 264 13744
rect 296 13712 336 13744
rect 368 13712 408 13744
rect 440 13712 480 13744
rect 512 13712 552 13744
rect 584 13712 624 13744
rect 656 13712 696 13744
rect 728 13712 768 13744
rect 800 13712 840 13744
rect 872 13712 912 13744
rect 944 13712 984 13744
rect 1016 13712 1056 13744
rect 1088 13712 1128 13744
rect 1160 13712 1200 13744
rect 1232 13712 1272 13744
rect 1304 13712 1344 13744
rect 1376 13712 1416 13744
rect 1448 13712 1488 13744
rect 1520 13712 1560 13744
rect 1592 13712 1632 13744
rect 1664 13712 1704 13744
rect 1736 13712 1776 13744
rect 1808 13712 1848 13744
rect 1880 13712 1950 13744
rect 50 13672 1950 13712
rect 50 13640 120 13672
rect 152 13640 192 13672
rect 224 13640 264 13672
rect 296 13640 336 13672
rect 368 13640 408 13672
rect 440 13640 480 13672
rect 512 13640 552 13672
rect 584 13640 624 13672
rect 656 13640 696 13672
rect 728 13640 768 13672
rect 800 13640 840 13672
rect 872 13640 912 13672
rect 944 13640 984 13672
rect 1016 13640 1056 13672
rect 1088 13640 1128 13672
rect 1160 13640 1200 13672
rect 1232 13640 1272 13672
rect 1304 13640 1344 13672
rect 1376 13640 1416 13672
rect 1448 13640 1488 13672
rect 1520 13640 1560 13672
rect 1592 13640 1632 13672
rect 1664 13640 1704 13672
rect 1736 13640 1776 13672
rect 1808 13640 1848 13672
rect 1880 13640 1950 13672
rect 50 13600 1950 13640
rect 50 13568 120 13600
rect 152 13568 192 13600
rect 224 13568 264 13600
rect 296 13568 336 13600
rect 368 13568 408 13600
rect 440 13568 480 13600
rect 512 13568 552 13600
rect 584 13568 624 13600
rect 656 13568 696 13600
rect 728 13568 768 13600
rect 800 13568 840 13600
rect 872 13568 912 13600
rect 944 13568 984 13600
rect 1016 13568 1056 13600
rect 1088 13568 1128 13600
rect 1160 13568 1200 13600
rect 1232 13568 1272 13600
rect 1304 13568 1344 13600
rect 1376 13568 1416 13600
rect 1448 13568 1488 13600
rect 1520 13568 1560 13600
rect 1592 13568 1632 13600
rect 1664 13568 1704 13600
rect 1736 13568 1776 13600
rect 1808 13568 1848 13600
rect 1880 13568 1950 13600
rect 50 13528 1950 13568
rect 50 13496 120 13528
rect 152 13496 192 13528
rect 224 13496 264 13528
rect 296 13496 336 13528
rect 368 13496 408 13528
rect 440 13496 480 13528
rect 512 13496 552 13528
rect 584 13496 624 13528
rect 656 13496 696 13528
rect 728 13496 768 13528
rect 800 13496 840 13528
rect 872 13496 912 13528
rect 944 13496 984 13528
rect 1016 13496 1056 13528
rect 1088 13496 1128 13528
rect 1160 13496 1200 13528
rect 1232 13496 1272 13528
rect 1304 13496 1344 13528
rect 1376 13496 1416 13528
rect 1448 13496 1488 13528
rect 1520 13496 1560 13528
rect 1592 13496 1632 13528
rect 1664 13496 1704 13528
rect 1736 13496 1776 13528
rect 1808 13496 1848 13528
rect 1880 13496 1950 13528
rect 50 13456 1950 13496
rect 50 13424 120 13456
rect 152 13424 192 13456
rect 224 13424 264 13456
rect 296 13424 336 13456
rect 368 13424 408 13456
rect 440 13424 480 13456
rect 512 13424 552 13456
rect 584 13424 624 13456
rect 656 13424 696 13456
rect 728 13424 768 13456
rect 800 13424 840 13456
rect 872 13424 912 13456
rect 944 13424 984 13456
rect 1016 13424 1056 13456
rect 1088 13424 1128 13456
rect 1160 13424 1200 13456
rect 1232 13424 1272 13456
rect 1304 13424 1344 13456
rect 1376 13424 1416 13456
rect 1448 13424 1488 13456
rect 1520 13424 1560 13456
rect 1592 13424 1632 13456
rect 1664 13424 1704 13456
rect 1736 13424 1776 13456
rect 1808 13424 1848 13456
rect 1880 13424 1950 13456
rect 50 13384 1950 13424
rect 50 13352 120 13384
rect 152 13352 192 13384
rect 224 13352 264 13384
rect 296 13352 336 13384
rect 368 13352 408 13384
rect 440 13352 480 13384
rect 512 13352 552 13384
rect 584 13352 624 13384
rect 656 13352 696 13384
rect 728 13352 768 13384
rect 800 13352 840 13384
rect 872 13352 912 13384
rect 944 13352 984 13384
rect 1016 13352 1056 13384
rect 1088 13352 1128 13384
rect 1160 13352 1200 13384
rect 1232 13352 1272 13384
rect 1304 13352 1344 13384
rect 1376 13352 1416 13384
rect 1448 13352 1488 13384
rect 1520 13352 1560 13384
rect 1592 13352 1632 13384
rect 1664 13352 1704 13384
rect 1736 13352 1776 13384
rect 1808 13352 1848 13384
rect 1880 13352 1950 13384
rect 50 13312 1950 13352
rect 50 13280 120 13312
rect 152 13280 192 13312
rect 224 13280 264 13312
rect 296 13280 336 13312
rect 368 13280 408 13312
rect 440 13280 480 13312
rect 512 13280 552 13312
rect 584 13280 624 13312
rect 656 13280 696 13312
rect 728 13280 768 13312
rect 800 13280 840 13312
rect 872 13280 912 13312
rect 944 13280 984 13312
rect 1016 13280 1056 13312
rect 1088 13280 1128 13312
rect 1160 13280 1200 13312
rect 1232 13280 1272 13312
rect 1304 13280 1344 13312
rect 1376 13280 1416 13312
rect 1448 13280 1488 13312
rect 1520 13280 1560 13312
rect 1592 13280 1632 13312
rect 1664 13280 1704 13312
rect 1736 13280 1776 13312
rect 1808 13280 1848 13312
rect 1880 13280 1950 13312
rect 50 13240 1950 13280
rect 50 13208 120 13240
rect 152 13208 192 13240
rect 224 13208 264 13240
rect 296 13208 336 13240
rect 368 13208 408 13240
rect 440 13208 480 13240
rect 512 13208 552 13240
rect 584 13208 624 13240
rect 656 13208 696 13240
rect 728 13208 768 13240
rect 800 13208 840 13240
rect 872 13208 912 13240
rect 944 13208 984 13240
rect 1016 13208 1056 13240
rect 1088 13208 1128 13240
rect 1160 13208 1200 13240
rect 1232 13208 1272 13240
rect 1304 13208 1344 13240
rect 1376 13208 1416 13240
rect 1448 13208 1488 13240
rect 1520 13208 1560 13240
rect 1592 13208 1632 13240
rect 1664 13208 1704 13240
rect 1736 13208 1776 13240
rect 1808 13208 1848 13240
rect 1880 13208 1950 13240
rect 50 13168 1950 13208
rect 50 13136 120 13168
rect 152 13136 192 13168
rect 224 13136 264 13168
rect 296 13136 336 13168
rect 368 13136 408 13168
rect 440 13136 480 13168
rect 512 13136 552 13168
rect 584 13136 624 13168
rect 656 13136 696 13168
rect 728 13136 768 13168
rect 800 13136 840 13168
rect 872 13136 912 13168
rect 944 13136 984 13168
rect 1016 13136 1056 13168
rect 1088 13136 1128 13168
rect 1160 13136 1200 13168
rect 1232 13136 1272 13168
rect 1304 13136 1344 13168
rect 1376 13136 1416 13168
rect 1448 13136 1488 13168
rect 1520 13136 1560 13168
rect 1592 13136 1632 13168
rect 1664 13136 1704 13168
rect 1736 13136 1776 13168
rect 1808 13136 1848 13168
rect 1880 13136 1950 13168
rect 50 13096 1950 13136
rect 50 13064 120 13096
rect 152 13064 192 13096
rect 224 13064 264 13096
rect 296 13064 336 13096
rect 368 13064 408 13096
rect 440 13064 480 13096
rect 512 13064 552 13096
rect 584 13064 624 13096
rect 656 13064 696 13096
rect 728 13064 768 13096
rect 800 13064 840 13096
rect 872 13064 912 13096
rect 944 13064 984 13096
rect 1016 13064 1056 13096
rect 1088 13064 1128 13096
rect 1160 13064 1200 13096
rect 1232 13064 1272 13096
rect 1304 13064 1344 13096
rect 1376 13064 1416 13096
rect 1448 13064 1488 13096
rect 1520 13064 1560 13096
rect 1592 13064 1632 13096
rect 1664 13064 1704 13096
rect 1736 13064 1776 13096
rect 1808 13064 1848 13096
rect 1880 13064 1950 13096
rect 50 13000 1950 13064
<< nsubdiff >>
rect 192 33384 224 33416
rect 264 33384 296 33416
rect 336 33384 368 33416
rect 408 33384 440 33416
rect 480 33384 512 33416
rect 552 33384 584 33416
rect 624 33384 656 33416
rect 696 33384 728 33416
rect 768 33384 800 33416
rect 840 33384 872 33416
rect 912 33384 944 33416
rect 984 33384 1016 33416
rect 1056 33384 1088 33416
rect 1128 33384 1160 33416
rect 1200 33384 1232 33416
rect 1272 33384 1304 33416
rect 1344 33384 1376 33416
rect 1416 33384 1448 33416
rect 1488 33384 1520 33416
rect 1560 33384 1592 33416
rect 1632 33384 1664 33416
rect 1704 33384 1736 33416
rect 1776 33384 1808 33416
rect 1848 33384 1880 33416
rect 192 29684 224 29716
rect 264 29684 296 29716
rect 336 29684 368 29716
rect 408 29684 440 29716
rect 480 29684 512 29716
rect 552 29684 584 29716
rect 624 29684 656 29716
rect 696 29684 728 29716
rect 768 29684 800 29716
rect 840 29684 872 29716
rect 912 29684 944 29716
rect 984 29684 1016 29716
rect 1056 29684 1088 29716
rect 1128 29684 1160 29716
rect 1200 29684 1232 29716
rect 1272 29684 1304 29716
rect 1344 29684 1376 29716
rect 1416 29684 1448 29716
rect 1488 29684 1520 29716
rect 1560 29684 1592 29716
rect 1632 29684 1664 29716
rect 1704 29684 1736 29716
rect 1776 29684 1808 29716
rect 1848 29684 1880 29716
rect 120 12112 152 12144
rect 192 12112 224 12144
rect 264 12112 296 12144
rect 336 12112 368 12144
rect 408 12112 440 12144
rect 480 12112 512 12144
rect 552 12112 584 12144
rect 624 12112 656 12144
rect 696 12112 728 12144
rect 768 12112 800 12144
rect 840 12112 872 12144
rect 912 12112 944 12144
rect 984 12112 1016 12144
rect 1056 12112 1088 12144
rect 1128 12112 1160 12144
rect 1200 12112 1232 12144
rect 1272 12112 1304 12144
rect 1344 12112 1376 12144
rect 1416 12112 1448 12144
rect 1488 12112 1520 12144
rect 1560 12112 1592 12144
rect 1632 12112 1664 12144
rect 1704 12112 1736 12144
rect 1776 12112 1808 12144
rect 1848 12112 1880 12144
rect 1920 12112 1952 12144
rect 48 12040 80 12072
rect 120 12040 152 12072
rect 192 12040 224 12072
rect 264 12040 296 12072
rect 336 12040 368 12072
rect 408 12040 440 12072
rect 480 12040 512 12072
rect 552 12040 584 12072
rect 624 12040 656 12072
rect 696 12040 728 12072
rect 768 12040 800 12072
rect 840 12040 872 12072
rect 912 12040 944 12072
rect 984 12040 1016 12072
rect 1056 12040 1088 12072
rect 1128 12040 1160 12072
rect 1200 12040 1232 12072
rect 1272 12040 1304 12072
rect 1344 12040 1376 12072
rect 1416 12040 1448 12072
rect 1488 12040 1520 12072
rect 1560 12040 1592 12072
rect 1632 12040 1664 12072
rect 1704 12040 1736 12072
rect 1776 12040 1808 12072
rect 1848 12040 1880 12072
rect 1920 12040 1952 12072
rect 48 11968 80 12000
rect 120 11968 152 12000
rect 192 11968 224 12000
rect 264 11968 296 12000
rect 336 11968 368 12000
rect 408 11968 440 12000
rect 480 11968 512 12000
rect 552 11968 584 12000
rect 624 11968 656 12000
rect 696 11968 728 12000
rect 768 11968 800 12000
rect 840 11968 872 12000
rect 912 11968 944 12000
rect 984 11968 1016 12000
rect 1056 11968 1088 12000
rect 1128 11968 1160 12000
rect 1200 11968 1232 12000
rect 1272 11968 1304 12000
rect 1344 11968 1376 12000
rect 1416 11968 1448 12000
rect 1488 11968 1520 12000
rect 1560 11968 1592 12000
rect 1632 11968 1664 12000
rect 1704 11968 1736 12000
rect 1776 11968 1808 12000
rect 1848 11968 1880 12000
rect 1920 11968 1952 12000
rect 48 11896 80 11928
rect 120 11896 152 11928
rect 192 11896 224 11928
rect 264 11896 296 11928
rect 336 11896 368 11928
rect 408 11896 440 11928
rect 480 11896 512 11928
rect 552 11896 584 11928
rect 624 11896 656 11928
rect 696 11896 728 11928
rect 768 11896 800 11928
rect 840 11896 872 11928
rect 912 11896 944 11928
rect 984 11896 1016 11928
rect 1056 11896 1088 11928
rect 1128 11896 1160 11928
rect 1200 11896 1232 11928
rect 1272 11896 1304 11928
rect 1344 11896 1376 11928
rect 1416 11896 1448 11928
rect 1488 11896 1520 11928
rect 1560 11896 1592 11928
rect 1632 11896 1664 11928
rect 1704 11896 1736 11928
rect 1776 11896 1808 11928
rect 1848 11896 1880 11928
rect 1920 11896 1952 11928
rect 48 11824 80 11856
rect 120 11824 152 11856
rect 192 11824 224 11856
rect 264 11824 296 11856
rect 336 11824 368 11856
rect 408 11824 440 11856
rect 480 11824 512 11856
rect 552 11824 584 11856
rect 624 11824 656 11856
rect 696 11824 728 11856
rect 768 11824 800 11856
rect 840 11824 872 11856
rect 912 11824 944 11856
rect 984 11824 1016 11856
rect 1056 11824 1088 11856
rect 1128 11824 1160 11856
rect 1200 11824 1232 11856
rect 1272 11824 1304 11856
rect 1344 11824 1376 11856
rect 1416 11824 1448 11856
rect 1488 11824 1520 11856
rect 1560 11824 1592 11856
rect 1632 11824 1664 11856
rect 1704 11824 1736 11856
rect 1776 11824 1808 11856
rect 1848 11824 1880 11856
rect 1920 11824 1952 11856
rect 48 11752 80 11784
rect 120 11752 152 11784
rect 192 11752 224 11784
rect 264 11752 296 11784
rect 336 11752 368 11784
rect 408 11752 440 11784
rect 480 11752 512 11784
rect 552 11752 584 11784
rect 624 11752 656 11784
rect 696 11752 728 11784
rect 768 11752 800 11784
rect 840 11752 872 11784
rect 912 11752 944 11784
rect 984 11752 1016 11784
rect 1056 11752 1088 11784
rect 1128 11752 1160 11784
rect 1200 11752 1232 11784
rect 1272 11752 1304 11784
rect 1344 11752 1376 11784
rect 1416 11752 1448 11784
rect 1488 11752 1520 11784
rect 1560 11752 1592 11784
rect 1632 11752 1664 11784
rect 1704 11752 1736 11784
rect 1776 11752 1808 11784
rect 1848 11752 1880 11784
rect 1920 11752 1952 11784
rect 48 11680 80 11712
rect 120 11680 152 11712
rect 192 11680 224 11712
rect 264 11680 296 11712
rect 336 11680 368 11712
rect 408 11680 440 11712
rect 480 11680 512 11712
rect 552 11680 584 11712
rect 624 11680 656 11712
rect 696 11680 728 11712
rect 768 11680 800 11712
rect 840 11680 872 11712
rect 912 11680 944 11712
rect 984 11680 1016 11712
rect 1056 11680 1088 11712
rect 1128 11680 1160 11712
rect 1200 11680 1232 11712
rect 1272 11680 1304 11712
rect 1344 11680 1376 11712
rect 1416 11680 1448 11712
rect 1488 11680 1520 11712
rect 1560 11680 1592 11712
rect 1632 11680 1664 11712
rect 1704 11680 1736 11712
rect 1776 11680 1808 11712
rect 1848 11680 1880 11712
rect 1920 11680 1952 11712
rect 48 11608 80 11640
rect 120 11608 152 11640
rect 192 11608 224 11640
rect 264 11608 296 11640
rect 336 11608 368 11640
rect 408 11608 440 11640
rect 480 11608 512 11640
rect 552 11608 584 11640
rect 624 11608 656 11640
rect 696 11608 728 11640
rect 768 11608 800 11640
rect 840 11608 872 11640
rect 912 11608 944 11640
rect 984 11608 1016 11640
rect 1056 11608 1088 11640
rect 1128 11608 1160 11640
rect 1200 11608 1232 11640
rect 1272 11608 1304 11640
rect 1344 11608 1376 11640
rect 1416 11608 1448 11640
rect 1488 11608 1520 11640
rect 1560 11608 1592 11640
rect 1632 11608 1664 11640
rect 1704 11608 1736 11640
rect 1776 11608 1808 11640
rect 1848 11608 1880 11640
rect 1920 11608 1952 11640
rect 48 11536 80 11568
rect 120 11536 152 11568
rect 192 11536 224 11568
rect 264 11536 296 11568
rect 336 11536 368 11568
rect 408 11536 440 11568
rect 480 11536 512 11568
rect 552 11536 584 11568
rect 624 11536 656 11568
rect 696 11536 728 11568
rect 768 11536 800 11568
rect 840 11536 872 11568
rect 912 11536 944 11568
rect 984 11536 1016 11568
rect 1056 11536 1088 11568
rect 1128 11536 1160 11568
rect 1200 11536 1232 11568
rect 1272 11536 1304 11568
rect 1344 11536 1376 11568
rect 1416 11536 1448 11568
rect 1488 11536 1520 11568
rect 1560 11536 1592 11568
rect 1632 11536 1664 11568
rect 1704 11536 1736 11568
rect 1776 11536 1808 11568
rect 1848 11536 1880 11568
rect 1920 11536 1952 11568
rect 48 11464 80 11496
rect 120 11464 152 11496
rect 192 11464 224 11496
rect 264 11464 296 11496
rect 336 11464 368 11496
rect 408 11464 440 11496
rect 480 11464 512 11496
rect 552 11464 584 11496
rect 624 11464 656 11496
rect 696 11464 728 11496
rect 768 11464 800 11496
rect 840 11464 872 11496
rect 912 11464 944 11496
rect 984 11464 1016 11496
rect 1056 11464 1088 11496
rect 1128 11464 1160 11496
rect 1200 11464 1232 11496
rect 1272 11464 1304 11496
rect 1344 11464 1376 11496
rect 1416 11464 1448 11496
rect 1488 11464 1520 11496
rect 1560 11464 1592 11496
rect 1632 11464 1664 11496
rect 1704 11464 1736 11496
rect 1776 11464 1808 11496
rect 1848 11464 1880 11496
rect 1920 11464 1952 11496
rect 48 11392 80 11424
rect 120 11392 152 11424
rect 192 11392 224 11424
rect 264 11392 296 11424
rect 336 11392 368 11424
rect 408 11392 440 11424
rect 480 11392 512 11424
rect 552 11392 584 11424
rect 624 11392 656 11424
rect 696 11392 728 11424
rect 768 11392 800 11424
rect 840 11392 872 11424
rect 912 11392 944 11424
rect 984 11392 1016 11424
rect 1056 11392 1088 11424
rect 1128 11392 1160 11424
rect 1200 11392 1232 11424
rect 1272 11392 1304 11424
rect 1344 11392 1376 11424
rect 1416 11392 1448 11424
rect 1488 11392 1520 11424
rect 1560 11392 1592 11424
rect 1632 11392 1664 11424
rect 1704 11392 1736 11424
rect 1776 11392 1808 11424
rect 1848 11392 1880 11424
rect 1920 11392 1952 11424
rect 48 11320 80 11352
rect 120 11320 152 11352
rect 192 11320 224 11352
rect 264 11320 296 11352
rect 336 11320 368 11352
rect 408 11320 440 11352
rect 480 11320 512 11352
rect 552 11320 584 11352
rect 624 11320 656 11352
rect 696 11320 728 11352
rect 768 11320 800 11352
rect 840 11320 872 11352
rect 912 11320 944 11352
rect 984 11320 1016 11352
rect 1056 11320 1088 11352
rect 1128 11320 1160 11352
rect 1200 11320 1232 11352
rect 1272 11320 1304 11352
rect 1344 11320 1376 11352
rect 1416 11320 1448 11352
rect 1488 11320 1520 11352
rect 1560 11320 1592 11352
rect 1632 11320 1664 11352
rect 1704 11320 1736 11352
rect 1776 11320 1808 11352
rect 1848 11320 1880 11352
rect 1920 11320 1952 11352
rect 48 11248 80 11280
rect 120 11248 152 11280
rect 192 11248 224 11280
rect 264 11248 296 11280
rect 336 11248 368 11280
rect 408 11248 440 11280
rect 480 11248 512 11280
rect 552 11248 584 11280
rect 624 11248 656 11280
rect 696 11248 728 11280
rect 768 11248 800 11280
rect 840 11248 872 11280
rect 912 11248 944 11280
rect 984 11248 1016 11280
rect 1056 11248 1088 11280
rect 1128 11248 1160 11280
rect 1200 11248 1232 11280
rect 1272 11248 1304 11280
rect 1344 11248 1376 11280
rect 1416 11248 1448 11280
rect 1488 11248 1520 11280
rect 1560 11248 1592 11280
rect 1632 11248 1664 11280
rect 1704 11248 1736 11280
rect 1776 11248 1808 11280
rect 1848 11248 1880 11280
rect 1920 11248 1952 11280
rect 48 11176 80 11208
rect 120 11176 152 11208
rect 192 11176 224 11208
rect 264 11176 296 11208
rect 336 11176 368 11208
rect 408 11176 440 11208
rect 480 11176 512 11208
rect 552 11176 584 11208
rect 624 11176 656 11208
rect 696 11176 728 11208
rect 768 11176 800 11208
rect 840 11176 872 11208
rect 912 11176 944 11208
rect 984 11176 1016 11208
rect 1056 11176 1088 11208
rect 1128 11176 1160 11208
rect 1200 11176 1232 11208
rect 1272 11176 1304 11208
rect 1344 11176 1376 11208
rect 1416 11176 1448 11208
rect 1488 11176 1520 11208
rect 1560 11176 1592 11208
rect 1632 11176 1664 11208
rect 1704 11176 1736 11208
rect 1776 11176 1808 11208
rect 1848 11176 1880 11208
rect 1920 11176 1952 11208
rect 48 11104 80 11136
rect 120 11104 152 11136
rect 192 11104 224 11136
rect 264 11104 296 11136
rect 336 11104 368 11136
rect 408 11104 440 11136
rect 480 11104 512 11136
rect 552 11104 584 11136
rect 624 11104 656 11136
rect 696 11104 728 11136
rect 768 11104 800 11136
rect 840 11104 872 11136
rect 912 11104 944 11136
rect 984 11104 1016 11136
rect 1056 11104 1088 11136
rect 1128 11104 1160 11136
rect 1200 11104 1232 11136
rect 1272 11104 1304 11136
rect 1344 11104 1376 11136
rect 1416 11104 1448 11136
rect 1488 11104 1520 11136
rect 1560 11104 1592 11136
rect 1632 11104 1664 11136
rect 1704 11104 1736 11136
rect 1776 11104 1808 11136
rect 1848 11104 1880 11136
rect 1920 11104 1952 11136
rect 48 11032 80 11064
rect 120 11032 152 11064
rect 192 11032 224 11064
rect 264 11032 296 11064
rect 336 11032 368 11064
rect 408 11032 440 11064
rect 480 11032 512 11064
rect 552 11032 584 11064
rect 624 11032 656 11064
rect 696 11032 728 11064
rect 768 11032 800 11064
rect 840 11032 872 11064
rect 912 11032 944 11064
rect 984 11032 1016 11064
rect 1056 11032 1088 11064
rect 1128 11032 1160 11064
rect 1200 11032 1232 11064
rect 1272 11032 1304 11064
rect 1344 11032 1376 11064
rect 1416 11032 1448 11064
rect 1488 11032 1520 11064
rect 1560 11032 1592 11064
rect 1632 11032 1664 11064
rect 1704 11032 1736 11064
rect 1776 11032 1808 11064
rect 1848 11032 1880 11064
rect 1920 11032 1952 11064
rect 48 10960 80 10992
rect 120 10960 152 10992
rect 192 10960 224 10992
rect 264 10960 296 10992
rect 336 10960 368 10992
rect 408 10960 440 10992
rect 480 10960 512 10992
rect 552 10960 584 10992
rect 624 10960 656 10992
rect 696 10960 728 10992
rect 768 10960 800 10992
rect 840 10960 872 10992
rect 912 10960 944 10992
rect 984 10960 1016 10992
rect 1056 10960 1088 10992
rect 1128 10960 1160 10992
rect 1200 10960 1232 10992
rect 1272 10960 1304 10992
rect 1344 10960 1376 10992
rect 1416 10960 1448 10992
rect 1488 10960 1520 10992
rect 1560 10960 1592 10992
rect 1632 10960 1664 10992
rect 1704 10960 1736 10992
rect 1776 10960 1808 10992
rect 1848 10960 1880 10992
rect 1920 10960 1952 10992
rect 48 10888 80 10920
rect 120 10888 152 10920
rect 192 10888 224 10920
rect 264 10888 296 10920
rect 336 10888 368 10920
rect 408 10888 440 10920
rect 480 10888 512 10920
rect 552 10888 584 10920
rect 624 10888 656 10920
rect 696 10888 728 10920
rect 768 10888 800 10920
rect 840 10888 872 10920
rect 912 10888 944 10920
rect 984 10888 1016 10920
rect 1056 10888 1088 10920
rect 1128 10888 1160 10920
rect 1200 10888 1232 10920
rect 1272 10888 1304 10920
rect 1344 10888 1376 10920
rect 1416 10888 1448 10920
rect 1488 10888 1520 10920
rect 1560 10888 1592 10920
rect 1632 10888 1664 10920
rect 1704 10888 1736 10920
rect 1776 10888 1808 10920
rect 1848 10888 1880 10920
rect 1920 10888 1952 10920
rect 48 10816 80 10848
rect 120 10816 152 10848
rect 192 10816 224 10848
rect 264 10816 296 10848
rect 336 10816 368 10848
rect 408 10816 440 10848
rect 480 10816 512 10848
rect 552 10816 584 10848
rect 624 10816 656 10848
rect 696 10816 728 10848
rect 768 10816 800 10848
rect 840 10816 872 10848
rect 912 10816 944 10848
rect 984 10816 1016 10848
rect 1056 10816 1088 10848
rect 1128 10816 1160 10848
rect 1200 10816 1232 10848
rect 1272 10816 1304 10848
rect 1344 10816 1376 10848
rect 1416 10816 1448 10848
rect 1488 10816 1520 10848
rect 1560 10816 1592 10848
rect 1632 10816 1664 10848
rect 1704 10816 1736 10848
rect 1776 10816 1808 10848
rect 1848 10816 1880 10848
rect 1920 10816 1952 10848
rect 48 10744 80 10776
rect 120 10744 152 10776
rect 192 10744 224 10776
rect 264 10744 296 10776
rect 336 10744 368 10776
rect 408 10744 440 10776
rect 480 10744 512 10776
rect 552 10744 584 10776
rect 624 10744 656 10776
rect 696 10744 728 10776
rect 768 10744 800 10776
rect 840 10744 872 10776
rect 912 10744 944 10776
rect 984 10744 1016 10776
rect 1056 10744 1088 10776
rect 1128 10744 1160 10776
rect 1200 10744 1232 10776
rect 1272 10744 1304 10776
rect 1344 10744 1376 10776
rect 1416 10744 1448 10776
rect 1488 10744 1520 10776
rect 1560 10744 1592 10776
rect 1632 10744 1664 10776
rect 1704 10744 1736 10776
rect 1776 10744 1808 10776
rect 1848 10744 1880 10776
rect 1920 10744 1952 10776
rect 48 10672 80 10704
rect 120 10672 152 10704
rect 192 10672 224 10704
rect 264 10672 296 10704
rect 336 10672 368 10704
rect 408 10672 440 10704
rect 480 10672 512 10704
rect 552 10672 584 10704
rect 624 10672 656 10704
rect 696 10672 728 10704
rect 768 10672 800 10704
rect 840 10672 872 10704
rect 912 10672 944 10704
rect 984 10672 1016 10704
rect 1056 10672 1088 10704
rect 1128 10672 1160 10704
rect 1200 10672 1232 10704
rect 1272 10672 1304 10704
rect 1344 10672 1376 10704
rect 1416 10672 1448 10704
rect 1488 10672 1520 10704
rect 1560 10672 1592 10704
rect 1632 10672 1664 10704
rect 1704 10672 1736 10704
rect 1776 10672 1808 10704
rect 1848 10672 1880 10704
rect 1920 10672 1952 10704
rect 48 10600 80 10632
rect 120 10600 152 10632
rect 192 10600 224 10632
rect 264 10600 296 10632
rect 336 10600 368 10632
rect 408 10600 440 10632
rect 480 10600 512 10632
rect 552 10600 584 10632
rect 624 10600 656 10632
rect 696 10600 728 10632
rect 768 10600 800 10632
rect 840 10600 872 10632
rect 912 10600 944 10632
rect 984 10600 1016 10632
rect 1056 10600 1088 10632
rect 1128 10600 1160 10632
rect 1200 10600 1232 10632
rect 1272 10600 1304 10632
rect 1344 10600 1376 10632
rect 1416 10600 1448 10632
rect 1488 10600 1520 10632
rect 1560 10600 1592 10632
rect 1632 10600 1664 10632
rect 1704 10600 1736 10632
rect 1776 10600 1808 10632
rect 1848 10600 1880 10632
rect 1920 10600 1952 10632
rect 48 10528 80 10560
rect 120 10528 152 10560
rect 192 10528 224 10560
rect 264 10528 296 10560
rect 336 10528 368 10560
rect 408 10528 440 10560
rect 480 10528 512 10560
rect 552 10528 584 10560
rect 624 10528 656 10560
rect 696 10528 728 10560
rect 768 10528 800 10560
rect 840 10528 872 10560
rect 912 10528 944 10560
rect 984 10528 1016 10560
rect 1056 10528 1088 10560
rect 1128 10528 1160 10560
rect 1200 10528 1232 10560
rect 1272 10528 1304 10560
rect 1344 10528 1376 10560
rect 1416 10528 1448 10560
rect 1488 10528 1520 10560
rect 1560 10528 1592 10560
rect 1632 10528 1664 10560
rect 1704 10528 1736 10560
rect 1776 10528 1808 10560
rect 1848 10528 1880 10560
rect 1920 10528 1952 10560
rect 48 10456 80 10488
rect 120 10456 152 10488
rect 192 10456 224 10488
rect 264 10456 296 10488
rect 336 10456 368 10488
rect 408 10456 440 10488
rect 480 10456 512 10488
rect 552 10456 584 10488
rect 624 10456 656 10488
rect 696 10456 728 10488
rect 768 10456 800 10488
rect 840 10456 872 10488
rect 912 10456 944 10488
rect 984 10456 1016 10488
rect 1056 10456 1088 10488
rect 1128 10456 1160 10488
rect 1200 10456 1232 10488
rect 1272 10456 1304 10488
rect 1344 10456 1376 10488
rect 1416 10456 1448 10488
rect 1488 10456 1520 10488
rect 1560 10456 1592 10488
rect 1632 10456 1664 10488
rect 1704 10456 1736 10488
rect 1776 10456 1808 10488
rect 1848 10456 1880 10488
rect 1920 10456 1952 10488
rect 48 10384 80 10416
rect 120 10384 152 10416
rect 192 10384 224 10416
rect 264 10384 296 10416
rect 336 10384 368 10416
rect 408 10384 440 10416
rect 480 10384 512 10416
rect 552 10384 584 10416
rect 624 10384 656 10416
rect 696 10384 728 10416
rect 768 10384 800 10416
rect 840 10384 872 10416
rect 912 10384 944 10416
rect 984 10384 1016 10416
rect 1056 10384 1088 10416
rect 1128 10384 1160 10416
rect 1200 10384 1232 10416
rect 1272 10384 1304 10416
rect 1344 10384 1376 10416
rect 1416 10384 1448 10416
rect 1488 10384 1520 10416
rect 1560 10384 1592 10416
rect 1632 10384 1664 10416
rect 1704 10384 1736 10416
rect 1776 10384 1808 10416
rect 1848 10384 1880 10416
rect 1920 10384 1952 10416
rect 48 10312 80 10344
rect 120 10312 152 10344
rect 192 10312 224 10344
rect 264 10312 296 10344
rect 336 10312 368 10344
rect 408 10312 440 10344
rect 480 10312 512 10344
rect 552 10312 584 10344
rect 624 10312 656 10344
rect 696 10312 728 10344
rect 768 10312 800 10344
rect 840 10312 872 10344
rect 912 10312 944 10344
rect 984 10312 1016 10344
rect 1056 10312 1088 10344
rect 1128 10312 1160 10344
rect 1200 10312 1232 10344
rect 1272 10312 1304 10344
rect 1344 10312 1376 10344
rect 1416 10312 1448 10344
rect 1488 10312 1520 10344
rect 1560 10312 1592 10344
rect 1632 10312 1664 10344
rect 1704 10312 1736 10344
rect 1776 10312 1808 10344
rect 1848 10312 1880 10344
rect 1920 10312 1952 10344
rect 48 10240 80 10272
rect 120 10240 152 10272
rect 192 10240 224 10272
rect 264 10240 296 10272
rect 336 10240 368 10272
rect 408 10240 440 10272
rect 480 10240 512 10272
rect 552 10240 584 10272
rect 624 10240 656 10272
rect 696 10240 728 10272
rect 768 10240 800 10272
rect 840 10240 872 10272
rect 912 10240 944 10272
rect 984 10240 1016 10272
rect 1056 10240 1088 10272
rect 1128 10240 1160 10272
rect 1200 10240 1232 10272
rect 1272 10240 1304 10272
rect 1344 10240 1376 10272
rect 1416 10240 1448 10272
rect 1488 10240 1520 10272
rect 1560 10240 1592 10272
rect 1632 10240 1664 10272
rect 1704 10240 1736 10272
rect 1776 10240 1808 10272
rect 1848 10240 1880 10272
rect 1920 10240 1952 10272
rect 48 10168 80 10200
rect 120 10168 152 10200
rect 192 10168 224 10200
rect 264 10168 296 10200
rect 336 10168 368 10200
rect 408 10168 440 10200
rect 480 10168 512 10200
rect 552 10168 584 10200
rect 624 10168 656 10200
rect 696 10168 728 10200
rect 768 10168 800 10200
rect 840 10168 872 10200
rect 912 10168 944 10200
rect 984 10168 1016 10200
rect 1056 10168 1088 10200
rect 1128 10168 1160 10200
rect 1200 10168 1232 10200
rect 1272 10168 1304 10200
rect 1344 10168 1376 10200
rect 1416 10168 1448 10200
rect 1488 10168 1520 10200
rect 1560 10168 1592 10200
rect 1632 10168 1664 10200
rect 1704 10168 1736 10200
rect 1776 10168 1808 10200
rect 1848 10168 1880 10200
rect 1920 10168 1952 10200
rect 48 10096 80 10128
rect 120 10096 152 10128
rect 192 10096 224 10128
rect 264 10096 296 10128
rect 336 10096 368 10128
rect 408 10096 440 10128
rect 480 10096 512 10128
rect 552 10096 584 10128
rect 624 10096 656 10128
rect 696 10096 728 10128
rect 768 10096 800 10128
rect 840 10096 872 10128
rect 912 10096 944 10128
rect 984 10096 1016 10128
rect 1056 10096 1088 10128
rect 1128 10096 1160 10128
rect 1200 10096 1232 10128
rect 1272 10096 1304 10128
rect 1344 10096 1376 10128
rect 1416 10096 1448 10128
rect 1488 10096 1520 10128
rect 1560 10096 1592 10128
rect 1632 10096 1664 10128
rect 1704 10096 1736 10128
rect 1776 10096 1808 10128
rect 1848 10096 1880 10128
rect 1920 10096 1952 10128
rect 48 10024 80 10056
rect 120 10024 152 10056
rect 192 10024 224 10056
rect 264 10024 296 10056
rect 336 10024 368 10056
rect 408 10024 440 10056
rect 480 10024 512 10056
rect 552 10024 584 10056
rect 624 10024 656 10056
rect 696 10024 728 10056
rect 768 10024 800 10056
rect 840 10024 872 10056
rect 912 10024 944 10056
rect 984 10024 1016 10056
rect 1056 10024 1088 10056
rect 1128 10024 1160 10056
rect 1200 10024 1232 10056
rect 1272 10024 1304 10056
rect 1344 10024 1376 10056
rect 1416 10024 1448 10056
rect 1488 10024 1520 10056
rect 1560 10024 1592 10056
rect 1632 10024 1664 10056
rect 1704 10024 1736 10056
rect 1776 10024 1808 10056
rect 1848 10024 1880 10056
rect 1920 10024 1952 10056
rect 48 9952 80 9984
rect 120 9952 152 9984
rect 192 9952 224 9984
rect 264 9952 296 9984
rect 336 9952 368 9984
rect 408 9952 440 9984
rect 480 9952 512 9984
rect 552 9952 584 9984
rect 624 9952 656 9984
rect 696 9952 728 9984
rect 768 9952 800 9984
rect 840 9952 872 9984
rect 912 9952 944 9984
rect 984 9952 1016 9984
rect 1056 9952 1088 9984
rect 1128 9952 1160 9984
rect 1200 9952 1232 9984
rect 1272 9952 1304 9984
rect 1344 9952 1376 9984
rect 1416 9952 1448 9984
rect 1488 9952 1520 9984
rect 1560 9952 1592 9984
rect 1632 9952 1664 9984
rect 1704 9952 1736 9984
rect 1776 9952 1808 9984
rect 1848 9952 1880 9984
rect 1920 9952 1952 9984
rect 48 9880 80 9912
rect 120 9880 152 9912
rect 192 9880 224 9912
rect 264 9880 296 9912
rect 336 9880 368 9912
rect 408 9880 440 9912
rect 480 9880 512 9912
rect 552 9880 584 9912
rect 624 9880 656 9912
rect 696 9880 728 9912
rect 768 9880 800 9912
rect 840 9880 872 9912
rect 912 9880 944 9912
rect 984 9880 1016 9912
rect 1056 9880 1088 9912
rect 1128 9880 1160 9912
rect 1200 9880 1232 9912
rect 1272 9880 1304 9912
rect 1344 9880 1376 9912
rect 1416 9880 1448 9912
rect 1488 9880 1520 9912
rect 1560 9880 1592 9912
rect 1632 9880 1664 9912
rect 1704 9880 1736 9912
rect 1776 9880 1808 9912
rect 1848 9880 1880 9912
rect 1920 9880 1952 9912
rect 48 9808 80 9840
rect 120 9808 152 9840
rect 192 9808 224 9840
rect 264 9808 296 9840
rect 336 9808 368 9840
rect 408 9808 440 9840
rect 480 9808 512 9840
rect 552 9808 584 9840
rect 624 9808 656 9840
rect 696 9808 728 9840
rect 768 9808 800 9840
rect 840 9808 872 9840
rect 912 9808 944 9840
rect 984 9808 1016 9840
rect 1056 9808 1088 9840
rect 1128 9808 1160 9840
rect 1200 9808 1232 9840
rect 1272 9808 1304 9840
rect 1344 9808 1376 9840
rect 1416 9808 1448 9840
rect 1488 9808 1520 9840
rect 1560 9808 1592 9840
rect 1632 9808 1664 9840
rect 1704 9808 1736 9840
rect 1776 9808 1808 9840
rect 1848 9808 1880 9840
rect 1920 9808 1952 9840
rect 48 9736 80 9768
rect 120 9736 152 9768
rect 192 9736 224 9768
rect 264 9736 296 9768
rect 336 9736 368 9768
rect 408 9736 440 9768
rect 480 9736 512 9768
rect 552 9736 584 9768
rect 624 9736 656 9768
rect 696 9736 728 9768
rect 768 9736 800 9768
rect 840 9736 872 9768
rect 912 9736 944 9768
rect 984 9736 1016 9768
rect 1056 9736 1088 9768
rect 1128 9736 1160 9768
rect 1200 9736 1232 9768
rect 1272 9736 1304 9768
rect 1344 9736 1376 9768
rect 1416 9736 1448 9768
rect 1488 9736 1520 9768
rect 1560 9736 1592 9768
rect 1632 9736 1664 9768
rect 1704 9736 1736 9768
rect 1776 9736 1808 9768
rect 1848 9736 1880 9768
rect 1920 9736 1952 9768
rect 48 9664 80 9696
rect 120 9664 152 9696
rect 192 9664 224 9696
rect 264 9664 296 9696
rect 336 9664 368 9696
rect 408 9664 440 9696
rect 480 9664 512 9696
rect 552 9664 584 9696
rect 624 9664 656 9696
rect 696 9664 728 9696
rect 768 9664 800 9696
rect 840 9664 872 9696
rect 912 9664 944 9696
rect 984 9664 1016 9696
rect 1056 9664 1088 9696
rect 1128 9664 1160 9696
rect 1200 9664 1232 9696
rect 1272 9664 1304 9696
rect 1344 9664 1376 9696
rect 1416 9664 1448 9696
rect 1488 9664 1520 9696
rect 1560 9664 1592 9696
rect 1632 9664 1664 9696
rect 1704 9664 1736 9696
rect 1776 9664 1808 9696
rect 1848 9664 1880 9696
rect 1920 9664 1952 9696
rect 48 9592 80 9624
rect 120 9592 152 9624
rect 192 9592 224 9624
rect 264 9592 296 9624
rect 336 9592 368 9624
rect 408 9592 440 9624
rect 480 9592 512 9624
rect 552 9592 584 9624
rect 624 9592 656 9624
rect 696 9592 728 9624
rect 768 9592 800 9624
rect 840 9592 872 9624
rect 912 9592 944 9624
rect 984 9592 1016 9624
rect 1056 9592 1088 9624
rect 1128 9592 1160 9624
rect 1200 9592 1232 9624
rect 1272 9592 1304 9624
rect 1344 9592 1376 9624
rect 1416 9592 1448 9624
rect 1488 9592 1520 9624
rect 1560 9592 1592 9624
rect 1632 9592 1664 9624
rect 1704 9592 1736 9624
rect 1776 9592 1808 9624
rect 1848 9592 1880 9624
rect 1920 9592 1952 9624
rect 48 9520 80 9552
rect 120 9520 152 9552
rect 192 9520 224 9552
rect 264 9520 296 9552
rect 336 9520 368 9552
rect 408 9520 440 9552
rect 480 9520 512 9552
rect 552 9520 584 9552
rect 624 9520 656 9552
rect 696 9520 728 9552
rect 768 9520 800 9552
rect 840 9520 872 9552
rect 912 9520 944 9552
rect 984 9520 1016 9552
rect 1056 9520 1088 9552
rect 1128 9520 1160 9552
rect 1200 9520 1232 9552
rect 1272 9520 1304 9552
rect 1344 9520 1376 9552
rect 1416 9520 1448 9552
rect 1488 9520 1520 9552
rect 1560 9520 1592 9552
rect 1632 9520 1664 9552
rect 1704 9520 1736 9552
rect 1776 9520 1808 9552
rect 1848 9520 1880 9552
rect 1920 9520 1952 9552
rect 48 9448 80 9480
rect 120 9448 152 9480
rect 192 9448 224 9480
rect 264 9448 296 9480
rect 336 9448 368 9480
rect 408 9448 440 9480
rect 480 9448 512 9480
rect 552 9448 584 9480
rect 624 9448 656 9480
rect 696 9448 728 9480
rect 768 9448 800 9480
rect 840 9448 872 9480
rect 912 9448 944 9480
rect 984 9448 1016 9480
rect 1056 9448 1088 9480
rect 1128 9448 1160 9480
rect 1200 9448 1232 9480
rect 1272 9448 1304 9480
rect 1344 9448 1376 9480
rect 1416 9448 1448 9480
rect 1488 9448 1520 9480
rect 1560 9448 1592 9480
rect 1632 9448 1664 9480
rect 1704 9448 1736 9480
rect 1776 9448 1808 9480
rect 1848 9448 1880 9480
rect 1920 9448 1952 9480
rect 48 9376 80 9408
rect 120 9376 152 9408
rect 192 9376 224 9408
rect 264 9376 296 9408
rect 336 9376 368 9408
rect 408 9376 440 9408
rect 480 9376 512 9408
rect 552 9376 584 9408
rect 624 9376 656 9408
rect 696 9376 728 9408
rect 768 9376 800 9408
rect 840 9376 872 9408
rect 912 9376 944 9408
rect 984 9376 1016 9408
rect 1056 9376 1088 9408
rect 1128 9376 1160 9408
rect 1200 9376 1232 9408
rect 1272 9376 1304 9408
rect 1344 9376 1376 9408
rect 1416 9376 1448 9408
rect 1488 9376 1520 9408
rect 1560 9376 1592 9408
rect 1632 9376 1664 9408
rect 1704 9376 1736 9408
rect 1776 9376 1808 9408
rect 1848 9376 1880 9408
rect 1920 9376 1952 9408
rect 48 9304 80 9336
rect 120 9304 152 9336
rect 192 9304 224 9336
rect 264 9304 296 9336
rect 336 9304 368 9336
rect 408 9304 440 9336
rect 480 9304 512 9336
rect 552 9304 584 9336
rect 624 9304 656 9336
rect 696 9304 728 9336
rect 768 9304 800 9336
rect 840 9304 872 9336
rect 912 9304 944 9336
rect 984 9304 1016 9336
rect 1056 9304 1088 9336
rect 1128 9304 1160 9336
rect 1200 9304 1232 9336
rect 1272 9304 1304 9336
rect 1344 9304 1376 9336
rect 1416 9304 1448 9336
rect 1488 9304 1520 9336
rect 1560 9304 1592 9336
rect 1632 9304 1664 9336
rect 1704 9304 1736 9336
rect 1776 9304 1808 9336
rect 1848 9304 1880 9336
rect 1920 9304 1952 9336
rect 48 9232 80 9264
rect 120 9232 152 9264
rect 192 9232 224 9264
rect 264 9232 296 9264
rect 336 9232 368 9264
rect 408 9232 440 9264
rect 480 9232 512 9264
rect 552 9232 584 9264
rect 624 9232 656 9264
rect 696 9232 728 9264
rect 768 9232 800 9264
rect 840 9232 872 9264
rect 912 9232 944 9264
rect 984 9232 1016 9264
rect 1056 9232 1088 9264
rect 1128 9232 1160 9264
rect 1200 9232 1232 9264
rect 1272 9232 1304 9264
rect 1344 9232 1376 9264
rect 1416 9232 1448 9264
rect 1488 9232 1520 9264
rect 1560 9232 1592 9264
rect 1632 9232 1664 9264
rect 1704 9232 1736 9264
rect 1776 9232 1808 9264
rect 1848 9232 1880 9264
rect 1920 9232 1952 9264
rect 48 9160 80 9192
rect 120 9160 152 9192
rect 192 9160 224 9192
rect 264 9160 296 9192
rect 336 9160 368 9192
rect 408 9160 440 9192
rect 480 9160 512 9192
rect 552 9160 584 9192
rect 624 9160 656 9192
rect 696 9160 728 9192
rect 768 9160 800 9192
rect 840 9160 872 9192
rect 912 9160 944 9192
rect 984 9160 1016 9192
rect 1056 9160 1088 9192
rect 1128 9160 1160 9192
rect 1200 9160 1232 9192
rect 1272 9160 1304 9192
rect 1344 9160 1376 9192
rect 1416 9160 1448 9192
rect 1488 9160 1520 9192
rect 1560 9160 1592 9192
rect 1632 9160 1664 9192
rect 1704 9160 1736 9192
rect 1776 9160 1808 9192
rect 1848 9160 1880 9192
rect 1920 9160 1952 9192
rect 48 9088 80 9120
rect 120 9088 152 9120
rect 192 9088 224 9120
rect 264 9088 296 9120
rect 336 9088 368 9120
rect 408 9088 440 9120
rect 480 9088 512 9120
rect 552 9088 584 9120
rect 624 9088 656 9120
rect 696 9088 728 9120
rect 768 9088 800 9120
rect 840 9088 872 9120
rect 912 9088 944 9120
rect 984 9088 1016 9120
rect 1056 9088 1088 9120
rect 1128 9088 1160 9120
rect 1200 9088 1232 9120
rect 1272 9088 1304 9120
rect 1344 9088 1376 9120
rect 1416 9088 1448 9120
rect 1488 9088 1520 9120
rect 1560 9088 1592 9120
rect 1632 9088 1664 9120
rect 1704 9088 1736 9120
rect 1776 9088 1808 9120
rect 1848 9088 1880 9120
rect 1920 9088 1952 9120
rect 48 9016 80 9048
rect 120 9016 152 9048
rect 192 9016 224 9048
rect 264 9016 296 9048
rect 336 9016 368 9048
rect 408 9016 440 9048
rect 480 9016 512 9048
rect 552 9016 584 9048
rect 624 9016 656 9048
rect 696 9016 728 9048
rect 768 9016 800 9048
rect 840 9016 872 9048
rect 912 9016 944 9048
rect 984 9016 1016 9048
rect 1056 9016 1088 9048
rect 1128 9016 1160 9048
rect 1200 9016 1232 9048
rect 1272 9016 1304 9048
rect 1344 9016 1376 9048
rect 1416 9016 1448 9048
rect 1488 9016 1520 9048
rect 1560 9016 1592 9048
rect 1632 9016 1664 9048
rect 1704 9016 1736 9048
rect 1776 9016 1808 9048
rect 1848 9016 1880 9048
rect 1920 9016 1952 9048
rect 48 8944 80 8976
rect 120 8944 152 8976
rect 192 8944 224 8976
rect 264 8944 296 8976
rect 336 8944 368 8976
rect 408 8944 440 8976
rect 480 8944 512 8976
rect 552 8944 584 8976
rect 624 8944 656 8976
rect 696 8944 728 8976
rect 768 8944 800 8976
rect 840 8944 872 8976
rect 912 8944 944 8976
rect 984 8944 1016 8976
rect 1056 8944 1088 8976
rect 1128 8944 1160 8976
rect 1200 8944 1232 8976
rect 1272 8944 1304 8976
rect 1344 8944 1376 8976
rect 1416 8944 1448 8976
rect 1488 8944 1520 8976
rect 1560 8944 1592 8976
rect 1632 8944 1664 8976
rect 1704 8944 1736 8976
rect 1776 8944 1808 8976
rect 1848 8944 1880 8976
rect 1920 8944 1952 8976
rect 48 8872 80 8904
rect 120 8872 152 8904
rect 192 8872 224 8904
rect 264 8872 296 8904
rect 336 8872 368 8904
rect 408 8872 440 8904
rect 480 8872 512 8904
rect 552 8872 584 8904
rect 624 8872 656 8904
rect 696 8872 728 8904
rect 768 8872 800 8904
rect 840 8872 872 8904
rect 912 8872 944 8904
rect 984 8872 1016 8904
rect 1056 8872 1088 8904
rect 1128 8872 1160 8904
rect 1200 8872 1232 8904
rect 1272 8872 1304 8904
rect 1344 8872 1376 8904
rect 1416 8872 1448 8904
rect 1488 8872 1520 8904
rect 1560 8872 1592 8904
rect 1632 8872 1664 8904
rect 1704 8872 1736 8904
rect 1776 8872 1808 8904
rect 1848 8872 1880 8904
rect 1920 8872 1952 8904
rect 48 8800 80 8832
rect 120 8800 152 8832
rect 192 8800 224 8832
rect 264 8800 296 8832
rect 336 8800 368 8832
rect 408 8800 440 8832
rect 480 8800 512 8832
rect 552 8800 584 8832
rect 624 8800 656 8832
rect 696 8800 728 8832
rect 768 8800 800 8832
rect 840 8800 872 8832
rect 912 8800 944 8832
rect 984 8800 1016 8832
rect 1056 8800 1088 8832
rect 1128 8800 1160 8832
rect 1200 8800 1232 8832
rect 1272 8800 1304 8832
rect 1344 8800 1376 8832
rect 1416 8800 1448 8832
rect 1488 8800 1520 8832
rect 1560 8800 1592 8832
rect 1632 8800 1664 8832
rect 1704 8800 1736 8832
rect 1776 8800 1808 8832
rect 1848 8800 1880 8832
rect 1920 8800 1952 8832
rect 48 8728 80 8760
rect 120 8728 152 8760
rect 192 8728 224 8760
rect 264 8728 296 8760
rect 336 8728 368 8760
rect 408 8728 440 8760
rect 480 8728 512 8760
rect 552 8728 584 8760
rect 624 8728 656 8760
rect 696 8728 728 8760
rect 768 8728 800 8760
rect 840 8728 872 8760
rect 912 8728 944 8760
rect 984 8728 1016 8760
rect 1056 8728 1088 8760
rect 1128 8728 1160 8760
rect 1200 8728 1232 8760
rect 1272 8728 1304 8760
rect 1344 8728 1376 8760
rect 1416 8728 1448 8760
rect 1488 8728 1520 8760
rect 1560 8728 1592 8760
rect 1632 8728 1664 8760
rect 1704 8728 1736 8760
rect 1776 8728 1808 8760
rect 1848 8728 1880 8760
rect 1920 8728 1952 8760
rect 48 8656 80 8688
rect 120 8656 152 8688
rect 192 8656 224 8688
rect 264 8656 296 8688
rect 336 8656 368 8688
rect 408 8656 440 8688
rect 480 8656 512 8688
rect 552 8656 584 8688
rect 624 8656 656 8688
rect 696 8656 728 8688
rect 768 8656 800 8688
rect 840 8656 872 8688
rect 912 8656 944 8688
rect 984 8656 1016 8688
rect 1056 8656 1088 8688
rect 1128 8656 1160 8688
rect 1200 8656 1232 8688
rect 1272 8656 1304 8688
rect 1344 8656 1376 8688
rect 1416 8656 1448 8688
rect 1488 8656 1520 8688
rect 1560 8656 1592 8688
rect 1632 8656 1664 8688
rect 1704 8656 1736 8688
rect 1776 8656 1808 8688
rect 1848 8656 1880 8688
rect 1920 8656 1952 8688
rect 48 8584 80 8616
rect 120 8584 152 8616
rect 192 8584 224 8616
rect 264 8584 296 8616
rect 336 8584 368 8616
rect 408 8584 440 8616
rect 480 8584 512 8616
rect 552 8584 584 8616
rect 624 8584 656 8616
rect 696 8584 728 8616
rect 768 8584 800 8616
rect 840 8584 872 8616
rect 912 8584 944 8616
rect 984 8584 1016 8616
rect 1056 8584 1088 8616
rect 1128 8584 1160 8616
rect 1200 8584 1232 8616
rect 1272 8584 1304 8616
rect 1344 8584 1376 8616
rect 1416 8584 1448 8616
rect 1488 8584 1520 8616
rect 1560 8584 1592 8616
rect 1632 8584 1664 8616
rect 1704 8584 1736 8616
rect 1776 8584 1808 8616
rect 1848 8584 1880 8616
rect 1920 8584 1952 8616
rect 48 8512 80 8544
rect 120 8512 152 8544
rect 192 8512 224 8544
rect 264 8512 296 8544
rect 336 8512 368 8544
rect 408 8512 440 8544
rect 480 8512 512 8544
rect 552 8512 584 8544
rect 624 8512 656 8544
rect 696 8512 728 8544
rect 768 8512 800 8544
rect 840 8512 872 8544
rect 912 8512 944 8544
rect 984 8512 1016 8544
rect 1056 8512 1088 8544
rect 1128 8512 1160 8544
rect 1200 8512 1232 8544
rect 1272 8512 1304 8544
rect 1344 8512 1376 8544
rect 1416 8512 1448 8544
rect 1488 8512 1520 8544
rect 1560 8512 1592 8544
rect 1632 8512 1664 8544
rect 1704 8512 1736 8544
rect 1776 8512 1808 8544
rect 1848 8512 1880 8544
rect 1920 8512 1952 8544
rect 48 8440 80 8472
rect 120 8440 152 8472
rect 192 8440 224 8472
rect 264 8440 296 8472
rect 336 8440 368 8472
rect 408 8440 440 8472
rect 480 8440 512 8472
rect 552 8440 584 8472
rect 624 8440 656 8472
rect 696 8440 728 8472
rect 768 8440 800 8472
rect 840 8440 872 8472
rect 912 8440 944 8472
rect 984 8440 1016 8472
rect 1056 8440 1088 8472
rect 1128 8440 1160 8472
rect 1200 8440 1232 8472
rect 1272 8440 1304 8472
rect 1344 8440 1376 8472
rect 1416 8440 1448 8472
rect 1488 8440 1520 8472
rect 1560 8440 1592 8472
rect 1632 8440 1664 8472
rect 1704 8440 1736 8472
rect 1776 8440 1808 8472
rect 1848 8440 1880 8472
rect 1920 8440 1952 8472
rect 48 8368 80 8400
rect 120 8368 152 8400
rect 192 8368 224 8400
rect 264 8368 296 8400
rect 336 8368 368 8400
rect 408 8368 440 8400
rect 480 8368 512 8400
rect 552 8368 584 8400
rect 624 8368 656 8400
rect 696 8368 728 8400
rect 768 8368 800 8400
rect 840 8368 872 8400
rect 912 8368 944 8400
rect 984 8368 1016 8400
rect 1056 8368 1088 8400
rect 1128 8368 1160 8400
rect 1200 8368 1232 8400
rect 1272 8368 1304 8400
rect 1344 8368 1376 8400
rect 1416 8368 1448 8400
rect 1488 8368 1520 8400
rect 1560 8368 1592 8400
rect 1632 8368 1664 8400
rect 1704 8368 1736 8400
rect 1776 8368 1808 8400
rect 1848 8368 1880 8400
rect 1920 8368 1952 8400
rect 48 8296 80 8328
rect 120 8296 152 8328
rect 192 8296 224 8328
rect 264 8296 296 8328
rect 336 8296 368 8328
rect 408 8296 440 8328
rect 480 8296 512 8328
rect 552 8296 584 8328
rect 624 8296 656 8328
rect 696 8296 728 8328
rect 768 8296 800 8328
rect 840 8296 872 8328
rect 912 8296 944 8328
rect 984 8296 1016 8328
rect 1056 8296 1088 8328
rect 1128 8296 1160 8328
rect 1200 8296 1232 8328
rect 1272 8296 1304 8328
rect 1344 8296 1376 8328
rect 1416 8296 1448 8328
rect 1488 8296 1520 8328
rect 1560 8296 1592 8328
rect 1632 8296 1664 8328
rect 1704 8296 1736 8328
rect 1776 8296 1808 8328
rect 1848 8296 1880 8328
rect 1920 8296 1952 8328
rect 48 8224 80 8256
rect 120 8224 152 8256
rect 192 8224 224 8256
rect 264 8224 296 8256
rect 336 8224 368 8256
rect 408 8224 440 8256
rect 480 8224 512 8256
rect 552 8224 584 8256
rect 624 8224 656 8256
rect 696 8224 728 8256
rect 768 8224 800 8256
rect 840 8224 872 8256
rect 912 8224 944 8256
rect 984 8224 1016 8256
rect 1056 8224 1088 8256
rect 1128 8224 1160 8256
rect 1200 8224 1232 8256
rect 1272 8224 1304 8256
rect 1344 8224 1376 8256
rect 1416 8224 1448 8256
rect 1488 8224 1520 8256
rect 1560 8224 1592 8256
rect 1632 8224 1664 8256
rect 1704 8224 1736 8256
rect 1776 8224 1808 8256
rect 1848 8224 1880 8256
rect 1920 8224 1952 8256
rect 48 8152 80 8184
rect 120 8152 152 8184
rect 192 8152 224 8184
rect 264 8152 296 8184
rect 336 8152 368 8184
rect 408 8152 440 8184
rect 480 8152 512 8184
rect 552 8152 584 8184
rect 624 8152 656 8184
rect 696 8152 728 8184
rect 768 8152 800 8184
rect 840 8152 872 8184
rect 912 8152 944 8184
rect 984 8152 1016 8184
rect 1056 8152 1088 8184
rect 1128 8152 1160 8184
rect 1200 8152 1232 8184
rect 1272 8152 1304 8184
rect 1344 8152 1376 8184
rect 1416 8152 1448 8184
rect 1488 8152 1520 8184
rect 1560 8152 1592 8184
rect 1632 8152 1664 8184
rect 1704 8152 1736 8184
rect 1776 8152 1808 8184
rect 1848 8152 1880 8184
rect 1920 8152 1952 8184
rect 48 8080 80 8112
rect 120 8080 152 8112
rect 192 8080 224 8112
rect 264 8080 296 8112
rect 336 8080 368 8112
rect 408 8080 440 8112
rect 480 8080 512 8112
rect 552 8080 584 8112
rect 624 8080 656 8112
rect 696 8080 728 8112
rect 768 8080 800 8112
rect 840 8080 872 8112
rect 912 8080 944 8112
rect 984 8080 1016 8112
rect 1056 8080 1088 8112
rect 1128 8080 1160 8112
rect 1200 8080 1232 8112
rect 1272 8080 1304 8112
rect 1344 8080 1376 8112
rect 1416 8080 1448 8112
rect 1488 8080 1520 8112
rect 1560 8080 1592 8112
rect 1632 8080 1664 8112
rect 1704 8080 1736 8112
rect 1776 8080 1808 8112
rect 1848 8080 1880 8112
rect 1920 8080 1952 8112
rect 48 8008 80 8040
rect 120 8008 152 8040
rect 192 8008 224 8040
rect 264 8008 296 8040
rect 336 8008 368 8040
rect 408 8008 440 8040
rect 480 8008 512 8040
rect 552 8008 584 8040
rect 624 8008 656 8040
rect 696 8008 728 8040
rect 768 8008 800 8040
rect 840 8008 872 8040
rect 912 8008 944 8040
rect 984 8008 1016 8040
rect 1056 8008 1088 8040
rect 1128 8008 1160 8040
rect 1200 8008 1232 8040
rect 1272 8008 1304 8040
rect 1344 8008 1376 8040
rect 1416 8008 1448 8040
rect 1488 8008 1520 8040
rect 1560 8008 1592 8040
rect 1632 8008 1664 8040
rect 1704 8008 1736 8040
rect 1776 8008 1808 8040
rect 1848 8008 1880 8040
rect 1920 8008 1952 8040
rect 48 7936 80 7968
rect 120 7936 152 7968
rect 192 7936 224 7968
rect 264 7936 296 7968
rect 336 7936 368 7968
rect 408 7936 440 7968
rect 480 7936 512 7968
rect 552 7936 584 7968
rect 624 7936 656 7968
rect 696 7936 728 7968
rect 768 7936 800 7968
rect 840 7936 872 7968
rect 912 7936 944 7968
rect 984 7936 1016 7968
rect 1056 7936 1088 7968
rect 1128 7936 1160 7968
rect 1200 7936 1232 7968
rect 1272 7936 1304 7968
rect 1344 7936 1376 7968
rect 1416 7936 1448 7968
rect 1488 7936 1520 7968
rect 1560 7936 1592 7968
rect 1632 7936 1664 7968
rect 1704 7936 1736 7968
rect 1776 7936 1808 7968
rect 1848 7936 1880 7968
rect 1920 7936 1952 7968
rect 48 7864 80 7896
rect 120 7864 152 7896
rect 192 7864 224 7896
rect 264 7864 296 7896
rect 336 7864 368 7896
rect 408 7864 440 7896
rect 480 7864 512 7896
rect 552 7864 584 7896
rect 624 7864 656 7896
rect 696 7864 728 7896
rect 768 7864 800 7896
rect 840 7864 872 7896
rect 912 7864 944 7896
rect 984 7864 1016 7896
rect 1056 7864 1088 7896
rect 1128 7864 1160 7896
rect 1200 7864 1232 7896
rect 1272 7864 1304 7896
rect 1344 7864 1376 7896
rect 1416 7864 1448 7896
rect 1488 7864 1520 7896
rect 1560 7864 1592 7896
rect 1632 7864 1664 7896
rect 1704 7864 1736 7896
rect 1776 7864 1808 7896
rect 1848 7864 1880 7896
rect 1920 7864 1952 7896
rect 48 7792 80 7824
rect 120 7792 152 7824
rect 192 7792 224 7824
rect 264 7792 296 7824
rect 336 7792 368 7824
rect 408 7792 440 7824
rect 480 7792 512 7824
rect 552 7792 584 7824
rect 624 7792 656 7824
rect 696 7792 728 7824
rect 768 7792 800 7824
rect 840 7792 872 7824
rect 912 7792 944 7824
rect 984 7792 1016 7824
rect 1056 7792 1088 7824
rect 1128 7792 1160 7824
rect 1200 7792 1232 7824
rect 1272 7792 1304 7824
rect 1344 7792 1376 7824
rect 1416 7792 1448 7824
rect 1488 7792 1520 7824
rect 1560 7792 1592 7824
rect 1632 7792 1664 7824
rect 1704 7792 1736 7824
rect 1776 7792 1808 7824
rect 1848 7792 1880 7824
rect 1920 7792 1952 7824
rect 48 7720 80 7752
rect 120 7720 152 7752
rect 192 7720 224 7752
rect 264 7720 296 7752
rect 336 7720 368 7752
rect 408 7720 440 7752
rect 480 7720 512 7752
rect 552 7720 584 7752
rect 624 7720 656 7752
rect 696 7720 728 7752
rect 768 7720 800 7752
rect 840 7720 872 7752
rect 912 7720 944 7752
rect 984 7720 1016 7752
rect 1056 7720 1088 7752
rect 1128 7720 1160 7752
rect 1200 7720 1232 7752
rect 1272 7720 1304 7752
rect 1344 7720 1376 7752
rect 1416 7720 1448 7752
rect 1488 7720 1520 7752
rect 1560 7720 1592 7752
rect 1632 7720 1664 7752
rect 1704 7720 1736 7752
rect 1776 7720 1808 7752
rect 1848 7720 1880 7752
rect 1920 7720 1952 7752
rect 48 7648 80 7680
rect 120 7648 152 7680
rect 192 7648 224 7680
rect 264 7648 296 7680
rect 336 7648 368 7680
rect 408 7648 440 7680
rect 480 7648 512 7680
rect 552 7648 584 7680
rect 624 7648 656 7680
rect 696 7648 728 7680
rect 768 7648 800 7680
rect 840 7648 872 7680
rect 912 7648 944 7680
rect 984 7648 1016 7680
rect 1056 7648 1088 7680
rect 1128 7648 1160 7680
rect 1200 7648 1232 7680
rect 1272 7648 1304 7680
rect 1344 7648 1376 7680
rect 1416 7648 1448 7680
rect 1488 7648 1520 7680
rect 1560 7648 1592 7680
rect 1632 7648 1664 7680
rect 1704 7648 1736 7680
rect 1776 7648 1808 7680
rect 1848 7648 1880 7680
rect 1920 7648 1952 7680
rect 48 7576 80 7608
rect 120 7576 152 7608
rect 192 7576 224 7608
rect 264 7576 296 7608
rect 336 7576 368 7608
rect 408 7576 440 7608
rect 480 7576 512 7608
rect 552 7576 584 7608
rect 624 7576 656 7608
rect 696 7576 728 7608
rect 768 7576 800 7608
rect 840 7576 872 7608
rect 912 7576 944 7608
rect 984 7576 1016 7608
rect 1056 7576 1088 7608
rect 1128 7576 1160 7608
rect 1200 7576 1232 7608
rect 1272 7576 1304 7608
rect 1344 7576 1376 7608
rect 1416 7576 1448 7608
rect 1488 7576 1520 7608
rect 1560 7576 1592 7608
rect 1632 7576 1664 7608
rect 1704 7576 1736 7608
rect 1776 7576 1808 7608
rect 1848 7576 1880 7608
rect 1920 7576 1952 7608
rect 48 7504 80 7536
rect 120 7504 152 7536
rect 192 7504 224 7536
rect 264 7504 296 7536
rect 336 7504 368 7536
rect 408 7504 440 7536
rect 480 7504 512 7536
rect 552 7504 584 7536
rect 624 7504 656 7536
rect 696 7504 728 7536
rect 768 7504 800 7536
rect 840 7504 872 7536
rect 912 7504 944 7536
rect 984 7504 1016 7536
rect 1056 7504 1088 7536
rect 1128 7504 1160 7536
rect 1200 7504 1232 7536
rect 1272 7504 1304 7536
rect 1344 7504 1376 7536
rect 1416 7504 1448 7536
rect 1488 7504 1520 7536
rect 1560 7504 1592 7536
rect 1632 7504 1664 7536
rect 1704 7504 1736 7536
rect 1776 7504 1808 7536
rect 1848 7504 1880 7536
rect 1920 7504 1952 7536
rect 48 7432 80 7464
rect 120 7432 152 7464
rect 192 7432 224 7464
rect 264 7432 296 7464
rect 336 7432 368 7464
rect 408 7432 440 7464
rect 480 7432 512 7464
rect 552 7432 584 7464
rect 624 7432 656 7464
rect 696 7432 728 7464
rect 768 7432 800 7464
rect 840 7432 872 7464
rect 912 7432 944 7464
rect 984 7432 1016 7464
rect 1056 7432 1088 7464
rect 1128 7432 1160 7464
rect 1200 7432 1232 7464
rect 1272 7432 1304 7464
rect 1344 7432 1376 7464
rect 1416 7432 1448 7464
rect 1488 7432 1520 7464
rect 1560 7432 1592 7464
rect 1632 7432 1664 7464
rect 1704 7432 1736 7464
rect 1776 7432 1808 7464
rect 1848 7432 1880 7464
rect 1920 7432 1952 7464
rect 48 7360 80 7392
rect 120 7360 152 7392
rect 192 7360 224 7392
rect 264 7360 296 7392
rect 336 7360 368 7392
rect 408 7360 440 7392
rect 480 7360 512 7392
rect 552 7360 584 7392
rect 624 7360 656 7392
rect 696 7360 728 7392
rect 768 7360 800 7392
rect 840 7360 872 7392
rect 912 7360 944 7392
rect 984 7360 1016 7392
rect 1056 7360 1088 7392
rect 1128 7360 1160 7392
rect 1200 7360 1232 7392
rect 1272 7360 1304 7392
rect 1344 7360 1376 7392
rect 1416 7360 1448 7392
rect 1488 7360 1520 7392
rect 1560 7360 1592 7392
rect 1632 7360 1664 7392
rect 1704 7360 1736 7392
rect 1776 7360 1808 7392
rect 1848 7360 1880 7392
rect 1920 7360 1952 7392
rect 48 7288 80 7320
rect 120 7288 152 7320
rect 192 7288 224 7320
rect 264 7288 296 7320
rect 336 7288 368 7320
rect 408 7288 440 7320
rect 480 7288 512 7320
rect 552 7288 584 7320
rect 624 7288 656 7320
rect 696 7288 728 7320
rect 768 7288 800 7320
rect 840 7288 872 7320
rect 912 7288 944 7320
rect 984 7288 1016 7320
rect 1056 7288 1088 7320
rect 1128 7288 1160 7320
rect 1200 7288 1232 7320
rect 1272 7288 1304 7320
rect 1344 7288 1376 7320
rect 1416 7288 1448 7320
rect 1488 7288 1520 7320
rect 1560 7288 1592 7320
rect 1632 7288 1664 7320
rect 1704 7288 1736 7320
rect 1776 7288 1808 7320
rect 1848 7288 1880 7320
rect 1920 7288 1952 7320
rect 48 7216 80 7248
rect 120 7216 152 7248
rect 192 7216 224 7248
rect 264 7216 296 7248
rect 336 7216 368 7248
rect 408 7216 440 7248
rect 480 7216 512 7248
rect 552 7216 584 7248
rect 624 7216 656 7248
rect 696 7216 728 7248
rect 768 7216 800 7248
rect 840 7216 872 7248
rect 912 7216 944 7248
rect 984 7216 1016 7248
rect 1056 7216 1088 7248
rect 1128 7216 1160 7248
rect 1200 7216 1232 7248
rect 1272 7216 1304 7248
rect 1344 7216 1376 7248
rect 1416 7216 1448 7248
rect 1488 7216 1520 7248
rect 1560 7216 1592 7248
rect 1632 7216 1664 7248
rect 1704 7216 1736 7248
rect 1776 7216 1808 7248
rect 1848 7216 1880 7248
rect 1920 7216 1952 7248
rect 48 7144 80 7176
rect 120 7144 152 7176
rect 192 7144 224 7176
rect 264 7144 296 7176
rect 336 7144 368 7176
rect 408 7144 440 7176
rect 480 7144 512 7176
rect 552 7144 584 7176
rect 624 7144 656 7176
rect 696 7144 728 7176
rect 768 7144 800 7176
rect 840 7144 872 7176
rect 912 7144 944 7176
rect 984 7144 1016 7176
rect 1056 7144 1088 7176
rect 1128 7144 1160 7176
rect 1200 7144 1232 7176
rect 1272 7144 1304 7176
rect 1344 7144 1376 7176
rect 1416 7144 1448 7176
rect 1488 7144 1520 7176
rect 1560 7144 1592 7176
rect 1632 7144 1664 7176
rect 1704 7144 1736 7176
rect 1776 7144 1808 7176
rect 1848 7144 1880 7176
rect 1920 7144 1952 7176
rect 48 7072 80 7104
rect 120 7072 152 7104
rect 192 7072 224 7104
rect 264 7072 296 7104
rect 336 7072 368 7104
rect 408 7072 440 7104
rect 480 7072 512 7104
rect 552 7072 584 7104
rect 624 7072 656 7104
rect 696 7072 728 7104
rect 768 7072 800 7104
rect 840 7072 872 7104
rect 912 7072 944 7104
rect 984 7072 1016 7104
rect 1056 7072 1088 7104
rect 1128 7072 1160 7104
rect 1200 7072 1232 7104
rect 1272 7072 1304 7104
rect 1344 7072 1376 7104
rect 1416 7072 1448 7104
rect 1488 7072 1520 7104
rect 1560 7072 1592 7104
rect 1632 7072 1664 7104
rect 1704 7072 1736 7104
rect 1776 7072 1808 7104
rect 1848 7072 1880 7104
rect 1920 7072 1952 7104
rect 48 7000 80 7032
rect 120 7000 152 7032
rect 192 7000 224 7032
rect 264 7000 296 7032
rect 336 7000 368 7032
rect 408 7000 440 7032
rect 480 7000 512 7032
rect 552 7000 584 7032
rect 624 7000 656 7032
rect 696 7000 728 7032
rect 768 7000 800 7032
rect 840 7000 872 7032
rect 912 7000 944 7032
rect 984 7000 1016 7032
rect 1056 7000 1088 7032
rect 1128 7000 1160 7032
rect 1200 7000 1232 7032
rect 1272 7000 1304 7032
rect 1344 7000 1376 7032
rect 1416 7000 1448 7032
rect 1488 7000 1520 7032
rect 1560 7000 1592 7032
rect 1632 7000 1664 7032
rect 1704 7000 1736 7032
rect 1776 7000 1808 7032
rect 1848 7000 1880 7032
rect 1920 7000 1952 7032
rect 48 6928 80 6960
rect 120 6928 152 6960
rect 192 6928 224 6960
rect 264 6928 296 6960
rect 336 6928 368 6960
rect 408 6928 440 6960
rect 480 6928 512 6960
rect 552 6928 584 6960
rect 624 6928 656 6960
rect 696 6928 728 6960
rect 768 6928 800 6960
rect 840 6928 872 6960
rect 912 6928 944 6960
rect 984 6928 1016 6960
rect 1056 6928 1088 6960
rect 1128 6928 1160 6960
rect 1200 6928 1232 6960
rect 1272 6928 1304 6960
rect 1344 6928 1376 6960
rect 1416 6928 1448 6960
rect 1488 6928 1520 6960
rect 1560 6928 1592 6960
rect 1632 6928 1664 6960
rect 1704 6928 1736 6960
rect 1776 6928 1808 6960
rect 1848 6928 1880 6960
rect 1920 6928 1952 6960
rect 48 6856 80 6888
rect 120 6856 152 6888
rect 192 6856 224 6888
rect 264 6856 296 6888
rect 336 6856 368 6888
rect 408 6856 440 6888
rect 480 6856 512 6888
rect 552 6856 584 6888
rect 624 6856 656 6888
rect 696 6856 728 6888
rect 768 6856 800 6888
rect 840 6856 872 6888
rect 912 6856 944 6888
rect 984 6856 1016 6888
rect 1056 6856 1088 6888
rect 1128 6856 1160 6888
rect 1200 6856 1232 6888
rect 1272 6856 1304 6888
rect 1344 6856 1376 6888
rect 1416 6856 1448 6888
rect 1488 6856 1520 6888
rect 1560 6856 1592 6888
rect 1632 6856 1664 6888
rect 1704 6856 1736 6888
rect 1776 6856 1808 6888
rect 1848 6856 1880 6888
rect 1920 6856 1952 6888
rect 120 6512 152 6544
rect 192 6512 224 6544
rect 264 6512 296 6544
rect 336 6512 368 6544
rect 408 6512 440 6544
rect 480 6512 512 6544
rect 552 6512 584 6544
rect 624 6512 656 6544
rect 696 6512 728 6544
rect 768 6512 800 6544
rect 840 6512 872 6544
rect 912 6512 944 6544
rect 984 6512 1016 6544
rect 1056 6512 1088 6544
rect 1128 6512 1160 6544
rect 1200 6512 1232 6544
rect 1272 6512 1304 6544
rect 1344 6512 1376 6544
rect 1416 6512 1448 6544
rect 1488 6512 1520 6544
rect 1560 6512 1592 6544
rect 1632 6512 1664 6544
rect 1704 6512 1736 6544
rect 1776 6512 1808 6544
rect 1848 6512 1880 6544
rect 1920 6512 1952 6544
rect 48 6440 80 6472
rect 120 6440 152 6472
rect 192 6440 224 6472
rect 264 6440 296 6472
rect 336 6440 368 6472
rect 408 6440 440 6472
rect 480 6440 512 6472
rect 552 6440 584 6472
rect 624 6440 656 6472
rect 696 6440 728 6472
rect 768 6440 800 6472
rect 840 6440 872 6472
rect 912 6440 944 6472
rect 984 6440 1016 6472
rect 1056 6440 1088 6472
rect 1128 6440 1160 6472
rect 1200 6440 1232 6472
rect 1272 6440 1304 6472
rect 1344 6440 1376 6472
rect 1416 6440 1448 6472
rect 1488 6440 1520 6472
rect 1560 6440 1592 6472
rect 1632 6440 1664 6472
rect 1704 6440 1736 6472
rect 1776 6440 1808 6472
rect 1848 6440 1880 6472
rect 1920 6440 1952 6472
rect 48 6368 80 6400
rect 120 6368 152 6400
rect 192 6368 224 6400
rect 264 6368 296 6400
rect 336 6368 368 6400
rect 408 6368 440 6400
rect 480 6368 512 6400
rect 552 6368 584 6400
rect 624 6368 656 6400
rect 696 6368 728 6400
rect 768 6368 800 6400
rect 840 6368 872 6400
rect 912 6368 944 6400
rect 984 6368 1016 6400
rect 1056 6368 1088 6400
rect 1128 6368 1160 6400
rect 1200 6368 1232 6400
rect 1272 6368 1304 6400
rect 1344 6368 1376 6400
rect 1416 6368 1448 6400
rect 1488 6368 1520 6400
rect 1560 6368 1592 6400
rect 1632 6368 1664 6400
rect 1704 6368 1736 6400
rect 1776 6368 1808 6400
rect 1848 6368 1880 6400
rect 1920 6368 1952 6400
rect 48 6296 80 6328
rect 120 6296 152 6328
rect 192 6296 224 6328
rect 264 6296 296 6328
rect 336 6296 368 6328
rect 408 6296 440 6328
rect 480 6296 512 6328
rect 552 6296 584 6328
rect 624 6296 656 6328
rect 696 6296 728 6328
rect 768 6296 800 6328
rect 840 6296 872 6328
rect 912 6296 944 6328
rect 984 6296 1016 6328
rect 1056 6296 1088 6328
rect 1128 6296 1160 6328
rect 1200 6296 1232 6328
rect 1272 6296 1304 6328
rect 1344 6296 1376 6328
rect 1416 6296 1448 6328
rect 1488 6296 1520 6328
rect 1560 6296 1592 6328
rect 1632 6296 1664 6328
rect 1704 6296 1736 6328
rect 1776 6296 1808 6328
rect 1848 6296 1880 6328
rect 1920 6296 1952 6328
rect 48 6224 80 6256
rect 120 6224 152 6256
rect 192 6224 224 6256
rect 264 6224 296 6256
rect 336 6224 368 6256
rect 408 6224 440 6256
rect 480 6224 512 6256
rect 552 6224 584 6256
rect 624 6224 656 6256
rect 696 6224 728 6256
rect 768 6224 800 6256
rect 840 6224 872 6256
rect 912 6224 944 6256
rect 984 6224 1016 6256
rect 1056 6224 1088 6256
rect 1128 6224 1160 6256
rect 1200 6224 1232 6256
rect 1272 6224 1304 6256
rect 1344 6224 1376 6256
rect 1416 6224 1448 6256
rect 1488 6224 1520 6256
rect 1560 6224 1592 6256
rect 1632 6224 1664 6256
rect 1704 6224 1736 6256
rect 1776 6224 1808 6256
rect 1848 6224 1880 6256
rect 1920 6224 1952 6256
rect 48 6152 80 6184
rect 120 6152 152 6184
rect 192 6152 224 6184
rect 264 6152 296 6184
rect 336 6152 368 6184
rect 408 6152 440 6184
rect 480 6152 512 6184
rect 552 6152 584 6184
rect 624 6152 656 6184
rect 696 6152 728 6184
rect 768 6152 800 6184
rect 840 6152 872 6184
rect 912 6152 944 6184
rect 984 6152 1016 6184
rect 1056 6152 1088 6184
rect 1128 6152 1160 6184
rect 1200 6152 1232 6184
rect 1272 6152 1304 6184
rect 1344 6152 1376 6184
rect 1416 6152 1448 6184
rect 1488 6152 1520 6184
rect 1560 6152 1592 6184
rect 1632 6152 1664 6184
rect 1704 6152 1736 6184
rect 1776 6152 1808 6184
rect 1848 6152 1880 6184
rect 1920 6152 1952 6184
rect 48 6080 80 6112
rect 120 6080 152 6112
rect 192 6080 224 6112
rect 264 6080 296 6112
rect 336 6080 368 6112
rect 408 6080 440 6112
rect 480 6080 512 6112
rect 552 6080 584 6112
rect 624 6080 656 6112
rect 696 6080 728 6112
rect 768 6080 800 6112
rect 840 6080 872 6112
rect 912 6080 944 6112
rect 984 6080 1016 6112
rect 1056 6080 1088 6112
rect 1128 6080 1160 6112
rect 1200 6080 1232 6112
rect 1272 6080 1304 6112
rect 1344 6080 1376 6112
rect 1416 6080 1448 6112
rect 1488 6080 1520 6112
rect 1560 6080 1592 6112
rect 1632 6080 1664 6112
rect 1704 6080 1736 6112
rect 1776 6080 1808 6112
rect 1848 6080 1880 6112
rect 1920 6080 1952 6112
rect 48 6008 80 6040
rect 120 6008 152 6040
rect 192 6008 224 6040
rect 264 6008 296 6040
rect 336 6008 368 6040
rect 408 6008 440 6040
rect 480 6008 512 6040
rect 552 6008 584 6040
rect 624 6008 656 6040
rect 696 6008 728 6040
rect 768 6008 800 6040
rect 840 6008 872 6040
rect 912 6008 944 6040
rect 984 6008 1016 6040
rect 1056 6008 1088 6040
rect 1128 6008 1160 6040
rect 1200 6008 1232 6040
rect 1272 6008 1304 6040
rect 1344 6008 1376 6040
rect 1416 6008 1448 6040
rect 1488 6008 1520 6040
rect 1560 6008 1592 6040
rect 1632 6008 1664 6040
rect 1704 6008 1736 6040
rect 1776 6008 1808 6040
rect 1848 6008 1880 6040
rect 1920 6008 1952 6040
rect 48 5936 80 5968
rect 120 5936 152 5968
rect 192 5936 224 5968
rect 264 5936 296 5968
rect 336 5936 368 5968
rect 408 5936 440 5968
rect 480 5936 512 5968
rect 552 5936 584 5968
rect 624 5936 656 5968
rect 696 5936 728 5968
rect 768 5936 800 5968
rect 840 5936 872 5968
rect 912 5936 944 5968
rect 984 5936 1016 5968
rect 1056 5936 1088 5968
rect 1128 5936 1160 5968
rect 1200 5936 1232 5968
rect 1272 5936 1304 5968
rect 1344 5936 1376 5968
rect 1416 5936 1448 5968
rect 1488 5936 1520 5968
rect 1560 5936 1592 5968
rect 1632 5936 1664 5968
rect 1704 5936 1736 5968
rect 1776 5936 1808 5968
rect 1848 5936 1880 5968
rect 1920 5936 1952 5968
rect 48 5864 80 5896
rect 120 5864 152 5896
rect 192 5864 224 5896
rect 264 5864 296 5896
rect 336 5864 368 5896
rect 408 5864 440 5896
rect 480 5864 512 5896
rect 552 5864 584 5896
rect 624 5864 656 5896
rect 696 5864 728 5896
rect 768 5864 800 5896
rect 840 5864 872 5896
rect 912 5864 944 5896
rect 984 5864 1016 5896
rect 1056 5864 1088 5896
rect 1128 5864 1160 5896
rect 1200 5864 1232 5896
rect 1272 5864 1304 5896
rect 1344 5864 1376 5896
rect 1416 5864 1448 5896
rect 1488 5864 1520 5896
rect 1560 5864 1592 5896
rect 1632 5864 1664 5896
rect 1704 5864 1736 5896
rect 1776 5864 1808 5896
rect 1848 5864 1880 5896
rect 1920 5864 1952 5896
rect 48 5792 80 5824
rect 120 5792 152 5824
rect 192 5792 224 5824
rect 264 5792 296 5824
rect 336 5792 368 5824
rect 408 5792 440 5824
rect 480 5792 512 5824
rect 552 5792 584 5824
rect 624 5792 656 5824
rect 696 5792 728 5824
rect 768 5792 800 5824
rect 840 5792 872 5824
rect 912 5792 944 5824
rect 984 5792 1016 5824
rect 1056 5792 1088 5824
rect 1128 5792 1160 5824
rect 1200 5792 1232 5824
rect 1272 5792 1304 5824
rect 1344 5792 1376 5824
rect 1416 5792 1448 5824
rect 1488 5792 1520 5824
rect 1560 5792 1592 5824
rect 1632 5792 1664 5824
rect 1704 5792 1736 5824
rect 1776 5792 1808 5824
rect 1848 5792 1880 5824
rect 1920 5792 1952 5824
rect 48 5720 80 5752
rect 120 5720 152 5752
rect 192 5720 224 5752
rect 264 5720 296 5752
rect 336 5720 368 5752
rect 408 5720 440 5752
rect 480 5720 512 5752
rect 552 5720 584 5752
rect 624 5720 656 5752
rect 696 5720 728 5752
rect 768 5720 800 5752
rect 840 5720 872 5752
rect 912 5720 944 5752
rect 984 5720 1016 5752
rect 1056 5720 1088 5752
rect 1128 5720 1160 5752
rect 1200 5720 1232 5752
rect 1272 5720 1304 5752
rect 1344 5720 1376 5752
rect 1416 5720 1448 5752
rect 1488 5720 1520 5752
rect 1560 5720 1592 5752
rect 1632 5720 1664 5752
rect 1704 5720 1736 5752
rect 1776 5720 1808 5752
rect 1848 5720 1880 5752
rect 1920 5720 1952 5752
rect 48 5648 80 5680
rect 120 5648 152 5680
rect 192 5648 224 5680
rect 264 5648 296 5680
rect 336 5648 368 5680
rect 408 5648 440 5680
rect 480 5648 512 5680
rect 552 5648 584 5680
rect 624 5648 656 5680
rect 696 5648 728 5680
rect 768 5648 800 5680
rect 840 5648 872 5680
rect 912 5648 944 5680
rect 984 5648 1016 5680
rect 1056 5648 1088 5680
rect 1128 5648 1160 5680
rect 1200 5648 1232 5680
rect 1272 5648 1304 5680
rect 1344 5648 1376 5680
rect 1416 5648 1448 5680
rect 1488 5648 1520 5680
rect 1560 5648 1592 5680
rect 1632 5648 1664 5680
rect 1704 5648 1736 5680
rect 1776 5648 1808 5680
rect 1848 5648 1880 5680
rect 1920 5648 1952 5680
rect 48 5576 80 5608
rect 120 5576 152 5608
rect 192 5576 224 5608
rect 264 5576 296 5608
rect 336 5576 368 5608
rect 408 5576 440 5608
rect 480 5576 512 5608
rect 552 5576 584 5608
rect 624 5576 656 5608
rect 696 5576 728 5608
rect 768 5576 800 5608
rect 840 5576 872 5608
rect 912 5576 944 5608
rect 984 5576 1016 5608
rect 1056 5576 1088 5608
rect 1128 5576 1160 5608
rect 1200 5576 1232 5608
rect 1272 5576 1304 5608
rect 1344 5576 1376 5608
rect 1416 5576 1448 5608
rect 1488 5576 1520 5608
rect 1560 5576 1592 5608
rect 1632 5576 1664 5608
rect 1704 5576 1736 5608
rect 1776 5576 1808 5608
rect 1848 5576 1880 5608
rect 1920 5576 1952 5608
rect 48 5504 80 5536
rect 120 5504 152 5536
rect 192 5504 224 5536
rect 264 5504 296 5536
rect 336 5504 368 5536
rect 408 5504 440 5536
rect 480 5504 512 5536
rect 552 5504 584 5536
rect 624 5504 656 5536
rect 696 5504 728 5536
rect 768 5504 800 5536
rect 840 5504 872 5536
rect 912 5504 944 5536
rect 984 5504 1016 5536
rect 1056 5504 1088 5536
rect 1128 5504 1160 5536
rect 1200 5504 1232 5536
rect 1272 5504 1304 5536
rect 1344 5504 1376 5536
rect 1416 5504 1448 5536
rect 1488 5504 1520 5536
rect 1560 5504 1592 5536
rect 1632 5504 1664 5536
rect 1704 5504 1736 5536
rect 1776 5504 1808 5536
rect 1848 5504 1880 5536
rect 1920 5504 1952 5536
rect 48 5432 80 5464
rect 120 5432 152 5464
rect 192 5432 224 5464
rect 264 5432 296 5464
rect 336 5432 368 5464
rect 408 5432 440 5464
rect 480 5432 512 5464
rect 552 5432 584 5464
rect 624 5432 656 5464
rect 696 5432 728 5464
rect 768 5432 800 5464
rect 840 5432 872 5464
rect 912 5432 944 5464
rect 984 5432 1016 5464
rect 1056 5432 1088 5464
rect 1128 5432 1160 5464
rect 1200 5432 1232 5464
rect 1272 5432 1304 5464
rect 1344 5432 1376 5464
rect 1416 5432 1448 5464
rect 1488 5432 1520 5464
rect 1560 5432 1592 5464
rect 1632 5432 1664 5464
rect 1704 5432 1736 5464
rect 1776 5432 1808 5464
rect 1848 5432 1880 5464
rect 1920 5432 1952 5464
rect 48 5360 80 5392
rect 120 5360 152 5392
rect 192 5360 224 5392
rect 264 5360 296 5392
rect 336 5360 368 5392
rect 408 5360 440 5392
rect 480 5360 512 5392
rect 552 5360 584 5392
rect 624 5360 656 5392
rect 696 5360 728 5392
rect 768 5360 800 5392
rect 840 5360 872 5392
rect 912 5360 944 5392
rect 984 5360 1016 5392
rect 1056 5360 1088 5392
rect 1128 5360 1160 5392
rect 1200 5360 1232 5392
rect 1272 5360 1304 5392
rect 1344 5360 1376 5392
rect 1416 5360 1448 5392
rect 1488 5360 1520 5392
rect 1560 5360 1592 5392
rect 1632 5360 1664 5392
rect 1704 5360 1736 5392
rect 1776 5360 1808 5392
rect 1848 5360 1880 5392
rect 1920 5360 1952 5392
rect 48 5288 80 5320
rect 120 5288 152 5320
rect 192 5288 224 5320
rect 264 5288 296 5320
rect 336 5288 368 5320
rect 408 5288 440 5320
rect 480 5288 512 5320
rect 552 5288 584 5320
rect 624 5288 656 5320
rect 696 5288 728 5320
rect 768 5288 800 5320
rect 840 5288 872 5320
rect 912 5288 944 5320
rect 984 5288 1016 5320
rect 1056 5288 1088 5320
rect 1128 5288 1160 5320
rect 1200 5288 1232 5320
rect 1272 5288 1304 5320
rect 1344 5288 1376 5320
rect 1416 5288 1448 5320
rect 1488 5288 1520 5320
rect 1560 5288 1592 5320
rect 1632 5288 1664 5320
rect 1704 5288 1736 5320
rect 1776 5288 1808 5320
rect 1848 5288 1880 5320
rect 1920 5288 1952 5320
rect 48 5216 80 5248
rect 120 5216 152 5248
rect 192 5216 224 5248
rect 264 5216 296 5248
rect 336 5216 368 5248
rect 408 5216 440 5248
rect 480 5216 512 5248
rect 552 5216 584 5248
rect 624 5216 656 5248
rect 696 5216 728 5248
rect 768 5216 800 5248
rect 840 5216 872 5248
rect 912 5216 944 5248
rect 984 5216 1016 5248
rect 1056 5216 1088 5248
rect 1128 5216 1160 5248
rect 1200 5216 1232 5248
rect 1272 5216 1304 5248
rect 1344 5216 1376 5248
rect 1416 5216 1448 5248
rect 1488 5216 1520 5248
rect 1560 5216 1592 5248
rect 1632 5216 1664 5248
rect 1704 5216 1736 5248
rect 1776 5216 1808 5248
rect 1848 5216 1880 5248
rect 1920 5216 1952 5248
rect 48 5144 80 5176
rect 120 5144 152 5176
rect 192 5144 224 5176
rect 264 5144 296 5176
rect 336 5144 368 5176
rect 408 5144 440 5176
rect 480 5144 512 5176
rect 552 5144 584 5176
rect 624 5144 656 5176
rect 696 5144 728 5176
rect 768 5144 800 5176
rect 840 5144 872 5176
rect 912 5144 944 5176
rect 984 5144 1016 5176
rect 1056 5144 1088 5176
rect 1128 5144 1160 5176
rect 1200 5144 1232 5176
rect 1272 5144 1304 5176
rect 1344 5144 1376 5176
rect 1416 5144 1448 5176
rect 1488 5144 1520 5176
rect 1560 5144 1592 5176
rect 1632 5144 1664 5176
rect 1704 5144 1736 5176
rect 1776 5144 1808 5176
rect 1848 5144 1880 5176
rect 1920 5144 1952 5176
rect 48 5072 80 5104
rect 120 5072 152 5104
rect 192 5072 224 5104
rect 264 5072 296 5104
rect 336 5072 368 5104
rect 408 5072 440 5104
rect 480 5072 512 5104
rect 552 5072 584 5104
rect 624 5072 656 5104
rect 696 5072 728 5104
rect 768 5072 800 5104
rect 840 5072 872 5104
rect 912 5072 944 5104
rect 984 5072 1016 5104
rect 1056 5072 1088 5104
rect 1128 5072 1160 5104
rect 1200 5072 1232 5104
rect 1272 5072 1304 5104
rect 1344 5072 1376 5104
rect 1416 5072 1448 5104
rect 1488 5072 1520 5104
rect 1560 5072 1592 5104
rect 1632 5072 1664 5104
rect 1704 5072 1736 5104
rect 1776 5072 1808 5104
rect 1848 5072 1880 5104
rect 1920 5072 1952 5104
rect 48 5000 80 5032
rect 120 5000 152 5032
rect 192 5000 224 5032
rect 264 5000 296 5032
rect 336 5000 368 5032
rect 408 5000 440 5032
rect 480 5000 512 5032
rect 552 5000 584 5032
rect 624 5000 656 5032
rect 696 5000 728 5032
rect 768 5000 800 5032
rect 840 5000 872 5032
rect 912 5000 944 5032
rect 984 5000 1016 5032
rect 1056 5000 1088 5032
rect 1128 5000 1160 5032
rect 1200 5000 1232 5032
rect 1272 5000 1304 5032
rect 1344 5000 1376 5032
rect 1416 5000 1448 5032
rect 1488 5000 1520 5032
rect 1560 5000 1592 5032
rect 1632 5000 1664 5032
rect 1704 5000 1736 5032
rect 1776 5000 1808 5032
rect 1848 5000 1880 5032
rect 1920 5000 1952 5032
rect 48 4928 80 4960
rect 120 4928 152 4960
rect 192 4928 224 4960
rect 264 4928 296 4960
rect 336 4928 368 4960
rect 408 4928 440 4960
rect 480 4928 512 4960
rect 552 4928 584 4960
rect 624 4928 656 4960
rect 696 4928 728 4960
rect 768 4928 800 4960
rect 840 4928 872 4960
rect 912 4928 944 4960
rect 984 4928 1016 4960
rect 1056 4928 1088 4960
rect 1128 4928 1160 4960
rect 1200 4928 1232 4960
rect 1272 4928 1304 4960
rect 1344 4928 1376 4960
rect 1416 4928 1448 4960
rect 1488 4928 1520 4960
rect 1560 4928 1592 4960
rect 1632 4928 1664 4960
rect 1704 4928 1736 4960
rect 1776 4928 1808 4960
rect 1848 4928 1880 4960
rect 1920 4928 1952 4960
rect 48 4856 80 4888
rect 120 4856 152 4888
rect 192 4856 224 4888
rect 264 4856 296 4888
rect 336 4856 368 4888
rect 408 4856 440 4888
rect 480 4856 512 4888
rect 552 4856 584 4888
rect 624 4856 656 4888
rect 696 4856 728 4888
rect 768 4856 800 4888
rect 840 4856 872 4888
rect 912 4856 944 4888
rect 984 4856 1016 4888
rect 1056 4856 1088 4888
rect 1128 4856 1160 4888
rect 1200 4856 1232 4888
rect 1272 4856 1304 4888
rect 1344 4856 1376 4888
rect 1416 4856 1448 4888
rect 1488 4856 1520 4888
rect 1560 4856 1592 4888
rect 1632 4856 1664 4888
rect 1704 4856 1736 4888
rect 1776 4856 1808 4888
rect 1848 4856 1880 4888
rect 1920 4856 1952 4888
rect 48 4784 80 4816
rect 120 4784 152 4816
rect 192 4784 224 4816
rect 264 4784 296 4816
rect 336 4784 368 4816
rect 408 4784 440 4816
rect 480 4784 512 4816
rect 552 4784 584 4816
rect 624 4784 656 4816
rect 696 4784 728 4816
rect 768 4784 800 4816
rect 840 4784 872 4816
rect 912 4784 944 4816
rect 984 4784 1016 4816
rect 1056 4784 1088 4816
rect 1128 4784 1160 4816
rect 1200 4784 1232 4816
rect 1272 4784 1304 4816
rect 1344 4784 1376 4816
rect 1416 4784 1448 4816
rect 1488 4784 1520 4816
rect 1560 4784 1592 4816
rect 1632 4784 1664 4816
rect 1704 4784 1736 4816
rect 1776 4784 1808 4816
rect 1848 4784 1880 4816
rect 1920 4784 1952 4816
rect 48 4712 80 4744
rect 120 4712 152 4744
rect 192 4712 224 4744
rect 264 4712 296 4744
rect 336 4712 368 4744
rect 408 4712 440 4744
rect 480 4712 512 4744
rect 552 4712 584 4744
rect 624 4712 656 4744
rect 696 4712 728 4744
rect 768 4712 800 4744
rect 840 4712 872 4744
rect 912 4712 944 4744
rect 984 4712 1016 4744
rect 1056 4712 1088 4744
rect 1128 4712 1160 4744
rect 1200 4712 1232 4744
rect 1272 4712 1304 4744
rect 1344 4712 1376 4744
rect 1416 4712 1448 4744
rect 1488 4712 1520 4744
rect 1560 4712 1592 4744
rect 1632 4712 1664 4744
rect 1704 4712 1736 4744
rect 1776 4712 1808 4744
rect 1848 4712 1880 4744
rect 1920 4712 1952 4744
rect 48 4640 80 4672
rect 120 4640 152 4672
rect 192 4640 224 4672
rect 264 4640 296 4672
rect 336 4640 368 4672
rect 408 4640 440 4672
rect 480 4640 512 4672
rect 552 4640 584 4672
rect 624 4640 656 4672
rect 696 4640 728 4672
rect 768 4640 800 4672
rect 840 4640 872 4672
rect 912 4640 944 4672
rect 984 4640 1016 4672
rect 1056 4640 1088 4672
rect 1128 4640 1160 4672
rect 1200 4640 1232 4672
rect 1272 4640 1304 4672
rect 1344 4640 1376 4672
rect 1416 4640 1448 4672
rect 1488 4640 1520 4672
rect 1560 4640 1592 4672
rect 1632 4640 1664 4672
rect 1704 4640 1736 4672
rect 1776 4640 1808 4672
rect 1848 4640 1880 4672
rect 1920 4640 1952 4672
rect 48 4568 80 4600
rect 120 4568 152 4600
rect 192 4568 224 4600
rect 264 4568 296 4600
rect 336 4568 368 4600
rect 408 4568 440 4600
rect 480 4568 512 4600
rect 552 4568 584 4600
rect 624 4568 656 4600
rect 696 4568 728 4600
rect 768 4568 800 4600
rect 840 4568 872 4600
rect 912 4568 944 4600
rect 984 4568 1016 4600
rect 1056 4568 1088 4600
rect 1128 4568 1160 4600
rect 1200 4568 1232 4600
rect 1272 4568 1304 4600
rect 1344 4568 1376 4600
rect 1416 4568 1448 4600
rect 1488 4568 1520 4600
rect 1560 4568 1592 4600
rect 1632 4568 1664 4600
rect 1704 4568 1736 4600
rect 1776 4568 1808 4600
rect 1848 4568 1880 4600
rect 1920 4568 1952 4600
rect 48 4496 80 4528
rect 120 4496 152 4528
rect 192 4496 224 4528
rect 264 4496 296 4528
rect 336 4496 368 4528
rect 408 4496 440 4528
rect 480 4496 512 4528
rect 552 4496 584 4528
rect 624 4496 656 4528
rect 696 4496 728 4528
rect 768 4496 800 4528
rect 840 4496 872 4528
rect 912 4496 944 4528
rect 984 4496 1016 4528
rect 1056 4496 1088 4528
rect 1128 4496 1160 4528
rect 1200 4496 1232 4528
rect 1272 4496 1304 4528
rect 1344 4496 1376 4528
rect 1416 4496 1448 4528
rect 1488 4496 1520 4528
rect 1560 4496 1592 4528
rect 1632 4496 1664 4528
rect 1704 4496 1736 4528
rect 1776 4496 1808 4528
rect 1848 4496 1880 4528
rect 1920 4496 1952 4528
rect 48 4424 80 4456
rect 120 4424 152 4456
rect 192 4424 224 4456
rect 264 4424 296 4456
rect 336 4424 368 4456
rect 408 4424 440 4456
rect 480 4424 512 4456
rect 552 4424 584 4456
rect 624 4424 656 4456
rect 696 4424 728 4456
rect 768 4424 800 4456
rect 840 4424 872 4456
rect 912 4424 944 4456
rect 984 4424 1016 4456
rect 1056 4424 1088 4456
rect 1128 4424 1160 4456
rect 1200 4424 1232 4456
rect 1272 4424 1304 4456
rect 1344 4424 1376 4456
rect 1416 4424 1448 4456
rect 1488 4424 1520 4456
rect 1560 4424 1592 4456
rect 1632 4424 1664 4456
rect 1704 4424 1736 4456
rect 1776 4424 1808 4456
rect 1848 4424 1880 4456
rect 1920 4424 1952 4456
rect 48 4352 80 4384
rect 120 4352 152 4384
rect 192 4352 224 4384
rect 264 4352 296 4384
rect 336 4352 368 4384
rect 408 4352 440 4384
rect 480 4352 512 4384
rect 552 4352 584 4384
rect 624 4352 656 4384
rect 696 4352 728 4384
rect 768 4352 800 4384
rect 840 4352 872 4384
rect 912 4352 944 4384
rect 984 4352 1016 4384
rect 1056 4352 1088 4384
rect 1128 4352 1160 4384
rect 1200 4352 1232 4384
rect 1272 4352 1304 4384
rect 1344 4352 1376 4384
rect 1416 4352 1448 4384
rect 1488 4352 1520 4384
rect 1560 4352 1592 4384
rect 1632 4352 1664 4384
rect 1704 4352 1736 4384
rect 1776 4352 1808 4384
rect 1848 4352 1880 4384
rect 1920 4352 1952 4384
rect 48 4280 80 4312
rect 120 4280 152 4312
rect 192 4280 224 4312
rect 264 4280 296 4312
rect 336 4280 368 4312
rect 408 4280 440 4312
rect 480 4280 512 4312
rect 552 4280 584 4312
rect 624 4280 656 4312
rect 696 4280 728 4312
rect 768 4280 800 4312
rect 840 4280 872 4312
rect 912 4280 944 4312
rect 984 4280 1016 4312
rect 1056 4280 1088 4312
rect 1128 4280 1160 4312
rect 1200 4280 1232 4312
rect 1272 4280 1304 4312
rect 1344 4280 1376 4312
rect 1416 4280 1448 4312
rect 1488 4280 1520 4312
rect 1560 4280 1592 4312
rect 1632 4280 1664 4312
rect 1704 4280 1736 4312
rect 1776 4280 1808 4312
rect 1848 4280 1880 4312
rect 1920 4280 1952 4312
rect 48 4208 80 4240
rect 120 4208 152 4240
rect 192 4208 224 4240
rect 264 4208 296 4240
rect 336 4208 368 4240
rect 408 4208 440 4240
rect 480 4208 512 4240
rect 552 4208 584 4240
rect 624 4208 656 4240
rect 696 4208 728 4240
rect 768 4208 800 4240
rect 840 4208 872 4240
rect 912 4208 944 4240
rect 984 4208 1016 4240
rect 1056 4208 1088 4240
rect 1128 4208 1160 4240
rect 1200 4208 1232 4240
rect 1272 4208 1304 4240
rect 1344 4208 1376 4240
rect 1416 4208 1448 4240
rect 1488 4208 1520 4240
rect 1560 4208 1592 4240
rect 1632 4208 1664 4240
rect 1704 4208 1736 4240
rect 1776 4208 1808 4240
rect 1848 4208 1880 4240
rect 1920 4208 1952 4240
rect 48 4136 80 4168
rect 120 4136 152 4168
rect 192 4136 224 4168
rect 264 4136 296 4168
rect 336 4136 368 4168
rect 408 4136 440 4168
rect 480 4136 512 4168
rect 552 4136 584 4168
rect 624 4136 656 4168
rect 696 4136 728 4168
rect 768 4136 800 4168
rect 840 4136 872 4168
rect 912 4136 944 4168
rect 984 4136 1016 4168
rect 1056 4136 1088 4168
rect 1128 4136 1160 4168
rect 1200 4136 1232 4168
rect 1272 4136 1304 4168
rect 1344 4136 1376 4168
rect 1416 4136 1448 4168
rect 1488 4136 1520 4168
rect 1560 4136 1592 4168
rect 1632 4136 1664 4168
rect 1704 4136 1736 4168
rect 1776 4136 1808 4168
rect 1848 4136 1880 4168
rect 1920 4136 1952 4168
rect 48 4064 80 4096
rect 120 4064 152 4096
rect 192 4064 224 4096
rect 264 4064 296 4096
rect 336 4064 368 4096
rect 408 4064 440 4096
rect 480 4064 512 4096
rect 552 4064 584 4096
rect 624 4064 656 4096
rect 696 4064 728 4096
rect 768 4064 800 4096
rect 840 4064 872 4096
rect 912 4064 944 4096
rect 984 4064 1016 4096
rect 1056 4064 1088 4096
rect 1128 4064 1160 4096
rect 1200 4064 1232 4096
rect 1272 4064 1304 4096
rect 1344 4064 1376 4096
rect 1416 4064 1448 4096
rect 1488 4064 1520 4096
rect 1560 4064 1592 4096
rect 1632 4064 1664 4096
rect 1704 4064 1736 4096
rect 1776 4064 1808 4096
rect 1848 4064 1880 4096
rect 1920 4064 1952 4096
rect 48 3992 80 4024
rect 120 3992 152 4024
rect 192 3992 224 4024
rect 264 3992 296 4024
rect 336 3992 368 4024
rect 408 3992 440 4024
rect 480 3992 512 4024
rect 552 3992 584 4024
rect 624 3992 656 4024
rect 696 3992 728 4024
rect 768 3992 800 4024
rect 840 3992 872 4024
rect 912 3992 944 4024
rect 984 3992 1016 4024
rect 1056 3992 1088 4024
rect 1128 3992 1160 4024
rect 1200 3992 1232 4024
rect 1272 3992 1304 4024
rect 1344 3992 1376 4024
rect 1416 3992 1448 4024
rect 1488 3992 1520 4024
rect 1560 3992 1592 4024
rect 1632 3992 1664 4024
rect 1704 3992 1736 4024
rect 1776 3992 1808 4024
rect 1848 3992 1880 4024
rect 1920 3992 1952 4024
rect 48 3920 80 3952
rect 120 3920 152 3952
rect 192 3920 224 3952
rect 264 3920 296 3952
rect 336 3920 368 3952
rect 408 3920 440 3952
rect 480 3920 512 3952
rect 552 3920 584 3952
rect 624 3920 656 3952
rect 696 3920 728 3952
rect 768 3920 800 3952
rect 840 3920 872 3952
rect 912 3920 944 3952
rect 984 3920 1016 3952
rect 1056 3920 1088 3952
rect 1128 3920 1160 3952
rect 1200 3920 1232 3952
rect 1272 3920 1304 3952
rect 1344 3920 1376 3952
rect 1416 3920 1448 3952
rect 1488 3920 1520 3952
rect 1560 3920 1592 3952
rect 1632 3920 1664 3952
rect 1704 3920 1736 3952
rect 1776 3920 1808 3952
rect 1848 3920 1880 3952
rect 1920 3920 1952 3952
rect 48 3848 80 3880
rect 120 3848 152 3880
rect 192 3848 224 3880
rect 264 3848 296 3880
rect 336 3848 368 3880
rect 408 3848 440 3880
rect 480 3848 512 3880
rect 552 3848 584 3880
rect 624 3848 656 3880
rect 696 3848 728 3880
rect 768 3848 800 3880
rect 840 3848 872 3880
rect 912 3848 944 3880
rect 984 3848 1016 3880
rect 1056 3848 1088 3880
rect 1128 3848 1160 3880
rect 1200 3848 1232 3880
rect 1272 3848 1304 3880
rect 1344 3848 1376 3880
rect 1416 3848 1448 3880
rect 1488 3848 1520 3880
rect 1560 3848 1592 3880
rect 1632 3848 1664 3880
rect 1704 3848 1736 3880
rect 1776 3848 1808 3880
rect 1848 3848 1880 3880
rect 1920 3848 1952 3880
rect 48 3776 80 3808
rect 120 3776 152 3808
rect 192 3776 224 3808
rect 264 3776 296 3808
rect 336 3776 368 3808
rect 408 3776 440 3808
rect 480 3776 512 3808
rect 552 3776 584 3808
rect 624 3776 656 3808
rect 696 3776 728 3808
rect 768 3776 800 3808
rect 840 3776 872 3808
rect 912 3776 944 3808
rect 984 3776 1016 3808
rect 1056 3776 1088 3808
rect 1128 3776 1160 3808
rect 1200 3776 1232 3808
rect 1272 3776 1304 3808
rect 1344 3776 1376 3808
rect 1416 3776 1448 3808
rect 1488 3776 1520 3808
rect 1560 3776 1592 3808
rect 1632 3776 1664 3808
rect 1704 3776 1736 3808
rect 1776 3776 1808 3808
rect 1848 3776 1880 3808
rect 1920 3776 1952 3808
rect 48 3704 80 3736
rect 120 3704 152 3736
rect 192 3704 224 3736
rect 264 3704 296 3736
rect 336 3704 368 3736
rect 408 3704 440 3736
rect 480 3704 512 3736
rect 552 3704 584 3736
rect 624 3704 656 3736
rect 696 3704 728 3736
rect 768 3704 800 3736
rect 840 3704 872 3736
rect 912 3704 944 3736
rect 984 3704 1016 3736
rect 1056 3704 1088 3736
rect 1128 3704 1160 3736
rect 1200 3704 1232 3736
rect 1272 3704 1304 3736
rect 1344 3704 1376 3736
rect 1416 3704 1448 3736
rect 1488 3704 1520 3736
rect 1560 3704 1592 3736
rect 1632 3704 1664 3736
rect 1704 3704 1736 3736
rect 1776 3704 1808 3736
rect 1848 3704 1880 3736
rect 1920 3704 1952 3736
rect 48 3632 80 3664
rect 120 3632 152 3664
rect 192 3632 224 3664
rect 264 3632 296 3664
rect 336 3632 368 3664
rect 408 3632 440 3664
rect 480 3632 512 3664
rect 552 3632 584 3664
rect 624 3632 656 3664
rect 696 3632 728 3664
rect 768 3632 800 3664
rect 840 3632 872 3664
rect 912 3632 944 3664
rect 984 3632 1016 3664
rect 1056 3632 1088 3664
rect 1128 3632 1160 3664
rect 1200 3632 1232 3664
rect 1272 3632 1304 3664
rect 1344 3632 1376 3664
rect 1416 3632 1448 3664
rect 1488 3632 1520 3664
rect 1560 3632 1592 3664
rect 1632 3632 1664 3664
rect 1704 3632 1736 3664
rect 1776 3632 1808 3664
rect 1848 3632 1880 3664
rect 1920 3632 1952 3664
rect 48 3560 80 3592
rect 120 3560 152 3592
rect 192 3560 224 3592
rect 264 3560 296 3592
rect 336 3560 368 3592
rect 408 3560 440 3592
rect 480 3560 512 3592
rect 552 3560 584 3592
rect 624 3560 656 3592
rect 696 3560 728 3592
rect 768 3560 800 3592
rect 840 3560 872 3592
rect 912 3560 944 3592
rect 984 3560 1016 3592
rect 1056 3560 1088 3592
rect 1128 3560 1160 3592
rect 1200 3560 1232 3592
rect 1272 3560 1304 3592
rect 1344 3560 1376 3592
rect 1416 3560 1448 3592
rect 1488 3560 1520 3592
rect 1560 3560 1592 3592
rect 1632 3560 1664 3592
rect 1704 3560 1736 3592
rect 1776 3560 1808 3592
rect 1848 3560 1880 3592
rect 1920 3560 1952 3592
rect 48 3488 80 3520
rect 120 3488 152 3520
rect 192 3488 224 3520
rect 264 3488 296 3520
rect 336 3488 368 3520
rect 408 3488 440 3520
rect 480 3488 512 3520
rect 552 3488 584 3520
rect 624 3488 656 3520
rect 696 3488 728 3520
rect 768 3488 800 3520
rect 840 3488 872 3520
rect 912 3488 944 3520
rect 984 3488 1016 3520
rect 1056 3488 1088 3520
rect 1128 3488 1160 3520
rect 1200 3488 1232 3520
rect 1272 3488 1304 3520
rect 1344 3488 1376 3520
rect 1416 3488 1448 3520
rect 1488 3488 1520 3520
rect 1560 3488 1592 3520
rect 1632 3488 1664 3520
rect 1704 3488 1736 3520
rect 1776 3488 1808 3520
rect 1848 3488 1880 3520
rect 1920 3488 1952 3520
rect 48 3416 80 3448
rect 120 3416 152 3448
rect 192 3416 224 3448
rect 264 3416 296 3448
rect 336 3416 368 3448
rect 408 3416 440 3448
rect 480 3416 512 3448
rect 552 3416 584 3448
rect 624 3416 656 3448
rect 696 3416 728 3448
rect 768 3416 800 3448
rect 840 3416 872 3448
rect 912 3416 944 3448
rect 984 3416 1016 3448
rect 1056 3416 1088 3448
rect 1128 3416 1160 3448
rect 1200 3416 1232 3448
rect 1272 3416 1304 3448
rect 1344 3416 1376 3448
rect 1416 3416 1448 3448
rect 1488 3416 1520 3448
rect 1560 3416 1592 3448
rect 1632 3416 1664 3448
rect 1704 3416 1736 3448
rect 1776 3416 1808 3448
rect 1848 3416 1880 3448
rect 1920 3416 1952 3448
rect 48 3344 80 3376
rect 120 3344 152 3376
rect 192 3344 224 3376
rect 264 3344 296 3376
rect 336 3344 368 3376
rect 408 3344 440 3376
rect 480 3344 512 3376
rect 552 3344 584 3376
rect 624 3344 656 3376
rect 696 3344 728 3376
rect 768 3344 800 3376
rect 840 3344 872 3376
rect 912 3344 944 3376
rect 984 3344 1016 3376
rect 1056 3344 1088 3376
rect 1128 3344 1160 3376
rect 1200 3344 1232 3376
rect 1272 3344 1304 3376
rect 1344 3344 1376 3376
rect 1416 3344 1448 3376
rect 1488 3344 1520 3376
rect 1560 3344 1592 3376
rect 1632 3344 1664 3376
rect 1704 3344 1736 3376
rect 1776 3344 1808 3376
rect 1848 3344 1880 3376
rect 1920 3344 1952 3376
rect 48 3272 80 3304
rect 120 3272 152 3304
rect 192 3272 224 3304
rect 264 3272 296 3304
rect 336 3272 368 3304
rect 408 3272 440 3304
rect 480 3272 512 3304
rect 552 3272 584 3304
rect 624 3272 656 3304
rect 696 3272 728 3304
rect 768 3272 800 3304
rect 840 3272 872 3304
rect 912 3272 944 3304
rect 984 3272 1016 3304
rect 1056 3272 1088 3304
rect 1128 3272 1160 3304
rect 1200 3272 1232 3304
rect 1272 3272 1304 3304
rect 1344 3272 1376 3304
rect 1416 3272 1448 3304
rect 1488 3272 1520 3304
rect 1560 3272 1592 3304
rect 1632 3272 1664 3304
rect 1704 3272 1736 3304
rect 1776 3272 1808 3304
rect 1848 3272 1880 3304
rect 1920 3272 1952 3304
rect 48 3200 80 3232
rect 120 3200 152 3232
rect 192 3200 224 3232
rect 264 3200 296 3232
rect 336 3200 368 3232
rect 408 3200 440 3232
rect 480 3200 512 3232
rect 552 3200 584 3232
rect 624 3200 656 3232
rect 696 3200 728 3232
rect 768 3200 800 3232
rect 840 3200 872 3232
rect 912 3200 944 3232
rect 984 3200 1016 3232
rect 1056 3200 1088 3232
rect 1128 3200 1160 3232
rect 1200 3200 1232 3232
rect 1272 3200 1304 3232
rect 1344 3200 1376 3232
rect 1416 3200 1448 3232
rect 1488 3200 1520 3232
rect 1560 3200 1592 3232
rect 1632 3200 1664 3232
rect 1704 3200 1736 3232
rect 1776 3200 1808 3232
rect 1848 3200 1880 3232
rect 1920 3200 1952 3232
rect 48 3128 80 3160
rect 120 3128 152 3160
rect 192 3128 224 3160
rect 264 3128 296 3160
rect 336 3128 368 3160
rect 408 3128 440 3160
rect 480 3128 512 3160
rect 552 3128 584 3160
rect 624 3128 656 3160
rect 696 3128 728 3160
rect 768 3128 800 3160
rect 840 3128 872 3160
rect 912 3128 944 3160
rect 984 3128 1016 3160
rect 1056 3128 1088 3160
rect 1128 3128 1160 3160
rect 1200 3128 1232 3160
rect 1272 3128 1304 3160
rect 1344 3128 1376 3160
rect 1416 3128 1448 3160
rect 1488 3128 1520 3160
rect 1560 3128 1592 3160
rect 1632 3128 1664 3160
rect 1704 3128 1736 3160
rect 1776 3128 1808 3160
rect 1848 3128 1880 3160
rect 1920 3128 1952 3160
rect 48 3056 80 3088
rect 120 3056 152 3088
rect 192 3056 224 3088
rect 264 3056 296 3088
rect 336 3056 368 3088
rect 408 3056 440 3088
rect 480 3056 512 3088
rect 552 3056 584 3088
rect 624 3056 656 3088
rect 696 3056 728 3088
rect 768 3056 800 3088
rect 840 3056 872 3088
rect 912 3056 944 3088
rect 984 3056 1016 3088
rect 1056 3056 1088 3088
rect 1128 3056 1160 3088
rect 1200 3056 1232 3088
rect 1272 3056 1304 3088
rect 1344 3056 1376 3088
rect 1416 3056 1448 3088
rect 1488 3056 1520 3088
rect 1560 3056 1592 3088
rect 1632 3056 1664 3088
rect 1704 3056 1736 3088
rect 1776 3056 1808 3088
rect 1848 3056 1880 3088
rect 1920 3056 1952 3088
rect 48 2984 80 3016
rect 120 2984 152 3016
rect 192 2984 224 3016
rect 264 2984 296 3016
rect 336 2984 368 3016
rect 408 2984 440 3016
rect 480 2984 512 3016
rect 552 2984 584 3016
rect 624 2984 656 3016
rect 696 2984 728 3016
rect 768 2984 800 3016
rect 840 2984 872 3016
rect 912 2984 944 3016
rect 984 2984 1016 3016
rect 1056 2984 1088 3016
rect 1128 2984 1160 3016
rect 1200 2984 1232 3016
rect 1272 2984 1304 3016
rect 1344 2984 1376 3016
rect 1416 2984 1448 3016
rect 1488 2984 1520 3016
rect 1560 2984 1592 3016
rect 1632 2984 1664 3016
rect 1704 2984 1736 3016
rect 1776 2984 1808 3016
rect 1848 2984 1880 3016
rect 1920 2984 1952 3016
rect 48 2912 80 2944
rect 120 2912 152 2944
rect 192 2912 224 2944
rect 264 2912 296 2944
rect 336 2912 368 2944
rect 408 2912 440 2944
rect 480 2912 512 2944
rect 552 2912 584 2944
rect 624 2912 656 2944
rect 696 2912 728 2944
rect 768 2912 800 2944
rect 840 2912 872 2944
rect 912 2912 944 2944
rect 984 2912 1016 2944
rect 1056 2912 1088 2944
rect 1128 2912 1160 2944
rect 1200 2912 1232 2944
rect 1272 2912 1304 2944
rect 1344 2912 1376 2944
rect 1416 2912 1448 2944
rect 1488 2912 1520 2944
rect 1560 2912 1592 2944
rect 1632 2912 1664 2944
rect 1704 2912 1736 2944
rect 1776 2912 1808 2944
rect 1848 2912 1880 2944
rect 1920 2912 1952 2944
rect 48 2840 80 2872
rect 120 2840 152 2872
rect 192 2840 224 2872
rect 264 2840 296 2872
rect 336 2840 368 2872
rect 408 2840 440 2872
rect 480 2840 512 2872
rect 552 2840 584 2872
rect 624 2840 656 2872
rect 696 2840 728 2872
rect 768 2840 800 2872
rect 840 2840 872 2872
rect 912 2840 944 2872
rect 984 2840 1016 2872
rect 1056 2840 1088 2872
rect 1128 2840 1160 2872
rect 1200 2840 1232 2872
rect 1272 2840 1304 2872
rect 1344 2840 1376 2872
rect 1416 2840 1448 2872
rect 1488 2840 1520 2872
rect 1560 2840 1592 2872
rect 1632 2840 1664 2872
rect 1704 2840 1736 2872
rect 1776 2840 1808 2872
rect 1848 2840 1880 2872
rect 1920 2840 1952 2872
rect 48 2768 80 2800
rect 120 2768 152 2800
rect 192 2768 224 2800
rect 264 2768 296 2800
rect 336 2768 368 2800
rect 408 2768 440 2800
rect 480 2768 512 2800
rect 552 2768 584 2800
rect 624 2768 656 2800
rect 696 2768 728 2800
rect 768 2768 800 2800
rect 840 2768 872 2800
rect 912 2768 944 2800
rect 984 2768 1016 2800
rect 1056 2768 1088 2800
rect 1128 2768 1160 2800
rect 1200 2768 1232 2800
rect 1272 2768 1304 2800
rect 1344 2768 1376 2800
rect 1416 2768 1448 2800
rect 1488 2768 1520 2800
rect 1560 2768 1592 2800
rect 1632 2768 1664 2800
rect 1704 2768 1736 2800
rect 1776 2768 1808 2800
rect 1848 2768 1880 2800
rect 1920 2768 1952 2800
rect 48 2696 80 2728
rect 120 2696 152 2728
rect 192 2696 224 2728
rect 264 2696 296 2728
rect 336 2696 368 2728
rect 408 2696 440 2728
rect 480 2696 512 2728
rect 552 2696 584 2728
rect 624 2696 656 2728
rect 696 2696 728 2728
rect 768 2696 800 2728
rect 840 2696 872 2728
rect 912 2696 944 2728
rect 984 2696 1016 2728
rect 1056 2696 1088 2728
rect 1128 2696 1160 2728
rect 1200 2696 1232 2728
rect 1272 2696 1304 2728
rect 1344 2696 1376 2728
rect 1416 2696 1448 2728
rect 1488 2696 1520 2728
rect 1560 2696 1592 2728
rect 1632 2696 1664 2728
rect 1704 2696 1736 2728
rect 1776 2696 1808 2728
rect 1848 2696 1880 2728
rect 1920 2696 1952 2728
rect 48 2624 80 2656
rect 120 2624 152 2656
rect 192 2624 224 2656
rect 264 2624 296 2656
rect 336 2624 368 2656
rect 408 2624 440 2656
rect 480 2624 512 2656
rect 552 2624 584 2656
rect 624 2624 656 2656
rect 696 2624 728 2656
rect 768 2624 800 2656
rect 840 2624 872 2656
rect 912 2624 944 2656
rect 984 2624 1016 2656
rect 1056 2624 1088 2656
rect 1128 2624 1160 2656
rect 1200 2624 1232 2656
rect 1272 2624 1304 2656
rect 1344 2624 1376 2656
rect 1416 2624 1448 2656
rect 1488 2624 1520 2656
rect 1560 2624 1592 2656
rect 1632 2624 1664 2656
rect 1704 2624 1736 2656
rect 1776 2624 1808 2656
rect 1848 2624 1880 2656
rect 1920 2624 1952 2656
rect 48 2552 80 2584
rect 120 2552 152 2584
rect 192 2552 224 2584
rect 264 2552 296 2584
rect 336 2552 368 2584
rect 408 2552 440 2584
rect 480 2552 512 2584
rect 552 2552 584 2584
rect 624 2552 656 2584
rect 696 2552 728 2584
rect 768 2552 800 2584
rect 840 2552 872 2584
rect 912 2552 944 2584
rect 984 2552 1016 2584
rect 1056 2552 1088 2584
rect 1128 2552 1160 2584
rect 1200 2552 1232 2584
rect 1272 2552 1304 2584
rect 1344 2552 1376 2584
rect 1416 2552 1448 2584
rect 1488 2552 1520 2584
rect 1560 2552 1592 2584
rect 1632 2552 1664 2584
rect 1704 2552 1736 2584
rect 1776 2552 1808 2584
rect 1848 2552 1880 2584
rect 1920 2552 1952 2584
rect 48 2480 80 2512
rect 120 2480 152 2512
rect 192 2480 224 2512
rect 264 2480 296 2512
rect 336 2480 368 2512
rect 408 2480 440 2512
rect 480 2480 512 2512
rect 552 2480 584 2512
rect 624 2480 656 2512
rect 696 2480 728 2512
rect 768 2480 800 2512
rect 840 2480 872 2512
rect 912 2480 944 2512
rect 984 2480 1016 2512
rect 1056 2480 1088 2512
rect 1128 2480 1160 2512
rect 1200 2480 1232 2512
rect 1272 2480 1304 2512
rect 1344 2480 1376 2512
rect 1416 2480 1448 2512
rect 1488 2480 1520 2512
rect 1560 2480 1592 2512
rect 1632 2480 1664 2512
rect 1704 2480 1736 2512
rect 1776 2480 1808 2512
rect 1848 2480 1880 2512
rect 1920 2480 1952 2512
rect 48 2408 80 2440
rect 120 2408 152 2440
rect 192 2408 224 2440
rect 264 2408 296 2440
rect 336 2408 368 2440
rect 408 2408 440 2440
rect 480 2408 512 2440
rect 552 2408 584 2440
rect 624 2408 656 2440
rect 696 2408 728 2440
rect 768 2408 800 2440
rect 840 2408 872 2440
rect 912 2408 944 2440
rect 984 2408 1016 2440
rect 1056 2408 1088 2440
rect 1128 2408 1160 2440
rect 1200 2408 1232 2440
rect 1272 2408 1304 2440
rect 1344 2408 1376 2440
rect 1416 2408 1448 2440
rect 1488 2408 1520 2440
rect 1560 2408 1592 2440
rect 1632 2408 1664 2440
rect 1704 2408 1736 2440
rect 1776 2408 1808 2440
rect 1848 2408 1880 2440
rect 1920 2408 1952 2440
rect 48 2336 80 2368
rect 120 2336 152 2368
rect 192 2336 224 2368
rect 264 2336 296 2368
rect 336 2336 368 2368
rect 408 2336 440 2368
rect 480 2336 512 2368
rect 552 2336 584 2368
rect 624 2336 656 2368
rect 696 2336 728 2368
rect 768 2336 800 2368
rect 840 2336 872 2368
rect 912 2336 944 2368
rect 984 2336 1016 2368
rect 1056 2336 1088 2368
rect 1128 2336 1160 2368
rect 1200 2336 1232 2368
rect 1272 2336 1304 2368
rect 1344 2336 1376 2368
rect 1416 2336 1448 2368
rect 1488 2336 1520 2368
rect 1560 2336 1592 2368
rect 1632 2336 1664 2368
rect 1704 2336 1736 2368
rect 1776 2336 1808 2368
rect 1848 2336 1880 2368
rect 1920 2336 1952 2368
rect 48 2264 80 2296
rect 120 2264 152 2296
rect 192 2264 224 2296
rect 264 2264 296 2296
rect 336 2264 368 2296
rect 408 2264 440 2296
rect 480 2264 512 2296
rect 552 2264 584 2296
rect 624 2264 656 2296
rect 696 2264 728 2296
rect 768 2264 800 2296
rect 840 2264 872 2296
rect 912 2264 944 2296
rect 984 2264 1016 2296
rect 1056 2264 1088 2296
rect 1128 2264 1160 2296
rect 1200 2264 1232 2296
rect 1272 2264 1304 2296
rect 1344 2264 1376 2296
rect 1416 2264 1448 2296
rect 1488 2264 1520 2296
rect 1560 2264 1592 2296
rect 1632 2264 1664 2296
rect 1704 2264 1736 2296
rect 1776 2264 1808 2296
rect 1848 2264 1880 2296
rect 1920 2264 1952 2296
rect 48 2192 80 2224
rect 120 2192 152 2224
rect 192 2192 224 2224
rect 264 2192 296 2224
rect 336 2192 368 2224
rect 408 2192 440 2224
rect 480 2192 512 2224
rect 552 2192 584 2224
rect 624 2192 656 2224
rect 696 2192 728 2224
rect 768 2192 800 2224
rect 840 2192 872 2224
rect 912 2192 944 2224
rect 984 2192 1016 2224
rect 1056 2192 1088 2224
rect 1128 2192 1160 2224
rect 1200 2192 1232 2224
rect 1272 2192 1304 2224
rect 1344 2192 1376 2224
rect 1416 2192 1448 2224
rect 1488 2192 1520 2224
rect 1560 2192 1592 2224
rect 1632 2192 1664 2224
rect 1704 2192 1736 2224
rect 1776 2192 1808 2224
rect 1848 2192 1880 2224
rect 1920 2192 1952 2224
rect 48 2120 80 2152
rect 120 2120 152 2152
rect 192 2120 224 2152
rect 264 2120 296 2152
rect 336 2120 368 2152
rect 408 2120 440 2152
rect 480 2120 512 2152
rect 552 2120 584 2152
rect 624 2120 656 2152
rect 696 2120 728 2152
rect 768 2120 800 2152
rect 840 2120 872 2152
rect 912 2120 944 2152
rect 984 2120 1016 2152
rect 1056 2120 1088 2152
rect 1128 2120 1160 2152
rect 1200 2120 1232 2152
rect 1272 2120 1304 2152
rect 1344 2120 1376 2152
rect 1416 2120 1448 2152
rect 1488 2120 1520 2152
rect 1560 2120 1592 2152
rect 1632 2120 1664 2152
rect 1704 2120 1736 2152
rect 1776 2120 1808 2152
rect 1848 2120 1880 2152
rect 1920 2120 1952 2152
rect 48 2048 80 2080
rect 120 2048 152 2080
rect 192 2048 224 2080
rect 264 2048 296 2080
rect 336 2048 368 2080
rect 408 2048 440 2080
rect 480 2048 512 2080
rect 552 2048 584 2080
rect 624 2048 656 2080
rect 696 2048 728 2080
rect 768 2048 800 2080
rect 840 2048 872 2080
rect 912 2048 944 2080
rect 984 2048 1016 2080
rect 1056 2048 1088 2080
rect 1128 2048 1160 2080
rect 1200 2048 1232 2080
rect 1272 2048 1304 2080
rect 1344 2048 1376 2080
rect 1416 2048 1448 2080
rect 1488 2048 1520 2080
rect 1560 2048 1592 2080
rect 1632 2048 1664 2080
rect 1704 2048 1736 2080
rect 1776 2048 1808 2080
rect 1848 2048 1880 2080
rect 1920 2048 1952 2080
rect 48 1976 80 2008
rect 120 1976 152 2008
rect 192 1976 224 2008
rect 264 1976 296 2008
rect 336 1976 368 2008
rect 408 1976 440 2008
rect 480 1976 512 2008
rect 552 1976 584 2008
rect 624 1976 656 2008
rect 696 1976 728 2008
rect 768 1976 800 2008
rect 840 1976 872 2008
rect 912 1976 944 2008
rect 984 1976 1016 2008
rect 1056 1976 1088 2008
rect 1128 1976 1160 2008
rect 1200 1976 1232 2008
rect 1272 1976 1304 2008
rect 1344 1976 1376 2008
rect 1416 1976 1448 2008
rect 1488 1976 1520 2008
rect 1560 1976 1592 2008
rect 1632 1976 1664 2008
rect 1704 1976 1736 2008
rect 1776 1976 1808 2008
rect 1848 1976 1880 2008
rect 1920 1976 1952 2008
rect 48 1904 80 1936
rect 120 1904 152 1936
rect 192 1904 224 1936
rect 264 1904 296 1936
rect 336 1904 368 1936
rect 408 1904 440 1936
rect 480 1904 512 1936
rect 552 1904 584 1936
rect 624 1904 656 1936
rect 696 1904 728 1936
rect 768 1904 800 1936
rect 840 1904 872 1936
rect 912 1904 944 1936
rect 984 1904 1016 1936
rect 1056 1904 1088 1936
rect 1128 1904 1160 1936
rect 1200 1904 1232 1936
rect 1272 1904 1304 1936
rect 1344 1904 1376 1936
rect 1416 1904 1448 1936
rect 1488 1904 1520 1936
rect 1560 1904 1592 1936
rect 1632 1904 1664 1936
rect 1704 1904 1736 1936
rect 1776 1904 1808 1936
rect 1848 1904 1880 1936
rect 1920 1904 1952 1936
rect 48 1832 80 1864
rect 120 1832 152 1864
rect 192 1832 224 1864
rect 264 1832 296 1864
rect 336 1832 368 1864
rect 408 1832 440 1864
rect 480 1832 512 1864
rect 552 1832 584 1864
rect 624 1832 656 1864
rect 696 1832 728 1864
rect 768 1832 800 1864
rect 840 1832 872 1864
rect 912 1832 944 1864
rect 984 1832 1016 1864
rect 1056 1832 1088 1864
rect 1128 1832 1160 1864
rect 1200 1832 1232 1864
rect 1272 1832 1304 1864
rect 1344 1832 1376 1864
rect 1416 1832 1448 1864
rect 1488 1832 1520 1864
rect 1560 1832 1592 1864
rect 1632 1832 1664 1864
rect 1704 1832 1736 1864
rect 1776 1832 1808 1864
rect 1848 1832 1880 1864
rect 1920 1832 1952 1864
rect 48 1760 80 1792
rect 120 1760 152 1792
rect 192 1760 224 1792
rect 264 1760 296 1792
rect 336 1760 368 1792
rect 408 1760 440 1792
rect 480 1760 512 1792
rect 552 1760 584 1792
rect 624 1760 656 1792
rect 696 1760 728 1792
rect 768 1760 800 1792
rect 840 1760 872 1792
rect 912 1760 944 1792
rect 984 1760 1016 1792
rect 1056 1760 1088 1792
rect 1128 1760 1160 1792
rect 1200 1760 1232 1792
rect 1272 1760 1304 1792
rect 1344 1760 1376 1792
rect 1416 1760 1448 1792
rect 1488 1760 1520 1792
rect 1560 1760 1592 1792
rect 1632 1760 1664 1792
rect 1704 1760 1736 1792
rect 1776 1760 1808 1792
rect 1848 1760 1880 1792
rect 1920 1760 1952 1792
rect 48 1688 80 1720
rect 120 1688 152 1720
rect 192 1688 224 1720
rect 264 1688 296 1720
rect 336 1688 368 1720
rect 408 1688 440 1720
rect 480 1688 512 1720
rect 552 1688 584 1720
rect 624 1688 656 1720
rect 696 1688 728 1720
rect 768 1688 800 1720
rect 840 1688 872 1720
rect 912 1688 944 1720
rect 984 1688 1016 1720
rect 1056 1688 1088 1720
rect 1128 1688 1160 1720
rect 1200 1688 1232 1720
rect 1272 1688 1304 1720
rect 1344 1688 1376 1720
rect 1416 1688 1448 1720
rect 1488 1688 1520 1720
rect 1560 1688 1592 1720
rect 1632 1688 1664 1720
rect 1704 1688 1736 1720
rect 1776 1688 1808 1720
rect 1848 1688 1880 1720
rect 1920 1688 1952 1720
rect 48 1616 80 1648
rect 120 1616 152 1648
rect 192 1616 224 1648
rect 264 1616 296 1648
rect 336 1616 368 1648
rect 408 1616 440 1648
rect 480 1616 512 1648
rect 552 1616 584 1648
rect 624 1616 656 1648
rect 696 1616 728 1648
rect 768 1616 800 1648
rect 840 1616 872 1648
rect 912 1616 944 1648
rect 984 1616 1016 1648
rect 1056 1616 1088 1648
rect 1128 1616 1160 1648
rect 1200 1616 1232 1648
rect 1272 1616 1304 1648
rect 1344 1616 1376 1648
rect 1416 1616 1448 1648
rect 1488 1616 1520 1648
rect 1560 1616 1592 1648
rect 1632 1616 1664 1648
rect 1704 1616 1736 1648
rect 1776 1616 1808 1648
rect 1848 1616 1880 1648
rect 1920 1616 1952 1648
rect 48 1544 80 1576
rect 120 1544 152 1576
rect 192 1544 224 1576
rect 264 1544 296 1576
rect 336 1544 368 1576
rect 408 1544 440 1576
rect 480 1544 512 1576
rect 552 1544 584 1576
rect 624 1544 656 1576
rect 696 1544 728 1576
rect 768 1544 800 1576
rect 840 1544 872 1576
rect 912 1544 944 1576
rect 984 1544 1016 1576
rect 1056 1544 1088 1576
rect 1128 1544 1160 1576
rect 1200 1544 1232 1576
rect 1272 1544 1304 1576
rect 1344 1544 1376 1576
rect 1416 1544 1448 1576
rect 1488 1544 1520 1576
rect 1560 1544 1592 1576
rect 1632 1544 1664 1576
rect 1704 1544 1736 1576
rect 1776 1544 1808 1576
rect 1848 1544 1880 1576
rect 1920 1544 1952 1576
rect 48 1472 80 1504
rect 120 1472 152 1504
rect 192 1472 224 1504
rect 264 1472 296 1504
rect 336 1472 368 1504
rect 408 1472 440 1504
rect 480 1472 512 1504
rect 552 1472 584 1504
rect 624 1472 656 1504
rect 696 1472 728 1504
rect 768 1472 800 1504
rect 840 1472 872 1504
rect 912 1472 944 1504
rect 984 1472 1016 1504
rect 1056 1472 1088 1504
rect 1128 1472 1160 1504
rect 1200 1472 1232 1504
rect 1272 1472 1304 1504
rect 1344 1472 1376 1504
rect 1416 1472 1448 1504
rect 1488 1472 1520 1504
rect 1560 1472 1592 1504
rect 1632 1472 1664 1504
rect 1704 1472 1736 1504
rect 1776 1472 1808 1504
rect 1848 1472 1880 1504
rect 1920 1472 1952 1504
rect 48 1400 80 1432
rect 120 1400 152 1432
rect 192 1400 224 1432
rect 264 1400 296 1432
rect 336 1400 368 1432
rect 408 1400 440 1432
rect 480 1400 512 1432
rect 552 1400 584 1432
rect 624 1400 656 1432
rect 696 1400 728 1432
rect 768 1400 800 1432
rect 840 1400 872 1432
rect 912 1400 944 1432
rect 984 1400 1016 1432
rect 1056 1400 1088 1432
rect 1128 1400 1160 1432
rect 1200 1400 1232 1432
rect 1272 1400 1304 1432
rect 1344 1400 1376 1432
rect 1416 1400 1448 1432
rect 1488 1400 1520 1432
rect 1560 1400 1592 1432
rect 1632 1400 1664 1432
rect 1704 1400 1736 1432
rect 1776 1400 1808 1432
rect 1848 1400 1880 1432
rect 1920 1400 1952 1432
rect 48 1328 80 1360
rect 120 1328 152 1360
rect 192 1328 224 1360
rect 264 1328 296 1360
rect 336 1328 368 1360
rect 408 1328 440 1360
rect 480 1328 512 1360
rect 552 1328 584 1360
rect 624 1328 656 1360
rect 696 1328 728 1360
rect 768 1328 800 1360
rect 840 1328 872 1360
rect 912 1328 944 1360
rect 984 1328 1016 1360
rect 1056 1328 1088 1360
rect 1128 1328 1160 1360
rect 1200 1328 1232 1360
rect 1272 1328 1304 1360
rect 1344 1328 1376 1360
rect 1416 1328 1448 1360
rect 1488 1328 1520 1360
rect 1560 1328 1592 1360
rect 1632 1328 1664 1360
rect 1704 1328 1736 1360
rect 1776 1328 1808 1360
rect 1848 1328 1880 1360
rect 1920 1328 1952 1360
rect 48 1256 80 1288
rect 120 1256 152 1288
rect 192 1256 224 1288
rect 264 1256 296 1288
rect 336 1256 368 1288
rect 408 1256 440 1288
rect 480 1256 512 1288
rect 552 1256 584 1288
rect 624 1256 656 1288
rect 696 1256 728 1288
rect 768 1256 800 1288
rect 840 1256 872 1288
rect 912 1256 944 1288
rect 984 1256 1016 1288
rect 1056 1256 1088 1288
rect 1128 1256 1160 1288
rect 1200 1256 1232 1288
rect 1272 1256 1304 1288
rect 1344 1256 1376 1288
rect 1416 1256 1448 1288
rect 1488 1256 1520 1288
rect 1560 1256 1592 1288
rect 1632 1256 1664 1288
rect 1704 1256 1736 1288
rect 1776 1256 1808 1288
rect 1848 1256 1880 1288
rect 1920 1256 1952 1288
rect 0 33416 2000 33430
rect 0 33384 120 33416
rect 152 33384 192 33416
rect 224 33384 264 33416
rect 296 33384 336 33416
rect 368 33384 408 33416
rect 440 33384 480 33416
rect 512 33384 552 33416
rect 584 33384 624 33416
rect 656 33384 696 33416
rect 728 33384 768 33416
rect 800 33384 840 33416
rect 872 33384 912 33416
rect 944 33384 984 33416
rect 1016 33384 1056 33416
rect 1088 33384 1128 33416
rect 1160 33384 1200 33416
rect 1232 33384 1272 33416
rect 1304 33384 1344 33416
rect 1376 33384 1416 33416
rect 1448 33384 1488 33416
rect 1520 33384 1560 33416
rect 1592 33384 1632 33416
rect 1664 33384 1704 33416
rect 1736 33384 1776 33416
rect 1808 33384 1848 33416
rect 1880 33384 2000 33416
rect 0 33370 2000 33384
rect 0 29716 2000 29730
rect 0 29684 120 29716
rect 152 29684 192 29716
rect 224 29684 264 29716
rect 296 29684 336 29716
rect 368 29684 408 29716
rect 440 29684 480 29716
rect 512 29684 552 29716
rect 584 29684 624 29716
rect 656 29684 696 29716
rect 728 29684 768 29716
rect 800 29684 840 29716
rect 872 29684 912 29716
rect 944 29684 984 29716
rect 1016 29684 1056 29716
rect 1088 29684 1128 29716
rect 1160 29684 1200 29716
rect 1232 29684 1272 29716
rect 1304 29684 1344 29716
rect 1376 29684 1416 29716
rect 1448 29684 1488 29716
rect 1520 29684 1560 29716
rect 1592 29684 1632 29716
rect 1664 29684 1704 29716
rect 1736 29684 1776 29716
rect 1808 29684 1848 29716
rect 1880 29684 2000 29716
rect 0 29670 2000 29684
rect 0 12144 2000 12200
rect 0 12112 48 12144
rect 80 12112 120 12144
rect 152 12112 192 12144
rect 224 12112 264 12144
rect 296 12112 336 12144
rect 368 12112 408 12144
rect 440 12112 480 12144
rect 512 12112 552 12144
rect 584 12112 624 12144
rect 656 12112 696 12144
rect 728 12112 768 12144
rect 800 12112 840 12144
rect 872 12112 912 12144
rect 944 12112 984 12144
rect 1016 12112 1056 12144
rect 1088 12112 1128 12144
rect 1160 12112 1200 12144
rect 1232 12112 1272 12144
rect 1304 12112 1344 12144
rect 1376 12112 1416 12144
rect 1448 12112 1488 12144
rect 1520 12112 1560 12144
rect 1592 12112 1632 12144
rect 1664 12112 1704 12144
rect 1736 12112 1776 12144
rect 1808 12112 1848 12144
rect 1880 12112 1920 12144
rect 1952 12112 2000 12144
rect 0 12072 2000 12112
rect 0 12040 48 12072
rect 80 12040 120 12072
rect 152 12040 192 12072
rect 224 12040 264 12072
rect 296 12040 336 12072
rect 368 12040 408 12072
rect 440 12040 480 12072
rect 512 12040 552 12072
rect 584 12040 624 12072
rect 656 12040 696 12072
rect 728 12040 768 12072
rect 800 12040 840 12072
rect 872 12040 912 12072
rect 944 12040 984 12072
rect 1016 12040 1056 12072
rect 1088 12040 1128 12072
rect 1160 12040 1200 12072
rect 1232 12040 1272 12072
rect 1304 12040 1344 12072
rect 1376 12040 1416 12072
rect 1448 12040 1488 12072
rect 1520 12040 1560 12072
rect 1592 12040 1632 12072
rect 1664 12040 1704 12072
rect 1736 12040 1776 12072
rect 1808 12040 1848 12072
rect 1880 12040 1920 12072
rect 1952 12040 2000 12072
rect 0 12000 2000 12040
rect 0 11968 48 12000
rect 80 11968 120 12000
rect 152 11968 192 12000
rect 224 11968 264 12000
rect 296 11968 336 12000
rect 368 11968 408 12000
rect 440 11968 480 12000
rect 512 11968 552 12000
rect 584 11968 624 12000
rect 656 11968 696 12000
rect 728 11968 768 12000
rect 800 11968 840 12000
rect 872 11968 912 12000
rect 944 11968 984 12000
rect 1016 11968 1056 12000
rect 1088 11968 1128 12000
rect 1160 11968 1200 12000
rect 1232 11968 1272 12000
rect 1304 11968 1344 12000
rect 1376 11968 1416 12000
rect 1448 11968 1488 12000
rect 1520 11968 1560 12000
rect 1592 11968 1632 12000
rect 1664 11968 1704 12000
rect 1736 11968 1776 12000
rect 1808 11968 1848 12000
rect 1880 11968 1920 12000
rect 1952 11968 2000 12000
rect 0 11928 2000 11968
rect 0 11896 48 11928
rect 80 11896 120 11928
rect 152 11896 192 11928
rect 224 11896 264 11928
rect 296 11896 336 11928
rect 368 11896 408 11928
rect 440 11896 480 11928
rect 512 11896 552 11928
rect 584 11896 624 11928
rect 656 11896 696 11928
rect 728 11896 768 11928
rect 800 11896 840 11928
rect 872 11896 912 11928
rect 944 11896 984 11928
rect 1016 11896 1056 11928
rect 1088 11896 1128 11928
rect 1160 11896 1200 11928
rect 1232 11896 1272 11928
rect 1304 11896 1344 11928
rect 1376 11896 1416 11928
rect 1448 11896 1488 11928
rect 1520 11896 1560 11928
rect 1592 11896 1632 11928
rect 1664 11896 1704 11928
rect 1736 11896 1776 11928
rect 1808 11896 1848 11928
rect 1880 11896 1920 11928
rect 1952 11896 2000 11928
rect 0 11856 2000 11896
rect 0 11824 48 11856
rect 80 11824 120 11856
rect 152 11824 192 11856
rect 224 11824 264 11856
rect 296 11824 336 11856
rect 368 11824 408 11856
rect 440 11824 480 11856
rect 512 11824 552 11856
rect 584 11824 624 11856
rect 656 11824 696 11856
rect 728 11824 768 11856
rect 800 11824 840 11856
rect 872 11824 912 11856
rect 944 11824 984 11856
rect 1016 11824 1056 11856
rect 1088 11824 1128 11856
rect 1160 11824 1200 11856
rect 1232 11824 1272 11856
rect 1304 11824 1344 11856
rect 1376 11824 1416 11856
rect 1448 11824 1488 11856
rect 1520 11824 1560 11856
rect 1592 11824 1632 11856
rect 1664 11824 1704 11856
rect 1736 11824 1776 11856
rect 1808 11824 1848 11856
rect 1880 11824 1920 11856
rect 1952 11824 2000 11856
rect 0 11784 2000 11824
rect 0 11752 48 11784
rect 80 11752 120 11784
rect 152 11752 192 11784
rect 224 11752 264 11784
rect 296 11752 336 11784
rect 368 11752 408 11784
rect 440 11752 480 11784
rect 512 11752 552 11784
rect 584 11752 624 11784
rect 656 11752 696 11784
rect 728 11752 768 11784
rect 800 11752 840 11784
rect 872 11752 912 11784
rect 944 11752 984 11784
rect 1016 11752 1056 11784
rect 1088 11752 1128 11784
rect 1160 11752 1200 11784
rect 1232 11752 1272 11784
rect 1304 11752 1344 11784
rect 1376 11752 1416 11784
rect 1448 11752 1488 11784
rect 1520 11752 1560 11784
rect 1592 11752 1632 11784
rect 1664 11752 1704 11784
rect 1736 11752 1776 11784
rect 1808 11752 1848 11784
rect 1880 11752 1920 11784
rect 1952 11752 2000 11784
rect 0 11712 2000 11752
rect 0 11680 48 11712
rect 80 11680 120 11712
rect 152 11680 192 11712
rect 224 11680 264 11712
rect 296 11680 336 11712
rect 368 11680 408 11712
rect 440 11680 480 11712
rect 512 11680 552 11712
rect 584 11680 624 11712
rect 656 11680 696 11712
rect 728 11680 768 11712
rect 800 11680 840 11712
rect 872 11680 912 11712
rect 944 11680 984 11712
rect 1016 11680 1056 11712
rect 1088 11680 1128 11712
rect 1160 11680 1200 11712
rect 1232 11680 1272 11712
rect 1304 11680 1344 11712
rect 1376 11680 1416 11712
rect 1448 11680 1488 11712
rect 1520 11680 1560 11712
rect 1592 11680 1632 11712
rect 1664 11680 1704 11712
rect 1736 11680 1776 11712
rect 1808 11680 1848 11712
rect 1880 11680 1920 11712
rect 1952 11680 2000 11712
rect 0 11640 2000 11680
rect 0 11608 48 11640
rect 80 11608 120 11640
rect 152 11608 192 11640
rect 224 11608 264 11640
rect 296 11608 336 11640
rect 368 11608 408 11640
rect 440 11608 480 11640
rect 512 11608 552 11640
rect 584 11608 624 11640
rect 656 11608 696 11640
rect 728 11608 768 11640
rect 800 11608 840 11640
rect 872 11608 912 11640
rect 944 11608 984 11640
rect 1016 11608 1056 11640
rect 1088 11608 1128 11640
rect 1160 11608 1200 11640
rect 1232 11608 1272 11640
rect 1304 11608 1344 11640
rect 1376 11608 1416 11640
rect 1448 11608 1488 11640
rect 1520 11608 1560 11640
rect 1592 11608 1632 11640
rect 1664 11608 1704 11640
rect 1736 11608 1776 11640
rect 1808 11608 1848 11640
rect 1880 11608 1920 11640
rect 1952 11608 2000 11640
rect 0 11568 2000 11608
rect 0 11536 48 11568
rect 80 11536 120 11568
rect 152 11536 192 11568
rect 224 11536 264 11568
rect 296 11536 336 11568
rect 368 11536 408 11568
rect 440 11536 480 11568
rect 512 11536 552 11568
rect 584 11536 624 11568
rect 656 11536 696 11568
rect 728 11536 768 11568
rect 800 11536 840 11568
rect 872 11536 912 11568
rect 944 11536 984 11568
rect 1016 11536 1056 11568
rect 1088 11536 1128 11568
rect 1160 11536 1200 11568
rect 1232 11536 1272 11568
rect 1304 11536 1344 11568
rect 1376 11536 1416 11568
rect 1448 11536 1488 11568
rect 1520 11536 1560 11568
rect 1592 11536 1632 11568
rect 1664 11536 1704 11568
rect 1736 11536 1776 11568
rect 1808 11536 1848 11568
rect 1880 11536 1920 11568
rect 1952 11536 2000 11568
rect 0 11496 2000 11536
rect 0 11464 48 11496
rect 80 11464 120 11496
rect 152 11464 192 11496
rect 224 11464 264 11496
rect 296 11464 336 11496
rect 368 11464 408 11496
rect 440 11464 480 11496
rect 512 11464 552 11496
rect 584 11464 624 11496
rect 656 11464 696 11496
rect 728 11464 768 11496
rect 800 11464 840 11496
rect 872 11464 912 11496
rect 944 11464 984 11496
rect 1016 11464 1056 11496
rect 1088 11464 1128 11496
rect 1160 11464 1200 11496
rect 1232 11464 1272 11496
rect 1304 11464 1344 11496
rect 1376 11464 1416 11496
rect 1448 11464 1488 11496
rect 1520 11464 1560 11496
rect 1592 11464 1632 11496
rect 1664 11464 1704 11496
rect 1736 11464 1776 11496
rect 1808 11464 1848 11496
rect 1880 11464 1920 11496
rect 1952 11464 2000 11496
rect 0 11424 2000 11464
rect 0 11392 48 11424
rect 80 11392 120 11424
rect 152 11392 192 11424
rect 224 11392 264 11424
rect 296 11392 336 11424
rect 368 11392 408 11424
rect 440 11392 480 11424
rect 512 11392 552 11424
rect 584 11392 624 11424
rect 656 11392 696 11424
rect 728 11392 768 11424
rect 800 11392 840 11424
rect 872 11392 912 11424
rect 944 11392 984 11424
rect 1016 11392 1056 11424
rect 1088 11392 1128 11424
rect 1160 11392 1200 11424
rect 1232 11392 1272 11424
rect 1304 11392 1344 11424
rect 1376 11392 1416 11424
rect 1448 11392 1488 11424
rect 1520 11392 1560 11424
rect 1592 11392 1632 11424
rect 1664 11392 1704 11424
rect 1736 11392 1776 11424
rect 1808 11392 1848 11424
rect 1880 11392 1920 11424
rect 1952 11392 2000 11424
rect 0 11352 2000 11392
rect 0 11320 48 11352
rect 80 11320 120 11352
rect 152 11320 192 11352
rect 224 11320 264 11352
rect 296 11320 336 11352
rect 368 11320 408 11352
rect 440 11320 480 11352
rect 512 11320 552 11352
rect 584 11320 624 11352
rect 656 11320 696 11352
rect 728 11320 768 11352
rect 800 11320 840 11352
rect 872 11320 912 11352
rect 944 11320 984 11352
rect 1016 11320 1056 11352
rect 1088 11320 1128 11352
rect 1160 11320 1200 11352
rect 1232 11320 1272 11352
rect 1304 11320 1344 11352
rect 1376 11320 1416 11352
rect 1448 11320 1488 11352
rect 1520 11320 1560 11352
rect 1592 11320 1632 11352
rect 1664 11320 1704 11352
rect 1736 11320 1776 11352
rect 1808 11320 1848 11352
rect 1880 11320 1920 11352
rect 1952 11320 2000 11352
rect 0 11280 2000 11320
rect 0 11248 48 11280
rect 80 11248 120 11280
rect 152 11248 192 11280
rect 224 11248 264 11280
rect 296 11248 336 11280
rect 368 11248 408 11280
rect 440 11248 480 11280
rect 512 11248 552 11280
rect 584 11248 624 11280
rect 656 11248 696 11280
rect 728 11248 768 11280
rect 800 11248 840 11280
rect 872 11248 912 11280
rect 944 11248 984 11280
rect 1016 11248 1056 11280
rect 1088 11248 1128 11280
rect 1160 11248 1200 11280
rect 1232 11248 1272 11280
rect 1304 11248 1344 11280
rect 1376 11248 1416 11280
rect 1448 11248 1488 11280
rect 1520 11248 1560 11280
rect 1592 11248 1632 11280
rect 1664 11248 1704 11280
rect 1736 11248 1776 11280
rect 1808 11248 1848 11280
rect 1880 11248 1920 11280
rect 1952 11248 2000 11280
rect 0 11208 2000 11248
rect 0 11176 48 11208
rect 80 11176 120 11208
rect 152 11176 192 11208
rect 224 11176 264 11208
rect 296 11176 336 11208
rect 368 11176 408 11208
rect 440 11176 480 11208
rect 512 11176 552 11208
rect 584 11176 624 11208
rect 656 11176 696 11208
rect 728 11176 768 11208
rect 800 11176 840 11208
rect 872 11176 912 11208
rect 944 11176 984 11208
rect 1016 11176 1056 11208
rect 1088 11176 1128 11208
rect 1160 11176 1200 11208
rect 1232 11176 1272 11208
rect 1304 11176 1344 11208
rect 1376 11176 1416 11208
rect 1448 11176 1488 11208
rect 1520 11176 1560 11208
rect 1592 11176 1632 11208
rect 1664 11176 1704 11208
rect 1736 11176 1776 11208
rect 1808 11176 1848 11208
rect 1880 11176 1920 11208
rect 1952 11176 2000 11208
rect 0 11136 2000 11176
rect 0 11104 48 11136
rect 80 11104 120 11136
rect 152 11104 192 11136
rect 224 11104 264 11136
rect 296 11104 336 11136
rect 368 11104 408 11136
rect 440 11104 480 11136
rect 512 11104 552 11136
rect 584 11104 624 11136
rect 656 11104 696 11136
rect 728 11104 768 11136
rect 800 11104 840 11136
rect 872 11104 912 11136
rect 944 11104 984 11136
rect 1016 11104 1056 11136
rect 1088 11104 1128 11136
rect 1160 11104 1200 11136
rect 1232 11104 1272 11136
rect 1304 11104 1344 11136
rect 1376 11104 1416 11136
rect 1448 11104 1488 11136
rect 1520 11104 1560 11136
rect 1592 11104 1632 11136
rect 1664 11104 1704 11136
rect 1736 11104 1776 11136
rect 1808 11104 1848 11136
rect 1880 11104 1920 11136
rect 1952 11104 2000 11136
rect 0 11064 2000 11104
rect 0 11032 48 11064
rect 80 11032 120 11064
rect 152 11032 192 11064
rect 224 11032 264 11064
rect 296 11032 336 11064
rect 368 11032 408 11064
rect 440 11032 480 11064
rect 512 11032 552 11064
rect 584 11032 624 11064
rect 656 11032 696 11064
rect 728 11032 768 11064
rect 800 11032 840 11064
rect 872 11032 912 11064
rect 944 11032 984 11064
rect 1016 11032 1056 11064
rect 1088 11032 1128 11064
rect 1160 11032 1200 11064
rect 1232 11032 1272 11064
rect 1304 11032 1344 11064
rect 1376 11032 1416 11064
rect 1448 11032 1488 11064
rect 1520 11032 1560 11064
rect 1592 11032 1632 11064
rect 1664 11032 1704 11064
rect 1736 11032 1776 11064
rect 1808 11032 1848 11064
rect 1880 11032 1920 11064
rect 1952 11032 2000 11064
rect 0 10992 2000 11032
rect 0 10960 48 10992
rect 80 10960 120 10992
rect 152 10960 192 10992
rect 224 10960 264 10992
rect 296 10960 336 10992
rect 368 10960 408 10992
rect 440 10960 480 10992
rect 512 10960 552 10992
rect 584 10960 624 10992
rect 656 10960 696 10992
rect 728 10960 768 10992
rect 800 10960 840 10992
rect 872 10960 912 10992
rect 944 10960 984 10992
rect 1016 10960 1056 10992
rect 1088 10960 1128 10992
rect 1160 10960 1200 10992
rect 1232 10960 1272 10992
rect 1304 10960 1344 10992
rect 1376 10960 1416 10992
rect 1448 10960 1488 10992
rect 1520 10960 1560 10992
rect 1592 10960 1632 10992
rect 1664 10960 1704 10992
rect 1736 10960 1776 10992
rect 1808 10960 1848 10992
rect 1880 10960 1920 10992
rect 1952 10960 2000 10992
rect 0 10920 2000 10960
rect 0 10888 48 10920
rect 80 10888 120 10920
rect 152 10888 192 10920
rect 224 10888 264 10920
rect 296 10888 336 10920
rect 368 10888 408 10920
rect 440 10888 480 10920
rect 512 10888 552 10920
rect 584 10888 624 10920
rect 656 10888 696 10920
rect 728 10888 768 10920
rect 800 10888 840 10920
rect 872 10888 912 10920
rect 944 10888 984 10920
rect 1016 10888 1056 10920
rect 1088 10888 1128 10920
rect 1160 10888 1200 10920
rect 1232 10888 1272 10920
rect 1304 10888 1344 10920
rect 1376 10888 1416 10920
rect 1448 10888 1488 10920
rect 1520 10888 1560 10920
rect 1592 10888 1632 10920
rect 1664 10888 1704 10920
rect 1736 10888 1776 10920
rect 1808 10888 1848 10920
rect 1880 10888 1920 10920
rect 1952 10888 2000 10920
rect 0 10848 2000 10888
rect 0 10816 48 10848
rect 80 10816 120 10848
rect 152 10816 192 10848
rect 224 10816 264 10848
rect 296 10816 336 10848
rect 368 10816 408 10848
rect 440 10816 480 10848
rect 512 10816 552 10848
rect 584 10816 624 10848
rect 656 10816 696 10848
rect 728 10816 768 10848
rect 800 10816 840 10848
rect 872 10816 912 10848
rect 944 10816 984 10848
rect 1016 10816 1056 10848
rect 1088 10816 1128 10848
rect 1160 10816 1200 10848
rect 1232 10816 1272 10848
rect 1304 10816 1344 10848
rect 1376 10816 1416 10848
rect 1448 10816 1488 10848
rect 1520 10816 1560 10848
rect 1592 10816 1632 10848
rect 1664 10816 1704 10848
rect 1736 10816 1776 10848
rect 1808 10816 1848 10848
rect 1880 10816 1920 10848
rect 1952 10816 2000 10848
rect 0 10776 2000 10816
rect 0 10744 48 10776
rect 80 10744 120 10776
rect 152 10744 192 10776
rect 224 10744 264 10776
rect 296 10744 336 10776
rect 368 10744 408 10776
rect 440 10744 480 10776
rect 512 10744 552 10776
rect 584 10744 624 10776
rect 656 10744 696 10776
rect 728 10744 768 10776
rect 800 10744 840 10776
rect 872 10744 912 10776
rect 944 10744 984 10776
rect 1016 10744 1056 10776
rect 1088 10744 1128 10776
rect 1160 10744 1200 10776
rect 1232 10744 1272 10776
rect 1304 10744 1344 10776
rect 1376 10744 1416 10776
rect 1448 10744 1488 10776
rect 1520 10744 1560 10776
rect 1592 10744 1632 10776
rect 1664 10744 1704 10776
rect 1736 10744 1776 10776
rect 1808 10744 1848 10776
rect 1880 10744 1920 10776
rect 1952 10744 2000 10776
rect 0 10704 2000 10744
rect 0 10672 48 10704
rect 80 10672 120 10704
rect 152 10672 192 10704
rect 224 10672 264 10704
rect 296 10672 336 10704
rect 368 10672 408 10704
rect 440 10672 480 10704
rect 512 10672 552 10704
rect 584 10672 624 10704
rect 656 10672 696 10704
rect 728 10672 768 10704
rect 800 10672 840 10704
rect 872 10672 912 10704
rect 944 10672 984 10704
rect 1016 10672 1056 10704
rect 1088 10672 1128 10704
rect 1160 10672 1200 10704
rect 1232 10672 1272 10704
rect 1304 10672 1344 10704
rect 1376 10672 1416 10704
rect 1448 10672 1488 10704
rect 1520 10672 1560 10704
rect 1592 10672 1632 10704
rect 1664 10672 1704 10704
rect 1736 10672 1776 10704
rect 1808 10672 1848 10704
rect 1880 10672 1920 10704
rect 1952 10672 2000 10704
rect 0 10632 2000 10672
rect 0 10600 48 10632
rect 80 10600 120 10632
rect 152 10600 192 10632
rect 224 10600 264 10632
rect 296 10600 336 10632
rect 368 10600 408 10632
rect 440 10600 480 10632
rect 512 10600 552 10632
rect 584 10600 624 10632
rect 656 10600 696 10632
rect 728 10600 768 10632
rect 800 10600 840 10632
rect 872 10600 912 10632
rect 944 10600 984 10632
rect 1016 10600 1056 10632
rect 1088 10600 1128 10632
rect 1160 10600 1200 10632
rect 1232 10600 1272 10632
rect 1304 10600 1344 10632
rect 1376 10600 1416 10632
rect 1448 10600 1488 10632
rect 1520 10600 1560 10632
rect 1592 10600 1632 10632
rect 1664 10600 1704 10632
rect 1736 10600 1776 10632
rect 1808 10600 1848 10632
rect 1880 10600 1920 10632
rect 1952 10600 2000 10632
rect 0 10560 2000 10600
rect 0 10528 48 10560
rect 80 10528 120 10560
rect 152 10528 192 10560
rect 224 10528 264 10560
rect 296 10528 336 10560
rect 368 10528 408 10560
rect 440 10528 480 10560
rect 512 10528 552 10560
rect 584 10528 624 10560
rect 656 10528 696 10560
rect 728 10528 768 10560
rect 800 10528 840 10560
rect 872 10528 912 10560
rect 944 10528 984 10560
rect 1016 10528 1056 10560
rect 1088 10528 1128 10560
rect 1160 10528 1200 10560
rect 1232 10528 1272 10560
rect 1304 10528 1344 10560
rect 1376 10528 1416 10560
rect 1448 10528 1488 10560
rect 1520 10528 1560 10560
rect 1592 10528 1632 10560
rect 1664 10528 1704 10560
rect 1736 10528 1776 10560
rect 1808 10528 1848 10560
rect 1880 10528 1920 10560
rect 1952 10528 2000 10560
rect 0 10488 2000 10528
rect 0 10456 48 10488
rect 80 10456 120 10488
rect 152 10456 192 10488
rect 224 10456 264 10488
rect 296 10456 336 10488
rect 368 10456 408 10488
rect 440 10456 480 10488
rect 512 10456 552 10488
rect 584 10456 624 10488
rect 656 10456 696 10488
rect 728 10456 768 10488
rect 800 10456 840 10488
rect 872 10456 912 10488
rect 944 10456 984 10488
rect 1016 10456 1056 10488
rect 1088 10456 1128 10488
rect 1160 10456 1200 10488
rect 1232 10456 1272 10488
rect 1304 10456 1344 10488
rect 1376 10456 1416 10488
rect 1448 10456 1488 10488
rect 1520 10456 1560 10488
rect 1592 10456 1632 10488
rect 1664 10456 1704 10488
rect 1736 10456 1776 10488
rect 1808 10456 1848 10488
rect 1880 10456 1920 10488
rect 1952 10456 2000 10488
rect 0 10416 2000 10456
rect 0 10384 48 10416
rect 80 10384 120 10416
rect 152 10384 192 10416
rect 224 10384 264 10416
rect 296 10384 336 10416
rect 368 10384 408 10416
rect 440 10384 480 10416
rect 512 10384 552 10416
rect 584 10384 624 10416
rect 656 10384 696 10416
rect 728 10384 768 10416
rect 800 10384 840 10416
rect 872 10384 912 10416
rect 944 10384 984 10416
rect 1016 10384 1056 10416
rect 1088 10384 1128 10416
rect 1160 10384 1200 10416
rect 1232 10384 1272 10416
rect 1304 10384 1344 10416
rect 1376 10384 1416 10416
rect 1448 10384 1488 10416
rect 1520 10384 1560 10416
rect 1592 10384 1632 10416
rect 1664 10384 1704 10416
rect 1736 10384 1776 10416
rect 1808 10384 1848 10416
rect 1880 10384 1920 10416
rect 1952 10384 2000 10416
rect 0 10344 2000 10384
rect 0 10312 48 10344
rect 80 10312 120 10344
rect 152 10312 192 10344
rect 224 10312 264 10344
rect 296 10312 336 10344
rect 368 10312 408 10344
rect 440 10312 480 10344
rect 512 10312 552 10344
rect 584 10312 624 10344
rect 656 10312 696 10344
rect 728 10312 768 10344
rect 800 10312 840 10344
rect 872 10312 912 10344
rect 944 10312 984 10344
rect 1016 10312 1056 10344
rect 1088 10312 1128 10344
rect 1160 10312 1200 10344
rect 1232 10312 1272 10344
rect 1304 10312 1344 10344
rect 1376 10312 1416 10344
rect 1448 10312 1488 10344
rect 1520 10312 1560 10344
rect 1592 10312 1632 10344
rect 1664 10312 1704 10344
rect 1736 10312 1776 10344
rect 1808 10312 1848 10344
rect 1880 10312 1920 10344
rect 1952 10312 2000 10344
rect 0 10272 2000 10312
rect 0 10240 48 10272
rect 80 10240 120 10272
rect 152 10240 192 10272
rect 224 10240 264 10272
rect 296 10240 336 10272
rect 368 10240 408 10272
rect 440 10240 480 10272
rect 512 10240 552 10272
rect 584 10240 624 10272
rect 656 10240 696 10272
rect 728 10240 768 10272
rect 800 10240 840 10272
rect 872 10240 912 10272
rect 944 10240 984 10272
rect 1016 10240 1056 10272
rect 1088 10240 1128 10272
rect 1160 10240 1200 10272
rect 1232 10240 1272 10272
rect 1304 10240 1344 10272
rect 1376 10240 1416 10272
rect 1448 10240 1488 10272
rect 1520 10240 1560 10272
rect 1592 10240 1632 10272
rect 1664 10240 1704 10272
rect 1736 10240 1776 10272
rect 1808 10240 1848 10272
rect 1880 10240 1920 10272
rect 1952 10240 2000 10272
rect 0 10200 2000 10240
rect 0 10168 48 10200
rect 80 10168 120 10200
rect 152 10168 192 10200
rect 224 10168 264 10200
rect 296 10168 336 10200
rect 368 10168 408 10200
rect 440 10168 480 10200
rect 512 10168 552 10200
rect 584 10168 624 10200
rect 656 10168 696 10200
rect 728 10168 768 10200
rect 800 10168 840 10200
rect 872 10168 912 10200
rect 944 10168 984 10200
rect 1016 10168 1056 10200
rect 1088 10168 1128 10200
rect 1160 10168 1200 10200
rect 1232 10168 1272 10200
rect 1304 10168 1344 10200
rect 1376 10168 1416 10200
rect 1448 10168 1488 10200
rect 1520 10168 1560 10200
rect 1592 10168 1632 10200
rect 1664 10168 1704 10200
rect 1736 10168 1776 10200
rect 1808 10168 1848 10200
rect 1880 10168 1920 10200
rect 1952 10168 2000 10200
rect 0 10128 2000 10168
rect 0 10096 48 10128
rect 80 10096 120 10128
rect 152 10096 192 10128
rect 224 10096 264 10128
rect 296 10096 336 10128
rect 368 10096 408 10128
rect 440 10096 480 10128
rect 512 10096 552 10128
rect 584 10096 624 10128
rect 656 10096 696 10128
rect 728 10096 768 10128
rect 800 10096 840 10128
rect 872 10096 912 10128
rect 944 10096 984 10128
rect 1016 10096 1056 10128
rect 1088 10096 1128 10128
rect 1160 10096 1200 10128
rect 1232 10096 1272 10128
rect 1304 10096 1344 10128
rect 1376 10096 1416 10128
rect 1448 10096 1488 10128
rect 1520 10096 1560 10128
rect 1592 10096 1632 10128
rect 1664 10096 1704 10128
rect 1736 10096 1776 10128
rect 1808 10096 1848 10128
rect 1880 10096 1920 10128
rect 1952 10096 2000 10128
rect 0 10056 2000 10096
rect 0 10024 48 10056
rect 80 10024 120 10056
rect 152 10024 192 10056
rect 224 10024 264 10056
rect 296 10024 336 10056
rect 368 10024 408 10056
rect 440 10024 480 10056
rect 512 10024 552 10056
rect 584 10024 624 10056
rect 656 10024 696 10056
rect 728 10024 768 10056
rect 800 10024 840 10056
rect 872 10024 912 10056
rect 944 10024 984 10056
rect 1016 10024 1056 10056
rect 1088 10024 1128 10056
rect 1160 10024 1200 10056
rect 1232 10024 1272 10056
rect 1304 10024 1344 10056
rect 1376 10024 1416 10056
rect 1448 10024 1488 10056
rect 1520 10024 1560 10056
rect 1592 10024 1632 10056
rect 1664 10024 1704 10056
rect 1736 10024 1776 10056
rect 1808 10024 1848 10056
rect 1880 10024 1920 10056
rect 1952 10024 2000 10056
rect 0 9984 2000 10024
rect 0 9952 48 9984
rect 80 9952 120 9984
rect 152 9952 192 9984
rect 224 9952 264 9984
rect 296 9952 336 9984
rect 368 9952 408 9984
rect 440 9952 480 9984
rect 512 9952 552 9984
rect 584 9952 624 9984
rect 656 9952 696 9984
rect 728 9952 768 9984
rect 800 9952 840 9984
rect 872 9952 912 9984
rect 944 9952 984 9984
rect 1016 9952 1056 9984
rect 1088 9952 1128 9984
rect 1160 9952 1200 9984
rect 1232 9952 1272 9984
rect 1304 9952 1344 9984
rect 1376 9952 1416 9984
rect 1448 9952 1488 9984
rect 1520 9952 1560 9984
rect 1592 9952 1632 9984
rect 1664 9952 1704 9984
rect 1736 9952 1776 9984
rect 1808 9952 1848 9984
rect 1880 9952 1920 9984
rect 1952 9952 2000 9984
rect 0 9912 2000 9952
rect 0 9880 48 9912
rect 80 9880 120 9912
rect 152 9880 192 9912
rect 224 9880 264 9912
rect 296 9880 336 9912
rect 368 9880 408 9912
rect 440 9880 480 9912
rect 512 9880 552 9912
rect 584 9880 624 9912
rect 656 9880 696 9912
rect 728 9880 768 9912
rect 800 9880 840 9912
rect 872 9880 912 9912
rect 944 9880 984 9912
rect 1016 9880 1056 9912
rect 1088 9880 1128 9912
rect 1160 9880 1200 9912
rect 1232 9880 1272 9912
rect 1304 9880 1344 9912
rect 1376 9880 1416 9912
rect 1448 9880 1488 9912
rect 1520 9880 1560 9912
rect 1592 9880 1632 9912
rect 1664 9880 1704 9912
rect 1736 9880 1776 9912
rect 1808 9880 1848 9912
rect 1880 9880 1920 9912
rect 1952 9880 2000 9912
rect 0 9840 2000 9880
rect 0 9808 48 9840
rect 80 9808 120 9840
rect 152 9808 192 9840
rect 224 9808 264 9840
rect 296 9808 336 9840
rect 368 9808 408 9840
rect 440 9808 480 9840
rect 512 9808 552 9840
rect 584 9808 624 9840
rect 656 9808 696 9840
rect 728 9808 768 9840
rect 800 9808 840 9840
rect 872 9808 912 9840
rect 944 9808 984 9840
rect 1016 9808 1056 9840
rect 1088 9808 1128 9840
rect 1160 9808 1200 9840
rect 1232 9808 1272 9840
rect 1304 9808 1344 9840
rect 1376 9808 1416 9840
rect 1448 9808 1488 9840
rect 1520 9808 1560 9840
rect 1592 9808 1632 9840
rect 1664 9808 1704 9840
rect 1736 9808 1776 9840
rect 1808 9808 1848 9840
rect 1880 9808 1920 9840
rect 1952 9808 2000 9840
rect 0 9768 2000 9808
rect 0 9736 48 9768
rect 80 9736 120 9768
rect 152 9736 192 9768
rect 224 9736 264 9768
rect 296 9736 336 9768
rect 368 9736 408 9768
rect 440 9736 480 9768
rect 512 9736 552 9768
rect 584 9736 624 9768
rect 656 9736 696 9768
rect 728 9736 768 9768
rect 800 9736 840 9768
rect 872 9736 912 9768
rect 944 9736 984 9768
rect 1016 9736 1056 9768
rect 1088 9736 1128 9768
rect 1160 9736 1200 9768
rect 1232 9736 1272 9768
rect 1304 9736 1344 9768
rect 1376 9736 1416 9768
rect 1448 9736 1488 9768
rect 1520 9736 1560 9768
rect 1592 9736 1632 9768
rect 1664 9736 1704 9768
rect 1736 9736 1776 9768
rect 1808 9736 1848 9768
rect 1880 9736 1920 9768
rect 1952 9736 2000 9768
rect 0 9696 2000 9736
rect 0 9664 48 9696
rect 80 9664 120 9696
rect 152 9664 192 9696
rect 224 9664 264 9696
rect 296 9664 336 9696
rect 368 9664 408 9696
rect 440 9664 480 9696
rect 512 9664 552 9696
rect 584 9664 624 9696
rect 656 9664 696 9696
rect 728 9664 768 9696
rect 800 9664 840 9696
rect 872 9664 912 9696
rect 944 9664 984 9696
rect 1016 9664 1056 9696
rect 1088 9664 1128 9696
rect 1160 9664 1200 9696
rect 1232 9664 1272 9696
rect 1304 9664 1344 9696
rect 1376 9664 1416 9696
rect 1448 9664 1488 9696
rect 1520 9664 1560 9696
rect 1592 9664 1632 9696
rect 1664 9664 1704 9696
rect 1736 9664 1776 9696
rect 1808 9664 1848 9696
rect 1880 9664 1920 9696
rect 1952 9664 2000 9696
rect 0 9624 2000 9664
rect 0 9592 48 9624
rect 80 9592 120 9624
rect 152 9592 192 9624
rect 224 9592 264 9624
rect 296 9592 336 9624
rect 368 9592 408 9624
rect 440 9592 480 9624
rect 512 9592 552 9624
rect 584 9592 624 9624
rect 656 9592 696 9624
rect 728 9592 768 9624
rect 800 9592 840 9624
rect 872 9592 912 9624
rect 944 9592 984 9624
rect 1016 9592 1056 9624
rect 1088 9592 1128 9624
rect 1160 9592 1200 9624
rect 1232 9592 1272 9624
rect 1304 9592 1344 9624
rect 1376 9592 1416 9624
rect 1448 9592 1488 9624
rect 1520 9592 1560 9624
rect 1592 9592 1632 9624
rect 1664 9592 1704 9624
rect 1736 9592 1776 9624
rect 1808 9592 1848 9624
rect 1880 9592 1920 9624
rect 1952 9592 2000 9624
rect 0 9552 2000 9592
rect 0 9520 48 9552
rect 80 9520 120 9552
rect 152 9520 192 9552
rect 224 9520 264 9552
rect 296 9520 336 9552
rect 368 9520 408 9552
rect 440 9520 480 9552
rect 512 9520 552 9552
rect 584 9520 624 9552
rect 656 9520 696 9552
rect 728 9520 768 9552
rect 800 9520 840 9552
rect 872 9520 912 9552
rect 944 9520 984 9552
rect 1016 9520 1056 9552
rect 1088 9520 1128 9552
rect 1160 9520 1200 9552
rect 1232 9520 1272 9552
rect 1304 9520 1344 9552
rect 1376 9520 1416 9552
rect 1448 9520 1488 9552
rect 1520 9520 1560 9552
rect 1592 9520 1632 9552
rect 1664 9520 1704 9552
rect 1736 9520 1776 9552
rect 1808 9520 1848 9552
rect 1880 9520 1920 9552
rect 1952 9520 2000 9552
rect 0 9480 2000 9520
rect 0 9448 48 9480
rect 80 9448 120 9480
rect 152 9448 192 9480
rect 224 9448 264 9480
rect 296 9448 336 9480
rect 368 9448 408 9480
rect 440 9448 480 9480
rect 512 9448 552 9480
rect 584 9448 624 9480
rect 656 9448 696 9480
rect 728 9448 768 9480
rect 800 9448 840 9480
rect 872 9448 912 9480
rect 944 9448 984 9480
rect 1016 9448 1056 9480
rect 1088 9448 1128 9480
rect 1160 9448 1200 9480
rect 1232 9448 1272 9480
rect 1304 9448 1344 9480
rect 1376 9448 1416 9480
rect 1448 9448 1488 9480
rect 1520 9448 1560 9480
rect 1592 9448 1632 9480
rect 1664 9448 1704 9480
rect 1736 9448 1776 9480
rect 1808 9448 1848 9480
rect 1880 9448 1920 9480
rect 1952 9448 2000 9480
rect 0 9408 2000 9448
rect 0 9376 48 9408
rect 80 9376 120 9408
rect 152 9376 192 9408
rect 224 9376 264 9408
rect 296 9376 336 9408
rect 368 9376 408 9408
rect 440 9376 480 9408
rect 512 9376 552 9408
rect 584 9376 624 9408
rect 656 9376 696 9408
rect 728 9376 768 9408
rect 800 9376 840 9408
rect 872 9376 912 9408
rect 944 9376 984 9408
rect 1016 9376 1056 9408
rect 1088 9376 1128 9408
rect 1160 9376 1200 9408
rect 1232 9376 1272 9408
rect 1304 9376 1344 9408
rect 1376 9376 1416 9408
rect 1448 9376 1488 9408
rect 1520 9376 1560 9408
rect 1592 9376 1632 9408
rect 1664 9376 1704 9408
rect 1736 9376 1776 9408
rect 1808 9376 1848 9408
rect 1880 9376 1920 9408
rect 1952 9376 2000 9408
rect 0 9336 2000 9376
rect 0 9304 48 9336
rect 80 9304 120 9336
rect 152 9304 192 9336
rect 224 9304 264 9336
rect 296 9304 336 9336
rect 368 9304 408 9336
rect 440 9304 480 9336
rect 512 9304 552 9336
rect 584 9304 624 9336
rect 656 9304 696 9336
rect 728 9304 768 9336
rect 800 9304 840 9336
rect 872 9304 912 9336
rect 944 9304 984 9336
rect 1016 9304 1056 9336
rect 1088 9304 1128 9336
rect 1160 9304 1200 9336
rect 1232 9304 1272 9336
rect 1304 9304 1344 9336
rect 1376 9304 1416 9336
rect 1448 9304 1488 9336
rect 1520 9304 1560 9336
rect 1592 9304 1632 9336
rect 1664 9304 1704 9336
rect 1736 9304 1776 9336
rect 1808 9304 1848 9336
rect 1880 9304 1920 9336
rect 1952 9304 2000 9336
rect 0 9264 2000 9304
rect 0 9232 48 9264
rect 80 9232 120 9264
rect 152 9232 192 9264
rect 224 9232 264 9264
rect 296 9232 336 9264
rect 368 9232 408 9264
rect 440 9232 480 9264
rect 512 9232 552 9264
rect 584 9232 624 9264
rect 656 9232 696 9264
rect 728 9232 768 9264
rect 800 9232 840 9264
rect 872 9232 912 9264
rect 944 9232 984 9264
rect 1016 9232 1056 9264
rect 1088 9232 1128 9264
rect 1160 9232 1200 9264
rect 1232 9232 1272 9264
rect 1304 9232 1344 9264
rect 1376 9232 1416 9264
rect 1448 9232 1488 9264
rect 1520 9232 1560 9264
rect 1592 9232 1632 9264
rect 1664 9232 1704 9264
rect 1736 9232 1776 9264
rect 1808 9232 1848 9264
rect 1880 9232 1920 9264
rect 1952 9232 2000 9264
rect 0 9192 2000 9232
rect 0 9160 48 9192
rect 80 9160 120 9192
rect 152 9160 192 9192
rect 224 9160 264 9192
rect 296 9160 336 9192
rect 368 9160 408 9192
rect 440 9160 480 9192
rect 512 9160 552 9192
rect 584 9160 624 9192
rect 656 9160 696 9192
rect 728 9160 768 9192
rect 800 9160 840 9192
rect 872 9160 912 9192
rect 944 9160 984 9192
rect 1016 9160 1056 9192
rect 1088 9160 1128 9192
rect 1160 9160 1200 9192
rect 1232 9160 1272 9192
rect 1304 9160 1344 9192
rect 1376 9160 1416 9192
rect 1448 9160 1488 9192
rect 1520 9160 1560 9192
rect 1592 9160 1632 9192
rect 1664 9160 1704 9192
rect 1736 9160 1776 9192
rect 1808 9160 1848 9192
rect 1880 9160 1920 9192
rect 1952 9160 2000 9192
rect 0 9120 2000 9160
rect 0 9088 48 9120
rect 80 9088 120 9120
rect 152 9088 192 9120
rect 224 9088 264 9120
rect 296 9088 336 9120
rect 368 9088 408 9120
rect 440 9088 480 9120
rect 512 9088 552 9120
rect 584 9088 624 9120
rect 656 9088 696 9120
rect 728 9088 768 9120
rect 800 9088 840 9120
rect 872 9088 912 9120
rect 944 9088 984 9120
rect 1016 9088 1056 9120
rect 1088 9088 1128 9120
rect 1160 9088 1200 9120
rect 1232 9088 1272 9120
rect 1304 9088 1344 9120
rect 1376 9088 1416 9120
rect 1448 9088 1488 9120
rect 1520 9088 1560 9120
rect 1592 9088 1632 9120
rect 1664 9088 1704 9120
rect 1736 9088 1776 9120
rect 1808 9088 1848 9120
rect 1880 9088 1920 9120
rect 1952 9088 2000 9120
rect 0 9048 2000 9088
rect 0 9016 48 9048
rect 80 9016 120 9048
rect 152 9016 192 9048
rect 224 9016 264 9048
rect 296 9016 336 9048
rect 368 9016 408 9048
rect 440 9016 480 9048
rect 512 9016 552 9048
rect 584 9016 624 9048
rect 656 9016 696 9048
rect 728 9016 768 9048
rect 800 9016 840 9048
rect 872 9016 912 9048
rect 944 9016 984 9048
rect 1016 9016 1056 9048
rect 1088 9016 1128 9048
rect 1160 9016 1200 9048
rect 1232 9016 1272 9048
rect 1304 9016 1344 9048
rect 1376 9016 1416 9048
rect 1448 9016 1488 9048
rect 1520 9016 1560 9048
rect 1592 9016 1632 9048
rect 1664 9016 1704 9048
rect 1736 9016 1776 9048
rect 1808 9016 1848 9048
rect 1880 9016 1920 9048
rect 1952 9016 2000 9048
rect 0 8976 2000 9016
rect 0 8944 48 8976
rect 80 8944 120 8976
rect 152 8944 192 8976
rect 224 8944 264 8976
rect 296 8944 336 8976
rect 368 8944 408 8976
rect 440 8944 480 8976
rect 512 8944 552 8976
rect 584 8944 624 8976
rect 656 8944 696 8976
rect 728 8944 768 8976
rect 800 8944 840 8976
rect 872 8944 912 8976
rect 944 8944 984 8976
rect 1016 8944 1056 8976
rect 1088 8944 1128 8976
rect 1160 8944 1200 8976
rect 1232 8944 1272 8976
rect 1304 8944 1344 8976
rect 1376 8944 1416 8976
rect 1448 8944 1488 8976
rect 1520 8944 1560 8976
rect 1592 8944 1632 8976
rect 1664 8944 1704 8976
rect 1736 8944 1776 8976
rect 1808 8944 1848 8976
rect 1880 8944 1920 8976
rect 1952 8944 2000 8976
rect 0 8904 2000 8944
rect 0 8872 48 8904
rect 80 8872 120 8904
rect 152 8872 192 8904
rect 224 8872 264 8904
rect 296 8872 336 8904
rect 368 8872 408 8904
rect 440 8872 480 8904
rect 512 8872 552 8904
rect 584 8872 624 8904
rect 656 8872 696 8904
rect 728 8872 768 8904
rect 800 8872 840 8904
rect 872 8872 912 8904
rect 944 8872 984 8904
rect 1016 8872 1056 8904
rect 1088 8872 1128 8904
rect 1160 8872 1200 8904
rect 1232 8872 1272 8904
rect 1304 8872 1344 8904
rect 1376 8872 1416 8904
rect 1448 8872 1488 8904
rect 1520 8872 1560 8904
rect 1592 8872 1632 8904
rect 1664 8872 1704 8904
rect 1736 8872 1776 8904
rect 1808 8872 1848 8904
rect 1880 8872 1920 8904
rect 1952 8872 2000 8904
rect 0 8832 2000 8872
rect 0 8800 48 8832
rect 80 8800 120 8832
rect 152 8800 192 8832
rect 224 8800 264 8832
rect 296 8800 336 8832
rect 368 8800 408 8832
rect 440 8800 480 8832
rect 512 8800 552 8832
rect 584 8800 624 8832
rect 656 8800 696 8832
rect 728 8800 768 8832
rect 800 8800 840 8832
rect 872 8800 912 8832
rect 944 8800 984 8832
rect 1016 8800 1056 8832
rect 1088 8800 1128 8832
rect 1160 8800 1200 8832
rect 1232 8800 1272 8832
rect 1304 8800 1344 8832
rect 1376 8800 1416 8832
rect 1448 8800 1488 8832
rect 1520 8800 1560 8832
rect 1592 8800 1632 8832
rect 1664 8800 1704 8832
rect 1736 8800 1776 8832
rect 1808 8800 1848 8832
rect 1880 8800 1920 8832
rect 1952 8800 2000 8832
rect 0 8760 2000 8800
rect 0 8728 48 8760
rect 80 8728 120 8760
rect 152 8728 192 8760
rect 224 8728 264 8760
rect 296 8728 336 8760
rect 368 8728 408 8760
rect 440 8728 480 8760
rect 512 8728 552 8760
rect 584 8728 624 8760
rect 656 8728 696 8760
rect 728 8728 768 8760
rect 800 8728 840 8760
rect 872 8728 912 8760
rect 944 8728 984 8760
rect 1016 8728 1056 8760
rect 1088 8728 1128 8760
rect 1160 8728 1200 8760
rect 1232 8728 1272 8760
rect 1304 8728 1344 8760
rect 1376 8728 1416 8760
rect 1448 8728 1488 8760
rect 1520 8728 1560 8760
rect 1592 8728 1632 8760
rect 1664 8728 1704 8760
rect 1736 8728 1776 8760
rect 1808 8728 1848 8760
rect 1880 8728 1920 8760
rect 1952 8728 2000 8760
rect 0 8688 2000 8728
rect 0 8656 48 8688
rect 80 8656 120 8688
rect 152 8656 192 8688
rect 224 8656 264 8688
rect 296 8656 336 8688
rect 368 8656 408 8688
rect 440 8656 480 8688
rect 512 8656 552 8688
rect 584 8656 624 8688
rect 656 8656 696 8688
rect 728 8656 768 8688
rect 800 8656 840 8688
rect 872 8656 912 8688
rect 944 8656 984 8688
rect 1016 8656 1056 8688
rect 1088 8656 1128 8688
rect 1160 8656 1200 8688
rect 1232 8656 1272 8688
rect 1304 8656 1344 8688
rect 1376 8656 1416 8688
rect 1448 8656 1488 8688
rect 1520 8656 1560 8688
rect 1592 8656 1632 8688
rect 1664 8656 1704 8688
rect 1736 8656 1776 8688
rect 1808 8656 1848 8688
rect 1880 8656 1920 8688
rect 1952 8656 2000 8688
rect 0 8616 2000 8656
rect 0 8584 48 8616
rect 80 8584 120 8616
rect 152 8584 192 8616
rect 224 8584 264 8616
rect 296 8584 336 8616
rect 368 8584 408 8616
rect 440 8584 480 8616
rect 512 8584 552 8616
rect 584 8584 624 8616
rect 656 8584 696 8616
rect 728 8584 768 8616
rect 800 8584 840 8616
rect 872 8584 912 8616
rect 944 8584 984 8616
rect 1016 8584 1056 8616
rect 1088 8584 1128 8616
rect 1160 8584 1200 8616
rect 1232 8584 1272 8616
rect 1304 8584 1344 8616
rect 1376 8584 1416 8616
rect 1448 8584 1488 8616
rect 1520 8584 1560 8616
rect 1592 8584 1632 8616
rect 1664 8584 1704 8616
rect 1736 8584 1776 8616
rect 1808 8584 1848 8616
rect 1880 8584 1920 8616
rect 1952 8584 2000 8616
rect 0 8544 2000 8584
rect 0 8512 48 8544
rect 80 8512 120 8544
rect 152 8512 192 8544
rect 224 8512 264 8544
rect 296 8512 336 8544
rect 368 8512 408 8544
rect 440 8512 480 8544
rect 512 8512 552 8544
rect 584 8512 624 8544
rect 656 8512 696 8544
rect 728 8512 768 8544
rect 800 8512 840 8544
rect 872 8512 912 8544
rect 944 8512 984 8544
rect 1016 8512 1056 8544
rect 1088 8512 1128 8544
rect 1160 8512 1200 8544
rect 1232 8512 1272 8544
rect 1304 8512 1344 8544
rect 1376 8512 1416 8544
rect 1448 8512 1488 8544
rect 1520 8512 1560 8544
rect 1592 8512 1632 8544
rect 1664 8512 1704 8544
rect 1736 8512 1776 8544
rect 1808 8512 1848 8544
rect 1880 8512 1920 8544
rect 1952 8512 2000 8544
rect 0 8472 2000 8512
rect 0 8440 48 8472
rect 80 8440 120 8472
rect 152 8440 192 8472
rect 224 8440 264 8472
rect 296 8440 336 8472
rect 368 8440 408 8472
rect 440 8440 480 8472
rect 512 8440 552 8472
rect 584 8440 624 8472
rect 656 8440 696 8472
rect 728 8440 768 8472
rect 800 8440 840 8472
rect 872 8440 912 8472
rect 944 8440 984 8472
rect 1016 8440 1056 8472
rect 1088 8440 1128 8472
rect 1160 8440 1200 8472
rect 1232 8440 1272 8472
rect 1304 8440 1344 8472
rect 1376 8440 1416 8472
rect 1448 8440 1488 8472
rect 1520 8440 1560 8472
rect 1592 8440 1632 8472
rect 1664 8440 1704 8472
rect 1736 8440 1776 8472
rect 1808 8440 1848 8472
rect 1880 8440 1920 8472
rect 1952 8440 2000 8472
rect 0 8400 2000 8440
rect 0 8368 48 8400
rect 80 8368 120 8400
rect 152 8368 192 8400
rect 224 8368 264 8400
rect 296 8368 336 8400
rect 368 8368 408 8400
rect 440 8368 480 8400
rect 512 8368 552 8400
rect 584 8368 624 8400
rect 656 8368 696 8400
rect 728 8368 768 8400
rect 800 8368 840 8400
rect 872 8368 912 8400
rect 944 8368 984 8400
rect 1016 8368 1056 8400
rect 1088 8368 1128 8400
rect 1160 8368 1200 8400
rect 1232 8368 1272 8400
rect 1304 8368 1344 8400
rect 1376 8368 1416 8400
rect 1448 8368 1488 8400
rect 1520 8368 1560 8400
rect 1592 8368 1632 8400
rect 1664 8368 1704 8400
rect 1736 8368 1776 8400
rect 1808 8368 1848 8400
rect 1880 8368 1920 8400
rect 1952 8368 2000 8400
rect 0 8328 2000 8368
rect 0 8296 48 8328
rect 80 8296 120 8328
rect 152 8296 192 8328
rect 224 8296 264 8328
rect 296 8296 336 8328
rect 368 8296 408 8328
rect 440 8296 480 8328
rect 512 8296 552 8328
rect 584 8296 624 8328
rect 656 8296 696 8328
rect 728 8296 768 8328
rect 800 8296 840 8328
rect 872 8296 912 8328
rect 944 8296 984 8328
rect 1016 8296 1056 8328
rect 1088 8296 1128 8328
rect 1160 8296 1200 8328
rect 1232 8296 1272 8328
rect 1304 8296 1344 8328
rect 1376 8296 1416 8328
rect 1448 8296 1488 8328
rect 1520 8296 1560 8328
rect 1592 8296 1632 8328
rect 1664 8296 1704 8328
rect 1736 8296 1776 8328
rect 1808 8296 1848 8328
rect 1880 8296 1920 8328
rect 1952 8296 2000 8328
rect 0 8256 2000 8296
rect 0 8224 48 8256
rect 80 8224 120 8256
rect 152 8224 192 8256
rect 224 8224 264 8256
rect 296 8224 336 8256
rect 368 8224 408 8256
rect 440 8224 480 8256
rect 512 8224 552 8256
rect 584 8224 624 8256
rect 656 8224 696 8256
rect 728 8224 768 8256
rect 800 8224 840 8256
rect 872 8224 912 8256
rect 944 8224 984 8256
rect 1016 8224 1056 8256
rect 1088 8224 1128 8256
rect 1160 8224 1200 8256
rect 1232 8224 1272 8256
rect 1304 8224 1344 8256
rect 1376 8224 1416 8256
rect 1448 8224 1488 8256
rect 1520 8224 1560 8256
rect 1592 8224 1632 8256
rect 1664 8224 1704 8256
rect 1736 8224 1776 8256
rect 1808 8224 1848 8256
rect 1880 8224 1920 8256
rect 1952 8224 2000 8256
rect 0 8184 2000 8224
rect 0 8152 48 8184
rect 80 8152 120 8184
rect 152 8152 192 8184
rect 224 8152 264 8184
rect 296 8152 336 8184
rect 368 8152 408 8184
rect 440 8152 480 8184
rect 512 8152 552 8184
rect 584 8152 624 8184
rect 656 8152 696 8184
rect 728 8152 768 8184
rect 800 8152 840 8184
rect 872 8152 912 8184
rect 944 8152 984 8184
rect 1016 8152 1056 8184
rect 1088 8152 1128 8184
rect 1160 8152 1200 8184
rect 1232 8152 1272 8184
rect 1304 8152 1344 8184
rect 1376 8152 1416 8184
rect 1448 8152 1488 8184
rect 1520 8152 1560 8184
rect 1592 8152 1632 8184
rect 1664 8152 1704 8184
rect 1736 8152 1776 8184
rect 1808 8152 1848 8184
rect 1880 8152 1920 8184
rect 1952 8152 2000 8184
rect 0 8112 2000 8152
rect 0 8080 48 8112
rect 80 8080 120 8112
rect 152 8080 192 8112
rect 224 8080 264 8112
rect 296 8080 336 8112
rect 368 8080 408 8112
rect 440 8080 480 8112
rect 512 8080 552 8112
rect 584 8080 624 8112
rect 656 8080 696 8112
rect 728 8080 768 8112
rect 800 8080 840 8112
rect 872 8080 912 8112
rect 944 8080 984 8112
rect 1016 8080 1056 8112
rect 1088 8080 1128 8112
rect 1160 8080 1200 8112
rect 1232 8080 1272 8112
rect 1304 8080 1344 8112
rect 1376 8080 1416 8112
rect 1448 8080 1488 8112
rect 1520 8080 1560 8112
rect 1592 8080 1632 8112
rect 1664 8080 1704 8112
rect 1736 8080 1776 8112
rect 1808 8080 1848 8112
rect 1880 8080 1920 8112
rect 1952 8080 2000 8112
rect 0 8040 2000 8080
rect 0 8008 48 8040
rect 80 8008 120 8040
rect 152 8008 192 8040
rect 224 8008 264 8040
rect 296 8008 336 8040
rect 368 8008 408 8040
rect 440 8008 480 8040
rect 512 8008 552 8040
rect 584 8008 624 8040
rect 656 8008 696 8040
rect 728 8008 768 8040
rect 800 8008 840 8040
rect 872 8008 912 8040
rect 944 8008 984 8040
rect 1016 8008 1056 8040
rect 1088 8008 1128 8040
rect 1160 8008 1200 8040
rect 1232 8008 1272 8040
rect 1304 8008 1344 8040
rect 1376 8008 1416 8040
rect 1448 8008 1488 8040
rect 1520 8008 1560 8040
rect 1592 8008 1632 8040
rect 1664 8008 1704 8040
rect 1736 8008 1776 8040
rect 1808 8008 1848 8040
rect 1880 8008 1920 8040
rect 1952 8008 2000 8040
rect 0 7968 2000 8008
rect 0 7936 48 7968
rect 80 7936 120 7968
rect 152 7936 192 7968
rect 224 7936 264 7968
rect 296 7936 336 7968
rect 368 7936 408 7968
rect 440 7936 480 7968
rect 512 7936 552 7968
rect 584 7936 624 7968
rect 656 7936 696 7968
rect 728 7936 768 7968
rect 800 7936 840 7968
rect 872 7936 912 7968
rect 944 7936 984 7968
rect 1016 7936 1056 7968
rect 1088 7936 1128 7968
rect 1160 7936 1200 7968
rect 1232 7936 1272 7968
rect 1304 7936 1344 7968
rect 1376 7936 1416 7968
rect 1448 7936 1488 7968
rect 1520 7936 1560 7968
rect 1592 7936 1632 7968
rect 1664 7936 1704 7968
rect 1736 7936 1776 7968
rect 1808 7936 1848 7968
rect 1880 7936 1920 7968
rect 1952 7936 2000 7968
rect 0 7896 2000 7936
rect 0 7864 48 7896
rect 80 7864 120 7896
rect 152 7864 192 7896
rect 224 7864 264 7896
rect 296 7864 336 7896
rect 368 7864 408 7896
rect 440 7864 480 7896
rect 512 7864 552 7896
rect 584 7864 624 7896
rect 656 7864 696 7896
rect 728 7864 768 7896
rect 800 7864 840 7896
rect 872 7864 912 7896
rect 944 7864 984 7896
rect 1016 7864 1056 7896
rect 1088 7864 1128 7896
rect 1160 7864 1200 7896
rect 1232 7864 1272 7896
rect 1304 7864 1344 7896
rect 1376 7864 1416 7896
rect 1448 7864 1488 7896
rect 1520 7864 1560 7896
rect 1592 7864 1632 7896
rect 1664 7864 1704 7896
rect 1736 7864 1776 7896
rect 1808 7864 1848 7896
rect 1880 7864 1920 7896
rect 1952 7864 2000 7896
rect 0 7824 2000 7864
rect 0 7792 48 7824
rect 80 7792 120 7824
rect 152 7792 192 7824
rect 224 7792 264 7824
rect 296 7792 336 7824
rect 368 7792 408 7824
rect 440 7792 480 7824
rect 512 7792 552 7824
rect 584 7792 624 7824
rect 656 7792 696 7824
rect 728 7792 768 7824
rect 800 7792 840 7824
rect 872 7792 912 7824
rect 944 7792 984 7824
rect 1016 7792 1056 7824
rect 1088 7792 1128 7824
rect 1160 7792 1200 7824
rect 1232 7792 1272 7824
rect 1304 7792 1344 7824
rect 1376 7792 1416 7824
rect 1448 7792 1488 7824
rect 1520 7792 1560 7824
rect 1592 7792 1632 7824
rect 1664 7792 1704 7824
rect 1736 7792 1776 7824
rect 1808 7792 1848 7824
rect 1880 7792 1920 7824
rect 1952 7792 2000 7824
rect 0 7752 2000 7792
rect 0 7720 48 7752
rect 80 7720 120 7752
rect 152 7720 192 7752
rect 224 7720 264 7752
rect 296 7720 336 7752
rect 368 7720 408 7752
rect 440 7720 480 7752
rect 512 7720 552 7752
rect 584 7720 624 7752
rect 656 7720 696 7752
rect 728 7720 768 7752
rect 800 7720 840 7752
rect 872 7720 912 7752
rect 944 7720 984 7752
rect 1016 7720 1056 7752
rect 1088 7720 1128 7752
rect 1160 7720 1200 7752
rect 1232 7720 1272 7752
rect 1304 7720 1344 7752
rect 1376 7720 1416 7752
rect 1448 7720 1488 7752
rect 1520 7720 1560 7752
rect 1592 7720 1632 7752
rect 1664 7720 1704 7752
rect 1736 7720 1776 7752
rect 1808 7720 1848 7752
rect 1880 7720 1920 7752
rect 1952 7720 2000 7752
rect 0 7680 2000 7720
rect 0 7648 48 7680
rect 80 7648 120 7680
rect 152 7648 192 7680
rect 224 7648 264 7680
rect 296 7648 336 7680
rect 368 7648 408 7680
rect 440 7648 480 7680
rect 512 7648 552 7680
rect 584 7648 624 7680
rect 656 7648 696 7680
rect 728 7648 768 7680
rect 800 7648 840 7680
rect 872 7648 912 7680
rect 944 7648 984 7680
rect 1016 7648 1056 7680
rect 1088 7648 1128 7680
rect 1160 7648 1200 7680
rect 1232 7648 1272 7680
rect 1304 7648 1344 7680
rect 1376 7648 1416 7680
rect 1448 7648 1488 7680
rect 1520 7648 1560 7680
rect 1592 7648 1632 7680
rect 1664 7648 1704 7680
rect 1736 7648 1776 7680
rect 1808 7648 1848 7680
rect 1880 7648 1920 7680
rect 1952 7648 2000 7680
rect 0 7608 2000 7648
rect 0 7576 48 7608
rect 80 7576 120 7608
rect 152 7576 192 7608
rect 224 7576 264 7608
rect 296 7576 336 7608
rect 368 7576 408 7608
rect 440 7576 480 7608
rect 512 7576 552 7608
rect 584 7576 624 7608
rect 656 7576 696 7608
rect 728 7576 768 7608
rect 800 7576 840 7608
rect 872 7576 912 7608
rect 944 7576 984 7608
rect 1016 7576 1056 7608
rect 1088 7576 1128 7608
rect 1160 7576 1200 7608
rect 1232 7576 1272 7608
rect 1304 7576 1344 7608
rect 1376 7576 1416 7608
rect 1448 7576 1488 7608
rect 1520 7576 1560 7608
rect 1592 7576 1632 7608
rect 1664 7576 1704 7608
rect 1736 7576 1776 7608
rect 1808 7576 1848 7608
rect 1880 7576 1920 7608
rect 1952 7576 2000 7608
rect 0 7536 2000 7576
rect 0 7504 48 7536
rect 80 7504 120 7536
rect 152 7504 192 7536
rect 224 7504 264 7536
rect 296 7504 336 7536
rect 368 7504 408 7536
rect 440 7504 480 7536
rect 512 7504 552 7536
rect 584 7504 624 7536
rect 656 7504 696 7536
rect 728 7504 768 7536
rect 800 7504 840 7536
rect 872 7504 912 7536
rect 944 7504 984 7536
rect 1016 7504 1056 7536
rect 1088 7504 1128 7536
rect 1160 7504 1200 7536
rect 1232 7504 1272 7536
rect 1304 7504 1344 7536
rect 1376 7504 1416 7536
rect 1448 7504 1488 7536
rect 1520 7504 1560 7536
rect 1592 7504 1632 7536
rect 1664 7504 1704 7536
rect 1736 7504 1776 7536
rect 1808 7504 1848 7536
rect 1880 7504 1920 7536
rect 1952 7504 2000 7536
rect 0 7464 2000 7504
rect 0 7432 48 7464
rect 80 7432 120 7464
rect 152 7432 192 7464
rect 224 7432 264 7464
rect 296 7432 336 7464
rect 368 7432 408 7464
rect 440 7432 480 7464
rect 512 7432 552 7464
rect 584 7432 624 7464
rect 656 7432 696 7464
rect 728 7432 768 7464
rect 800 7432 840 7464
rect 872 7432 912 7464
rect 944 7432 984 7464
rect 1016 7432 1056 7464
rect 1088 7432 1128 7464
rect 1160 7432 1200 7464
rect 1232 7432 1272 7464
rect 1304 7432 1344 7464
rect 1376 7432 1416 7464
rect 1448 7432 1488 7464
rect 1520 7432 1560 7464
rect 1592 7432 1632 7464
rect 1664 7432 1704 7464
rect 1736 7432 1776 7464
rect 1808 7432 1848 7464
rect 1880 7432 1920 7464
rect 1952 7432 2000 7464
rect 0 7392 2000 7432
rect 0 7360 48 7392
rect 80 7360 120 7392
rect 152 7360 192 7392
rect 224 7360 264 7392
rect 296 7360 336 7392
rect 368 7360 408 7392
rect 440 7360 480 7392
rect 512 7360 552 7392
rect 584 7360 624 7392
rect 656 7360 696 7392
rect 728 7360 768 7392
rect 800 7360 840 7392
rect 872 7360 912 7392
rect 944 7360 984 7392
rect 1016 7360 1056 7392
rect 1088 7360 1128 7392
rect 1160 7360 1200 7392
rect 1232 7360 1272 7392
rect 1304 7360 1344 7392
rect 1376 7360 1416 7392
rect 1448 7360 1488 7392
rect 1520 7360 1560 7392
rect 1592 7360 1632 7392
rect 1664 7360 1704 7392
rect 1736 7360 1776 7392
rect 1808 7360 1848 7392
rect 1880 7360 1920 7392
rect 1952 7360 2000 7392
rect 0 7320 2000 7360
rect 0 7288 48 7320
rect 80 7288 120 7320
rect 152 7288 192 7320
rect 224 7288 264 7320
rect 296 7288 336 7320
rect 368 7288 408 7320
rect 440 7288 480 7320
rect 512 7288 552 7320
rect 584 7288 624 7320
rect 656 7288 696 7320
rect 728 7288 768 7320
rect 800 7288 840 7320
rect 872 7288 912 7320
rect 944 7288 984 7320
rect 1016 7288 1056 7320
rect 1088 7288 1128 7320
rect 1160 7288 1200 7320
rect 1232 7288 1272 7320
rect 1304 7288 1344 7320
rect 1376 7288 1416 7320
rect 1448 7288 1488 7320
rect 1520 7288 1560 7320
rect 1592 7288 1632 7320
rect 1664 7288 1704 7320
rect 1736 7288 1776 7320
rect 1808 7288 1848 7320
rect 1880 7288 1920 7320
rect 1952 7288 2000 7320
rect 0 7248 2000 7288
rect 0 7216 48 7248
rect 80 7216 120 7248
rect 152 7216 192 7248
rect 224 7216 264 7248
rect 296 7216 336 7248
rect 368 7216 408 7248
rect 440 7216 480 7248
rect 512 7216 552 7248
rect 584 7216 624 7248
rect 656 7216 696 7248
rect 728 7216 768 7248
rect 800 7216 840 7248
rect 872 7216 912 7248
rect 944 7216 984 7248
rect 1016 7216 1056 7248
rect 1088 7216 1128 7248
rect 1160 7216 1200 7248
rect 1232 7216 1272 7248
rect 1304 7216 1344 7248
rect 1376 7216 1416 7248
rect 1448 7216 1488 7248
rect 1520 7216 1560 7248
rect 1592 7216 1632 7248
rect 1664 7216 1704 7248
rect 1736 7216 1776 7248
rect 1808 7216 1848 7248
rect 1880 7216 1920 7248
rect 1952 7216 2000 7248
rect 0 7176 2000 7216
rect 0 7144 48 7176
rect 80 7144 120 7176
rect 152 7144 192 7176
rect 224 7144 264 7176
rect 296 7144 336 7176
rect 368 7144 408 7176
rect 440 7144 480 7176
rect 512 7144 552 7176
rect 584 7144 624 7176
rect 656 7144 696 7176
rect 728 7144 768 7176
rect 800 7144 840 7176
rect 872 7144 912 7176
rect 944 7144 984 7176
rect 1016 7144 1056 7176
rect 1088 7144 1128 7176
rect 1160 7144 1200 7176
rect 1232 7144 1272 7176
rect 1304 7144 1344 7176
rect 1376 7144 1416 7176
rect 1448 7144 1488 7176
rect 1520 7144 1560 7176
rect 1592 7144 1632 7176
rect 1664 7144 1704 7176
rect 1736 7144 1776 7176
rect 1808 7144 1848 7176
rect 1880 7144 1920 7176
rect 1952 7144 2000 7176
rect 0 7104 2000 7144
rect 0 7072 48 7104
rect 80 7072 120 7104
rect 152 7072 192 7104
rect 224 7072 264 7104
rect 296 7072 336 7104
rect 368 7072 408 7104
rect 440 7072 480 7104
rect 512 7072 552 7104
rect 584 7072 624 7104
rect 656 7072 696 7104
rect 728 7072 768 7104
rect 800 7072 840 7104
rect 872 7072 912 7104
rect 944 7072 984 7104
rect 1016 7072 1056 7104
rect 1088 7072 1128 7104
rect 1160 7072 1200 7104
rect 1232 7072 1272 7104
rect 1304 7072 1344 7104
rect 1376 7072 1416 7104
rect 1448 7072 1488 7104
rect 1520 7072 1560 7104
rect 1592 7072 1632 7104
rect 1664 7072 1704 7104
rect 1736 7072 1776 7104
rect 1808 7072 1848 7104
rect 1880 7072 1920 7104
rect 1952 7072 2000 7104
rect 0 7032 2000 7072
rect 0 7000 48 7032
rect 80 7000 120 7032
rect 152 7000 192 7032
rect 224 7000 264 7032
rect 296 7000 336 7032
rect 368 7000 408 7032
rect 440 7000 480 7032
rect 512 7000 552 7032
rect 584 7000 624 7032
rect 656 7000 696 7032
rect 728 7000 768 7032
rect 800 7000 840 7032
rect 872 7000 912 7032
rect 944 7000 984 7032
rect 1016 7000 1056 7032
rect 1088 7000 1128 7032
rect 1160 7000 1200 7032
rect 1232 7000 1272 7032
rect 1304 7000 1344 7032
rect 1376 7000 1416 7032
rect 1448 7000 1488 7032
rect 1520 7000 1560 7032
rect 1592 7000 1632 7032
rect 1664 7000 1704 7032
rect 1736 7000 1776 7032
rect 1808 7000 1848 7032
rect 1880 7000 1920 7032
rect 1952 7000 2000 7032
rect 0 6960 2000 7000
rect 0 6928 48 6960
rect 80 6928 120 6960
rect 152 6928 192 6960
rect 224 6928 264 6960
rect 296 6928 336 6960
rect 368 6928 408 6960
rect 440 6928 480 6960
rect 512 6928 552 6960
rect 584 6928 624 6960
rect 656 6928 696 6960
rect 728 6928 768 6960
rect 800 6928 840 6960
rect 872 6928 912 6960
rect 944 6928 984 6960
rect 1016 6928 1056 6960
rect 1088 6928 1128 6960
rect 1160 6928 1200 6960
rect 1232 6928 1272 6960
rect 1304 6928 1344 6960
rect 1376 6928 1416 6960
rect 1448 6928 1488 6960
rect 1520 6928 1560 6960
rect 1592 6928 1632 6960
rect 1664 6928 1704 6960
rect 1736 6928 1776 6960
rect 1808 6928 1848 6960
rect 1880 6928 1920 6960
rect 1952 6928 2000 6960
rect 0 6888 2000 6928
rect 0 6856 48 6888
rect 80 6856 120 6888
rect 152 6856 192 6888
rect 224 6856 264 6888
rect 296 6856 336 6888
rect 368 6856 408 6888
rect 440 6856 480 6888
rect 512 6856 552 6888
rect 584 6856 624 6888
rect 656 6856 696 6888
rect 728 6856 768 6888
rect 800 6856 840 6888
rect 872 6856 912 6888
rect 944 6856 984 6888
rect 1016 6856 1056 6888
rect 1088 6856 1128 6888
rect 1160 6856 1200 6888
rect 1232 6856 1272 6888
rect 1304 6856 1344 6888
rect 1376 6856 1416 6888
rect 1448 6856 1488 6888
rect 1520 6856 1560 6888
rect 1592 6856 1632 6888
rect 1664 6856 1704 6888
rect 1736 6856 1776 6888
rect 1808 6856 1848 6888
rect 1880 6856 1920 6888
rect 1952 6856 2000 6888
rect 0 6800 2000 6856
rect 0 6544 2000 6600
rect 0 6512 48 6544
rect 80 6512 120 6544
rect 152 6512 192 6544
rect 224 6512 264 6544
rect 296 6512 336 6544
rect 368 6512 408 6544
rect 440 6512 480 6544
rect 512 6512 552 6544
rect 584 6512 624 6544
rect 656 6512 696 6544
rect 728 6512 768 6544
rect 800 6512 840 6544
rect 872 6512 912 6544
rect 944 6512 984 6544
rect 1016 6512 1056 6544
rect 1088 6512 1128 6544
rect 1160 6512 1200 6544
rect 1232 6512 1272 6544
rect 1304 6512 1344 6544
rect 1376 6512 1416 6544
rect 1448 6512 1488 6544
rect 1520 6512 1560 6544
rect 1592 6512 1632 6544
rect 1664 6512 1704 6544
rect 1736 6512 1776 6544
rect 1808 6512 1848 6544
rect 1880 6512 1920 6544
rect 1952 6512 2000 6544
rect 0 6472 2000 6512
rect 0 6440 48 6472
rect 80 6440 120 6472
rect 152 6440 192 6472
rect 224 6440 264 6472
rect 296 6440 336 6472
rect 368 6440 408 6472
rect 440 6440 480 6472
rect 512 6440 552 6472
rect 584 6440 624 6472
rect 656 6440 696 6472
rect 728 6440 768 6472
rect 800 6440 840 6472
rect 872 6440 912 6472
rect 944 6440 984 6472
rect 1016 6440 1056 6472
rect 1088 6440 1128 6472
rect 1160 6440 1200 6472
rect 1232 6440 1272 6472
rect 1304 6440 1344 6472
rect 1376 6440 1416 6472
rect 1448 6440 1488 6472
rect 1520 6440 1560 6472
rect 1592 6440 1632 6472
rect 1664 6440 1704 6472
rect 1736 6440 1776 6472
rect 1808 6440 1848 6472
rect 1880 6440 1920 6472
rect 1952 6440 2000 6472
rect 0 6400 2000 6440
rect 0 6368 48 6400
rect 80 6368 120 6400
rect 152 6368 192 6400
rect 224 6368 264 6400
rect 296 6368 336 6400
rect 368 6368 408 6400
rect 440 6368 480 6400
rect 512 6368 552 6400
rect 584 6368 624 6400
rect 656 6368 696 6400
rect 728 6368 768 6400
rect 800 6368 840 6400
rect 872 6368 912 6400
rect 944 6368 984 6400
rect 1016 6368 1056 6400
rect 1088 6368 1128 6400
rect 1160 6368 1200 6400
rect 1232 6368 1272 6400
rect 1304 6368 1344 6400
rect 1376 6368 1416 6400
rect 1448 6368 1488 6400
rect 1520 6368 1560 6400
rect 1592 6368 1632 6400
rect 1664 6368 1704 6400
rect 1736 6368 1776 6400
rect 1808 6368 1848 6400
rect 1880 6368 1920 6400
rect 1952 6368 2000 6400
rect 0 6328 2000 6368
rect 0 6296 48 6328
rect 80 6296 120 6328
rect 152 6296 192 6328
rect 224 6296 264 6328
rect 296 6296 336 6328
rect 368 6296 408 6328
rect 440 6296 480 6328
rect 512 6296 552 6328
rect 584 6296 624 6328
rect 656 6296 696 6328
rect 728 6296 768 6328
rect 800 6296 840 6328
rect 872 6296 912 6328
rect 944 6296 984 6328
rect 1016 6296 1056 6328
rect 1088 6296 1128 6328
rect 1160 6296 1200 6328
rect 1232 6296 1272 6328
rect 1304 6296 1344 6328
rect 1376 6296 1416 6328
rect 1448 6296 1488 6328
rect 1520 6296 1560 6328
rect 1592 6296 1632 6328
rect 1664 6296 1704 6328
rect 1736 6296 1776 6328
rect 1808 6296 1848 6328
rect 1880 6296 1920 6328
rect 1952 6296 2000 6328
rect 0 6256 2000 6296
rect 0 6224 48 6256
rect 80 6224 120 6256
rect 152 6224 192 6256
rect 224 6224 264 6256
rect 296 6224 336 6256
rect 368 6224 408 6256
rect 440 6224 480 6256
rect 512 6224 552 6256
rect 584 6224 624 6256
rect 656 6224 696 6256
rect 728 6224 768 6256
rect 800 6224 840 6256
rect 872 6224 912 6256
rect 944 6224 984 6256
rect 1016 6224 1056 6256
rect 1088 6224 1128 6256
rect 1160 6224 1200 6256
rect 1232 6224 1272 6256
rect 1304 6224 1344 6256
rect 1376 6224 1416 6256
rect 1448 6224 1488 6256
rect 1520 6224 1560 6256
rect 1592 6224 1632 6256
rect 1664 6224 1704 6256
rect 1736 6224 1776 6256
rect 1808 6224 1848 6256
rect 1880 6224 1920 6256
rect 1952 6224 2000 6256
rect 0 6184 2000 6224
rect 0 6152 48 6184
rect 80 6152 120 6184
rect 152 6152 192 6184
rect 224 6152 264 6184
rect 296 6152 336 6184
rect 368 6152 408 6184
rect 440 6152 480 6184
rect 512 6152 552 6184
rect 584 6152 624 6184
rect 656 6152 696 6184
rect 728 6152 768 6184
rect 800 6152 840 6184
rect 872 6152 912 6184
rect 944 6152 984 6184
rect 1016 6152 1056 6184
rect 1088 6152 1128 6184
rect 1160 6152 1200 6184
rect 1232 6152 1272 6184
rect 1304 6152 1344 6184
rect 1376 6152 1416 6184
rect 1448 6152 1488 6184
rect 1520 6152 1560 6184
rect 1592 6152 1632 6184
rect 1664 6152 1704 6184
rect 1736 6152 1776 6184
rect 1808 6152 1848 6184
rect 1880 6152 1920 6184
rect 1952 6152 2000 6184
rect 0 6112 2000 6152
rect 0 6080 48 6112
rect 80 6080 120 6112
rect 152 6080 192 6112
rect 224 6080 264 6112
rect 296 6080 336 6112
rect 368 6080 408 6112
rect 440 6080 480 6112
rect 512 6080 552 6112
rect 584 6080 624 6112
rect 656 6080 696 6112
rect 728 6080 768 6112
rect 800 6080 840 6112
rect 872 6080 912 6112
rect 944 6080 984 6112
rect 1016 6080 1056 6112
rect 1088 6080 1128 6112
rect 1160 6080 1200 6112
rect 1232 6080 1272 6112
rect 1304 6080 1344 6112
rect 1376 6080 1416 6112
rect 1448 6080 1488 6112
rect 1520 6080 1560 6112
rect 1592 6080 1632 6112
rect 1664 6080 1704 6112
rect 1736 6080 1776 6112
rect 1808 6080 1848 6112
rect 1880 6080 1920 6112
rect 1952 6080 2000 6112
rect 0 6040 2000 6080
rect 0 6008 48 6040
rect 80 6008 120 6040
rect 152 6008 192 6040
rect 224 6008 264 6040
rect 296 6008 336 6040
rect 368 6008 408 6040
rect 440 6008 480 6040
rect 512 6008 552 6040
rect 584 6008 624 6040
rect 656 6008 696 6040
rect 728 6008 768 6040
rect 800 6008 840 6040
rect 872 6008 912 6040
rect 944 6008 984 6040
rect 1016 6008 1056 6040
rect 1088 6008 1128 6040
rect 1160 6008 1200 6040
rect 1232 6008 1272 6040
rect 1304 6008 1344 6040
rect 1376 6008 1416 6040
rect 1448 6008 1488 6040
rect 1520 6008 1560 6040
rect 1592 6008 1632 6040
rect 1664 6008 1704 6040
rect 1736 6008 1776 6040
rect 1808 6008 1848 6040
rect 1880 6008 1920 6040
rect 1952 6008 2000 6040
rect 0 5968 2000 6008
rect 0 5936 48 5968
rect 80 5936 120 5968
rect 152 5936 192 5968
rect 224 5936 264 5968
rect 296 5936 336 5968
rect 368 5936 408 5968
rect 440 5936 480 5968
rect 512 5936 552 5968
rect 584 5936 624 5968
rect 656 5936 696 5968
rect 728 5936 768 5968
rect 800 5936 840 5968
rect 872 5936 912 5968
rect 944 5936 984 5968
rect 1016 5936 1056 5968
rect 1088 5936 1128 5968
rect 1160 5936 1200 5968
rect 1232 5936 1272 5968
rect 1304 5936 1344 5968
rect 1376 5936 1416 5968
rect 1448 5936 1488 5968
rect 1520 5936 1560 5968
rect 1592 5936 1632 5968
rect 1664 5936 1704 5968
rect 1736 5936 1776 5968
rect 1808 5936 1848 5968
rect 1880 5936 1920 5968
rect 1952 5936 2000 5968
rect 0 5896 2000 5936
rect 0 5864 48 5896
rect 80 5864 120 5896
rect 152 5864 192 5896
rect 224 5864 264 5896
rect 296 5864 336 5896
rect 368 5864 408 5896
rect 440 5864 480 5896
rect 512 5864 552 5896
rect 584 5864 624 5896
rect 656 5864 696 5896
rect 728 5864 768 5896
rect 800 5864 840 5896
rect 872 5864 912 5896
rect 944 5864 984 5896
rect 1016 5864 1056 5896
rect 1088 5864 1128 5896
rect 1160 5864 1200 5896
rect 1232 5864 1272 5896
rect 1304 5864 1344 5896
rect 1376 5864 1416 5896
rect 1448 5864 1488 5896
rect 1520 5864 1560 5896
rect 1592 5864 1632 5896
rect 1664 5864 1704 5896
rect 1736 5864 1776 5896
rect 1808 5864 1848 5896
rect 1880 5864 1920 5896
rect 1952 5864 2000 5896
rect 0 5824 2000 5864
rect 0 5792 48 5824
rect 80 5792 120 5824
rect 152 5792 192 5824
rect 224 5792 264 5824
rect 296 5792 336 5824
rect 368 5792 408 5824
rect 440 5792 480 5824
rect 512 5792 552 5824
rect 584 5792 624 5824
rect 656 5792 696 5824
rect 728 5792 768 5824
rect 800 5792 840 5824
rect 872 5792 912 5824
rect 944 5792 984 5824
rect 1016 5792 1056 5824
rect 1088 5792 1128 5824
rect 1160 5792 1200 5824
rect 1232 5792 1272 5824
rect 1304 5792 1344 5824
rect 1376 5792 1416 5824
rect 1448 5792 1488 5824
rect 1520 5792 1560 5824
rect 1592 5792 1632 5824
rect 1664 5792 1704 5824
rect 1736 5792 1776 5824
rect 1808 5792 1848 5824
rect 1880 5792 1920 5824
rect 1952 5792 2000 5824
rect 0 5752 2000 5792
rect 0 5720 48 5752
rect 80 5720 120 5752
rect 152 5720 192 5752
rect 224 5720 264 5752
rect 296 5720 336 5752
rect 368 5720 408 5752
rect 440 5720 480 5752
rect 512 5720 552 5752
rect 584 5720 624 5752
rect 656 5720 696 5752
rect 728 5720 768 5752
rect 800 5720 840 5752
rect 872 5720 912 5752
rect 944 5720 984 5752
rect 1016 5720 1056 5752
rect 1088 5720 1128 5752
rect 1160 5720 1200 5752
rect 1232 5720 1272 5752
rect 1304 5720 1344 5752
rect 1376 5720 1416 5752
rect 1448 5720 1488 5752
rect 1520 5720 1560 5752
rect 1592 5720 1632 5752
rect 1664 5720 1704 5752
rect 1736 5720 1776 5752
rect 1808 5720 1848 5752
rect 1880 5720 1920 5752
rect 1952 5720 2000 5752
rect 0 5680 2000 5720
rect 0 5648 48 5680
rect 80 5648 120 5680
rect 152 5648 192 5680
rect 224 5648 264 5680
rect 296 5648 336 5680
rect 368 5648 408 5680
rect 440 5648 480 5680
rect 512 5648 552 5680
rect 584 5648 624 5680
rect 656 5648 696 5680
rect 728 5648 768 5680
rect 800 5648 840 5680
rect 872 5648 912 5680
rect 944 5648 984 5680
rect 1016 5648 1056 5680
rect 1088 5648 1128 5680
rect 1160 5648 1200 5680
rect 1232 5648 1272 5680
rect 1304 5648 1344 5680
rect 1376 5648 1416 5680
rect 1448 5648 1488 5680
rect 1520 5648 1560 5680
rect 1592 5648 1632 5680
rect 1664 5648 1704 5680
rect 1736 5648 1776 5680
rect 1808 5648 1848 5680
rect 1880 5648 1920 5680
rect 1952 5648 2000 5680
rect 0 5608 2000 5648
rect 0 5576 48 5608
rect 80 5576 120 5608
rect 152 5576 192 5608
rect 224 5576 264 5608
rect 296 5576 336 5608
rect 368 5576 408 5608
rect 440 5576 480 5608
rect 512 5576 552 5608
rect 584 5576 624 5608
rect 656 5576 696 5608
rect 728 5576 768 5608
rect 800 5576 840 5608
rect 872 5576 912 5608
rect 944 5576 984 5608
rect 1016 5576 1056 5608
rect 1088 5576 1128 5608
rect 1160 5576 1200 5608
rect 1232 5576 1272 5608
rect 1304 5576 1344 5608
rect 1376 5576 1416 5608
rect 1448 5576 1488 5608
rect 1520 5576 1560 5608
rect 1592 5576 1632 5608
rect 1664 5576 1704 5608
rect 1736 5576 1776 5608
rect 1808 5576 1848 5608
rect 1880 5576 1920 5608
rect 1952 5576 2000 5608
rect 0 5536 2000 5576
rect 0 5504 48 5536
rect 80 5504 120 5536
rect 152 5504 192 5536
rect 224 5504 264 5536
rect 296 5504 336 5536
rect 368 5504 408 5536
rect 440 5504 480 5536
rect 512 5504 552 5536
rect 584 5504 624 5536
rect 656 5504 696 5536
rect 728 5504 768 5536
rect 800 5504 840 5536
rect 872 5504 912 5536
rect 944 5504 984 5536
rect 1016 5504 1056 5536
rect 1088 5504 1128 5536
rect 1160 5504 1200 5536
rect 1232 5504 1272 5536
rect 1304 5504 1344 5536
rect 1376 5504 1416 5536
rect 1448 5504 1488 5536
rect 1520 5504 1560 5536
rect 1592 5504 1632 5536
rect 1664 5504 1704 5536
rect 1736 5504 1776 5536
rect 1808 5504 1848 5536
rect 1880 5504 1920 5536
rect 1952 5504 2000 5536
rect 0 5464 2000 5504
rect 0 5432 48 5464
rect 80 5432 120 5464
rect 152 5432 192 5464
rect 224 5432 264 5464
rect 296 5432 336 5464
rect 368 5432 408 5464
rect 440 5432 480 5464
rect 512 5432 552 5464
rect 584 5432 624 5464
rect 656 5432 696 5464
rect 728 5432 768 5464
rect 800 5432 840 5464
rect 872 5432 912 5464
rect 944 5432 984 5464
rect 1016 5432 1056 5464
rect 1088 5432 1128 5464
rect 1160 5432 1200 5464
rect 1232 5432 1272 5464
rect 1304 5432 1344 5464
rect 1376 5432 1416 5464
rect 1448 5432 1488 5464
rect 1520 5432 1560 5464
rect 1592 5432 1632 5464
rect 1664 5432 1704 5464
rect 1736 5432 1776 5464
rect 1808 5432 1848 5464
rect 1880 5432 1920 5464
rect 1952 5432 2000 5464
rect 0 5392 2000 5432
rect 0 5360 48 5392
rect 80 5360 120 5392
rect 152 5360 192 5392
rect 224 5360 264 5392
rect 296 5360 336 5392
rect 368 5360 408 5392
rect 440 5360 480 5392
rect 512 5360 552 5392
rect 584 5360 624 5392
rect 656 5360 696 5392
rect 728 5360 768 5392
rect 800 5360 840 5392
rect 872 5360 912 5392
rect 944 5360 984 5392
rect 1016 5360 1056 5392
rect 1088 5360 1128 5392
rect 1160 5360 1200 5392
rect 1232 5360 1272 5392
rect 1304 5360 1344 5392
rect 1376 5360 1416 5392
rect 1448 5360 1488 5392
rect 1520 5360 1560 5392
rect 1592 5360 1632 5392
rect 1664 5360 1704 5392
rect 1736 5360 1776 5392
rect 1808 5360 1848 5392
rect 1880 5360 1920 5392
rect 1952 5360 2000 5392
rect 0 5320 2000 5360
rect 0 5288 48 5320
rect 80 5288 120 5320
rect 152 5288 192 5320
rect 224 5288 264 5320
rect 296 5288 336 5320
rect 368 5288 408 5320
rect 440 5288 480 5320
rect 512 5288 552 5320
rect 584 5288 624 5320
rect 656 5288 696 5320
rect 728 5288 768 5320
rect 800 5288 840 5320
rect 872 5288 912 5320
rect 944 5288 984 5320
rect 1016 5288 1056 5320
rect 1088 5288 1128 5320
rect 1160 5288 1200 5320
rect 1232 5288 1272 5320
rect 1304 5288 1344 5320
rect 1376 5288 1416 5320
rect 1448 5288 1488 5320
rect 1520 5288 1560 5320
rect 1592 5288 1632 5320
rect 1664 5288 1704 5320
rect 1736 5288 1776 5320
rect 1808 5288 1848 5320
rect 1880 5288 1920 5320
rect 1952 5288 2000 5320
rect 0 5248 2000 5288
rect 0 5216 48 5248
rect 80 5216 120 5248
rect 152 5216 192 5248
rect 224 5216 264 5248
rect 296 5216 336 5248
rect 368 5216 408 5248
rect 440 5216 480 5248
rect 512 5216 552 5248
rect 584 5216 624 5248
rect 656 5216 696 5248
rect 728 5216 768 5248
rect 800 5216 840 5248
rect 872 5216 912 5248
rect 944 5216 984 5248
rect 1016 5216 1056 5248
rect 1088 5216 1128 5248
rect 1160 5216 1200 5248
rect 1232 5216 1272 5248
rect 1304 5216 1344 5248
rect 1376 5216 1416 5248
rect 1448 5216 1488 5248
rect 1520 5216 1560 5248
rect 1592 5216 1632 5248
rect 1664 5216 1704 5248
rect 1736 5216 1776 5248
rect 1808 5216 1848 5248
rect 1880 5216 1920 5248
rect 1952 5216 2000 5248
rect 0 5176 2000 5216
rect 0 5144 48 5176
rect 80 5144 120 5176
rect 152 5144 192 5176
rect 224 5144 264 5176
rect 296 5144 336 5176
rect 368 5144 408 5176
rect 440 5144 480 5176
rect 512 5144 552 5176
rect 584 5144 624 5176
rect 656 5144 696 5176
rect 728 5144 768 5176
rect 800 5144 840 5176
rect 872 5144 912 5176
rect 944 5144 984 5176
rect 1016 5144 1056 5176
rect 1088 5144 1128 5176
rect 1160 5144 1200 5176
rect 1232 5144 1272 5176
rect 1304 5144 1344 5176
rect 1376 5144 1416 5176
rect 1448 5144 1488 5176
rect 1520 5144 1560 5176
rect 1592 5144 1632 5176
rect 1664 5144 1704 5176
rect 1736 5144 1776 5176
rect 1808 5144 1848 5176
rect 1880 5144 1920 5176
rect 1952 5144 2000 5176
rect 0 5104 2000 5144
rect 0 5072 48 5104
rect 80 5072 120 5104
rect 152 5072 192 5104
rect 224 5072 264 5104
rect 296 5072 336 5104
rect 368 5072 408 5104
rect 440 5072 480 5104
rect 512 5072 552 5104
rect 584 5072 624 5104
rect 656 5072 696 5104
rect 728 5072 768 5104
rect 800 5072 840 5104
rect 872 5072 912 5104
rect 944 5072 984 5104
rect 1016 5072 1056 5104
rect 1088 5072 1128 5104
rect 1160 5072 1200 5104
rect 1232 5072 1272 5104
rect 1304 5072 1344 5104
rect 1376 5072 1416 5104
rect 1448 5072 1488 5104
rect 1520 5072 1560 5104
rect 1592 5072 1632 5104
rect 1664 5072 1704 5104
rect 1736 5072 1776 5104
rect 1808 5072 1848 5104
rect 1880 5072 1920 5104
rect 1952 5072 2000 5104
rect 0 5032 2000 5072
rect 0 5000 48 5032
rect 80 5000 120 5032
rect 152 5000 192 5032
rect 224 5000 264 5032
rect 296 5000 336 5032
rect 368 5000 408 5032
rect 440 5000 480 5032
rect 512 5000 552 5032
rect 584 5000 624 5032
rect 656 5000 696 5032
rect 728 5000 768 5032
rect 800 5000 840 5032
rect 872 5000 912 5032
rect 944 5000 984 5032
rect 1016 5000 1056 5032
rect 1088 5000 1128 5032
rect 1160 5000 1200 5032
rect 1232 5000 1272 5032
rect 1304 5000 1344 5032
rect 1376 5000 1416 5032
rect 1448 5000 1488 5032
rect 1520 5000 1560 5032
rect 1592 5000 1632 5032
rect 1664 5000 1704 5032
rect 1736 5000 1776 5032
rect 1808 5000 1848 5032
rect 1880 5000 1920 5032
rect 1952 5000 2000 5032
rect 0 4960 2000 5000
rect 0 4928 48 4960
rect 80 4928 120 4960
rect 152 4928 192 4960
rect 224 4928 264 4960
rect 296 4928 336 4960
rect 368 4928 408 4960
rect 440 4928 480 4960
rect 512 4928 552 4960
rect 584 4928 624 4960
rect 656 4928 696 4960
rect 728 4928 768 4960
rect 800 4928 840 4960
rect 872 4928 912 4960
rect 944 4928 984 4960
rect 1016 4928 1056 4960
rect 1088 4928 1128 4960
rect 1160 4928 1200 4960
rect 1232 4928 1272 4960
rect 1304 4928 1344 4960
rect 1376 4928 1416 4960
rect 1448 4928 1488 4960
rect 1520 4928 1560 4960
rect 1592 4928 1632 4960
rect 1664 4928 1704 4960
rect 1736 4928 1776 4960
rect 1808 4928 1848 4960
rect 1880 4928 1920 4960
rect 1952 4928 2000 4960
rect 0 4888 2000 4928
rect 0 4856 48 4888
rect 80 4856 120 4888
rect 152 4856 192 4888
rect 224 4856 264 4888
rect 296 4856 336 4888
rect 368 4856 408 4888
rect 440 4856 480 4888
rect 512 4856 552 4888
rect 584 4856 624 4888
rect 656 4856 696 4888
rect 728 4856 768 4888
rect 800 4856 840 4888
rect 872 4856 912 4888
rect 944 4856 984 4888
rect 1016 4856 1056 4888
rect 1088 4856 1128 4888
rect 1160 4856 1200 4888
rect 1232 4856 1272 4888
rect 1304 4856 1344 4888
rect 1376 4856 1416 4888
rect 1448 4856 1488 4888
rect 1520 4856 1560 4888
rect 1592 4856 1632 4888
rect 1664 4856 1704 4888
rect 1736 4856 1776 4888
rect 1808 4856 1848 4888
rect 1880 4856 1920 4888
rect 1952 4856 2000 4888
rect 0 4816 2000 4856
rect 0 4784 48 4816
rect 80 4784 120 4816
rect 152 4784 192 4816
rect 224 4784 264 4816
rect 296 4784 336 4816
rect 368 4784 408 4816
rect 440 4784 480 4816
rect 512 4784 552 4816
rect 584 4784 624 4816
rect 656 4784 696 4816
rect 728 4784 768 4816
rect 800 4784 840 4816
rect 872 4784 912 4816
rect 944 4784 984 4816
rect 1016 4784 1056 4816
rect 1088 4784 1128 4816
rect 1160 4784 1200 4816
rect 1232 4784 1272 4816
rect 1304 4784 1344 4816
rect 1376 4784 1416 4816
rect 1448 4784 1488 4816
rect 1520 4784 1560 4816
rect 1592 4784 1632 4816
rect 1664 4784 1704 4816
rect 1736 4784 1776 4816
rect 1808 4784 1848 4816
rect 1880 4784 1920 4816
rect 1952 4784 2000 4816
rect 0 4744 2000 4784
rect 0 4712 48 4744
rect 80 4712 120 4744
rect 152 4712 192 4744
rect 224 4712 264 4744
rect 296 4712 336 4744
rect 368 4712 408 4744
rect 440 4712 480 4744
rect 512 4712 552 4744
rect 584 4712 624 4744
rect 656 4712 696 4744
rect 728 4712 768 4744
rect 800 4712 840 4744
rect 872 4712 912 4744
rect 944 4712 984 4744
rect 1016 4712 1056 4744
rect 1088 4712 1128 4744
rect 1160 4712 1200 4744
rect 1232 4712 1272 4744
rect 1304 4712 1344 4744
rect 1376 4712 1416 4744
rect 1448 4712 1488 4744
rect 1520 4712 1560 4744
rect 1592 4712 1632 4744
rect 1664 4712 1704 4744
rect 1736 4712 1776 4744
rect 1808 4712 1848 4744
rect 1880 4712 1920 4744
rect 1952 4712 2000 4744
rect 0 4672 2000 4712
rect 0 4640 48 4672
rect 80 4640 120 4672
rect 152 4640 192 4672
rect 224 4640 264 4672
rect 296 4640 336 4672
rect 368 4640 408 4672
rect 440 4640 480 4672
rect 512 4640 552 4672
rect 584 4640 624 4672
rect 656 4640 696 4672
rect 728 4640 768 4672
rect 800 4640 840 4672
rect 872 4640 912 4672
rect 944 4640 984 4672
rect 1016 4640 1056 4672
rect 1088 4640 1128 4672
rect 1160 4640 1200 4672
rect 1232 4640 1272 4672
rect 1304 4640 1344 4672
rect 1376 4640 1416 4672
rect 1448 4640 1488 4672
rect 1520 4640 1560 4672
rect 1592 4640 1632 4672
rect 1664 4640 1704 4672
rect 1736 4640 1776 4672
rect 1808 4640 1848 4672
rect 1880 4640 1920 4672
rect 1952 4640 2000 4672
rect 0 4600 2000 4640
rect 0 4568 48 4600
rect 80 4568 120 4600
rect 152 4568 192 4600
rect 224 4568 264 4600
rect 296 4568 336 4600
rect 368 4568 408 4600
rect 440 4568 480 4600
rect 512 4568 552 4600
rect 584 4568 624 4600
rect 656 4568 696 4600
rect 728 4568 768 4600
rect 800 4568 840 4600
rect 872 4568 912 4600
rect 944 4568 984 4600
rect 1016 4568 1056 4600
rect 1088 4568 1128 4600
rect 1160 4568 1200 4600
rect 1232 4568 1272 4600
rect 1304 4568 1344 4600
rect 1376 4568 1416 4600
rect 1448 4568 1488 4600
rect 1520 4568 1560 4600
rect 1592 4568 1632 4600
rect 1664 4568 1704 4600
rect 1736 4568 1776 4600
rect 1808 4568 1848 4600
rect 1880 4568 1920 4600
rect 1952 4568 2000 4600
rect 0 4528 2000 4568
rect 0 4496 48 4528
rect 80 4496 120 4528
rect 152 4496 192 4528
rect 224 4496 264 4528
rect 296 4496 336 4528
rect 368 4496 408 4528
rect 440 4496 480 4528
rect 512 4496 552 4528
rect 584 4496 624 4528
rect 656 4496 696 4528
rect 728 4496 768 4528
rect 800 4496 840 4528
rect 872 4496 912 4528
rect 944 4496 984 4528
rect 1016 4496 1056 4528
rect 1088 4496 1128 4528
rect 1160 4496 1200 4528
rect 1232 4496 1272 4528
rect 1304 4496 1344 4528
rect 1376 4496 1416 4528
rect 1448 4496 1488 4528
rect 1520 4496 1560 4528
rect 1592 4496 1632 4528
rect 1664 4496 1704 4528
rect 1736 4496 1776 4528
rect 1808 4496 1848 4528
rect 1880 4496 1920 4528
rect 1952 4496 2000 4528
rect 0 4456 2000 4496
rect 0 4424 48 4456
rect 80 4424 120 4456
rect 152 4424 192 4456
rect 224 4424 264 4456
rect 296 4424 336 4456
rect 368 4424 408 4456
rect 440 4424 480 4456
rect 512 4424 552 4456
rect 584 4424 624 4456
rect 656 4424 696 4456
rect 728 4424 768 4456
rect 800 4424 840 4456
rect 872 4424 912 4456
rect 944 4424 984 4456
rect 1016 4424 1056 4456
rect 1088 4424 1128 4456
rect 1160 4424 1200 4456
rect 1232 4424 1272 4456
rect 1304 4424 1344 4456
rect 1376 4424 1416 4456
rect 1448 4424 1488 4456
rect 1520 4424 1560 4456
rect 1592 4424 1632 4456
rect 1664 4424 1704 4456
rect 1736 4424 1776 4456
rect 1808 4424 1848 4456
rect 1880 4424 1920 4456
rect 1952 4424 2000 4456
rect 0 4384 2000 4424
rect 0 4352 48 4384
rect 80 4352 120 4384
rect 152 4352 192 4384
rect 224 4352 264 4384
rect 296 4352 336 4384
rect 368 4352 408 4384
rect 440 4352 480 4384
rect 512 4352 552 4384
rect 584 4352 624 4384
rect 656 4352 696 4384
rect 728 4352 768 4384
rect 800 4352 840 4384
rect 872 4352 912 4384
rect 944 4352 984 4384
rect 1016 4352 1056 4384
rect 1088 4352 1128 4384
rect 1160 4352 1200 4384
rect 1232 4352 1272 4384
rect 1304 4352 1344 4384
rect 1376 4352 1416 4384
rect 1448 4352 1488 4384
rect 1520 4352 1560 4384
rect 1592 4352 1632 4384
rect 1664 4352 1704 4384
rect 1736 4352 1776 4384
rect 1808 4352 1848 4384
rect 1880 4352 1920 4384
rect 1952 4352 2000 4384
rect 0 4312 2000 4352
rect 0 4280 48 4312
rect 80 4280 120 4312
rect 152 4280 192 4312
rect 224 4280 264 4312
rect 296 4280 336 4312
rect 368 4280 408 4312
rect 440 4280 480 4312
rect 512 4280 552 4312
rect 584 4280 624 4312
rect 656 4280 696 4312
rect 728 4280 768 4312
rect 800 4280 840 4312
rect 872 4280 912 4312
rect 944 4280 984 4312
rect 1016 4280 1056 4312
rect 1088 4280 1128 4312
rect 1160 4280 1200 4312
rect 1232 4280 1272 4312
rect 1304 4280 1344 4312
rect 1376 4280 1416 4312
rect 1448 4280 1488 4312
rect 1520 4280 1560 4312
rect 1592 4280 1632 4312
rect 1664 4280 1704 4312
rect 1736 4280 1776 4312
rect 1808 4280 1848 4312
rect 1880 4280 1920 4312
rect 1952 4280 2000 4312
rect 0 4240 2000 4280
rect 0 4208 48 4240
rect 80 4208 120 4240
rect 152 4208 192 4240
rect 224 4208 264 4240
rect 296 4208 336 4240
rect 368 4208 408 4240
rect 440 4208 480 4240
rect 512 4208 552 4240
rect 584 4208 624 4240
rect 656 4208 696 4240
rect 728 4208 768 4240
rect 800 4208 840 4240
rect 872 4208 912 4240
rect 944 4208 984 4240
rect 1016 4208 1056 4240
rect 1088 4208 1128 4240
rect 1160 4208 1200 4240
rect 1232 4208 1272 4240
rect 1304 4208 1344 4240
rect 1376 4208 1416 4240
rect 1448 4208 1488 4240
rect 1520 4208 1560 4240
rect 1592 4208 1632 4240
rect 1664 4208 1704 4240
rect 1736 4208 1776 4240
rect 1808 4208 1848 4240
rect 1880 4208 1920 4240
rect 1952 4208 2000 4240
rect 0 4168 2000 4208
rect 0 4136 48 4168
rect 80 4136 120 4168
rect 152 4136 192 4168
rect 224 4136 264 4168
rect 296 4136 336 4168
rect 368 4136 408 4168
rect 440 4136 480 4168
rect 512 4136 552 4168
rect 584 4136 624 4168
rect 656 4136 696 4168
rect 728 4136 768 4168
rect 800 4136 840 4168
rect 872 4136 912 4168
rect 944 4136 984 4168
rect 1016 4136 1056 4168
rect 1088 4136 1128 4168
rect 1160 4136 1200 4168
rect 1232 4136 1272 4168
rect 1304 4136 1344 4168
rect 1376 4136 1416 4168
rect 1448 4136 1488 4168
rect 1520 4136 1560 4168
rect 1592 4136 1632 4168
rect 1664 4136 1704 4168
rect 1736 4136 1776 4168
rect 1808 4136 1848 4168
rect 1880 4136 1920 4168
rect 1952 4136 2000 4168
rect 0 4096 2000 4136
rect 0 4064 48 4096
rect 80 4064 120 4096
rect 152 4064 192 4096
rect 224 4064 264 4096
rect 296 4064 336 4096
rect 368 4064 408 4096
rect 440 4064 480 4096
rect 512 4064 552 4096
rect 584 4064 624 4096
rect 656 4064 696 4096
rect 728 4064 768 4096
rect 800 4064 840 4096
rect 872 4064 912 4096
rect 944 4064 984 4096
rect 1016 4064 1056 4096
rect 1088 4064 1128 4096
rect 1160 4064 1200 4096
rect 1232 4064 1272 4096
rect 1304 4064 1344 4096
rect 1376 4064 1416 4096
rect 1448 4064 1488 4096
rect 1520 4064 1560 4096
rect 1592 4064 1632 4096
rect 1664 4064 1704 4096
rect 1736 4064 1776 4096
rect 1808 4064 1848 4096
rect 1880 4064 1920 4096
rect 1952 4064 2000 4096
rect 0 4024 2000 4064
rect 0 3992 48 4024
rect 80 3992 120 4024
rect 152 3992 192 4024
rect 224 3992 264 4024
rect 296 3992 336 4024
rect 368 3992 408 4024
rect 440 3992 480 4024
rect 512 3992 552 4024
rect 584 3992 624 4024
rect 656 3992 696 4024
rect 728 3992 768 4024
rect 800 3992 840 4024
rect 872 3992 912 4024
rect 944 3992 984 4024
rect 1016 3992 1056 4024
rect 1088 3992 1128 4024
rect 1160 3992 1200 4024
rect 1232 3992 1272 4024
rect 1304 3992 1344 4024
rect 1376 3992 1416 4024
rect 1448 3992 1488 4024
rect 1520 3992 1560 4024
rect 1592 3992 1632 4024
rect 1664 3992 1704 4024
rect 1736 3992 1776 4024
rect 1808 3992 1848 4024
rect 1880 3992 1920 4024
rect 1952 3992 2000 4024
rect 0 3952 2000 3992
rect 0 3920 48 3952
rect 80 3920 120 3952
rect 152 3920 192 3952
rect 224 3920 264 3952
rect 296 3920 336 3952
rect 368 3920 408 3952
rect 440 3920 480 3952
rect 512 3920 552 3952
rect 584 3920 624 3952
rect 656 3920 696 3952
rect 728 3920 768 3952
rect 800 3920 840 3952
rect 872 3920 912 3952
rect 944 3920 984 3952
rect 1016 3920 1056 3952
rect 1088 3920 1128 3952
rect 1160 3920 1200 3952
rect 1232 3920 1272 3952
rect 1304 3920 1344 3952
rect 1376 3920 1416 3952
rect 1448 3920 1488 3952
rect 1520 3920 1560 3952
rect 1592 3920 1632 3952
rect 1664 3920 1704 3952
rect 1736 3920 1776 3952
rect 1808 3920 1848 3952
rect 1880 3920 1920 3952
rect 1952 3920 2000 3952
rect 0 3880 2000 3920
rect 0 3848 48 3880
rect 80 3848 120 3880
rect 152 3848 192 3880
rect 224 3848 264 3880
rect 296 3848 336 3880
rect 368 3848 408 3880
rect 440 3848 480 3880
rect 512 3848 552 3880
rect 584 3848 624 3880
rect 656 3848 696 3880
rect 728 3848 768 3880
rect 800 3848 840 3880
rect 872 3848 912 3880
rect 944 3848 984 3880
rect 1016 3848 1056 3880
rect 1088 3848 1128 3880
rect 1160 3848 1200 3880
rect 1232 3848 1272 3880
rect 1304 3848 1344 3880
rect 1376 3848 1416 3880
rect 1448 3848 1488 3880
rect 1520 3848 1560 3880
rect 1592 3848 1632 3880
rect 1664 3848 1704 3880
rect 1736 3848 1776 3880
rect 1808 3848 1848 3880
rect 1880 3848 1920 3880
rect 1952 3848 2000 3880
rect 0 3808 2000 3848
rect 0 3776 48 3808
rect 80 3776 120 3808
rect 152 3776 192 3808
rect 224 3776 264 3808
rect 296 3776 336 3808
rect 368 3776 408 3808
rect 440 3776 480 3808
rect 512 3776 552 3808
rect 584 3776 624 3808
rect 656 3776 696 3808
rect 728 3776 768 3808
rect 800 3776 840 3808
rect 872 3776 912 3808
rect 944 3776 984 3808
rect 1016 3776 1056 3808
rect 1088 3776 1128 3808
rect 1160 3776 1200 3808
rect 1232 3776 1272 3808
rect 1304 3776 1344 3808
rect 1376 3776 1416 3808
rect 1448 3776 1488 3808
rect 1520 3776 1560 3808
rect 1592 3776 1632 3808
rect 1664 3776 1704 3808
rect 1736 3776 1776 3808
rect 1808 3776 1848 3808
rect 1880 3776 1920 3808
rect 1952 3776 2000 3808
rect 0 3736 2000 3776
rect 0 3704 48 3736
rect 80 3704 120 3736
rect 152 3704 192 3736
rect 224 3704 264 3736
rect 296 3704 336 3736
rect 368 3704 408 3736
rect 440 3704 480 3736
rect 512 3704 552 3736
rect 584 3704 624 3736
rect 656 3704 696 3736
rect 728 3704 768 3736
rect 800 3704 840 3736
rect 872 3704 912 3736
rect 944 3704 984 3736
rect 1016 3704 1056 3736
rect 1088 3704 1128 3736
rect 1160 3704 1200 3736
rect 1232 3704 1272 3736
rect 1304 3704 1344 3736
rect 1376 3704 1416 3736
rect 1448 3704 1488 3736
rect 1520 3704 1560 3736
rect 1592 3704 1632 3736
rect 1664 3704 1704 3736
rect 1736 3704 1776 3736
rect 1808 3704 1848 3736
rect 1880 3704 1920 3736
rect 1952 3704 2000 3736
rect 0 3664 2000 3704
rect 0 3632 48 3664
rect 80 3632 120 3664
rect 152 3632 192 3664
rect 224 3632 264 3664
rect 296 3632 336 3664
rect 368 3632 408 3664
rect 440 3632 480 3664
rect 512 3632 552 3664
rect 584 3632 624 3664
rect 656 3632 696 3664
rect 728 3632 768 3664
rect 800 3632 840 3664
rect 872 3632 912 3664
rect 944 3632 984 3664
rect 1016 3632 1056 3664
rect 1088 3632 1128 3664
rect 1160 3632 1200 3664
rect 1232 3632 1272 3664
rect 1304 3632 1344 3664
rect 1376 3632 1416 3664
rect 1448 3632 1488 3664
rect 1520 3632 1560 3664
rect 1592 3632 1632 3664
rect 1664 3632 1704 3664
rect 1736 3632 1776 3664
rect 1808 3632 1848 3664
rect 1880 3632 1920 3664
rect 1952 3632 2000 3664
rect 0 3592 2000 3632
rect 0 3560 48 3592
rect 80 3560 120 3592
rect 152 3560 192 3592
rect 224 3560 264 3592
rect 296 3560 336 3592
rect 368 3560 408 3592
rect 440 3560 480 3592
rect 512 3560 552 3592
rect 584 3560 624 3592
rect 656 3560 696 3592
rect 728 3560 768 3592
rect 800 3560 840 3592
rect 872 3560 912 3592
rect 944 3560 984 3592
rect 1016 3560 1056 3592
rect 1088 3560 1128 3592
rect 1160 3560 1200 3592
rect 1232 3560 1272 3592
rect 1304 3560 1344 3592
rect 1376 3560 1416 3592
rect 1448 3560 1488 3592
rect 1520 3560 1560 3592
rect 1592 3560 1632 3592
rect 1664 3560 1704 3592
rect 1736 3560 1776 3592
rect 1808 3560 1848 3592
rect 1880 3560 1920 3592
rect 1952 3560 2000 3592
rect 0 3520 2000 3560
rect 0 3488 48 3520
rect 80 3488 120 3520
rect 152 3488 192 3520
rect 224 3488 264 3520
rect 296 3488 336 3520
rect 368 3488 408 3520
rect 440 3488 480 3520
rect 512 3488 552 3520
rect 584 3488 624 3520
rect 656 3488 696 3520
rect 728 3488 768 3520
rect 800 3488 840 3520
rect 872 3488 912 3520
rect 944 3488 984 3520
rect 1016 3488 1056 3520
rect 1088 3488 1128 3520
rect 1160 3488 1200 3520
rect 1232 3488 1272 3520
rect 1304 3488 1344 3520
rect 1376 3488 1416 3520
rect 1448 3488 1488 3520
rect 1520 3488 1560 3520
rect 1592 3488 1632 3520
rect 1664 3488 1704 3520
rect 1736 3488 1776 3520
rect 1808 3488 1848 3520
rect 1880 3488 1920 3520
rect 1952 3488 2000 3520
rect 0 3448 2000 3488
rect 0 3416 48 3448
rect 80 3416 120 3448
rect 152 3416 192 3448
rect 224 3416 264 3448
rect 296 3416 336 3448
rect 368 3416 408 3448
rect 440 3416 480 3448
rect 512 3416 552 3448
rect 584 3416 624 3448
rect 656 3416 696 3448
rect 728 3416 768 3448
rect 800 3416 840 3448
rect 872 3416 912 3448
rect 944 3416 984 3448
rect 1016 3416 1056 3448
rect 1088 3416 1128 3448
rect 1160 3416 1200 3448
rect 1232 3416 1272 3448
rect 1304 3416 1344 3448
rect 1376 3416 1416 3448
rect 1448 3416 1488 3448
rect 1520 3416 1560 3448
rect 1592 3416 1632 3448
rect 1664 3416 1704 3448
rect 1736 3416 1776 3448
rect 1808 3416 1848 3448
rect 1880 3416 1920 3448
rect 1952 3416 2000 3448
rect 0 3376 2000 3416
rect 0 3344 48 3376
rect 80 3344 120 3376
rect 152 3344 192 3376
rect 224 3344 264 3376
rect 296 3344 336 3376
rect 368 3344 408 3376
rect 440 3344 480 3376
rect 512 3344 552 3376
rect 584 3344 624 3376
rect 656 3344 696 3376
rect 728 3344 768 3376
rect 800 3344 840 3376
rect 872 3344 912 3376
rect 944 3344 984 3376
rect 1016 3344 1056 3376
rect 1088 3344 1128 3376
rect 1160 3344 1200 3376
rect 1232 3344 1272 3376
rect 1304 3344 1344 3376
rect 1376 3344 1416 3376
rect 1448 3344 1488 3376
rect 1520 3344 1560 3376
rect 1592 3344 1632 3376
rect 1664 3344 1704 3376
rect 1736 3344 1776 3376
rect 1808 3344 1848 3376
rect 1880 3344 1920 3376
rect 1952 3344 2000 3376
rect 0 3304 2000 3344
rect 0 3272 48 3304
rect 80 3272 120 3304
rect 152 3272 192 3304
rect 224 3272 264 3304
rect 296 3272 336 3304
rect 368 3272 408 3304
rect 440 3272 480 3304
rect 512 3272 552 3304
rect 584 3272 624 3304
rect 656 3272 696 3304
rect 728 3272 768 3304
rect 800 3272 840 3304
rect 872 3272 912 3304
rect 944 3272 984 3304
rect 1016 3272 1056 3304
rect 1088 3272 1128 3304
rect 1160 3272 1200 3304
rect 1232 3272 1272 3304
rect 1304 3272 1344 3304
rect 1376 3272 1416 3304
rect 1448 3272 1488 3304
rect 1520 3272 1560 3304
rect 1592 3272 1632 3304
rect 1664 3272 1704 3304
rect 1736 3272 1776 3304
rect 1808 3272 1848 3304
rect 1880 3272 1920 3304
rect 1952 3272 2000 3304
rect 0 3232 2000 3272
rect 0 3200 48 3232
rect 80 3200 120 3232
rect 152 3200 192 3232
rect 224 3200 264 3232
rect 296 3200 336 3232
rect 368 3200 408 3232
rect 440 3200 480 3232
rect 512 3200 552 3232
rect 584 3200 624 3232
rect 656 3200 696 3232
rect 728 3200 768 3232
rect 800 3200 840 3232
rect 872 3200 912 3232
rect 944 3200 984 3232
rect 1016 3200 1056 3232
rect 1088 3200 1128 3232
rect 1160 3200 1200 3232
rect 1232 3200 1272 3232
rect 1304 3200 1344 3232
rect 1376 3200 1416 3232
rect 1448 3200 1488 3232
rect 1520 3200 1560 3232
rect 1592 3200 1632 3232
rect 1664 3200 1704 3232
rect 1736 3200 1776 3232
rect 1808 3200 1848 3232
rect 1880 3200 1920 3232
rect 1952 3200 2000 3232
rect 0 3160 2000 3200
rect 0 3128 48 3160
rect 80 3128 120 3160
rect 152 3128 192 3160
rect 224 3128 264 3160
rect 296 3128 336 3160
rect 368 3128 408 3160
rect 440 3128 480 3160
rect 512 3128 552 3160
rect 584 3128 624 3160
rect 656 3128 696 3160
rect 728 3128 768 3160
rect 800 3128 840 3160
rect 872 3128 912 3160
rect 944 3128 984 3160
rect 1016 3128 1056 3160
rect 1088 3128 1128 3160
rect 1160 3128 1200 3160
rect 1232 3128 1272 3160
rect 1304 3128 1344 3160
rect 1376 3128 1416 3160
rect 1448 3128 1488 3160
rect 1520 3128 1560 3160
rect 1592 3128 1632 3160
rect 1664 3128 1704 3160
rect 1736 3128 1776 3160
rect 1808 3128 1848 3160
rect 1880 3128 1920 3160
rect 1952 3128 2000 3160
rect 0 3088 2000 3128
rect 0 3056 48 3088
rect 80 3056 120 3088
rect 152 3056 192 3088
rect 224 3056 264 3088
rect 296 3056 336 3088
rect 368 3056 408 3088
rect 440 3056 480 3088
rect 512 3056 552 3088
rect 584 3056 624 3088
rect 656 3056 696 3088
rect 728 3056 768 3088
rect 800 3056 840 3088
rect 872 3056 912 3088
rect 944 3056 984 3088
rect 1016 3056 1056 3088
rect 1088 3056 1128 3088
rect 1160 3056 1200 3088
rect 1232 3056 1272 3088
rect 1304 3056 1344 3088
rect 1376 3056 1416 3088
rect 1448 3056 1488 3088
rect 1520 3056 1560 3088
rect 1592 3056 1632 3088
rect 1664 3056 1704 3088
rect 1736 3056 1776 3088
rect 1808 3056 1848 3088
rect 1880 3056 1920 3088
rect 1952 3056 2000 3088
rect 0 3016 2000 3056
rect 0 2984 48 3016
rect 80 2984 120 3016
rect 152 2984 192 3016
rect 224 2984 264 3016
rect 296 2984 336 3016
rect 368 2984 408 3016
rect 440 2984 480 3016
rect 512 2984 552 3016
rect 584 2984 624 3016
rect 656 2984 696 3016
rect 728 2984 768 3016
rect 800 2984 840 3016
rect 872 2984 912 3016
rect 944 2984 984 3016
rect 1016 2984 1056 3016
rect 1088 2984 1128 3016
rect 1160 2984 1200 3016
rect 1232 2984 1272 3016
rect 1304 2984 1344 3016
rect 1376 2984 1416 3016
rect 1448 2984 1488 3016
rect 1520 2984 1560 3016
rect 1592 2984 1632 3016
rect 1664 2984 1704 3016
rect 1736 2984 1776 3016
rect 1808 2984 1848 3016
rect 1880 2984 1920 3016
rect 1952 2984 2000 3016
rect 0 2944 2000 2984
rect 0 2912 48 2944
rect 80 2912 120 2944
rect 152 2912 192 2944
rect 224 2912 264 2944
rect 296 2912 336 2944
rect 368 2912 408 2944
rect 440 2912 480 2944
rect 512 2912 552 2944
rect 584 2912 624 2944
rect 656 2912 696 2944
rect 728 2912 768 2944
rect 800 2912 840 2944
rect 872 2912 912 2944
rect 944 2912 984 2944
rect 1016 2912 1056 2944
rect 1088 2912 1128 2944
rect 1160 2912 1200 2944
rect 1232 2912 1272 2944
rect 1304 2912 1344 2944
rect 1376 2912 1416 2944
rect 1448 2912 1488 2944
rect 1520 2912 1560 2944
rect 1592 2912 1632 2944
rect 1664 2912 1704 2944
rect 1736 2912 1776 2944
rect 1808 2912 1848 2944
rect 1880 2912 1920 2944
rect 1952 2912 2000 2944
rect 0 2872 2000 2912
rect 0 2840 48 2872
rect 80 2840 120 2872
rect 152 2840 192 2872
rect 224 2840 264 2872
rect 296 2840 336 2872
rect 368 2840 408 2872
rect 440 2840 480 2872
rect 512 2840 552 2872
rect 584 2840 624 2872
rect 656 2840 696 2872
rect 728 2840 768 2872
rect 800 2840 840 2872
rect 872 2840 912 2872
rect 944 2840 984 2872
rect 1016 2840 1056 2872
rect 1088 2840 1128 2872
rect 1160 2840 1200 2872
rect 1232 2840 1272 2872
rect 1304 2840 1344 2872
rect 1376 2840 1416 2872
rect 1448 2840 1488 2872
rect 1520 2840 1560 2872
rect 1592 2840 1632 2872
rect 1664 2840 1704 2872
rect 1736 2840 1776 2872
rect 1808 2840 1848 2872
rect 1880 2840 1920 2872
rect 1952 2840 2000 2872
rect 0 2800 2000 2840
rect 0 2768 48 2800
rect 80 2768 120 2800
rect 152 2768 192 2800
rect 224 2768 264 2800
rect 296 2768 336 2800
rect 368 2768 408 2800
rect 440 2768 480 2800
rect 512 2768 552 2800
rect 584 2768 624 2800
rect 656 2768 696 2800
rect 728 2768 768 2800
rect 800 2768 840 2800
rect 872 2768 912 2800
rect 944 2768 984 2800
rect 1016 2768 1056 2800
rect 1088 2768 1128 2800
rect 1160 2768 1200 2800
rect 1232 2768 1272 2800
rect 1304 2768 1344 2800
rect 1376 2768 1416 2800
rect 1448 2768 1488 2800
rect 1520 2768 1560 2800
rect 1592 2768 1632 2800
rect 1664 2768 1704 2800
rect 1736 2768 1776 2800
rect 1808 2768 1848 2800
rect 1880 2768 1920 2800
rect 1952 2768 2000 2800
rect 0 2728 2000 2768
rect 0 2696 48 2728
rect 80 2696 120 2728
rect 152 2696 192 2728
rect 224 2696 264 2728
rect 296 2696 336 2728
rect 368 2696 408 2728
rect 440 2696 480 2728
rect 512 2696 552 2728
rect 584 2696 624 2728
rect 656 2696 696 2728
rect 728 2696 768 2728
rect 800 2696 840 2728
rect 872 2696 912 2728
rect 944 2696 984 2728
rect 1016 2696 1056 2728
rect 1088 2696 1128 2728
rect 1160 2696 1200 2728
rect 1232 2696 1272 2728
rect 1304 2696 1344 2728
rect 1376 2696 1416 2728
rect 1448 2696 1488 2728
rect 1520 2696 1560 2728
rect 1592 2696 1632 2728
rect 1664 2696 1704 2728
rect 1736 2696 1776 2728
rect 1808 2696 1848 2728
rect 1880 2696 1920 2728
rect 1952 2696 2000 2728
rect 0 2656 2000 2696
rect 0 2624 48 2656
rect 80 2624 120 2656
rect 152 2624 192 2656
rect 224 2624 264 2656
rect 296 2624 336 2656
rect 368 2624 408 2656
rect 440 2624 480 2656
rect 512 2624 552 2656
rect 584 2624 624 2656
rect 656 2624 696 2656
rect 728 2624 768 2656
rect 800 2624 840 2656
rect 872 2624 912 2656
rect 944 2624 984 2656
rect 1016 2624 1056 2656
rect 1088 2624 1128 2656
rect 1160 2624 1200 2656
rect 1232 2624 1272 2656
rect 1304 2624 1344 2656
rect 1376 2624 1416 2656
rect 1448 2624 1488 2656
rect 1520 2624 1560 2656
rect 1592 2624 1632 2656
rect 1664 2624 1704 2656
rect 1736 2624 1776 2656
rect 1808 2624 1848 2656
rect 1880 2624 1920 2656
rect 1952 2624 2000 2656
rect 0 2584 2000 2624
rect 0 2552 48 2584
rect 80 2552 120 2584
rect 152 2552 192 2584
rect 224 2552 264 2584
rect 296 2552 336 2584
rect 368 2552 408 2584
rect 440 2552 480 2584
rect 512 2552 552 2584
rect 584 2552 624 2584
rect 656 2552 696 2584
rect 728 2552 768 2584
rect 800 2552 840 2584
rect 872 2552 912 2584
rect 944 2552 984 2584
rect 1016 2552 1056 2584
rect 1088 2552 1128 2584
rect 1160 2552 1200 2584
rect 1232 2552 1272 2584
rect 1304 2552 1344 2584
rect 1376 2552 1416 2584
rect 1448 2552 1488 2584
rect 1520 2552 1560 2584
rect 1592 2552 1632 2584
rect 1664 2552 1704 2584
rect 1736 2552 1776 2584
rect 1808 2552 1848 2584
rect 1880 2552 1920 2584
rect 1952 2552 2000 2584
rect 0 2512 2000 2552
rect 0 2480 48 2512
rect 80 2480 120 2512
rect 152 2480 192 2512
rect 224 2480 264 2512
rect 296 2480 336 2512
rect 368 2480 408 2512
rect 440 2480 480 2512
rect 512 2480 552 2512
rect 584 2480 624 2512
rect 656 2480 696 2512
rect 728 2480 768 2512
rect 800 2480 840 2512
rect 872 2480 912 2512
rect 944 2480 984 2512
rect 1016 2480 1056 2512
rect 1088 2480 1128 2512
rect 1160 2480 1200 2512
rect 1232 2480 1272 2512
rect 1304 2480 1344 2512
rect 1376 2480 1416 2512
rect 1448 2480 1488 2512
rect 1520 2480 1560 2512
rect 1592 2480 1632 2512
rect 1664 2480 1704 2512
rect 1736 2480 1776 2512
rect 1808 2480 1848 2512
rect 1880 2480 1920 2512
rect 1952 2480 2000 2512
rect 0 2440 2000 2480
rect 0 2408 48 2440
rect 80 2408 120 2440
rect 152 2408 192 2440
rect 224 2408 264 2440
rect 296 2408 336 2440
rect 368 2408 408 2440
rect 440 2408 480 2440
rect 512 2408 552 2440
rect 584 2408 624 2440
rect 656 2408 696 2440
rect 728 2408 768 2440
rect 800 2408 840 2440
rect 872 2408 912 2440
rect 944 2408 984 2440
rect 1016 2408 1056 2440
rect 1088 2408 1128 2440
rect 1160 2408 1200 2440
rect 1232 2408 1272 2440
rect 1304 2408 1344 2440
rect 1376 2408 1416 2440
rect 1448 2408 1488 2440
rect 1520 2408 1560 2440
rect 1592 2408 1632 2440
rect 1664 2408 1704 2440
rect 1736 2408 1776 2440
rect 1808 2408 1848 2440
rect 1880 2408 1920 2440
rect 1952 2408 2000 2440
rect 0 2368 2000 2408
rect 0 2336 48 2368
rect 80 2336 120 2368
rect 152 2336 192 2368
rect 224 2336 264 2368
rect 296 2336 336 2368
rect 368 2336 408 2368
rect 440 2336 480 2368
rect 512 2336 552 2368
rect 584 2336 624 2368
rect 656 2336 696 2368
rect 728 2336 768 2368
rect 800 2336 840 2368
rect 872 2336 912 2368
rect 944 2336 984 2368
rect 1016 2336 1056 2368
rect 1088 2336 1128 2368
rect 1160 2336 1200 2368
rect 1232 2336 1272 2368
rect 1304 2336 1344 2368
rect 1376 2336 1416 2368
rect 1448 2336 1488 2368
rect 1520 2336 1560 2368
rect 1592 2336 1632 2368
rect 1664 2336 1704 2368
rect 1736 2336 1776 2368
rect 1808 2336 1848 2368
rect 1880 2336 1920 2368
rect 1952 2336 2000 2368
rect 0 2296 2000 2336
rect 0 2264 48 2296
rect 80 2264 120 2296
rect 152 2264 192 2296
rect 224 2264 264 2296
rect 296 2264 336 2296
rect 368 2264 408 2296
rect 440 2264 480 2296
rect 512 2264 552 2296
rect 584 2264 624 2296
rect 656 2264 696 2296
rect 728 2264 768 2296
rect 800 2264 840 2296
rect 872 2264 912 2296
rect 944 2264 984 2296
rect 1016 2264 1056 2296
rect 1088 2264 1128 2296
rect 1160 2264 1200 2296
rect 1232 2264 1272 2296
rect 1304 2264 1344 2296
rect 1376 2264 1416 2296
rect 1448 2264 1488 2296
rect 1520 2264 1560 2296
rect 1592 2264 1632 2296
rect 1664 2264 1704 2296
rect 1736 2264 1776 2296
rect 1808 2264 1848 2296
rect 1880 2264 1920 2296
rect 1952 2264 2000 2296
rect 0 2224 2000 2264
rect 0 2192 48 2224
rect 80 2192 120 2224
rect 152 2192 192 2224
rect 224 2192 264 2224
rect 296 2192 336 2224
rect 368 2192 408 2224
rect 440 2192 480 2224
rect 512 2192 552 2224
rect 584 2192 624 2224
rect 656 2192 696 2224
rect 728 2192 768 2224
rect 800 2192 840 2224
rect 872 2192 912 2224
rect 944 2192 984 2224
rect 1016 2192 1056 2224
rect 1088 2192 1128 2224
rect 1160 2192 1200 2224
rect 1232 2192 1272 2224
rect 1304 2192 1344 2224
rect 1376 2192 1416 2224
rect 1448 2192 1488 2224
rect 1520 2192 1560 2224
rect 1592 2192 1632 2224
rect 1664 2192 1704 2224
rect 1736 2192 1776 2224
rect 1808 2192 1848 2224
rect 1880 2192 1920 2224
rect 1952 2192 2000 2224
rect 0 2152 2000 2192
rect 0 2120 48 2152
rect 80 2120 120 2152
rect 152 2120 192 2152
rect 224 2120 264 2152
rect 296 2120 336 2152
rect 368 2120 408 2152
rect 440 2120 480 2152
rect 512 2120 552 2152
rect 584 2120 624 2152
rect 656 2120 696 2152
rect 728 2120 768 2152
rect 800 2120 840 2152
rect 872 2120 912 2152
rect 944 2120 984 2152
rect 1016 2120 1056 2152
rect 1088 2120 1128 2152
rect 1160 2120 1200 2152
rect 1232 2120 1272 2152
rect 1304 2120 1344 2152
rect 1376 2120 1416 2152
rect 1448 2120 1488 2152
rect 1520 2120 1560 2152
rect 1592 2120 1632 2152
rect 1664 2120 1704 2152
rect 1736 2120 1776 2152
rect 1808 2120 1848 2152
rect 1880 2120 1920 2152
rect 1952 2120 2000 2152
rect 0 2080 2000 2120
rect 0 2048 48 2080
rect 80 2048 120 2080
rect 152 2048 192 2080
rect 224 2048 264 2080
rect 296 2048 336 2080
rect 368 2048 408 2080
rect 440 2048 480 2080
rect 512 2048 552 2080
rect 584 2048 624 2080
rect 656 2048 696 2080
rect 728 2048 768 2080
rect 800 2048 840 2080
rect 872 2048 912 2080
rect 944 2048 984 2080
rect 1016 2048 1056 2080
rect 1088 2048 1128 2080
rect 1160 2048 1200 2080
rect 1232 2048 1272 2080
rect 1304 2048 1344 2080
rect 1376 2048 1416 2080
rect 1448 2048 1488 2080
rect 1520 2048 1560 2080
rect 1592 2048 1632 2080
rect 1664 2048 1704 2080
rect 1736 2048 1776 2080
rect 1808 2048 1848 2080
rect 1880 2048 1920 2080
rect 1952 2048 2000 2080
rect 0 2008 2000 2048
rect 0 1976 48 2008
rect 80 1976 120 2008
rect 152 1976 192 2008
rect 224 1976 264 2008
rect 296 1976 336 2008
rect 368 1976 408 2008
rect 440 1976 480 2008
rect 512 1976 552 2008
rect 584 1976 624 2008
rect 656 1976 696 2008
rect 728 1976 768 2008
rect 800 1976 840 2008
rect 872 1976 912 2008
rect 944 1976 984 2008
rect 1016 1976 1056 2008
rect 1088 1976 1128 2008
rect 1160 1976 1200 2008
rect 1232 1976 1272 2008
rect 1304 1976 1344 2008
rect 1376 1976 1416 2008
rect 1448 1976 1488 2008
rect 1520 1976 1560 2008
rect 1592 1976 1632 2008
rect 1664 1976 1704 2008
rect 1736 1976 1776 2008
rect 1808 1976 1848 2008
rect 1880 1976 1920 2008
rect 1952 1976 2000 2008
rect 0 1936 2000 1976
rect 0 1904 48 1936
rect 80 1904 120 1936
rect 152 1904 192 1936
rect 224 1904 264 1936
rect 296 1904 336 1936
rect 368 1904 408 1936
rect 440 1904 480 1936
rect 512 1904 552 1936
rect 584 1904 624 1936
rect 656 1904 696 1936
rect 728 1904 768 1936
rect 800 1904 840 1936
rect 872 1904 912 1936
rect 944 1904 984 1936
rect 1016 1904 1056 1936
rect 1088 1904 1128 1936
rect 1160 1904 1200 1936
rect 1232 1904 1272 1936
rect 1304 1904 1344 1936
rect 1376 1904 1416 1936
rect 1448 1904 1488 1936
rect 1520 1904 1560 1936
rect 1592 1904 1632 1936
rect 1664 1904 1704 1936
rect 1736 1904 1776 1936
rect 1808 1904 1848 1936
rect 1880 1904 1920 1936
rect 1952 1904 2000 1936
rect 0 1864 2000 1904
rect 0 1832 48 1864
rect 80 1832 120 1864
rect 152 1832 192 1864
rect 224 1832 264 1864
rect 296 1832 336 1864
rect 368 1832 408 1864
rect 440 1832 480 1864
rect 512 1832 552 1864
rect 584 1832 624 1864
rect 656 1832 696 1864
rect 728 1832 768 1864
rect 800 1832 840 1864
rect 872 1832 912 1864
rect 944 1832 984 1864
rect 1016 1832 1056 1864
rect 1088 1832 1128 1864
rect 1160 1832 1200 1864
rect 1232 1832 1272 1864
rect 1304 1832 1344 1864
rect 1376 1832 1416 1864
rect 1448 1832 1488 1864
rect 1520 1832 1560 1864
rect 1592 1832 1632 1864
rect 1664 1832 1704 1864
rect 1736 1832 1776 1864
rect 1808 1832 1848 1864
rect 1880 1832 1920 1864
rect 1952 1832 2000 1864
rect 0 1792 2000 1832
rect 0 1760 48 1792
rect 80 1760 120 1792
rect 152 1760 192 1792
rect 224 1760 264 1792
rect 296 1760 336 1792
rect 368 1760 408 1792
rect 440 1760 480 1792
rect 512 1760 552 1792
rect 584 1760 624 1792
rect 656 1760 696 1792
rect 728 1760 768 1792
rect 800 1760 840 1792
rect 872 1760 912 1792
rect 944 1760 984 1792
rect 1016 1760 1056 1792
rect 1088 1760 1128 1792
rect 1160 1760 1200 1792
rect 1232 1760 1272 1792
rect 1304 1760 1344 1792
rect 1376 1760 1416 1792
rect 1448 1760 1488 1792
rect 1520 1760 1560 1792
rect 1592 1760 1632 1792
rect 1664 1760 1704 1792
rect 1736 1760 1776 1792
rect 1808 1760 1848 1792
rect 1880 1760 1920 1792
rect 1952 1760 2000 1792
rect 0 1720 2000 1760
rect 0 1688 48 1720
rect 80 1688 120 1720
rect 152 1688 192 1720
rect 224 1688 264 1720
rect 296 1688 336 1720
rect 368 1688 408 1720
rect 440 1688 480 1720
rect 512 1688 552 1720
rect 584 1688 624 1720
rect 656 1688 696 1720
rect 728 1688 768 1720
rect 800 1688 840 1720
rect 872 1688 912 1720
rect 944 1688 984 1720
rect 1016 1688 1056 1720
rect 1088 1688 1128 1720
rect 1160 1688 1200 1720
rect 1232 1688 1272 1720
rect 1304 1688 1344 1720
rect 1376 1688 1416 1720
rect 1448 1688 1488 1720
rect 1520 1688 1560 1720
rect 1592 1688 1632 1720
rect 1664 1688 1704 1720
rect 1736 1688 1776 1720
rect 1808 1688 1848 1720
rect 1880 1688 1920 1720
rect 1952 1688 2000 1720
rect 0 1648 2000 1688
rect 0 1616 48 1648
rect 80 1616 120 1648
rect 152 1616 192 1648
rect 224 1616 264 1648
rect 296 1616 336 1648
rect 368 1616 408 1648
rect 440 1616 480 1648
rect 512 1616 552 1648
rect 584 1616 624 1648
rect 656 1616 696 1648
rect 728 1616 768 1648
rect 800 1616 840 1648
rect 872 1616 912 1648
rect 944 1616 984 1648
rect 1016 1616 1056 1648
rect 1088 1616 1128 1648
rect 1160 1616 1200 1648
rect 1232 1616 1272 1648
rect 1304 1616 1344 1648
rect 1376 1616 1416 1648
rect 1448 1616 1488 1648
rect 1520 1616 1560 1648
rect 1592 1616 1632 1648
rect 1664 1616 1704 1648
rect 1736 1616 1776 1648
rect 1808 1616 1848 1648
rect 1880 1616 1920 1648
rect 1952 1616 2000 1648
rect 0 1576 2000 1616
rect 0 1544 48 1576
rect 80 1544 120 1576
rect 152 1544 192 1576
rect 224 1544 264 1576
rect 296 1544 336 1576
rect 368 1544 408 1576
rect 440 1544 480 1576
rect 512 1544 552 1576
rect 584 1544 624 1576
rect 656 1544 696 1576
rect 728 1544 768 1576
rect 800 1544 840 1576
rect 872 1544 912 1576
rect 944 1544 984 1576
rect 1016 1544 1056 1576
rect 1088 1544 1128 1576
rect 1160 1544 1200 1576
rect 1232 1544 1272 1576
rect 1304 1544 1344 1576
rect 1376 1544 1416 1576
rect 1448 1544 1488 1576
rect 1520 1544 1560 1576
rect 1592 1544 1632 1576
rect 1664 1544 1704 1576
rect 1736 1544 1776 1576
rect 1808 1544 1848 1576
rect 1880 1544 1920 1576
rect 1952 1544 2000 1576
rect 0 1504 2000 1544
rect 0 1472 48 1504
rect 80 1472 120 1504
rect 152 1472 192 1504
rect 224 1472 264 1504
rect 296 1472 336 1504
rect 368 1472 408 1504
rect 440 1472 480 1504
rect 512 1472 552 1504
rect 584 1472 624 1504
rect 656 1472 696 1504
rect 728 1472 768 1504
rect 800 1472 840 1504
rect 872 1472 912 1504
rect 944 1472 984 1504
rect 1016 1472 1056 1504
rect 1088 1472 1128 1504
rect 1160 1472 1200 1504
rect 1232 1472 1272 1504
rect 1304 1472 1344 1504
rect 1376 1472 1416 1504
rect 1448 1472 1488 1504
rect 1520 1472 1560 1504
rect 1592 1472 1632 1504
rect 1664 1472 1704 1504
rect 1736 1472 1776 1504
rect 1808 1472 1848 1504
rect 1880 1472 1920 1504
rect 1952 1472 2000 1504
rect 0 1432 2000 1472
rect 0 1400 48 1432
rect 80 1400 120 1432
rect 152 1400 192 1432
rect 224 1400 264 1432
rect 296 1400 336 1432
rect 368 1400 408 1432
rect 440 1400 480 1432
rect 512 1400 552 1432
rect 584 1400 624 1432
rect 656 1400 696 1432
rect 728 1400 768 1432
rect 800 1400 840 1432
rect 872 1400 912 1432
rect 944 1400 984 1432
rect 1016 1400 1056 1432
rect 1088 1400 1128 1432
rect 1160 1400 1200 1432
rect 1232 1400 1272 1432
rect 1304 1400 1344 1432
rect 1376 1400 1416 1432
rect 1448 1400 1488 1432
rect 1520 1400 1560 1432
rect 1592 1400 1632 1432
rect 1664 1400 1704 1432
rect 1736 1400 1776 1432
rect 1808 1400 1848 1432
rect 1880 1400 1920 1432
rect 1952 1400 2000 1432
rect 0 1360 2000 1400
rect 0 1328 48 1360
rect 80 1328 120 1360
rect 152 1328 192 1360
rect 224 1328 264 1360
rect 296 1328 336 1360
rect 368 1328 408 1360
rect 440 1328 480 1360
rect 512 1328 552 1360
rect 584 1328 624 1360
rect 656 1328 696 1360
rect 728 1328 768 1360
rect 800 1328 840 1360
rect 872 1328 912 1360
rect 944 1328 984 1360
rect 1016 1328 1056 1360
rect 1088 1328 1128 1360
rect 1160 1328 1200 1360
rect 1232 1328 1272 1360
rect 1304 1328 1344 1360
rect 1376 1328 1416 1360
rect 1448 1328 1488 1360
rect 1520 1328 1560 1360
rect 1592 1328 1632 1360
rect 1664 1328 1704 1360
rect 1736 1328 1776 1360
rect 1808 1328 1848 1360
rect 1880 1328 1920 1360
rect 1952 1328 2000 1360
rect 0 1288 2000 1328
rect 0 1256 48 1288
rect 80 1256 120 1288
rect 152 1256 192 1288
rect 224 1256 264 1288
rect 296 1256 336 1288
rect 368 1256 408 1288
rect 440 1256 480 1288
rect 512 1256 552 1288
rect 584 1256 624 1288
rect 656 1256 696 1288
rect 728 1256 768 1288
rect 800 1256 840 1288
rect 872 1256 912 1288
rect 944 1256 984 1288
rect 1016 1256 1056 1288
rect 1088 1256 1128 1288
rect 1160 1256 1200 1288
rect 1232 1256 1272 1288
rect 1304 1256 1344 1288
rect 1376 1256 1416 1288
rect 1448 1256 1488 1288
rect 1520 1256 1560 1288
rect 1592 1256 1632 1288
rect 1664 1256 1704 1288
rect 1736 1256 1776 1288
rect 1808 1256 1848 1288
rect 1880 1256 1920 1288
rect 1952 1256 2000 1288
rect 0 1200 2000 1256
<< psubdiffcont >>
rect 699 31384 731 31416
rect 120 27939 152 27971
rect 120 22842 152 22874
rect 120 17816 152 17848
<< nsubdiffcont >>
rect 120 33384 152 33416
rect 120 29684 152 29716
rect 48 12112 80 12144
rect 48 6512 80 6544
<< metal1 >>
rect 192 33384 224 33416
rect 264 33384 296 33416
rect 336 33384 368 33416
rect 408 33384 440 33416
rect 480 33384 512 33416
rect 552 33384 584 33416
rect 624 33384 656 33416
rect 696 33384 728 33416
rect 768 33384 800 33416
rect 840 33384 872 33416
rect 912 33384 944 33416
rect 984 33384 1016 33416
rect 1056 33384 1088 33416
rect 1128 33384 1160 33416
rect 1200 33384 1232 33416
rect 1272 33384 1304 33416
rect 1344 33384 1376 33416
rect 1416 33384 1448 33416
rect 1488 33384 1520 33416
rect 1560 33384 1592 33416
rect 1632 33384 1664 33416
rect 1704 33384 1736 33416
rect 1776 33384 1808 33416
rect 1848 33384 1880 33416
rect 192 29684 224 29716
rect 264 29684 296 29716
rect 336 29684 368 29716
rect 408 29684 440 29716
rect 480 29684 512 29716
rect 552 29684 584 29716
rect 624 29684 656 29716
rect 696 29684 728 29716
rect 768 29684 800 29716
rect 840 29684 872 29716
rect 912 29684 944 29716
rect 984 29684 1016 29716
rect 1056 29684 1088 29716
rect 1128 29684 1160 29716
rect 1200 29684 1232 29716
rect 1272 29684 1304 29716
rect 1344 29684 1376 29716
rect 1416 29684 1448 29716
rect 1488 29684 1520 29716
rect 1560 29684 1592 29716
rect 1632 29684 1664 29716
rect 1704 29684 1736 29716
rect 1776 29684 1808 29716
rect 1848 29684 1880 29716
rect 120 12112 152 12144
rect 192 12112 224 12144
rect 264 12112 296 12144
rect 336 12112 368 12144
rect 408 12112 440 12144
rect 480 12112 512 12144
rect 552 12112 584 12144
rect 624 12112 656 12144
rect 696 12112 728 12144
rect 768 12112 800 12144
rect 840 12112 872 12144
rect 912 12112 944 12144
rect 984 12112 1016 12144
rect 1056 12112 1088 12144
rect 1128 12112 1160 12144
rect 1200 12112 1232 12144
rect 1272 12112 1304 12144
rect 1344 12112 1376 12144
rect 1416 12112 1448 12144
rect 1488 12112 1520 12144
rect 1560 12112 1592 12144
rect 1632 12112 1664 12144
rect 1704 12112 1736 12144
rect 1776 12112 1808 12144
rect 1848 12112 1880 12144
rect 1920 12112 1952 12144
rect 48 12040 80 12072
rect 120 12040 152 12072
rect 192 12040 224 12072
rect 264 12040 296 12072
rect 336 12040 368 12072
rect 408 12040 440 12072
rect 480 12040 512 12072
rect 552 12040 584 12072
rect 624 12040 656 12072
rect 696 12040 728 12072
rect 768 12040 800 12072
rect 840 12040 872 12072
rect 912 12040 944 12072
rect 984 12040 1016 12072
rect 1056 12040 1088 12072
rect 1128 12040 1160 12072
rect 1200 12040 1232 12072
rect 1272 12040 1304 12072
rect 1344 12040 1376 12072
rect 1416 12040 1448 12072
rect 1488 12040 1520 12072
rect 1560 12040 1592 12072
rect 1632 12040 1664 12072
rect 1704 12040 1736 12072
rect 1776 12040 1808 12072
rect 1848 12040 1880 12072
rect 1920 12040 1952 12072
rect 48 11968 80 12000
rect 120 11968 152 12000
rect 192 11968 224 12000
rect 264 11968 296 12000
rect 336 11968 368 12000
rect 408 11968 440 12000
rect 480 11968 512 12000
rect 552 11968 584 12000
rect 624 11968 656 12000
rect 696 11968 728 12000
rect 768 11968 800 12000
rect 840 11968 872 12000
rect 912 11968 944 12000
rect 984 11968 1016 12000
rect 1056 11968 1088 12000
rect 1128 11968 1160 12000
rect 1200 11968 1232 12000
rect 1272 11968 1304 12000
rect 1344 11968 1376 12000
rect 1416 11968 1448 12000
rect 1488 11968 1520 12000
rect 1560 11968 1592 12000
rect 1632 11968 1664 12000
rect 1704 11968 1736 12000
rect 1776 11968 1808 12000
rect 1848 11968 1880 12000
rect 1920 11968 1952 12000
rect 48 11896 80 11928
rect 120 11896 152 11928
rect 192 11896 224 11928
rect 264 11896 296 11928
rect 336 11896 368 11928
rect 408 11896 440 11928
rect 480 11896 512 11928
rect 552 11896 584 11928
rect 624 11896 656 11928
rect 696 11896 728 11928
rect 768 11896 800 11928
rect 840 11896 872 11928
rect 912 11896 944 11928
rect 984 11896 1016 11928
rect 1056 11896 1088 11928
rect 1128 11896 1160 11928
rect 1200 11896 1232 11928
rect 1272 11896 1304 11928
rect 1344 11896 1376 11928
rect 1416 11896 1448 11928
rect 1488 11896 1520 11928
rect 1560 11896 1592 11928
rect 1632 11896 1664 11928
rect 1704 11896 1736 11928
rect 1776 11896 1808 11928
rect 1848 11896 1880 11928
rect 1920 11896 1952 11928
rect 48 11824 80 11856
rect 120 11824 152 11856
rect 192 11824 224 11856
rect 264 11824 296 11856
rect 336 11824 368 11856
rect 408 11824 440 11856
rect 480 11824 512 11856
rect 552 11824 584 11856
rect 624 11824 656 11856
rect 696 11824 728 11856
rect 768 11824 800 11856
rect 840 11824 872 11856
rect 912 11824 944 11856
rect 984 11824 1016 11856
rect 1056 11824 1088 11856
rect 1128 11824 1160 11856
rect 1200 11824 1232 11856
rect 1272 11824 1304 11856
rect 1344 11824 1376 11856
rect 1416 11824 1448 11856
rect 1488 11824 1520 11856
rect 1560 11824 1592 11856
rect 1632 11824 1664 11856
rect 1704 11824 1736 11856
rect 1776 11824 1808 11856
rect 1848 11824 1880 11856
rect 1920 11824 1952 11856
rect 48 11752 80 11784
rect 120 11752 152 11784
rect 192 11752 224 11784
rect 264 11752 296 11784
rect 336 11752 368 11784
rect 408 11752 440 11784
rect 480 11752 512 11784
rect 552 11752 584 11784
rect 624 11752 656 11784
rect 696 11752 728 11784
rect 768 11752 800 11784
rect 840 11752 872 11784
rect 912 11752 944 11784
rect 984 11752 1016 11784
rect 1056 11752 1088 11784
rect 1128 11752 1160 11784
rect 1200 11752 1232 11784
rect 1272 11752 1304 11784
rect 1344 11752 1376 11784
rect 1416 11752 1448 11784
rect 1488 11752 1520 11784
rect 1560 11752 1592 11784
rect 1632 11752 1664 11784
rect 1704 11752 1736 11784
rect 1776 11752 1808 11784
rect 1848 11752 1880 11784
rect 1920 11752 1952 11784
rect 48 11680 80 11712
rect 120 11680 152 11712
rect 192 11680 224 11712
rect 264 11680 296 11712
rect 336 11680 368 11712
rect 408 11680 440 11712
rect 480 11680 512 11712
rect 552 11680 584 11712
rect 624 11680 656 11712
rect 696 11680 728 11712
rect 768 11680 800 11712
rect 840 11680 872 11712
rect 912 11680 944 11712
rect 984 11680 1016 11712
rect 1056 11680 1088 11712
rect 1128 11680 1160 11712
rect 1200 11680 1232 11712
rect 1272 11680 1304 11712
rect 1344 11680 1376 11712
rect 1416 11680 1448 11712
rect 1488 11680 1520 11712
rect 1560 11680 1592 11712
rect 1632 11680 1664 11712
rect 1704 11680 1736 11712
rect 1776 11680 1808 11712
rect 1848 11680 1880 11712
rect 1920 11680 1952 11712
rect 48 11608 80 11640
rect 120 11608 152 11640
rect 192 11608 224 11640
rect 264 11608 296 11640
rect 336 11608 368 11640
rect 408 11608 440 11640
rect 480 11608 512 11640
rect 552 11608 584 11640
rect 624 11608 656 11640
rect 696 11608 728 11640
rect 768 11608 800 11640
rect 840 11608 872 11640
rect 912 11608 944 11640
rect 984 11608 1016 11640
rect 1056 11608 1088 11640
rect 1128 11608 1160 11640
rect 1200 11608 1232 11640
rect 1272 11608 1304 11640
rect 1344 11608 1376 11640
rect 1416 11608 1448 11640
rect 1488 11608 1520 11640
rect 1560 11608 1592 11640
rect 1632 11608 1664 11640
rect 1704 11608 1736 11640
rect 1776 11608 1808 11640
rect 1848 11608 1880 11640
rect 1920 11608 1952 11640
rect 48 11536 80 11568
rect 120 11536 152 11568
rect 192 11536 224 11568
rect 264 11536 296 11568
rect 336 11536 368 11568
rect 408 11536 440 11568
rect 480 11536 512 11568
rect 552 11536 584 11568
rect 624 11536 656 11568
rect 696 11536 728 11568
rect 768 11536 800 11568
rect 840 11536 872 11568
rect 912 11536 944 11568
rect 984 11536 1016 11568
rect 1056 11536 1088 11568
rect 1128 11536 1160 11568
rect 1200 11536 1232 11568
rect 1272 11536 1304 11568
rect 1344 11536 1376 11568
rect 1416 11536 1448 11568
rect 1488 11536 1520 11568
rect 1560 11536 1592 11568
rect 1632 11536 1664 11568
rect 1704 11536 1736 11568
rect 1776 11536 1808 11568
rect 1848 11536 1880 11568
rect 1920 11536 1952 11568
rect 48 11464 80 11496
rect 120 11464 152 11496
rect 192 11464 224 11496
rect 264 11464 296 11496
rect 336 11464 368 11496
rect 408 11464 440 11496
rect 480 11464 512 11496
rect 552 11464 584 11496
rect 624 11464 656 11496
rect 696 11464 728 11496
rect 768 11464 800 11496
rect 840 11464 872 11496
rect 912 11464 944 11496
rect 984 11464 1016 11496
rect 1056 11464 1088 11496
rect 1128 11464 1160 11496
rect 1200 11464 1232 11496
rect 1272 11464 1304 11496
rect 1344 11464 1376 11496
rect 1416 11464 1448 11496
rect 1488 11464 1520 11496
rect 1560 11464 1592 11496
rect 1632 11464 1664 11496
rect 1704 11464 1736 11496
rect 1776 11464 1808 11496
rect 1848 11464 1880 11496
rect 1920 11464 1952 11496
rect 48 11392 80 11424
rect 120 11392 152 11424
rect 192 11392 224 11424
rect 264 11392 296 11424
rect 336 11392 368 11424
rect 408 11392 440 11424
rect 480 11392 512 11424
rect 552 11392 584 11424
rect 624 11392 656 11424
rect 696 11392 728 11424
rect 768 11392 800 11424
rect 840 11392 872 11424
rect 912 11392 944 11424
rect 984 11392 1016 11424
rect 1056 11392 1088 11424
rect 1128 11392 1160 11424
rect 1200 11392 1232 11424
rect 1272 11392 1304 11424
rect 1344 11392 1376 11424
rect 1416 11392 1448 11424
rect 1488 11392 1520 11424
rect 1560 11392 1592 11424
rect 1632 11392 1664 11424
rect 1704 11392 1736 11424
rect 1776 11392 1808 11424
rect 1848 11392 1880 11424
rect 1920 11392 1952 11424
rect 48 11320 80 11352
rect 120 11320 152 11352
rect 192 11320 224 11352
rect 264 11320 296 11352
rect 336 11320 368 11352
rect 408 11320 440 11352
rect 480 11320 512 11352
rect 552 11320 584 11352
rect 624 11320 656 11352
rect 696 11320 728 11352
rect 768 11320 800 11352
rect 840 11320 872 11352
rect 912 11320 944 11352
rect 984 11320 1016 11352
rect 1056 11320 1088 11352
rect 1128 11320 1160 11352
rect 1200 11320 1232 11352
rect 1272 11320 1304 11352
rect 1344 11320 1376 11352
rect 1416 11320 1448 11352
rect 1488 11320 1520 11352
rect 1560 11320 1592 11352
rect 1632 11320 1664 11352
rect 1704 11320 1736 11352
rect 1776 11320 1808 11352
rect 1848 11320 1880 11352
rect 1920 11320 1952 11352
rect 48 11248 80 11280
rect 120 11248 152 11280
rect 192 11248 224 11280
rect 264 11248 296 11280
rect 336 11248 368 11280
rect 408 11248 440 11280
rect 480 11248 512 11280
rect 552 11248 584 11280
rect 624 11248 656 11280
rect 696 11248 728 11280
rect 768 11248 800 11280
rect 840 11248 872 11280
rect 912 11248 944 11280
rect 984 11248 1016 11280
rect 1056 11248 1088 11280
rect 1128 11248 1160 11280
rect 1200 11248 1232 11280
rect 1272 11248 1304 11280
rect 1344 11248 1376 11280
rect 1416 11248 1448 11280
rect 1488 11248 1520 11280
rect 1560 11248 1592 11280
rect 1632 11248 1664 11280
rect 1704 11248 1736 11280
rect 1776 11248 1808 11280
rect 1848 11248 1880 11280
rect 1920 11248 1952 11280
rect 48 11176 80 11208
rect 120 11176 152 11208
rect 192 11176 224 11208
rect 264 11176 296 11208
rect 336 11176 368 11208
rect 408 11176 440 11208
rect 480 11176 512 11208
rect 552 11176 584 11208
rect 624 11176 656 11208
rect 696 11176 728 11208
rect 768 11176 800 11208
rect 840 11176 872 11208
rect 912 11176 944 11208
rect 984 11176 1016 11208
rect 1056 11176 1088 11208
rect 1128 11176 1160 11208
rect 1200 11176 1232 11208
rect 1272 11176 1304 11208
rect 1344 11176 1376 11208
rect 1416 11176 1448 11208
rect 1488 11176 1520 11208
rect 1560 11176 1592 11208
rect 1632 11176 1664 11208
rect 1704 11176 1736 11208
rect 1776 11176 1808 11208
rect 1848 11176 1880 11208
rect 1920 11176 1952 11208
rect 48 11104 80 11136
rect 120 11104 152 11136
rect 192 11104 224 11136
rect 264 11104 296 11136
rect 336 11104 368 11136
rect 408 11104 440 11136
rect 480 11104 512 11136
rect 552 11104 584 11136
rect 624 11104 656 11136
rect 696 11104 728 11136
rect 768 11104 800 11136
rect 840 11104 872 11136
rect 912 11104 944 11136
rect 984 11104 1016 11136
rect 1056 11104 1088 11136
rect 1128 11104 1160 11136
rect 1200 11104 1232 11136
rect 1272 11104 1304 11136
rect 1344 11104 1376 11136
rect 1416 11104 1448 11136
rect 1488 11104 1520 11136
rect 1560 11104 1592 11136
rect 1632 11104 1664 11136
rect 1704 11104 1736 11136
rect 1776 11104 1808 11136
rect 1848 11104 1880 11136
rect 1920 11104 1952 11136
rect 48 11032 80 11064
rect 120 11032 152 11064
rect 192 11032 224 11064
rect 264 11032 296 11064
rect 336 11032 368 11064
rect 408 11032 440 11064
rect 480 11032 512 11064
rect 552 11032 584 11064
rect 624 11032 656 11064
rect 696 11032 728 11064
rect 768 11032 800 11064
rect 840 11032 872 11064
rect 912 11032 944 11064
rect 984 11032 1016 11064
rect 1056 11032 1088 11064
rect 1128 11032 1160 11064
rect 1200 11032 1232 11064
rect 1272 11032 1304 11064
rect 1344 11032 1376 11064
rect 1416 11032 1448 11064
rect 1488 11032 1520 11064
rect 1560 11032 1592 11064
rect 1632 11032 1664 11064
rect 1704 11032 1736 11064
rect 1776 11032 1808 11064
rect 1848 11032 1880 11064
rect 1920 11032 1952 11064
rect 48 10960 80 10992
rect 120 10960 152 10992
rect 192 10960 224 10992
rect 264 10960 296 10992
rect 336 10960 368 10992
rect 408 10960 440 10992
rect 480 10960 512 10992
rect 552 10960 584 10992
rect 624 10960 656 10992
rect 696 10960 728 10992
rect 768 10960 800 10992
rect 840 10960 872 10992
rect 912 10960 944 10992
rect 984 10960 1016 10992
rect 1056 10960 1088 10992
rect 1128 10960 1160 10992
rect 1200 10960 1232 10992
rect 1272 10960 1304 10992
rect 1344 10960 1376 10992
rect 1416 10960 1448 10992
rect 1488 10960 1520 10992
rect 1560 10960 1592 10992
rect 1632 10960 1664 10992
rect 1704 10960 1736 10992
rect 1776 10960 1808 10992
rect 1848 10960 1880 10992
rect 1920 10960 1952 10992
rect 48 10888 80 10920
rect 120 10888 152 10920
rect 192 10888 224 10920
rect 264 10888 296 10920
rect 336 10888 368 10920
rect 408 10888 440 10920
rect 480 10888 512 10920
rect 552 10888 584 10920
rect 624 10888 656 10920
rect 696 10888 728 10920
rect 768 10888 800 10920
rect 840 10888 872 10920
rect 912 10888 944 10920
rect 984 10888 1016 10920
rect 1056 10888 1088 10920
rect 1128 10888 1160 10920
rect 1200 10888 1232 10920
rect 1272 10888 1304 10920
rect 1344 10888 1376 10920
rect 1416 10888 1448 10920
rect 1488 10888 1520 10920
rect 1560 10888 1592 10920
rect 1632 10888 1664 10920
rect 1704 10888 1736 10920
rect 1776 10888 1808 10920
rect 1848 10888 1880 10920
rect 1920 10888 1952 10920
rect 48 10816 80 10848
rect 120 10816 152 10848
rect 192 10816 224 10848
rect 264 10816 296 10848
rect 336 10816 368 10848
rect 408 10816 440 10848
rect 480 10816 512 10848
rect 552 10816 584 10848
rect 624 10816 656 10848
rect 696 10816 728 10848
rect 768 10816 800 10848
rect 840 10816 872 10848
rect 912 10816 944 10848
rect 984 10816 1016 10848
rect 1056 10816 1088 10848
rect 1128 10816 1160 10848
rect 1200 10816 1232 10848
rect 1272 10816 1304 10848
rect 1344 10816 1376 10848
rect 1416 10816 1448 10848
rect 1488 10816 1520 10848
rect 1560 10816 1592 10848
rect 1632 10816 1664 10848
rect 1704 10816 1736 10848
rect 1776 10816 1808 10848
rect 1848 10816 1880 10848
rect 1920 10816 1952 10848
rect 48 10744 80 10776
rect 120 10744 152 10776
rect 192 10744 224 10776
rect 264 10744 296 10776
rect 336 10744 368 10776
rect 408 10744 440 10776
rect 480 10744 512 10776
rect 552 10744 584 10776
rect 624 10744 656 10776
rect 696 10744 728 10776
rect 768 10744 800 10776
rect 840 10744 872 10776
rect 912 10744 944 10776
rect 984 10744 1016 10776
rect 1056 10744 1088 10776
rect 1128 10744 1160 10776
rect 1200 10744 1232 10776
rect 1272 10744 1304 10776
rect 1344 10744 1376 10776
rect 1416 10744 1448 10776
rect 1488 10744 1520 10776
rect 1560 10744 1592 10776
rect 1632 10744 1664 10776
rect 1704 10744 1736 10776
rect 1776 10744 1808 10776
rect 1848 10744 1880 10776
rect 1920 10744 1952 10776
rect 48 10672 80 10704
rect 120 10672 152 10704
rect 192 10672 224 10704
rect 264 10672 296 10704
rect 336 10672 368 10704
rect 408 10672 440 10704
rect 480 10672 512 10704
rect 552 10672 584 10704
rect 624 10672 656 10704
rect 696 10672 728 10704
rect 768 10672 800 10704
rect 840 10672 872 10704
rect 912 10672 944 10704
rect 984 10672 1016 10704
rect 1056 10672 1088 10704
rect 1128 10672 1160 10704
rect 1200 10672 1232 10704
rect 1272 10672 1304 10704
rect 1344 10672 1376 10704
rect 1416 10672 1448 10704
rect 1488 10672 1520 10704
rect 1560 10672 1592 10704
rect 1632 10672 1664 10704
rect 1704 10672 1736 10704
rect 1776 10672 1808 10704
rect 1848 10672 1880 10704
rect 1920 10672 1952 10704
rect 48 10600 80 10632
rect 120 10600 152 10632
rect 192 10600 224 10632
rect 264 10600 296 10632
rect 336 10600 368 10632
rect 408 10600 440 10632
rect 480 10600 512 10632
rect 552 10600 584 10632
rect 624 10600 656 10632
rect 696 10600 728 10632
rect 768 10600 800 10632
rect 840 10600 872 10632
rect 912 10600 944 10632
rect 984 10600 1016 10632
rect 1056 10600 1088 10632
rect 1128 10600 1160 10632
rect 1200 10600 1232 10632
rect 1272 10600 1304 10632
rect 1344 10600 1376 10632
rect 1416 10600 1448 10632
rect 1488 10600 1520 10632
rect 1560 10600 1592 10632
rect 1632 10600 1664 10632
rect 1704 10600 1736 10632
rect 1776 10600 1808 10632
rect 1848 10600 1880 10632
rect 1920 10600 1952 10632
rect 48 10528 80 10560
rect 120 10528 152 10560
rect 192 10528 224 10560
rect 264 10528 296 10560
rect 336 10528 368 10560
rect 408 10528 440 10560
rect 480 10528 512 10560
rect 552 10528 584 10560
rect 624 10528 656 10560
rect 696 10528 728 10560
rect 768 10528 800 10560
rect 840 10528 872 10560
rect 912 10528 944 10560
rect 984 10528 1016 10560
rect 1056 10528 1088 10560
rect 1128 10528 1160 10560
rect 1200 10528 1232 10560
rect 1272 10528 1304 10560
rect 1344 10528 1376 10560
rect 1416 10528 1448 10560
rect 1488 10528 1520 10560
rect 1560 10528 1592 10560
rect 1632 10528 1664 10560
rect 1704 10528 1736 10560
rect 1776 10528 1808 10560
rect 1848 10528 1880 10560
rect 1920 10528 1952 10560
rect 48 10456 80 10488
rect 120 10456 152 10488
rect 192 10456 224 10488
rect 264 10456 296 10488
rect 336 10456 368 10488
rect 408 10456 440 10488
rect 480 10456 512 10488
rect 552 10456 584 10488
rect 624 10456 656 10488
rect 696 10456 728 10488
rect 768 10456 800 10488
rect 840 10456 872 10488
rect 912 10456 944 10488
rect 984 10456 1016 10488
rect 1056 10456 1088 10488
rect 1128 10456 1160 10488
rect 1200 10456 1232 10488
rect 1272 10456 1304 10488
rect 1344 10456 1376 10488
rect 1416 10456 1448 10488
rect 1488 10456 1520 10488
rect 1560 10456 1592 10488
rect 1632 10456 1664 10488
rect 1704 10456 1736 10488
rect 1776 10456 1808 10488
rect 1848 10456 1880 10488
rect 1920 10456 1952 10488
rect 48 10384 80 10416
rect 120 10384 152 10416
rect 192 10384 224 10416
rect 264 10384 296 10416
rect 336 10384 368 10416
rect 408 10384 440 10416
rect 480 10384 512 10416
rect 552 10384 584 10416
rect 624 10384 656 10416
rect 696 10384 728 10416
rect 768 10384 800 10416
rect 840 10384 872 10416
rect 912 10384 944 10416
rect 984 10384 1016 10416
rect 1056 10384 1088 10416
rect 1128 10384 1160 10416
rect 1200 10384 1232 10416
rect 1272 10384 1304 10416
rect 1344 10384 1376 10416
rect 1416 10384 1448 10416
rect 1488 10384 1520 10416
rect 1560 10384 1592 10416
rect 1632 10384 1664 10416
rect 1704 10384 1736 10416
rect 1776 10384 1808 10416
rect 1848 10384 1880 10416
rect 1920 10384 1952 10416
rect 48 10312 80 10344
rect 120 10312 152 10344
rect 192 10312 224 10344
rect 264 10312 296 10344
rect 336 10312 368 10344
rect 408 10312 440 10344
rect 480 10312 512 10344
rect 552 10312 584 10344
rect 624 10312 656 10344
rect 696 10312 728 10344
rect 768 10312 800 10344
rect 840 10312 872 10344
rect 912 10312 944 10344
rect 984 10312 1016 10344
rect 1056 10312 1088 10344
rect 1128 10312 1160 10344
rect 1200 10312 1232 10344
rect 1272 10312 1304 10344
rect 1344 10312 1376 10344
rect 1416 10312 1448 10344
rect 1488 10312 1520 10344
rect 1560 10312 1592 10344
rect 1632 10312 1664 10344
rect 1704 10312 1736 10344
rect 1776 10312 1808 10344
rect 1848 10312 1880 10344
rect 1920 10312 1952 10344
rect 48 10240 80 10272
rect 120 10240 152 10272
rect 192 10240 224 10272
rect 264 10240 296 10272
rect 336 10240 368 10272
rect 408 10240 440 10272
rect 480 10240 512 10272
rect 552 10240 584 10272
rect 624 10240 656 10272
rect 696 10240 728 10272
rect 768 10240 800 10272
rect 840 10240 872 10272
rect 912 10240 944 10272
rect 984 10240 1016 10272
rect 1056 10240 1088 10272
rect 1128 10240 1160 10272
rect 1200 10240 1232 10272
rect 1272 10240 1304 10272
rect 1344 10240 1376 10272
rect 1416 10240 1448 10272
rect 1488 10240 1520 10272
rect 1560 10240 1592 10272
rect 1632 10240 1664 10272
rect 1704 10240 1736 10272
rect 1776 10240 1808 10272
rect 1848 10240 1880 10272
rect 1920 10240 1952 10272
rect 48 10168 80 10200
rect 120 10168 152 10200
rect 192 10168 224 10200
rect 264 10168 296 10200
rect 336 10168 368 10200
rect 408 10168 440 10200
rect 480 10168 512 10200
rect 552 10168 584 10200
rect 624 10168 656 10200
rect 696 10168 728 10200
rect 768 10168 800 10200
rect 840 10168 872 10200
rect 912 10168 944 10200
rect 984 10168 1016 10200
rect 1056 10168 1088 10200
rect 1128 10168 1160 10200
rect 1200 10168 1232 10200
rect 1272 10168 1304 10200
rect 1344 10168 1376 10200
rect 1416 10168 1448 10200
rect 1488 10168 1520 10200
rect 1560 10168 1592 10200
rect 1632 10168 1664 10200
rect 1704 10168 1736 10200
rect 1776 10168 1808 10200
rect 1848 10168 1880 10200
rect 1920 10168 1952 10200
rect 48 10096 80 10128
rect 120 10096 152 10128
rect 192 10096 224 10128
rect 264 10096 296 10128
rect 336 10096 368 10128
rect 408 10096 440 10128
rect 480 10096 512 10128
rect 552 10096 584 10128
rect 624 10096 656 10128
rect 696 10096 728 10128
rect 768 10096 800 10128
rect 840 10096 872 10128
rect 912 10096 944 10128
rect 984 10096 1016 10128
rect 1056 10096 1088 10128
rect 1128 10096 1160 10128
rect 1200 10096 1232 10128
rect 1272 10096 1304 10128
rect 1344 10096 1376 10128
rect 1416 10096 1448 10128
rect 1488 10096 1520 10128
rect 1560 10096 1592 10128
rect 1632 10096 1664 10128
rect 1704 10096 1736 10128
rect 1776 10096 1808 10128
rect 1848 10096 1880 10128
rect 1920 10096 1952 10128
rect 48 10024 80 10056
rect 120 10024 152 10056
rect 192 10024 224 10056
rect 264 10024 296 10056
rect 336 10024 368 10056
rect 408 10024 440 10056
rect 480 10024 512 10056
rect 552 10024 584 10056
rect 624 10024 656 10056
rect 696 10024 728 10056
rect 768 10024 800 10056
rect 840 10024 872 10056
rect 912 10024 944 10056
rect 984 10024 1016 10056
rect 1056 10024 1088 10056
rect 1128 10024 1160 10056
rect 1200 10024 1232 10056
rect 1272 10024 1304 10056
rect 1344 10024 1376 10056
rect 1416 10024 1448 10056
rect 1488 10024 1520 10056
rect 1560 10024 1592 10056
rect 1632 10024 1664 10056
rect 1704 10024 1736 10056
rect 1776 10024 1808 10056
rect 1848 10024 1880 10056
rect 1920 10024 1952 10056
rect 48 9952 80 9984
rect 120 9952 152 9984
rect 192 9952 224 9984
rect 264 9952 296 9984
rect 336 9952 368 9984
rect 408 9952 440 9984
rect 480 9952 512 9984
rect 552 9952 584 9984
rect 624 9952 656 9984
rect 696 9952 728 9984
rect 768 9952 800 9984
rect 840 9952 872 9984
rect 912 9952 944 9984
rect 984 9952 1016 9984
rect 1056 9952 1088 9984
rect 1128 9952 1160 9984
rect 1200 9952 1232 9984
rect 1272 9952 1304 9984
rect 1344 9952 1376 9984
rect 1416 9952 1448 9984
rect 1488 9952 1520 9984
rect 1560 9952 1592 9984
rect 1632 9952 1664 9984
rect 1704 9952 1736 9984
rect 1776 9952 1808 9984
rect 1848 9952 1880 9984
rect 1920 9952 1952 9984
rect 48 9880 80 9912
rect 120 9880 152 9912
rect 192 9880 224 9912
rect 264 9880 296 9912
rect 336 9880 368 9912
rect 408 9880 440 9912
rect 480 9880 512 9912
rect 552 9880 584 9912
rect 624 9880 656 9912
rect 696 9880 728 9912
rect 768 9880 800 9912
rect 840 9880 872 9912
rect 912 9880 944 9912
rect 984 9880 1016 9912
rect 1056 9880 1088 9912
rect 1128 9880 1160 9912
rect 1200 9880 1232 9912
rect 1272 9880 1304 9912
rect 1344 9880 1376 9912
rect 1416 9880 1448 9912
rect 1488 9880 1520 9912
rect 1560 9880 1592 9912
rect 1632 9880 1664 9912
rect 1704 9880 1736 9912
rect 1776 9880 1808 9912
rect 1848 9880 1880 9912
rect 1920 9880 1952 9912
rect 48 9808 80 9840
rect 120 9808 152 9840
rect 192 9808 224 9840
rect 264 9808 296 9840
rect 336 9808 368 9840
rect 408 9808 440 9840
rect 480 9808 512 9840
rect 552 9808 584 9840
rect 624 9808 656 9840
rect 696 9808 728 9840
rect 768 9808 800 9840
rect 840 9808 872 9840
rect 912 9808 944 9840
rect 984 9808 1016 9840
rect 1056 9808 1088 9840
rect 1128 9808 1160 9840
rect 1200 9808 1232 9840
rect 1272 9808 1304 9840
rect 1344 9808 1376 9840
rect 1416 9808 1448 9840
rect 1488 9808 1520 9840
rect 1560 9808 1592 9840
rect 1632 9808 1664 9840
rect 1704 9808 1736 9840
rect 1776 9808 1808 9840
rect 1848 9808 1880 9840
rect 1920 9808 1952 9840
rect 48 9736 80 9768
rect 120 9736 152 9768
rect 192 9736 224 9768
rect 264 9736 296 9768
rect 336 9736 368 9768
rect 408 9736 440 9768
rect 480 9736 512 9768
rect 552 9736 584 9768
rect 624 9736 656 9768
rect 696 9736 728 9768
rect 768 9736 800 9768
rect 840 9736 872 9768
rect 912 9736 944 9768
rect 984 9736 1016 9768
rect 1056 9736 1088 9768
rect 1128 9736 1160 9768
rect 1200 9736 1232 9768
rect 1272 9736 1304 9768
rect 1344 9736 1376 9768
rect 1416 9736 1448 9768
rect 1488 9736 1520 9768
rect 1560 9736 1592 9768
rect 1632 9736 1664 9768
rect 1704 9736 1736 9768
rect 1776 9736 1808 9768
rect 1848 9736 1880 9768
rect 1920 9736 1952 9768
rect 48 9664 80 9696
rect 120 9664 152 9696
rect 192 9664 224 9696
rect 264 9664 296 9696
rect 336 9664 368 9696
rect 408 9664 440 9696
rect 480 9664 512 9696
rect 552 9664 584 9696
rect 624 9664 656 9696
rect 696 9664 728 9696
rect 768 9664 800 9696
rect 840 9664 872 9696
rect 912 9664 944 9696
rect 984 9664 1016 9696
rect 1056 9664 1088 9696
rect 1128 9664 1160 9696
rect 1200 9664 1232 9696
rect 1272 9664 1304 9696
rect 1344 9664 1376 9696
rect 1416 9664 1448 9696
rect 1488 9664 1520 9696
rect 1560 9664 1592 9696
rect 1632 9664 1664 9696
rect 1704 9664 1736 9696
rect 1776 9664 1808 9696
rect 1848 9664 1880 9696
rect 1920 9664 1952 9696
rect 48 9592 80 9624
rect 120 9592 152 9624
rect 192 9592 224 9624
rect 264 9592 296 9624
rect 336 9592 368 9624
rect 408 9592 440 9624
rect 480 9592 512 9624
rect 552 9592 584 9624
rect 624 9592 656 9624
rect 696 9592 728 9624
rect 768 9592 800 9624
rect 840 9592 872 9624
rect 912 9592 944 9624
rect 984 9592 1016 9624
rect 1056 9592 1088 9624
rect 1128 9592 1160 9624
rect 1200 9592 1232 9624
rect 1272 9592 1304 9624
rect 1344 9592 1376 9624
rect 1416 9592 1448 9624
rect 1488 9592 1520 9624
rect 1560 9592 1592 9624
rect 1632 9592 1664 9624
rect 1704 9592 1736 9624
rect 1776 9592 1808 9624
rect 1848 9592 1880 9624
rect 1920 9592 1952 9624
rect 48 9520 80 9552
rect 120 9520 152 9552
rect 192 9520 224 9552
rect 264 9520 296 9552
rect 336 9520 368 9552
rect 408 9520 440 9552
rect 480 9520 512 9552
rect 552 9520 584 9552
rect 624 9520 656 9552
rect 696 9520 728 9552
rect 768 9520 800 9552
rect 840 9520 872 9552
rect 912 9520 944 9552
rect 984 9520 1016 9552
rect 1056 9520 1088 9552
rect 1128 9520 1160 9552
rect 1200 9520 1232 9552
rect 1272 9520 1304 9552
rect 1344 9520 1376 9552
rect 1416 9520 1448 9552
rect 1488 9520 1520 9552
rect 1560 9520 1592 9552
rect 1632 9520 1664 9552
rect 1704 9520 1736 9552
rect 1776 9520 1808 9552
rect 1848 9520 1880 9552
rect 1920 9520 1952 9552
rect 48 9448 80 9480
rect 120 9448 152 9480
rect 192 9448 224 9480
rect 264 9448 296 9480
rect 336 9448 368 9480
rect 408 9448 440 9480
rect 480 9448 512 9480
rect 552 9448 584 9480
rect 624 9448 656 9480
rect 696 9448 728 9480
rect 768 9448 800 9480
rect 840 9448 872 9480
rect 912 9448 944 9480
rect 984 9448 1016 9480
rect 1056 9448 1088 9480
rect 1128 9448 1160 9480
rect 1200 9448 1232 9480
rect 1272 9448 1304 9480
rect 1344 9448 1376 9480
rect 1416 9448 1448 9480
rect 1488 9448 1520 9480
rect 1560 9448 1592 9480
rect 1632 9448 1664 9480
rect 1704 9448 1736 9480
rect 1776 9448 1808 9480
rect 1848 9448 1880 9480
rect 1920 9448 1952 9480
rect 48 9376 80 9408
rect 120 9376 152 9408
rect 192 9376 224 9408
rect 264 9376 296 9408
rect 336 9376 368 9408
rect 408 9376 440 9408
rect 480 9376 512 9408
rect 552 9376 584 9408
rect 624 9376 656 9408
rect 696 9376 728 9408
rect 768 9376 800 9408
rect 840 9376 872 9408
rect 912 9376 944 9408
rect 984 9376 1016 9408
rect 1056 9376 1088 9408
rect 1128 9376 1160 9408
rect 1200 9376 1232 9408
rect 1272 9376 1304 9408
rect 1344 9376 1376 9408
rect 1416 9376 1448 9408
rect 1488 9376 1520 9408
rect 1560 9376 1592 9408
rect 1632 9376 1664 9408
rect 1704 9376 1736 9408
rect 1776 9376 1808 9408
rect 1848 9376 1880 9408
rect 1920 9376 1952 9408
rect 48 9304 80 9336
rect 120 9304 152 9336
rect 192 9304 224 9336
rect 264 9304 296 9336
rect 336 9304 368 9336
rect 408 9304 440 9336
rect 480 9304 512 9336
rect 552 9304 584 9336
rect 624 9304 656 9336
rect 696 9304 728 9336
rect 768 9304 800 9336
rect 840 9304 872 9336
rect 912 9304 944 9336
rect 984 9304 1016 9336
rect 1056 9304 1088 9336
rect 1128 9304 1160 9336
rect 1200 9304 1232 9336
rect 1272 9304 1304 9336
rect 1344 9304 1376 9336
rect 1416 9304 1448 9336
rect 1488 9304 1520 9336
rect 1560 9304 1592 9336
rect 1632 9304 1664 9336
rect 1704 9304 1736 9336
rect 1776 9304 1808 9336
rect 1848 9304 1880 9336
rect 1920 9304 1952 9336
rect 48 9232 80 9264
rect 120 9232 152 9264
rect 192 9232 224 9264
rect 264 9232 296 9264
rect 336 9232 368 9264
rect 408 9232 440 9264
rect 480 9232 512 9264
rect 552 9232 584 9264
rect 624 9232 656 9264
rect 696 9232 728 9264
rect 768 9232 800 9264
rect 840 9232 872 9264
rect 912 9232 944 9264
rect 984 9232 1016 9264
rect 1056 9232 1088 9264
rect 1128 9232 1160 9264
rect 1200 9232 1232 9264
rect 1272 9232 1304 9264
rect 1344 9232 1376 9264
rect 1416 9232 1448 9264
rect 1488 9232 1520 9264
rect 1560 9232 1592 9264
rect 1632 9232 1664 9264
rect 1704 9232 1736 9264
rect 1776 9232 1808 9264
rect 1848 9232 1880 9264
rect 1920 9232 1952 9264
rect 48 9160 80 9192
rect 120 9160 152 9192
rect 192 9160 224 9192
rect 264 9160 296 9192
rect 336 9160 368 9192
rect 408 9160 440 9192
rect 480 9160 512 9192
rect 552 9160 584 9192
rect 624 9160 656 9192
rect 696 9160 728 9192
rect 768 9160 800 9192
rect 840 9160 872 9192
rect 912 9160 944 9192
rect 984 9160 1016 9192
rect 1056 9160 1088 9192
rect 1128 9160 1160 9192
rect 1200 9160 1232 9192
rect 1272 9160 1304 9192
rect 1344 9160 1376 9192
rect 1416 9160 1448 9192
rect 1488 9160 1520 9192
rect 1560 9160 1592 9192
rect 1632 9160 1664 9192
rect 1704 9160 1736 9192
rect 1776 9160 1808 9192
rect 1848 9160 1880 9192
rect 1920 9160 1952 9192
rect 48 9088 80 9120
rect 120 9088 152 9120
rect 192 9088 224 9120
rect 264 9088 296 9120
rect 336 9088 368 9120
rect 408 9088 440 9120
rect 480 9088 512 9120
rect 552 9088 584 9120
rect 624 9088 656 9120
rect 696 9088 728 9120
rect 768 9088 800 9120
rect 840 9088 872 9120
rect 912 9088 944 9120
rect 984 9088 1016 9120
rect 1056 9088 1088 9120
rect 1128 9088 1160 9120
rect 1200 9088 1232 9120
rect 1272 9088 1304 9120
rect 1344 9088 1376 9120
rect 1416 9088 1448 9120
rect 1488 9088 1520 9120
rect 1560 9088 1592 9120
rect 1632 9088 1664 9120
rect 1704 9088 1736 9120
rect 1776 9088 1808 9120
rect 1848 9088 1880 9120
rect 1920 9088 1952 9120
rect 48 9016 80 9048
rect 120 9016 152 9048
rect 192 9016 224 9048
rect 264 9016 296 9048
rect 336 9016 368 9048
rect 408 9016 440 9048
rect 480 9016 512 9048
rect 552 9016 584 9048
rect 624 9016 656 9048
rect 696 9016 728 9048
rect 768 9016 800 9048
rect 840 9016 872 9048
rect 912 9016 944 9048
rect 984 9016 1016 9048
rect 1056 9016 1088 9048
rect 1128 9016 1160 9048
rect 1200 9016 1232 9048
rect 1272 9016 1304 9048
rect 1344 9016 1376 9048
rect 1416 9016 1448 9048
rect 1488 9016 1520 9048
rect 1560 9016 1592 9048
rect 1632 9016 1664 9048
rect 1704 9016 1736 9048
rect 1776 9016 1808 9048
rect 1848 9016 1880 9048
rect 1920 9016 1952 9048
rect 48 8944 80 8976
rect 120 8944 152 8976
rect 192 8944 224 8976
rect 264 8944 296 8976
rect 336 8944 368 8976
rect 408 8944 440 8976
rect 480 8944 512 8976
rect 552 8944 584 8976
rect 624 8944 656 8976
rect 696 8944 728 8976
rect 768 8944 800 8976
rect 840 8944 872 8976
rect 912 8944 944 8976
rect 984 8944 1016 8976
rect 1056 8944 1088 8976
rect 1128 8944 1160 8976
rect 1200 8944 1232 8976
rect 1272 8944 1304 8976
rect 1344 8944 1376 8976
rect 1416 8944 1448 8976
rect 1488 8944 1520 8976
rect 1560 8944 1592 8976
rect 1632 8944 1664 8976
rect 1704 8944 1736 8976
rect 1776 8944 1808 8976
rect 1848 8944 1880 8976
rect 1920 8944 1952 8976
rect 48 8872 80 8904
rect 120 8872 152 8904
rect 192 8872 224 8904
rect 264 8872 296 8904
rect 336 8872 368 8904
rect 408 8872 440 8904
rect 480 8872 512 8904
rect 552 8872 584 8904
rect 624 8872 656 8904
rect 696 8872 728 8904
rect 768 8872 800 8904
rect 840 8872 872 8904
rect 912 8872 944 8904
rect 984 8872 1016 8904
rect 1056 8872 1088 8904
rect 1128 8872 1160 8904
rect 1200 8872 1232 8904
rect 1272 8872 1304 8904
rect 1344 8872 1376 8904
rect 1416 8872 1448 8904
rect 1488 8872 1520 8904
rect 1560 8872 1592 8904
rect 1632 8872 1664 8904
rect 1704 8872 1736 8904
rect 1776 8872 1808 8904
rect 1848 8872 1880 8904
rect 1920 8872 1952 8904
rect 48 8800 80 8832
rect 120 8800 152 8832
rect 192 8800 224 8832
rect 264 8800 296 8832
rect 336 8800 368 8832
rect 408 8800 440 8832
rect 480 8800 512 8832
rect 552 8800 584 8832
rect 624 8800 656 8832
rect 696 8800 728 8832
rect 768 8800 800 8832
rect 840 8800 872 8832
rect 912 8800 944 8832
rect 984 8800 1016 8832
rect 1056 8800 1088 8832
rect 1128 8800 1160 8832
rect 1200 8800 1232 8832
rect 1272 8800 1304 8832
rect 1344 8800 1376 8832
rect 1416 8800 1448 8832
rect 1488 8800 1520 8832
rect 1560 8800 1592 8832
rect 1632 8800 1664 8832
rect 1704 8800 1736 8832
rect 1776 8800 1808 8832
rect 1848 8800 1880 8832
rect 1920 8800 1952 8832
rect 48 8728 80 8760
rect 120 8728 152 8760
rect 192 8728 224 8760
rect 264 8728 296 8760
rect 336 8728 368 8760
rect 408 8728 440 8760
rect 480 8728 512 8760
rect 552 8728 584 8760
rect 624 8728 656 8760
rect 696 8728 728 8760
rect 768 8728 800 8760
rect 840 8728 872 8760
rect 912 8728 944 8760
rect 984 8728 1016 8760
rect 1056 8728 1088 8760
rect 1128 8728 1160 8760
rect 1200 8728 1232 8760
rect 1272 8728 1304 8760
rect 1344 8728 1376 8760
rect 1416 8728 1448 8760
rect 1488 8728 1520 8760
rect 1560 8728 1592 8760
rect 1632 8728 1664 8760
rect 1704 8728 1736 8760
rect 1776 8728 1808 8760
rect 1848 8728 1880 8760
rect 1920 8728 1952 8760
rect 48 8656 80 8688
rect 120 8656 152 8688
rect 192 8656 224 8688
rect 264 8656 296 8688
rect 336 8656 368 8688
rect 408 8656 440 8688
rect 480 8656 512 8688
rect 552 8656 584 8688
rect 624 8656 656 8688
rect 696 8656 728 8688
rect 768 8656 800 8688
rect 840 8656 872 8688
rect 912 8656 944 8688
rect 984 8656 1016 8688
rect 1056 8656 1088 8688
rect 1128 8656 1160 8688
rect 1200 8656 1232 8688
rect 1272 8656 1304 8688
rect 1344 8656 1376 8688
rect 1416 8656 1448 8688
rect 1488 8656 1520 8688
rect 1560 8656 1592 8688
rect 1632 8656 1664 8688
rect 1704 8656 1736 8688
rect 1776 8656 1808 8688
rect 1848 8656 1880 8688
rect 1920 8656 1952 8688
rect 48 8584 80 8616
rect 120 8584 152 8616
rect 192 8584 224 8616
rect 264 8584 296 8616
rect 336 8584 368 8616
rect 408 8584 440 8616
rect 480 8584 512 8616
rect 552 8584 584 8616
rect 624 8584 656 8616
rect 696 8584 728 8616
rect 768 8584 800 8616
rect 840 8584 872 8616
rect 912 8584 944 8616
rect 984 8584 1016 8616
rect 1056 8584 1088 8616
rect 1128 8584 1160 8616
rect 1200 8584 1232 8616
rect 1272 8584 1304 8616
rect 1344 8584 1376 8616
rect 1416 8584 1448 8616
rect 1488 8584 1520 8616
rect 1560 8584 1592 8616
rect 1632 8584 1664 8616
rect 1704 8584 1736 8616
rect 1776 8584 1808 8616
rect 1848 8584 1880 8616
rect 1920 8584 1952 8616
rect 48 8512 80 8544
rect 120 8512 152 8544
rect 192 8512 224 8544
rect 264 8512 296 8544
rect 336 8512 368 8544
rect 408 8512 440 8544
rect 480 8512 512 8544
rect 552 8512 584 8544
rect 624 8512 656 8544
rect 696 8512 728 8544
rect 768 8512 800 8544
rect 840 8512 872 8544
rect 912 8512 944 8544
rect 984 8512 1016 8544
rect 1056 8512 1088 8544
rect 1128 8512 1160 8544
rect 1200 8512 1232 8544
rect 1272 8512 1304 8544
rect 1344 8512 1376 8544
rect 1416 8512 1448 8544
rect 1488 8512 1520 8544
rect 1560 8512 1592 8544
rect 1632 8512 1664 8544
rect 1704 8512 1736 8544
rect 1776 8512 1808 8544
rect 1848 8512 1880 8544
rect 1920 8512 1952 8544
rect 48 8440 80 8472
rect 120 8440 152 8472
rect 192 8440 224 8472
rect 264 8440 296 8472
rect 336 8440 368 8472
rect 408 8440 440 8472
rect 480 8440 512 8472
rect 552 8440 584 8472
rect 624 8440 656 8472
rect 696 8440 728 8472
rect 768 8440 800 8472
rect 840 8440 872 8472
rect 912 8440 944 8472
rect 984 8440 1016 8472
rect 1056 8440 1088 8472
rect 1128 8440 1160 8472
rect 1200 8440 1232 8472
rect 1272 8440 1304 8472
rect 1344 8440 1376 8472
rect 1416 8440 1448 8472
rect 1488 8440 1520 8472
rect 1560 8440 1592 8472
rect 1632 8440 1664 8472
rect 1704 8440 1736 8472
rect 1776 8440 1808 8472
rect 1848 8440 1880 8472
rect 1920 8440 1952 8472
rect 48 8368 80 8400
rect 120 8368 152 8400
rect 192 8368 224 8400
rect 264 8368 296 8400
rect 336 8368 368 8400
rect 408 8368 440 8400
rect 480 8368 512 8400
rect 552 8368 584 8400
rect 624 8368 656 8400
rect 696 8368 728 8400
rect 768 8368 800 8400
rect 840 8368 872 8400
rect 912 8368 944 8400
rect 984 8368 1016 8400
rect 1056 8368 1088 8400
rect 1128 8368 1160 8400
rect 1200 8368 1232 8400
rect 1272 8368 1304 8400
rect 1344 8368 1376 8400
rect 1416 8368 1448 8400
rect 1488 8368 1520 8400
rect 1560 8368 1592 8400
rect 1632 8368 1664 8400
rect 1704 8368 1736 8400
rect 1776 8368 1808 8400
rect 1848 8368 1880 8400
rect 1920 8368 1952 8400
rect 48 8296 80 8328
rect 120 8296 152 8328
rect 192 8296 224 8328
rect 264 8296 296 8328
rect 336 8296 368 8328
rect 408 8296 440 8328
rect 480 8296 512 8328
rect 552 8296 584 8328
rect 624 8296 656 8328
rect 696 8296 728 8328
rect 768 8296 800 8328
rect 840 8296 872 8328
rect 912 8296 944 8328
rect 984 8296 1016 8328
rect 1056 8296 1088 8328
rect 1128 8296 1160 8328
rect 1200 8296 1232 8328
rect 1272 8296 1304 8328
rect 1344 8296 1376 8328
rect 1416 8296 1448 8328
rect 1488 8296 1520 8328
rect 1560 8296 1592 8328
rect 1632 8296 1664 8328
rect 1704 8296 1736 8328
rect 1776 8296 1808 8328
rect 1848 8296 1880 8328
rect 1920 8296 1952 8328
rect 48 8224 80 8256
rect 120 8224 152 8256
rect 192 8224 224 8256
rect 264 8224 296 8256
rect 336 8224 368 8256
rect 408 8224 440 8256
rect 480 8224 512 8256
rect 552 8224 584 8256
rect 624 8224 656 8256
rect 696 8224 728 8256
rect 768 8224 800 8256
rect 840 8224 872 8256
rect 912 8224 944 8256
rect 984 8224 1016 8256
rect 1056 8224 1088 8256
rect 1128 8224 1160 8256
rect 1200 8224 1232 8256
rect 1272 8224 1304 8256
rect 1344 8224 1376 8256
rect 1416 8224 1448 8256
rect 1488 8224 1520 8256
rect 1560 8224 1592 8256
rect 1632 8224 1664 8256
rect 1704 8224 1736 8256
rect 1776 8224 1808 8256
rect 1848 8224 1880 8256
rect 1920 8224 1952 8256
rect 48 8152 80 8184
rect 120 8152 152 8184
rect 192 8152 224 8184
rect 264 8152 296 8184
rect 336 8152 368 8184
rect 408 8152 440 8184
rect 480 8152 512 8184
rect 552 8152 584 8184
rect 624 8152 656 8184
rect 696 8152 728 8184
rect 768 8152 800 8184
rect 840 8152 872 8184
rect 912 8152 944 8184
rect 984 8152 1016 8184
rect 1056 8152 1088 8184
rect 1128 8152 1160 8184
rect 1200 8152 1232 8184
rect 1272 8152 1304 8184
rect 1344 8152 1376 8184
rect 1416 8152 1448 8184
rect 1488 8152 1520 8184
rect 1560 8152 1592 8184
rect 1632 8152 1664 8184
rect 1704 8152 1736 8184
rect 1776 8152 1808 8184
rect 1848 8152 1880 8184
rect 1920 8152 1952 8184
rect 48 8080 80 8112
rect 120 8080 152 8112
rect 192 8080 224 8112
rect 264 8080 296 8112
rect 336 8080 368 8112
rect 408 8080 440 8112
rect 480 8080 512 8112
rect 552 8080 584 8112
rect 624 8080 656 8112
rect 696 8080 728 8112
rect 768 8080 800 8112
rect 840 8080 872 8112
rect 912 8080 944 8112
rect 984 8080 1016 8112
rect 1056 8080 1088 8112
rect 1128 8080 1160 8112
rect 1200 8080 1232 8112
rect 1272 8080 1304 8112
rect 1344 8080 1376 8112
rect 1416 8080 1448 8112
rect 1488 8080 1520 8112
rect 1560 8080 1592 8112
rect 1632 8080 1664 8112
rect 1704 8080 1736 8112
rect 1776 8080 1808 8112
rect 1848 8080 1880 8112
rect 1920 8080 1952 8112
rect 48 8008 80 8040
rect 120 8008 152 8040
rect 192 8008 224 8040
rect 264 8008 296 8040
rect 336 8008 368 8040
rect 408 8008 440 8040
rect 480 8008 512 8040
rect 552 8008 584 8040
rect 624 8008 656 8040
rect 696 8008 728 8040
rect 768 8008 800 8040
rect 840 8008 872 8040
rect 912 8008 944 8040
rect 984 8008 1016 8040
rect 1056 8008 1088 8040
rect 1128 8008 1160 8040
rect 1200 8008 1232 8040
rect 1272 8008 1304 8040
rect 1344 8008 1376 8040
rect 1416 8008 1448 8040
rect 1488 8008 1520 8040
rect 1560 8008 1592 8040
rect 1632 8008 1664 8040
rect 1704 8008 1736 8040
rect 1776 8008 1808 8040
rect 1848 8008 1880 8040
rect 1920 8008 1952 8040
rect 48 7936 80 7968
rect 120 7936 152 7968
rect 192 7936 224 7968
rect 264 7936 296 7968
rect 336 7936 368 7968
rect 408 7936 440 7968
rect 480 7936 512 7968
rect 552 7936 584 7968
rect 624 7936 656 7968
rect 696 7936 728 7968
rect 768 7936 800 7968
rect 840 7936 872 7968
rect 912 7936 944 7968
rect 984 7936 1016 7968
rect 1056 7936 1088 7968
rect 1128 7936 1160 7968
rect 1200 7936 1232 7968
rect 1272 7936 1304 7968
rect 1344 7936 1376 7968
rect 1416 7936 1448 7968
rect 1488 7936 1520 7968
rect 1560 7936 1592 7968
rect 1632 7936 1664 7968
rect 1704 7936 1736 7968
rect 1776 7936 1808 7968
rect 1848 7936 1880 7968
rect 1920 7936 1952 7968
rect 48 7864 80 7896
rect 120 7864 152 7896
rect 192 7864 224 7896
rect 264 7864 296 7896
rect 336 7864 368 7896
rect 408 7864 440 7896
rect 480 7864 512 7896
rect 552 7864 584 7896
rect 624 7864 656 7896
rect 696 7864 728 7896
rect 768 7864 800 7896
rect 840 7864 872 7896
rect 912 7864 944 7896
rect 984 7864 1016 7896
rect 1056 7864 1088 7896
rect 1128 7864 1160 7896
rect 1200 7864 1232 7896
rect 1272 7864 1304 7896
rect 1344 7864 1376 7896
rect 1416 7864 1448 7896
rect 1488 7864 1520 7896
rect 1560 7864 1592 7896
rect 1632 7864 1664 7896
rect 1704 7864 1736 7896
rect 1776 7864 1808 7896
rect 1848 7864 1880 7896
rect 1920 7864 1952 7896
rect 48 7792 80 7824
rect 120 7792 152 7824
rect 192 7792 224 7824
rect 264 7792 296 7824
rect 336 7792 368 7824
rect 408 7792 440 7824
rect 480 7792 512 7824
rect 552 7792 584 7824
rect 624 7792 656 7824
rect 696 7792 728 7824
rect 768 7792 800 7824
rect 840 7792 872 7824
rect 912 7792 944 7824
rect 984 7792 1016 7824
rect 1056 7792 1088 7824
rect 1128 7792 1160 7824
rect 1200 7792 1232 7824
rect 1272 7792 1304 7824
rect 1344 7792 1376 7824
rect 1416 7792 1448 7824
rect 1488 7792 1520 7824
rect 1560 7792 1592 7824
rect 1632 7792 1664 7824
rect 1704 7792 1736 7824
rect 1776 7792 1808 7824
rect 1848 7792 1880 7824
rect 1920 7792 1952 7824
rect 48 7720 80 7752
rect 120 7720 152 7752
rect 192 7720 224 7752
rect 264 7720 296 7752
rect 336 7720 368 7752
rect 408 7720 440 7752
rect 480 7720 512 7752
rect 552 7720 584 7752
rect 624 7720 656 7752
rect 696 7720 728 7752
rect 768 7720 800 7752
rect 840 7720 872 7752
rect 912 7720 944 7752
rect 984 7720 1016 7752
rect 1056 7720 1088 7752
rect 1128 7720 1160 7752
rect 1200 7720 1232 7752
rect 1272 7720 1304 7752
rect 1344 7720 1376 7752
rect 1416 7720 1448 7752
rect 1488 7720 1520 7752
rect 1560 7720 1592 7752
rect 1632 7720 1664 7752
rect 1704 7720 1736 7752
rect 1776 7720 1808 7752
rect 1848 7720 1880 7752
rect 1920 7720 1952 7752
rect 48 7648 80 7680
rect 120 7648 152 7680
rect 192 7648 224 7680
rect 264 7648 296 7680
rect 336 7648 368 7680
rect 408 7648 440 7680
rect 480 7648 512 7680
rect 552 7648 584 7680
rect 624 7648 656 7680
rect 696 7648 728 7680
rect 768 7648 800 7680
rect 840 7648 872 7680
rect 912 7648 944 7680
rect 984 7648 1016 7680
rect 1056 7648 1088 7680
rect 1128 7648 1160 7680
rect 1200 7648 1232 7680
rect 1272 7648 1304 7680
rect 1344 7648 1376 7680
rect 1416 7648 1448 7680
rect 1488 7648 1520 7680
rect 1560 7648 1592 7680
rect 1632 7648 1664 7680
rect 1704 7648 1736 7680
rect 1776 7648 1808 7680
rect 1848 7648 1880 7680
rect 1920 7648 1952 7680
rect 48 7576 80 7608
rect 120 7576 152 7608
rect 192 7576 224 7608
rect 264 7576 296 7608
rect 336 7576 368 7608
rect 408 7576 440 7608
rect 480 7576 512 7608
rect 552 7576 584 7608
rect 624 7576 656 7608
rect 696 7576 728 7608
rect 768 7576 800 7608
rect 840 7576 872 7608
rect 912 7576 944 7608
rect 984 7576 1016 7608
rect 1056 7576 1088 7608
rect 1128 7576 1160 7608
rect 1200 7576 1232 7608
rect 1272 7576 1304 7608
rect 1344 7576 1376 7608
rect 1416 7576 1448 7608
rect 1488 7576 1520 7608
rect 1560 7576 1592 7608
rect 1632 7576 1664 7608
rect 1704 7576 1736 7608
rect 1776 7576 1808 7608
rect 1848 7576 1880 7608
rect 1920 7576 1952 7608
rect 48 7504 80 7536
rect 120 7504 152 7536
rect 192 7504 224 7536
rect 264 7504 296 7536
rect 336 7504 368 7536
rect 408 7504 440 7536
rect 480 7504 512 7536
rect 552 7504 584 7536
rect 624 7504 656 7536
rect 696 7504 728 7536
rect 768 7504 800 7536
rect 840 7504 872 7536
rect 912 7504 944 7536
rect 984 7504 1016 7536
rect 1056 7504 1088 7536
rect 1128 7504 1160 7536
rect 1200 7504 1232 7536
rect 1272 7504 1304 7536
rect 1344 7504 1376 7536
rect 1416 7504 1448 7536
rect 1488 7504 1520 7536
rect 1560 7504 1592 7536
rect 1632 7504 1664 7536
rect 1704 7504 1736 7536
rect 1776 7504 1808 7536
rect 1848 7504 1880 7536
rect 1920 7504 1952 7536
rect 48 7432 80 7464
rect 120 7432 152 7464
rect 192 7432 224 7464
rect 264 7432 296 7464
rect 336 7432 368 7464
rect 408 7432 440 7464
rect 480 7432 512 7464
rect 552 7432 584 7464
rect 624 7432 656 7464
rect 696 7432 728 7464
rect 768 7432 800 7464
rect 840 7432 872 7464
rect 912 7432 944 7464
rect 984 7432 1016 7464
rect 1056 7432 1088 7464
rect 1128 7432 1160 7464
rect 1200 7432 1232 7464
rect 1272 7432 1304 7464
rect 1344 7432 1376 7464
rect 1416 7432 1448 7464
rect 1488 7432 1520 7464
rect 1560 7432 1592 7464
rect 1632 7432 1664 7464
rect 1704 7432 1736 7464
rect 1776 7432 1808 7464
rect 1848 7432 1880 7464
rect 1920 7432 1952 7464
rect 48 7360 80 7392
rect 120 7360 152 7392
rect 192 7360 224 7392
rect 264 7360 296 7392
rect 336 7360 368 7392
rect 408 7360 440 7392
rect 480 7360 512 7392
rect 552 7360 584 7392
rect 624 7360 656 7392
rect 696 7360 728 7392
rect 768 7360 800 7392
rect 840 7360 872 7392
rect 912 7360 944 7392
rect 984 7360 1016 7392
rect 1056 7360 1088 7392
rect 1128 7360 1160 7392
rect 1200 7360 1232 7392
rect 1272 7360 1304 7392
rect 1344 7360 1376 7392
rect 1416 7360 1448 7392
rect 1488 7360 1520 7392
rect 1560 7360 1592 7392
rect 1632 7360 1664 7392
rect 1704 7360 1736 7392
rect 1776 7360 1808 7392
rect 1848 7360 1880 7392
rect 1920 7360 1952 7392
rect 48 7288 80 7320
rect 120 7288 152 7320
rect 192 7288 224 7320
rect 264 7288 296 7320
rect 336 7288 368 7320
rect 408 7288 440 7320
rect 480 7288 512 7320
rect 552 7288 584 7320
rect 624 7288 656 7320
rect 696 7288 728 7320
rect 768 7288 800 7320
rect 840 7288 872 7320
rect 912 7288 944 7320
rect 984 7288 1016 7320
rect 1056 7288 1088 7320
rect 1128 7288 1160 7320
rect 1200 7288 1232 7320
rect 1272 7288 1304 7320
rect 1344 7288 1376 7320
rect 1416 7288 1448 7320
rect 1488 7288 1520 7320
rect 1560 7288 1592 7320
rect 1632 7288 1664 7320
rect 1704 7288 1736 7320
rect 1776 7288 1808 7320
rect 1848 7288 1880 7320
rect 1920 7288 1952 7320
rect 48 7216 80 7248
rect 120 7216 152 7248
rect 192 7216 224 7248
rect 264 7216 296 7248
rect 336 7216 368 7248
rect 408 7216 440 7248
rect 480 7216 512 7248
rect 552 7216 584 7248
rect 624 7216 656 7248
rect 696 7216 728 7248
rect 768 7216 800 7248
rect 840 7216 872 7248
rect 912 7216 944 7248
rect 984 7216 1016 7248
rect 1056 7216 1088 7248
rect 1128 7216 1160 7248
rect 1200 7216 1232 7248
rect 1272 7216 1304 7248
rect 1344 7216 1376 7248
rect 1416 7216 1448 7248
rect 1488 7216 1520 7248
rect 1560 7216 1592 7248
rect 1632 7216 1664 7248
rect 1704 7216 1736 7248
rect 1776 7216 1808 7248
rect 1848 7216 1880 7248
rect 1920 7216 1952 7248
rect 48 7144 80 7176
rect 120 7144 152 7176
rect 192 7144 224 7176
rect 264 7144 296 7176
rect 336 7144 368 7176
rect 408 7144 440 7176
rect 480 7144 512 7176
rect 552 7144 584 7176
rect 624 7144 656 7176
rect 696 7144 728 7176
rect 768 7144 800 7176
rect 840 7144 872 7176
rect 912 7144 944 7176
rect 984 7144 1016 7176
rect 1056 7144 1088 7176
rect 1128 7144 1160 7176
rect 1200 7144 1232 7176
rect 1272 7144 1304 7176
rect 1344 7144 1376 7176
rect 1416 7144 1448 7176
rect 1488 7144 1520 7176
rect 1560 7144 1592 7176
rect 1632 7144 1664 7176
rect 1704 7144 1736 7176
rect 1776 7144 1808 7176
rect 1848 7144 1880 7176
rect 1920 7144 1952 7176
rect 48 7072 80 7104
rect 120 7072 152 7104
rect 192 7072 224 7104
rect 264 7072 296 7104
rect 336 7072 368 7104
rect 408 7072 440 7104
rect 480 7072 512 7104
rect 552 7072 584 7104
rect 624 7072 656 7104
rect 696 7072 728 7104
rect 768 7072 800 7104
rect 840 7072 872 7104
rect 912 7072 944 7104
rect 984 7072 1016 7104
rect 1056 7072 1088 7104
rect 1128 7072 1160 7104
rect 1200 7072 1232 7104
rect 1272 7072 1304 7104
rect 1344 7072 1376 7104
rect 1416 7072 1448 7104
rect 1488 7072 1520 7104
rect 1560 7072 1592 7104
rect 1632 7072 1664 7104
rect 1704 7072 1736 7104
rect 1776 7072 1808 7104
rect 1848 7072 1880 7104
rect 1920 7072 1952 7104
rect 48 7000 80 7032
rect 120 7000 152 7032
rect 192 7000 224 7032
rect 264 7000 296 7032
rect 336 7000 368 7032
rect 408 7000 440 7032
rect 480 7000 512 7032
rect 552 7000 584 7032
rect 624 7000 656 7032
rect 696 7000 728 7032
rect 768 7000 800 7032
rect 840 7000 872 7032
rect 912 7000 944 7032
rect 984 7000 1016 7032
rect 1056 7000 1088 7032
rect 1128 7000 1160 7032
rect 1200 7000 1232 7032
rect 1272 7000 1304 7032
rect 1344 7000 1376 7032
rect 1416 7000 1448 7032
rect 1488 7000 1520 7032
rect 1560 7000 1592 7032
rect 1632 7000 1664 7032
rect 1704 7000 1736 7032
rect 1776 7000 1808 7032
rect 1848 7000 1880 7032
rect 1920 7000 1952 7032
rect 48 6928 80 6960
rect 120 6928 152 6960
rect 192 6928 224 6960
rect 264 6928 296 6960
rect 336 6928 368 6960
rect 408 6928 440 6960
rect 480 6928 512 6960
rect 552 6928 584 6960
rect 624 6928 656 6960
rect 696 6928 728 6960
rect 768 6928 800 6960
rect 840 6928 872 6960
rect 912 6928 944 6960
rect 984 6928 1016 6960
rect 1056 6928 1088 6960
rect 1128 6928 1160 6960
rect 1200 6928 1232 6960
rect 1272 6928 1304 6960
rect 1344 6928 1376 6960
rect 1416 6928 1448 6960
rect 1488 6928 1520 6960
rect 1560 6928 1592 6960
rect 1632 6928 1664 6960
rect 1704 6928 1736 6960
rect 1776 6928 1808 6960
rect 1848 6928 1880 6960
rect 1920 6928 1952 6960
rect 48 6856 80 6888
rect 120 6856 152 6888
rect 192 6856 224 6888
rect 264 6856 296 6888
rect 336 6856 368 6888
rect 408 6856 440 6888
rect 480 6856 512 6888
rect 552 6856 584 6888
rect 624 6856 656 6888
rect 696 6856 728 6888
rect 768 6856 800 6888
rect 840 6856 872 6888
rect 912 6856 944 6888
rect 984 6856 1016 6888
rect 1056 6856 1088 6888
rect 1128 6856 1160 6888
rect 1200 6856 1232 6888
rect 1272 6856 1304 6888
rect 1344 6856 1376 6888
rect 1416 6856 1448 6888
rect 1488 6856 1520 6888
rect 1560 6856 1592 6888
rect 1632 6856 1664 6888
rect 1704 6856 1736 6888
rect 1776 6856 1808 6888
rect 1848 6856 1880 6888
rect 1920 6856 1952 6888
rect 120 6512 152 6544
rect 192 6512 224 6544
rect 264 6512 296 6544
rect 336 6512 368 6544
rect 408 6512 440 6544
rect 480 6512 512 6544
rect 552 6512 584 6544
rect 624 6512 656 6544
rect 696 6512 728 6544
rect 768 6512 800 6544
rect 840 6512 872 6544
rect 912 6512 944 6544
rect 984 6512 1016 6544
rect 1056 6512 1088 6544
rect 1128 6512 1160 6544
rect 1200 6512 1232 6544
rect 1272 6512 1304 6544
rect 1344 6512 1376 6544
rect 1416 6512 1448 6544
rect 1488 6512 1520 6544
rect 1560 6512 1592 6544
rect 1632 6512 1664 6544
rect 1704 6512 1736 6544
rect 1776 6512 1808 6544
rect 1848 6512 1880 6544
rect 1920 6512 1952 6544
rect 48 6440 80 6472
rect 120 6440 152 6472
rect 192 6440 224 6472
rect 264 6440 296 6472
rect 336 6440 368 6472
rect 408 6440 440 6472
rect 480 6440 512 6472
rect 552 6440 584 6472
rect 624 6440 656 6472
rect 696 6440 728 6472
rect 768 6440 800 6472
rect 840 6440 872 6472
rect 912 6440 944 6472
rect 984 6440 1016 6472
rect 1056 6440 1088 6472
rect 1128 6440 1160 6472
rect 1200 6440 1232 6472
rect 1272 6440 1304 6472
rect 1344 6440 1376 6472
rect 1416 6440 1448 6472
rect 1488 6440 1520 6472
rect 1560 6440 1592 6472
rect 1632 6440 1664 6472
rect 1704 6440 1736 6472
rect 1776 6440 1808 6472
rect 1848 6440 1880 6472
rect 1920 6440 1952 6472
rect 48 6368 80 6400
rect 120 6368 152 6400
rect 192 6368 224 6400
rect 264 6368 296 6400
rect 336 6368 368 6400
rect 408 6368 440 6400
rect 480 6368 512 6400
rect 552 6368 584 6400
rect 624 6368 656 6400
rect 696 6368 728 6400
rect 768 6368 800 6400
rect 840 6368 872 6400
rect 912 6368 944 6400
rect 984 6368 1016 6400
rect 1056 6368 1088 6400
rect 1128 6368 1160 6400
rect 1200 6368 1232 6400
rect 1272 6368 1304 6400
rect 1344 6368 1376 6400
rect 1416 6368 1448 6400
rect 1488 6368 1520 6400
rect 1560 6368 1592 6400
rect 1632 6368 1664 6400
rect 1704 6368 1736 6400
rect 1776 6368 1808 6400
rect 1848 6368 1880 6400
rect 1920 6368 1952 6400
rect 48 6296 80 6328
rect 120 6296 152 6328
rect 192 6296 224 6328
rect 264 6296 296 6328
rect 336 6296 368 6328
rect 408 6296 440 6328
rect 480 6296 512 6328
rect 552 6296 584 6328
rect 624 6296 656 6328
rect 696 6296 728 6328
rect 768 6296 800 6328
rect 840 6296 872 6328
rect 912 6296 944 6328
rect 984 6296 1016 6328
rect 1056 6296 1088 6328
rect 1128 6296 1160 6328
rect 1200 6296 1232 6328
rect 1272 6296 1304 6328
rect 1344 6296 1376 6328
rect 1416 6296 1448 6328
rect 1488 6296 1520 6328
rect 1560 6296 1592 6328
rect 1632 6296 1664 6328
rect 1704 6296 1736 6328
rect 1776 6296 1808 6328
rect 1848 6296 1880 6328
rect 1920 6296 1952 6328
rect 48 6224 80 6256
rect 120 6224 152 6256
rect 192 6224 224 6256
rect 264 6224 296 6256
rect 336 6224 368 6256
rect 408 6224 440 6256
rect 480 6224 512 6256
rect 552 6224 584 6256
rect 624 6224 656 6256
rect 696 6224 728 6256
rect 768 6224 800 6256
rect 840 6224 872 6256
rect 912 6224 944 6256
rect 984 6224 1016 6256
rect 1056 6224 1088 6256
rect 1128 6224 1160 6256
rect 1200 6224 1232 6256
rect 1272 6224 1304 6256
rect 1344 6224 1376 6256
rect 1416 6224 1448 6256
rect 1488 6224 1520 6256
rect 1560 6224 1592 6256
rect 1632 6224 1664 6256
rect 1704 6224 1736 6256
rect 1776 6224 1808 6256
rect 1848 6224 1880 6256
rect 1920 6224 1952 6256
rect 48 6152 80 6184
rect 120 6152 152 6184
rect 192 6152 224 6184
rect 264 6152 296 6184
rect 336 6152 368 6184
rect 408 6152 440 6184
rect 480 6152 512 6184
rect 552 6152 584 6184
rect 624 6152 656 6184
rect 696 6152 728 6184
rect 768 6152 800 6184
rect 840 6152 872 6184
rect 912 6152 944 6184
rect 984 6152 1016 6184
rect 1056 6152 1088 6184
rect 1128 6152 1160 6184
rect 1200 6152 1232 6184
rect 1272 6152 1304 6184
rect 1344 6152 1376 6184
rect 1416 6152 1448 6184
rect 1488 6152 1520 6184
rect 1560 6152 1592 6184
rect 1632 6152 1664 6184
rect 1704 6152 1736 6184
rect 1776 6152 1808 6184
rect 1848 6152 1880 6184
rect 1920 6152 1952 6184
rect 48 6080 80 6112
rect 120 6080 152 6112
rect 192 6080 224 6112
rect 264 6080 296 6112
rect 336 6080 368 6112
rect 408 6080 440 6112
rect 480 6080 512 6112
rect 552 6080 584 6112
rect 624 6080 656 6112
rect 696 6080 728 6112
rect 768 6080 800 6112
rect 840 6080 872 6112
rect 912 6080 944 6112
rect 984 6080 1016 6112
rect 1056 6080 1088 6112
rect 1128 6080 1160 6112
rect 1200 6080 1232 6112
rect 1272 6080 1304 6112
rect 1344 6080 1376 6112
rect 1416 6080 1448 6112
rect 1488 6080 1520 6112
rect 1560 6080 1592 6112
rect 1632 6080 1664 6112
rect 1704 6080 1736 6112
rect 1776 6080 1808 6112
rect 1848 6080 1880 6112
rect 1920 6080 1952 6112
rect 48 6008 80 6040
rect 120 6008 152 6040
rect 192 6008 224 6040
rect 264 6008 296 6040
rect 336 6008 368 6040
rect 408 6008 440 6040
rect 480 6008 512 6040
rect 552 6008 584 6040
rect 624 6008 656 6040
rect 696 6008 728 6040
rect 768 6008 800 6040
rect 840 6008 872 6040
rect 912 6008 944 6040
rect 984 6008 1016 6040
rect 1056 6008 1088 6040
rect 1128 6008 1160 6040
rect 1200 6008 1232 6040
rect 1272 6008 1304 6040
rect 1344 6008 1376 6040
rect 1416 6008 1448 6040
rect 1488 6008 1520 6040
rect 1560 6008 1592 6040
rect 1632 6008 1664 6040
rect 1704 6008 1736 6040
rect 1776 6008 1808 6040
rect 1848 6008 1880 6040
rect 1920 6008 1952 6040
rect 48 5936 80 5968
rect 120 5936 152 5968
rect 192 5936 224 5968
rect 264 5936 296 5968
rect 336 5936 368 5968
rect 408 5936 440 5968
rect 480 5936 512 5968
rect 552 5936 584 5968
rect 624 5936 656 5968
rect 696 5936 728 5968
rect 768 5936 800 5968
rect 840 5936 872 5968
rect 912 5936 944 5968
rect 984 5936 1016 5968
rect 1056 5936 1088 5968
rect 1128 5936 1160 5968
rect 1200 5936 1232 5968
rect 1272 5936 1304 5968
rect 1344 5936 1376 5968
rect 1416 5936 1448 5968
rect 1488 5936 1520 5968
rect 1560 5936 1592 5968
rect 1632 5936 1664 5968
rect 1704 5936 1736 5968
rect 1776 5936 1808 5968
rect 1848 5936 1880 5968
rect 1920 5936 1952 5968
rect 48 5864 80 5896
rect 120 5864 152 5896
rect 192 5864 224 5896
rect 264 5864 296 5896
rect 336 5864 368 5896
rect 408 5864 440 5896
rect 480 5864 512 5896
rect 552 5864 584 5896
rect 624 5864 656 5896
rect 696 5864 728 5896
rect 768 5864 800 5896
rect 840 5864 872 5896
rect 912 5864 944 5896
rect 984 5864 1016 5896
rect 1056 5864 1088 5896
rect 1128 5864 1160 5896
rect 1200 5864 1232 5896
rect 1272 5864 1304 5896
rect 1344 5864 1376 5896
rect 1416 5864 1448 5896
rect 1488 5864 1520 5896
rect 1560 5864 1592 5896
rect 1632 5864 1664 5896
rect 1704 5864 1736 5896
rect 1776 5864 1808 5896
rect 1848 5864 1880 5896
rect 1920 5864 1952 5896
rect 48 5792 80 5824
rect 120 5792 152 5824
rect 192 5792 224 5824
rect 264 5792 296 5824
rect 336 5792 368 5824
rect 408 5792 440 5824
rect 480 5792 512 5824
rect 552 5792 584 5824
rect 624 5792 656 5824
rect 696 5792 728 5824
rect 768 5792 800 5824
rect 840 5792 872 5824
rect 912 5792 944 5824
rect 984 5792 1016 5824
rect 1056 5792 1088 5824
rect 1128 5792 1160 5824
rect 1200 5792 1232 5824
rect 1272 5792 1304 5824
rect 1344 5792 1376 5824
rect 1416 5792 1448 5824
rect 1488 5792 1520 5824
rect 1560 5792 1592 5824
rect 1632 5792 1664 5824
rect 1704 5792 1736 5824
rect 1776 5792 1808 5824
rect 1848 5792 1880 5824
rect 1920 5792 1952 5824
rect 48 5720 80 5752
rect 120 5720 152 5752
rect 192 5720 224 5752
rect 264 5720 296 5752
rect 336 5720 368 5752
rect 408 5720 440 5752
rect 480 5720 512 5752
rect 552 5720 584 5752
rect 624 5720 656 5752
rect 696 5720 728 5752
rect 768 5720 800 5752
rect 840 5720 872 5752
rect 912 5720 944 5752
rect 984 5720 1016 5752
rect 1056 5720 1088 5752
rect 1128 5720 1160 5752
rect 1200 5720 1232 5752
rect 1272 5720 1304 5752
rect 1344 5720 1376 5752
rect 1416 5720 1448 5752
rect 1488 5720 1520 5752
rect 1560 5720 1592 5752
rect 1632 5720 1664 5752
rect 1704 5720 1736 5752
rect 1776 5720 1808 5752
rect 1848 5720 1880 5752
rect 1920 5720 1952 5752
rect 48 5648 80 5680
rect 120 5648 152 5680
rect 192 5648 224 5680
rect 264 5648 296 5680
rect 336 5648 368 5680
rect 408 5648 440 5680
rect 480 5648 512 5680
rect 552 5648 584 5680
rect 624 5648 656 5680
rect 696 5648 728 5680
rect 768 5648 800 5680
rect 840 5648 872 5680
rect 912 5648 944 5680
rect 984 5648 1016 5680
rect 1056 5648 1088 5680
rect 1128 5648 1160 5680
rect 1200 5648 1232 5680
rect 1272 5648 1304 5680
rect 1344 5648 1376 5680
rect 1416 5648 1448 5680
rect 1488 5648 1520 5680
rect 1560 5648 1592 5680
rect 1632 5648 1664 5680
rect 1704 5648 1736 5680
rect 1776 5648 1808 5680
rect 1848 5648 1880 5680
rect 1920 5648 1952 5680
rect 48 5576 80 5608
rect 120 5576 152 5608
rect 192 5576 224 5608
rect 264 5576 296 5608
rect 336 5576 368 5608
rect 408 5576 440 5608
rect 480 5576 512 5608
rect 552 5576 584 5608
rect 624 5576 656 5608
rect 696 5576 728 5608
rect 768 5576 800 5608
rect 840 5576 872 5608
rect 912 5576 944 5608
rect 984 5576 1016 5608
rect 1056 5576 1088 5608
rect 1128 5576 1160 5608
rect 1200 5576 1232 5608
rect 1272 5576 1304 5608
rect 1344 5576 1376 5608
rect 1416 5576 1448 5608
rect 1488 5576 1520 5608
rect 1560 5576 1592 5608
rect 1632 5576 1664 5608
rect 1704 5576 1736 5608
rect 1776 5576 1808 5608
rect 1848 5576 1880 5608
rect 1920 5576 1952 5608
rect 48 5504 80 5536
rect 120 5504 152 5536
rect 192 5504 224 5536
rect 264 5504 296 5536
rect 336 5504 368 5536
rect 408 5504 440 5536
rect 480 5504 512 5536
rect 552 5504 584 5536
rect 624 5504 656 5536
rect 696 5504 728 5536
rect 768 5504 800 5536
rect 840 5504 872 5536
rect 912 5504 944 5536
rect 984 5504 1016 5536
rect 1056 5504 1088 5536
rect 1128 5504 1160 5536
rect 1200 5504 1232 5536
rect 1272 5504 1304 5536
rect 1344 5504 1376 5536
rect 1416 5504 1448 5536
rect 1488 5504 1520 5536
rect 1560 5504 1592 5536
rect 1632 5504 1664 5536
rect 1704 5504 1736 5536
rect 1776 5504 1808 5536
rect 1848 5504 1880 5536
rect 1920 5504 1952 5536
rect 48 5432 80 5464
rect 120 5432 152 5464
rect 192 5432 224 5464
rect 264 5432 296 5464
rect 336 5432 368 5464
rect 408 5432 440 5464
rect 480 5432 512 5464
rect 552 5432 584 5464
rect 624 5432 656 5464
rect 696 5432 728 5464
rect 768 5432 800 5464
rect 840 5432 872 5464
rect 912 5432 944 5464
rect 984 5432 1016 5464
rect 1056 5432 1088 5464
rect 1128 5432 1160 5464
rect 1200 5432 1232 5464
rect 1272 5432 1304 5464
rect 1344 5432 1376 5464
rect 1416 5432 1448 5464
rect 1488 5432 1520 5464
rect 1560 5432 1592 5464
rect 1632 5432 1664 5464
rect 1704 5432 1736 5464
rect 1776 5432 1808 5464
rect 1848 5432 1880 5464
rect 1920 5432 1952 5464
rect 48 5360 80 5392
rect 120 5360 152 5392
rect 192 5360 224 5392
rect 264 5360 296 5392
rect 336 5360 368 5392
rect 408 5360 440 5392
rect 480 5360 512 5392
rect 552 5360 584 5392
rect 624 5360 656 5392
rect 696 5360 728 5392
rect 768 5360 800 5392
rect 840 5360 872 5392
rect 912 5360 944 5392
rect 984 5360 1016 5392
rect 1056 5360 1088 5392
rect 1128 5360 1160 5392
rect 1200 5360 1232 5392
rect 1272 5360 1304 5392
rect 1344 5360 1376 5392
rect 1416 5360 1448 5392
rect 1488 5360 1520 5392
rect 1560 5360 1592 5392
rect 1632 5360 1664 5392
rect 1704 5360 1736 5392
rect 1776 5360 1808 5392
rect 1848 5360 1880 5392
rect 1920 5360 1952 5392
rect 48 5288 80 5320
rect 120 5288 152 5320
rect 192 5288 224 5320
rect 264 5288 296 5320
rect 336 5288 368 5320
rect 408 5288 440 5320
rect 480 5288 512 5320
rect 552 5288 584 5320
rect 624 5288 656 5320
rect 696 5288 728 5320
rect 768 5288 800 5320
rect 840 5288 872 5320
rect 912 5288 944 5320
rect 984 5288 1016 5320
rect 1056 5288 1088 5320
rect 1128 5288 1160 5320
rect 1200 5288 1232 5320
rect 1272 5288 1304 5320
rect 1344 5288 1376 5320
rect 1416 5288 1448 5320
rect 1488 5288 1520 5320
rect 1560 5288 1592 5320
rect 1632 5288 1664 5320
rect 1704 5288 1736 5320
rect 1776 5288 1808 5320
rect 1848 5288 1880 5320
rect 1920 5288 1952 5320
rect 48 5216 80 5248
rect 120 5216 152 5248
rect 192 5216 224 5248
rect 264 5216 296 5248
rect 336 5216 368 5248
rect 408 5216 440 5248
rect 480 5216 512 5248
rect 552 5216 584 5248
rect 624 5216 656 5248
rect 696 5216 728 5248
rect 768 5216 800 5248
rect 840 5216 872 5248
rect 912 5216 944 5248
rect 984 5216 1016 5248
rect 1056 5216 1088 5248
rect 1128 5216 1160 5248
rect 1200 5216 1232 5248
rect 1272 5216 1304 5248
rect 1344 5216 1376 5248
rect 1416 5216 1448 5248
rect 1488 5216 1520 5248
rect 1560 5216 1592 5248
rect 1632 5216 1664 5248
rect 1704 5216 1736 5248
rect 1776 5216 1808 5248
rect 1848 5216 1880 5248
rect 1920 5216 1952 5248
rect 48 5144 80 5176
rect 120 5144 152 5176
rect 192 5144 224 5176
rect 264 5144 296 5176
rect 336 5144 368 5176
rect 408 5144 440 5176
rect 480 5144 512 5176
rect 552 5144 584 5176
rect 624 5144 656 5176
rect 696 5144 728 5176
rect 768 5144 800 5176
rect 840 5144 872 5176
rect 912 5144 944 5176
rect 984 5144 1016 5176
rect 1056 5144 1088 5176
rect 1128 5144 1160 5176
rect 1200 5144 1232 5176
rect 1272 5144 1304 5176
rect 1344 5144 1376 5176
rect 1416 5144 1448 5176
rect 1488 5144 1520 5176
rect 1560 5144 1592 5176
rect 1632 5144 1664 5176
rect 1704 5144 1736 5176
rect 1776 5144 1808 5176
rect 1848 5144 1880 5176
rect 1920 5144 1952 5176
rect 48 5072 80 5104
rect 120 5072 152 5104
rect 192 5072 224 5104
rect 264 5072 296 5104
rect 336 5072 368 5104
rect 408 5072 440 5104
rect 480 5072 512 5104
rect 552 5072 584 5104
rect 624 5072 656 5104
rect 696 5072 728 5104
rect 768 5072 800 5104
rect 840 5072 872 5104
rect 912 5072 944 5104
rect 984 5072 1016 5104
rect 1056 5072 1088 5104
rect 1128 5072 1160 5104
rect 1200 5072 1232 5104
rect 1272 5072 1304 5104
rect 1344 5072 1376 5104
rect 1416 5072 1448 5104
rect 1488 5072 1520 5104
rect 1560 5072 1592 5104
rect 1632 5072 1664 5104
rect 1704 5072 1736 5104
rect 1776 5072 1808 5104
rect 1848 5072 1880 5104
rect 1920 5072 1952 5104
rect 48 5000 80 5032
rect 120 5000 152 5032
rect 192 5000 224 5032
rect 264 5000 296 5032
rect 336 5000 368 5032
rect 408 5000 440 5032
rect 480 5000 512 5032
rect 552 5000 584 5032
rect 624 5000 656 5032
rect 696 5000 728 5032
rect 768 5000 800 5032
rect 840 5000 872 5032
rect 912 5000 944 5032
rect 984 5000 1016 5032
rect 1056 5000 1088 5032
rect 1128 5000 1160 5032
rect 1200 5000 1232 5032
rect 1272 5000 1304 5032
rect 1344 5000 1376 5032
rect 1416 5000 1448 5032
rect 1488 5000 1520 5032
rect 1560 5000 1592 5032
rect 1632 5000 1664 5032
rect 1704 5000 1736 5032
rect 1776 5000 1808 5032
rect 1848 5000 1880 5032
rect 1920 5000 1952 5032
rect 48 4928 80 4960
rect 120 4928 152 4960
rect 192 4928 224 4960
rect 264 4928 296 4960
rect 336 4928 368 4960
rect 408 4928 440 4960
rect 480 4928 512 4960
rect 552 4928 584 4960
rect 624 4928 656 4960
rect 696 4928 728 4960
rect 768 4928 800 4960
rect 840 4928 872 4960
rect 912 4928 944 4960
rect 984 4928 1016 4960
rect 1056 4928 1088 4960
rect 1128 4928 1160 4960
rect 1200 4928 1232 4960
rect 1272 4928 1304 4960
rect 1344 4928 1376 4960
rect 1416 4928 1448 4960
rect 1488 4928 1520 4960
rect 1560 4928 1592 4960
rect 1632 4928 1664 4960
rect 1704 4928 1736 4960
rect 1776 4928 1808 4960
rect 1848 4928 1880 4960
rect 1920 4928 1952 4960
rect 48 4856 80 4888
rect 120 4856 152 4888
rect 192 4856 224 4888
rect 264 4856 296 4888
rect 336 4856 368 4888
rect 408 4856 440 4888
rect 480 4856 512 4888
rect 552 4856 584 4888
rect 624 4856 656 4888
rect 696 4856 728 4888
rect 768 4856 800 4888
rect 840 4856 872 4888
rect 912 4856 944 4888
rect 984 4856 1016 4888
rect 1056 4856 1088 4888
rect 1128 4856 1160 4888
rect 1200 4856 1232 4888
rect 1272 4856 1304 4888
rect 1344 4856 1376 4888
rect 1416 4856 1448 4888
rect 1488 4856 1520 4888
rect 1560 4856 1592 4888
rect 1632 4856 1664 4888
rect 1704 4856 1736 4888
rect 1776 4856 1808 4888
rect 1848 4856 1880 4888
rect 1920 4856 1952 4888
rect 48 4784 80 4816
rect 120 4784 152 4816
rect 192 4784 224 4816
rect 264 4784 296 4816
rect 336 4784 368 4816
rect 408 4784 440 4816
rect 480 4784 512 4816
rect 552 4784 584 4816
rect 624 4784 656 4816
rect 696 4784 728 4816
rect 768 4784 800 4816
rect 840 4784 872 4816
rect 912 4784 944 4816
rect 984 4784 1016 4816
rect 1056 4784 1088 4816
rect 1128 4784 1160 4816
rect 1200 4784 1232 4816
rect 1272 4784 1304 4816
rect 1344 4784 1376 4816
rect 1416 4784 1448 4816
rect 1488 4784 1520 4816
rect 1560 4784 1592 4816
rect 1632 4784 1664 4816
rect 1704 4784 1736 4816
rect 1776 4784 1808 4816
rect 1848 4784 1880 4816
rect 1920 4784 1952 4816
rect 48 4712 80 4744
rect 120 4712 152 4744
rect 192 4712 224 4744
rect 264 4712 296 4744
rect 336 4712 368 4744
rect 408 4712 440 4744
rect 480 4712 512 4744
rect 552 4712 584 4744
rect 624 4712 656 4744
rect 696 4712 728 4744
rect 768 4712 800 4744
rect 840 4712 872 4744
rect 912 4712 944 4744
rect 984 4712 1016 4744
rect 1056 4712 1088 4744
rect 1128 4712 1160 4744
rect 1200 4712 1232 4744
rect 1272 4712 1304 4744
rect 1344 4712 1376 4744
rect 1416 4712 1448 4744
rect 1488 4712 1520 4744
rect 1560 4712 1592 4744
rect 1632 4712 1664 4744
rect 1704 4712 1736 4744
rect 1776 4712 1808 4744
rect 1848 4712 1880 4744
rect 1920 4712 1952 4744
rect 48 4640 80 4672
rect 120 4640 152 4672
rect 192 4640 224 4672
rect 264 4640 296 4672
rect 336 4640 368 4672
rect 408 4640 440 4672
rect 480 4640 512 4672
rect 552 4640 584 4672
rect 624 4640 656 4672
rect 696 4640 728 4672
rect 768 4640 800 4672
rect 840 4640 872 4672
rect 912 4640 944 4672
rect 984 4640 1016 4672
rect 1056 4640 1088 4672
rect 1128 4640 1160 4672
rect 1200 4640 1232 4672
rect 1272 4640 1304 4672
rect 1344 4640 1376 4672
rect 1416 4640 1448 4672
rect 1488 4640 1520 4672
rect 1560 4640 1592 4672
rect 1632 4640 1664 4672
rect 1704 4640 1736 4672
rect 1776 4640 1808 4672
rect 1848 4640 1880 4672
rect 1920 4640 1952 4672
rect 48 4568 80 4600
rect 120 4568 152 4600
rect 192 4568 224 4600
rect 264 4568 296 4600
rect 336 4568 368 4600
rect 408 4568 440 4600
rect 480 4568 512 4600
rect 552 4568 584 4600
rect 624 4568 656 4600
rect 696 4568 728 4600
rect 768 4568 800 4600
rect 840 4568 872 4600
rect 912 4568 944 4600
rect 984 4568 1016 4600
rect 1056 4568 1088 4600
rect 1128 4568 1160 4600
rect 1200 4568 1232 4600
rect 1272 4568 1304 4600
rect 1344 4568 1376 4600
rect 1416 4568 1448 4600
rect 1488 4568 1520 4600
rect 1560 4568 1592 4600
rect 1632 4568 1664 4600
rect 1704 4568 1736 4600
rect 1776 4568 1808 4600
rect 1848 4568 1880 4600
rect 1920 4568 1952 4600
rect 48 4496 80 4528
rect 120 4496 152 4528
rect 192 4496 224 4528
rect 264 4496 296 4528
rect 336 4496 368 4528
rect 408 4496 440 4528
rect 480 4496 512 4528
rect 552 4496 584 4528
rect 624 4496 656 4528
rect 696 4496 728 4528
rect 768 4496 800 4528
rect 840 4496 872 4528
rect 912 4496 944 4528
rect 984 4496 1016 4528
rect 1056 4496 1088 4528
rect 1128 4496 1160 4528
rect 1200 4496 1232 4528
rect 1272 4496 1304 4528
rect 1344 4496 1376 4528
rect 1416 4496 1448 4528
rect 1488 4496 1520 4528
rect 1560 4496 1592 4528
rect 1632 4496 1664 4528
rect 1704 4496 1736 4528
rect 1776 4496 1808 4528
rect 1848 4496 1880 4528
rect 1920 4496 1952 4528
rect 48 4424 80 4456
rect 120 4424 152 4456
rect 192 4424 224 4456
rect 264 4424 296 4456
rect 336 4424 368 4456
rect 408 4424 440 4456
rect 480 4424 512 4456
rect 552 4424 584 4456
rect 624 4424 656 4456
rect 696 4424 728 4456
rect 768 4424 800 4456
rect 840 4424 872 4456
rect 912 4424 944 4456
rect 984 4424 1016 4456
rect 1056 4424 1088 4456
rect 1128 4424 1160 4456
rect 1200 4424 1232 4456
rect 1272 4424 1304 4456
rect 1344 4424 1376 4456
rect 1416 4424 1448 4456
rect 1488 4424 1520 4456
rect 1560 4424 1592 4456
rect 1632 4424 1664 4456
rect 1704 4424 1736 4456
rect 1776 4424 1808 4456
rect 1848 4424 1880 4456
rect 1920 4424 1952 4456
rect 48 4352 80 4384
rect 120 4352 152 4384
rect 192 4352 224 4384
rect 264 4352 296 4384
rect 336 4352 368 4384
rect 408 4352 440 4384
rect 480 4352 512 4384
rect 552 4352 584 4384
rect 624 4352 656 4384
rect 696 4352 728 4384
rect 768 4352 800 4384
rect 840 4352 872 4384
rect 912 4352 944 4384
rect 984 4352 1016 4384
rect 1056 4352 1088 4384
rect 1128 4352 1160 4384
rect 1200 4352 1232 4384
rect 1272 4352 1304 4384
rect 1344 4352 1376 4384
rect 1416 4352 1448 4384
rect 1488 4352 1520 4384
rect 1560 4352 1592 4384
rect 1632 4352 1664 4384
rect 1704 4352 1736 4384
rect 1776 4352 1808 4384
rect 1848 4352 1880 4384
rect 1920 4352 1952 4384
rect 48 4280 80 4312
rect 120 4280 152 4312
rect 192 4280 224 4312
rect 264 4280 296 4312
rect 336 4280 368 4312
rect 408 4280 440 4312
rect 480 4280 512 4312
rect 552 4280 584 4312
rect 624 4280 656 4312
rect 696 4280 728 4312
rect 768 4280 800 4312
rect 840 4280 872 4312
rect 912 4280 944 4312
rect 984 4280 1016 4312
rect 1056 4280 1088 4312
rect 1128 4280 1160 4312
rect 1200 4280 1232 4312
rect 1272 4280 1304 4312
rect 1344 4280 1376 4312
rect 1416 4280 1448 4312
rect 1488 4280 1520 4312
rect 1560 4280 1592 4312
rect 1632 4280 1664 4312
rect 1704 4280 1736 4312
rect 1776 4280 1808 4312
rect 1848 4280 1880 4312
rect 1920 4280 1952 4312
rect 48 4208 80 4240
rect 120 4208 152 4240
rect 192 4208 224 4240
rect 264 4208 296 4240
rect 336 4208 368 4240
rect 408 4208 440 4240
rect 480 4208 512 4240
rect 552 4208 584 4240
rect 624 4208 656 4240
rect 696 4208 728 4240
rect 768 4208 800 4240
rect 840 4208 872 4240
rect 912 4208 944 4240
rect 984 4208 1016 4240
rect 1056 4208 1088 4240
rect 1128 4208 1160 4240
rect 1200 4208 1232 4240
rect 1272 4208 1304 4240
rect 1344 4208 1376 4240
rect 1416 4208 1448 4240
rect 1488 4208 1520 4240
rect 1560 4208 1592 4240
rect 1632 4208 1664 4240
rect 1704 4208 1736 4240
rect 1776 4208 1808 4240
rect 1848 4208 1880 4240
rect 1920 4208 1952 4240
rect 48 4136 80 4168
rect 120 4136 152 4168
rect 192 4136 224 4168
rect 264 4136 296 4168
rect 336 4136 368 4168
rect 408 4136 440 4168
rect 480 4136 512 4168
rect 552 4136 584 4168
rect 624 4136 656 4168
rect 696 4136 728 4168
rect 768 4136 800 4168
rect 840 4136 872 4168
rect 912 4136 944 4168
rect 984 4136 1016 4168
rect 1056 4136 1088 4168
rect 1128 4136 1160 4168
rect 1200 4136 1232 4168
rect 1272 4136 1304 4168
rect 1344 4136 1376 4168
rect 1416 4136 1448 4168
rect 1488 4136 1520 4168
rect 1560 4136 1592 4168
rect 1632 4136 1664 4168
rect 1704 4136 1736 4168
rect 1776 4136 1808 4168
rect 1848 4136 1880 4168
rect 1920 4136 1952 4168
rect 48 4064 80 4096
rect 120 4064 152 4096
rect 192 4064 224 4096
rect 264 4064 296 4096
rect 336 4064 368 4096
rect 408 4064 440 4096
rect 480 4064 512 4096
rect 552 4064 584 4096
rect 624 4064 656 4096
rect 696 4064 728 4096
rect 768 4064 800 4096
rect 840 4064 872 4096
rect 912 4064 944 4096
rect 984 4064 1016 4096
rect 1056 4064 1088 4096
rect 1128 4064 1160 4096
rect 1200 4064 1232 4096
rect 1272 4064 1304 4096
rect 1344 4064 1376 4096
rect 1416 4064 1448 4096
rect 1488 4064 1520 4096
rect 1560 4064 1592 4096
rect 1632 4064 1664 4096
rect 1704 4064 1736 4096
rect 1776 4064 1808 4096
rect 1848 4064 1880 4096
rect 1920 4064 1952 4096
rect 48 3992 80 4024
rect 120 3992 152 4024
rect 192 3992 224 4024
rect 264 3992 296 4024
rect 336 3992 368 4024
rect 408 3992 440 4024
rect 480 3992 512 4024
rect 552 3992 584 4024
rect 624 3992 656 4024
rect 696 3992 728 4024
rect 768 3992 800 4024
rect 840 3992 872 4024
rect 912 3992 944 4024
rect 984 3992 1016 4024
rect 1056 3992 1088 4024
rect 1128 3992 1160 4024
rect 1200 3992 1232 4024
rect 1272 3992 1304 4024
rect 1344 3992 1376 4024
rect 1416 3992 1448 4024
rect 1488 3992 1520 4024
rect 1560 3992 1592 4024
rect 1632 3992 1664 4024
rect 1704 3992 1736 4024
rect 1776 3992 1808 4024
rect 1848 3992 1880 4024
rect 1920 3992 1952 4024
rect 48 3920 80 3952
rect 120 3920 152 3952
rect 192 3920 224 3952
rect 264 3920 296 3952
rect 336 3920 368 3952
rect 408 3920 440 3952
rect 480 3920 512 3952
rect 552 3920 584 3952
rect 624 3920 656 3952
rect 696 3920 728 3952
rect 768 3920 800 3952
rect 840 3920 872 3952
rect 912 3920 944 3952
rect 984 3920 1016 3952
rect 1056 3920 1088 3952
rect 1128 3920 1160 3952
rect 1200 3920 1232 3952
rect 1272 3920 1304 3952
rect 1344 3920 1376 3952
rect 1416 3920 1448 3952
rect 1488 3920 1520 3952
rect 1560 3920 1592 3952
rect 1632 3920 1664 3952
rect 1704 3920 1736 3952
rect 1776 3920 1808 3952
rect 1848 3920 1880 3952
rect 1920 3920 1952 3952
rect 48 3848 80 3880
rect 120 3848 152 3880
rect 192 3848 224 3880
rect 264 3848 296 3880
rect 336 3848 368 3880
rect 408 3848 440 3880
rect 480 3848 512 3880
rect 552 3848 584 3880
rect 624 3848 656 3880
rect 696 3848 728 3880
rect 768 3848 800 3880
rect 840 3848 872 3880
rect 912 3848 944 3880
rect 984 3848 1016 3880
rect 1056 3848 1088 3880
rect 1128 3848 1160 3880
rect 1200 3848 1232 3880
rect 1272 3848 1304 3880
rect 1344 3848 1376 3880
rect 1416 3848 1448 3880
rect 1488 3848 1520 3880
rect 1560 3848 1592 3880
rect 1632 3848 1664 3880
rect 1704 3848 1736 3880
rect 1776 3848 1808 3880
rect 1848 3848 1880 3880
rect 1920 3848 1952 3880
rect 48 3776 80 3808
rect 120 3776 152 3808
rect 192 3776 224 3808
rect 264 3776 296 3808
rect 336 3776 368 3808
rect 408 3776 440 3808
rect 480 3776 512 3808
rect 552 3776 584 3808
rect 624 3776 656 3808
rect 696 3776 728 3808
rect 768 3776 800 3808
rect 840 3776 872 3808
rect 912 3776 944 3808
rect 984 3776 1016 3808
rect 1056 3776 1088 3808
rect 1128 3776 1160 3808
rect 1200 3776 1232 3808
rect 1272 3776 1304 3808
rect 1344 3776 1376 3808
rect 1416 3776 1448 3808
rect 1488 3776 1520 3808
rect 1560 3776 1592 3808
rect 1632 3776 1664 3808
rect 1704 3776 1736 3808
rect 1776 3776 1808 3808
rect 1848 3776 1880 3808
rect 1920 3776 1952 3808
rect 48 3704 80 3736
rect 120 3704 152 3736
rect 192 3704 224 3736
rect 264 3704 296 3736
rect 336 3704 368 3736
rect 408 3704 440 3736
rect 480 3704 512 3736
rect 552 3704 584 3736
rect 624 3704 656 3736
rect 696 3704 728 3736
rect 768 3704 800 3736
rect 840 3704 872 3736
rect 912 3704 944 3736
rect 984 3704 1016 3736
rect 1056 3704 1088 3736
rect 1128 3704 1160 3736
rect 1200 3704 1232 3736
rect 1272 3704 1304 3736
rect 1344 3704 1376 3736
rect 1416 3704 1448 3736
rect 1488 3704 1520 3736
rect 1560 3704 1592 3736
rect 1632 3704 1664 3736
rect 1704 3704 1736 3736
rect 1776 3704 1808 3736
rect 1848 3704 1880 3736
rect 1920 3704 1952 3736
rect 48 3632 80 3664
rect 120 3632 152 3664
rect 192 3632 224 3664
rect 264 3632 296 3664
rect 336 3632 368 3664
rect 408 3632 440 3664
rect 480 3632 512 3664
rect 552 3632 584 3664
rect 624 3632 656 3664
rect 696 3632 728 3664
rect 768 3632 800 3664
rect 840 3632 872 3664
rect 912 3632 944 3664
rect 984 3632 1016 3664
rect 1056 3632 1088 3664
rect 1128 3632 1160 3664
rect 1200 3632 1232 3664
rect 1272 3632 1304 3664
rect 1344 3632 1376 3664
rect 1416 3632 1448 3664
rect 1488 3632 1520 3664
rect 1560 3632 1592 3664
rect 1632 3632 1664 3664
rect 1704 3632 1736 3664
rect 1776 3632 1808 3664
rect 1848 3632 1880 3664
rect 1920 3632 1952 3664
rect 48 3560 80 3592
rect 120 3560 152 3592
rect 192 3560 224 3592
rect 264 3560 296 3592
rect 336 3560 368 3592
rect 408 3560 440 3592
rect 480 3560 512 3592
rect 552 3560 584 3592
rect 624 3560 656 3592
rect 696 3560 728 3592
rect 768 3560 800 3592
rect 840 3560 872 3592
rect 912 3560 944 3592
rect 984 3560 1016 3592
rect 1056 3560 1088 3592
rect 1128 3560 1160 3592
rect 1200 3560 1232 3592
rect 1272 3560 1304 3592
rect 1344 3560 1376 3592
rect 1416 3560 1448 3592
rect 1488 3560 1520 3592
rect 1560 3560 1592 3592
rect 1632 3560 1664 3592
rect 1704 3560 1736 3592
rect 1776 3560 1808 3592
rect 1848 3560 1880 3592
rect 1920 3560 1952 3592
rect 48 3488 80 3520
rect 120 3488 152 3520
rect 192 3488 224 3520
rect 264 3488 296 3520
rect 336 3488 368 3520
rect 408 3488 440 3520
rect 480 3488 512 3520
rect 552 3488 584 3520
rect 624 3488 656 3520
rect 696 3488 728 3520
rect 768 3488 800 3520
rect 840 3488 872 3520
rect 912 3488 944 3520
rect 984 3488 1016 3520
rect 1056 3488 1088 3520
rect 1128 3488 1160 3520
rect 1200 3488 1232 3520
rect 1272 3488 1304 3520
rect 1344 3488 1376 3520
rect 1416 3488 1448 3520
rect 1488 3488 1520 3520
rect 1560 3488 1592 3520
rect 1632 3488 1664 3520
rect 1704 3488 1736 3520
rect 1776 3488 1808 3520
rect 1848 3488 1880 3520
rect 1920 3488 1952 3520
rect 48 3416 80 3448
rect 120 3416 152 3448
rect 192 3416 224 3448
rect 264 3416 296 3448
rect 336 3416 368 3448
rect 408 3416 440 3448
rect 480 3416 512 3448
rect 552 3416 584 3448
rect 624 3416 656 3448
rect 696 3416 728 3448
rect 768 3416 800 3448
rect 840 3416 872 3448
rect 912 3416 944 3448
rect 984 3416 1016 3448
rect 1056 3416 1088 3448
rect 1128 3416 1160 3448
rect 1200 3416 1232 3448
rect 1272 3416 1304 3448
rect 1344 3416 1376 3448
rect 1416 3416 1448 3448
rect 1488 3416 1520 3448
rect 1560 3416 1592 3448
rect 1632 3416 1664 3448
rect 1704 3416 1736 3448
rect 1776 3416 1808 3448
rect 1848 3416 1880 3448
rect 1920 3416 1952 3448
rect 48 3344 80 3376
rect 120 3344 152 3376
rect 192 3344 224 3376
rect 264 3344 296 3376
rect 336 3344 368 3376
rect 408 3344 440 3376
rect 480 3344 512 3376
rect 552 3344 584 3376
rect 624 3344 656 3376
rect 696 3344 728 3376
rect 768 3344 800 3376
rect 840 3344 872 3376
rect 912 3344 944 3376
rect 984 3344 1016 3376
rect 1056 3344 1088 3376
rect 1128 3344 1160 3376
rect 1200 3344 1232 3376
rect 1272 3344 1304 3376
rect 1344 3344 1376 3376
rect 1416 3344 1448 3376
rect 1488 3344 1520 3376
rect 1560 3344 1592 3376
rect 1632 3344 1664 3376
rect 1704 3344 1736 3376
rect 1776 3344 1808 3376
rect 1848 3344 1880 3376
rect 1920 3344 1952 3376
rect 48 3272 80 3304
rect 120 3272 152 3304
rect 192 3272 224 3304
rect 264 3272 296 3304
rect 336 3272 368 3304
rect 408 3272 440 3304
rect 480 3272 512 3304
rect 552 3272 584 3304
rect 624 3272 656 3304
rect 696 3272 728 3304
rect 768 3272 800 3304
rect 840 3272 872 3304
rect 912 3272 944 3304
rect 984 3272 1016 3304
rect 1056 3272 1088 3304
rect 1128 3272 1160 3304
rect 1200 3272 1232 3304
rect 1272 3272 1304 3304
rect 1344 3272 1376 3304
rect 1416 3272 1448 3304
rect 1488 3272 1520 3304
rect 1560 3272 1592 3304
rect 1632 3272 1664 3304
rect 1704 3272 1736 3304
rect 1776 3272 1808 3304
rect 1848 3272 1880 3304
rect 1920 3272 1952 3304
rect 48 3200 80 3232
rect 120 3200 152 3232
rect 192 3200 224 3232
rect 264 3200 296 3232
rect 336 3200 368 3232
rect 408 3200 440 3232
rect 480 3200 512 3232
rect 552 3200 584 3232
rect 624 3200 656 3232
rect 696 3200 728 3232
rect 768 3200 800 3232
rect 840 3200 872 3232
rect 912 3200 944 3232
rect 984 3200 1016 3232
rect 1056 3200 1088 3232
rect 1128 3200 1160 3232
rect 1200 3200 1232 3232
rect 1272 3200 1304 3232
rect 1344 3200 1376 3232
rect 1416 3200 1448 3232
rect 1488 3200 1520 3232
rect 1560 3200 1592 3232
rect 1632 3200 1664 3232
rect 1704 3200 1736 3232
rect 1776 3200 1808 3232
rect 1848 3200 1880 3232
rect 1920 3200 1952 3232
rect 48 3128 80 3160
rect 120 3128 152 3160
rect 192 3128 224 3160
rect 264 3128 296 3160
rect 336 3128 368 3160
rect 408 3128 440 3160
rect 480 3128 512 3160
rect 552 3128 584 3160
rect 624 3128 656 3160
rect 696 3128 728 3160
rect 768 3128 800 3160
rect 840 3128 872 3160
rect 912 3128 944 3160
rect 984 3128 1016 3160
rect 1056 3128 1088 3160
rect 1128 3128 1160 3160
rect 1200 3128 1232 3160
rect 1272 3128 1304 3160
rect 1344 3128 1376 3160
rect 1416 3128 1448 3160
rect 1488 3128 1520 3160
rect 1560 3128 1592 3160
rect 1632 3128 1664 3160
rect 1704 3128 1736 3160
rect 1776 3128 1808 3160
rect 1848 3128 1880 3160
rect 1920 3128 1952 3160
rect 48 3056 80 3088
rect 120 3056 152 3088
rect 192 3056 224 3088
rect 264 3056 296 3088
rect 336 3056 368 3088
rect 408 3056 440 3088
rect 480 3056 512 3088
rect 552 3056 584 3088
rect 624 3056 656 3088
rect 696 3056 728 3088
rect 768 3056 800 3088
rect 840 3056 872 3088
rect 912 3056 944 3088
rect 984 3056 1016 3088
rect 1056 3056 1088 3088
rect 1128 3056 1160 3088
rect 1200 3056 1232 3088
rect 1272 3056 1304 3088
rect 1344 3056 1376 3088
rect 1416 3056 1448 3088
rect 1488 3056 1520 3088
rect 1560 3056 1592 3088
rect 1632 3056 1664 3088
rect 1704 3056 1736 3088
rect 1776 3056 1808 3088
rect 1848 3056 1880 3088
rect 1920 3056 1952 3088
rect 48 2984 80 3016
rect 120 2984 152 3016
rect 192 2984 224 3016
rect 264 2984 296 3016
rect 336 2984 368 3016
rect 408 2984 440 3016
rect 480 2984 512 3016
rect 552 2984 584 3016
rect 624 2984 656 3016
rect 696 2984 728 3016
rect 768 2984 800 3016
rect 840 2984 872 3016
rect 912 2984 944 3016
rect 984 2984 1016 3016
rect 1056 2984 1088 3016
rect 1128 2984 1160 3016
rect 1200 2984 1232 3016
rect 1272 2984 1304 3016
rect 1344 2984 1376 3016
rect 1416 2984 1448 3016
rect 1488 2984 1520 3016
rect 1560 2984 1592 3016
rect 1632 2984 1664 3016
rect 1704 2984 1736 3016
rect 1776 2984 1808 3016
rect 1848 2984 1880 3016
rect 1920 2984 1952 3016
rect 48 2912 80 2944
rect 120 2912 152 2944
rect 192 2912 224 2944
rect 264 2912 296 2944
rect 336 2912 368 2944
rect 408 2912 440 2944
rect 480 2912 512 2944
rect 552 2912 584 2944
rect 624 2912 656 2944
rect 696 2912 728 2944
rect 768 2912 800 2944
rect 840 2912 872 2944
rect 912 2912 944 2944
rect 984 2912 1016 2944
rect 1056 2912 1088 2944
rect 1128 2912 1160 2944
rect 1200 2912 1232 2944
rect 1272 2912 1304 2944
rect 1344 2912 1376 2944
rect 1416 2912 1448 2944
rect 1488 2912 1520 2944
rect 1560 2912 1592 2944
rect 1632 2912 1664 2944
rect 1704 2912 1736 2944
rect 1776 2912 1808 2944
rect 1848 2912 1880 2944
rect 1920 2912 1952 2944
rect 48 2840 80 2872
rect 120 2840 152 2872
rect 192 2840 224 2872
rect 264 2840 296 2872
rect 336 2840 368 2872
rect 408 2840 440 2872
rect 480 2840 512 2872
rect 552 2840 584 2872
rect 624 2840 656 2872
rect 696 2840 728 2872
rect 768 2840 800 2872
rect 840 2840 872 2872
rect 912 2840 944 2872
rect 984 2840 1016 2872
rect 1056 2840 1088 2872
rect 1128 2840 1160 2872
rect 1200 2840 1232 2872
rect 1272 2840 1304 2872
rect 1344 2840 1376 2872
rect 1416 2840 1448 2872
rect 1488 2840 1520 2872
rect 1560 2840 1592 2872
rect 1632 2840 1664 2872
rect 1704 2840 1736 2872
rect 1776 2840 1808 2872
rect 1848 2840 1880 2872
rect 1920 2840 1952 2872
rect 48 2768 80 2800
rect 120 2768 152 2800
rect 192 2768 224 2800
rect 264 2768 296 2800
rect 336 2768 368 2800
rect 408 2768 440 2800
rect 480 2768 512 2800
rect 552 2768 584 2800
rect 624 2768 656 2800
rect 696 2768 728 2800
rect 768 2768 800 2800
rect 840 2768 872 2800
rect 912 2768 944 2800
rect 984 2768 1016 2800
rect 1056 2768 1088 2800
rect 1128 2768 1160 2800
rect 1200 2768 1232 2800
rect 1272 2768 1304 2800
rect 1344 2768 1376 2800
rect 1416 2768 1448 2800
rect 1488 2768 1520 2800
rect 1560 2768 1592 2800
rect 1632 2768 1664 2800
rect 1704 2768 1736 2800
rect 1776 2768 1808 2800
rect 1848 2768 1880 2800
rect 1920 2768 1952 2800
rect 48 2696 80 2728
rect 120 2696 152 2728
rect 192 2696 224 2728
rect 264 2696 296 2728
rect 336 2696 368 2728
rect 408 2696 440 2728
rect 480 2696 512 2728
rect 552 2696 584 2728
rect 624 2696 656 2728
rect 696 2696 728 2728
rect 768 2696 800 2728
rect 840 2696 872 2728
rect 912 2696 944 2728
rect 984 2696 1016 2728
rect 1056 2696 1088 2728
rect 1128 2696 1160 2728
rect 1200 2696 1232 2728
rect 1272 2696 1304 2728
rect 1344 2696 1376 2728
rect 1416 2696 1448 2728
rect 1488 2696 1520 2728
rect 1560 2696 1592 2728
rect 1632 2696 1664 2728
rect 1704 2696 1736 2728
rect 1776 2696 1808 2728
rect 1848 2696 1880 2728
rect 1920 2696 1952 2728
rect 48 2624 80 2656
rect 120 2624 152 2656
rect 192 2624 224 2656
rect 264 2624 296 2656
rect 336 2624 368 2656
rect 408 2624 440 2656
rect 480 2624 512 2656
rect 552 2624 584 2656
rect 624 2624 656 2656
rect 696 2624 728 2656
rect 768 2624 800 2656
rect 840 2624 872 2656
rect 912 2624 944 2656
rect 984 2624 1016 2656
rect 1056 2624 1088 2656
rect 1128 2624 1160 2656
rect 1200 2624 1232 2656
rect 1272 2624 1304 2656
rect 1344 2624 1376 2656
rect 1416 2624 1448 2656
rect 1488 2624 1520 2656
rect 1560 2624 1592 2656
rect 1632 2624 1664 2656
rect 1704 2624 1736 2656
rect 1776 2624 1808 2656
rect 1848 2624 1880 2656
rect 1920 2624 1952 2656
rect 48 2552 80 2584
rect 120 2552 152 2584
rect 192 2552 224 2584
rect 264 2552 296 2584
rect 336 2552 368 2584
rect 408 2552 440 2584
rect 480 2552 512 2584
rect 552 2552 584 2584
rect 624 2552 656 2584
rect 696 2552 728 2584
rect 768 2552 800 2584
rect 840 2552 872 2584
rect 912 2552 944 2584
rect 984 2552 1016 2584
rect 1056 2552 1088 2584
rect 1128 2552 1160 2584
rect 1200 2552 1232 2584
rect 1272 2552 1304 2584
rect 1344 2552 1376 2584
rect 1416 2552 1448 2584
rect 1488 2552 1520 2584
rect 1560 2552 1592 2584
rect 1632 2552 1664 2584
rect 1704 2552 1736 2584
rect 1776 2552 1808 2584
rect 1848 2552 1880 2584
rect 1920 2552 1952 2584
rect 48 2480 80 2512
rect 120 2480 152 2512
rect 192 2480 224 2512
rect 264 2480 296 2512
rect 336 2480 368 2512
rect 408 2480 440 2512
rect 480 2480 512 2512
rect 552 2480 584 2512
rect 624 2480 656 2512
rect 696 2480 728 2512
rect 768 2480 800 2512
rect 840 2480 872 2512
rect 912 2480 944 2512
rect 984 2480 1016 2512
rect 1056 2480 1088 2512
rect 1128 2480 1160 2512
rect 1200 2480 1232 2512
rect 1272 2480 1304 2512
rect 1344 2480 1376 2512
rect 1416 2480 1448 2512
rect 1488 2480 1520 2512
rect 1560 2480 1592 2512
rect 1632 2480 1664 2512
rect 1704 2480 1736 2512
rect 1776 2480 1808 2512
rect 1848 2480 1880 2512
rect 1920 2480 1952 2512
rect 48 2408 80 2440
rect 120 2408 152 2440
rect 192 2408 224 2440
rect 264 2408 296 2440
rect 336 2408 368 2440
rect 408 2408 440 2440
rect 480 2408 512 2440
rect 552 2408 584 2440
rect 624 2408 656 2440
rect 696 2408 728 2440
rect 768 2408 800 2440
rect 840 2408 872 2440
rect 912 2408 944 2440
rect 984 2408 1016 2440
rect 1056 2408 1088 2440
rect 1128 2408 1160 2440
rect 1200 2408 1232 2440
rect 1272 2408 1304 2440
rect 1344 2408 1376 2440
rect 1416 2408 1448 2440
rect 1488 2408 1520 2440
rect 1560 2408 1592 2440
rect 1632 2408 1664 2440
rect 1704 2408 1736 2440
rect 1776 2408 1808 2440
rect 1848 2408 1880 2440
rect 1920 2408 1952 2440
rect 48 2336 80 2368
rect 120 2336 152 2368
rect 192 2336 224 2368
rect 264 2336 296 2368
rect 336 2336 368 2368
rect 408 2336 440 2368
rect 480 2336 512 2368
rect 552 2336 584 2368
rect 624 2336 656 2368
rect 696 2336 728 2368
rect 768 2336 800 2368
rect 840 2336 872 2368
rect 912 2336 944 2368
rect 984 2336 1016 2368
rect 1056 2336 1088 2368
rect 1128 2336 1160 2368
rect 1200 2336 1232 2368
rect 1272 2336 1304 2368
rect 1344 2336 1376 2368
rect 1416 2336 1448 2368
rect 1488 2336 1520 2368
rect 1560 2336 1592 2368
rect 1632 2336 1664 2368
rect 1704 2336 1736 2368
rect 1776 2336 1808 2368
rect 1848 2336 1880 2368
rect 1920 2336 1952 2368
rect 48 2264 80 2296
rect 120 2264 152 2296
rect 192 2264 224 2296
rect 264 2264 296 2296
rect 336 2264 368 2296
rect 408 2264 440 2296
rect 480 2264 512 2296
rect 552 2264 584 2296
rect 624 2264 656 2296
rect 696 2264 728 2296
rect 768 2264 800 2296
rect 840 2264 872 2296
rect 912 2264 944 2296
rect 984 2264 1016 2296
rect 1056 2264 1088 2296
rect 1128 2264 1160 2296
rect 1200 2264 1232 2296
rect 1272 2264 1304 2296
rect 1344 2264 1376 2296
rect 1416 2264 1448 2296
rect 1488 2264 1520 2296
rect 1560 2264 1592 2296
rect 1632 2264 1664 2296
rect 1704 2264 1736 2296
rect 1776 2264 1808 2296
rect 1848 2264 1880 2296
rect 1920 2264 1952 2296
rect 48 2192 80 2224
rect 120 2192 152 2224
rect 192 2192 224 2224
rect 264 2192 296 2224
rect 336 2192 368 2224
rect 408 2192 440 2224
rect 480 2192 512 2224
rect 552 2192 584 2224
rect 624 2192 656 2224
rect 696 2192 728 2224
rect 768 2192 800 2224
rect 840 2192 872 2224
rect 912 2192 944 2224
rect 984 2192 1016 2224
rect 1056 2192 1088 2224
rect 1128 2192 1160 2224
rect 1200 2192 1232 2224
rect 1272 2192 1304 2224
rect 1344 2192 1376 2224
rect 1416 2192 1448 2224
rect 1488 2192 1520 2224
rect 1560 2192 1592 2224
rect 1632 2192 1664 2224
rect 1704 2192 1736 2224
rect 1776 2192 1808 2224
rect 1848 2192 1880 2224
rect 1920 2192 1952 2224
rect 48 2120 80 2152
rect 120 2120 152 2152
rect 192 2120 224 2152
rect 264 2120 296 2152
rect 336 2120 368 2152
rect 408 2120 440 2152
rect 480 2120 512 2152
rect 552 2120 584 2152
rect 624 2120 656 2152
rect 696 2120 728 2152
rect 768 2120 800 2152
rect 840 2120 872 2152
rect 912 2120 944 2152
rect 984 2120 1016 2152
rect 1056 2120 1088 2152
rect 1128 2120 1160 2152
rect 1200 2120 1232 2152
rect 1272 2120 1304 2152
rect 1344 2120 1376 2152
rect 1416 2120 1448 2152
rect 1488 2120 1520 2152
rect 1560 2120 1592 2152
rect 1632 2120 1664 2152
rect 1704 2120 1736 2152
rect 1776 2120 1808 2152
rect 1848 2120 1880 2152
rect 1920 2120 1952 2152
rect 48 2048 80 2080
rect 120 2048 152 2080
rect 192 2048 224 2080
rect 264 2048 296 2080
rect 336 2048 368 2080
rect 408 2048 440 2080
rect 480 2048 512 2080
rect 552 2048 584 2080
rect 624 2048 656 2080
rect 696 2048 728 2080
rect 768 2048 800 2080
rect 840 2048 872 2080
rect 912 2048 944 2080
rect 984 2048 1016 2080
rect 1056 2048 1088 2080
rect 1128 2048 1160 2080
rect 1200 2048 1232 2080
rect 1272 2048 1304 2080
rect 1344 2048 1376 2080
rect 1416 2048 1448 2080
rect 1488 2048 1520 2080
rect 1560 2048 1592 2080
rect 1632 2048 1664 2080
rect 1704 2048 1736 2080
rect 1776 2048 1808 2080
rect 1848 2048 1880 2080
rect 1920 2048 1952 2080
rect 48 1976 80 2008
rect 120 1976 152 2008
rect 192 1976 224 2008
rect 264 1976 296 2008
rect 336 1976 368 2008
rect 408 1976 440 2008
rect 480 1976 512 2008
rect 552 1976 584 2008
rect 624 1976 656 2008
rect 696 1976 728 2008
rect 768 1976 800 2008
rect 840 1976 872 2008
rect 912 1976 944 2008
rect 984 1976 1016 2008
rect 1056 1976 1088 2008
rect 1128 1976 1160 2008
rect 1200 1976 1232 2008
rect 1272 1976 1304 2008
rect 1344 1976 1376 2008
rect 1416 1976 1448 2008
rect 1488 1976 1520 2008
rect 1560 1976 1592 2008
rect 1632 1976 1664 2008
rect 1704 1976 1736 2008
rect 1776 1976 1808 2008
rect 1848 1976 1880 2008
rect 1920 1976 1952 2008
rect 48 1904 80 1936
rect 120 1904 152 1936
rect 192 1904 224 1936
rect 264 1904 296 1936
rect 336 1904 368 1936
rect 408 1904 440 1936
rect 480 1904 512 1936
rect 552 1904 584 1936
rect 624 1904 656 1936
rect 696 1904 728 1936
rect 768 1904 800 1936
rect 840 1904 872 1936
rect 912 1904 944 1936
rect 984 1904 1016 1936
rect 1056 1904 1088 1936
rect 1128 1904 1160 1936
rect 1200 1904 1232 1936
rect 1272 1904 1304 1936
rect 1344 1904 1376 1936
rect 1416 1904 1448 1936
rect 1488 1904 1520 1936
rect 1560 1904 1592 1936
rect 1632 1904 1664 1936
rect 1704 1904 1736 1936
rect 1776 1904 1808 1936
rect 1848 1904 1880 1936
rect 1920 1904 1952 1936
rect 48 1832 80 1864
rect 120 1832 152 1864
rect 192 1832 224 1864
rect 264 1832 296 1864
rect 336 1832 368 1864
rect 408 1832 440 1864
rect 480 1832 512 1864
rect 552 1832 584 1864
rect 624 1832 656 1864
rect 696 1832 728 1864
rect 768 1832 800 1864
rect 840 1832 872 1864
rect 912 1832 944 1864
rect 984 1832 1016 1864
rect 1056 1832 1088 1864
rect 1128 1832 1160 1864
rect 1200 1832 1232 1864
rect 1272 1832 1304 1864
rect 1344 1832 1376 1864
rect 1416 1832 1448 1864
rect 1488 1832 1520 1864
rect 1560 1832 1592 1864
rect 1632 1832 1664 1864
rect 1704 1832 1736 1864
rect 1776 1832 1808 1864
rect 1848 1832 1880 1864
rect 1920 1832 1952 1864
rect 48 1760 80 1792
rect 120 1760 152 1792
rect 192 1760 224 1792
rect 264 1760 296 1792
rect 336 1760 368 1792
rect 408 1760 440 1792
rect 480 1760 512 1792
rect 552 1760 584 1792
rect 624 1760 656 1792
rect 696 1760 728 1792
rect 768 1760 800 1792
rect 840 1760 872 1792
rect 912 1760 944 1792
rect 984 1760 1016 1792
rect 1056 1760 1088 1792
rect 1128 1760 1160 1792
rect 1200 1760 1232 1792
rect 1272 1760 1304 1792
rect 1344 1760 1376 1792
rect 1416 1760 1448 1792
rect 1488 1760 1520 1792
rect 1560 1760 1592 1792
rect 1632 1760 1664 1792
rect 1704 1760 1736 1792
rect 1776 1760 1808 1792
rect 1848 1760 1880 1792
rect 1920 1760 1952 1792
rect 48 1688 80 1720
rect 120 1688 152 1720
rect 192 1688 224 1720
rect 264 1688 296 1720
rect 336 1688 368 1720
rect 408 1688 440 1720
rect 480 1688 512 1720
rect 552 1688 584 1720
rect 624 1688 656 1720
rect 696 1688 728 1720
rect 768 1688 800 1720
rect 840 1688 872 1720
rect 912 1688 944 1720
rect 984 1688 1016 1720
rect 1056 1688 1088 1720
rect 1128 1688 1160 1720
rect 1200 1688 1232 1720
rect 1272 1688 1304 1720
rect 1344 1688 1376 1720
rect 1416 1688 1448 1720
rect 1488 1688 1520 1720
rect 1560 1688 1592 1720
rect 1632 1688 1664 1720
rect 1704 1688 1736 1720
rect 1776 1688 1808 1720
rect 1848 1688 1880 1720
rect 1920 1688 1952 1720
rect 48 1616 80 1648
rect 120 1616 152 1648
rect 192 1616 224 1648
rect 264 1616 296 1648
rect 336 1616 368 1648
rect 408 1616 440 1648
rect 480 1616 512 1648
rect 552 1616 584 1648
rect 624 1616 656 1648
rect 696 1616 728 1648
rect 768 1616 800 1648
rect 840 1616 872 1648
rect 912 1616 944 1648
rect 984 1616 1016 1648
rect 1056 1616 1088 1648
rect 1128 1616 1160 1648
rect 1200 1616 1232 1648
rect 1272 1616 1304 1648
rect 1344 1616 1376 1648
rect 1416 1616 1448 1648
rect 1488 1616 1520 1648
rect 1560 1616 1592 1648
rect 1632 1616 1664 1648
rect 1704 1616 1736 1648
rect 1776 1616 1808 1648
rect 1848 1616 1880 1648
rect 1920 1616 1952 1648
rect 48 1544 80 1576
rect 120 1544 152 1576
rect 192 1544 224 1576
rect 264 1544 296 1576
rect 336 1544 368 1576
rect 408 1544 440 1576
rect 480 1544 512 1576
rect 552 1544 584 1576
rect 624 1544 656 1576
rect 696 1544 728 1576
rect 768 1544 800 1576
rect 840 1544 872 1576
rect 912 1544 944 1576
rect 984 1544 1016 1576
rect 1056 1544 1088 1576
rect 1128 1544 1160 1576
rect 1200 1544 1232 1576
rect 1272 1544 1304 1576
rect 1344 1544 1376 1576
rect 1416 1544 1448 1576
rect 1488 1544 1520 1576
rect 1560 1544 1592 1576
rect 1632 1544 1664 1576
rect 1704 1544 1736 1576
rect 1776 1544 1808 1576
rect 1848 1544 1880 1576
rect 1920 1544 1952 1576
rect 48 1472 80 1504
rect 120 1472 152 1504
rect 192 1472 224 1504
rect 264 1472 296 1504
rect 336 1472 368 1504
rect 408 1472 440 1504
rect 480 1472 512 1504
rect 552 1472 584 1504
rect 624 1472 656 1504
rect 696 1472 728 1504
rect 768 1472 800 1504
rect 840 1472 872 1504
rect 912 1472 944 1504
rect 984 1472 1016 1504
rect 1056 1472 1088 1504
rect 1128 1472 1160 1504
rect 1200 1472 1232 1504
rect 1272 1472 1304 1504
rect 1344 1472 1376 1504
rect 1416 1472 1448 1504
rect 1488 1472 1520 1504
rect 1560 1472 1592 1504
rect 1632 1472 1664 1504
rect 1704 1472 1736 1504
rect 1776 1472 1808 1504
rect 1848 1472 1880 1504
rect 1920 1472 1952 1504
rect 48 1400 80 1432
rect 120 1400 152 1432
rect 192 1400 224 1432
rect 264 1400 296 1432
rect 336 1400 368 1432
rect 408 1400 440 1432
rect 480 1400 512 1432
rect 552 1400 584 1432
rect 624 1400 656 1432
rect 696 1400 728 1432
rect 768 1400 800 1432
rect 840 1400 872 1432
rect 912 1400 944 1432
rect 984 1400 1016 1432
rect 1056 1400 1088 1432
rect 1128 1400 1160 1432
rect 1200 1400 1232 1432
rect 1272 1400 1304 1432
rect 1344 1400 1376 1432
rect 1416 1400 1448 1432
rect 1488 1400 1520 1432
rect 1560 1400 1592 1432
rect 1632 1400 1664 1432
rect 1704 1400 1736 1432
rect 1776 1400 1808 1432
rect 1848 1400 1880 1432
rect 1920 1400 1952 1432
rect 48 1328 80 1360
rect 120 1328 152 1360
rect 192 1328 224 1360
rect 264 1328 296 1360
rect 336 1328 368 1360
rect 408 1328 440 1360
rect 480 1328 512 1360
rect 552 1328 584 1360
rect 624 1328 656 1360
rect 696 1328 728 1360
rect 768 1328 800 1360
rect 840 1328 872 1360
rect 912 1328 944 1360
rect 984 1328 1016 1360
rect 1056 1328 1088 1360
rect 1128 1328 1160 1360
rect 1200 1328 1232 1360
rect 1272 1328 1304 1360
rect 1344 1328 1376 1360
rect 1416 1328 1448 1360
rect 1488 1328 1520 1360
rect 1560 1328 1592 1360
rect 1632 1328 1664 1360
rect 1704 1328 1736 1360
rect 1776 1328 1808 1360
rect 1848 1328 1880 1360
rect 1920 1328 1952 1360
rect 48 1256 80 1288
rect 120 1256 152 1288
rect 192 1256 224 1288
rect 264 1256 296 1288
rect 336 1256 368 1288
rect 408 1256 440 1288
rect 480 1256 512 1288
rect 552 1256 584 1288
rect 624 1256 656 1288
rect 696 1256 728 1288
rect 768 1256 800 1288
rect 840 1256 872 1288
rect 912 1256 944 1288
rect 984 1256 1016 1288
rect 1056 1256 1088 1288
rect 1128 1256 1160 1288
rect 1200 1256 1232 1288
rect 1272 1256 1304 1288
rect 1344 1256 1376 1288
rect 1416 1256 1448 1288
rect 1488 1256 1520 1288
rect 1560 1256 1592 1288
rect 1632 1256 1664 1288
rect 1704 1256 1736 1288
rect 1776 1256 1808 1288
rect 1848 1256 1880 1288
rect 1920 1256 1952 1288
rect 768 31384 800 31416
rect 838 31384 870 31416
rect 907 31384 939 31416
rect 978 31384 1010 31416
rect 1048 31384 1080 31416
rect 1116 31384 1148 31416
rect 1186 31384 1218 31416
rect 192 27939 224 27971
rect 264 27939 296 27971
rect 336 27939 368 27971
rect 408 27939 440 27971
rect 480 27939 512 27971
rect 552 27939 584 27971
rect 624 27939 656 27971
rect 696 27939 728 27971
rect 768 27939 800 27971
rect 840 27939 872 27971
rect 912 27939 944 27971
rect 984 27939 1016 27971
rect 1056 27939 1088 27971
rect 1128 27939 1160 27971
rect 1200 27939 1232 27971
rect 1272 27939 1304 27971
rect 1344 27939 1376 27971
rect 1416 27939 1448 27971
rect 1488 27939 1520 27971
rect 1560 27939 1592 27971
rect 1632 27939 1664 27971
rect 1704 27939 1736 27971
rect 1776 27939 1808 27971
rect 1848 27939 1880 27971
rect 120 27867 152 27899
rect 192 27867 224 27899
rect 264 27867 296 27899
rect 336 27867 368 27899
rect 408 27867 440 27899
rect 480 27867 512 27899
rect 552 27867 584 27899
rect 624 27867 656 27899
rect 696 27867 728 27899
rect 768 27867 800 27899
rect 840 27867 872 27899
rect 912 27867 944 27899
rect 984 27867 1016 27899
rect 1056 27867 1088 27899
rect 1128 27867 1160 27899
rect 1200 27867 1232 27899
rect 1272 27867 1304 27899
rect 1344 27867 1376 27899
rect 1416 27867 1448 27899
rect 1488 27867 1520 27899
rect 1560 27867 1592 27899
rect 1632 27867 1664 27899
rect 1704 27867 1736 27899
rect 1776 27867 1808 27899
rect 1848 27867 1880 27899
rect 120 27795 152 27827
rect 192 27795 224 27827
rect 264 27795 296 27827
rect 336 27795 368 27827
rect 408 27795 440 27827
rect 480 27795 512 27827
rect 552 27795 584 27827
rect 624 27795 656 27827
rect 696 27795 728 27827
rect 768 27795 800 27827
rect 840 27795 872 27827
rect 912 27795 944 27827
rect 984 27795 1016 27827
rect 1056 27795 1088 27827
rect 1128 27795 1160 27827
rect 1200 27795 1232 27827
rect 1272 27795 1304 27827
rect 1344 27795 1376 27827
rect 1416 27795 1448 27827
rect 1488 27795 1520 27827
rect 1560 27795 1592 27827
rect 1632 27795 1664 27827
rect 1704 27795 1736 27827
rect 1776 27795 1808 27827
rect 1848 27795 1880 27827
rect 120 27723 152 27755
rect 192 27723 224 27755
rect 264 27723 296 27755
rect 336 27723 368 27755
rect 408 27723 440 27755
rect 480 27723 512 27755
rect 552 27723 584 27755
rect 624 27723 656 27755
rect 696 27723 728 27755
rect 768 27723 800 27755
rect 840 27723 872 27755
rect 912 27723 944 27755
rect 984 27723 1016 27755
rect 1056 27723 1088 27755
rect 1128 27723 1160 27755
rect 1200 27723 1232 27755
rect 1272 27723 1304 27755
rect 1344 27723 1376 27755
rect 1416 27723 1448 27755
rect 1488 27723 1520 27755
rect 1560 27723 1592 27755
rect 1632 27723 1664 27755
rect 1704 27723 1736 27755
rect 1776 27723 1808 27755
rect 1848 27723 1880 27755
rect 120 27651 152 27683
rect 192 27651 224 27683
rect 264 27651 296 27683
rect 336 27651 368 27683
rect 408 27651 440 27683
rect 480 27651 512 27683
rect 552 27651 584 27683
rect 624 27651 656 27683
rect 696 27651 728 27683
rect 768 27651 800 27683
rect 840 27651 872 27683
rect 912 27651 944 27683
rect 984 27651 1016 27683
rect 1056 27651 1088 27683
rect 1128 27651 1160 27683
rect 1200 27651 1232 27683
rect 1272 27651 1304 27683
rect 1344 27651 1376 27683
rect 1416 27651 1448 27683
rect 1488 27651 1520 27683
rect 1560 27651 1592 27683
rect 1632 27651 1664 27683
rect 1704 27651 1736 27683
rect 1776 27651 1808 27683
rect 1848 27651 1880 27683
rect 120 27579 152 27611
rect 192 27579 224 27611
rect 264 27579 296 27611
rect 336 27579 368 27611
rect 408 27579 440 27611
rect 480 27579 512 27611
rect 552 27579 584 27611
rect 624 27579 656 27611
rect 696 27579 728 27611
rect 768 27579 800 27611
rect 840 27579 872 27611
rect 912 27579 944 27611
rect 984 27579 1016 27611
rect 1056 27579 1088 27611
rect 1128 27579 1160 27611
rect 1200 27579 1232 27611
rect 1272 27579 1304 27611
rect 1344 27579 1376 27611
rect 1416 27579 1448 27611
rect 1488 27579 1520 27611
rect 1560 27579 1592 27611
rect 1632 27579 1664 27611
rect 1704 27579 1736 27611
rect 1776 27579 1808 27611
rect 1848 27579 1880 27611
rect 120 27507 152 27539
rect 192 27507 224 27539
rect 264 27507 296 27539
rect 336 27507 368 27539
rect 408 27507 440 27539
rect 480 27507 512 27539
rect 552 27507 584 27539
rect 624 27507 656 27539
rect 696 27507 728 27539
rect 768 27507 800 27539
rect 840 27507 872 27539
rect 912 27507 944 27539
rect 984 27507 1016 27539
rect 1056 27507 1088 27539
rect 1128 27507 1160 27539
rect 1200 27507 1232 27539
rect 1272 27507 1304 27539
rect 1344 27507 1376 27539
rect 1416 27507 1448 27539
rect 1488 27507 1520 27539
rect 1560 27507 1592 27539
rect 1632 27507 1664 27539
rect 1704 27507 1736 27539
rect 1776 27507 1808 27539
rect 1848 27507 1880 27539
rect 120 27435 152 27467
rect 192 27435 224 27467
rect 264 27435 296 27467
rect 336 27435 368 27467
rect 408 27435 440 27467
rect 480 27435 512 27467
rect 552 27435 584 27467
rect 624 27435 656 27467
rect 696 27435 728 27467
rect 768 27435 800 27467
rect 840 27435 872 27467
rect 912 27435 944 27467
rect 984 27435 1016 27467
rect 1056 27435 1088 27467
rect 1128 27435 1160 27467
rect 1200 27435 1232 27467
rect 1272 27435 1304 27467
rect 1344 27435 1376 27467
rect 1416 27435 1448 27467
rect 1488 27435 1520 27467
rect 1560 27435 1592 27467
rect 1632 27435 1664 27467
rect 1704 27435 1736 27467
rect 1776 27435 1808 27467
rect 1848 27435 1880 27467
rect 120 27363 152 27395
rect 192 27363 224 27395
rect 264 27363 296 27395
rect 336 27363 368 27395
rect 408 27363 440 27395
rect 480 27363 512 27395
rect 552 27363 584 27395
rect 624 27363 656 27395
rect 696 27363 728 27395
rect 768 27363 800 27395
rect 840 27363 872 27395
rect 912 27363 944 27395
rect 984 27363 1016 27395
rect 1056 27363 1088 27395
rect 1128 27363 1160 27395
rect 1200 27363 1232 27395
rect 1272 27363 1304 27395
rect 1344 27363 1376 27395
rect 1416 27363 1448 27395
rect 1488 27363 1520 27395
rect 1560 27363 1592 27395
rect 1632 27363 1664 27395
rect 1704 27363 1736 27395
rect 1776 27363 1808 27395
rect 1848 27363 1880 27395
rect 120 27291 152 27323
rect 192 27291 224 27323
rect 264 27291 296 27323
rect 336 27291 368 27323
rect 408 27291 440 27323
rect 480 27291 512 27323
rect 552 27291 584 27323
rect 624 27291 656 27323
rect 696 27291 728 27323
rect 768 27291 800 27323
rect 840 27291 872 27323
rect 912 27291 944 27323
rect 984 27291 1016 27323
rect 1056 27291 1088 27323
rect 1128 27291 1160 27323
rect 1200 27291 1232 27323
rect 1272 27291 1304 27323
rect 1344 27291 1376 27323
rect 1416 27291 1448 27323
rect 1488 27291 1520 27323
rect 1560 27291 1592 27323
rect 1632 27291 1664 27323
rect 1704 27291 1736 27323
rect 1776 27291 1808 27323
rect 1848 27291 1880 27323
rect 120 27219 152 27251
rect 192 27219 224 27251
rect 264 27219 296 27251
rect 336 27219 368 27251
rect 408 27219 440 27251
rect 480 27219 512 27251
rect 552 27219 584 27251
rect 624 27219 656 27251
rect 696 27219 728 27251
rect 768 27219 800 27251
rect 840 27219 872 27251
rect 912 27219 944 27251
rect 984 27219 1016 27251
rect 1056 27219 1088 27251
rect 1128 27219 1160 27251
rect 1200 27219 1232 27251
rect 1272 27219 1304 27251
rect 1344 27219 1376 27251
rect 1416 27219 1448 27251
rect 1488 27219 1520 27251
rect 1560 27219 1592 27251
rect 1632 27219 1664 27251
rect 1704 27219 1736 27251
rect 1776 27219 1808 27251
rect 1848 27219 1880 27251
rect 120 27147 152 27179
rect 192 27147 224 27179
rect 264 27147 296 27179
rect 336 27147 368 27179
rect 408 27147 440 27179
rect 480 27147 512 27179
rect 552 27147 584 27179
rect 624 27147 656 27179
rect 696 27147 728 27179
rect 768 27147 800 27179
rect 840 27147 872 27179
rect 912 27147 944 27179
rect 984 27147 1016 27179
rect 1056 27147 1088 27179
rect 1128 27147 1160 27179
rect 1200 27147 1232 27179
rect 1272 27147 1304 27179
rect 1344 27147 1376 27179
rect 1416 27147 1448 27179
rect 1488 27147 1520 27179
rect 1560 27147 1592 27179
rect 1632 27147 1664 27179
rect 1704 27147 1736 27179
rect 1776 27147 1808 27179
rect 1848 27147 1880 27179
rect 120 27075 152 27107
rect 192 27075 224 27107
rect 264 27075 296 27107
rect 336 27075 368 27107
rect 408 27075 440 27107
rect 480 27075 512 27107
rect 552 27075 584 27107
rect 624 27075 656 27107
rect 696 27075 728 27107
rect 768 27075 800 27107
rect 840 27075 872 27107
rect 912 27075 944 27107
rect 984 27075 1016 27107
rect 1056 27075 1088 27107
rect 1128 27075 1160 27107
rect 1200 27075 1232 27107
rect 1272 27075 1304 27107
rect 1344 27075 1376 27107
rect 1416 27075 1448 27107
rect 1488 27075 1520 27107
rect 1560 27075 1592 27107
rect 1632 27075 1664 27107
rect 1704 27075 1736 27107
rect 1776 27075 1808 27107
rect 1848 27075 1880 27107
rect 120 27003 152 27035
rect 192 27003 224 27035
rect 264 27003 296 27035
rect 336 27003 368 27035
rect 408 27003 440 27035
rect 480 27003 512 27035
rect 552 27003 584 27035
rect 624 27003 656 27035
rect 696 27003 728 27035
rect 768 27003 800 27035
rect 840 27003 872 27035
rect 912 27003 944 27035
rect 984 27003 1016 27035
rect 1056 27003 1088 27035
rect 1128 27003 1160 27035
rect 1200 27003 1232 27035
rect 1272 27003 1304 27035
rect 1344 27003 1376 27035
rect 1416 27003 1448 27035
rect 1488 27003 1520 27035
rect 1560 27003 1592 27035
rect 1632 27003 1664 27035
rect 1704 27003 1736 27035
rect 1776 27003 1808 27035
rect 1848 27003 1880 27035
rect 120 26931 152 26963
rect 192 26931 224 26963
rect 264 26931 296 26963
rect 336 26931 368 26963
rect 408 26931 440 26963
rect 480 26931 512 26963
rect 552 26931 584 26963
rect 624 26931 656 26963
rect 696 26931 728 26963
rect 768 26931 800 26963
rect 840 26931 872 26963
rect 912 26931 944 26963
rect 984 26931 1016 26963
rect 1056 26931 1088 26963
rect 1128 26931 1160 26963
rect 1200 26931 1232 26963
rect 1272 26931 1304 26963
rect 1344 26931 1376 26963
rect 1416 26931 1448 26963
rect 1488 26931 1520 26963
rect 1560 26931 1592 26963
rect 1632 26931 1664 26963
rect 1704 26931 1736 26963
rect 1776 26931 1808 26963
rect 1848 26931 1880 26963
rect 120 26859 152 26891
rect 192 26859 224 26891
rect 264 26859 296 26891
rect 336 26859 368 26891
rect 408 26859 440 26891
rect 480 26859 512 26891
rect 552 26859 584 26891
rect 624 26859 656 26891
rect 696 26859 728 26891
rect 768 26859 800 26891
rect 840 26859 872 26891
rect 912 26859 944 26891
rect 984 26859 1016 26891
rect 1056 26859 1088 26891
rect 1128 26859 1160 26891
rect 1200 26859 1232 26891
rect 1272 26859 1304 26891
rect 1344 26859 1376 26891
rect 1416 26859 1448 26891
rect 1488 26859 1520 26891
rect 1560 26859 1592 26891
rect 1632 26859 1664 26891
rect 1704 26859 1736 26891
rect 1776 26859 1808 26891
rect 1848 26859 1880 26891
rect 120 26787 152 26819
rect 192 26787 224 26819
rect 264 26787 296 26819
rect 336 26787 368 26819
rect 408 26787 440 26819
rect 480 26787 512 26819
rect 552 26787 584 26819
rect 624 26787 656 26819
rect 696 26787 728 26819
rect 768 26787 800 26819
rect 840 26787 872 26819
rect 912 26787 944 26819
rect 984 26787 1016 26819
rect 1056 26787 1088 26819
rect 1128 26787 1160 26819
rect 1200 26787 1232 26819
rect 1272 26787 1304 26819
rect 1344 26787 1376 26819
rect 1416 26787 1448 26819
rect 1488 26787 1520 26819
rect 1560 26787 1592 26819
rect 1632 26787 1664 26819
rect 1704 26787 1736 26819
rect 1776 26787 1808 26819
rect 1848 26787 1880 26819
rect 120 26715 152 26747
rect 192 26715 224 26747
rect 264 26715 296 26747
rect 336 26715 368 26747
rect 408 26715 440 26747
rect 480 26715 512 26747
rect 552 26715 584 26747
rect 624 26715 656 26747
rect 696 26715 728 26747
rect 768 26715 800 26747
rect 840 26715 872 26747
rect 912 26715 944 26747
rect 984 26715 1016 26747
rect 1056 26715 1088 26747
rect 1128 26715 1160 26747
rect 1200 26715 1232 26747
rect 1272 26715 1304 26747
rect 1344 26715 1376 26747
rect 1416 26715 1448 26747
rect 1488 26715 1520 26747
rect 1560 26715 1592 26747
rect 1632 26715 1664 26747
rect 1704 26715 1736 26747
rect 1776 26715 1808 26747
rect 1848 26715 1880 26747
rect 120 26643 152 26675
rect 192 26643 224 26675
rect 264 26643 296 26675
rect 336 26643 368 26675
rect 408 26643 440 26675
rect 480 26643 512 26675
rect 552 26643 584 26675
rect 624 26643 656 26675
rect 696 26643 728 26675
rect 768 26643 800 26675
rect 840 26643 872 26675
rect 912 26643 944 26675
rect 984 26643 1016 26675
rect 1056 26643 1088 26675
rect 1128 26643 1160 26675
rect 1200 26643 1232 26675
rect 1272 26643 1304 26675
rect 1344 26643 1376 26675
rect 1416 26643 1448 26675
rect 1488 26643 1520 26675
rect 1560 26643 1592 26675
rect 1632 26643 1664 26675
rect 1704 26643 1736 26675
rect 1776 26643 1808 26675
rect 1848 26643 1880 26675
rect 120 26571 152 26603
rect 192 26571 224 26603
rect 264 26571 296 26603
rect 336 26571 368 26603
rect 408 26571 440 26603
rect 480 26571 512 26603
rect 552 26571 584 26603
rect 624 26571 656 26603
rect 696 26571 728 26603
rect 768 26571 800 26603
rect 840 26571 872 26603
rect 912 26571 944 26603
rect 984 26571 1016 26603
rect 1056 26571 1088 26603
rect 1128 26571 1160 26603
rect 1200 26571 1232 26603
rect 1272 26571 1304 26603
rect 1344 26571 1376 26603
rect 1416 26571 1448 26603
rect 1488 26571 1520 26603
rect 1560 26571 1592 26603
rect 1632 26571 1664 26603
rect 1704 26571 1736 26603
rect 1776 26571 1808 26603
rect 1848 26571 1880 26603
rect 120 26499 152 26531
rect 192 26499 224 26531
rect 264 26499 296 26531
rect 336 26499 368 26531
rect 408 26499 440 26531
rect 480 26499 512 26531
rect 552 26499 584 26531
rect 624 26499 656 26531
rect 696 26499 728 26531
rect 768 26499 800 26531
rect 840 26499 872 26531
rect 912 26499 944 26531
rect 984 26499 1016 26531
rect 1056 26499 1088 26531
rect 1128 26499 1160 26531
rect 1200 26499 1232 26531
rect 1272 26499 1304 26531
rect 1344 26499 1376 26531
rect 1416 26499 1448 26531
rect 1488 26499 1520 26531
rect 1560 26499 1592 26531
rect 1632 26499 1664 26531
rect 1704 26499 1736 26531
rect 1776 26499 1808 26531
rect 1848 26499 1880 26531
rect 120 26427 152 26459
rect 192 26427 224 26459
rect 264 26427 296 26459
rect 336 26427 368 26459
rect 408 26427 440 26459
rect 480 26427 512 26459
rect 552 26427 584 26459
rect 624 26427 656 26459
rect 696 26427 728 26459
rect 768 26427 800 26459
rect 840 26427 872 26459
rect 912 26427 944 26459
rect 984 26427 1016 26459
rect 1056 26427 1088 26459
rect 1128 26427 1160 26459
rect 1200 26427 1232 26459
rect 1272 26427 1304 26459
rect 1344 26427 1376 26459
rect 1416 26427 1448 26459
rect 1488 26427 1520 26459
rect 1560 26427 1592 26459
rect 1632 26427 1664 26459
rect 1704 26427 1736 26459
rect 1776 26427 1808 26459
rect 1848 26427 1880 26459
rect 120 26355 152 26387
rect 192 26355 224 26387
rect 264 26355 296 26387
rect 336 26355 368 26387
rect 408 26355 440 26387
rect 480 26355 512 26387
rect 552 26355 584 26387
rect 624 26355 656 26387
rect 696 26355 728 26387
rect 768 26355 800 26387
rect 840 26355 872 26387
rect 912 26355 944 26387
rect 984 26355 1016 26387
rect 1056 26355 1088 26387
rect 1128 26355 1160 26387
rect 1200 26355 1232 26387
rect 1272 26355 1304 26387
rect 1344 26355 1376 26387
rect 1416 26355 1448 26387
rect 1488 26355 1520 26387
rect 1560 26355 1592 26387
rect 1632 26355 1664 26387
rect 1704 26355 1736 26387
rect 1776 26355 1808 26387
rect 1848 26355 1880 26387
rect 120 26283 152 26315
rect 192 26283 224 26315
rect 264 26283 296 26315
rect 336 26283 368 26315
rect 408 26283 440 26315
rect 480 26283 512 26315
rect 552 26283 584 26315
rect 624 26283 656 26315
rect 696 26283 728 26315
rect 768 26283 800 26315
rect 840 26283 872 26315
rect 912 26283 944 26315
rect 984 26283 1016 26315
rect 1056 26283 1088 26315
rect 1128 26283 1160 26315
rect 1200 26283 1232 26315
rect 1272 26283 1304 26315
rect 1344 26283 1376 26315
rect 1416 26283 1448 26315
rect 1488 26283 1520 26315
rect 1560 26283 1592 26315
rect 1632 26283 1664 26315
rect 1704 26283 1736 26315
rect 1776 26283 1808 26315
rect 1848 26283 1880 26315
rect 120 26211 152 26243
rect 192 26211 224 26243
rect 264 26211 296 26243
rect 336 26211 368 26243
rect 408 26211 440 26243
rect 480 26211 512 26243
rect 552 26211 584 26243
rect 624 26211 656 26243
rect 696 26211 728 26243
rect 768 26211 800 26243
rect 840 26211 872 26243
rect 912 26211 944 26243
rect 984 26211 1016 26243
rect 1056 26211 1088 26243
rect 1128 26211 1160 26243
rect 1200 26211 1232 26243
rect 1272 26211 1304 26243
rect 1344 26211 1376 26243
rect 1416 26211 1448 26243
rect 1488 26211 1520 26243
rect 1560 26211 1592 26243
rect 1632 26211 1664 26243
rect 1704 26211 1736 26243
rect 1776 26211 1808 26243
rect 1848 26211 1880 26243
rect 120 26139 152 26171
rect 192 26139 224 26171
rect 264 26139 296 26171
rect 336 26139 368 26171
rect 408 26139 440 26171
rect 480 26139 512 26171
rect 552 26139 584 26171
rect 624 26139 656 26171
rect 696 26139 728 26171
rect 768 26139 800 26171
rect 840 26139 872 26171
rect 912 26139 944 26171
rect 984 26139 1016 26171
rect 1056 26139 1088 26171
rect 1128 26139 1160 26171
rect 1200 26139 1232 26171
rect 1272 26139 1304 26171
rect 1344 26139 1376 26171
rect 1416 26139 1448 26171
rect 1488 26139 1520 26171
rect 1560 26139 1592 26171
rect 1632 26139 1664 26171
rect 1704 26139 1736 26171
rect 1776 26139 1808 26171
rect 1848 26139 1880 26171
rect 120 26067 152 26099
rect 192 26067 224 26099
rect 264 26067 296 26099
rect 336 26067 368 26099
rect 408 26067 440 26099
rect 480 26067 512 26099
rect 552 26067 584 26099
rect 624 26067 656 26099
rect 696 26067 728 26099
rect 768 26067 800 26099
rect 840 26067 872 26099
rect 912 26067 944 26099
rect 984 26067 1016 26099
rect 1056 26067 1088 26099
rect 1128 26067 1160 26099
rect 1200 26067 1232 26099
rect 1272 26067 1304 26099
rect 1344 26067 1376 26099
rect 1416 26067 1448 26099
rect 1488 26067 1520 26099
rect 1560 26067 1592 26099
rect 1632 26067 1664 26099
rect 1704 26067 1736 26099
rect 1776 26067 1808 26099
rect 1848 26067 1880 26099
rect 120 25995 152 26027
rect 192 25995 224 26027
rect 264 25995 296 26027
rect 336 25995 368 26027
rect 408 25995 440 26027
rect 480 25995 512 26027
rect 552 25995 584 26027
rect 624 25995 656 26027
rect 696 25995 728 26027
rect 768 25995 800 26027
rect 840 25995 872 26027
rect 912 25995 944 26027
rect 984 25995 1016 26027
rect 1056 25995 1088 26027
rect 1128 25995 1160 26027
rect 1200 25995 1232 26027
rect 1272 25995 1304 26027
rect 1344 25995 1376 26027
rect 1416 25995 1448 26027
rect 1488 25995 1520 26027
rect 1560 25995 1592 26027
rect 1632 25995 1664 26027
rect 1704 25995 1736 26027
rect 1776 25995 1808 26027
rect 1848 25995 1880 26027
rect 120 25923 152 25955
rect 192 25923 224 25955
rect 264 25923 296 25955
rect 336 25923 368 25955
rect 408 25923 440 25955
rect 480 25923 512 25955
rect 552 25923 584 25955
rect 624 25923 656 25955
rect 696 25923 728 25955
rect 768 25923 800 25955
rect 840 25923 872 25955
rect 912 25923 944 25955
rect 984 25923 1016 25955
rect 1056 25923 1088 25955
rect 1128 25923 1160 25955
rect 1200 25923 1232 25955
rect 1272 25923 1304 25955
rect 1344 25923 1376 25955
rect 1416 25923 1448 25955
rect 1488 25923 1520 25955
rect 1560 25923 1592 25955
rect 1632 25923 1664 25955
rect 1704 25923 1736 25955
rect 1776 25923 1808 25955
rect 1848 25923 1880 25955
rect 120 25851 152 25883
rect 192 25851 224 25883
rect 264 25851 296 25883
rect 336 25851 368 25883
rect 408 25851 440 25883
rect 480 25851 512 25883
rect 552 25851 584 25883
rect 624 25851 656 25883
rect 696 25851 728 25883
rect 768 25851 800 25883
rect 840 25851 872 25883
rect 912 25851 944 25883
rect 984 25851 1016 25883
rect 1056 25851 1088 25883
rect 1128 25851 1160 25883
rect 1200 25851 1232 25883
rect 1272 25851 1304 25883
rect 1344 25851 1376 25883
rect 1416 25851 1448 25883
rect 1488 25851 1520 25883
rect 1560 25851 1592 25883
rect 1632 25851 1664 25883
rect 1704 25851 1736 25883
rect 1776 25851 1808 25883
rect 1848 25851 1880 25883
rect 120 25779 152 25811
rect 192 25779 224 25811
rect 264 25779 296 25811
rect 336 25779 368 25811
rect 408 25779 440 25811
rect 480 25779 512 25811
rect 552 25779 584 25811
rect 624 25779 656 25811
rect 696 25779 728 25811
rect 768 25779 800 25811
rect 840 25779 872 25811
rect 912 25779 944 25811
rect 984 25779 1016 25811
rect 1056 25779 1088 25811
rect 1128 25779 1160 25811
rect 1200 25779 1232 25811
rect 1272 25779 1304 25811
rect 1344 25779 1376 25811
rect 1416 25779 1448 25811
rect 1488 25779 1520 25811
rect 1560 25779 1592 25811
rect 1632 25779 1664 25811
rect 1704 25779 1736 25811
rect 1776 25779 1808 25811
rect 1848 25779 1880 25811
rect 120 25707 152 25739
rect 192 25707 224 25739
rect 264 25707 296 25739
rect 336 25707 368 25739
rect 408 25707 440 25739
rect 480 25707 512 25739
rect 552 25707 584 25739
rect 624 25707 656 25739
rect 696 25707 728 25739
rect 768 25707 800 25739
rect 840 25707 872 25739
rect 912 25707 944 25739
rect 984 25707 1016 25739
rect 1056 25707 1088 25739
rect 1128 25707 1160 25739
rect 1200 25707 1232 25739
rect 1272 25707 1304 25739
rect 1344 25707 1376 25739
rect 1416 25707 1448 25739
rect 1488 25707 1520 25739
rect 1560 25707 1592 25739
rect 1632 25707 1664 25739
rect 1704 25707 1736 25739
rect 1776 25707 1808 25739
rect 1848 25707 1880 25739
rect 120 25635 152 25667
rect 192 25635 224 25667
rect 264 25635 296 25667
rect 336 25635 368 25667
rect 408 25635 440 25667
rect 480 25635 512 25667
rect 552 25635 584 25667
rect 624 25635 656 25667
rect 696 25635 728 25667
rect 768 25635 800 25667
rect 840 25635 872 25667
rect 912 25635 944 25667
rect 984 25635 1016 25667
rect 1056 25635 1088 25667
rect 1128 25635 1160 25667
rect 1200 25635 1232 25667
rect 1272 25635 1304 25667
rect 1344 25635 1376 25667
rect 1416 25635 1448 25667
rect 1488 25635 1520 25667
rect 1560 25635 1592 25667
rect 1632 25635 1664 25667
rect 1704 25635 1736 25667
rect 1776 25635 1808 25667
rect 1848 25635 1880 25667
rect 120 25563 152 25595
rect 192 25563 224 25595
rect 264 25563 296 25595
rect 336 25563 368 25595
rect 408 25563 440 25595
rect 480 25563 512 25595
rect 552 25563 584 25595
rect 624 25563 656 25595
rect 696 25563 728 25595
rect 768 25563 800 25595
rect 840 25563 872 25595
rect 912 25563 944 25595
rect 984 25563 1016 25595
rect 1056 25563 1088 25595
rect 1128 25563 1160 25595
rect 1200 25563 1232 25595
rect 1272 25563 1304 25595
rect 1344 25563 1376 25595
rect 1416 25563 1448 25595
rect 1488 25563 1520 25595
rect 1560 25563 1592 25595
rect 1632 25563 1664 25595
rect 1704 25563 1736 25595
rect 1776 25563 1808 25595
rect 1848 25563 1880 25595
rect 120 25491 152 25523
rect 192 25491 224 25523
rect 264 25491 296 25523
rect 336 25491 368 25523
rect 408 25491 440 25523
rect 480 25491 512 25523
rect 552 25491 584 25523
rect 624 25491 656 25523
rect 696 25491 728 25523
rect 768 25491 800 25523
rect 840 25491 872 25523
rect 912 25491 944 25523
rect 984 25491 1016 25523
rect 1056 25491 1088 25523
rect 1128 25491 1160 25523
rect 1200 25491 1232 25523
rect 1272 25491 1304 25523
rect 1344 25491 1376 25523
rect 1416 25491 1448 25523
rect 1488 25491 1520 25523
rect 1560 25491 1592 25523
rect 1632 25491 1664 25523
rect 1704 25491 1736 25523
rect 1776 25491 1808 25523
rect 1848 25491 1880 25523
rect 120 25419 152 25451
rect 192 25419 224 25451
rect 264 25419 296 25451
rect 336 25419 368 25451
rect 408 25419 440 25451
rect 480 25419 512 25451
rect 552 25419 584 25451
rect 624 25419 656 25451
rect 696 25419 728 25451
rect 768 25419 800 25451
rect 840 25419 872 25451
rect 912 25419 944 25451
rect 984 25419 1016 25451
rect 1056 25419 1088 25451
rect 1128 25419 1160 25451
rect 1200 25419 1232 25451
rect 1272 25419 1304 25451
rect 1344 25419 1376 25451
rect 1416 25419 1448 25451
rect 1488 25419 1520 25451
rect 1560 25419 1592 25451
rect 1632 25419 1664 25451
rect 1704 25419 1736 25451
rect 1776 25419 1808 25451
rect 1848 25419 1880 25451
rect 120 25347 152 25379
rect 192 25347 224 25379
rect 264 25347 296 25379
rect 336 25347 368 25379
rect 408 25347 440 25379
rect 480 25347 512 25379
rect 552 25347 584 25379
rect 624 25347 656 25379
rect 696 25347 728 25379
rect 768 25347 800 25379
rect 840 25347 872 25379
rect 912 25347 944 25379
rect 984 25347 1016 25379
rect 1056 25347 1088 25379
rect 1128 25347 1160 25379
rect 1200 25347 1232 25379
rect 1272 25347 1304 25379
rect 1344 25347 1376 25379
rect 1416 25347 1448 25379
rect 1488 25347 1520 25379
rect 1560 25347 1592 25379
rect 1632 25347 1664 25379
rect 1704 25347 1736 25379
rect 1776 25347 1808 25379
rect 1848 25347 1880 25379
rect 120 25275 152 25307
rect 192 25275 224 25307
rect 264 25275 296 25307
rect 336 25275 368 25307
rect 408 25275 440 25307
rect 480 25275 512 25307
rect 552 25275 584 25307
rect 624 25275 656 25307
rect 696 25275 728 25307
rect 768 25275 800 25307
rect 840 25275 872 25307
rect 912 25275 944 25307
rect 984 25275 1016 25307
rect 1056 25275 1088 25307
rect 1128 25275 1160 25307
rect 1200 25275 1232 25307
rect 1272 25275 1304 25307
rect 1344 25275 1376 25307
rect 1416 25275 1448 25307
rect 1488 25275 1520 25307
rect 1560 25275 1592 25307
rect 1632 25275 1664 25307
rect 1704 25275 1736 25307
rect 1776 25275 1808 25307
rect 1848 25275 1880 25307
rect 120 25203 152 25235
rect 192 25203 224 25235
rect 264 25203 296 25235
rect 336 25203 368 25235
rect 408 25203 440 25235
rect 480 25203 512 25235
rect 552 25203 584 25235
rect 624 25203 656 25235
rect 696 25203 728 25235
rect 768 25203 800 25235
rect 840 25203 872 25235
rect 912 25203 944 25235
rect 984 25203 1016 25235
rect 1056 25203 1088 25235
rect 1128 25203 1160 25235
rect 1200 25203 1232 25235
rect 1272 25203 1304 25235
rect 1344 25203 1376 25235
rect 1416 25203 1448 25235
rect 1488 25203 1520 25235
rect 1560 25203 1592 25235
rect 1632 25203 1664 25235
rect 1704 25203 1736 25235
rect 1776 25203 1808 25235
rect 1848 25203 1880 25235
rect 120 25131 152 25163
rect 192 25131 224 25163
rect 264 25131 296 25163
rect 336 25131 368 25163
rect 408 25131 440 25163
rect 480 25131 512 25163
rect 552 25131 584 25163
rect 624 25131 656 25163
rect 696 25131 728 25163
rect 768 25131 800 25163
rect 840 25131 872 25163
rect 912 25131 944 25163
rect 984 25131 1016 25163
rect 1056 25131 1088 25163
rect 1128 25131 1160 25163
rect 1200 25131 1232 25163
rect 1272 25131 1304 25163
rect 1344 25131 1376 25163
rect 1416 25131 1448 25163
rect 1488 25131 1520 25163
rect 1560 25131 1592 25163
rect 1632 25131 1664 25163
rect 1704 25131 1736 25163
rect 1776 25131 1808 25163
rect 1848 25131 1880 25163
rect 120 25059 152 25091
rect 192 25059 224 25091
rect 264 25059 296 25091
rect 336 25059 368 25091
rect 408 25059 440 25091
rect 480 25059 512 25091
rect 552 25059 584 25091
rect 624 25059 656 25091
rect 696 25059 728 25091
rect 768 25059 800 25091
rect 840 25059 872 25091
rect 912 25059 944 25091
rect 984 25059 1016 25091
rect 1056 25059 1088 25091
rect 1128 25059 1160 25091
rect 1200 25059 1232 25091
rect 1272 25059 1304 25091
rect 1344 25059 1376 25091
rect 1416 25059 1448 25091
rect 1488 25059 1520 25091
rect 1560 25059 1592 25091
rect 1632 25059 1664 25091
rect 1704 25059 1736 25091
rect 1776 25059 1808 25091
rect 1848 25059 1880 25091
rect 120 24987 152 25019
rect 192 24987 224 25019
rect 264 24987 296 25019
rect 336 24987 368 25019
rect 408 24987 440 25019
rect 480 24987 512 25019
rect 552 24987 584 25019
rect 624 24987 656 25019
rect 696 24987 728 25019
rect 768 24987 800 25019
rect 840 24987 872 25019
rect 912 24987 944 25019
rect 984 24987 1016 25019
rect 1056 24987 1088 25019
rect 1128 24987 1160 25019
rect 1200 24987 1232 25019
rect 1272 24987 1304 25019
rect 1344 24987 1376 25019
rect 1416 24987 1448 25019
rect 1488 24987 1520 25019
rect 1560 24987 1592 25019
rect 1632 24987 1664 25019
rect 1704 24987 1736 25019
rect 1776 24987 1808 25019
rect 1848 24987 1880 25019
rect 120 24915 152 24947
rect 192 24915 224 24947
rect 264 24915 296 24947
rect 336 24915 368 24947
rect 408 24915 440 24947
rect 480 24915 512 24947
rect 552 24915 584 24947
rect 624 24915 656 24947
rect 696 24915 728 24947
rect 768 24915 800 24947
rect 840 24915 872 24947
rect 912 24915 944 24947
rect 984 24915 1016 24947
rect 1056 24915 1088 24947
rect 1128 24915 1160 24947
rect 1200 24915 1232 24947
rect 1272 24915 1304 24947
rect 1344 24915 1376 24947
rect 1416 24915 1448 24947
rect 1488 24915 1520 24947
rect 1560 24915 1592 24947
rect 1632 24915 1664 24947
rect 1704 24915 1736 24947
rect 1776 24915 1808 24947
rect 1848 24915 1880 24947
rect 120 24843 152 24875
rect 192 24843 224 24875
rect 264 24843 296 24875
rect 336 24843 368 24875
rect 408 24843 440 24875
rect 480 24843 512 24875
rect 552 24843 584 24875
rect 624 24843 656 24875
rect 696 24843 728 24875
rect 768 24843 800 24875
rect 840 24843 872 24875
rect 912 24843 944 24875
rect 984 24843 1016 24875
rect 1056 24843 1088 24875
rect 1128 24843 1160 24875
rect 1200 24843 1232 24875
rect 1272 24843 1304 24875
rect 1344 24843 1376 24875
rect 1416 24843 1448 24875
rect 1488 24843 1520 24875
rect 1560 24843 1592 24875
rect 1632 24843 1664 24875
rect 1704 24843 1736 24875
rect 1776 24843 1808 24875
rect 1848 24843 1880 24875
rect 120 24771 152 24803
rect 192 24771 224 24803
rect 264 24771 296 24803
rect 336 24771 368 24803
rect 408 24771 440 24803
rect 480 24771 512 24803
rect 552 24771 584 24803
rect 624 24771 656 24803
rect 696 24771 728 24803
rect 768 24771 800 24803
rect 840 24771 872 24803
rect 912 24771 944 24803
rect 984 24771 1016 24803
rect 1056 24771 1088 24803
rect 1128 24771 1160 24803
rect 1200 24771 1232 24803
rect 1272 24771 1304 24803
rect 1344 24771 1376 24803
rect 1416 24771 1448 24803
rect 1488 24771 1520 24803
rect 1560 24771 1592 24803
rect 1632 24771 1664 24803
rect 1704 24771 1736 24803
rect 1776 24771 1808 24803
rect 1848 24771 1880 24803
rect 120 24699 152 24731
rect 192 24699 224 24731
rect 264 24699 296 24731
rect 336 24699 368 24731
rect 408 24699 440 24731
rect 480 24699 512 24731
rect 552 24699 584 24731
rect 624 24699 656 24731
rect 696 24699 728 24731
rect 768 24699 800 24731
rect 840 24699 872 24731
rect 912 24699 944 24731
rect 984 24699 1016 24731
rect 1056 24699 1088 24731
rect 1128 24699 1160 24731
rect 1200 24699 1232 24731
rect 1272 24699 1304 24731
rect 1344 24699 1376 24731
rect 1416 24699 1448 24731
rect 1488 24699 1520 24731
rect 1560 24699 1592 24731
rect 1632 24699 1664 24731
rect 1704 24699 1736 24731
rect 1776 24699 1808 24731
rect 1848 24699 1880 24731
rect 120 24627 152 24659
rect 192 24627 224 24659
rect 264 24627 296 24659
rect 336 24627 368 24659
rect 408 24627 440 24659
rect 480 24627 512 24659
rect 552 24627 584 24659
rect 624 24627 656 24659
rect 696 24627 728 24659
rect 768 24627 800 24659
rect 840 24627 872 24659
rect 912 24627 944 24659
rect 984 24627 1016 24659
rect 1056 24627 1088 24659
rect 1128 24627 1160 24659
rect 1200 24627 1232 24659
rect 1272 24627 1304 24659
rect 1344 24627 1376 24659
rect 1416 24627 1448 24659
rect 1488 24627 1520 24659
rect 1560 24627 1592 24659
rect 1632 24627 1664 24659
rect 1704 24627 1736 24659
rect 1776 24627 1808 24659
rect 1848 24627 1880 24659
rect 120 24555 152 24587
rect 192 24555 224 24587
rect 264 24555 296 24587
rect 336 24555 368 24587
rect 408 24555 440 24587
rect 480 24555 512 24587
rect 552 24555 584 24587
rect 624 24555 656 24587
rect 696 24555 728 24587
rect 768 24555 800 24587
rect 840 24555 872 24587
rect 912 24555 944 24587
rect 984 24555 1016 24587
rect 1056 24555 1088 24587
rect 1128 24555 1160 24587
rect 1200 24555 1232 24587
rect 1272 24555 1304 24587
rect 1344 24555 1376 24587
rect 1416 24555 1448 24587
rect 1488 24555 1520 24587
rect 1560 24555 1592 24587
rect 1632 24555 1664 24587
rect 1704 24555 1736 24587
rect 1776 24555 1808 24587
rect 1848 24555 1880 24587
rect 120 24483 152 24515
rect 192 24483 224 24515
rect 264 24483 296 24515
rect 336 24483 368 24515
rect 408 24483 440 24515
rect 480 24483 512 24515
rect 552 24483 584 24515
rect 624 24483 656 24515
rect 696 24483 728 24515
rect 768 24483 800 24515
rect 840 24483 872 24515
rect 912 24483 944 24515
rect 984 24483 1016 24515
rect 1056 24483 1088 24515
rect 1128 24483 1160 24515
rect 1200 24483 1232 24515
rect 1272 24483 1304 24515
rect 1344 24483 1376 24515
rect 1416 24483 1448 24515
rect 1488 24483 1520 24515
rect 1560 24483 1592 24515
rect 1632 24483 1664 24515
rect 1704 24483 1736 24515
rect 1776 24483 1808 24515
rect 1848 24483 1880 24515
rect 120 24411 152 24443
rect 192 24411 224 24443
rect 264 24411 296 24443
rect 336 24411 368 24443
rect 408 24411 440 24443
rect 480 24411 512 24443
rect 552 24411 584 24443
rect 624 24411 656 24443
rect 696 24411 728 24443
rect 768 24411 800 24443
rect 840 24411 872 24443
rect 912 24411 944 24443
rect 984 24411 1016 24443
rect 1056 24411 1088 24443
rect 1128 24411 1160 24443
rect 1200 24411 1232 24443
rect 1272 24411 1304 24443
rect 1344 24411 1376 24443
rect 1416 24411 1448 24443
rect 1488 24411 1520 24443
rect 1560 24411 1592 24443
rect 1632 24411 1664 24443
rect 1704 24411 1736 24443
rect 1776 24411 1808 24443
rect 1848 24411 1880 24443
rect 120 24339 152 24371
rect 192 24339 224 24371
rect 264 24339 296 24371
rect 336 24339 368 24371
rect 408 24339 440 24371
rect 480 24339 512 24371
rect 552 24339 584 24371
rect 624 24339 656 24371
rect 696 24339 728 24371
rect 768 24339 800 24371
rect 840 24339 872 24371
rect 912 24339 944 24371
rect 984 24339 1016 24371
rect 1056 24339 1088 24371
rect 1128 24339 1160 24371
rect 1200 24339 1232 24371
rect 1272 24339 1304 24371
rect 1344 24339 1376 24371
rect 1416 24339 1448 24371
rect 1488 24339 1520 24371
rect 1560 24339 1592 24371
rect 1632 24339 1664 24371
rect 1704 24339 1736 24371
rect 1776 24339 1808 24371
rect 1848 24339 1880 24371
rect 120 24267 152 24299
rect 192 24267 224 24299
rect 264 24267 296 24299
rect 336 24267 368 24299
rect 408 24267 440 24299
rect 480 24267 512 24299
rect 552 24267 584 24299
rect 624 24267 656 24299
rect 696 24267 728 24299
rect 768 24267 800 24299
rect 840 24267 872 24299
rect 912 24267 944 24299
rect 984 24267 1016 24299
rect 1056 24267 1088 24299
rect 1128 24267 1160 24299
rect 1200 24267 1232 24299
rect 1272 24267 1304 24299
rect 1344 24267 1376 24299
rect 1416 24267 1448 24299
rect 1488 24267 1520 24299
rect 1560 24267 1592 24299
rect 1632 24267 1664 24299
rect 1704 24267 1736 24299
rect 1776 24267 1808 24299
rect 1848 24267 1880 24299
rect 120 24195 152 24227
rect 192 24195 224 24227
rect 264 24195 296 24227
rect 336 24195 368 24227
rect 408 24195 440 24227
rect 480 24195 512 24227
rect 552 24195 584 24227
rect 624 24195 656 24227
rect 696 24195 728 24227
rect 768 24195 800 24227
rect 840 24195 872 24227
rect 912 24195 944 24227
rect 984 24195 1016 24227
rect 1056 24195 1088 24227
rect 1128 24195 1160 24227
rect 1200 24195 1232 24227
rect 1272 24195 1304 24227
rect 1344 24195 1376 24227
rect 1416 24195 1448 24227
rect 1488 24195 1520 24227
rect 1560 24195 1592 24227
rect 1632 24195 1664 24227
rect 1704 24195 1736 24227
rect 1776 24195 1808 24227
rect 1848 24195 1880 24227
rect 120 24123 152 24155
rect 192 24123 224 24155
rect 264 24123 296 24155
rect 336 24123 368 24155
rect 408 24123 440 24155
rect 480 24123 512 24155
rect 552 24123 584 24155
rect 624 24123 656 24155
rect 696 24123 728 24155
rect 768 24123 800 24155
rect 840 24123 872 24155
rect 912 24123 944 24155
rect 984 24123 1016 24155
rect 1056 24123 1088 24155
rect 1128 24123 1160 24155
rect 1200 24123 1232 24155
rect 1272 24123 1304 24155
rect 1344 24123 1376 24155
rect 1416 24123 1448 24155
rect 1488 24123 1520 24155
rect 1560 24123 1592 24155
rect 1632 24123 1664 24155
rect 1704 24123 1736 24155
rect 1776 24123 1808 24155
rect 1848 24123 1880 24155
rect 120 24051 152 24083
rect 192 24051 224 24083
rect 264 24051 296 24083
rect 336 24051 368 24083
rect 408 24051 440 24083
rect 480 24051 512 24083
rect 552 24051 584 24083
rect 624 24051 656 24083
rect 696 24051 728 24083
rect 768 24051 800 24083
rect 840 24051 872 24083
rect 912 24051 944 24083
rect 984 24051 1016 24083
rect 1056 24051 1088 24083
rect 1128 24051 1160 24083
rect 1200 24051 1232 24083
rect 1272 24051 1304 24083
rect 1344 24051 1376 24083
rect 1416 24051 1448 24083
rect 1488 24051 1520 24083
rect 1560 24051 1592 24083
rect 1632 24051 1664 24083
rect 1704 24051 1736 24083
rect 1776 24051 1808 24083
rect 1848 24051 1880 24083
rect 120 23979 152 24011
rect 192 23979 224 24011
rect 264 23979 296 24011
rect 336 23979 368 24011
rect 408 23979 440 24011
rect 480 23979 512 24011
rect 552 23979 584 24011
rect 624 23979 656 24011
rect 696 23979 728 24011
rect 768 23979 800 24011
rect 840 23979 872 24011
rect 912 23979 944 24011
rect 984 23979 1016 24011
rect 1056 23979 1088 24011
rect 1128 23979 1160 24011
rect 1200 23979 1232 24011
rect 1272 23979 1304 24011
rect 1344 23979 1376 24011
rect 1416 23979 1448 24011
rect 1488 23979 1520 24011
rect 1560 23979 1592 24011
rect 1632 23979 1664 24011
rect 1704 23979 1736 24011
rect 1776 23979 1808 24011
rect 1848 23979 1880 24011
rect 120 23907 152 23939
rect 192 23907 224 23939
rect 264 23907 296 23939
rect 336 23907 368 23939
rect 408 23907 440 23939
rect 480 23907 512 23939
rect 552 23907 584 23939
rect 624 23907 656 23939
rect 696 23907 728 23939
rect 768 23907 800 23939
rect 840 23907 872 23939
rect 912 23907 944 23939
rect 984 23907 1016 23939
rect 1056 23907 1088 23939
rect 1128 23907 1160 23939
rect 1200 23907 1232 23939
rect 1272 23907 1304 23939
rect 1344 23907 1376 23939
rect 1416 23907 1448 23939
rect 1488 23907 1520 23939
rect 1560 23907 1592 23939
rect 1632 23907 1664 23939
rect 1704 23907 1736 23939
rect 1776 23907 1808 23939
rect 1848 23907 1880 23939
rect 120 23835 152 23867
rect 192 23835 224 23867
rect 264 23835 296 23867
rect 336 23835 368 23867
rect 408 23835 440 23867
rect 480 23835 512 23867
rect 552 23835 584 23867
rect 624 23835 656 23867
rect 696 23835 728 23867
rect 768 23835 800 23867
rect 840 23835 872 23867
rect 912 23835 944 23867
rect 984 23835 1016 23867
rect 1056 23835 1088 23867
rect 1128 23835 1160 23867
rect 1200 23835 1232 23867
rect 1272 23835 1304 23867
rect 1344 23835 1376 23867
rect 1416 23835 1448 23867
rect 1488 23835 1520 23867
rect 1560 23835 1592 23867
rect 1632 23835 1664 23867
rect 1704 23835 1736 23867
rect 1776 23835 1808 23867
rect 1848 23835 1880 23867
rect 120 23763 152 23795
rect 192 23763 224 23795
rect 264 23763 296 23795
rect 336 23763 368 23795
rect 408 23763 440 23795
rect 480 23763 512 23795
rect 552 23763 584 23795
rect 624 23763 656 23795
rect 696 23763 728 23795
rect 768 23763 800 23795
rect 840 23763 872 23795
rect 912 23763 944 23795
rect 984 23763 1016 23795
rect 1056 23763 1088 23795
rect 1128 23763 1160 23795
rect 1200 23763 1232 23795
rect 1272 23763 1304 23795
rect 1344 23763 1376 23795
rect 1416 23763 1448 23795
rect 1488 23763 1520 23795
rect 1560 23763 1592 23795
rect 1632 23763 1664 23795
rect 1704 23763 1736 23795
rect 1776 23763 1808 23795
rect 1848 23763 1880 23795
rect 120 23691 152 23723
rect 192 23691 224 23723
rect 264 23691 296 23723
rect 336 23691 368 23723
rect 408 23691 440 23723
rect 480 23691 512 23723
rect 552 23691 584 23723
rect 624 23691 656 23723
rect 696 23691 728 23723
rect 768 23691 800 23723
rect 840 23691 872 23723
rect 912 23691 944 23723
rect 984 23691 1016 23723
rect 1056 23691 1088 23723
rect 1128 23691 1160 23723
rect 1200 23691 1232 23723
rect 1272 23691 1304 23723
rect 1344 23691 1376 23723
rect 1416 23691 1448 23723
rect 1488 23691 1520 23723
rect 1560 23691 1592 23723
rect 1632 23691 1664 23723
rect 1704 23691 1736 23723
rect 1776 23691 1808 23723
rect 1848 23691 1880 23723
rect 120 23619 152 23651
rect 192 23619 224 23651
rect 264 23619 296 23651
rect 336 23619 368 23651
rect 408 23619 440 23651
rect 480 23619 512 23651
rect 552 23619 584 23651
rect 624 23619 656 23651
rect 696 23619 728 23651
rect 768 23619 800 23651
rect 840 23619 872 23651
rect 912 23619 944 23651
rect 984 23619 1016 23651
rect 1056 23619 1088 23651
rect 1128 23619 1160 23651
rect 1200 23619 1232 23651
rect 1272 23619 1304 23651
rect 1344 23619 1376 23651
rect 1416 23619 1448 23651
rect 1488 23619 1520 23651
rect 1560 23619 1592 23651
rect 1632 23619 1664 23651
rect 1704 23619 1736 23651
rect 1776 23619 1808 23651
rect 1848 23619 1880 23651
rect 120 23547 152 23579
rect 192 23547 224 23579
rect 264 23547 296 23579
rect 336 23547 368 23579
rect 408 23547 440 23579
rect 480 23547 512 23579
rect 552 23547 584 23579
rect 624 23547 656 23579
rect 696 23547 728 23579
rect 768 23547 800 23579
rect 840 23547 872 23579
rect 912 23547 944 23579
rect 984 23547 1016 23579
rect 1056 23547 1088 23579
rect 1128 23547 1160 23579
rect 1200 23547 1232 23579
rect 1272 23547 1304 23579
rect 1344 23547 1376 23579
rect 1416 23547 1448 23579
rect 1488 23547 1520 23579
rect 1560 23547 1592 23579
rect 1632 23547 1664 23579
rect 1704 23547 1736 23579
rect 1776 23547 1808 23579
rect 1848 23547 1880 23579
rect 120 23475 152 23507
rect 192 23475 224 23507
rect 264 23475 296 23507
rect 336 23475 368 23507
rect 408 23475 440 23507
rect 480 23475 512 23507
rect 552 23475 584 23507
rect 624 23475 656 23507
rect 696 23475 728 23507
rect 768 23475 800 23507
rect 840 23475 872 23507
rect 912 23475 944 23507
rect 984 23475 1016 23507
rect 1056 23475 1088 23507
rect 1128 23475 1160 23507
rect 1200 23475 1232 23507
rect 1272 23475 1304 23507
rect 1344 23475 1376 23507
rect 1416 23475 1448 23507
rect 1488 23475 1520 23507
rect 1560 23475 1592 23507
rect 1632 23475 1664 23507
rect 1704 23475 1736 23507
rect 1776 23475 1808 23507
rect 1848 23475 1880 23507
rect 120 23403 152 23435
rect 192 23403 224 23435
rect 264 23403 296 23435
rect 336 23403 368 23435
rect 408 23403 440 23435
rect 480 23403 512 23435
rect 552 23403 584 23435
rect 624 23403 656 23435
rect 696 23403 728 23435
rect 768 23403 800 23435
rect 840 23403 872 23435
rect 912 23403 944 23435
rect 984 23403 1016 23435
rect 1056 23403 1088 23435
rect 1128 23403 1160 23435
rect 1200 23403 1232 23435
rect 1272 23403 1304 23435
rect 1344 23403 1376 23435
rect 1416 23403 1448 23435
rect 1488 23403 1520 23435
rect 1560 23403 1592 23435
rect 1632 23403 1664 23435
rect 1704 23403 1736 23435
rect 1776 23403 1808 23435
rect 1848 23403 1880 23435
rect 120 23331 152 23363
rect 192 23331 224 23363
rect 264 23331 296 23363
rect 336 23331 368 23363
rect 408 23331 440 23363
rect 480 23331 512 23363
rect 552 23331 584 23363
rect 624 23331 656 23363
rect 696 23331 728 23363
rect 768 23331 800 23363
rect 840 23331 872 23363
rect 912 23331 944 23363
rect 984 23331 1016 23363
rect 1056 23331 1088 23363
rect 1128 23331 1160 23363
rect 1200 23331 1232 23363
rect 1272 23331 1304 23363
rect 1344 23331 1376 23363
rect 1416 23331 1448 23363
rect 1488 23331 1520 23363
rect 1560 23331 1592 23363
rect 1632 23331 1664 23363
rect 1704 23331 1736 23363
rect 1776 23331 1808 23363
rect 1848 23331 1880 23363
rect 120 23259 152 23291
rect 192 23259 224 23291
rect 264 23259 296 23291
rect 336 23259 368 23291
rect 408 23259 440 23291
rect 480 23259 512 23291
rect 552 23259 584 23291
rect 624 23259 656 23291
rect 696 23259 728 23291
rect 768 23259 800 23291
rect 840 23259 872 23291
rect 912 23259 944 23291
rect 984 23259 1016 23291
rect 1056 23259 1088 23291
rect 1128 23259 1160 23291
rect 1200 23259 1232 23291
rect 1272 23259 1304 23291
rect 1344 23259 1376 23291
rect 1416 23259 1448 23291
rect 1488 23259 1520 23291
rect 1560 23259 1592 23291
rect 1632 23259 1664 23291
rect 1704 23259 1736 23291
rect 1776 23259 1808 23291
rect 1848 23259 1880 23291
rect 120 23187 152 23219
rect 192 23187 224 23219
rect 264 23187 296 23219
rect 336 23187 368 23219
rect 408 23187 440 23219
rect 480 23187 512 23219
rect 552 23187 584 23219
rect 624 23187 656 23219
rect 696 23187 728 23219
rect 768 23187 800 23219
rect 840 23187 872 23219
rect 912 23187 944 23219
rect 984 23187 1016 23219
rect 1056 23187 1088 23219
rect 1128 23187 1160 23219
rect 1200 23187 1232 23219
rect 1272 23187 1304 23219
rect 1344 23187 1376 23219
rect 1416 23187 1448 23219
rect 1488 23187 1520 23219
rect 1560 23187 1592 23219
rect 1632 23187 1664 23219
rect 1704 23187 1736 23219
rect 1776 23187 1808 23219
rect 1848 23187 1880 23219
rect 192 22842 224 22874
rect 264 22842 296 22874
rect 336 22842 368 22874
rect 408 22842 440 22874
rect 480 22842 512 22874
rect 552 22842 584 22874
rect 624 22842 656 22874
rect 696 22842 728 22874
rect 768 22842 800 22874
rect 840 22842 872 22874
rect 912 22842 944 22874
rect 984 22842 1016 22874
rect 1056 22842 1088 22874
rect 1128 22842 1160 22874
rect 1200 22842 1232 22874
rect 1272 22842 1304 22874
rect 1344 22842 1376 22874
rect 1416 22842 1448 22874
rect 1488 22842 1520 22874
rect 1560 22842 1592 22874
rect 1632 22842 1664 22874
rect 1704 22842 1736 22874
rect 1776 22842 1808 22874
rect 1848 22842 1880 22874
rect 120 22770 152 22802
rect 192 22770 224 22802
rect 264 22770 296 22802
rect 336 22770 368 22802
rect 408 22770 440 22802
rect 480 22770 512 22802
rect 552 22770 584 22802
rect 624 22770 656 22802
rect 696 22770 728 22802
rect 768 22770 800 22802
rect 840 22770 872 22802
rect 912 22770 944 22802
rect 984 22770 1016 22802
rect 1056 22770 1088 22802
rect 1128 22770 1160 22802
rect 1200 22770 1232 22802
rect 1272 22770 1304 22802
rect 1344 22770 1376 22802
rect 1416 22770 1448 22802
rect 1488 22770 1520 22802
rect 1560 22770 1592 22802
rect 1632 22770 1664 22802
rect 1704 22770 1736 22802
rect 1776 22770 1808 22802
rect 1848 22770 1880 22802
rect 120 22698 152 22730
rect 192 22698 224 22730
rect 264 22698 296 22730
rect 336 22698 368 22730
rect 408 22698 440 22730
rect 480 22698 512 22730
rect 552 22698 584 22730
rect 624 22698 656 22730
rect 696 22698 728 22730
rect 768 22698 800 22730
rect 840 22698 872 22730
rect 912 22698 944 22730
rect 984 22698 1016 22730
rect 1056 22698 1088 22730
rect 1128 22698 1160 22730
rect 1200 22698 1232 22730
rect 1272 22698 1304 22730
rect 1344 22698 1376 22730
rect 1416 22698 1448 22730
rect 1488 22698 1520 22730
rect 1560 22698 1592 22730
rect 1632 22698 1664 22730
rect 1704 22698 1736 22730
rect 1776 22698 1808 22730
rect 1848 22698 1880 22730
rect 120 22626 152 22658
rect 192 22626 224 22658
rect 264 22626 296 22658
rect 336 22626 368 22658
rect 408 22626 440 22658
rect 480 22626 512 22658
rect 552 22626 584 22658
rect 624 22626 656 22658
rect 696 22626 728 22658
rect 768 22626 800 22658
rect 840 22626 872 22658
rect 912 22626 944 22658
rect 984 22626 1016 22658
rect 1056 22626 1088 22658
rect 1128 22626 1160 22658
rect 1200 22626 1232 22658
rect 1272 22626 1304 22658
rect 1344 22626 1376 22658
rect 1416 22626 1448 22658
rect 1488 22626 1520 22658
rect 1560 22626 1592 22658
rect 1632 22626 1664 22658
rect 1704 22626 1736 22658
rect 1776 22626 1808 22658
rect 1848 22626 1880 22658
rect 120 22554 152 22586
rect 192 22554 224 22586
rect 264 22554 296 22586
rect 336 22554 368 22586
rect 408 22554 440 22586
rect 480 22554 512 22586
rect 552 22554 584 22586
rect 624 22554 656 22586
rect 696 22554 728 22586
rect 768 22554 800 22586
rect 840 22554 872 22586
rect 912 22554 944 22586
rect 984 22554 1016 22586
rect 1056 22554 1088 22586
rect 1128 22554 1160 22586
rect 1200 22554 1232 22586
rect 1272 22554 1304 22586
rect 1344 22554 1376 22586
rect 1416 22554 1448 22586
rect 1488 22554 1520 22586
rect 1560 22554 1592 22586
rect 1632 22554 1664 22586
rect 1704 22554 1736 22586
rect 1776 22554 1808 22586
rect 1848 22554 1880 22586
rect 120 22482 152 22514
rect 192 22482 224 22514
rect 264 22482 296 22514
rect 336 22482 368 22514
rect 408 22482 440 22514
rect 480 22482 512 22514
rect 552 22482 584 22514
rect 624 22482 656 22514
rect 696 22482 728 22514
rect 768 22482 800 22514
rect 840 22482 872 22514
rect 912 22482 944 22514
rect 984 22482 1016 22514
rect 1056 22482 1088 22514
rect 1128 22482 1160 22514
rect 1200 22482 1232 22514
rect 1272 22482 1304 22514
rect 1344 22482 1376 22514
rect 1416 22482 1448 22514
rect 1488 22482 1520 22514
rect 1560 22482 1592 22514
rect 1632 22482 1664 22514
rect 1704 22482 1736 22514
rect 1776 22482 1808 22514
rect 1848 22482 1880 22514
rect 120 22410 152 22442
rect 192 22410 224 22442
rect 264 22410 296 22442
rect 336 22410 368 22442
rect 408 22410 440 22442
rect 480 22410 512 22442
rect 552 22410 584 22442
rect 624 22410 656 22442
rect 696 22410 728 22442
rect 768 22410 800 22442
rect 840 22410 872 22442
rect 912 22410 944 22442
rect 984 22410 1016 22442
rect 1056 22410 1088 22442
rect 1128 22410 1160 22442
rect 1200 22410 1232 22442
rect 1272 22410 1304 22442
rect 1344 22410 1376 22442
rect 1416 22410 1448 22442
rect 1488 22410 1520 22442
rect 1560 22410 1592 22442
rect 1632 22410 1664 22442
rect 1704 22410 1736 22442
rect 1776 22410 1808 22442
rect 1848 22410 1880 22442
rect 120 22338 152 22370
rect 192 22338 224 22370
rect 264 22338 296 22370
rect 336 22338 368 22370
rect 408 22338 440 22370
rect 480 22338 512 22370
rect 552 22338 584 22370
rect 624 22338 656 22370
rect 696 22338 728 22370
rect 768 22338 800 22370
rect 840 22338 872 22370
rect 912 22338 944 22370
rect 984 22338 1016 22370
rect 1056 22338 1088 22370
rect 1128 22338 1160 22370
rect 1200 22338 1232 22370
rect 1272 22338 1304 22370
rect 1344 22338 1376 22370
rect 1416 22338 1448 22370
rect 1488 22338 1520 22370
rect 1560 22338 1592 22370
rect 1632 22338 1664 22370
rect 1704 22338 1736 22370
rect 1776 22338 1808 22370
rect 1848 22338 1880 22370
rect 120 22266 152 22298
rect 192 22266 224 22298
rect 264 22266 296 22298
rect 336 22266 368 22298
rect 408 22266 440 22298
rect 480 22266 512 22298
rect 552 22266 584 22298
rect 624 22266 656 22298
rect 696 22266 728 22298
rect 768 22266 800 22298
rect 840 22266 872 22298
rect 912 22266 944 22298
rect 984 22266 1016 22298
rect 1056 22266 1088 22298
rect 1128 22266 1160 22298
rect 1200 22266 1232 22298
rect 1272 22266 1304 22298
rect 1344 22266 1376 22298
rect 1416 22266 1448 22298
rect 1488 22266 1520 22298
rect 1560 22266 1592 22298
rect 1632 22266 1664 22298
rect 1704 22266 1736 22298
rect 1776 22266 1808 22298
rect 1848 22266 1880 22298
rect 120 22194 152 22226
rect 192 22194 224 22226
rect 264 22194 296 22226
rect 336 22194 368 22226
rect 408 22194 440 22226
rect 480 22194 512 22226
rect 552 22194 584 22226
rect 624 22194 656 22226
rect 696 22194 728 22226
rect 768 22194 800 22226
rect 840 22194 872 22226
rect 912 22194 944 22226
rect 984 22194 1016 22226
rect 1056 22194 1088 22226
rect 1128 22194 1160 22226
rect 1200 22194 1232 22226
rect 1272 22194 1304 22226
rect 1344 22194 1376 22226
rect 1416 22194 1448 22226
rect 1488 22194 1520 22226
rect 1560 22194 1592 22226
rect 1632 22194 1664 22226
rect 1704 22194 1736 22226
rect 1776 22194 1808 22226
rect 1848 22194 1880 22226
rect 120 22122 152 22154
rect 192 22122 224 22154
rect 264 22122 296 22154
rect 336 22122 368 22154
rect 408 22122 440 22154
rect 480 22122 512 22154
rect 552 22122 584 22154
rect 624 22122 656 22154
rect 696 22122 728 22154
rect 768 22122 800 22154
rect 840 22122 872 22154
rect 912 22122 944 22154
rect 984 22122 1016 22154
rect 1056 22122 1088 22154
rect 1128 22122 1160 22154
rect 1200 22122 1232 22154
rect 1272 22122 1304 22154
rect 1344 22122 1376 22154
rect 1416 22122 1448 22154
rect 1488 22122 1520 22154
rect 1560 22122 1592 22154
rect 1632 22122 1664 22154
rect 1704 22122 1736 22154
rect 1776 22122 1808 22154
rect 1848 22122 1880 22154
rect 120 22050 152 22082
rect 192 22050 224 22082
rect 264 22050 296 22082
rect 336 22050 368 22082
rect 408 22050 440 22082
rect 480 22050 512 22082
rect 552 22050 584 22082
rect 624 22050 656 22082
rect 696 22050 728 22082
rect 768 22050 800 22082
rect 840 22050 872 22082
rect 912 22050 944 22082
rect 984 22050 1016 22082
rect 1056 22050 1088 22082
rect 1128 22050 1160 22082
rect 1200 22050 1232 22082
rect 1272 22050 1304 22082
rect 1344 22050 1376 22082
rect 1416 22050 1448 22082
rect 1488 22050 1520 22082
rect 1560 22050 1592 22082
rect 1632 22050 1664 22082
rect 1704 22050 1736 22082
rect 1776 22050 1808 22082
rect 1848 22050 1880 22082
rect 120 21978 152 22010
rect 192 21978 224 22010
rect 264 21978 296 22010
rect 336 21978 368 22010
rect 408 21978 440 22010
rect 480 21978 512 22010
rect 552 21978 584 22010
rect 624 21978 656 22010
rect 696 21978 728 22010
rect 768 21978 800 22010
rect 840 21978 872 22010
rect 912 21978 944 22010
rect 984 21978 1016 22010
rect 1056 21978 1088 22010
rect 1128 21978 1160 22010
rect 1200 21978 1232 22010
rect 1272 21978 1304 22010
rect 1344 21978 1376 22010
rect 1416 21978 1448 22010
rect 1488 21978 1520 22010
rect 1560 21978 1592 22010
rect 1632 21978 1664 22010
rect 1704 21978 1736 22010
rect 1776 21978 1808 22010
rect 1848 21978 1880 22010
rect 120 21906 152 21938
rect 192 21906 224 21938
rect 264 21906 296 21938
rect 336 21906 368 21938
rect 408 21906 440 21938
rect 480 21906 512 21938
rect 552 21906 584 21938
rect 624 21906 656 21938
rect 696 21906 728 21938
rect 768 21906 800 21938
rect 840 21906 872 21938
rect 912 21906 944 21938
rect 984 21906 1016 21938
rect 1056 21906 1088 21938
rect 1128 21906 1160 21938
rect 1200 21906 1232 21938
rect 1272 21906 1304 21938
rect 1344 21906 1376 21938
rect 1416 21906 1448 21938
rect 1488 21906 1520 21938
rect 1560 21906 1592 21938
rect 1632 21906 1664 21938
rect 1704 21906 1736 21938
rect 1776 21906 1808 21938
rect 1848 21906 1880 21938
rect 120 21834 152 21866
rect 192 21834 224 21866
rect 264 21834 296 21866
rect 336 21834 368 21866
rect 408 21834 440 21866
rect 480 21834 512 21866
rect 552 21834 584 21866
rect 624 21834 656 21866
rect 696 21834 728 21866
rect 768 21834 800 21866
rect 840 21834 872 21866
rect 912 21834 944 21866
rect 984 21834 1016 21866
rect 1056 21834 1088 21866
rect 1128 21834 1160 21866
rect 1200 21834 1232 21866
rect 1272 21834 1304 21866
rect 1344 21834 1376 21866
rect 1416 21834 1448 21866
rect 1488 21834 1520 21866
rect 1560 21834 1592 21866
rect 1632 21834 1664 21866
rect 1704 21834 1736 21866
rect 1776 21834 1808 21866
rect 1848 21834 1880 21866
rect 120 21762 152 21794
rect 192 21762 224 21794
rect 264 21762 296 21794
rect 336 21762 368 21794
rect 408 21762 440 21794
rect 480 21762 512 21794
rect 552 21762 584 21794
rect 624 21762 656 21794
rect 696 21762 728 21794
rect 768 21762 800 21794
rect 840 21762 872 21794
rect 912 21762 944 21794
rect 984 21762 1016 21794
rect 1056 21762 1088 21794
rect 1128 21762 1160 21794
rect 1200 21762 1232 21794
rect 1272 21762 1304 21794
rect 1344 21762 1376 21794
rect 1416 21762 1448 21794
rect 1488 21762 1520 21794
rect 1560 21762 1592 21794
rect 1632 21762 1664 21794
rect 1704 21762 1736 21794
rect 1776 21762 1808 21794
rect 1848 21762 1880 21794
rect 120 21690 152 21722
rect 192 21690 224 21722
rect 264 21690 296 21722
rect 336 21690 368 21722
rect 408 21690 440 21722
rect 480 21690 512 21722
rect 552 21690 584 21722
rect 624 21690 656 21722
rect 696 21690 728 21722
rect 768 21690 800 21722
rect 840 21690 872 21722
rect 912 21690 944 21722
rect 984 21690 1016 21722
rect 1056 21690 1088 21722
rect 1128 21690 1160 21722
rect 1200 21690 1232 21722
rect 1272 21690 1304 21722
rect 1344 21690 1376 21722
rect 1416 21690 1448 21722
rect 1488 21690 1520 21722
rect 1560 21690 1592 21722
rect 1632 21690 1664 21722
rect 1704 21690 1736 21722
rect 1776 21690 1808 21722
rect 1848 21690 1880 21722
rect 120 21618 152 21650
rect 192 21618 224 21650
rect 264 21618 296 21650
rect 336 21618 368 21650
rect 408 21618 440 21650
rect 480 21618 512 21650
rect 552 21618 584 21650
rect 624 21618 656 21650
rect 696 21618 728 21650
rect 768 21618 800 21650
rect 840 21618 872 21650
rect 912 21618 944 21650
rect 984 21618 1016 21650
rect 1056 21618 1088 21650
rect 1128 21618 1160 21650
rect 1200 21618 1232 21650
rect 1272 21618 1304 21650
rect 1344 21618 1376 21650
rect 1416 21618 1448 21650
rect 1488 21618 1520 21650
rect 1560 21618 1592 21650
rect 1632 21618 1664 21650
rect 1704 21618 1736 21650
rect 1776 21618 1808 21650
rect 1848 21618 1880 21650
rect 120 21546 152 21578
rect 192 21546 224 21578
rect 264 21546 296 21578
rect 336 21546 368 21578
rect 408 21546 440 21578
rect 480 21546 512 21578
rect 552 21546 584 21578
rect 624 21546 656 21578
rect 696 21546 728 21578
rect 768 21546 800 21578
rect 840 21546 872 21578
rect 912 21546 944 21578
rect 984 21546 1016 21578
rect 1056 21546 1088 21578
rect 1128 21546 1160 21578
rect 1200 21546 1232 21578
rect 1272 21546 1304 21578
rect 1344 21546 1376 21578
rect 1416 21546 1448 21578
rect 1488 21546 1520 21578
rect 1560 21546 1592 21578
rect 1632 21546 1664 21578
rect 1704 21546 1736 21578
rect 1776 21546 1808 21578
rect 1848 21546 1880 21578
rect 120 21474 152 21506
rect 192 21474 224 21506
rect 264 21474 296 21506
rect 336 21474 368 21506
rect 408 21474 440 21506
rect 480 21474 512 21506
rect 552 21474 584 21506
rect 624 21474 656 21506
rect 696 21474 728 21506
rect 768 21474 800 21506
rect 840 21474 872 21506
rect 912 21474 944 21506
rect 984 21474 1016 21506
rect 1056 21474 1088 21506
rect 1128 21474 1160 21506
rect 1200 21474 1232 21506
rect 1272 21474 1304 21506
rect 1344 21474 1376 21506
rect 1416 21474 1448 21506
rect 1488 21474 1520 21506
rect 1560 21474 1592 21506
rect 1632 21474 1664 21506
rect 1704 21474 1736 21506
rect 1776 21474 1808 21506
rect 1848 21474 1880 21506
rect 120 21402 152 21434
rect 192 21402 224 21434
rect 264 21402 296 21434
rect 336 21402 368 21434
rect 408 21402 440 21434
rect 480 21402 512 21434
rect 552 21402 584 21434
rect 624 21402 656 21434
rect 696 21402 728 21434
rect 768 21402 800 21434
rect 840 21402 872 21434
rect 912 21402 944 21434
rect 984 21402 1016 21434
rect 1056 21402 1088 21434
rect 1128 21402 1160 21434
rect 1200 21402 1232 21434
rect 1272 21402 1304 21434
rect 1344 21402 1376 21434
rect 1416 21402 1448 21434
rect 1488 21402 1520 21434
rect 1560 21402 1592 21434
rect 1632 21402 1664 21434
rect 1704 21402 1736 21434
rect 1776 21402 1808 21434
rect 1848 21402 1880 21434
rect 120 21330 152 21362
rect 192 21330 224 21362
rect 264 21330 296 21362
rect 336 21330 368 21362
rect 408 21330 440 21362
rect 480 21330 512 21362
rect 552 21330 584 21362
rect 624 21330 656 21362
rect 696 21330 728 21362
rect 768 21330 800 21362
rect 840 21330 872 21362
rect 912 21330 944 21362
rect 984 21330 1016 21362
rect 1056 21330 1088 21362
rect 1128 21330 1160 21362
rect 1200 21330 1232 21362
rect 1272 21330 1304 21362
rect 1344 21330 1376 21362
rect 1416 21330 1448 21362
rect 1488 21330 1520 21362
rect 1560 21330 1592 21362
rect 1632 21330 1664 21362
rect 1704 21330 1736 21362
rect 1776 21330 1808 21362
rect 1848 21330 1880 21362
rect 120 21258 152 21290
rect 192 21258 224 21290
rect 264 21258 296 21290
rect 336 21258 368 21290
rect 408 21258 440 21290
rect 480 21258 512 21290
rect 552 21258 584 21290
rect 624 21258 656 21290
rect 696 21258 728 21290
rect 768 21258 800 21290
rect 840 21258 872 21290
rect 912 21258 944 21290
rect 984 21258 1016 21290
rect 1056 21258 1088 21290
rect 1128 21258 1160 21290
rect 1200 21258 1232 21290
rect 1272 21258 1304 21290
rect 1344 21258 1376 21290
rect 1416 21258 1448 21290
rect 1488 21258 1520 21290
rect 1560 21258 1592 21290
rect 1632 21258 1664 21290
rect 1704 21258 1736 21290
rect 1776 21258 1808 21290
rect 1848 21258 1880 21290
rect 120 21186 152 21218
rect 192 21186 224 21218
rect 264 21186 296 21218
rect 336 21186 368 21218
rect 408 21186 440 21218
rect 480 21186 512 21218
rect 552 21186 584 21218
rect 624 21186 656 21218
rect 696 21186 728 21218
rect 768 21186 800 21218
rect 840 21186 872 21218
rect 912 21186 944 21218
rect 984 21186 1016 21218
rect 1056 21186 1088 21218
rect 1128 21186 1160 21218
rect 1200 21186 1232 21218
rect 1272 21186 1304 21218
rect 1344 21186 1376 21218
rect 1416 21186 1448 21218
rect 1488 21186 1520 21218
rect 1560 21186 1592 21218
rect 1632 21186 1664 21218
rect 1704 21186 1736 21218
rect 1776 21186 1808 21218
rect 1848 21186 1880 21218
rect 120 21114 152 21146
rect 192 21114 224 21146
rect 264 21114 296 21146
rect 336 21114 368 21146
rect 408 21114 440 21146
rect 480 21114 512 21146
rect 552 21114 584 21146
rect 624 21114 656 21146
rect 696 21114 728 21146
rect 768 21114 800 21146
rect 840 21114 872 21146
rect 912 21114 944 21146
rect 984 21114 1016 21146
rect 1056 21114 1088 21146
rect 1128 21114 1160 21146
rect 1200 21114 1232 21146
rect 1272 21114 1304 21146
rect 1344 21114 1376 21146
rect 1416 21114 1448 21146
rect 1488 21114 1520 21146
rect 1560 21114 1592 21146
rect 1632 21114 1664 21146
rect 1704 21114 1736 21146
rect 1776 21114 1808 21146
rect 1848 21114 1880 21146
rect 120 21042 152 21074
rect 192 21042 224 21074
rect 264 21042 296 21074
rect 336 21042 368 21074
rect 408 21042 440 21074
rect 480 21042 512 21074
rect 552 21042 584 21074
rect 624 21042 656 21074
rect 696 21042 728 21074
rect 768 21042 800 21074
rect 840 21042 872 21074
rect 912 21042 944 21074
rect 984 21042 1016 21074
rect 1056 21042 1088 21074
rect 1128 21042 1160 21074
rect 1200 21042 1232 21074
rect 1272 21042 1304 21074
rect 1344 21042 1376 21074
rect 1416 21042 1448 21074
rect 1488 21042 1520 21074
rect 1560 21042 1592 21074
rect 1632 21042 1664 21074
rect 1704 21042 1736 21074
rect 1776 21042 1808 21074
rect 1848 21042 1880 21074
rect 120 20970 152 21002
rect 192 20970 224 21002
rect 264 20970 296 21002
rect 336 20970 368 21002
rect 408 20970 440 21002
rect 480 20970 512 21002
rect 552 20970 584 21002
rect 624 20970 656 21002
rect 696 20970 728 21002
rect 768 20970 800 21002
rect 840 20970 872 21002
rect 912 20970 944 21002
rect 984 20970 1016 21002
rect 1056 20970 1088 21002
rect 1128 20970 1160 21002
rect 1200 20970 1232 21002
rect 1272 20970 1304 21002
rect 1344 20970 1376 21002
rect 1416 20970 1448 21002
rect 1488 20970 1520 21002
rect 1560 20970 1592 21002
rect 1632 20970 1664 21002
rect 1704 20970 1736 21002
rect 1776 20970 1808 21002
rect 1848 20970 1880 21002
rect 120 20898 152 20930
rect 192 20898 224 20930
rect 264 20898 296 20930
rect 336 20898 368 20930
rect 408 20898 440 20930
rect 480 20898 512 20930
rect 552 20898 584 20930
rect 624 20898 656 20930
rect 696 20898 728 20930
rect 768 20898 800 20930
rect 840 20898 872 20930
rect 912 20898 944 20930
rect 984 20898 1016 20930
rect 1056 20898 1088 20930
rect 1128 20898 1160 20930
rect 1200 20898 1232 20930
rect 1272 20898 1304 20930
rect 1344 20898 1376 20930
rect 1416 20898 1448 20930
rect 1488 20898 1520 20930
rect 1560 20898 1592 20930
rect 1632 20898 1664 20930
rect 1704 20898 1736 20930
rect 1776 20898 1808 20930
rect 1848 20898 1880 20930
rect 120 20826 152 20858
rect 192 20826 224 20858
rect 264 20826 296 20858
rect 336 20826 368 20858
rect 408 20826 440 20858
rect 480 20826 512 20858
rect 552 20826 584 20858
rect 624 20826 656 20858
rect 696 20826 728 20858
rect 768 20826 800 20858
rect 840 20826 872 20858
rect 912 20826 944 20858
rect 984 20826 1016 20858
rect 1056 20826 1088 20858
rect 1128 20826 1160 20858
rect 1200 20826 1232 20858
rect 1272 20826 1304 20858
rect 1344 20826 1376 20858
rect 1416 20826 1448 20858
rect 1488 20826 1520 20858
rect 1560 20826 1592 20858
rect 1632 20826 1664 20858
rect 1704 20826 1736 20858
rect 1776 20826 1808 20858
rect 1848 20826 1880 20858
rect 120 20754 152 20786
rect 192 20754 224 20786
rect 264 20754 296 20786
rect 336 20754 368 20786
rect 408 20754 440 20786
rect 480 20754 512 20786
rect 552 20754 584 20786
rect 624 20754 656 20786
rect 696 20754 728 20786
rect 768 20754 800 20786
rect 840 20754 872 20786
rect 912 20754 944 20786
rect 984 20754 1016 20786
rect 1056 20754 1088 20786
rect 1128 20754 1160 20786
rect 1200 20754 1232 20786
rect 1272 20754 1304 20786
rect 1344 20754 1376 20786
rect 1416 20754 1448 20786
rect 1488 20754 1520 20786
rect 1560 20754 1592 20786
rect 1632 20754 1664 20786
rect 1704 20754 1736 20786
rect 1776 20754 1808 20786
rect 1848 20754 1880 20786
rect 120 20682 152 20714
rect 192 20682 224 20714
rect 264 20682 296 20714
rect 336 20682 368 20714
rect 408 20682 440 20714
rect 480 20682 512 20714
rect 552 20682 584 20714
rect 624 20682 656 20714
rect 696 20682 728 20714
rect 768 20682 800 20714
rect 840 20682 872 20714
rect 912 20682 944 20714
rect 984 20682 1016 20714
rect 1056 20682 1088 20714
rect 1128 20682 1160 20714
rect 1200 20682 1232 20714
rect 1272 20682 1304 20714
rect 1344 20682 1376 20714
rect 1416 20682 1448 20714
rect 1488 20682 1520 20714
rect 1560 20682 1592 20714
rect 1632 20682 1664 20714
rect 1704 20682 1736 20714
rect 1776 20682 1808 20714
rect 1848 20682 1880 20714
rect 120 20610 152 20642
rect 192 20610 224 20642
rect 264 20610 296 20642
rect 336 20610 368 20642
rect 408 20610 440 20642
rect 480 20610 512 20642
rect 552 20610 584 20642
rect 624 20610 656 20642
rect 696 20610 728 20642
rect 768 20610 800 20642
rect 840 20610 872 20642
rect 912 20610 944 20642
rect 984 20610 1016 20642
rect 1056 20610 1088 20642
rect 1128 20610 1160 20642
rect 1200 20610 1232 20642
rect 1272 20610 1304 20642
rect 1344 20610 1376 20642
rect 1416 20610 1448 20642
rect 1488 20610 1520 20642
rect 1560 20610 1592 20642
rect 1632 20610 1664 20642
rect 1704 20610 1736 20642
rect 1776 20610 1808 20642
rect 1848 20610 1880 20642
rect 120 20538 152 20570
rect 192 20538 224 20570
rect 264 20538 296 20570
rect 336 20538 368 20570
rect 408 20538 440 20570
rect 480 20538 512 20570
rect 552 20538 584 20570
rect 624 20538 656 20570
rect 696 20538 728 20570
rect 768 20538 800 20570
rect 840 20538 872 20570
rect 912 20538 944 20570
rect 984 20538 1016 20570
rect 1056 20538 1088 20570
rect 1128 20538 1160 20570
rect 1200 20538 1232 20570
rect 1272 20538 1304 20570
rect 1344 20538 1376 20570
rect 1416 20538 1448 20570
rect 1488 20538 1520 20570
rect 1560 20538 1592 20570
rect 1632 20538 1664 20570
rect 1704 20538 1736 20570
rect 1776 20538 1808 20570
rect 1848 20538 1880 20570
rect 120 20466 152 20498
rect 192 20466 224 20498
rect 264 20466 296 20498
rect 336 20466 368 20498
rect 408 20466 440 20498
rect 480 20466 512 20498
rect 552 20466 584 20498
rect 624 20466 656 20498
rect 696 20466 728 20498
rect 768 20466 800 20498
rect 840 20466 872 20498
rect 912 20466 944 20498
rect 984 20466 1016 20498
rect 1056 20466 1088 20498
rect 1128 20466 1160 20498
rect 1200 20466 1232 20498
rect 1272 20466 1304 20498
rect 1344 20466 1376 20498
rect 1416 20466 1448 20498
rect 1488 20466 1520 20498
rect 1560 20466 1592 20498
rect 1632 20466 1664 20498
rect 1704 20466 1736 20498
rect 1776 20466 1808 20498
rect 1848 20466 1880 20498
rect 120 20394 152 20426
rect 192 20394 224 20426
rect 264 20394 296 20426
rect 336 20394 368 20426
rect 408 20394 440 20426
rect 480 20394 512 20426
rect 552 20394 584 20426
rect 624 20394 656 20426
rect 696 20394 728 20426
rect 768 20394 800 20426
rect 840 20394 872 20426
rect 912 20394 944 20426
rect 984 20394 1016 20426
rect 1056 20394 1088 20426
rect 1128 20394 1160 20426
rect 1200 20394 1232 20426
rect 1272 20394 1304 20426
rect 1344 20394 1376 20426
rect 1416 20394 1448 20426
rect 1488 20394 1520 20426
rect 1560 20394 1592 20426
rect 1632 20394 1664 20426
rect 1704 20394 1736 20426
rect 1776 20394 1808 20426
rect 1848 20394 1880 20426
rect 120 20322 152 20354
rect 192 20322 224 20354
rect 264 20322 296 20354
rect 336 20322 368 20354
rect 408 20322 440 20354
rect 480 20322 512 20354
rect 552 20322 584 20354
rect 624 20322 656 20354
rect 696 20322 728 20354
rect 768 20322 800 20354
rect 840 20322 872 20354
rect 912 20322 944 20354
rect 984 20322 1016 20354
rect 1056 20322 1088 20354
rect 1128 20322 1160 20354
rect 1200 20322 1232 20354
rect 1272 20322 1304 20354
rect 1344 20322 1376 20354
rect 1416 20322 1448 20354
rect 1488 20322 1520 20354
rect 1560 20322 1592 20354
rect 1632 20322 1664 20354
rect 1704 20322 1736 20354
rect 1776 20322 1808 20354
rect 1848 20322 1880 20354
rect 120 20250 152 20282
rect 192 20250 224 20282
rect 264 20250 296 20282
rect 336 20250 368 20282
rect 408 20250 440 20282
rect 480 20250 512 20282
rect 552 20250 584 20282
rect 624 20250 656 20282
rect 696 20250 728 20282
rect 768 20250 800 20282
rect 840 20250 872 20282
rect 912 20250 944 20282
rect 984 20250 1016 20282
rect 1056 20250 1088 20282
rect 1128 20250 1160 20282
rect 1200 20250 1232 20282
rect 1272 20250 1304 20282
rect 1344 20250 1376 20282
rect 1416 20250 1448 20282
rect 1488 20250 1520 20282
rect 1560 20250 1592 20282
rect 1632 20250 1664 20282
rect 1704 20250 1736 20282
rect 1776 20250 1808 20282
rect 1848 20250 1880 20282
rect 120 20178 152 20210
rect 192 20178 224 20210
rect 264 20178 296 20210
rect 336 20178 368 20210
rect 408 20178 440 20210
rect 480 20178 512 20210
rect 552 20178 584 20210
rect 624 20178 656 20210
rect 696 20178 728 20210
rect 768 20178 800 20210
rect 840 20178 872 20210
rect 912 20178 944 20210
rect 984 20178 1016 20210
rect 1056 20178 1088 20210
rect 1128 20178 1160 20210
rect 1200 20178 1232 20210
rect 1272 20178 1304 20210
rect 1344 20178 1376 20210
rect 1416 20178 1448 20210
rect 1488 20178 1520 20210
rect 1560 20178 1592 20210
rect 1632 20178 1664 20210
rect 1704 20178 1736 20210
rect 1776 20178 1808 20210
rect 1848 20178 1880 20210
rect 120 20106 152 20138
rect 192 20106 224 20138
rect 264 20106 296 20138
rect 336 20106 368 20138
rect 408 20106 440 20138
rect 480 20106 512 20138
rect 552 20106 584 20138
rect 624 20106 656 20138
rect 696 20106 728 20138
rect 768 20106 800 20138
rect 840 20106 872 20138
rect 912 20106 944 20138
rect 984 20106 1016 20138
rect 1056 20106 1088 20138
rect 1128 20106 1160 20138
rect 1200 20106 1232 20138
rect 1272 20106 1304 20138
rect 1344 20106 1376 20138
rect 1416 20106 1448 20138
rect 1488 20106 1520 20138
rect 1560 20106 1592 20138
rect 1632 20106 1664 20138
rect 1704 20106 1736 20138
rect 1776 20106 1808 20138
rect 1848 20106 1880 20138
rect 120 20034 152 20066
rect 192 20034 224 20066
rect 264 20034 296 20066
rect 336 20034 368 20066
rect 408 20034 440 20066
rect 480 20034 512 20066
rect 552 20034 584 20066
rect 624 20034 656 20066
rect 696 20034 728 20066
rect 768 20034 800 20066
rect 840 20034 872 20066
rect 912 20034 944 20066
rect 984 20034 1016 20066
rect 1056 20034 1088 20066
rect 1128 20034 1160 20066
rect 1200 20034 1232 20066
rect 1272 20034 1304 20066
rect 1344 20034 1376 20066
rect 1416 20034 1448 20066
rect 1488 20034 1520 20066
rect 1560 20034 1592 20066
rect 1632 20034 1664 20066
rect 1704 20034 1736 20066
rect 1776 20034 1808 20066
rect 1848 20034 1880 20066
rect 120 19962 152 19994
rect 192 19962 224 19994
rect 264 19962 296 19994
rect 336 19962 368 19994
rect 408 19962 440 19994
rect 480 19962 512 19994
rect 552 19962 584 19994
rect 624 19962 656 19994
rect 696 19962 728 19994
rect 768 19962 800 19994
rect 840 19962 872 19994
rect 912 19962 944 19994
rect 984 19962 1016 19994
rect 1056 19962 1088 19994
rect 1128 19962 1160 19994
rect 1200 19962 1232 19994
rect 1272 19962 1304 19994
rect 1344 19962 1376 19994
rect 1416 19962 1448 19994
rect 1488 19962 1520 19994
rect 1560 19962 1592 19994
rect 1632 19962 1664 19994
rect 1704 19962 1736 19994
rect 1776 19962 1808 19994
rect 1848 19962 1880 19994
rect 120 19890 152 19922
rect 192 19890 224 19922
rect 264 19890 296 19922
rect 336 19890 368 19922
rect 408 19890 440 19922
rect 480 19890 512 19922
rect 552 19890 584 19922
rect 624 19890 656 19922
rect 696 19890 728 19922
rect 768 19890 800 19922
rect 840 19890 872 19922
rect 912 19890 944 19922
rect 984 19890 1016 19922
rect 1056 19890 1088 19922
rect 1128 19890 1160 19922
rect 1200 19890 1232 19922
rect 1272 19890 1304 19922
rect 1344 19890 1376 19922
rect 1416 19890 1448 19922
rect 1488 19890 1520 19922
rect 1560 19890 1592 19922
rect 1632 19890 1664 19922
rect 1704 19890 1736 19922
rect 1776 19890 1808 19922
rect 1848 19890 1880 19922
rect 120 19818 152 19850
rect 192 19818 224 19850
rect 264 19818 296 19850
rect 336 19818 368 19850
rect 408 19818 440 19850
rect 480 19818 512 19850
rect 552 19818 584 19850
rect 624 19818 656 19850
rect 696 19818 728 19850
rect 768 19818 800 19850
rect 840 19818 872 19850
rect 912 19818 944 19850
rect 984 19818 1016 19850
rect 1056 19818 1088 19850
rect 1128 19818 1160 19850
rect 1200 19818 1232 19850
rect 1272 19818 1304 19850
rect 1344 19818 1376 19850
rect 1416 19818 1448 19850
rect 1488 19818 1520 19850
rect 1560 19818 1592 19850
rect 1632 19818 1664 19850
rect 1704 19818 1736 19850
rect 1776 19818 1808 19850
rect 1848 19818 1880 19850
rect 120 19746 152 19778
rect 192 19746 224 19778
rect 264 19746 296 19778
rect 336 19746 368 19778
rect 408 19746 440 19778
rect 480 19746 512 19778
rect 552 19746 584 19778
rect 624 19746 656 19778
rect 696 19746 728 19778
rect 768 19746 800 19778
rect 840 19746 872 19778
rect 912 19746 944 19778
rect 984 19746 1016 19778
rect 1056 19746 1088 19778
rect 1128 19746 1160 19778
rect 1200 19746 1232 19778
rect 1272 19746 1304 19778
rect 1344 19746 1376 19778
rect 1416 19746 1448 19778
rect 1488 19746 1520 19778
rect 1560 19746 1592 19778
rect 1632 19746 1664 19778
rect 1704 19746 1736 19778
rect 1776 19746 1808 19778
rect 1848 19746 1880 19778
rect 120 19674 152 19706
rect 192 19674 224 19706
rect 264 19674 296 19706
rect 336 19674 368 19706
rect 408 19674 440 19706
rect 480 19674 512 19706
rect 552 19674 584 19706
rect 624 19674 656 19706
rect 696 19674 728 19706
rect 768 19674 800 19706
rect 840 19674 872 19706
rect 912 19674 944 19706
rect 984 19674 1016 19706
rect 1056 19674 1088 19706
rect 1128 19674 1160 19706
rect 1200 19674 1232 19706
rect 1272 19674 1304 19706
rect 1344 19674 1376 19706
rect 1416 19674 1448 19706
rect 1488 19674 1520 19706
rect 1560 19674 1592 19706
rect 1632 19674 1664 19706
rect 1704 19674 1736 19706
rect 1776 19674 1808 19706
rect 1848 19674 1880 19706
rect 120 19602 152 19634
rect 192 19602 224 19634
rect 264 19602 296 19634
rect 336 19602 368 19634
rect 408 19602 440 19634
rect 480 19602 512 19634
rect 552 19602 584 19634
rect 624 19602 656 19634
rect 696 19602 728 19634
rect 768 19602 800 19634
rect 840 19602 872 19634
rect 912 19602 944 19634
rect 984 19602 1016 19634
rect 1056 19602 1088 19634
rect 1128 19602 1160 19634
rect 1200 19602 1232 19634
rect 1272 19602 1304 19634
rect 1344 19602 1376 19634
rect 1416 19602 1448 19634
rect 1488 19602 1520 19634
rect 1560 19602 1592 19634
rect 1632 19602 1664 19634
rect 1704 19602 1736 19634
rect 1776 19602 1808 19634
rect 1848 19602 1880 19634
rect 120 19530 152 19562
rect 192 19530 224 19562
rect 264 19530 296 19562
rect 336 19530 368 19562
rect 408 19530 440 19562
rect 480 19530 512 19562
rect 552 19530 584 19562
rect 624 19530 656 19562
rect 696 19530 728 19562
rect 768 19530 800 19562
rect 840 19530 872 19562
rect 912 19530 944 19562
rect 984 19530 1016 19562
rect 1056 19530 1088 19562
rect 1128 19530 1160 19562
rect 1200 19530 1232 19562
rect 1272 19530 1304 19562
rect 1344 19530 1376 19562
rect 1416 19530 1448 19562
rect 1488 19530 1520 19562
rect 1560 19530 1592 19562
rect 1632 19530 1664 19562
rect 1704 19530 1736 19562
rect 1776 19530 1808 19562
rect 1848 19530 1880 19562
rect 120 19458 152 19490
rect 192 19458 224 19490
rect 264 19458 296 19490
rect 336 19458 368 19490
rect 408 19458 440 19490
rect 480 19458 512 19490
rect 552 19458 584 19490
rect 624 19458 656 19490
rect 696 19458 728 19490
rect 768 19458 800 19490
rect 840 19458 872 19490
rect 912 19458 944 19490
rect 984 19458 1016 19490
rect 1056 19458 1088 19490
rect 1128 19458 1160 19490
rect 1200 19458 1232 19490
rect 1272 19458 1304 19490
rect 1344 19458 1376 19490
rect 1416 19458 1448 19490
rect 1488 19458 1520 19490
rect 1560 19458 1592 19490
rect 1632 19458 1664 19490
rect 1704 19458 1736 19490
rect 1776 19458 1808 19490
rect 1848 19458 1880 19490
rect 120 19386 152 19418
rect 192 19386 224 19418
rect 264 19386 296 19418
rect 336 19386 368 19418
rect 408 19386 440 19418
rect 480 19386 512 19418
rect 552 19386 584 19418
rect 624 19386 656 19418
rect 696 19386 728 19418
rect 768 19386 800 19418
rect 840 19386 872 19418
rect 912 19386 944 19418
rect 984 19386 1016 19418
rect 1056 19386 1088 19418
rect 1128 19386 1160 19418
rect 1200 19386 1232 19418
rect 1272 19386 1304 19418
rect 1344 19386 1376 19418
rect 1416 19386 1448 19418
rect 1488 19386 1520 19418
rect 1560 19386 1592 19418
rect 1632 19386 1664 19418
rect 1704 19386 1736 19418
rect 1776 19386 1808 19418
rect 1848 19386 1880 19418
rect 120 19314 152 19346
rect 192 19314 224 19346
rect 264 19314 296 19346
rect 336 19314 368 19346
rect 408 19314 440 19346
rect 480 19314 512 19346
rect 552 19314 584 19346
rect 624 19314 656 19346
rect 696 19314 728 19346
rect 768 19314 800 19346
rect 840 19314 872 19346
rect 912 19314 944 19346
rect 984 19314 1016 19346
rect 1056 19314 1088 19346
rect 1128 19314 1160 19346
rect 1200 19314 1232 19346
rect 1272 19314 1304 19346
rect 1344 19314 1376 19346
rect 1416 19314 1448 19346
rect 1488 19314 1520 19346
rect 1560 19314 1592 19346
rect 1632 19314 1664 19346
rect 1704 19314 1736 19346
rect 1776 19314 1808 19346
rect 1848 19314 1880 19346
rect 120 19242 152 19274
rect 192 19242 224 19274
rect 264 19242 296 19274
rect 336 19242 368 19274
rect 408 19242 440 19274
rect 480 19242 512 19274
rect 552 19242 584 19274
rect 624 19242 656 19274
rect 696 19242 728 19274
rect 768 19242 800 19274
rect 840 19242 872 19274
rect 912 19242 944 19274
rect 984 19242 1016 19274
rect 1056 19242 1088 19274
rect 1128 19242 1160 19274
rect 1200 19242 1232 19274
rect 1272 19242 1304 19274
rect 1344 19242 1376 19274
rect 1416 19242 1448 19274
rect 1488 19242 1520 19274
rect 1560 19242 1592 19274
rect 1632 19242 1664 19274
rect 1704 19242 1736 19274
rect 1776 19242 1808 19274
rect 1848 19242 1880 19274
rect 120 19170 152 19202
rect 192 19170 224 19202
rect 264 19170 296 19202
rect 336 19170 368 19202
rect 408 19170 440 19202
rect 480 19170 512 19202
rect 552 19170 584 19202
rect 624 19170 656 19202
rect 696 19170 728 19202
rect 768 19170 800 19202
rect 840 19170 872 19202
rect 912 19170 944 19202
rect 984 19170 1016 19202
rect 1056 19170 1088 19202
rect 1128 19170 1160 19202
rect 1200 19170 1232 19202
rect 1272 19170 1304 19202
rect 1344 19170 1376 19202
rect 1416 19170 1448 19202
rect 1488 19170 1520 19202
rect 1560 19170 1592 19202
rect 1632 19170 1664 19202
rect 1704 19170 1736 19202
rect 1776 19170 1808 19202
rect 1848 19170 1880 19202
rect 120 19098 152 19130
rect 192 19098 224 19130
rect 264 19098 296 19130
rect 336 19098 368 19130
rect 408 19098 440 19130
rect 480 19098 512 19130
rect 552 19098 584 19130
rect 624 19098 656 19130
rect 696 19098 728 19130
rect 768 19098 800 19130
rect 840 19098 872 19130
rect 912 19098 944 19130
rect 984 19098 1016 19130
rect 1056 19098 1088 19130
rect 1128 19098 1160 19130
rect 1200 19098 1232 19130
rect 1272 19098 1304 19130
rect 1344 19098 1376 19130
rect 1416 19098 1448 19130
rect 1488 19098 1520 19130
rect 1560 19098 1592 19130
rect 1632 19098 1664 19130
rect 1704 19098 1736 19130
rect 1776 19098 1808 19130
rect 1848 19098 1880 19130
rect 120 19026 152 19058
rect 192 19026 224 19058
rect 264 19026 296 19058
rect 336 19026 368 19058
rect 408 19026 440 19058
rect 480 19026 512 19058
rect 552 19026 584 19058
rect 624 19026 656 19058
rect 696 19026 728 19058
rect 768 19026 800 19058
rect 840 19026 872 19058
rect 912 19026 944 19058
rect 984 19026 1016 19058
rect 1056 19026 1088 19058
rect 1128 19026 1160 19058
rect 1200 19026 1232 19058
rect 1272 19026 1304 19058
rect 1344 19026 1376 19058
rect 1416 19026 1448 19058
rect 1488 19026 1520 19058
rect 1560 19026 1592 19058
rect 1632 19026 1664 19058
rect 1704 19026 1736 19058
rect 1776 19026 1808 19058
rect 1848 19026 1880 19058
rect 120 18954 152 18986
rect 192 18954 224 18986
rect 264 18954 296 18986
rect 336 18954 368 18986
rect 408 18954 440 18986
rect 480 18954 512 18986
rect 552 18954 584 18986
rect 624 18954 656 18986
rect 696 18954 728 18986
rect 768 18954 800 18986
rect 840 18954 872 18986
rect 912 18954 944 18986
rect 984 18954 1016 18986
rect 1056 18954 1088 18986
rect 1128 18954 1160 18986
rect 1200 18954 1232 18986
rect 1272 18954 1304 18986
rect 1344 18954 1376 18986
rect 1416 18954 1448 18986
rect 1488 18954 1520 18986
rect 1560 18954 1592 18986
rect 1632 18954 1664 18986
rect 1704 18954 1736 18986
rect 1776 18954 1808 18986
rect 1848 18954 1880 18986
rect 120 18882 152 18914
rect 192 18882 224 18914
rect 264 18882 296 18914
rect 336 18882 368 18914
rect 408 18882 440 18914
rect 480 18882 512 18914
rect 552 18882 584 18914
rect 624 18882 656 18914
rect 696 18882 728 18914
rect 768 18882 800 18914
rect 840 18882 872 18914
rect 912 18882 944 18914
rect 984 18882 1016 18914
rect 1056 18882 1088 18914
rect 1128 18882 1160 18914
rect 1200 18882 1232 18914
rect 1272 18882 1304 18914
rect 1344 18882 1376 18914
rect 1416 18882 1448 18914
rect 1488 18882 1520 18914
rect 1560 18882 1592 18914
rect 1632 18882 1664 18914
rect 1704 18882 1736 18914
rect 1776 18882 1808 18914
rect 1848 18882 1880 18914
rect 120 18810 152 18842
rect 192 18810 224 18842
rect 264 18810 296 18842
rect 336 18810 368 18842
rect 408 18810 440 18842
rect 480 18810 512 18842
rect 552 18810 584 18842
rect 624 18810 656 18842
rect 696 18810 728 18842
rect 768 18810 800 18842
rect 840 18810 872 18842
rect 912 18810 944 18842
rect 984 18810 1016 18842
rect 1056 18810 1088 18842
rect 1128 18810 1160 18842
rect 1200 18810 1232 18842
rect 1272 18810 1304 18842
rect 1344 18810 1376 18842
rect 1416 18810 1448 18842
rect 1488 18810 1520 18842
rect 1560 18810 1592 18842
rect 1632 18810 1664 18842
rect 1704 18810 1736 18842
rect 1776 18810 1808 18842
rect 1848 18810 1880 18842
rect 120 18738 152 18770
rect 192 18738 224 18770
rect 264 18738 296 18770
rect 336 18738 368 18770
rect 408 18738 440 18770
rect 480 18738 512 18770
rect 552 18738 584 18770
rect 624 18738 656 18770
rect 696 18738 728 18770
rect 768 18738 800 18770
rect 840 18738 872 18770
rect 912 18738 944 18770
rect 984 18738 1016 18770
rect 1056 18738 1088 18770
rect 1128 18738 1160 18770
rect 1200 18738 1232 18770
rect 1272 18738 1304 18770
rect 1344 18738 1376 18770
rect 1416 18738 1448 18770
rect 1488 18738 1520 18770
rect 1560 18738 1592 18770
rect 1632 18738 1664 18770
rect 1704 18738 1736 18770
rect 1776 18738 1808 18770
rect 1848 18738 1880 18770
rect 120 18666 152 18698
rect 192 18666 224 18698
rect 264 18666 296 18698
rect 336 18666 368 18698
rect 408 18666 440 18698
rect 480 18666 512 18698
rect 552 18666 584 18698
rect 624 18666 656 18698
rect 696 18666 728 18698
rect 768 18666 800 18698
rect 840 18666 872 18698
rect 912 18666 944 18698
rect 984 18666 1016 18698
rect 1056 18666 1088 18698
rect 1128 18666 1160 18698
rect 1200 18666 1232 18698
rect 1272 18666 1304 18698
rect 1344 18666 1376 18698
rect 1416 18666 1448 18698
rect 1488 18666 1520 18698
rect 1560 18666 1592 18698
rect 1632 18666 1664 18698
rect 1704 18666 1736 18698
rect 1776 18666 1808 18698
rect 1848 18666 1880 18698
rect 120 18594 152 18626
rect 192 18594 224 18626
rect 264 18594 296 18626
rect 336 18594 368 18626
rect 408 18594 440 18626
rect 480 18594 512 18626
rect 552 18594 584 18626
rect 624 18594 656 18626
rect 696 18594 728 18626
rect 768 18594 800 18626
rect 840 18594 872 18626
rect 912 18594 944 18626
rect 984 18594 1016 18626
rect 1056 18594 1088 18626
rect 1128 18594 1160 18626
rect 1200 18594 1232 18626
rect 1272 18594 1304 18626
rect 1344 18594 1376 18626
rect 1416 18594 1448 18626
rect 1488 18594 1520 18626
rect 1560 18594 1592 18626
rect 1632 18594 1664 18626
rect 1704 18594 1736 18626
rect 1776 18594 1808 18626
rect 1848 18594 1880 18626
rect 120 18522 152 18554
rect 192 18522 224 18554
rect 264 18522 296 18554
rect 336 18522 368 18554
rect 408 18522 440 18554
rect 480 18522 512 18554
rect 552 18522 584 18554
rect 624 18522 656 18554
rect 696 18522 728 18554
rect 768 18522 800 18554
rect 840 18522 872 18554
rect 912 18522 944 18554
rect 984 18522 1016 18554
rect 1056 18522 1088 18554
rect 1128 18522 1160 18554
rect 1200 18522 1232 18554
rect 1272 18522 1304 18554
rect 1344 18522 1376 18554
rect 1416 18522 1448 18554
rect 1488 18522 1520 18554
rect 1560 18522 1592 18554
rect 1632 18522 1664 18554
rect 1704 18522 1736 18554
rect 1776 18522 1808 18554
rect 1848 18522 1880 18554
rect 120 18450 152 18482
rect 192 18450 224 18482
rect 264 18450 296 18482
rect 336 18450 368 18482
rect 408 18450 440 18482
rect 480 18450 512 18482
rect 552 18450 584 18482
rect 624 18450 656 18482
rect 696 18450 728 18482
rect 768 18450 800 18482
rect 840 18450 872 18482
rect 912 18450 944 18482
rect 984 18450 1016 18482
rect 1056 18450 1088 18482
rect 1128 18450 1160 18482
rect 1200 18450 1232 18482
rect 1272 18450 1304 18482
rect 1344 18450 1376 18482
rect 1416 18450 1448 18482
rect 1488 18450 1520 18482
rect 1560 18450 1592 18482
rect 1632 18450 1664 18482
rect 1704 18450 1736 18482
rect 1776 18450 1808 18482
rect 1848 18450 1880 18482
rect 120 18378 152 18410
rect 192 18378 224 18410
rect 264 18378 296 18410
rect 336 18378 368 18410
rect 408 18378 440 18410
rect 480 18378 512 18410
rect 552 18378 584 18410
rect 624 18378 656 18410
rect 696 18378 728 18410
rect 768 18378 800 18410
rect 840 18378 872 18410
rect 912 18378 944 18410
rect 984 18378 1016 18410
rect 1056 18378 1088 18410
rect 1128 18378 1160 18410
rect 1200 18378 1232 18410
rect 1272 18378 1304 18410
rect 1344 18378 1376 18410
rect 1416 18378 1448 18410
rect 1488 18378 1520 18410
rect 1560 18378 1592 18410
rect 1632 18378 1664 18410
rect 1704 18378 1736 18410
rect 1776 18378 1808 18410
rect 1848 18378 1880 18410
rect 120 18306 152 18338
rect 192 18306 224 18338
rect 264 18306 296 18338
rect 336 18306 368 18338
rect 408 18306 440 18338
rect 480 18306 512 18338
rect 552 18306 584 18338
rect 624 18306 656 18338
rect 696 18306 728 18338
rect 768 18306 800 18338
rect 840 18306 872 18338
rect 912 18306 944 18338
rect 984 18306 1016 18338
rect 1056 18306 1088 18338
rect 1128 18306 1160 18338
rect 1200 18306 1232 18338
rect 1272 18306 1304 18338
rect 1344 18306 1376 18338
rect 1416 18306 1448 18338
rect 1488 18306 1520 18338
rect 1560 18306 1592 18338
rect 1632 18306 1664 18338
rect 1704 18306 1736 18338
rect 1776 18306 1808 18338
rect 1848 18306 1880 18338
rect 120 18234 152 18266
rect 192 18234 224 18266
rect 264 18234 296 18266
rect 336 18234 368 18266
rect 408 18234 440 18266
rect 480 18234 512 18266
rect 552 18234 584 18266
rect 624 18234 656 18266
rect 696 18234 728 18266
rect 768 18234 800 18266
rect 840 18234 872 18266
rect 912 18234 944 18266
rect 984 18234 1016 18266
rect 1056 18234 1088 18266
rect 1128 18234 1160 18266
rect 1200 18234 1232 18266
rect 1272 18234 1304 18266
rect 1344 18234 1376 18266
rect 1416 18234 1448 18266
rect 1488 18234 1520 18266
rect 1560 18234 1592 18266
rect 1632 18234 1664 18266
rect 1704 18234 1736 18266
rect 1776 18234 1808 18266
rect 1848 18234 1880 18266
rect 120 18162 152 18194
rect 192 18162 224 18194
rect 264 18162 296 18194
rect 336 18162 368 18194
rect 408 18162 440 18194
rect 480 18162 512 18194
rect 552 18162 584 18194
rect 624 18162 656 18194
rect 696 18162 728 18194
rect 768 18162 800 18194
rect 840 18162 872 18194
rect 912 18162 944 18194
rect 984 18162 1016 18194
rect 1056 18162 1088 18194
rect 1128 18162 1160 18194
rect 1200 18162 1232 18194
rect 1272 18162 1304 18194
rect 1344 18162 1376 18194
rect 1416 18162 1448 18194
rect 1488 18162 1520 18194
rect 1560 18162 1592 18194
rect 1632 18162 1664 18194
rect 1704 18162 1736 18194
rect 1776 18162 1808 18194
rect 1848 18162 1880 18194
rect 192 17816 224 17848
rect 264 17816 296 17848
rect 336 17816 368 17848
rect 408 17816 440 17848
rect 480 17816 512 17848
rect 552 17816 584 17848
rect 624 17816 656 17848
rect 696 17816 728 17848
rect 768 17816 800 17848
rect 840 17816 872 17848
rect 912 17816 944 17848
rect 984 17816 1016 17848
rect 1056 17816 1088 17848
rect 1128 17816 1160 17848
rect 1200 17816 1232 17848
rect 1272 17816 1304 17848
rect 1344 17816 1376 17848
rect 1416 17816 1448 17848
rect 1488 17816 1520 17848
rect 1560 17816 1592 17848
rect 1632 17816 1664 17848
rect 1704 17816 1736 17848
rect 1776 17816 1808 17848
rect 1848 17816 1880 17848
rect 120 17744 152 17776
rect 192 17744 224 17776
rect 264 17744 296 17776
rect 336 17744 368 17776
rect 408 17744 440 17776
rect 480 17744 512 17776
rect 552 17744 584 17776
rect 624 17744 656 17776
rect 696 17744 728 17776
rect 768 17744 800 17776
rect 840 17744 872 17776
rect 912 17744 944 17776
rect 984 17744 1016 17776
rect 1056 17744 1088 17776
rect 1128 17744 1160 17776
rect 1200 17744 1232 17776
rect 1272 17744 1304 17776
rect 1344 17744 1376 17776
rect 1416 17744 1448 17776
rect 1488 17744 1520 17776
rect 1560 17744 1592 17776
rect 1632 17744 1664 17776
rect 1704 17744 1736 17776
rect 1776 17744 1808 17776
rect 1848 17744 1880 17776
rect 120 17672 152 17704
rect 192 17672 224 17704
rect 264 17672 296 17704
rect 336 17672 368 17704
rect 408 17672 440 17704
rect 480 17672 512 17704
rect 552 17672 584 17704
rect 624 17672 656 17704
rect 696 17672 728 17704
rect 768 17672 800 17704
rect 840 17672 872 17704
rect 912 17672 944 17704
rect 984 17672 1016 17704
rect 1056 17672 1088 17704
rect 1128 17672 1160 17704
rect 1200 17672 1232 17704
rect 1272 17672 1304 17704
rect 1344 17672 1376 17704
rect 1416 17672 1448 17704
rect 1488 17672 1520 17704
rect 1560 17672 1592 17704
rect 1632 17672 1664 17704
rect 1704 17672 1736 17704
rect 1776 17672 1808 17704
rect 1848 17672 1880 17704
rect 120 17600 152 17632
rect 192 17600 224 17632
rect 264 17600 296 17632
rect 336 17600 368 17632
rect 408 17600 440 17632
rect 480 17600 512 17632
rect 552 17600 584 17632
rect 624 17600 656 17632
rect 696 17600 728 17632
rect 768 17600 800 17632
rect 840 17600 872 17632
rect 912 17600 944 17632
rect 984 17600 1016 17632
rect 1056 17600 1088 17632
rect 1128 17600 1160 17632
rect 1200 17600 1232 17632
rect 1272 17600 1304 17632
rect 1344 17600 1376 17632
rect 1416 17600 1448 17632
rect 1488 17600 1520 17632
rect 1560 17600 1592 17632
rect 1632 17600 1664 17632
rect 1704 17600 1736 17632
rect 1776 17600 1808 17632
rect 1848 17600 1880 17632
rect 120 17528 152 17560
rect 192 17528 224 17560
rect 264 17528 296 17560
rect 336 17528 368 17560
rect 408 17528 440 17560
rect 480 17528 512 17560
rect 552 17528 584 17560
rect 624 17528 656 17560
rect 696 17528 728 17560
rect 768 17528 800 17560
rect 840 17528 872 17560
rect 912 17528 944 17560
rect 984 17528 1016 17560
rect 1056 17528 1088 17560
rect 1128 17528 1160 17560
rect 1200 17528 1232 17560
rect 1272 17528 1304 17560
rect 1344 17528 1376 17560
rect 1416 17528 1448 17560
rect 1488 17528 1520 17560
rect 1560 17528 1592 17560
rect 1632 17528 1664 17560
rect 1704 17528 1736 17560
rect 1776 17528 1808 17560
rect 1848 17528 1880 17560
rect 120 17456 152 17488
rect 192 17456 224 17488
rect 264 17456 296 17488
rect 336 17456 368 17488
rect 408 17456 440 17488
rect 480 17456 512 17488
rect 552 17456 584 17488
rect 624 17456 656 17488
rect 696 17456 728 17488
rect 768 17456 800 17488
rect 840 17456 872 17488
rect 912 17456 944 17488
rect 984 17456 1016 17488
rect 1056 17456 1088 17488
rect 1128 17456 1160 17488
rect 1200 17456 1232 17488
rect 1272 17456 1304 17488
rect 1344 17456 1376 17488
rect 1416 17456 1448 17488
rect 1488 17456 1520 17488
rect 1560 17456 1592 17488
rect 1632 17456 1664 17488
rect 1704 17456 1736 17488
rect 1776 17456 1808 17488
rect 1848 17456 1880 17488
rect 120 17384 152 17416
rect 192 17384 224 17416
rect 264 17384 296 17416
rect 336 17384 368 17416
rect 408 17384 440 17416
rect 480 17384 512 17416
rect 552 17384 584 17416
rect 624 17384 656 17416
rect 696 17384 728 17416
rect 768 17384 800 17416
rect 840 17384 872 17416
rect 912 17384 944 17416
rect 984 17384 1016 17416
rect 1056 17384 1088 17416
rect 1128 17384 1160 17416
rect 1200 17384 1232 17416
rect 1272 17384 1304 17416
rect 1344 17384 1376 17416
rect 1416 17384 1448 17416
rect 1488 17384 1520 17416
rect 1560 17384 1592 17416
rect 1632 17384 1664 17416
rect 1704 17384 1736 17416
rect 1776 17384 1808 17416
rect 1848 17384 1880 17416
rect 120 17312 152 17344
rect 192 17312 224 17344
rect 264 17312 296 17344
rect 336 17312 368 17344
rect 408 17312 440 17344
rect 480 17312 512 17344
rect 552 17312 584 17344
rect 624 17312 656 17344
rect 696 17312 728 17344
rect 768 17312 800 17344
rect 840 17312 872 17344
rect 912 17312 944 17344
rect 984 17312 1016 17344
rect 1056 17312 1088 17344
rect 1128 17312 1160 17344
rect 1200 17312 1232 17344
rect 1272 17312 1304 17344
rect 1344 17312 1376 17344
rect 1416 17312 1448 17344
rect 1488 17312 1520 17344
rect 1560 17312 1592 17344
rect 1632 17312 1664 17344
rect 1704 17312 1736 17344
rect 1776 17312 1808 17344
rect 1848 17312 1880 17344
rect 120 17240 152 17272
rect 192 17240 224 17272
rect 264 17240 296 17272
rect 336 17240 368 17272
rect 408 17240 440 17272
rect 480 17240 512 17272
rect 552 17240 584 17272
rect 624 17240 656 17272
rect 696 17240 728 17272
rect 768 17240 800 17272
rect 840 17240 872 17272
rect 912 17240 944 17272
rect 984 17240 1016 17272
rect 1056 17240 1088 17272
rect 1128 17240 1160 17272
rect 1200 17240 1232 17272
rect 1272 17240 1304 17272
rect 1344 17240 1376 17272
rect 1416 17240 1448 17272
rect 1488 17240 1520 17272
rect 1560 17240 1592 17272
rect 1632 17240 1664 17272
rect 1704 17240 1736 17272
rect 1776 17240 1808 17272
rect 1848 17240 1880 17272
rect 120 17168 152 17200
rect 192 17168 224 17200
rect 264 17168 296 17200
rect 336 17168 368 17200
rect 408 17168 440 17200
rect 480 17168 512 17200
rect 552 17168 584 17200
rect 624 17168 656 17200
rect 696 17168 728 17200
rect 768 17168 800 17200
rect 840 17168 872 17200
rect 912 17168 944 17200
rect 984 17168 1016 17200
rect 1056 17168 1088 17200
rect 1128 17168 1160 17200
rect 1200 17168 1232 17200
rect 1272 17168 1304 17200
rect 1344 17168 1376 17200
rect 1416 17168 1448 17200
rect 1488 17168 1520 17200
rect 1560 17168 1592 17200
rect 1632 17168 1664 17200
rect 1704 17168 1736 17200
rect 1776 17168 1808 17200
rect 1848 17168 1880 17200
rect 120 17096 152 17128
rect 192 17096 224 17128
rect 264 17096 296 17128
rect 336 17096 368 17128
rect 408 17096 440 17128
rect 480 17096 512 17128
rect 552 17096 584 17128
rect 624 17096 656 17128
rect 696 17096 728 17128
rect 768 17096 800 17128
rect 840 17096 872 17128
rect 912 17096 944 17128
rect 984 17096 1016 17128
rect 1056 17096 1088 17128
rect 1128 17096 1160 17128
rect 1200 17096 1232 17128
rect 1272 17096 1304 17128
rect 1344 17096 1376 17128
rect 1416 17096 1448 17128
rect 1488 17096 1520 17128
rect 1560 17096 1592 17128
rect 1632 17096 1664 17128
rect 1704 17096 1736 17128
rect 1776 17096 1808 17128
rect 1848 17096 1880 17128
rect 120 17024 152 17056
rect 192 17024 224 17056
rect 264 17024 296 17056
rect 336 17024 368 17056
rect 408 17024 440 17056
rect 480 17024 512 17056
rect 552 17024 584 17056
rect 624 17024 656 17056
rect 696 17024 728 17056
rect 768 17024 800 17056
rect 840 17024 872 17056
rect 912 17024 944 17056
rect 984 17024 1016 17056
rect 1056 17024 1088 17056
rect 1128 17024 1160 17056
rect 1200 17024 1232 17056
rect 1272 17024 1304 17056
rect 1344 17024 1376 17056
rect 1416 17024 1448 17056
rect 1488 17024 1520 17056
rect 1560 17024 1592 17056
rect 1632 17024 1664 17056
rect 1704 17024 1736 17056
rect 1776 17024 1808 17056
rect 1848 17024 1880 17056
rect 120 16952 152 16984
rect 192 16952 224 16984
rect 264 16952 296 16984
rect 336 16952 368 16984
rect 408 16952 440 16984
rect 480 16952 512 16984
rect 552 16952 584 16984
rect 624 16952 656 16984
rect 696 16952 728 16984
rect 768 16952 800 16984
rect 840 16952 872 16984
rect 912 16952 944 16984
rect 984 16952 1016 16984
rect 1056 16952 1088 16984
rect 1128 16952 1160 16984
rect 1200 16952 1232 16984
rect 1272 16952 1304 16984
rect 1344 16952 1376 16984
rect 1416 16952 1448 16984
rect 1488 16952 1520 16984
rect 1560 16952 1592 16984
rect 1632 16952 1664 16984
rect 1704 16952 1736 16984
rect 1776 16952 1808 16984
rect 1848 16952 1880 16984
rect 120 16880 152 16912
rect 192 16880 224 16912
rect 264 16880 296 16912
rect 336 16880 368 16912
rect 408 16880 440 16912
rect 480 16880 512 16912
rect 552 16880 584 16912
rect 624 16880 656 16912
rect 696 16880 728 16912
rect 768 16880 800 16912
rect 840 16880 872 16912
rect 912 16880 944 16912
rect 984 16880 1016 16912
rect 1056 16880 1088 16912
rect 1128 16880 1160 16912
rect 1200 16880 1232 16912
rect 1272 16880 1304 16912
rect 1344 16880 1376 16912
rect 1416 16880 1448 16912
rect 1488 16880 1520 16912
rect 1560 16880 1592 16912
rect 1632 16880 1664 16912
rect 1704 16880 1736 16912
rect 1776 16880 1808 16912
rect 1848 16880 1880 16912
rect 120 16808 152 16840
rect 192 16808 224 16840
rect 264 16808 296 16840
rect 336 16808 368 16840
rect 408 16808 440 16840
rect 480 16808 512 16840
rect 552 16808 584 16840
rect 624 16808 656 16840
rect 696 16808 728 16840
rect 768 16808 800 16840
rect 840 16808 872 16840
rect 912 16808 944 16840
rect 984 16808 1016 16840
rect 1056 16808 1088 16840
rect 1128 16808 1160 16840
rect 1200 16808 1232 16840
rect 1272 16808 1304 16840
rect 1344 16808 1376 16840
rect 1416 16808 1448 16840
rect 1488 16808 1520 16840
rect 1560 16808 1592 16840
rect 1632 16808 1664 16840
rect 1704 16808 1736 16840
rect 1776 16808 1808 16840
rect 1848 16808 1880 16840
rect 120 16736 152 16768
rect 192 16736 224 16768
rect 264 16736 296 16768
rect 336 16736 368 16768
rect 408 16736 440 16768
rect 480 16736 512 16768
rect 552 16736 584 16768
rect 624 16736 656 16768
rect 696 16736 728 16768
rect 768 16736 800 16768
rect 840 16736 872 16768
rect 912 16736 944 16768
rect 984 16736 1016 16768
rect 1056 16736 1088 16768
rect 1128 16736 1160 16768
rect 1200 16736 1232 16768
rect 1272 16736 1304 16768
rect 1344 16736 1376 16768
rect 1416 16736 1448 16768
rect 1488 16736 1520 16768
rect 1560 16736 1592 16768
rect 1632 16736 1664 16768
rect 1704 16736 1736 16768
rect 1776 16736 1808 16768
rect 1848 16736 1880 16768
rect 120 16664 152 16696
rect 192 16664 224 16696
rect 264 16664 296 16696
rect 336 16664 368 16696
rect 408 16664 440 16696
rect 480 16664 512 16696
rect 552 16664 584 16696
rect 624 16664 656 16696
rect 696 16664 728 16696
rect 768 16664 800 16696
rect 840 16664 872 16696
rect 912 16664 944 16696
rect 984 16664 1016 16696
rect 1056 16664 1088 16696
rect 1128 16664 1160 16696
rect 1200 16664 1232 16696
rect 1272 16664 1304 16696
rect 1344 16664 1376 16696
rect 1416 16664 1448 16696
rect 1488 16664 1520 16696
rect 1560 16664 1592 16696
rect 1632 16664 1664 16696
rect 1704 16664 1736 16696
rect 1776 16664 1808 16696
rect 1848 16664 1880 16696
rect 120 16592 152 16624
rect 192 16592 224 16624
rect 264 16592 296 16624
rect 336 16592 368 16624
rect 408 16592 440 16624
rect 480 16592 512 16624
rect 552 16592 584 16624
rect 624 16592 656 16624
rect 696 16592 728 16624
rect 768 16592 800 16624
rect 840 16592 872 16624
rect 912 16592 944 16624
rect 984 16592 1016 16624
rect 1056 16592 1088 16624
rect 1128 16592 1160 16624
rect 1200 16592 1232 16624
rect 1272 16592 1304 16624
rect 1344 16592 1376 16624
rect 1416 16592 1448 16624
rect 1488 16592 1520 16624
rect 1560 16592 1592 16624
rect 1632 16592 1664 16624
rect 1704 16592 1736 16624
rect 1776 16592 1808 16624
rect 1848 16592 1880 16624
rect 120 16520 152 16552
rect 192 16520 224 16552
rect 264 16520 296 16552
rect 336 16520 368 16552
rect 408 16520 440 16552
rect 480 16520 512 16552
rect 552 16520 584 16552
rect 624 16520 656 16552
rect 696 16520 728 16552
rect 768 16520 800 16552
rect 840 16520 872 16552
rect 912 16520 944 16552
rect 984 16520 1016 16552
rect 1056 16520 1088 16552
rect 1128 16520 1160 16552
rect 1200 16520 1232 16552
rect 1272 16520 1304 16552
rect 1344 16520 1376 16552
rect 1416 16520 1448 16552
rect 1488 16520 1520 16552
rect 1560 16520 1592 16552
rect 1632 16520 1664 16552
rect 1704 16520 1736 16552
rect 1776 16520 1808 16552
rect 1848 16520 1880 16552
rect 120 16448 152 16480
rect 192 16448 224 16480
rect 264 16448 296 16480
rect 336 16448 368 16480
rect 408 16448 440 16480
rect 480 16448 512 16480
rect 552 16448 584 16480
rect 624 16448 656 16480
rect 696 16448 728 16480
rect 768 16448 800 16480
rect 840 16448 872 16480
rect 912 16448 944 16480
rect 984 16448 1016 16480
rect 1056 16448 1088 16480
rect 1128 16448 1160 16480
rect 1200 16448 1232 16480
rect 1272 16448 1304 16480
rect 1344 16448 1376 16480
rect 1416 16448 1448 16480
rect 1488 16448 1520 16480
rect 1560 16448 1592 16480
rect 1632 16448 1664 16480
rect 1704 16448 1736 16480
rect 1776 16448 1808 16480
rect 1848 16448 1880 16480
rect 120 16376 152 16408
rect 192 16376 224 16408
rect 264 16376 296 16408
rect 336 16376 368 16408
rect 408 16376 440 16408
rect 480 16376 512 16408
rect 552 16376 584 16408
rect 624 16376 656 16408
rect 696 16376 728 16408
rect 768 16376 800 16408
rect 840 16376 872 16408
rect 912 16376 944 16408
rect 984 16376 1016 16408
rect 1056 16376 1088 16408
rect 1128 16376 1160 16408
rect 1200 16376 1232 16408
rect 1272 16376 1304 16408
rect 1344 16376 1376 16408
rect 1416 16376 1448 16408
rect 1488 16376 1520 16408
rect 1560 16376 1592 16408
rect 1632 16376 1664 16408
rect 1704 16376 1736 16408
rect 1776 16376 1808 16408
rect 1848 16376 1880 16408
rect 120 16304 152 16336
rect 192 16304 224 16336
rect 264 16304 296 16336
rect 336 16304 368 16336
rect 408 16304 440 16336
rect 480 16304 512 16336
rect 552 16304 584 16336
rect 624 16304 656 16336
rect 696 16304 728 16336
rect 768 16304 800 16336
rect 840 16304 872 16336
rect 912 16304 944 16336
rect 984 16304 1016 16336
rect 1056 16304 1088 16336
rect 1128 16304 1160 16336
rect 1200 16304 1232 16336
rect 1272 16304 1304 16336
rect 1344 16304 1376 16336
rect 1416 16304 1448 16336
rect 1488 16304 1520 16336
rect 1560 16304 1592 16336
rect 1632 16304 1664 16336
rect 1704 16304 1736 16336
rect 1776 16304 1808 16336
rect 1848 16304 1880 16336
rect 120 16232 152 16264
rect 192 16232 224 16264
rect 264 16232 296 16264
rect 336 16232 368 16264
rect 408 16232 440 16264
rect 480 16232 512 16264
rect 552 16232 584 16264
rect 624 16232 656 16264
rect 696 16232 728 16264
rect 768 16232 800 16264
rect 840 16232 872 16264
rect 912 16232 944 16264
rect 984 16232 1016 16264
rect 1056 16232 1088 16264
rect 1128 16232 1160 16264
rect 1200 16232 1232 16264
rect 1272 16232 1304 16264
rect 1344 16232 1376 16264
rect 1416 16232 1448 16264
rect 1488 16232 1520 16264
rect 1560 16232 1592 16264
rect 1632 16232 1664 16264
rect 1704 16232 1736 16264
rect 1776 16232 1808 16264
rect 1848 16232 1880 16264
rect 120 16160 152 16192
rect 192 16160 224 16192
rect 264 16160 296 16192
rect 336 16160 368 16192
rect 408 16160 440 16192
rect 480 16160 512 16192
rect 552 16160 584 16192
rect 624 16160 656 16192
rect 696 16160 728 16192
rect 768 16160 800 16192
rect 840 16160 872 16192
rect 912 16160 944 16192
rect 984 16160 1016 16192
rect 1056 16160 1088 16192
rect 1128 16160 1160 16192
rect 1200 16160 1232 16192
rect 1272 16160 1304 16192
rect 1344 16160 1376 16192
rect 1416 16160 1448 16192
rect 1488 16160 1520 16192
rect 1560 16160 1592 16192
rect 1632 16160 1664 16192
rect 1704 16160 1736 16192
rect 1776 16160 1808 16192
rect 1848 16160 1880 16192
rect 120 16088 152 16120
rect 192 16088 224 16120
rect 264 16088 296 16120
rect 336 16088 368 16120
rect 408 16088 440 16120
rect 480 16088 512 16120
rect 552 16088 584 16120
rect 624 16088 656 16120
rect 696 16088 728 16120
rect 768 16088 800 16120
rect 840 16088 872 16120
rect 912 16088 944 16120
rect 984 16088 1016 16120
rect 1056 16088 1088 16120
rect 1128 16088 1160 16120
rect 1200 16088 1232 16120
rect 1272 16088 1304 16120
rect 1344 16088 1376 16120
rect 1416 16088 1448 16120
rect 1488 16088 1520 16120
rect 1560 16088 1592 16120
rect 1632 16088 1664 16120
rect 1704 16088 1736 16120
rect 1776 16088 1808 16120
rect 1848 16088 1880 16120
rect 120 16016 152 16048
rect 192 16016 224 16048
rect 264 16016 296 16048
rect 336 16016 368 16048
rect 408 16016 440 16048
rect 480 16016 512 16048
rect 552 16016 584 16048
rect 624 16016 656 16048
rect 696 16016 728 16048
rect 768 16016 800 16048
rect 840 16016 872 16048
rect 912 16016 944 16048
rect 984 16016 1016 16048
rect 1056 16016 1088 16048
rect 1128 16016 1160 16048
rect 1200 16016 1232 16048
rect 1272 16016 1304 16048
rect 1344 16016 1376 16048
rect 1416 16016 1448 16048
rect 1488 16016 1520 16048
rect 1560 16016 1592 16048
rect 1632 16016 1664 16048
rect 1704 16016 1736 16048
rect 1776 16016 1808 16048
rect 1848 16016 1880 16048
rect 120 15944 152 15976
rect 192 15944 224 15976
rect 264 15944 296 15976
rect 336 15944 368 15976
rect 408 15944 440 15976
rect 480 15944 512 15976
rect 552 15944 584 15976
rect 624 15944 656 15976
rect 696 15944 728 15976
rect 768 15944 800 15976
rect 840 15944 872 15976
rect 912 15944 944 15976
rect 984 15944 1016 15976
rect 1056 15944 1088 15976
rect 1128 15944 1160 15976
rect 1200 15944 1232 15976
rect 1272 15944 1304 15976
rect 1344 15944 1376 15976
rect 1416 15944 1448 15976
rect 1488 15944 1520 15976
rect 1560 15944 1592 15976
rect 1632 15944 1664 15976
rect 1704 15944 1736 15976
rect 1776 15944 1808 15976
rect 1848 15944 1880 15976
rect 120 15872 152 15904
rect 192 15872 224 15904
rect 264 15872 296 15904
rect 336 15872 368 15904
rect 408 15872 440 15904
rect 480 15872 512 15904
rect 552 15872 584 15904
rect 624 15872 656 15904
rect 696 15872 728 15904
rect 768 15872 800 15904
rect 840 15872 872 15904
rect 912 15872 944 15904
rect 984 15872 1016 15904
rect 1056 15872 1088 15904
rect 1128 15872 1160 15904
rect 1200 15872 1232 15904
rect 1272 15872 1304 15904
rect 1344 15872 1376 15904
rect 1416 15872 1448 15904
rect 1488 15872 1520 15904
rect 1560 15872 1592 15904
rect 1632 15872 1664 15904
rect 1704 15872 1736 15904
rect 1776 15872 1808 15904
rect 1848 15872 1880 15904
rect 120 15800 152 15832
rect 192 15800 224 15832
rect 264 15800 296 15832
rect 336 15800 368 15832
rect 408 15800 440 15832
rect 480 15800 512 15832
rect 552 15800 584 15832
rect 624 15800 656 15832
rect 696 15800 728 15832
rect 768 15800 800 15832
rect 840 15800 872 15832
rect 912 15800 944 15832
rect 984 15800 1016 15832
rect 1056 15800 1088 15832
rect 1128 15800 1160 15832
rect 1200 15800 1232 15832
rect 1272 15800 1304 15832
rect 1344 15800 1376 15832
rect 1416 15800 1448 15832
rect 1488 15800 1520 15832
rect 1560 15800 1592 15832
rect 1632 15800 1664 15832
rect 1704 15800 1736 15832
rect 1776 15800 1808 15832
rect 1848 15800 1880 15832
rect 120 15728 152 15760
rect 192 15728 224 15760
rect 264 15728 296 15760
rect 336 15728 368 15760
rect 408 15728 440 15760
rect 480 15728 512 15760
rect 552 15728 584 15760
rect 624 15728 656 15760
rect 696 15728 728 15760
rect 768 15728 800 15760
rect 840 15728 872 15760
rect 912 15728 944 15760
rect 984 15728 1016 15760
rect 1056 15728 1088 15760
rect 1128 15728 1160 15760
rect 1200 15728 1232 15760
rect 1272 15728 1304 15760
rect 1344 15728 1376 15760
rect 1416 15728 1448 15760
rect 1488 15728 1520 15760
rect 1560 15728 1592 15760
rect 1632 15728 1664 15760
rect 1704 15728 1736 15760
rect 1776 15728 1808 15760
rect 1848 15728 1880 15760
rect 120 15656 152 15688
rect 192 15656 224 15688
rect 264 15656 296 15688
rect 336 15656 368 15688
rect 408 15656 440 15688
rect 480 15656 512 15688
rect 552 15656 584 15688
rect 624 15656 656 15688
rect 696 15656 728 15688
rect 768 15656 800 15688
rect 840 15656 872 15688
rect 912 15656 944 15688
rect 984 15656 1016 15688
rect 1056 15656 1088 15688
rect 1128 15656 1160 15688
rect 1200 15656 1232 15688
rect 1272 15656 1304 15688
rect 1344 15656 1376 15688
rect 1416 15656 1448 15688
rect 1488 15656 1520 15688
rect 1560 15656 1592 15688
rect 1632 15656 1664 15688
rect 1704 15656 1736 15688
rect 1776 15656 1808 15688
rect 1848 15656 1880 15688
rect 120 15584 152 15616
rect 192 15584 224 15616
rect 264 15584 296 15616
rect 336 15584 368 15616
rect 408 15584 440 15616
rect 480 15584 512 15616
rect 552 15584 584 15616
rect 624 15584 656 15616
rect 696 15584 728 15616
rect 768 15584 800 15616
rect 840 15584 872 15616
rect 912 15584 944 15616
rect 984 15584 1016 15616
rect 1056 15584 1088 15616
rect 1128 15584 1160 15616
rect 1200 15584 1232 15616
rect 1272 15584 1304 15616
rect 1344 15584 1376 15616
rect 1416 15584 1448 15616
rect 1488 15584 1520 15616
rect 1560 15584 1592 15616
rect 1632 15584 1664 15616
rect 1704 15584 1736 15616
rect 1776 15584 1808 15616
rect 1848 15584 1880 15616
rect 120 15512 152 15544
rect 192 15512 224 15544
rect 264 15512 296 15544
rect 336 15512 368 15544
rect 408 15512 440 15544
rect 480 15512 512 15544
rect 552 15512 584 15544
rect 624 15512 656 15544
rect 696 15512 728 15544
rect 768 15512 800 15544
rect 840 15512 872 15544
rect 912 15512 944 15544
rect 984 15512 1016 15544
rect 1056 15512 1088 15544
rect 1128 15512 1160 15544
rect 1200 15512 1232 15544
rect 1272 15512 1304 15544
rect 1344 15512 1376 15544
rect 1416 15512 1448 15544
rect 1488 15512 1520 15544
rect 1560 15512 1592 15544
rect 1632 15512 1664 15544
rect 1704 15512 1736 15544
rect 1776 15512 1808 15544
rect 1848 15512 1880 15544
rect 120 15440 152 15472
rect 192 15440 224 15472
rect 264 15440 296 15472
rect 336 15440 368 15472
rect 408 15440 440 15472
rect 480 15440 512 15472
rect 552 15440 584 15472
rect 624 15440 656 15472
rect 696 15440 728 15472
rect 768 15440 800 15472
rect 840 15440 872 15472
rect 912 15440 944 15472
rect 984 15440 1016 15472
rect 1056 15440 1088 15472
rect 1128 15440 1160 15472
rect 1200 15440 1232 15472
rect 1272 15440 1304 15472
rect 1344 15440 1376 15472
rect 1416 15440 1448 15472
rect 1488 15440 1520 15472
rect 1560 15440 1592 15472
rect 1632 15440 1664 15472
rect 1704 15440 1736 15472
rect 1776 15440 1808 15472
rect 1848 15440 1880 15472
rect 120 15368 152 15400
rect 192 15368 224 15400
rect 264 15368 296 15400
rect 336 15368 368 15400
rect 408 15368 440 15400
rect 480 15368 512 15400
rect 552 15368 584 15400
rect 624 15368 656 15400
rect 696 15368 728 15400
rect 768 15368 800 15400
rect 840 15368 872 15400
rect 912 15368 944 15400
rect 984 15368 1016 15400
rect 1056 15368 1088 15400
rect 1128 15368 1160 15400
rect 1200 15368 1232 15400
rect 1272 15368 1304 15400
rect 1344 15368 1376 15400
rect 1416 15368 1448 15400
rect 1488 15368 1520 15400
rect 1560 15368 1592 15400
rect 1632 15368 1664 15400
rect 1704 15368 1736 15400
rect 1776 15368 1808 15400
rect 1848 15368 1880 15400
rect 120 15296 152 15328
rect 192 15296 224 15328
rect 264 15296 296 15328
rect 336 15296 368 15328
rect 408 15296 440 15328
rect 480 15296 512 15328
rect 552 15296 584 15328
rect 624 15296 656 15328
rect 696 15296 728 15328
rect 768 15296 800 15328
rect 840 15296 872 15328
rect 912 15296 944 15328
rect 984 15296 1016 15328
rect 1056 15296 1088 15328
rect 1128 15296 1160 15328
rect 1200 15296 1232 15328
rect 1272 15296 1304 15328
rect 1344 15296 1376 15328
rect 1416 15296 1448 15328
rect 1488 15296 1520 15328
rect 1560 15296 1592 15328
rect 1632 15296 1664 15328
rect 1704 15296 1736 15328
rect 1776 15296 1808 15328
rect 1848 15296 1880 15328
rect 120 15224 152 15256
rect 192 15224 224 15256
rect 264 15224 296 15256
rect 336 15224 368 15256
rect 408 15224 440 15256
rect 480 15224 512 15256
rect 552 15224 584 15256
rect 624 15224 656 15256
rect 696 15224 728 15256
rect 768 15224 800 15256
rect 840 15224 872 15256
rect 912 15224 944 15256
rect 984 15224 1016 15256
rect 1056 15224 1088 15256
rect 1128 15224 1160 15256
rect 1200 15224 1232 15256
rect 1272 15224 1304 15256
rect 1344 15224 1376 15256
rect 1416 15224 1448 15256
rect 1488 15224 1520 15256
rect 1560 15224 1592 15256
rect 1632 15224 1664 15256
rect 1704 15224 1736 15256
rect 1776 15224 1808 15256
rect 1848 15224 1880 15256
rect 120 15152 152 15184
rect 192 15152 224 15184
rect 264 15152 296 15184
rect 336 15152 368 15184
rect 408 15152 440 15184
rect 480 15152 512 15184
rect 552 15152 584 15184
rect 624 15152 656 15184
rect 696 15152 728 15184
rect 768 15152 800 15184
rect 840 15152 872 15184
rect 912 15152 944 15184
rect 984 15152 1016 15184
rect 1056 15152 1088 15184
rect 1128 15152 1160 15184
rect 1200 15152 1232 15184
rect 1272 15152 1304 15184
rect 1344 15152 1376 15184
rect 1416 15152 1448 15184
rect 1488 15152 1520 15184
rect 1560 15152 1592 15184
rect 1632 15152 1664 15184
rect 1704 15152 1736 15184
rect 1776 15152 1808 15184
rect 1848 15152 1880 15184
rect 120 15080 152 15112
rect 192 15080 224 15112
rect 264 15080 296 15112
rect 336 15080 368 15112
rect 408 15080 440 15112
rect 480 15080 512 15112
rect 552 15080 584 15112
rect 624 15080 656 15112
rect 696 15080 728 15112
rect 768 15080 800 15112
rect 840 15080 872 15112
rect 912 15080 944 15112
rect 984 15080 1016 15112
rect 1056 15080 1088 15112
rect 1128 15080 1160 15112
rect 1200 15080 1232 15112
rect 1272 15080 1304 15112
rect 1344 15080 1376 15112
rect 1416 15080 1448 15112
rect 1488 15080 1520 15112
rect 1560 15080 1592 15112
rect 1632 15080 1664 15112
rect 1704 15080 1736 15112
rect 1776 15080 1808 15112
rect 1848 15080 1880 15112
rect 120 15008 152 15040
rect 192 15008 224 15040
rect 264 15008 296 15040
rect 336 15008 368 15040
rect 408 15008 440 15040
rect 480 15008 512 15040
rect 552 15008 584 15040
rect 624 15008 656 15040
rect 696 15008 728 15040
rect 768 15008 800 15040
rect 840 15008 872 15040
rect 912 15008 944 15040
rect 984 15008 1016 15040
rect 1056 15008 1088 15040
rect 1128 15008 1160 15040
rect 1200 15008 1232 15040
rect 1272 15008 1304 15040
rect 1344 15008 1376 15040
rect 1416 15008 1448 15040
rect 1488 15008 1520 15040
rect 1560 15008 1592 15040
rect 1632 15008 1664 15040
rect 1704 15008 1736 15040
rect 1776 15008 1808 15040
rect 1848 15008 1880 15040
rect 120 14936 152 14968
rect 192 14936 224 14968
rect 264 14936 296 14968
rect 336 14936 368 14968
rect 408 14936 440 14968
rect 480 14936 512 14968
rect 552 14936 584 14968
rect 624 14936 656 14968
rect 696 14936 728 14968
rect 768 14936 800 14968
rect 840 14936 872 14968
rect 912 14936 944 14968
rect 984 14936 1016 14968
rect 1056 14936 1088 14968
rect 1128 14936 1160 14968
rect 1200 14936 1232 14968
rect 1272 14936 1304 14968
rect 1344 14936 1376 14968
rect 1416 14936 1448 14968
rect 1488 14936 1520 14968
rect 1560 14936 1592 14968
rect 1632 14936 1664 14968
rect 1704 14936 1736 14968
rect 1776 14936 1808 14968
rect 1848 14936 1880 14968
rect 120 14864 152 14896
rect 192 14864 224 14896
rect 264 14864 296 14896
rect 336 14864 368 14896
rect 408 14864 440 14896
rect 480 14864 512 14896
rect 552 14864 584 14896
rect 624 14864 656 14896
rect 696 14864 728 14896
rect 768 14864 800 14896
rect 840 14864 872 14896
rect 912 14864 944 14896
rect 984 14864 1016 14896
rect 1056 14864 1088 14896
rect 1128 14864 1160 14896
rect 1200 14864 1232 14896
rect 1272 14864 1304 14896
rect 1344 14864 1376 14896
rect 1416 14864 1448 14896
rect 1488 14864 1520 14896
rect 1560 14864 1592 14896
rect 1632 14864 1664 14896
rect 1704 14864 1736 14896
rect 1776 14864 1808 14896
rect 1848 14864 1880 14896
rect 120 14792 152 14824
rect 192 14792 224 14824
rect 264 14792 296 14824
rect 336 14792 368 14824
rect 408 14792 440 14824
rect 480 14792 512 14824
rect 552 14792 584 14824
rect 624 14792 656 14824
rect 696 14792 728 14824
rect 768 14792 800 14824
rect 840 14792 872 14824
rect 912 14792 944 14824
rect 984 14792 1016 14824
rect 1056 14792 1088 14824
rect 1128 14792 1160 14824
rect 1200 14792 1232 14824
rect 1272 14792 1304 14824
rect 1344 14792 1376 14824
rect 1416 14792 1448 14824
rect 1488 14792 1520 14824
rect 1560 14792 1592 14824
rect 1632 14792 1664 14824
rect 1704 14792 1736 14824
rect 1776 14792 1808 14824
rect 1848 14792 1880 14824
rect 120 14720 152 14752
rect 192 14720 224 14752
rect 264 14720 296 14752
rect 336 14720 368 14752
rect 408 14720 440 14752
rect 480 14720 512 14752
rect 552 14720 584 14752
rect 624 14720 656 14752
rect 696 14720 728 14752
rect 768 14720 800 14752
rect 840 14720 872 14752
rect 912 14720 944 14752
rect 984 14720 1016 14752
rect 1056 14720 1088 14752
rect 1128 14720 1160 14752
rect 1200 14720 1232 14752
rect 1272 14720 1304 14752
rect 1344 14720 1376 14752
rect 1416 14720 1448 14752
rect 1488 14720 1520 14752
rect 1560 14720 1592 14752
rect 1632 14720 1664 14752
rect 1704 14720 1736 14752
rect 1776 14720 1808 14752
rect 1848 14720 1880 14752
rect 120 14648 152 14680
rect 192 14648 224 14680
rect 264 14648 296 14680
rect 336 14648 368 14680
rect 408 14648 440 14680
rect 480 14648 512 14680
rect 552 14648 584 14680
rect 624 14648 656 14680
rect 696 14648 728 14680
rect 768 14648 800 14680
rect 840 14648 872 14680
rect 912 14648 944 14680
rect 984 14648 1016 14680
rect 1056 14648 1088 14680
rect 1128 14648 1160 14680
rect 1200 14648 1232 14680
rect 1272 14648 1304 14680
rect 1344 14648 1376 14680
rect 1416 14648 1448 14680
rect 1488 14648 1520 14680
rect 1560 14648 1592 14680
rect 1632 14648 1664 14680
rect 1704 14648 1736 14680
rect 1776 14648 1808 14680
rect 1848 14648 1880 14680
rect 120 14576 152 14608
rect 192 14576 224 14608
rect 264 14576 296 14608
rect 336 14576 368 14608
rect 408 14576 440 14608
rect 480 14576 512 14608
rect 552 14576 584 14608
rect 624 14576 656 14608
rect 696 14576 728 14608
rect 768 14576 800 14608
rect 840 14576 872 14608
rect 912 14576 944 14608
rect 984 14576 1016 14608
rect 1056 14576 1088 14608
rect 1128 14576 1160 14608
rect 1200 14576 1232 14608
rect 1272 14576 1304 14608
rect 1344 14576 1376 14608
rect 1416 14576 1448 14608
rect 1488 14576 1520 14608
rect 1560 14576 1592 14608
rect 1632 14576 1664 14608
rect 1704 14576 1736 14608
rect 1776 14576 1808 14608
rect 1848 14576 1880 14608
rect 120 14504 152 14536
rect 192 14504 224 14536
rect 264 14504 296 14536
rect 336 14504 368 14536
rect 408 14504 440 14536
rect 480 14504 512 14536
rect 552 14504 584 14536
rect 624 14504 656 14536
rect 696 14504 728 14536
rect 768 14504 800 14536
rect 840 14504 872 14536
rect 912 14504 944 14536
rect 984 14504 1016 14536
rect 1056 14504 1088 14536
rect 1128 14504 1160 14536
rect 1200 14504 1232 14536
rect 1272 14504 1304 14536
rect 1344 14504 1376 14536
rect 1416 14504 1448 14536
rect 1488 14504 1520 14536
rect 1560 14504 1592 14536
rect 1632 14504 1664 14536
rect 1704 14504 1736 14536
rect 1776 14504 1808 14536
rect 1848 14504 1880 14536
rect 120 14432 152 14464
rect 192 14432 224 14464
rect 264 14432 296 14464
rect 336 14432 368 14464
rect 408 14432 440 14464
rect 480 14432 512 14464
rect 552 14432 584 14464
rect 624 14432 656 14464
rect 696 14432 728 14464
rect 768 14432 800 14464
rect 840 14432 872 14464
rect 912 14432 944 14464
rect 984 14432 1016 14464
rect 1056 14432 1088 14464
rect 1128 14432 1160 14464
rect 1200 14432 1232 14464
rect 1272 14432 1304 14464
rect 1344 14432 1376 14464
rect 1416 14432 1448 14464
rect 1488 14432 1520 14464
rect 1560 14432 1592 14464
rect 1632 14432 1664 14464
rect 1704 14432 1736 14464
rect 1776 14432 1808 14464
rect 1848 14432 1880 14464
rect 120 14360 152 14392
rect 192 14360 224 14392
rect 264 14360 296 14392
rect 336 14360 368 14392
rect 408 14360 440 14392
rect 480 14360 512 14392
rect 552 14360 584 14392
rect 624 14360 656 14392
rect 696 14360 728 14392
rect 768 14360 800 14392
rect 840 14360 872 14392
rect 912 14360 944 14392
rect 984 14360 1016 14392
rect 1056 14360 1088 14392
rect 1128 14360 1160 14392
rect 1200 14360 1232 14392
rect 1272 14360 1304 14392
rect 1344 14360 1376 14392
rect 1416 14360 1448 14392
rect 1488 14360 1520 14392
rect 1560 14360 1592 14392
rect 1632 14360 1664 14392
rect 1704 14360 1736 14392
rect 1776 14360 1808 14392
rect 1848 14360 1880 14392
rect 120 14288 152 14320
rect 192 14288 224 14320
rect 264 14288 296 14320
rect 336 14288 368 14320
rect 408 14288 440 14320
rect 480 14288 512 14320
rect 552 14288 584 14320
rect 624 14288 656 14320
rect 696 14288 728 14320
rect 768 14288 800 14320
rect 840 14288 872 14320
rect 912 14288 944 14320
rect 984 14288 1016 14320
rect 1056 14288 1088 14320
rect 1128 14288 1160 14320
rect 1200 14288 1232 14320
rect 1272 14288 1304 14320
rect 1344 14288 1376 14320
rect 1416 14288 1448 14320
rect 1488 14288 1520 14320
rect 1560 14288 1592 14320
rect 1632 14288 1664 14320
rect 1704 14288 1736 14320
rect 1776 14288 1808 14320
rect 1848 14288 1880 14320
rect 120 14216 152 14248
rect 192 14216 224 14248
rect 264 14216 296 14248
rect 336 14216 368 14248
rect 408 14216 440 14248
rect 480 14216 512 14248
rect 552 14216 584 14248
rect 624 14216 656 14248
rect 696 14216 728 14248
rect 768 14216 800 14248
rect 840 14216 872 14248
rect 912 14216 944 14248
rect 984 14216 1016 14248
rect 1056 14216 1088 14248
rect 1128 14216 1160 14248
rect 1200 14216 1232 14248
rect 1272 14216 1304 14248
rect 1344 14216 1376 14248
rect 1416 14216 1448 14248
rect 1488 14216 1520 14248
rect 1560 14216 1592 14248
rect 1632 14216 1664 14248
rect 1704 14216 1736 14248
rect 1776 14216 1808 14248
rect 1848 14216 1880 14248
rect 120 14144 152 14176
rect 192 14144 224 14176
rect 264 14144 296 14176
rect 336 14144 368 14176
rect 408 14144 440 14176
rect 480 14144 512 14176
rect 552 14144 584 14176
rect 624 14144 656 14176
rect 696 14144 728 14176
rect 768 14144 800 14176
rect 840 14144 872 14176
rect 912 14144 944 14176
rect 984 14144 1016 14176
rect 1056 14144 1088 14176
rect 1128 14144 1160 14176
rect 1200 14144 1232 14176
rect 1272 14144 1304 14176
rect 1344 14144 1376 14176
rect 1416 14144 1448 14176
rect 1488 14144 1520 14176
rect 1560 14144 1592 14176
rect 1632 14144 1664 14176
rect 1704 14144 1736 14176
rect 1776 14144 1808 14176
rect 1848 14144 1880 14176
rect 120 14072 152 14104
rect 192 14072 224 14104
rect 264 14072 296 14104
rect 336 14072 368 14104
rect 408 14072 440 14104
rect 480 14072 512 14104
rect 552 14072 584 14104
rect 624 14072 656 14104
rect 696 14072 728 14104
rect 768 14072 800 14104
rect 840 14072 872 14104
rect 912 14072 944 14104
rect 984 14072 1016 14104
rect 1056 14072 1088 14104
rect 1128 14072 1160 14104
rect 1200 14072 1232 14104
rect 1272 14072 1304 14104
rect 1344 14072 1376 14104
rect 1416 14072 1448 14104
rect 1488 14072 1520 14104
rect 1560 14072 1592 14104
rect 1632 14072 1664 14104
rect 1704 14072 1736 14104
rect 1776 14072 1808 14104
rect 1848 14072 1880 14104
rect 120 14000 152 14032
rect 192 14000 224 14032
rect 264 14000 296 14032
rect 336 14000 368 14032
rect 408 14000 440 14032
rect 480 14000 512 14032
rect 552 14000 584 14032
rect 624 14000 656 14032
rect 696 14000 728 14032
rect 768 14000 800 14032
rect 840 14000 872 14032
rect 912 14000 944 14032
rect 984 14000 1016 14032
rect 1056 14000 1088 14032
rect 1128 14000 1160 14032
rect 1200 14000 1232 14032
rect 1272 14000 1304 14032
rect 1344 14000 1376 14032
rect 1416 14000 1448 14032
rect 1488 14000 1520 14032
rect 1560 14000 1592 14032
rect 1632 14000 1664 14032
rect 1704 14000 1736 14032
rect 1776 14000 1808 14032
rect 1848 14000 1880 14032
rect 120 13928 152 13960
rect 192 13928 224 13960
rect 264 13928 296 13960
rect 336 13928 368 13960
rect 408 13928 440 13960
rect 480 13928 512 13960
rect 552 13928 584 13960
rect 624 13928 656 13960
rect 696 13928 728 13960
rect 768 13928 800 13960
rect 840 13928 872 13960
rect 912 13928 944 13960
rect 984 13928 1016 13960
rect 1056 13928 1088 13960
rect 1128 13928 1160 13960
rect 1200 13928 1232 13960
rect 1272 13928 1304 13960
rect 1344 13928 1376 13960
rect 1416 13928 1448 13960
rect 1488 13928 1520 13960
rect 1560 13928 1592 13960
rect 1632 13928 1664 13960
rect 1704 13928 1736 13960
rect 1776 13928 1808 13960
rect 1848 13928 1880 13960
rect 120 13856 152 13888
rect 192 13856 224 13888
rect 264 13856 296 13888
rect 336 13856 368 13888
rect 408 13856 440 13888
rect 480 13856 512 13888
rect 552 13856 584 13888
rect 624 13856 656 13888
rect 696 13856 728 13888
rect 768 13856 800 13888
rect 840 13856 872 13888
rect 912 13856 944 13888
rect 984 13856 1016 13888
rect 1056 13856 1088 13888
rect 1128 13856 1160 13888
rect 1200 13856 1232 13888
rect 1272 13856 1304 13888
rect 1344 13856 1376 13888
rect 1416 13856 1448 13888
rect 1488 13856 1520 13888
rect 1560 13856 1592 13888
rect 1632 13856 1664 13888
rect 1704 13856 1736 13888
rect 1776 13856 1808 13888
rect 1848 13856 1880 13888
rect 120 13784 152 13816
rect 192 13784 224 13816
rect 264 13784 296 13816
rect 336 13784 368 13816
rect 408 13784 440 13816
rect 480 13784 512 13816
rect 552 13784 584 13816
rect 624 13784 656 13816
rect 696 13784 728 13816
rect 768 13784 800 13816
rect 840 13784 872 13816
rect 912 13784 944 13816
rect 984 13784 1016 13816
rect 1056 13784 1088 13816
rect 1128 13784 1160 13816
rect 1200 13784 1232 13816
rect 1272 13784 1304 13816
rect 1344 13784 1376 13816
rect 1416 13784 1448 13816
rect 1488 13784 1520 13816
rect 1560 13784 1592 13816
rect 1632 13784 1664 13816
rect 1704 13784 1736 13816
rect 1776 13784 1808 13816
rect 1848 13784 1880 13816
rect 120 13712 152 13744
rect 192 13712 224 13744
rect 264 13712 296 13744
rect 336 13712 368 13744
rect 408 13712 440 13744
rect 480 13712 512 13744
rect 552 13712 584 13744
rect 624 13712 656 13744
rect 696 13712 728 13744
rect 768 13712 800 13744
rect 840 13712 872 13744
rect 912 13712 944 13744
rect 984 13712 1016 13744
rect 1056 13712 1088 13744
rect 1128 13712 1160 13744
rect 1200 13712 1232 13744
rect 1272 13712 1304 13744
rect 1344 13712 1376 13744
rect 1416 13712 1448 13744
rect 1488 13712 1520 13744
rect 1560 13712 1592 13744
rect 1632 13712 1664 13744
rect 1704 13712 1736 13744
rect 1776 13712 1808 13744
rect 1848 13712 1880 13744
rect 120 13640 152 13672
rect 192 13640 224 13672
rect 264 13640 296 13672
rect 336 13640 368 13672
rect 408 13640 440 13672
rect 480 13640 512 13672
rect 552 13640 584 13672
rect 624 13640 656 13672
rect 696 13640 728 13672
rect 768 13640 800 13672
rect 840 13640 872 13672
rect 912 13640 944 13672
rect 984 13640 1016 13672
rect 1056 13640 1088 13672
rect 1128 13640 1160 13672
rect 1200 13640 1232 13672
rect 1272 13640 1304 13672
rect 1344 13640 1376 13672
rect 1416 13640 1448 13672
rect 1488 13640 1520 13672
rect 1560 13640 1592 13672
rect 1632 13640 1664 13672
rect 1704 13640 1736 13672
rect 1776 13640 1808 13672
rect 1848 13640 1880 13672
rect 120 13568 152 13600
rect 192 13568 224 13600
rect 264 13568 296 13600
rect 336 13568 368 13600
rect 408 13568 440 13600
rect 480 13568 512 13600
rect 552 13568 584 13600
rect 624 13568 656 13600
rect 696 13568 728 13600
rect 768 13568 800 13600
rect 840 13568 872 13600
rect 912 13568 944 13600
rect 984 13568 1016 13600
rect 1056 13568 1088 13600
rect 1128 13568 1160 13600
rect 1200 13568 1232 13600
rect 1272 13568 1304 13600
rect 1344 13568 1376 13600
rect 1416 13568 1448 13600
rect 1488 13568 1520 13600
rect 1560 13568 1592 13600
rect 1632 13568 1664 13600
rect 1704 13568 1736 13600
rect 1776 13568 1808 13600
rect 1848 13568 1880 13600
rect 120 13496 152 13528
rect 192 13496 224 13528
rect 264 13496 296 13528
rect 336 13496 368 13528
rect 408 13496 440 13528
rect 480 13496 512 13528
rect 552 13496 584 13528
rect 624 13496 656 13528
rect 696 13496 728 13528
rect 768 13496 800 13528
rect 840 13496 872 13528
rect 912 13496 944 13528
rect 984 13496 1016 13528
rect 1056 13496 1088 13528
rect 1128 13496 1160 13528
rect 1200 13496 1232 13528
rect 1272 13496 1304 13528
rect 1344 13496 1376 13528
rect 1416 13496 1448 13528
rect 1488 13496 1520 13528
rect 1560 13496 1592 13528
rect 1632 13496 1664 13528
rect 1704 13496 1736 13528
rect 1776 13496 1808 13528
rect 1848 13496 1880 13528
rect 120 13424 152 13456
rect 192 13424 224 13456
rect 264 13424 296 13456
rect 336 13424 368 13456
rect 408 13424 440 13456
rect 480 13424 512 13456
rect 552 13424 584 13456
rect 624 13424 656 13456
rect 696 13424 728 13456
rect 768 13424 800 13456
rect 840 13424 872 13456
rect 912 13424 944 13456
rect 984 13424 1016 13456
rect 1056 13424 1088 13456
rect 1128 13424 1160 13456
rect 1200 13424 1232 13456
rect 1272 13424 1304 13456
rect 1344 13424 1376 13456
rect 1416 13424 1448 13456
rect 1488 13424 1520 13456
rect 1560 13424 1592 13456
rect 1632 13424 1664 13456
rect 1704 13424 1736 13456
rect 1776 13424 1808 13456
rect 1848 13424 1880 13456
rect 120 13352 152 13384
rect 192 13352 224 13384
rect 264 13352 296 13384
rect 336 13352 368 13384
rect 408 13352 440 13384
rect 480 13352 512 13384
rect 552 13352 584 13384
rect 624 13352 656 13384
rect 696 13352 728 13384
rect 768 13352 800 13384
rect 840 13352 872 13384
rect 912 13352 944 13384
rect 984 13352 1016 13384
rect 1056 13352 1088 13384
rect 1128 13352 1160 13384
rect 1200 13352 1232 13384
rect 1272 13352 1304 13384
rect 1344 13352 1376 13384
rect 1416 13352 1448 13384
rect 1488 13352 1520 13384
rect 1560 13352 1592 13384
rect 1632 13352 1664 13384
rect 1704 13352 1736 13384
rect 1776 13352 1808 13384
rect 1848 13352 1880 13384
rect 120 13280 152 13312
rect 192 13280 224 13312
rect 264 13280 296 13312
rect 336 13280 368 13312
rect 408 13280 440 13312
rect 480 13280 512 13312
rect 552 13280 584 13312
rect 624 13280 656 13312
rect 696 13280 728 13312
rect 768 13280 800 13312
rect 840 13280 872 13312
rect 912 13280 944 13312
rect 984 13280 1016 13312
rect 1056 13280 1088 13312
rect 1128 13280 1160 13312
rect 1200 13280 1232 13312
rect 1272 13280 1304 13312
rect 1344 13280 1376 13312
rect 1416 13280 1448 13312
rect 1488 13280 1520 13312
rect 1560 13280 1592 13312
rect 1632 13280 1664 13312
rect 1704 13280 1736 13312
rect 1776 13280 1808 13312
rect 1848 13280 1880 13312
rect 120 13208 152 13240
rect 192 13208 224 13240
rect 264 13208 296 13240
rect 336 13208 368 13240
rect 408 13208 440 13240
rect 480 13208 512 13240
rect 552 13208 584 13240
rect 624 13208 656 13240
rect 696 13208 728 13240
rect 768 13208 800 13240
rect 840 13208 872 13240
rect 912 13208 944 13240
rect 984 13208 1016 13240
rect 1056 13208 1088 13240
rect 1128 13208 1160 13240
rect 1200 13208 1232 13240
rect 1272 13208 1304 13240
rect 1344 13208 1376 13240
rect 1416 13208 1448 13240
rect 1488 13208 1520 13240
rect 1560 13208 1592 13240
rect 1632 13208 1664 13240
rect 1704 13208 1736 13240
rect 1776 13208 1808 13240
rect 1848 13208 1880 13240
rect 120 13136 152 13168
rect 192 13136 224 13168
rect 264 13136 296 13168
rect 336 13136 368 13168
rect 408 13136 440 13168
rect 480 13136 512 13168
rect 552 13136 584 13168
rect 624 13136 656 13168
rect 696 13136 728 13168
rect 768 13136 800 13168
rect 840 13136 872 13168
rect 912 13136 944 13168
rect 984 13136 1016 13168
rect 1056 13136 1088 13168
rect 1128 13136 1160 13168
rect 1200 13136 1232 13168
rect 1272 13136 1304 13168
rect 1344 13136 1376 13168
rect 1416 13136 1448 13168
rect 1488 13136 1520 13168
rect 1560 13136 1592 13168
rect 1632 13136 1664 13168
rect 1704 13136 1736 13168
rect 1776 13136 1808 13168
rect 1848 13136 1880 13168
rect 120 13064 152 13096
rect 192 13064 224 13096
rect 264 13064 296 13096
rect 336 13064 368 13096
rect 408 13064 440 13096
rect 480 13064 512 13096
rect 552 13064 584 13096
rect 624 13064 656 13096
rect 696 13064 728 13096
rect 768 13064 800 13096
rect 840 13064 872 13096
rect 912 13064 944 13096
rect 984 13064 1016 13096
rect 1056 13064 1088 13096
rect 1128 13064 1160 13096
rect 1200 13064 1232 13096
rect 1272 13064 1304 13096
rect 1344 13064 1376 13096
rect 1416 13064 1448 13096
rect 1488 13064 1520 13096
rect 1560 13064 1592 13096
rect 1632 13064 1664 13096
rect 1704 13064 1736 13096
rect 1776 13064 1808 13096
rect 1848 13064 1880 13096
rect 0 33384 120 33416
rect 152 33384 192 33416
rect 224 33384 264 33416
rect 296 33384 336 33416
rect 368 33384 408 33416
rect 440 33384 480 33416
rect 512 33384 552 33416
rect 584 33384 624 33416
rect 656 33384 696 33416
rect 728 33384 768 33416
rect 800 33384 840 33416
rect 872 33384 912 33416
rect 944 33384 984 33416
rect 1016 33384 1056 33416
rect 1088 33384 1128 33416
rect 1160 33384 1200 33416
rect 1232 33384 1272 33416
rect 1304 33384 1344 33416
rect 1376 33384 1416 33416
rect 1448 33384 1488 33416
rect 1520 33384 1560 33416
rect 1592 33384 1632 33416
rect 1664 33384 1704 33416
rect 1736 33384 1776 33416
rect 1808 33384 1848 33416
rect 1880 33384 2000 33416
rect 0 31384 699 31416
rect 731 31384 768 31416
rect 800 31384 838 31416
rect 870 31384 907 31416
rect 939 31384 978 31416
rect 1010 31384 1048 31416
rect 1080 31384 1116 31416
rect 1148 31384 1186 31416
rect 1218 31384 2000 31416
rect 0 29684 120 29716
rect 152 29684 192 29716
rect 224 29684 264 29716
rect 296 29684 336 29716
rect 368 29684 408 29716
rect 440 29684 480 29716
rect 512 29684 552 29716
rect 584 29684 624 29716
rect 656 29684 696 29716
rect 728 29684 768 29716
rect 800 29684 840 29716
rect 872 29684 912 29716
rect 944 29684 984 29716
rect 1016 29684 1056 29716
rect 1088 29684 1128 29716
rect 1160 29684 1200 29716
rect 1232 29684 1272 29716
rect 1304 29684 1344 29716
rect 1376 29684 1416 29716
rect 1448 29684 1488 29716
rect 1520 29684 1560 29716
rect 1592 29684 1632 29716
rect 1664 29684 1704 29716
rect 1736 29684 1776 29716
rect 1808 29684 1848 29716
rect 1880 29684 2000 29716
rect 0 27971 2000 28034
rect 0 27939 120 27971
rect 152 27939 192 27971
rect 224 27939 264 27971
rect 296 27939 336 27971
rect 368 27939 408 27971
rect 440 27939 480 27971
rect 512 27939 552 27971
rect 584 27939 624 27971
rect 656 27939 696 27971
rect 728 27939 768 27971
rect 800 27939 840 27971
rect 872 27939 912 27971
rect 944 27939 984 27971
rect 1016 27939 1056 27971
rect 1088 27939 1128 27971
rect 1160 27939 1200 27971
rect 1232 27939 1272 27971
rect 1304 27939 1344 27971
rect 1376 27939 1416 27971
rect 1448 27939 1488 27971
rect 1520 27939 1560 27971
rect 1592 27939 1632 27971
rect 1664 27939 1704 27971
rect 1736 27939 1776 27971
rect 1808 27939 1848 27971
rect 1880 27939 2000 27971
rect 0 27899 2000 27939
rect 0 27867 120 27899
rect 152 27867 192 27899
rect 224 27867 264 27899
rect 296 27867 336 27899
rect 368 27867 408 27899
rect 440 27867 480 27899
rect 512 27867 552 27899
rect 584 27867 624 27899
rect 656 27867 696 27899
rect 728 27867 768 27899
rect 800 27867 840 27899
rect 872 27867 912 27899
rect 944 27867 984 27899
rect 1016 27867 1056 27899
rect 1088 27867 1128 27899
rect 1160 27867 1200 27899
rect 1232 27867 1272 27899
rect 1304 27867 1344 27899
rect 1376 27867 1416 27899
rect 1448 27867 1488 27899
rect 1520 27867 1560 27899
rect 1592 27867 1632 27899
rect 1664 27867 1704 27899
rect 1736 27867 1776 27899
rect 1808 27867 1848 27899
rect 1880 27867 2000 27899
rect 0 27827 2000 27867
rect 0 27795 120 27827
rect 152 27795 192 27827
rect 224 27795 264 27827
rect 296 27795 336 27827
rect 368 27795 408 27827
rect 440 27795 480 27827
rect 512 27795 552 27827
rect 584 27795 624 27827
rect 656 27795 696 27827
rect 728 27795 768 27827
rect 800 27795 840 27827
rect 872 27795 912 27827
rect 944 27795 984 27827
rect 1016 27795 1056 27827
rect 1088 27795 1128 27827
rect 1160 27795 1200 27827
rect 1232 27795 1272 27827
rect 1304 27795 1344 27827
rect 1376 27795 1416 27827
rect 1448 27795 1488 27827
rect 1520 27795 1560 27827
rect 1592 27795 1632 27827
rect 1664 27795 1704 27827
rect 1736 27795 1776 27827
rect 1808 27795 1848 27827
rect 1880 27795 2000 27827
rect 0 27755 2000 27795
rect 0 27723 120 27755
rect 152 27723 192 27755
rect 224 27723 264 27755
rect 296 27723 336 27755
rect 368 27723 408 27755
rect 440 27723 480 27755
rect 512 27723 552 27755
rect 584 27723 624 27755
rect 656 27723 696 27755
rect 728 27723 768 27755
rect 800 27723 840 27755
rect 872 27723 912 27755
rect 944 27723 984 27755
rect 1016 27723 1056 27755
rect 1088 27723 1128 27755
rect 1160 27723 1200 27755
rect 1232 27723 1272 27755
rect 1304 27723 1344 27755
rect 1376 27723 1416 27755
rect 1448 27723 1488 27755
rect 1520 27723 1560 27755
rect 1592 27723 1632 27755
rect 1664 27723 1704 27755
rect 1736 27723 1776 27755
rect 1808 27723 1848 27755
rect 1880 27723 2000 27755
rect 0 27683 2000 27723
rect 0 27651 120 27683
rect 152 27651 192 27683
rect 224 27651 264 27683
rect 296 27651 336 27683
rect 368 27651 408 27683
rect 440 27651 480 27683
rect 512 27651 552 27683
rect 584 27651 624 27683
rect 656 27651 696 27683
rect 728 27651 768 27683
rect 800 27651 840 27683
rect 872 27651 912 27683
rect 944 27651 984 27683
rect 1016 27651 1056 27683
rect 1088 27651 1128 27683
rect 1160 27651 1200 27683
rect 1232 27651 1272 27683
rect 1304 27651 1344 27683
rect 1376 27651 1416 27683
rect 1448 27651 1488 27683
rect 1520 27651 1560 27683
rect 1592 27651 1632 27683
rect 1664 27651 1704 27683
rect 1736 27651 1776 27683
rect 1808 27651 1848 27683
rect 1880 27651 2000 27683
rect 0 27611 2000 27651
rect 0 27579 120 27611
rect 152 27579 192 27611
rect 224 27579 264 27611
rect 296 27579 336 27611
rect 368 27579 408 27611
rect 440 27579 480 27611
rect 512 27579 552 27611
rect 584 27579 624 27611
rect 656 27579 696 27611
rect 728 27579 768 27611
rect 800 27579 840 27611
rect 872 27579 912 27611
rect 944 27579 984 27611
rect 1016 27579 1056 27611
rect 1088 27579 1128 27611
rect 1160 27579 1200 27611
rect 1232 27579 1272 27611
rect 1304 27579 1344 27611
rect 1376 27579 1416 27611
rect 1448 27579 1488 27611
rect 1520 27579 1560 27611
rect 1592 27579 1632 27611
rect 1664 27579 1704 27611
rect 1736 27579 1776 27611
rect 1808 27579 1848 27611
rect 1880 27579 2000 27611
rect 0 27539 2000 27579
rect 0 27507 120 27539
rect 152 27507 192 27539
rect 224 27507 264 27539
rect 296 27507 336 27539
rect 368 27507 408 27539
rect 440 27507 480 27539
rect 512 27507 552 27539
rect 584 27507 624 27539
rect 656 27507 696 27539
rect 728 27507 768 27539
rect 800 27507 840 27539
rect 872 27507 912 27539
rect 944 27507 984 27539
rect 1016 27507 1056 27539
rect 1088 27507 1128 27539
rect 1160 27507 1200 27539
rect 1232 27507 1272 27539
rect 1304 27507 1344 27539
rect 1376 27507 1416 27539
rect 1448 27507 1488 27539
rect 1520 27507 1560 27539
rect 1592 27507 1632 27539
rect 1664 27507 1704 27539
rect 1736 27507 1776 27539
rect 1808 27507 1848 27539
rect 1880 27507 2000 27539
rect 0 27467 2000 27507
rect 0 27435 120 27467
rect 152 27435 192 27467
rect 224 27435 264 27467
rect 296 27435 336 27467
rect 368 27435 408 27467
rect 440 27435 480 27467
rect 512 27435 552 27467
rect 584 27435 624 27467
rect 656 27435 696 27467
rect 728 27435 768 27467
rect 800 27435 840 27467
rect 872 27435 912 27467
rect 944 27435 984 27467
rect 1016 27435 1056 27467
rect 1088 27435 1128 27467
rect 1160 27435 1200 27467
rect 1232 27435 1272 27467
rect 1304 27435 1344 27467
rect 1376 27435 1416 27467
rect 1448 27435 1488 27467
rect 1520 27435 1560 27467
rect 1592 27435 1632 27467
rect 1664 27435 1704 27467
rect 1736 27435 1776 27467
rect 1808 27435 1848 27467
rect 1880 27435 2000 27467
rect 0 27395 2000 27435
rect 0 27363 120 27395
rect 152 27363 192 27395
rect 224 27363 264 27395
rect 296 27363 336 27395
rect 368 27363 408 27395
rect 440 27363 480 27395
rect 512 27363 552 27395
rect 584 27363 624 27395
rect 656 27363 696 27395
rect 728 27363 768 27395
rect 800 27363 840 27395
rect 872 27363 912 27395
rect 944 27363 984 27395
rect 1016 27363 1056 27395
rect 1088 27363 1128 27395
rect 1160 27363 1200 27395
rect 1232 27363 1272 27395
rect 1304 27363 1344 27395
rect 1376 27363 1416 27395
rect 1448 27363 1488 27395
rect 1520 27363 1560 27395
rect 1592 27363 1632 27395
rect 1664 27363 1704 27395
rect 1736 27363 1776 27395
rect 1808 27363 1848 27395
rect 1880 27363 2000 27395
rect 0 27323 2000 27363
rect 0 27291 120 27323
rect 152 27291 192 27323
rect 224 27291 264 27323
rect 296 27291 336 27323
rect 368 27291 408 27323
rect 440 27291 480 27323
rect 512 27291 552 27323
rect 584 27291 624 27323
rect 656 27291 696 27323
rect 728 27291 768 27323
rect 800 27291 840 27323
rect 872 27291 912 27323
rect 944 27291 984 27323
rect 1016 27291 1056 27323
rect 1088 27291 1128 27323
rect 1160 27291 1200 27323
rect 1232 27291 1272 27323
rect 1304 27291 1344 27323
rect 1376 27291 1416 27323
rect 1448 27291 1488 27323
rect 1520 27291 1560 27323
rect 1592 27291 1632 27323
rect 1664 27291 1704 27323
rect 1736 27291 1776 27323
rect 1808 27291 1848 27323
rect 1880 27291 2000 27323
rect 0 27251 2000 27291
rect 0 27219 120 27251
rect 152 27219 192 27251
rect 224 27219 264 27251
rect 296 27219 336 27251
rect 368 27219 408 27251
rect 440 27219 480 27251
rect 512 27219 552 27251
rect 584 27219 624 27251
rect 656 27219 696 27251
rect 728 27219 768 27251
rect 800 27219 840 27251
rect 872 27219 912 27251
rect 944 27219 984 27251
rect 1016 27219 1056 27251
rect 1088 27219 1128 27251
rect 1160 27219 1200 27251
rect 1232 27219 1272 27251
rect 1304 27219 1344 27251
rect 1376 27219 1416 27251
rect 1448 27219 1488 27251
rect 1520 27219 1560 27251
rect 1592 27219 1632 27251
rect 1664 27219 1704 27251
rect 1736 27219 1776 27251
rect 1808 27219 1848 27251
rect 1880 27219 2000 27251
rect 0 27179 2000 27219
rect 0 27147 120 27179
rect 152 27147 192 27179
rect 224 27147 264 27179
rect 296 27147 336 27179
rect 368 27147 408 27179
rect 440 27147 480 27179
rect 512 27147 552 27179
rect 584 27147 624 27179
rect 656 27147 696 27179
rect 728 27147 768 27179
rect 800 27147 840 27179
rect 872 27147 912 27179
rect 944 27147 984 27179
rect 1016 27147 1056 27179
rect 1088 27147 1128 27179
rect 1160 27147 1200 27179
rect 1232 27147 1272 27179
rect 1304 27147 1344 27179
rect 1376 27147 1416 27179
rect 1448 27147 1488 27179
rect 1520 27147 1560 27179
rect 1592 27147 1632 27179
rect 1664 27147 1704 27179
rect 1736 27147 1776 27179
rect 1808 27147 1848 27179
rect 1880 27147 2000 27179
rect 0 27107 2000 27147
rect 0 27075 120 27107
rect 152 27075 192 27107
rect 224 27075 264 27107
rect 296 27075 336 27107
rect 368 27075 408 27107
rect 440 27075 480 27107
rect 512 27075 552 27107
rect 584 27075 624 27107
rect 656 27075 696 27107
rect 728 27075 768 27107
rect 800 27075 840 27107
rect 872 27075 912 27107
rect 944 27075 984 27107
rect 1016 27075 1056 27107
rect 1088 27075 1128 27107
rect 1160 27075 1200 27107
rect 1232 27075 1272 27107
rect 1304 27075 1344 27107
rect 1376 27075 1416 27107
rect 1448 27075 1488 27107
rect 1520 27075 1560 27107
rect 1592 27075 1632 27107
rect 1664 27075 1704 27107
rect 1736 27075 1776 27107
rect 1808 27075 1848 27107
rect 1880 27075 2000 27107
rect 0 27035 2000 27075
rect 0 27003 120 27035
rect 152 27003 192 27035
rect 224 27003 264 27035
rect 296 27003 336 27035
rect 368 27003 408 27035
rect 440 27003 480 27035
rect 512 27003 552 27035
rect 584 27003 624 27035
rect 656 27003 696 27035
rect 728 27003 768 27035
rect 800 27003 840 27035
rect 872 27003 912 27035
rect 944 27003 984 27035
rect 1016 27003 1056 27035
rect 1088 27003 1128 27035
rect 1160 27003 1200 27035
rect 1232 27003 1272 27035
rect 1304 27003 1344 27035
rect 1376 27003 1416 27035
rect 1448 27003 1488 27035
rect 1520 27003 1560 27035
rect 1592 27003 1632 27035
rect 1664 27003 1704 27035
rect 1736 27003 1776 27035
rect 1808 27003 1848 27035
rect 1880 27003 2000 27035
rect 0 26963 2000 27003
rect 0 26931 120 26963
rect 152 26931 192 26963
rect 224 26931 264 26963
rect 296 26931 336 26963
rect 368 26931 408 26963
rect 440 26931 480 26963
rect 512 26931 552 26963
rect 584 26931 624 26963
rect 656 26931 696 26963
rect 728 26931 768 26963
rect 800 26931 840 26963
rect 872 26931 912 26963
rect 944 26931 984 26963
rect 1016 26931 1056 26963
rect 1088 26931 1128 26963
rect 1160 26931 1200 26963
rect 1232 26931 1272 26963
rect 1304 26931 1344 26963
rect 1376 26931 1416 26963
rect 1448 26931 1488 26963
rect 1520 26931 1560 26963
rect 1592 26931 1632 26963
rect 1664 26931 1704 26963
rect 1736 26931 1776 26963
rect 1808 26931 1848 26963
rect 1880 26931 2000 26963
rect 0 26891 2000 26931
rect 0 26859 120 26891
rect 152 26859 192 26891
rect 224 26859 264 26891
rect 296 26859 336 26891
rect 368 26859 408 26891
rect 440 26859 480 26891
rect 512 26859 552 26891
rect 584 26859 624 26891
rect 656 26859 696 26891
rect 728 26859 768 26891
rect 800 26859 840 26891
rect 872 26859 912 26891
rect 944 26859 984 26891
rect 1016 26859 1056 26891
rect 1088 26859 1128 26891
rect 1160 26859 1200 26891
rect 1232 26859 1272 26891
rect 1304 26859 1344 26891
rect 1376 26859 1416 26891
rect 1448 26859 1488 26891
rect 1520 26859 1560 26891
rect 1592 26859 1632 26891
rect 1664 26859 1704 26891
rect 1736 26859 1776 26891
rect 1808 26859 1848 26891
rect 1880 26859 2000 26891
rect 0 26819 2000 26859
rect 0 26787 120 26819
rect 152 26787 192 26819
rect 224 26787 264 26819
rect 296 26787 336 26819
rect 368 26787 408 26819
rect 440 26787 480 26819
rect 512 26787 552 26819
rect 584 26787 624 26819
rect 656 26787 696 26819
rect 728 26787 768 26819
rect 800 26787 840 26819
rect 872 26787 912 26819
rect 944 26787 984 26819
rect 1016 26787 1056 26819
rect 1088 26787 1128 26819
rect 1160 26787 1200 26819
rect 1232 26787 1272 26819
rect 1304 26787 1344 26819
rect 1376 26787 1416 26819
rect 1448 26787 1488 26819
rect 1520 26787 1560 26819
rect 1592 26787 1632 26819
rect 1664 26787 1704 26819
rect 1736 26787 1776 26819
rect 1808 26787 1848 26819
rect 1880 26787 2000 26819
rect 0 26747 2000 26787
rect 0 26715 120 26747
rect 152 26715 192 26747
rect 224 26715 264 26747
rect 296 26715 336 26747
rect 368 26715 408 26747
rect 440 26715 480 26747
rect 512 26715 552 26747
rect 584 26715 624 26747
rect 656 26715 696 26747
rect 728 26715 768 26747
rect 800 26715 840 26747
rect 872 26715 912 26747
rect 944 26715 984 26747
rect 1016 26715 1056 26747
rect 1088 26715 1128 26747
rect 1160 26715 1200 26747
rect 1232 26715 1272 26747
rect 1304 26715 1344 26747
rect 1376 26715 1416 26747
rect 1448 26715 1488 26747
rect 1520 26715 1560 26747
rect 1592 26715 1632 26747
rect 1664 26715 1704 26747
rect 1736 26715 1776 26747
rect 1808 26715 1848 26747
rect 1880 26715 2000 26747
rect 0 26675 2000 26715
rect 0 26643 120 26675
rect 152 26643 192 26675
rect 224 26643 264 26675
rect 296 26643 336 26675
rect 368 26643 408 26675
rect 440 26643 480 26675
rect 512 26643 552 26675
rect 584 26643 624 26675
rect 656 26643 696 26675
rect 728 26643 768 26675
rect 800 26643 840 26675
rect 872 26643 912 26675
rect 944 26643 984 26675
rect 1016 26643 1056 26675
rect 1088 26643 1128 26675
rect 1160 26643 1200 26675
rect 1232 26643 1272 26675
rect 1304 26643 1344 26675
rect 1376 26643 1416 26675
rect 1448 26643 1488 26675
rect 1520 26643 1560 26675
rect 1592 26643 1632 26675
rect 1664 26643 1704 26675
rect 1736 26643 1776 26675
rect 1808 26643 1848 26675
rect 1880 26643 2000 26675
rect 0 26603 2000 26643
rect 0 26571 120 26603
rect 152 26571 192 26603
rect 224 26571 264 26603
rect 296 26571 336 26603
rect 368 26571 408 26603
rect 440 26571 480 26603
rect 512 26571 552 26603
rect 584 26571 624 26603
rect 656 26571 696 26603
rect 728 26571 768 26603
rect 800 26571 840 26603
rect 872 26571 912 26603
rect 944 26571 984 26603
rect 1016 26571 1056 26603
rect 1088 26571 1128 26603
rect 1160 26571 1200 26603
rect 1232 26571 1272 26603
rect 1304 26571 1344 26603
rect 1376 26571 1416 26603
rect 1448 26571 1488 26603
rect 1520 26571 1560 26603
rect 1592 26571 1632 26603
rect 1664 26571 1704 26603
rect 1736 26571 1776 26603
rect 1808 26571 1848 26603
rect 1880 26571 2000 26603
rect 0 26531 2000 26571
rect 0 26499 120 26531
rect 152 26499 192 26531
rect 224 26499 264 26531
rect 296 26499 336 26531
rect 368 26499 408 26531
rect 440 26499 480 26531
rect 512 26499 552 26531
rect 584 26499 624 26531
rect 656 26499 696 26531
rect 728 26499 768 26531
rect 800 26499 840 26531
rect 872 26499 912 26531
rect 944 26499 984 26531
rect 1016 26499 1056 26531
rect 1088 26499 1128 26531
rect 1160 26499 1200 26531
rect 1232 26499 1272 26531
rect 1304 26499 1344 26531
rect 1376 26499 1416 26531
rect 1448 26499 1488 26531
rect 1520 26499 1560 26531
rect 1592 26499 1632 26531
rect 1664 26499 1704 26531
rect 1736 26499 1776 26531
rect 1808 26499 1848 26531
rect 1880 26499 2000 26531
rect 0 26459 2000 26499
rect 0 26427 120 26459
rect 152 26427 192 26459
rect 224 26427 264 26459
rect 296 26427 336 26459
rect 368 26427 408 26459
rect 440 26427 480 26459
rect 512 26427 552 26459
rect 584 26427 624 26459
rect 656 26427 696 26459
rect 728 26427 768 26459
rect 800 26427 840 26459
rect 872 26427 912 26459
rect 944 26427 984 26459
rect 1016 26427 1056 26459
rect 1088 26427 1128 26459
rect 1160 26427 1200 26459
rect 1232 26427 1272 26459
rect 1304 26427 1344 26459
rect 1376 26427 1416 26459
rect 1448 26427 1488 26459
rect 1520 26427 1560 26459
rect 1592 26427 1632 26459
rect 1664 26427 1704 26459
rect 1736 26427 1776 26459
rect 1808 26427 1848 26459
rect 1880 26427 2000 26459
rect 0 26387 2000 26427
rect 0 26355 120 26387
rect 152 26355 192 26387
rect 224 26355 264 26387
rect 296 26355 336 26387
rect 368 26355 408 26387
rect 440 26355 480 26387
rect 512 26355 552 26387
rect 584 26355 624 26387
rect 656 26355 696 26387
rect 728 26355 768 26387
rect 800 26355 840 26387
rect 872 26355 912 26387
rect 944 26355 984 26387
rect 1016 26355 1056 26387
rect 1088 26355 1128 26387
rect 1160 26355 1200 26387
rect 1232 26355 1272 26387
rect 1304 26355 1344 26387
rect 1376 26355 1416 26387
rect 1448 26355 1488 26387
rect 1520 26355 1560 26387
rect 1592 26355 1632 26387
rect 1664 26355 1704 26387
rect 1736 26355 1776 26387
rect 1808 26355 1848 26387
rect 1880 26355 2000 26387
rect 0 26315 2000 26355
rect 0 26283 120 26315
rect 152 26283 192 26315
rect 224 26283 264 26315
rect 296 26283 336 26315
rect 368 26283 408 26315
rect 440 26283 480 26315
rect 512 26283 552 26315
rect 584 26283 624 26315
rect 656 26283 696 26315
rect 728 26283 768 26315
rect 800 26283 840 26315
rect 872 26283 912 26315
rect 944 26283 984 26315
rect 1016 26283 1056 26315
rect 1088 26283 1128 26315
rect 1160 26283 1200 26315
rect 1232 26283 1272 26315
rect 1304 26283 1344 26315
rect 1376 26283 1416 26315
rect 1448 26283 1488 26315
rect 1520 26283 1560 26315
rect 1592 26283 1632 26315
rect 1664 26283 1704 26315
rect 1736 26283 1776 26315
rect 1808 26283 1848 26315
rect 1880 26283 2000 26315
rect 0 26243 2000 26283
rect 0 26211 120 26243
rect 152 26211 192 26243
rect 224 26211 264 26243
rect 296 26211 336 26243
rect 368 26211 408 26243
rect 440 26211 480 26243
rect 512 26211 552 26243
rect 584 26211 624 26243
rect 656 26211 696 26243
rect 728 26211 768 26243
rect 800 26211 840 26243
rect 872 26211 912 26243
rect 944 26211 984 26243
rect 1016 26211 1056 26243
rect 1088 26211 1128 26243
rect 1160 26211 1200 26243
rect 1232 26211 1272 26243
rect 1304 26211 1344 26243
rect 1376 26211 1416 26243
rect 1448 26211 1488 26243
rect 1520 26211 1560 26243
rect 1592 26211 1632 26243
rect 1664 26211 1704 26243
rect 1736 26211 1776 26243
rect 1808 26211 1848 26243
rect 1880 26211 2000 26243
rect 0 26171 2000 26211
rect 0 26139 120 26171
rect 152 26139 192 26171
rect 224 26139 264 26171
rect 296 26139 336 26171
rect 368 26139 408 26171
rect 440 26139 480 26171
rect 512 26139 552 26171
rect 584 26139 624 26171
rect 656 26139 696 26171
rect 728 26139 768 26171
rect 800 26139 840 26171
rect 872 26139 912 26171
rect 944 26139 984 26171
rect 1016 26139 1056 26171
rect 1088 26139 1128 26171
rect 1160 26139 1200 26171
rect 1232 26139 1272 26171
rect 1304 26139 1344 26171
rect 1376 26139 1416 26171
rect 1448 26139 1488 26171
rect 1520 26139 1560 26171
rect 1592 26139 1632 26171
rect 1664 26139 1704 26171
rect 1736 26139 1776 26171
rect 1808 26139 1848 26171
rect 1880 26139 2000 26171
rect 0 26099 2000 26139
rect 0 26067 120 26099
rect 152 26067 192 26099
rect 224 26067 264 26099
rect 296 26067 336 26099
rect 368 26067 408 26099
rect 440 26067 480 26099
rect 512 26067 552 26099
rect 584 26067 624 26099
rect 656 26067 696 26099
rect 728 26067 768 26099
rect 800 26067 840 26099
rect 872 26067 912 26099
rect 944 26067 984 26099
rect 1016 26067 1056 26099
rect 1088 26067 1128 26099
rect 1160 26067 1200 26099
rect 1232 26067 1272 26099
rect 1304 26067 1344 26099
rect 1376 26067 1416 26099
rect 1448 26067 1488 26099
rect 1520 26067 1560 26099
rect 1592 26067 1632 26099
rect 1664 26067 1704 26099
rect 1736 26067 1776 26099
rect 1808 26067 1848 26099
rect 1880 26067 2000 26099
rect 0 26027 2000 26067
rect 0 25995 120 26027
rect 152 25995 192 26027
rect 224 25995 264 26027
rect 296 25995 336 26027
rect 368 25995 408 26027
rect 440 25995 480 26027
rect 512 25995 552 26027
rect 584 25995 624 26027
rect 656 25995 696 26027
rect 728 25995 768 26027
rect 800 25995 840 26027
rect 872 25995 912 26027
rect 944 25995 984 26027
rect 1016 25995 1056 26027
rect 1088 25995 1128 26027
rect 1160 25995 1200 26027
rect 1232 25995 1272 26027
rect 1304 25995 1344 26027
rect 1376 25995 1416 26027
rect 1448 25995 1488 26027
rect 1520 25995 1560 26027
rect 1592 25995 1632 26027
rect 1664 25995 1704 26027
rect 1736 25995 1776 26027
rect 1808 25995 1848 26027
rect 1880 25995 2000 26027
rect 0 25955 2000 25995
rect 0 25923 120 25955
rect 152 25923 192 25955
rect 224 25923 264 25955
rect 296 25923 336 25955
rect 368 25923 408 25955
rect 440 25923 480 25955
rect 512 25923 552 25955
rect 584 25923 624 25955
rect 656 25923 696 25955
rect 728 25923 768 25955
rect 800 25923 840 25955
rect 872 25923 912 25955
rect 944 25923 984 25955
rect 1016 25923 1056 25955
rect 1088 25923 1128 25955
rect 1160 25923 1200 25955
rect 1232 25923 1272 25955
rect 1304 25923 1344 25955
rect 1376 25923 1416 25955
rect 1448 25923 1488 25955
rect 1520 25923 1560 25955
rect 1592 25923 1632 25955
rect 1664 25923 1704 25955
rect 1736 25923 1776 25955
rect 1808 25923 1848 25955
rect 1880 25923 2000 25955
rect 0 25883 2000 25923
rect 0 25851 120 25883
rect 152 25851 192 25883
rect 224 25851 264 25883
rect 296 25851 336 25883
rect 368 25851 408 25883
rect 440 25851 480 25883
rect 512 25851 552 25883
rect 584 25851 624 25883
rect 656 25851 696 25883
rect 728 25851 768 25883
rect 800 25851 840 25883
rect 872 25851 912 25883
rect 944 25851 984 25883
rect 1016 25851 1056 25883
rect 1088 25851 1128 25883
rect 1160 25851 1200 25883
rect 1232 25851 1272 25883
rect 1304 25851 1344 25883
rect 1376 25851 1416 25883
rect 1448 25851 1488 25883
rect 1520 25851 1560 25883
rect 1592 25851 1632 25883
rect 1664 25851 1704 25883
rect 1736 25851 1776 25883
rect 1808 25851 1848 25883
rect 1880 25851 2000 25883
rect 0 25811 2000 25851
rect 0 25779 120 25811
rect 152 25779 192 25811
rect 224 25779 264 25811
rect 296 25779 336 25811
rect 368 25779 408 25811
rect 440 25779 480 25811
rect 512 25779 552 25811
rect 584 25779 624 25811
rect 656 25779 696 25811
rect 728 25779 768 25811
rect 800 25779 840 25811
rect 872 25779 912 25811
rect 944 25779 984 25811
rect 1016 25779 1056 25811
rect 1088 25779 1128 25811
rect 1160 25779 1200 25811
rect 1232 25779 1272 25811
rect 1304 25779 1344 25811
rect 1376 25779 1416 25811
rect 1448 25779 1488 25811
rect 1520 25779 1560 25811
rect 1592 25779 1632 25811
rect 1664 25779 1704 25811
rect 1736 25779 1776 25811
rect 1808 25779 1848 25811
rect 1880 25779 2000 25811
rect 0 25739 2000 25779
rect 0 25707 120 25739
rect 152 25707 192 25739
rect 224 25707 264 25739
rect 296 25707 336 25739
rect 368 25707 408 25739
rect 440 25707 480 25739
rect 512 25707 552 25739
rect 584 25707 624 25739
rect 656 25707 696 25739
rect 728 25707 768 25739
rect 800 25707 840 25739
rect 872 25707 912 25739
rect 944 25707 984 25739
rect 1016 25707 1056 25739
rect 1088 25707 1128 25739
rect 1160 25707 1200 25739
rect 1232 25707 1272 25739
rect 1304 25707 1344 25739
rect 1376 25707 1416 25739
rect 1448 25707 1488 25739
rect 1520 25707 1560 25739
rect 1592 25707 1632 25739
rect 1664 25707 1704 25739
rect 1736 25707 1776 25739
rect 1808 25707 1848 25739
rect 1880 25707 2000 25739
rect 0 25667 2000 25707
rect 0 25635 120 25667
rect 152 25635 192 25667
rect 224 25635 264 25667
rect 296 25635 336 25667
rect 368 25635 408 25667
rect 440 25635 480 25667
rect 512 25635 552 25667
rect 584 25635 624 25667
rect 656 25635 696 25667
rect 728 25635 768 25667
rect 800 25635 840 25667
rect 872 25635 912 25667
rect 944 25635 984 25667
rect 1016 25635 1056 25667
rect 1088 25635 1128 25667
rect 1160 25635 1200 25667
rect 1232 25635 1272 25667
rect 1304 25635 1344 25667
rect 1376 25635 1416 25667
rect 1448 25635 1488 25667
rect 1520 25635 1560 25667
rect 1592 25635 1632 25667
rect 1664 25635 1704 25667
rect 1736 25635 1776 25667
rect 1808 25635 1848 25667
rect 1880 25635 2000 25667
rect 0 25595 2000 25635
rect 0 25563 120 25595
rect 152 25563 192 25595
rect 224 25563 264 25595
rect 296 25563 336 25595
rect 368 25563 408 25595
rect 440 25563 480 25595
rect 512 25563 552 25595
rect 584 25563 624 25595
rect 656 25563 696 25595
rect 728 25563 768 25595
rect 800 25563 840 25595
rect 872 25563 912 25595
rect 944 25563 984 25595
rect 1016 25563 1056 25595
rect 1088 25563 1128 25595
rect 1160 25563 1200 25595
rect 1232 25563 1272 25595
rect 1304 25563 1344 25595
rect 1376 25563 1416 25595
rect 1448 25563 1488 25595
rect 1520 25563 1560 25595
rect 1592 25563 1632 25595
rect 1664 25563 1704 25595
rect 1736 25563 1776 25595
rect 1808 25563 1848 25595
rect 1880 25563 2000 25595
rect 0 25523 2000 25563
rect 0 25491 120 25523
rect 152 25491 192 25523
rect 224 25491 264 25523
rect 296 25491 336 25523
rect 368 25491 408 25523
rect 440 25491 480 25523
rect 512 25491 552 25523
rect 584 25491 624 25523
rect 656 25491 696 25523
rect 728 25491 768 25523
rect 800 25491 840 25523
rect 872 25491 912 25523
rect 944 25491 984 25523
rect 1016 25491 1056 25523
rect 1088 25491 1128 25523
rect 1160 25491 1200 25523
rect 1232 25491 1272 25523
rect 1304 25491 1344 25523
rect 1376 25491 1416 25523
rect 1448 25491 1488 25523
rect 1520 25491 1560 25523
rect 1592 25491 1632 25523
rect 1664 25491 1704 25523
rect 1736 25491 1776 25523
rect 1808 25491 1848 25523
rect 1880 25491 2000 25523
rect 0 25451 2000 25491
rect 0 25419 120 25451
rect 152 25419 192 25451
rect 224 25419 264 25451
rect 296 25419 336 25451
rect 368 25419 408 25451
rect 440 25419 480 25451
rect 512 25419 552 25451
rect 584 25419 624 25451
rect 656 25419 696 25451
rect 728 25419 768 25451
rect 800 25419 840 25451
rect 872 25419 912 25451
rect 944 25419 984 25451
rect 1016 25419 1056 25451
rect 1088 25419 1128 25451
rect 1160 25419 1200 25451
rect 1232 25419 1272 25451
rect 1304 25419 1344 25451
rect 1376 25419 1416 25451
rect 1448 25419 1488 25451
rect 1520 25419 1560 25451
rect 1592 25419 1632 25451
rect 1664 25419 1704 25451
rect 1736 25419 1776 25451
rect 1808 25419 1848 25451
rect 1880 25419 2000 25451
rect 0 25379 2000 25419
rect 0 25347 120 25379
rect 152 25347 192 25379
rect 224 25347 264 25379
rect 296 25347 336 25379
rect 368 25347 408 25379
rect 440 25347 480 25379
rect 512 25347 552 25379
rect 584 25347 624 25379
rect 656 25347 696 25379
rect 728 25347 768 25379
rect 800 25347 840 25379
rect 872 25347 912 25379
rect 944 25347 984 25379
rect 1016 25347 1056 25379
rect 1088 25347 1128 25379
rect 1160 25347 1200 25379
rect 1232 25347 1272 25379
rect 1304 25347 1344 25379
rect 1376 25347 1416 25379
rect 1448 25347 1488 25379
rect 1520 25347 1560 25379
rect 1592 25347 1632 25379
rect 1664 25347 1704 25379
rect 1736 25347 1776 25379
rect 1808 25347 1848 25379
rect 1880 25347 2000 25379
rect 0 25307 2000 25347
rect 0 25275 120 25307
rect 152 25275 192 25307
rect 224 25275 264 25307
rect 296 25275 336 25307
rect 368 25275 408 25307
rect 440 25275 480 25307
rect 512 25275 552 25307
rect 584 25275 624 25307
rect 656 25275 696 25307
rect 728 25275 768 25307
rect 800 25275 840 25307
rect 872 25275 912 25307
rect 944 25275 984 25307
rect 1016 25275 1056 25307
rect 1088 25275 1128 25307
rect 1160 25275 1200 25307
rect 1232 25275 1272 25307
rect 1304 25275 1344 25307
rect 1376 25275 1416 25307
rect 1448 25275 1488 25307
rect 1520 25275 1560 25307
rect 1592 25275 1632 25307
rect 1664 25275 1704 25307
rect 1736 25275 1776 25307
rect 1808 25275 1848 25307
rect 1880 25275 2000 25307
rect 0 25235 2000 25275
rect 0 25203 120 25235
rect 152 25203 192 25235
rect 224 25203 264 25235
rect 296 25203 336 25235
rect 368 25203 408 25235
rect 440 25203 480 25235
rect 512 25203 552 25235
rect 584 25203 624 25235
rect 656 25203 696 25235
rect 728 25203 768 25235
rect 800 25203 840 25235
rect 872 25203 912 25235
rect 944 25203 984 25235
rect 1016 25203 1056 25235
rect 1088 25203 1128 25235
rect 1160 25203 1200 25235
rect 1232 25203 1272 25235
rect 1304 25203 1344 25235
rect 1376 25203 1416 25235
rect 1448 25203 1488 25235
rect 1520 25203 1560 25235
rect 1592 25203 1632 25235
rect 1664 25203 1704 25235
rect 1736 25203 1776 25235
rect 1808 25203 1848 25235
rect 1880 25203 2000 25235
rect 0 25163 2000 25203
rect 0 25131 120 25163
rect 152 25131 192 25163
rect 224 25131 264 25163
rect 296 25131 336 25163
rect 368 25131 408 25163
rect 440 25131 480 25163
rect 512 25131 552 25163
rect 584 25131 624 25163
rect 656 25131 696 25163
rect 728 25131 768 25163
rect 800 25131 840 25163
rect 872 25131 912 25163
rect 944 25131 984 25163
rect 1016 25131 1056 25163
rect 1088 25131 1128 25163
rect 1160 25131 1200 25163
rect 1232 25131 1272 25163
rect 1304 25131 1344 25163
rect 1376 25131 1416 25163
rect 1448 25131 1488 25163
rect 1520 25131 1560 25163
rect 1592 25131 1632 25163
rect 1664 25131 1704 25163
rect 1736 25131 1776 25163
rect 1808 25131 1848 25163
rect 1880 25131 2000 25163
rect 0 25091 2000 25131
rect 0 25059 120 25091
rect 152 25059 192 25091
rect 224 25059 264 25091
rect 296 25059 336 25091
rect 368 25059 408 25091
rect 440 25059 480 25091
rect 512 25059 552 25091
rect 584 25059 624 25091
rect 656 25059 696 25091
rect 728 25059 768 25091
rect 800 25059 840 25091
rect 872 25059 912 25091
rect 944 25059 984 25091
rect 1016 25059 1056 25091
rect 1088 25059 1128 25091
rect 1160 25059 1200 25091
rect 1232 25059 1272 25091
rect 1304 25059 1344 25091
rect 1376 25059 1416 25091
rect 1448 25059 1488 25091
rect 1520 25059 1560 25091
rect 1592 25059 1632 25091
rect 1664 25059 1704 25091
rect 1736 25059 1776 25091
rect 1808 25059 1848 25091
rect 1880 25059 2000 25091
rect 0 25019 2000 25059
rect 0 24987 120 25019
rect 152 24987 192 25019
rect 224 24987 264 25019
rect 296 24987 336 25019
rect 368 24987 408 25019
rect 440 24987 480 25019
rect 512 24987 552 25019
rect 584 24987 624 25019
rect 656 24987 696 25019
rect 728 24987 768 25019
rect 800 24987 840 25019
rect 872 24987 912 25019
rect 944 24987 984 25019
rect 1016 24987 1056 25019
rect 1088 24987 1128 25019
rect 1160 24987 1200 25019
rect 1232 24987 1272 25019
rect 1304 24987 1344 25019
rect 1376 24987 1416 25019
rect 1448 24987 1488 25019
rect 1520 24987 1560 25019
rect 1592 24987 1632 25019
rect 1664 24987 1704 25019
rect 1736 24987 1776 25019
rect 1808 24987 1848 25019
rect 1880 24987 2000 25019
rect 0 24947 2000 24987
rect 0 24915 120 24947
rect 152 24915 192 24947
rect 224 24915 264 24947
rect 296 24915 336 24947
rect 368 24915 408 24947
rect 440 24915 480 24947
rect 512 24915 552 24947
rect 584 24915 624 24947
rect 656 24915 696 24947
rect 728 24915 768 24947
rect 800 24915 840 24947
rect 872 24915 912 24947
rect 944 24915 984 24947
rect 1016 24915 1056 24947
rect 1088 24915 1128 24947
rect 1160 24915 1200 24947
rect 1232 24915 1272 24947
rect 1304 24915 1344 24947
rect 1376 24915 1416 24947
rect 1448 24915 1488 24947
rect 1520 24915 1560 24947
rect 1592 24915 1632 24947
rect 1664 24915 1704 24947
rect 1736 24915 1776 24947
rect 1808 24915 1848 24947
rect 1880 24915 2000 24947
rect 0 24875 2000 24915
rect 0 24843 120 24875
rect 152 24843 192 24875
rect 224 24843 264 24875
rect 296 24843 336 24875
rect 368 24843 408 24875
rect 440 24843 480 24875
rect 512 24843 552 24875
rect 584 24843 624 24875
rect 656 24843 696 24875
rect 728 24843 768 24875
rect 800 24843 840 24875
rect 872 24843 912 24875
rect 944 24843 984 24875
rect 1016 24843 1056 24875
rect 1088 24843 1128 24875
rect 1160 24843 1200 24875
rect 1232 24843 1272 24875
rect 1304 24843 1344 24875
rect 1376 24843 1416 24875
rect 1448 24843 1488 24875
rect 1520 24843 1560 24875
rect 1592 24843 1632 24875
rect 1664 24843 1704 24875
rect 1736 24843 1776 24875
rect 1808 24843 1848 24875
rect 1880 24843 2000 24875
rect 0 24803 2000 24843
rect 0 24771 120 24803
rect 152 24771 192 24803
rect 224 24771 264 24803
rect 296 24771 336 24803
rect 368 24771 408 24803
rect 440 24771 480 24803
rect 512 24771 552 24803
rect 584 24771 624 24803
rect 656 24771 696 24803
rect 728 24771 768 24803
rect 800 24771 840 24803
rect 872 24771 912 24803
rect 944 24771 984 24803
rect 1016 24771 1056 24803
rect 1088 24771 1128 24803
rect 1160 24771 1200 24803
rect 1232 24771 1272 24803
rect 1304 24771 1344 24803
rect 1376 24771 1416 24803
rect 1448 24771 1488 24803
rect 1520 24771 1560 24803
rect 1592 24771 1632 24803
rect 1664 24771 1704 24803
rect 1736 24771 1776 24803
rect 1808 24771 1848 24803
rect 1880 24771 2000 24803
rect 0 24731 2000 24771
rect 0 24699 120 24731
rect 152 24699 192 24731
rect 224 24699 264 24731
rect 296 24699 336 24731
rect 368 24699 408 24731
rect 440 24699 480 24731
rect 512 24699 552 24731
rect 584 24699 624 24731
rect 656 24699 696 24731
rect 728 24699 768 24731
rect 800 24699 840 24731
rect 872 24699 912 24731
rect 944 24699 984 24731
rect 1016 24699 1056 24731
rect 1088 24699 1128 24731
rect 1160 24699 1200 24731
rect 1232 24699 1272 24731
rect 1304 24699 1344 24731
rect 1376 24699 1416 24731
rect 1448 24699 1488 24731
rect 1520 24699 1560 24731
rect 1592 24699 1632 24731
rect 1664 24699 1704 24731
rect 1736 24699 1776 24731
rect 1808 24699 1848 24731
rect 1880 24699 2000 24731
rect 0 24659 2000 24699
rect 0 24627 120 24659
rect 152 24627 192 24659
rect 224 24627 264 24659
rect 296 24627 336 24659
rect 368 24627 408 24659
rect 440 24627 480 24659
rect 512 24627 552 24659
rect 584 24627 624 24659
rect 656 24627 696 24659
rect 728 24627 768 24659
rect 800 24627 840 24659
rect 872 24627 912 24659
rect 944 24627 984 24659
rect 1016 24627 1056 24659
rect 1088 24627 1128 24659
rect 1160 24627 1200 24659
rect 1232 24627 1272 24659
rect 1304 24627 1344 24659
rect 1376 24627 1416 24659
rect 1448 24627 1488 24659
rect 1520 24627 1560 24659
rect 1592 24627 1632 24659
rect 1664 24627 1704 24659
rect 1736 24627 1776 24659
rect 1808 24627 1848 24659
rect 1880 24627 2000 24659
rect 0 24587 2000 24627
rect 0 24555 120 24587
rect 152 24555 192 24587
rect 224 24555 264 24587
rect 296 24555 336 24587
rect 368 24555 408 24587
rect 440 24555 480 24587
rect 512 24555 552 24587
rect 584 24555 624 24587
rect 656 24555 696 24587
rect 728 24555 768 24587
rect 800 24555 840 24587
rect 872 24555 912 24587
rect 944 24555 984 24587
rect 1016 24555 1056 24587
rect 1088 24555 1128 24587
rect 1160 24555 1200 24587
rect 1232 24555 1272 24587
rect 1304 24555 1344 24587
rect 1376 24555 1416 24587
rect 1448 24555 1488 24587
rect 1520 24555 1560 24587
rect 1592 24555 1632 24587
rect 1664 24555 1704 24587
rect 1736 24555 1776 24587
rect 1808 24555 1848 24587
rect 1880 24555 2000 24587
rect 0 24515 2000 24555
rect 0 24483 120 24515
rect 152 24483 192 24515
rect 224 24483 264 24515
rect 296 24483 336 24515
rect 368 24483 408 24515
rect 440 24483 480 24515
rect 512 24483 552 24515
rect 584 24483 624 24515
rect 656 24483 696 24515
rect 728 24483 768 24515
rect 800 24483 840 24515
rect 872 24483 912 24515
rect 944 24483 984 24515
rect 1016 24483 1056 24515
rect 1088 24483 1128 24515
rect 1160 24483 1200 24515
rect 1232 24483 1272 24515
rect 1304 24483 1344 24515
rect 1376 24483 1416 24515
rect 1448 24483 1488 24515
rect 1520 24483 1560 24515
rect 1592 24483 1632 24515
rect 1664 24483 1704 24515
rect 1736 24483 1776 24515
rect 1808 24483 1848 24515
rect 1880 24483 2000 24515
rect 0 24443 2000 24483
rect 0 24411 120 24443
rect 152 24411 192 24443
rect 224 24411 264 24443
rect 296 24411 336 24443
rect 368 24411 408 24443
rect 440 24411 480 24443
rect 512 24411 552 24443
rect 584 24411 624 24443
rect 656 24411 696 24443
rect 728 24411 768 24443
rect 800 24411 840 24443
rect 872 24411 912 24443
rect 944 24411 984 24443
rect 1016 24411 1056 24443
rect 1088 24411 1128 24443
rect 1160 24411 1200 24443
rect 1232 24411 1272 24443
rect 1304 24411 1344 24443
rect 1376 24411 1416 24443
rect 1448 24411 1488 24443
rect 1520 24411 1560 24443
rect 1592 24411 1632 24443
rect 1664 24411 1704 24443
rect 1736 24411 1776 24443
rect 1808 24411 1848 24443
rect 1880 24411 2000 24443
rect 0 24371 2000 24411
rect 0 24339 120 24371
rect 152 24339 192 24371
rect 224 24339 264 24371
rect 296 24339 336 24371
rect 368 24339 408 24371
rect 440 24339 480 24371
rect 512 24339 552 24371
rect 584 24339 624 24371
rect 656 24339 696 24371
rect 728 24339 768 24371
rect 800 24339 840 24371
rect 872 24339 912 24371
rect 944 24339 984 24371
rect 1016 24339 1056 24371
rect 1088 24339 1128 24371
rect 1160 24339 1200 24371
rect 1232 24339 1272 24371
rect 1304 24339 1344 24371
rect 1376 24339 1416 24371
rect 1448 24339 1488 24371
rect 1520 24339 1560 24371
rect 1592 24339 1632 24371
rect 1664 24339 1704 24371
rect 1736 24339 1776 24371
rect 1808 24339 1848 24371
rect 1880 24339 2000 24371
rect 0 24299 2000 24339
rect 0 24267 120 24299
rect 152 24267 192 24299
rect 224 24267 264 24299
rect 296 24267 336 24299
rect 368 24267 408 24299
rect 440 24267 480 24299
rect 512 24267 552 24299
rect 584 24267 624 24299
rect 656 24267 696 24299
rect 728 24267 768 24299
rect 800 24267 840 24299
rect 872 24267 912 24299
rect 944 24267 984 24299
rect 1016 24267 1056 24299
rect 1088 24267 1128 24299
rect 1160 24267 1200 24299
rect 1232 24267 1272 24299
rect 1304 24267 1344 24299
rect 1376 24267 1416 24299
rect 1448 24267 1488 24299
rect 1520 24267 1560 24299
rect 1592 24267 1632 24299
rect 1664 24267 1704 24299
rect 1736 24267 1776 24299
rect 1808 24267 1848 24299
rect 1880 24267 2000 24299
rect 0 24227 2000 24267
rect 0 24195 120 24227
rect 152 24195 192 24227
rect 224 24195 264 24227
rect 296 24195 336 24227
rect 368 24195 408 24227
rect 440 24195 480 24227
rect 512 24195 552 24227
rect 584 24195 624 24227
rect 656 24195 696 24227
rect 728 24195 768 24227
rect 800 24195 840 24227
rect 872 24195 912 24227
rect 944 24195 984 24227
rect 1016 24195 1056 24227
rect 1088 24195 1128 24227
rect 1160 24195 1200 24227
rect 1232 24195 1272 24227
rect 1304 24195 1344 24227
rect 1376 24195 1416 24227
rect 1448 24195 1488 24227
rect 1520 24195 1560 24227
rect 1592 24195 1632 24227
rect 1664 24195 1704 24227
rect 1736 24195 1776 24227
rect 1808 24195 1848 24227
rect 1880 24195 2000 24227
rect 0 24155 2000 24195
rect 0 24123 120 24155
rect 152 24123 192 24155
rect 224 24123 264 24155
rect 296 24123 336 24155
rect 368 24123 408 24155
rect 440 24123 480 24155
rect 512 24123 552 24155
rect 584 24123 624 24155
rect 656 24123 696 24155
rect 728 24123 768 24155
rect 800 24123 840 24155
rect 872 24123 912 24155
rect 944 24123 984 24155
rect 1016 24123 1056 24155
rect 1088 24123 1128 24155
rect 1160 24123 1200 24155
rect 1232 24123 1272 24155
rect 1304 24123 1344 24155
rect 1376 24123 1416 24155
rect 1448 24123 1488 24155
rect 1520 24123 1560 24155
rect 1592 24123 1632 24155
rect 1664 24123 1704 24155
rect 1736 24123 1776 24155
rect 1808 24123 1848 24155
rect 1880 24123 2000 24155
rect 0 24083 2000 24123
rect 0 24051 120 24083
rect 152 24051 192 24083
rect 224 24051 264 24083
rect 296 24051 336 24083
rect 368 24051 408 24083
rect 440 24051 480 24083
rect 512 24051 552 24083
rect 584 24051 624 24083
rect 656 24051 696 24083
rect 728 24051 768 24083
rect 800 24051 840 24083
rect 872 24051 912 24083
rect 944 24051 984 24083
rect 1016 24051 1056 24083
rect 1088 24051 1128 24083
rect 1160 24051 1200 24083
rect 1232 24051 1272 24083
rect 1304 24051 1344 24083
rect 1376 24051 1416 24083
rect 1448 24051 1488 24083
rect 1520 24051 1560 24083
rect 1592 24051 1632 24083
rect 1664 24051 1704 24083
rect 1736 24051 1776 24083
rect 1808 24051 1848 24083
rect 1880 24051 2000 24083
rect 0 24011 2000 24051
rect 0 23979 120 24011
rect 152 23979 192 24011
rect 224 23979 264 24011
rect 296 23979 336 24011
rect 368 23979 408 24011
rect 440 23979 480 24011
rect 512 23979 552 24011
rect 584 23979 624 24011
rect 656 23979 696 24011
rect 728 23979 768 24011
rect 800 23979 840 24011
rect 872 23979 912 24011
rect 944 23979 984 24011
rect 1016 23979 1056 24011
rect 1088 23979 1128 24011
rect 1160 23979 1200 24011
rect 1232 23979 1272 24011
rect 1304 23979 1344 24011
rect 1376 23979 1416 24011
rect 1448 23979 1488 24011
rect 1520 23979 1560 24011
rect 1592 23979 1632 24011
rect 1664 23979 1704 24011
rect 1736 23979 1776 24011
rect 1808 23979 1848 24011
rect 1880 23979 2000 24011
rect 0 23939 2000 23979
rect 0 23907 120 23939
rect 152 23907 192 23939
rect 224 23907 264 23939
rect 296 23907 336 23939
rect 368 23907 408 23939
rect 440 23907 480 23939
rect 512 23907 552 23939
rect 584 23907 624 23939
rect 656 23907 696 23939
rect 728 23907 768 23939
rect 800 23907 840 23939
rect 872 23907 912 23939
rect 944 23907 984 23939
rect 1016 23907 1056 23939
rect 1088 23907 1128 23939
rect 1160 23907 1200 23939
rect 1232 23907 1272 23939
rect 1304 23907 1344 23939
rect 1376 23907 1416 23939
rect 1448 23907 1488 23939
rect 1520 23907 1560 23939
rect 1592 23907 1632 23939
rect 1664 23907 1704 23939
rect 1736 23907 1776 23939
rect 1808 23907 1848 23939
rect 1880 23907 2000 23939
rect 0 23867 2000 23907
rect 0 23835 120 23867
rect 152 23835 192 23867
rect 224 23835 264 23867
rect 296 23835 336 23867
rect 368 23835 408 23867
rect 440 23835 480 23867
rect 512 23835 552 23867
rect 584 23835 624 23867
rect 656 23835 696 23867
rect 728 23835 768 23867
rect 800 23835 840 23867
rect 872 23835 912 23867
rect 944 23835 984 23867
rect 1016 23835 1056 23867
rect 1088 23835 1128 23867
rect 1160 23835 1200 23867
rect 1232 23835 1272 23867
rect 1304 23835 1344 23867
rect 1376 23835 1416 23867
rect 1448 23835 1488 23867
rect 1520 23835 1560 23867
rect 1592 23835 1632 23867
rect 1664 23835 1704 23867
rect 1736 23835 1776 23867
rect 1808 23835 1848 23867
rect 1880 23835 2000 23867
rect 0 23795 2000 23835
rect 0 23763 120 23795
rect 152 23763 192 23795
rect 224 23763 264 23795
rect 296 23763 336 23795
rect 368 23763 408 23795
rect 440 23763 480 23795
rect 512 23763 552 23795
rect 584 23763 624 23795
rect 656 23763 696 23795
rect 728 23763 768 23795
rect 800 23763 840 23795
rect 872 23763 912 23795
rect 944 23763 984 23795
rect 1016 23763 1056 23795
rect 1088 23763 1128 23795
rect 1160 23763 1200 23795
rect 1232 23763 1272 23795
rect 1304 23763 1344 23795
rect 1376 23763 1416 23795
rect 1448 23763 1488 23795
rect 1520 23763 1560 23795
rect 1592 23763 1632 23795
rect 1664 23763 1704 23795
rect 1736 23763 1776 23795
rect 1808 23763 1848 23795
rect 1880 23763 2000 23795
rect 0 23723 2000 23763
rect 0 23691 120 23723
rect 152 23691 192 23723
rect 224 23691 264 23723
rect 296 23691 336 23723
rect 368 23691 408 23723
rect 440 23691 480 23723
rect 512 23691 552 23723
rect 584 23691 624 23723
rect 656 23691 696 23723
rect 728 23691 768 23723
rect 800 23691 840 23723
rect 872 23691 912 23723
rect 944 23691 984 23723
rect 1016 23691 1056 23723
rect 1088 23691 1128 23723
rect 1160 23691 1200 23723
rect 1232 23691 1272 23723
rect 1304 23691 1344 23723
rect 1376 23691 1416 23723
rect 1448 23691 1488 23723
rect 1520 23691 1560 23723
rect 1592 23691 1632 23723
rect 1664 23691 1704 23723
rect 1736 23691 1776 23723
rect 1808 23691 1848 23723
rect 1880 23691 2000 23723
rect 0 23651 2000 23691
rect 0 23619 120 23651
rect 152 23619 192 23651
rect 224 23619 264 23651
rect 296 23619 336 23651
rect 368 23619 408 23651
rect 440 23619 480 23651
rect 512 23619 552 23651
rect 584 23619 624 23651
rect 656 23619 696 23651
rect 728 23619 768 23651
rect 800 23619 840 23651
rect 872 23619 912 23651
rect 944 23619 984 23651
rect 1016 23619 1056 23651
rect 1088 23619 1128 23651
rect 1160 23619 1200 23651
rect 1232 23619 1272 23651
rect 1304 23619 1344 23651
rect 1376 23619 1416 23651
rect 1448 23619 1488 23651
rect 1520 23619 1560 23651
rect 1592 23619 1632 23651
rect 1664 23619 1704 23651
rect 1736 23619 1776 23651
rect 1808 23619 1848 23651
rect 1880 23619 2000 23651
rect 0 23579 2000 23619
rect 0 23547 120 23579
rect 152 23547 192 23579
rect 224 23547 264 23579
rect 296 23547 336 23579
rect 368 23547 408 23579
rect 440 23547 480 23579
rect 512 23547 552 23579
rect 584 23547 624 23579
rect 656 23547 696 23579
rect 728 23547 768 23579
rect 800 23547 840 23579
rect 872 23547 912 23579
rect 944 23547 984 23579
rect 1016 23547 1056 23579
rect 1088 23547 1128 23579
rect 1160 23547 1200 23579
rect 1232 23547 1272 23579
rect 1304 23547 1344 23579
rect 1376 23547 1416 23579
rect 1448 23547 1488 23579
rect 1520 23547 1560 23579
rect 1592 23547 1632 23579
rect 1664 23547 1704 23579
rect 1736 23547 1776 23579
rect 1808 23547 1848 23579
rect 1880 23547 2000 23579
rect 0 23507 2000 23547
rect 0 23475 120 23507
rect 152 23475 192 23507
rect 224 23475 264 23507
rect 296 23475 336 23507
rect 368 23475 408 23507
rect 440 23475 480 23507
rect 512 23475 552 23507
rect 584 23475 624 23507
rect 656 23475 696 23507
rect 728 23475 768 23507
rect 800 23475 840 23507
rect 872 23475 912 23507
rect 944 23475 984 23507
rect 1016 23475 1056 23507
rect 1088 23475 1128 23507
rect 1160 23475 1200 23507
rect 1232 23475 1272 23507
rect 1304 23475 1344 23507
rect 1376 23475 1416 23507
rect 1448 23475 1488 23507
rect 1520 23475 1560 23507
rect 1592 23475 1632 23507
rect 1664 23475 1704 23507
rect 1736 23475 1776 23507
rect 1808 23475 1848 23507
rect 1880 23475 2000 23507
rect 0 23435 2000 23475
rect 0 23403 120 23435
rect 152 23403 192 23435
rect 224 23403 264 23435
rect 296 23403 336 23435
rect 368 23403 408 23435
rect 440 23403 480 23435
rect 512 23403 552 23435
rect 584 23403 624 23435
rect 656 23403 696 23435
rect 728 23403 768 23435
rect 800 23403 840 23435
rect 872 23403 912 23435
rect 944 23403 984 23435
rect 1016 23403 1056 23435
rect 1088 23403 1128 23435
rect 1160 23403 1200 23435
rect 1232 23403 1272 23435
rect 1304 23403 1344 23435
rect 1376 23403 1416 23435
rect 1448 23403 1488 23435
rect 1520 23403 1560 23435
rect 1592 23403 1632 23435
rect 1664 23403 1704 23435
rect 1736 23403 1776 23435
rect 1808 23403 1848 23435
rect 1880 23403 2000 23435
rect 0 23363 2000 23403
rect 0 23331 120 23363
rect 152 23331 192 23363
rect 224 23331 264 23363
rect 296 23331 336 23363
rect 368 23331 408 23363
rect 440 23331 480 23363
rect 512 23331 552 23363
rect 584 23331 624 23363
rect 656 23331 696 23363
rect 728 23331 768 23363
rect 800 23331 840 23363
rect 872 23331 912 23363
rect 944 23331 984 23363
rect 1016 23331 1056 23363
rect 1088 23331 1128 23363
rect 1160 23331 1200 23363
rect 1232 23331 1272 23363
rect 1304 23331 1344 23363
rect 1376 23331 1416 23363
rect 1448 23331 1488 23363
rect 1520 23331 1560 23363
rect 1592 23331 1632 23363
rect 1664 23331 1704 23363
rect 1736 23331 1776 23363
rect 1808 23331 1848 23363
rect 1880 23331 2000 23363
rect 0 23291 2000 23331
rect 0 23259 120 23291
rect 152 23259 192 23291
rect 224 23259 264 23291
rect 296 23259 336 23291
rect 368 23259 408 23291
rect 440 23259 480 23291
rect 512 23259 552 23291
rect 584 23259 624 23291
rect 656 23259 696 23291
rect 728 23259 768 23291
rect 800 23259 840 23291
rect 872 23259 912 23291
rect 944 23259 984 23291
rect 1016 23259 1056 23291
rect 1088 23259 1128 23291
rect 1160 23259 1200 23291
rect 1232 23259 1272 23291
rect 1304 23259 1344 23291
rect 1376 23259 1416 23291
rect 1448 23259 1488 23291
rect 1520 23259 1560 23291
rect 1592 23259 1632 23291
rect 1664 23259 1704 23291
rect 1736 23259 1776 23291
rect 1808 23259 1848 23291
rect 1880 23259 2000 23291
rect 0 23219 2000 23259
rect 0 23187 120 23219
rect 152 23187 192 23219
rect 224 23187 264 23219
rect 296 23187 336 23219
rect 368 23187 408 23219
rect 440 23187 480 23219
rect 512 23187 552 23219
rect 584 23187 624 23219
rect 656 23187 696 23219
rect 728 23187 768 23219
rect 800 23187 840 23219
rect 872 23187 912 23219
rect 944 23187 984 23219
rect 1016 23187 1056 23219
rect 1088 23187 1128 23219
rect 1160 23187 1200 23219
rect 1232 23187 1272 23219
rect 1304 23187 1344 23219
rect 1376 23187 1416 23219
rect 1448 23187 1488 23219
rect 1520 23187 1560 23219
rect 1592 23187 1632 23219
rect 1664 23187 1704 23219
rect 1736 23187 1776 23219
rect 1808 23187 1848 23219
rect 1880 23187 2000 23219
rect 0 23124 2000 23187
rect 0 22874 2000 22924
rect 0 22842 120 22874
rect 152 22842 192 22874
rect 224 22842 264 22874
rect 296 22842 336 22874
rect 368 22842 408 22874
rect 440 22842 480 22874
rect 512 22842 552 22874
rect 584 22842 624 22874
rect 656 22842 696 22874
rect 728 22842 768 22874
rect 800 22842 840 22874
rect 872 22842 912 22874
rect 944 22842 984 22874
rect 1016 22842 1056 22874
rect 1088 22842 1128 22874
rect 1160 22842 1200 22874
rect 1232 22842 1272 22874
rect 1304 22842 1344 22874
rect 1376 22842 1416 22874
rect 1448 22842 1488 22874
rect 1520 22842 1560 22874
rect 1592 22842 1632 22874
rect 1664 22842 1704 22874
rect 1736 22842 1776 22874
rect 1808 22842 1848 22874
rect 1880 22842 2000 22874
rect 0 22802 2000 22842
rect 0 22770 120 22802
rect 152 22770 192 22802
rect 224 22770 264 22802
rect 296 22770 336 22802
rect 368 22770 408 22802
rect 440 22770 480 22802
rect 512 22770 552 22802
rect 584 22770 624 22802
rect 656 22770 696 22802
rect 728 22770 768 22802
rect 800 22770 840 22802
rect 872 22770 912 22802
rect 944 22770 984 22802
rect 1016 22770 1056 22802
rect 1088 22770 1128 22802
rect 1160 22770 1200 22802
rect 1232 22770 1272 22802
rect 1304 22770 1344 22802
rect 1376 22770 1416 22802
rect 1448 22770 1488 22802
rect 1520 22770 1560 22802
rect 1592 22770 1632 22802
rect 1664 22770 1704 22802
rect 1736 22770 1776 22802
rect 1808 22770 1848 22802
rect 1880 22770 2000 22802
rect 0 22730 2000 22770
rect 0 22698 120 22730
rect 152 22698 192 22730
rect 224 22698 264 22730
rect 296 22698 336 22730
rect 368 22698 408 22730
rect 440 22698 480 22730
rect 512 22698 552 22730
rect 584 22698 624 22730
rect 656 22698 696 22730
rect 728 22698 768 22730
rect 800 22698 840 22730
rect 872 22698 912 22730
rect 944 22698 984 22730
rect 1016 22698 1056 22730
rect 1088 22698 1128 22730
rect 1160 22698 1200 22730
rect 1232 22698 1272 22730
rect 1304 22698 1344 22730
rect 1376 22698 1416 22730
rect 1448 22698 1488 22730
rect 1520 22698 1560 22730
rect 1592 22698 1632 22730
rect 1664 22698 1704 22730
rect 1736 22698 1776 22730
rect 1808 22698 1848 22730
rect 1880 22698 2000 22730
rect 0 22658 2000 22698
rect 0 22626 120 22658
rect 152 22626 192 22658
rect 224 22626 264 22658
rect 296 22626 336 22658
rect 368 22626 408 22658
rect 440 22626 480 22658
rect 512 22626 552 22658
rect 584 22626 624 22658
rect 656 22626 696 22658
rect 728 22626 768 22658
rect 800 22626 840 22658
rect 872 22626 912 22658
rect 944 22626 984 22658
rect 1016 22626 1056 22658
rect 1088 22626 1128 22658
rect 1160 22626 1200 22658
rect 1232 22626 1272 22658
rect 1304 22626 1344 22658
rect 1376 22626 1416 22658
rect 1448 22626 1488 22658
rect 1520 22626 1560 22658
rect 1592 22626 1632 22658
rect 1664 22626 1704 22658
rect 1736 22626 1776 22658
rect 1808 22626 1848 22658
rect 1880 22626 2000 22658
rect 0 22586 2000 22626
rect 0 22554 120 22586
rect 152 22554 192 22586
rect 224 22554 264 22586
rect 296 22554 336 22586
rect 368 22554 408 22586
rect 440 22554 480 22586
rect 512 22554 552 22586
rect 584 22554 624 22586
rect 656 22554 696 22586
rect 728 22554 768 22586
rect 800 22554 840 22586
rect 872 22554 912 22586
rect 944 22554 984 22586
rect 1016 22554 1056 22586
rect 1088 22554 1128 22586
rect 1160 22554 1200 22586
rect 1232 22554 1272 22586
rect 1304 22554 1344 22586
rect 1376 22554 1416 22586
rect 1448 22554 1488 22586
rect 1520 22554 1560 22586
rect 1592 22554 1632 22586
rect 1664 22554 1704 22586
rect 1736 22554 1776 22586
rect 1808 22554 1848 22586
rect 1880 22554 2000 22586
rect 0 22514 2000 22554
rect 0 22482 120 22514
rect 152 22482 192 22514
rect 224 22482 264 22514
rect 296 22482 336 22514
rect 368 22482 408 22514
rect 440 22482 480 22514
rect 512 22482 552 22514
rect 584 22482 624 22514
rect 656 22482 696 22514
rect 728 22482 768 22514
rect 800 22482 840 22514
rect 872 22482 912 22514
rect 944 22482 984 22514
rect 1016 22482 1056 22514
rect 1088 22482 1128 22514
rect 1160 22482 1200 22514
rect 1232 22482 1272 22514
rect 1304 22482 1344 22514
rect 1376 22482 1416 22514
rect 1448 22482 1488 22514
rect 1520 22482 1560 22514
rect 1592 22482 1632 22514
rect 1664 22482 1704 22514
rect 1736 22482 1776 22514
rect 1808 22482 1848 22514
rect 1880 22482 2000 22514
rect 0 22442 2000 22482
rect 0 22410 120 22442
rect 152 22410 192 22442
rect 224 22410 264 22442
rect 296 22410 336 22442
rect 368 22410 408 22442
rect 440 22410 480 22442
rect 512 22410 552 22442
rect 584 22410 624 22442
rect 656 22410 696 22442
rect 728 22410 768 22442
rect 800 22410 840 22442
rect 872 22410 912 22442
rect 944 22410 984 22442
rect 1016 22410 1056 22442
rect 1088 22410 1128 22442
rect 1160 22410 1200 22442
rect 1232 22410 1272 22442
rect 1304 22410 1344 22442
rect 1376 22410 1416 22442
rect 1448 22410 1488 22442
rect 1520 22410 1560 22442
rect 1592 22410 1632 22442
rect 1664 22410 1704 22442
rect 1736 22410 1776 22442
rect 1808 22410 1848 22442
rect 1880 22410 2000 22442
rect 0 22370 2000 22410
rect 0 22338 120 22370
rect 152 22338 192 22370
rect 224 22338 264 22370
rect 296 22338 336 22370
rect 368 22338 408 22370
rect 440 22338 480 22370
rect 512 22338 552 22370
rect 584 22338 624 22370
rect 656 22338 696 22370
rect 728 22338 768 22370
rect 800 22338 840 22370
rect 872 22338 912 22370
rect 944 22338 984 22370
rect 1016 22338 1056 22370
rect 1088 22338 1128 22370
rect 1160 22338 1200 22370
rect 1232 22338 1272 22370
rect 1304 22338 1344 22370
rect 1376 22338 1416 22370
rect 1448 22338 1488 22370
rect 1520 22338 1560 22370
rect 1592 22338 1632 22370
rect 1664 22338 1704 22370
rect 1736 22338 1776 22370
rect 1808 22338 1848 22370
rect 1880 22338 2000 22370
rect 0 22298 2000 22338
rect 0 22266 120 22298
rect 152 22266 192 22298
rect 224 22266 264 22298
rect 296 22266 336 22298
rect 368 22266 408 22298
rect 440 22266 480 22298
rect 512 22266 552 22298
rect 584 22266 624 22298
rect 656 22266 696 22298
rect 728 22266 768 22298
rect 800 22266 840 22298
rect 872 22266 912 22298
rect 944 22266 984 22298
rect 1016 22266 1056 22298
rect 1088 22266 1128 22298
rect 1160 22266 1200 22298
rect 1232 22266 1272 22298
rect 1304 22266 1344 22298
rect 1376 22266 1416 22298
rect 1448 22266 1488 22298
rect 1520 22266 1560 22298
rect 1592 22266 1632 22298
rect 1664 22266 1704 22298
rect 1736 22266 1776 22298
rect 1808 22266 1848 22298
rect 1880 22266 2000 22298
rect 0 22226 2000 22266
rect 0 22194 120 22226
rect 152 22194 192 22226
rect 224 22194 264 22226
rect 296 22194 336 22226
rect 368 22194 408 22226
rect 440 22194 480 22226
rect 512 22194 552 22226
rect 584 22194 624 22226
rect 656 22194 696 22226
rect 728 22194 768 22226
rect 800 22194 840 22226
rect 872 22194 912 22226
rect 944 22194 984 22226
rect 1016 22194 1056 22226
rect 1088 22194 1128 22226
rect 1160 22194 1200 22226
rect 1232 22194 1272 22226
rect 1304 22194 1344 22226
rect 1376 22194 1416 22226
rect 1448 22194 1488 22226
rect 1520 22194 1560 22226
rect 1592 22194 1632 22226
rect 1664 22194 1704 22226
rect 1736 22194 1776 22226
rect 1808 22194 1848 22226
rect 1880 22194 2000 22226
rect 0 22154 2000 22194
rect 0 22122 120 22154
rect 152 22122 192 22154
rect 224 22122 264 22154
rect 296 22122 336 22154
rect 368 22122 408 22154
rect 440 22122 480 22154
rect 512 22122 552 22154
rect 584 22122 624 22154
rect 656 22122 696 22154
rect 728 22122 768 22154
rect 800 22122 840 22154
rect 872 22122 912 22154
rect 944 22122 984 22154
rect 1016 22122 1056 22154
rect 1088 22122 1128 22154
rect 1160 22122 1200 22154
rect 1232 22122 1272 22154
rect 1304 22122 1344 22154
rect 1376 22122 1416 22154
rect 1448 22122 1488 22154
rect 1520 22122 1560 22154
rect 1592 22122 1632 22154
rect 1664 22122 1704 22154
rect 1736 22122 1776 22154
rect 1808 22122 1848 22154
rect 1880 22122 2000 22154
rect 0 22082 2000 22122
rect 0 22050 120 22082
rect 152 22050 192 22082
rect 224 22050 264 22082
rect 296 22050 336 22082
rect 368 22050 408 22082
rect 440 22050 480 22082
rect 512 22050 552 22082
rect 584 22050 624 22082
rect 656 22050 696 22082
rect 728 22050 768 22082
rect 800 22050 840 22082
rect 872 22050 912 22082
rect 944 22050 984 22082
rect 1016 22050 1056 22082
rect 1088 22050 1128 22082
rect 1160 22050 1200 22082
rect 1232 22050 1272 22082
rect 1304 22050 1344 22082
rect 1376 22050 1416 22082
rect 1448 22050 1488 22082
rect 1520 22050 1560 22082
rect 1592 22050 1632 22082
rect 1664 22050 1704 22082
rect 1736 22050 1776 22082
rect 1808 22050 1848 22082
rect 1880 22050 2000 22082
rect 0 22010 2000 22050
rect 0 21978 120 22010
rect 152 21978 192 22010
rect 224 21978 264 22010
rect 296 21978 336 22010
rect 368 21978 408 22010
rect 440 21978 480 22010
rect 512 21978 552 22010
rect 584 21978 624 22010
rect 656 21978 696 22010
rect 728 21978 768 22010
rect 800 21978 840 22010
rect 872 21978 912 22010
rect 944 21978 984 22010
rect 1016 21978 1056 22010
rect 1088 21978 1128 22010
rect 1160 21978 1200 22010
rect 1232 21978 1272 22010
rect 1304 21978 1344 22010
rect 1376 21978 1416 22010
rect 1448 21978 1488 22010
rect 1520 21978 1560 22010
rect 1592 21978 1632 22010
rect 1664 21978 1704 22010
rect 1736 21978 1776 22010
rect 1808 21978 1848 22010
rect 1880 21978 2000 22010
rect 0 21938 2000 21978
rect 0 21906 120 21938
rect 152 21906 192 21938
rect 224 21906 264 21938
rect 296 21906 336 21938
rect 368 21906 408 21938
rect 440 21906 480 21938
rect 512 21906 552 21938
rect 584 21906 624 21938
rect 656 21906 696 21938
rect 728 21906 768 21938
rect 800 21906 840 21938
rect 872 21906 912 21938
rect 944 21906 984 21938
rect 1016 21906 1056 21938
rect 1088 21906 1128 21938
rect 1160 21906 1200 21938
rect 1232 21906 1272 21938
rect 1304 21906 1344 21938
rect 1376 21906 1416 21938
rect 1448 21906 1488 21938
rect 1520 21906 1560 21938
rect 1592 21906 1632 21938
rect 1664 21906 1704 21938
rect 1736 21906 1776 21938
rect 1808 21906 1848 21938
rect 1880 21906 2000 21938
rect 0 21866 2000 21906
rect 0 21834 120 21866
rect 152 21834 192 21866
rect 224 21834 264 21866
rect 296 21834 336 21866
rect 368 21834 408 21866
rect 440 21834 480 21866
rect 512 21834 552 21866
rect 584 21834 624 21866
rect 656 21834 696 21866
rect 728 21834 768 21866
rect 800 21834 840 21866
rect 872 21834 912 21866
rect 944 21834 984 21866
rect 1016 21834 1056 21866
rect 1088 21834 1128 21866
rect 1160 21834 1200 21866
rect 1232 21834 1272 21866
rect 1304 21834 1344 21866
rect 1376 21834 1416 21866
rect 1448 21834 1488 21866
rect 1520 21834 1560 21866
rect 1592 21834 1632 21866
rect 1664 21834 1704 21866
rect 1736 21834 1776 21866
rect 1808 21834 1848 21866
rect 1880 21834 2000 21866
rect 0 21794 2000 21834
rect 0 21762 120 21794
rect 152 21762 192 21794
rect 224 21762 264 21794
rect 296 21762 336 21794
rect 368 21762 408 21794
rect 440 21762 480 21794
rect 512 21762 552 21794
rect 584 21762 624 21794
rect 656 21762 696 21794
rect 728 21762 768 21794
rect 800 21762 840 21794
rect 872 21762 912 21794
rect 944 21762 984 21794
rect 1016 21762 1056 21794
rect 1088 21762 1128 21794
rect 1160 21762 1200 21794
rect 1232 21762 1272 21794
rect 1304 21762 1344 21794
rect 1376 21762 1416 21794
rect 1448 21762 1488 21794
rect 1520 21762 1560 21794
rect 1592 21762 1632 21794
rect 1664 21762 1704 21794
rect 1736 21762 1776 21794
rect 1808 21762 1848 21794
rect 1880 21762 2000 21794
rect 0 21722 2000 21762
rect 0 21690 120 21722
rect 152 21690 192 21722
rect 224 21690 264 21722
rect 296 21690 336 21722
rect 368 21690 408 21722
rect 440 21690 480 21722
rect 512 21690 552 21722
rect 584 21690 624 21722
rect 656 21690 696 21722
rect 728 21690 768 21722
rect 800 21690 840 21722
rect 872 21690 912 21722
rect 944 21690 984 21722
rect 1016 21690 1056 21722
rect 1088 21690 1128 21722
rect 1160 21690 1200 21722
rect 1232 21690 1272 21722
rect 1304 21690 1344 21722
rect 1376 21690 1416 21722
rect 1448 21690 1488 21722
rect 1520 21690 1560 21722
rect 1592 21690 1632 21722
rect 1664 21690 1704 21722
rect 1736 21690 1776 21722
rect 1808 21690 1848 21722
rect 1880 21690 2000 21722
rect 0 21650 2000 21690
rect 0 21618 120 21650
rect 152 21618 192 21650
rect 224 21618 264 21650
rect 296 21618 336 21650
rect 368 21618 408 21650
rect 440 21618 480 21650
rect 512 21618 552 21650
rect 584 21618 624 21650
rect 656 21618 696 21650
rect 728 21618 768 21650
rect 800 21618 840 21650
rect 872 21618 912 21650
rect 944 21618 984 21650
rect 1016 21618 1056 21650
rect 1088 21618 1128 21650
rect 1160 21618 1200 21650
rect 1232 21618 1272 21650
rect 1304 21618 1344 21650
rect 1376 21618 1416 21650
rect 1448 21618 1488 21650
rect 1520 21618 1560 21650
rect 1592 21618 1632 21650
rect 1664 21618 1704 21650
rect 1736 21618 1776 21650
rect 1808 21618 1848 21650
rect 1880 21618 2000 21650
rect 0 21578 2000 21618
rect 0 21546 120 21578
rect 152 21546 192 21578
rect 224 21546 264 21578
rect 296 21546 336 21578
rect 368 21546 408 21578
rect 440 21546 480 21578
rect 512 21546 552 21578
rect 584 21546 624 21578
rect 656 21546 696 21578
rect 728 21546 768 21578
rect 800 21546 840 21578
rect 872 21546 912 21578
rect 944 21546 984 21578
rect 1016 21546 1056 21578
rect 1088 21546 1128 21578
rect 1160 21546 1200 21578
rect 1232 21546 1272 21578
rect 1304 21546 1344 21578
rect 1376 21546 1416 21578
rect 1448 21546 1488 21578
rect 1520 21546 1560 21578
rect 1592 21546 1632 21578
rect 1664 21546 1704 21578
rect 1736 21546 1776 21578
rect 1808 21546 1848 21578
rect 1880 21546 2000 21578
rect 0 21506 2000 21546
rect 0 21474 120 21506
rect 152 21474 192 21506
rect 224 21474 264 21506
rect 296 21474 336 21506
rect 368 21474 408 21506
rect 440 21474 480 21506
rect 512 21474 552 21506
rect 584 21474 624 21506
rect 656 21474 696 21506
rect 728 21474 768 21506
rect 800 21474 840 21506
rect 872 21474 912 21506
rect 944 21474 984 21506
rect 1016 21474 1056 21506
rect 1088 21474 1128 21506
rect 1160 21474 1200 21506
rect 1232 21474 1272 21506
rect 1304 21474 1344 21506
rect 1376 21474 1416 21506
rect 1448 21474 1488 21506
rect 1520 21474 1560 21506
rect 1592 21474 1632 21506
rect 1664 21474 1704 21506
rect 1736 21474 1776 21506
rect 1808 21474 1848 21506
rect 1880 21474 2000 21506
rect 0 21434 2000 21474
rect 0 21402 120 21434
rect 152 21402 192 21434
rect 224 21402 264 21434
rect 296 21402 336 21434
rect 368 21402 408 21434
rect 440 21402 480 21434
rect 512 21402 552 21434
rect 584 21402 624 21434
rect 656 21402 696 21434
rect 728 21402 768 21434
rect 800 21402 840 21434
rect 872 21402 912 21434
rect 944 21402 984 21434
rect 1016 21402 1056 21434
rect 1088 21402 1128 21434
rect 1160 21402 1200 21434
rect 1232 21402 1272 21434
rect 1304 21402 1344 21434
rect 1376 21402 1416 21434
rect 1448 21402 1488 21434
rect 1520 21402 1560 21434
rect 1592 21402 1632 21434
rect 1664 21402 1704 21434
rect 1736 21402 1776 21434
rect 1808 21402 1848 21434
rect 1880 21402 2000 21434
rect 0 21362 2000 21402
rect 0 21330 120 21362
rect 152 21330 192 21362
rect 224 21330 264 21362
rect 296 21330 336 21362
rect 368 21330 408 21362
rect 440 21330 480 21362
rect 512 21330 552 21362
rect 584 21330 624 21362
rect 656 21330 696 21362
rect 728 21330 768 21362
rect 800 21330 840 21362
rect 872 21330 912 21362
rect 944 21330 984 21362
rect 1016 21330 1056 21362
rect 1088 21330 1128 21362
rect 1160 21330 1200 21362
rect 1232 21330 1272 21362
rect 1304 21330 1344 21362
rect 1376 21330 1416 21362
rect 1448 21330 1488 21362
rect 1520 21330 1560 21362
rect 1592 21330 1632 21362
rect 1664 21330 1704 21362
rect 1736 21330 1776 21362
rect 1808 21330 1848 21362
rect 1880 21330 2000 21362
rect 0 21290 2000 21330
rect 0 21258 120 21290
rect 152 21258 192 21290
rect 224 21258 264 21290
rect 296 21258 336 21290
rect 368 21258 408 21290
rect 440 21258 480 21290
rect 512 21258 552 21290
rect 584 21258 624 21290
rect 656 21258 696 21290
rect 728 21258 768 21290
rect 800 21258 840 21290
rect 872 21258 912 21290
rect 944 21258 984 21290
rect 1016 21258 1056 21290
rect 1088 21258 1128 21290
rect 1160 21258 1200 21290
rect 1232 21258 1272 21290
rect 1304 21258 1344 21290
rect 1376 21258 1416 21290
rect 1448 21258 1488 21290
rect 1520 21258 1560 21290
rect 1592 21258 1632 21290
rect 1664 21258 1704 21290
rect 1736 21258 1776 21290
rect 1808 21258 1848 21290
rect 1880 21258 2000 21290
rect 0 21218 2000 21258
rect 0 21186 120 21218
rect 152 21186 192 21218
rect 224 21186 264 21218
rect 296 21186 336 21218
rect 368 21186 408 21218
rect 440 21186 480 21218
rect 512 21186 552 21218
rect 584 21186 624 21218
rect 656 21186 696 21218
rect 728 21186 768 21218
rect 800 21186 840 21218
rect 872 21186 912 21218
rect 944 21186 984 21218
rect 1016 21186 1056 21218
rect 1088 21186 1128 21218
rect 1160 21186 1200 21218
rect 1232 21186 1272 21218
rect 1304 21186 1344 21218
rect 1376 21186 1416 21218
rect 1448 21186 1488 21218
rect 1520 21186 1560 21218
rect 1592 21186 1632 21218
rect 1664 21186 1704 21218
rect 1736 21186 1776 21218
rect 1808 21186 1848 21218
rect 1880 21186 2000 21218
rect 0 21146 2000 21186
rect 0 21114 120 21146
rect 152 21114 192 21146
rect 224 21114 264 21146
rect 296 21114 336 21146
rect 368 21114 408 21146
rect 440 21114 480 21146
rect 512 21114 552 21146
rect 584 21114 624 21146
rect 656 21114 696 21146
rect 728 21114 768 21146
rect 800 21114 840 21146
rect 872 21114 912 21146
rect 944 21114 984 21146
rect 1016 21114 1056 21146
rect 1088 21114 1128 21146
rect 1160 21114 1200 21146
rect 1232 21114 1272 21146
rect 1304 21114 1344 21146
rect 1376 21114 1416 21146
rect 1448 21114 1488 21146
rect 1520 21114 1560 21146
rect 1592 21114 1632 21146
rect 1664 21114 1704 21146
rect 1736 21114 1776 21146
rect 1808 21114 1848 21146
rect 1880 21114 2000 21146
rect 0 21074 2000 21114
rect 0 21042 120 21074
rect 152 21042 192 21074
rect 224 21042 264 21074
rect 296 21042 336 21074
rect 368 21042 408 21074
rect 440 21042 480 21074
rect 512 21042 552 21074
rect 584 21042 624 21074
rect 656 21042 696 21074
rect 728 21042 768 21074
rect 800 21042 840 21074
rect 872 21042 912 21074
rect 944 21042 984 21074
rect 1016 21042 1056 21074
rect 1088 21042 1128 21074
rect 1160 21042 1200 21074
rect 1232 21042 1272 21074
rect 1304 21042 1344 21074
rect 1376 21042 1416 21074
rect 1448 21042 1488 21074
rect 1520 21042 1560 21074
rect 1592 21042 1632 21074
rect 1664 21042 1704 21074
rect 1736 21042 1776 21074
rect 1808 21042 1848 21074
rect 1880 21042 2000 21074
rect 0 21002 2000 21042
rect 0 20970 120 21002
rect 152 20970 192 21002
rect 224 20970 264 21002
rect 296 20970 336 21002
rect 368 20970 408 21002
rect 440 20970 480 21002
rect 512 20970 552 21002
rect 584 20970 624 21002
rect 656 20970 696 21002
rect 728 20970 768 21002
rect 800 20970 840 21002
rect 872 20970 912 21002
rect 944 20970 984 21002
rect 1016 20970 1056 21002
rect 1088 20970 1128 21002
rect 1160 20970 1200 21002
rect 1232 20970 1272 21002
rect 1304 20970 1344 21002
rect 1376 20970 1416 21002
rect 1448 20970 1488 21002
rect 1520 20970 1560 21002
rect 1592 20970 1632 21002
rect 1664 20970 1704 21002
rect 1736 20970 1776 21002
rect 1808 20970 1848 21002
rect 1880 20970 2000 21002
rect 0 20930 2000 20970
rect 0 20898 120 20930
rect 152 20898 192 20930
rect 224 20898 264 20930
rect 296 20898 336 20930
rect 368 20898 408 20930
rect 440 20898 480 20930
rect 512 20898 552 20930
rect 584 20898 624 20930
rect 656 20898 696 20930
rect 728 20898 768 20930
rect 800 20898 840 20930
rect 872 20898 912 20930
rect 944 20898 984 20930
rect 1016 20898 1056 20930
rect 1088 20898 1128 20930
rect 1160 20898 1200 20930
rect 1232 20898 1272 20930
rect 1304 20898 1344 20930
rect 1376 20898 1416 20930
rect 1448 20898 1488 20930
rect 1520 20898 1560 20930
rect 1592 20898 1632 20930
rect 1664 20898 1704 20930
rect 1736 20898 1776 20930
rect 1808 20898 1848 20930
rect 1880 20898 2000 20930
rect 0 20858 2000 20898
rect 0 20826 120 20858
rect 152 20826 192 20858
rect 224 20826 264 20858
rect 296 20826 336 20858
rect 368 20826 408 20858
rect 440 20826 480 20858
rect 512 20826 552 20858
rect 584 20826 624 20858
rect 656 20826 696 20858
rect 728 20826 768 20858
rect 800 20826 840 20858
rect 872 20826 912 20858
rect 944 20826 984 20858
rect 1016 20826 1056 20858
rect 1088 20826 1128 20858
rect 1160 20826 1200 20858
rect 1232 20826 1272 20858
rect 1304 20826 1344 20858
rect 1376 20826 1416 20858
rect 1448 20826 1488 20858
rect 1520 20826 1560 20858
rect 1592 20826 1632 20858
rect 1664 20826 1704 20858
rect 1736 20826 1776 20858
rect 1808 20826 1848 20858
rect 1880 20826 2000 20858
rect 0 20786 2000 20826
rect 0 20754 120 20786
rect 152 20754 192 20786
rect 224 20754 264 20786
rect 296 20754 336 20786
rect 368 20754 408 20786
rect 440 20754 480 20786
rect 512 20754 552 20786
rect 584 20754 624 20786
rect 656 20754 696 20786
rect 728 20754 768 20786
rect 800 20754 840 20786
rect 872 20754 912 20786
rect 944 20754 984 20786
rect 1016 20754 1056 20786
rect 1088 20754 1128 20786
rect 1160 20754 1200 20786
rect 1232 20754 1272 20786
rect 1304 20754 1344 20786
rect 1376 20754 1416 20786
rect 1448 20754 1488 20786
rect 1520 20754 1560 20786
rect 1592 20754 1632 20786
rect 1664 20754 1704 20786
rect 1736 20754 1776 20786
rect 1808 20754 1848 20786
rect 1880 20754 2000 20786
rect 0 20714 2000 20754
rect 0 20682 120 20714
rect 152 20682 192 20714
rect 224 20682 264 20714
rect 296 20682 336 20714
rect 368 20682 408 20714
rect 440 20682 480 20714
rect 512 20682 552 20714
rect 584 20682 624 20714
rect 656 20682 696 20714
rect 728 20682 768 20714
rect 800 20682 840 20714
rect 872 20682 912 20714
rect 944 20682 984 20714
rect 1016 20682 1056 20714
rect 1088 20682 1128 20714
rect 1160 20682 1200 20714
rect 1232 20682 1272 20714
rect 1304 20682 1344 20714
rect 1376 20682 1416 20714
rect 1448 20682 1488 20714
rect 1520 20682 1560 20714
rect 1592 20682 1632 20714
rect 1664 20682 1704 20714
rect 1736 20682 1776 20714
rect 1808 20682 1848 20714
rect 1880 20682 2000 20714
rect 0 20642 2000 20682
rect 0 20610 120 20642
rect 152 20610 192 20642
rect 224 20610 264 20642
rect 296 20610 336 20642
rect 368 20610 408 20642
rect 440 20610 480 20642
rect 512 20610 552 20642
rect 584 20610 624 20642
rect 656 20610 696 20642
rect 728 20610 768 20642
rect 800 20610 840 20642
rect 872 20610 912 20642
rect 944 20610 984 20642
rect 1016 20610 1056 20642
rect 1088 20610 1128 20642
rect 1160 20610 1200 20642
rect 1232 20610 1272 20642
rect 1304 20610 1344 20642
rect 1376 20610 1416 20642
rect 1448 20610 1488 20642
rect 1520 20610 1560 20642
rect 1592 20610 1632 20642
rect 1664 20610 1704 20642
rect 1736 20610 1776 20642
rect 1808 20610 1848 20642
rect 1880 20610 2000 20642
rect 0 20570 2000 20610
rect 0 20538 120 20570
rect 152 20538 192 20570
rect 224 20538 264 20570
rect 296 20538 336 20570
rect 368 20538 408 20570
rect 440 20538 480 20570
rect 512 20538 552 20570
rect 584 20538 624 20570
rect 656 20538 696 20570
rect 728 20538 768 20570
rect 800 20538 840 20570
rect 872 20538 912 20570
rect 944 20538 984 20570
rect 1016 20538 1056 20570
rect 1088 20538 1128 20570
rect 1160 20538 1200 20570
rect 1232 20538 1272 20570
rect 1304 20538 1344 20570
rect 1376 20538 1416 20570
rect 1448 20538 1488 20570
rect 1520 20538 1560 20570
rect 1592 20538 1632 20570
rect 1664 20538 1704 20570
rect 1736 20538 1776 20570
rect 1808 20538 1848 20570
rect 1880 20538 2000 20570
rect 0 20498 2000 20538
rect 0 20466 120 20498
rect 152 20466 192 20498
rect 224 20466 264 20498
rect 296 20466 336 20498
rect 368 20466 408 20498
rect 440 20466 480 20498
rect 512 20466 552 20498
rect 584 20466 624 20498
rect 656 20466 696 20498
rect 728 20466 768 20498
rect 800 20466 840 20498
rect 872 20466 912 20498
rect 944 20466 984 20498
rect 1016 20466 1056 20498
rect 1088 20466 1128 20498
rect 1160 20466 1200 20498
rect 1232 20466 1272 20498
rect 1304 20466 1344 20498
rect 1376 20466 1416 20498
rect 1448 20466 1488 20498
rect 1520 20466 1560 20498
rect 1592 20466 1632 20498
rect 1664 20466 1704 20498
rect 1736 20466 1776 20498
rect 1808 20466 1848 20498
rect 1880 20466 2000 20498
rect 0 20426 2000 20466
rect 0 20394 120 20426
rect 152 20394 192 20426
rect 224 20394 264 20426
rect 296 20394 336 20426
rect 368 20394 408 20426
rect 440 20394 480 20426
rect 512 20394 552 20426
rect 584 20394 624 20426
rect 656 20394 696 20426
rect 728 20394 768 20426
rect 800 20394 840 20426
rect 872 20394 912 20426
rect 944 20394 984 20426
rect 1016 20394 1056 20426
rect 1088 20394 1128 20426
rect 1160 20394 1200 20426
rect 1232 20394 1272 20426
rect 1304 20394 1344 20426
rect 1376 20394 1416 20426
rect 1448 20394 1488 20426
rect 1520 20394 1560 20426
rect 1592 20394 1632 20426
rect 1664 20394 1704 20426
rect 1736 20394 1776 20426
rect 1808 20394 1848 20426
rect 1880 20394 2000 20426
rect 0 20354 2000 20394
rect 0 20322 120 20354
rect 152 20322 192 20354
rect 224 20322 264 20354
rect 296 20322 336 20354
rect 368 20322 408 20354
rect 440 20322 480 20354
rect 512 20322 552 20354
rect 584 20322 624 20354
rect 656 20322 696 20354
rect 728 20322 768 20354
rect 800 20322 840 20354
rect 872 20322 912 20354
rect 944 20322 984 20354
rect 1016 20322 1056 20354
rect 1088 20322 1128 20354
rect 1160 20322 1200 20354
rect 1232 20322 1272 20354
rect 1304 20322 1344 20354
rect 1376 20322 1416 20354
rect 1448 20322 1488 20354
rect 1520 20322 1560 20354
rect 1592 20322 1632 20354
rect 1664 20322 1704 20354
rect 1736 20322 1776 20354
rect 1808 20322 1848 20354
rect 1880 20322 2000 20354
rect 0 20282 2000 20322
rect 0 20250 120 20282
rect 152 20250 192 20282
rect 224 20250 264 20282
rect 296 20250 336 20282
rect 368 20250 408 20282
rect 440 20250 480 20282
rect 512 20250 552 20282
rect 584 20250 624 20282
rect 656 20250 696 20282
rect 728 20250 768 20282
rect 800 20250 840 20282
rect 872 20250 912 20282
rect 944 20250 984 20282
rect 1016 20250 1056 20282
rect 1088 20250 1128 20282
rect 1160 20250 1200 20282
rect 1232 20250 1272 20282
rect 1304 20250 1344 20282
rect 1376 20250 1416 20282
rect 1448 20250 1488 20282
rect 1520 20250 1560 20282
rect 1592 20250 1632 20282
rect 1664 20250 1704 20282
rect 1736 20250 1776 20282
rect 1808 20250 1848 20282
rect 1880 20250 2000 20282
rect 0 20210 2000 20250
rect 0 20178 120 20210
rect 152 20178 192 20210
rect 224 20178 264 20210
rect 296 20178 336 20210
rect 368 20178 408 20210
rect 440 20178 480 20210
rect 512 20178 552 20210
rect 584 20178 624 20210
rect 656 20178 696 20210
rect 728 20178 768 20210
rect 800 20178 840 20210
rect 872 20178 912 20210
rect 944 20178 984 20210
rect 1016 20178 1056 20210
rect 1088 20178 1128 20210
rect 1160 20178 1200 20210
rect 1232 20178 1272 20210
rect 1304 20178 1344 20210
rect 1376 20178 1416 20210
rect 1448 20178 1488 20210
rect 1520 20178 1560 20210
rect 1592 20178 1632 20210
rect 1664 20178 1704 20210
rect 1736 20178 1776 20210
rect 1808 20178 1848 20210
rect 1880 20178 2000 20210
rect 0 20138 2000 20178
rect 0 20106 120 20138
rect 152 20106 192 20138
rect 224 20106 264 20138
rect 296 20106 336 20138
rect 368 20106 408 20138
rect 440 20106 480 20138
rect 512 20106 552 20138
rect 584 20106 624 20138
rect 656 20106 696 20138
rect 728 20106 768 20138
rect 800 20106 840 20138
rect 872 20106 912 20138
rect 944 20106 984 20138
rect 1016 20106 1056 20138
rect 1088 20106 1128 20138
rect 1160 20106 1200 20138
rect 1232 20106 1272 20138
rect 1304 20106 1344 20138
rect 1376 20106 1416 20138
rect 1448 20106 1488 20138
rect 1520 20106 1560 20138
rect 1592 20106 1632 20138
rect 1664 20106 1704 20138
rect 1736 20106 1776 20138
rect 1808 20106 1848 20138
rect 1880 20106 2000 20138
rect 0 20066 2000 20106
rect 0 20034 120 20066
rect 152 20034 192 20066
rect 224 20034 264 20066
rect 296 20034 336 20066
rect 368 20034 408 20066
rect 440 20034 480 20066
rect 512 20034 552 20066
rect 584 20034 624 20066
rect 656 20034 696 20066
rect 728 20034 768 20066
rect 800 20034 840 20066
rect 872 20034 912 20066
rect 944 20034 984 20066
rect 1016 20034 1056 20066
rect 1088 20034 1128 20066
rect 1160 20034 1200 20066
rect 1232 20034 1272 20066
rect 1304 20034 1344 20066
rect 1376 20034 1416 20066
rect 1448 20034 1488 20066
rect 1520 20034 1560 20066
rect 1592 20034 1632 20066
rect 1664 20034 1704 20066
rect 1736 20034 1776 20066
rect 1808 20034 1848 20066
rect 1880 20034 2000 20066
rect 0 19994 2000 20034
rect 0 19962 120 19994
rect 152 19962 192 19994
rect 224 19962 264 19994
rect 296 19962 336 19994
rect 368 19962 408 19994
rect 440 19962 480 19994
rect 512 19962 552 19994
rect 584 19962 624 19994
rect 656 19962 696 19994
rect 728 19962 768 19994
rect 800 19962 840 19994
rect 872 19962 912 19994
rect 944 19962 984 19994
rect 1016 19962 1056 19994
rect 1088 19962 1128 19994
rect 1160 19962 1200 19994
rect 1232 19962 1272 19994
rect 1304 19962 1344 19994
rect 1376 19962 1416 19994
rect 1448 19962 1488 19994
rect 1520 19962 1560 19994
rect 1592 19962 1632 19994
rect 1664 19962 1704 19994
rect 1736 19962 1776 19994
rect 1808 19962 1848 19994
rect 1880 19962 2000 19994
rect 0 19922 2000 19962
rect 0 19890 120 19922
rect 152 19890 192 19922
rect 224 19890 264 19922
rect 296 19890 336 19922
rect 368 19890 408 19922
rect 440 19890 480 19922
rect 512 19890 552 19922
rect 584 19890 624 19922
rect 656 19890 696 19922
rect 728 19890 768 19922
rect 800 19890 840 19922
rect 872 19890 912 19922
rect 944 19890 984 19922
rect 1016 19890 1056 19922
rect 1088 19890 1128 19922
rect 1160 19890 1200 19922
rect 1232 19890 1272 19922
rect 1304 19890 1344 19922
rect 1376 19890 1416 19922
rect 1448 19890 1488 19922
rect 1520 19890 1560 19922
rect 1592 19890 1632 19922
rect 1664 19890 1704 19922
rect 1736 19890 1776 19922
rect 1808 19890 1848 19922
rect 1880 19890 2000 19922
rect 0 19850 2000 19890
rect 0 19818 120 19850
rect 152 19818 192 19850
rect 224 19818 264 19850
rect 296 19818 336 19850
rect 368 19818 408 19850
rect 440 19818 480 19850
rect 512 19818 552 19850
rect 584 19818 624 19850
rect 656 19818 696 19850
rect 728 19818 768 19850
rect 800 19818 840 19850
rect 872 19818 912 19850
rect 944 19818 984 19850
rect 1016 19818 1056 19850
rect 1088 19818 1128 19850
rect 1160 19818 1200 19850
rect 1232 19818 1272 19850
rect 1304 19818 1344 19850
rect 1376 19818 1416 19850
rect 1448 19818 1488 19850
rect 1520 19818 1560 19850
rect 1592 19818 1632 19850
rect 1664 19818 1704 19850
rect 1736 19818 1776 19850
rect 1808 19818 1848 19850
rect 1880 19818 2000 19850
rect 0 19778 2000 19818
rect 0 19746 120 19778
rect 152 19746 192 19778
rect 224 19746 264 19778
rect 296 19746 336 19778
rect 368 19746 408 19778
rect 440 19746 480 19778
rect 512 19746 552 19778
rect 584 19746 624 19778
rect 656 19746 696 19778
rect 728 19746 768 19778
rect 800 19746 840 19778
rect 872 19746 912 19778
rect 944 19746 984 19778
rect 1016 19746 1056 19778
rect 1088 19746 1128 19778
rect 1160 19746 1200 19778
rect 1232 19746 1272 19778
rect 1304 19746 1344 19778
rect 1376 19746 1416 19778
rect 1448 19746 1488 19778
rect 1520 19746 1560 19778
rect 1592 19746 1632 19778
rect 1664 19746 1704 19778
rect 1736 19746 1776 19778
rect 1808 19746 1848 19778
rect 1880 19746 2000 19778
rect 0 19706 2000 19746
rect 0 19674 120 19706
rect 152 19674 192 19706
rect 224 19674 264 19706
rect 296 19674 336 19706
rect 368 19674 408 19706
rect 440 19674 480 19706
rect 512 19674 552 19706
rect 584 19674 624 19706
rect 656 19674 696 19706
rect 728 19674 768 19706
rect 800 19674 840 19706
rect 872 19674 912 19706
rect 944 19674 984 19706
rect 1016 19674 1056 19706
rect 1088 19674 1128 19706
rect 1160 19674 1200 19706
rect 1232 19674 1272 19706
rect 1304 19674 1344 19706
rect 1376 19674 1416 19706
rect 1448 19674 1488 19706
rect 1520 19674 1560 19706
rect 1592 19674 1632 19706
rect 1664 19674 1704 19706
rect 1736 19674 1776 19706
rect 1808 19674 1848 19706
rect 1880 19674 2000 19706
rect 0 19634 2000 19674
rect 0 19602 120 19634
rect 152 19602 192 19634
rect 224 19602 264 19634
rect 296 19602 336 19634
rect 368 19602 408 19634
rect 440 19602 480 19634
rect 512 19602 552 19634
rect 584 19602 624 19634
rect 656 19602 696 19634
rect 728 19602 768 19634
rect 800 19602 840 19634
rect 872 19602 912 19634
rect 944 19602 984 19634
rect 1016 19602 1056 19634
rect 1088 19602 1128 19634
rect 1160 19602 1200 19634
rect 1232 19602 1272 19634
rect 1304 19602 1344 19634
rect 1376 19602 1416 19634
rect 1448 19602 1488 19634
rect 1520 19602 1560 19634
rect 1592 19602 1632 19634
rect 1664 19602 1704 19634
rect 1736 19602 1776 19634
rect 1808 19602 1848 19634
rect 1880 19602 2000 19634
rect 0 19562 2000 19602
rect 0 19530 120 19562
rect 152 19530 192 19562
rect 224 19530 264 19562
rect 296 19530 336 19562
rect 368 19530 408 19562
rect 440 19530 480 19562
rect 512 19530 552 19562
rect 584 19530 624 19562
rect 656 19530 696 19562
rect 728 19530 768 19562
rect 800 19530 840 19562
rect 872 19530 912 19562
rect 944 19530 984 19562
rect 1016 19530 1056 19562
rect 1088 19530 1128 19562
rect 1160 19530 1200 19562
rect 1232 19530 1272 19562
rect 1304 19530 1344 19562
rect 1376 19530 1416 19562
rect 1448 19530 1488 19562
rect 1520 19530 1560 19562
rect 1592 19530 1632 19562
rect 1664 19530 1704 19562
rect 1736 19530 1776 19562
rect 1808 19530 1848 19562
rect 1880 19530 2000 19562
rect 0 19490 2000 19530
rect 0 19458 120 19490
rect 152 19458 192 19490
rect 224 19458 264 19490
rect 296 19458 336 19490
rect 368 19458 408 19490
rect 440 19458 480 19490
rect 512 19458 552 19490
rect 584 19458 624 19490
rect 656 19458 696 19490
rect 728 19458 768 19490
rect 800 19458 840 19490
rect 872 19458 912 19490
rect 944 19458 984 19490
rect 1016 19458 1056 19490
rect 1088 19458 1128 19490
rect 1160 19458 1200 19490
rect 1232 19458 1272 19490
rect 1304 19458 1344 19490
rect 1376 19458 1416 19490
rect 1448 19458 1488 19490
rect 1520 19458 1560 19490
rect 1592 19458 1632 19490
rect 1664 19458 1704 19490
rect 1736 19458 1776 19490
rect 1808 19458 1848 19490
rect 1880 19458 2000 19490
rect 0 19418 2000 19458
rect 0 19386 120 19418
rect 152 19386 192 19418
rect 224 19386 264 19418
rect 296 19386 336 19418
rect 368 19386 408 19418
rect 440 19386 480 19418
rect 512 19386 552 19418
rect 584 19386 624 19418
rect 656 19386 696 19418
rect 728 19386 768 19418
rect 800 19386 840 19418
rect 872 19386 912 19418
rect 944 19386 984 19418
rect 1016 19386 1056 19418
rect 1088 19386 1128 19418
rect 1160 19386 1200 19418
rect 1232 19386 1272 19418
rect 1304 19386 1344 19418
rect 1376 19386 1416 19418
rect 1448 19386 1488 19418
rect 1520 19386 1560 19418
rect 1592 19386 1632 19418
rect 1664 19386 1704 19418
rect 1736 19386 1776 19418
rect 1808 19386 1848 19418
rect 1880 19386 2000 19418
rect 0 19346 2000 19386
rect 0 19314 120 19346
rect 152 19314 192 19346
rect 224 19314 264 19346
rect 296 19314 336 19346
rect 368 19314 408 19346
rect 440 19314 480 19346
rect 512 19314 552 19346
rect 584 19314 624 19346
rect 656 19314 696 19346
rect 728 19314 768 19346
rect 800 19314 840 19346
rect 872 19314 912 19346
rect 944 19314 984 19346
rect 1016 19314 1056 19346
rect 1088 19314 1128 19346
rect 1160 19314 1200 19346
rect 1232 19314 1272 19346
rect 1304 19314 1344 19346
rect 1376 19314 1416 19346
rect 1448 19314 1488 19346
rect 1520 19314 1560 19346
rect 1592 19314 1632 19346
rect 1664 19314 1704 19346
rect 1736 19314 1776 19346
rect 1808 19314 1848 19346
rect 1880 19314 2000 19346
rect 0 19274 2000 19314
rect 0 19242 120 19274
rect 152 19242 192 19274
rect 224 19242 264 19274
rect 296 19242 336 19274
rect 368 19242 408 19274
rect 440 19242 480 19274
rect 512 19242 552 19274
rect 584 19242 624 19274
rect 656 19242 696 19274
rect 728 19242 768 19274
rect 800 19242 840 19274
rect 872 19242 912 19274
rect 944 19242 984 19274
rect 1016 19242 1056 19274
rect 1088 19242 1128 19274
rect 1160 19242 1200 19274
rect 1232 19242 1272 19274
rect 1304 19242 1344 19274
rect 1376 19242 1416 19274
rect 1448 19242 1488 19274
rect 1520 19242 1560 19274
rect 1592 19242 1632 19274
rect 1664 19242 1704 19274
rect 1736 19242 1776 19274
rect 1808 19242 1848 19274
rect 1880 19242 2000 19274
rect 0 19202 2000 19242
rect 0 19170 120 19202
rect 152 19170 192 19202
rect 224 19170 264 19202
rect 296 19170 336 19202
rect 368 19170 408 19202
rect 440 19170 480 19202
rect 512 19170 552 19202
rect 584 19170 624 19202
rect 656 19170 696 19202
rect 728 19170 768 19202
rect 800 19170 840 19202
rect 872 19170 912 19202
rect 944 19170 984 19202
rect 1016 19170 1056 19202
rect 1088 19170 1128 19202
rect 1160 19170 1200 19202
rect 1232 19170 1272 19202
rect 1304 19170 1344 19202
rect 1376 19170 1416 19202
rect 1448 19170 1488 19202
rect 1520 19170 1560 19202
rect 1592 19170 1632 19202
rect 1664 19170 1704 19202
rect 1736 19170 1776 19202
rect 1808 19170 1848 19202
rect 1880 19170 2000 19202
rect 0 19130 2000 19170
rect 0 19098 120 19130
rect 152 19098 192 19130
rect 224 19098 264 19130
rect 296 19098 336 19130
rect 368 19098 408 19130
rect 440 19098 480 19130
rect 512 19098 552 19130
rect 584 19098 624 19130
rect 656 19098 696 19130
rect 728 19098 768 19130
rect 800 19098 840 19130
rect 872 19098 912 19130
rect 944 19098 984 19130
rect 1016 19098 1056 19130
rect 1088 19098 1128 19130
rect 1160 19098 1200 19130
rect 1232 19098 1272 19130
rect 1304 19098 1344 19130
rect 1376 19098 1416 19130
rect 1448 19098 1488 19130
rect 1520 19098 1560 19130
rect 1592 19098 1632 19130
rect 1664 19098 1704 19130
rect 1736 19098 1776 19130
rect 1808 19098 1848 19130
rect 1880 19098 2000 19130
rect 0 19058 2000 19098
rect 0 19026 120 19058
rect 152 19026 192 19058
rect 224 19026 264 19058
rect 296 19026 336 19058
rect 368 19026 408 19058
rect 440 19026 480 19058
rect 512 19026 552 19058
rect 584 19026 624 19058
rect 656 19026 696 19058
rect 728 19026 768 19058
rect 800 19026 840 19058
rect 872 19026 912 19058
rect 944 19026 984 19058
rect 1016 19026 1056 19058
rect 1088 19026 1128 19058
rect 1160 19026 1200 19058
rect 1232 19026 1272 19058
rect 1304 19026 1344 19058
rect 1376 19026 1416 19058
rect 1448 19026 1488 19058
rect 1520 19026 1560 19058
rect 1592 19026 1632 19058
rect 1664 19026 1704 19058
rect 1736 19026 1776 19058
rect 1808 19026 1848 19058
rect 1880 19026 2000 19058
rect 0 18986 2000 19026
rect 0 18954 120 18986
rect 152 18954 192 18986
rect 224 18954 264 18986
rect 296 18954 336 18986
rect 368 18954 408 18986
rect 440 18954 480 18986
rect 512 18954 552 18986
rect 584 18954 624 18986
rect 656 18954 696 18986
rect 728 18954 768 18986
rect 800 18954 840 18986
rect 872 18954 912 18986
rect 944 18954 984 18986
rect 1016 18954 1056 18986
rect 1088 18954 1128 18986
rect 1160 18954 1200 18986
rect 1232 18954 1272 18986
rect 1304 18954 1344 18986
rect 1376 18954 1416 18986
rect 1448 18954 1488 18986
rect 1520 18954 1560 18986
rect 1592 18954 1632 18986
rect 1664 18954 1704 18986
rect 1736 18954 1776 18986
rect 1808 18954 1848 18986
rect 1880 18954 2000 18986
rect 0 18914 2000 18954
rect 0 18882 120 18914
rect 152 18882 192 18914
rect 224 18882 264 18914
rect 296 18882 336 18914
rect 368 18882 408 18914
rect 440 18882 480 18914
rect 512 18882 552 18914
rect 584 18882 624 18914
rect 656 18882 696 18914
rect 728 18882 768 18914
rect 800 18882 840 18914
rect 872 18882 912 18914
rect 944 18882 984 18914
rect 1016 18882 1056 18914
rect 1088 18882 1128 18914
rect 1160 18882 1200 18914
rect 1232 18882 1272 18914
rect 1304 18882 1344 18914
rect 1376 18882 1416 18914
rect 1448 18882 1488 18914
rect 1520 18882 1560 18914
rect 1592 18882 1632 18914
rect 1664 18882 1704 18914
rect 1736 18882 1776 18914
rect 1808 18882 1848 18914
rect 1880 18882 2000 18914
rect 0 18842 2000 18882
rect 0 18810 120 18842
rect 152 18810 192 18842
rect 224 18810 264 18842
rect 296 18810 336 18842
rect 368 18810 408 18842
rect 440 18810 480 18842
rect 512 18810 552 18842
rect 584 18810 624 18842
rect 656 18810 696 18842
rect 728 18810 768 18842
rect 800 18810 840 18842
rect 872 18810 912 18842
rect 944 18810 984 18842
rect 1016 18810 1056 18842
rect 1088 18810 1128 18842
rect 1160 18810 1200 18842
rect 1232 18810 1272 18842
rect 1304 18810 1344 18842
rect 1376 18810 1416 18842
rect 1448 18810 1488 18842
rect 1520 18810 1560 18842
rect 1592 18810 1632 18842
rect 1664 18810 1704 18842
rect 1736 18810 1776 18842
rect 1808 18810 1848 18842
rect 1880 18810 2000 18842
rect 0 18770 2000 18810
rect 0 18738 120 18770
rect 152 18738 192 18770
rect 224 18738 264 18770
rect 296 18738 336 18770
rect 368 18738 408 18770
rect 440 18738 480 18770
rect 512 18738 552 18770
rect 584 18738 624 18770
rect 656 18738 696 18770
rect 728 18738 768 18770
rect 800 18738 840 18770
rect 872 18738 912 18770
rect 944 18738 984 18770
rect 1016 18738 1056 18770
rect 1088 18738 1128 18770
rect 1160 18738 1200 18770
rect 1232 18738 1272 18770
rect 1304 18738 1344 18770
rect 1376 18738 1416 18770
rect 1448 18738 1488 18770
rect 1520 18738 1560 18770
rect 1592 18738 1632 18770
rect 1664 18738 1704 18770
rect 1736 18738 1776 18770
rect 1808 18738 1848 18770
rect 1880 18738 2000 18770
rect 0 18698 2000 18738
rect 0 18666 120 18698
rect 152 18666 192 18698
rect 224 18666 264 18698
rect 296 18666 336 18698
rect 368 18666 408 18698
rect 440 18666 480 18698
rect 512 18666 552 18698
rect 584 18666 624 18698
rect 656 18666 696 18698
rect 728 18666 768 18698
rect 800 18666 840 18698
rect 872 18666 912 18698
rect 944 18666 984 18698
rect 1016 18666 1056 18698
rect 1088 18666 1128 18698
rect 1160 18666 1200 18698
rect 1232 18666 1272 18698
rect 1304 18666 1344 18698
rect 1376 18666 1416 18698
rect 1448 18666 1488 18698
rect 1520 18666 1560 18698
rect 1592 18666 1632 18698
rect 1664 18666 1704 18698
rect 1736 18666 1776 18698
rect 1808 18666 1848 18698
rect 1880 18666 2000 18698
rect 0 18626 2000 18666
rect 0 18594 120 18626
rect 152 18594 192 18626
rect 224 18594 264 18626
rect 296 18594 336 18626
rect 368 18594 408 18626
rect 440 18594 480 18626
rect 512 18594 552 18626
rect 584 18594 624 18626
rect 656 18594 696 18626
rect 728 18594 768 18626
rect 800 18594 840 18626
rect 872 18594 912 18626
rect 944 18594 984 18626
rect 1016 18594 1056 18626
rect 1088 18594 1128 18626
rect 1160 18594 1200 18626
rect 1232 18594 1272 18626
rect 1304 18594 1344 18626
rect 1376 18594 1416 18626
rect 1448 18594 1488 18626
rect 1520 18594 1560 18626
rect 1592 18594 1632 18626
rect 1664 18594 1704 18626
rect 1736 18594 1776 18626
rect 1808 18594 1848 18626
rect 1880 18594 2000 18626
rect 0 18554 2000 18594
rect 0 18522 120 18554
rect 152 18522 192 18554
rect 224 18522 264 18554
rect 296 18522 336 18554
rect 368 18522 408 18554
rect 440 18522 480 18554
rect 512 18522 552 18554
rect 584 18522 624 18554
rect 656 18522 696 18554
rect 728 18522 768 18554
rect 800 18522 840 18554
rect 872 18522 912 18554
rect 944 18522 984 18554
rect 1016 18522 1056 18554
rect 1088 18522 1128 18554
rect 1160 18522 1200 18554
rect 1232 18522 1272 18554
rect 1304 18522 1344 18554
rect 1376 18522 1416 18554
rect 1448 18522 1488 18554
rect 1520 18522 1560 18554
rect 1592 18522 1632 18554
rect 1664 18522 1704 18554
rect 1736 18522 1776 18554
rect 1808 18522 1848 18554
rect 1880 18522 2000 18554
rect 0 18482 2000 18522
rect 0 18450 120 18482
rect 152 18450 192 18482
rect 224 18450 264 18482
rect 296 18450 336 18482
rect 368 18450 408 18482
rect 440 18450 480 18482
rect 512 18450 552 18482
rect 584 18450 624 18482
rect 656 18450 696 18482
rect 728 18450 768 18482
rect 800 18450 840 18482
rect 872 18450 912 18482
rect 944 18450 984 18482
rect 1016 18450 1056 18482
rect 1088 18450 1128 18482
rect 1160 18450 1200 18482
rect 1232 18450 1272 18482
rect 1304 18450 1344 18482
rect 1376 18450 1416 18482
rect 1448 18450 1488 18482
rect 1520 18450 1560 18482
rect 1592 18450 1632 18482
rect 1664 18450 1704 18482
rect 1736 18450 1776 18482
rect 1808 18450 1848 18482
rect 1880 18450 2000 18482
rect 0 18410 2000 18450
rect 0 18378 120 18410
rect 152 18378 192 18410
rect 224 18378 264 18410
rect 296 18378 336 18410
rect 368 18378 408 18410
rect 440 18378 480 18410
rect 512 18378 552 18410
rect 584 18378 624 18410
rect 656 18378 696 18410
rect 728 18378 768 18410
rect 800 18378 840 18410
rect 872 18378 912 18410
rect 944 18378 984 18410
rect 1016 18378 1056 18410
rect 1088 18378 1128 18410
rect 1160 18378 1200 18410
rect 1232 18378 1272 18410
rect 1304 18378 1344 18410
rect 1376 18378 1416 18410
rect 1448 18378 1488 18410
rect 1520 18378 1560 18410
rect 1592 18378 1632 18410
rect 1664 18378 1704 18410
rect 1736 18378 1776 18410
rect 1808 18378 1848 18410
rect 1880 18378 2000 18410
rect 0 18338 2000 18378
rect 0 18306 120 18338
rect 152 18306 192 18338
rect 224 18306 264 18338
rect 296 18306 336 18338
rect 368 18306 408 18338
rect 440 18306 480 18338
rect 512 18306 552 18338
rect 584 18306 624 18338
rect 656 18306 696 18338
rect 728 18306 768 18338
rect 800 18306 840 18338
rect 872 18306 912 18338
rect 944 18306 984 18338
rect 1016 18306 1056 18338
rect 1088 18306 1128 18338
rect 1160 18306 1200 18338
rect 1232 18306 1272 18338
rect 1304 18306 1344 18338
rect 1376 18306 1416 18338
rect 1448 18306 1488 18338
rect 1520 18306 1560 18338
rect 1592 18306 1632 18338
rect 1664 18306 1704 18338
rect 1736 18306 1776 18338
rect 1808 18306 1848 18338
rect 1880 18306 2000 18338
rect 0 18266 2000 18306
rect 0 18234 120 18266
rect 152 18234 192 18266
rect 224 18234 264 18266
rect 296 18234 336 18266
rect 368 18234 408 18266
rect 440 18234 480 18266
rect 512 18234 552 18266
rect 584 18234 624 18266
rect 656 18234 696 18266
rect 728 18234 768 18266
rect 800 18234 840 18266
rect 872 18234 912 18266
rect 944 18234 984 18266
rect 1016 18234 1056 18266
rect 1088 18234 1128 18266
rect 1160 18234 1200 18266
rect 1232 18234 1272 18266
rect 1304 18234 1344 18266
rect 1376 18234 1416 18266
rect 1448 18234 1488 18266
rect 1520 18234 1560 18266
rect 1592 18234 1632 18266
rect 1664 18234 1704 18266
rect 1736 18234 1776 18266
rect 1808 18234 1848 18266
rect 1880 18234 2000 18266
rect 0 18194 2000 18234
rect 0 18162 120 18194
rect 152 18162 192 18194
rect 224 18162 264 18194
rect 296 18162 336 18194
rect 368 18162 408 18194
rect 440 18162 480 18194
rect 512 18162 552 18194
rect 584 18162 624 18194
rect 656 18162 696 18194
rect 728 18162 768 18194
rect 800 18162 840 18194
rect 872 18162 912 18194
rect 944 18162 984 18194
rect 1016 18162 1056 18194
rect 1088 18162 1128 18194
rect 1160 18162 1200 18194
rect 1232 18162 1272 18194
rect 1304 18162 1344 18194
rect 1376 18162 1416 18194
rect 1448 18162 1488 18194
rect 1520 18162 1560 18194
rect 1592 18162 1632 18194
rect 1664 18162 1704 18194
rect 1736 18162 1776 18194
rect 1808 18162 1848 18194
rect 1880 18162 2000 18194
rect 0 18112 2000 18162
rect 0 17848 2000 17912
rect 0 17816 120 17848
rect 152 17816 192 17848
rect 224 17816 264 17848
rect 296 17816 336 17848
rect 368 17816 408 17848
rect 440 17816 480 17848
rect 512 17816 552 17848
rect 584 17816 624 17848
rect 656 17816 696 17848
rect 728 17816 768 17848
rect 800 17816 840 17848
rect 872 17816 912 17848
rect 944 17816 984 17848
rect 1016 17816 1056 17848
rect 1088 17816 1128 17848
rect 1160 17816 1200 17848
rect 1232 17816 1272 17848
rect 1304 17816 1344 17848
rect 1376 17816 1416 17848
rect 1448 17816 1488 17848
rect 1520 17816 1560 17848
rect 1592 17816 1632 17848
rect 1664 17816 1704 17848
rect 1736 17816 1776 17848
rect 1808 17816 1848 17848
rect 1880 17816 2000 17848
rect 0 17776 2000 17816
rect 0 17744 120 17776
rect 152 17744 192 17776
rect 224 17744 264 17776
rect 296 17744 336 17776
rect 368 17744 408 17776
rect 440 17744 480 17776
rect 512 17744 552 17776
rect 584 17744 624 17776
rect 656 17744 696 17776
rect 728 17744 768 17776
rect 800 17744 840 17776
rect 872 17744 912 17776
rect 944 17744 984 17776
rect 1016 17744 1056 17776
rect 1088 17744 1128 17776
rect 1160 17744 1200 17776
rect 1232 17744 1272 17776
rect 1304 17744 1344 17776
rect 1376 17744 1416 17776
rect 1448 17744 1488 17776
rect 1520 17744 1560 17776
rect 1592 17744 1632 17776
rect 1664 17744 1704 17776
rect 1736 17744 1776 17776
rect 1808 17744 1848 17776
rect 1880 17744 2000 17776
rect 0 17704 2000 17744
rect 0 17672 120 17704
rect 152 17672 192 17704
rect 224 17672 264 17704
rect 296 17672 336 17704
rect 368 17672 408 17704
rect 440 17672 480 17704
rect 512 17672 552 17704
rect 584 17672 624 17704
rect 656 17672 696 17704
rect 728 17672 768 17704
rect 800 17672 840 17704
rect 872 17672 912 17704
rect 944 17672 984 17704
rect 1016 17672 1056 17704
rect 1088 17672 1128 17704
rect 1160 17672 1200 17704
rect 1232 17672 1272 17704
rect 1304 17672 1344 17704
rect 1376 17672 1416 17704
rect 1448 17672 1488 17704
rect 1520 17672 1560 17704
rect 1592 17672 1632 17704
rect 1664 17672 1704 17704
rect 1736 17672 1776 17704
rect 1808 17672 1848 17704
rect 1880 17672 2000 17704
rect 0 17632 2000 17672
rect 0 17600 120 17632
rect 152 17600 192 17632
rect 224 17600 264 17632
rect 296 17600 336 17632
rect 368 17600 408 17632
rect 440 17600 480 17632
rect 512 17600 552 17632
rect 584 17600 624 17632
rect 656 17600 696 17632
rect 728 17600 768 17632
rect 800 17600 840 17632
rect 872 17600 912 17632
rect 944 17600 984 17632
rect 1016 17600 1056 17632
rect 1088 17600 1128 17632
rect 1160 17600 1200 17632
rect 1232 17600 1272 17632
rect 1304 17600 1344 17632
rect 1376 17600 1416 17632
rect 1448 17600 1488 17632
rect 1520 17600 1560 17632
rect 1592 17600 1632 17632
rect 1664 17600 1704 17632
rect 1736 17600 1776 17632
rect 1808 17600 1848 17632
rect 1880 17600 2000 17632
rect 0 17560 2000 17600
rect 0 17528 120 17560
rect 152 17528 192 17560
rect 224 17528 264 17560
rect 296 17528 336 17560
rect 368 17528 408 17560
rect 440 17528 480 17560
rect 512 17528 552 17560
rect 584 17528 624 17560
rect 656 17528 696 17560
rect 728 17528 768 17560
rect 800 17528 840 17560
rect 872 17528 912 17560
rect 944 17528 984 17560
rect 1016 17528 1056 17560
rect 1088 17528 1128 17560
rect 1160 17528 1200 17560
rect 1232 17528 1272 17560
rect 1304 17528 1344 17560
rect 1376 17528 1416 17560
rect 1448 17528 1488 17560
rect 1520 17528 1560 17560
rect 1592 17528 1632 17560
rect 1664 17528 1704 17560
rect 1736 17528 1776 17560
rect 1808 17528 1848 17560
rect 1880 17528 2000 17560
rect 0 17488 2000 17528
rect 0 17456 120 17488
rect 152 17456 192 17488
rect 224 17456 264 17488
rect 296 17456 336 17488
rect 368 17456 408 17488
rect 440 17456 480 17488
rect 512 17456 552 17488
rect 584 17456 624 17488
rect 656 17456 696 17488
rect 728 17456 768 17488
rect 800 17456 840 17488
rect 872 17456 912 17488
rect 944 17456 984 17488
rect 1016 17456 1056 17488
rect 1088 17456 1128 17488
rect 1160 17456 1200 17488
rect 1232 17456 1272 17488
rect 1304 17456 1344 17488
rect 1376 17456 1416 17488
rect 1448 17456 1488 17488
rect 1520 17456 1560 17488
rect 1592 17456 1632 17488
rect 1664 17456 1704 17488
rect 1736 17456 1776 17488
rect 1808 17456 1848 17488
rect 1880 17456 2000 17488
rect 0 17416 2000 17456
rect 0 17384 120 17416
rect 152 17384 192 17416
rect 224 17384 264 17416
rect 296 17384 336 17416
rect 368 17384 408 17416
rect 440 17384 480 17416
rect 512 17384 552 17416
rect 584 17384 624 17416
rect 656 17384 696 17416
rect 728 17384 768 17416
rect 800 17384 840 17416
rect 872 17384 912 17416
rect 944 17384 984 17416
rect 1016 17384 1056 17416
rect 1088 17384 1128 17416
rect 1160 17384 1200 17416
rect 1232 17384 1272 17416
rect 1304 17384 1344 17416
rect 1376 17384 1416 17416
rect 1448 17384 1488 17416
rect 1520 17384 1560 17416
rect 1592 17384 1632 17416
rect 1664 17384 1704 17416
rect 1736 17384 1776 17416
rect 1808 17384 1848 17416
rect 1880 17384 2000 17416
rect 0 17344 2000 17384
rect 0 17312 120 17344
rect 152 17312 192 17344
rect 224 17312 264 17344
rect 296 17312 336 17344
rect 368 17312 408 17344
rect 440 17312 480 17344
rect 512 17312 552 17344
rect 584 17312 624 17344
rect 656 17312 696 17344
rect 728 17312 768 17344
rect 800 17312 840 17344
rect 872 17312 912 17344
rect 944 17312 984 17344
rect 1016 17312 1056 17344
rect 1088 17312 1128 17344
rect 1160 17312 1200 17344
rect 1232 17312 1272 17344
rect 1304 17312 1344 17344
rect 1376 17312 1416 17344
rect 1448 17312 1488 17344
rect 1520 17312 1560 17344
rect 1592 17312 1632 17344
rect 1664 17312 1704 17344
rect 1736 17312 1776 17344
rect 1808 17312 1848 17344
rect 1880 17312 2000 17344
rect 0 17272 2000 17312
rect 0 17240 120 17272
rect 152 17240 192 17272
rect 224 17240 264 17272
rect 296 17240 336 17272
rect 368 17240 408 17272
rect 440 17240 480 17272
rect 512 17240 552 17272
rect 584 17240 624 17272
rect 656 17240 696 17272
rect 728 17240 768 17272
rect 800 17240 840 17272
rect 872 17240 912 17272
rect 944 17240 984 17272
rect 1016 17240 1056 17272
rect 1088 17240 1128 17272
rect 1160 17240 1200 17272
rect 1232 17240 1272 17272
rect 1304 17240 1344 17272
rect 1376 17240 1416 17272
rect 1448 17240 1488 17272
rect 1520 17240 1560 17272
rect 1592 17240 1632 17272
rect 1664 17240 1704 17272
rect 1736 17240 1776 17272
rect 1808 17240 1848 17272
rect 1880 17240 2000 17272
rect 0 17200 2000 17240
rect 0 17168 120 17200
rect 152 17168 192 17200
rect 224 17168 264 17200
rect 296 17168 336 17200
rect 368 17168 408 17200
rect 440 17168 480 17200
rect 512 17168 552 17200
rect 584 17168 624 17200
rect 656 17168 696 17200
rect 728 17168 768 17200
rect 800 17168 840 17200
rect 872 17168 912 17200
rect 944 17168 984 17200
rect 1016 17168 1056 17200
rect 1088 17168 1128 17200
rect 1160 17168 1200 17200
rect 1232 17168 1272 17200
rect 1304 17168 1344 17200
rect 1376 17168 1416 17200
rect 1448 17168 1488 17200
rect 1520 17168 1560 17200
rect 1592 17168 1632 17200
rect 1664 17168 1704 17200
rect 1736 17168 1776 17200
rect 1808 17168 1848 17200
rect 1880 17168 2000 17200
rect 0 17128 2000 17168
rect 0 17096 120 17128
rect 152 17096 192 17128
rect 224 17096 264 17128
rect 296 17096 336 17128
rect 368 17096 408 17128
rect 440 17096 480 17128
rect 512 17096 552 17128
rect 584 17096 624 17128
rect 656 17096 696 17128
rect 728 17096 768 17128
rect 800 17096 840 17128
rect 872 17096 912 17128
rect 944 17096 984 17128
rect 1016 17096 1056 17128
rect 1088 17096 1128 17128
rect 1160 17096 1200 17128
rect 1232 17096 1272 17128
rect 1304 17096 1344 17128
rect 1376 17096 1416 17128
rect 1448 17096 1488 17128
rect 1520 17096 1560 17128
rect 1592 17096 1632 17128
rect 1664 17096 1704 17128
rect 1736 17096 1776 17128
rect 1808 17096 1848 17128
rect 1880 17096 2000 17128
rect 0 17056 2000 17096
rect 0 17024 120 17056
rect 152 17024 192 17056
rect 224 17024 264 17056
rect 296 17024 336 17056
rect 368 17024 408 17056
rect 440 17024 480 17056
rect 512 17024 552 17056
rect 584 17024 624 17056
rect 656 17024 696 17056
rect 728 17024 768 17056
rect 800 17024 840 17056
rect 872 17024 912 17056
rect 944 17024 984 17056
rect 1016 17024 1056 17056
rect 1088 17024 1128 17056
rect 1160 17024 1200 17056
rect 1232 17024 1272 17056
rect 1304 17024 1344 17056
rect 1376 17024 1416 17056
rect 1448 17024 1488 17056
rect 1520 17024 1560 17056
rect 1592 17024 1632 17056
rect 1664 17024 1704 17056
rect 1736 17024 1776 17056
rect 1808 17024 1848 17056
rect 1880 17024 2000 17056
rect 0 16984 2000 17024
rect 0 16952 120 16984
rect 152 16952 192 16984
rect 224 16952 264 16984
rect 296 16952 336 16984
rect 368 16952 408 16984
rect 440 16952 480 16984
rect 512 16952 552 16984
rect 584 16952 624 16984
rect 656 16952 696 16984
rect 728 16952 768 16984
rect 800 16952 840 16984
rect 872 16952 912 16984
rect 944 16952 984 16984
rect 1016 16952 1056 16984
rect 1088 16952 1128 16984
rect 1160 16952 1200 16984
rect 1232 16952 1272 16984
rect 1304 16952 1344 16984
rect 1376 16952 1416 16984
rect 1448 16952 1488 16984
rect 1520 16952 1560 16984
rect 1592 16952 1632 16984
rect 1664 16952 1704 16984
rect 1736 16952 1776 16984
rect 1808 16952 1848 16984
rect 1880 16952 2000 16984
rect 0 16912 2000 16952
rect 0 16880 120 16912
rect 152 16880 192 16912
rect 224 16880 264 16912
rect 296 16880 336 16912
rect 368 16880 408 16912
rect 440 16880 480 16912
rect 512 16880 552 16912
rect 584 16880 624 16912
rect 656 16880 696 16912
rect 728 16880 768 16912
rect 800 16880 840 16912
rect 872 16880 912 16912
rect 944 16880 984 16912
rect 1016 16880 1056 16912
rect 1088 16880 1128 16912
rect 1160 16880 1200 16912
rect 1232 16880 1272 16912
rect 1304 16880 1344 16912
rect 1376 16880 1416 16912
rect 1448 16880 1488 16912
rect 1520 16880 1560 16912
rect 1592 16880 1632 16912
rect 1664 16880 1704 16912
rect 1736 16880 1776 16912
rect 1808 16880 1848 16912
rect 1880 16880 2000 16912
rect 0 16840 2000 16880
rect 0 16808 120 16840
rect 152 16808 192 16840
rect 224 16808 264 16840
rect 296 16808 336 16840
rect 368 16808 408 16840
rect 440 16808 480 16840
rect 512 16808 552 16840
rect 584 16808 624 16840
rect 656 16808 696 16840
rect 728 16808 768 16840
rect 800 16808 840 16840
rect 872 16808 912 16840
rect 944 16808 984 16840
rect 1016 16808 1056 16840
rect 1088 16808 1128 16840
rect 1160 16808 1200 16840
rect 1232 16808 1272 16840
rect 1304 16808 1344 16840
rect 1376 16808 1416 16840
rect 1448 16808 1488 16840
rect 1520 16808 1560 16840
rect 1592 16808 1632 16840
rect 1664 16808 1704 16840
rect 1736 16808 1776 16840
rect 1808 16808 1848 16840
rect 1880 16808 2000 16840
rect 0 16768 2000 16808
rect 0 16736 120 16768
rect 152 16736 192 16768
rect 224 16736 264 16768
rect 296 16736 336 16768
rect 368 16736 408 16768
rect 440 16736 480 16768
rect 512 16736 552 16768
rect 584 16736 624 16768
rect 656 16736 696 16768
rect 728 16736 768 16768
rect 800 16736 840 16768
rect 872 16736 912 16768
rect 944 16736 984 16768
rect 1016 16736 1056 16768
rect 1088 16736 1128 16768
rect 1160 16736 1200 16768
rect 1232 16736 1272 16768
rect 1304 16736 1344 16768
rect 1376 16736 1416 16768
rect 1448 16736 1488 16768
rect 1520 16736 1560 16768
rect 1592 16736 1632 16768
rect 1664 16736 1704 16768
rect 1736 16736 1776 16768
rect 1808 16736 1848 16768
rect 1880 16736 2000 16768
rect 0 16696 2000 16736
rect 0 16664 120 16696
rect 152 16664 192 16696
rect 224 16664 264 16696
rect 296 16664 336 16696
rect 368 16664 408 16696
rect 440 16664 480 16696
rect 512 16664 552 16696
rect 584 16664 624 16696
rect 656 16664 696 16696
rect 728 16664 768 16696
rect 800 16664 840 16696
rect 872 16664 912 16696
rect 944 16664 984 16696
rect 1016 16664 1056 16696
rect 1088 16664 1128 16696
rect 1160 16664 1200 16696
rect 1232 16664 1272 16696
rect 1304 16664 1344 16696
rect 1376 16664 1416 16696
rect 1448 16664 1488 16696
rect 1520 16664 1560 16696
rect 1592 16664 1632 16696
rect 1664 16664 1704 16696
rect 1736 16664 1776 16696
rect 1808 16664 1848 16696
rect 1880 16664 2000 16696
rect 0 16624 2000 16664
rect 0 16592 120 16624
rect 152 16592 192 16624
rect 224 16592 264 16624
rect 296 16592 336 16624
rect 368 16592 408 16624
rect 440 16592 480 16624
rect 512 16592 552 16624
rect 584 16592 624 16624
rect 656 16592 696 16624
rect 728 16592 768 16624
rect 800 16592 840 16624
rect 872 16592 912 16624
rect 944 16592 984 16624
rect 1016 16592 1056 16624
rect 1088 16592 1128 16624
rect 1160 16592 1200 16624
rect 1232 16592 1272 16624
rect 1304 16592 1344 16624
rect 1376 16592 1416 16624
rect 1448 16592 1488 16624
rect 1520 16592 1560 16624
rect 1592 16592 1632 16624
rect 1664 16592 1704 16624
rect 1736 16592 1776 16624
rect 1808 16592 1848 16624
rect 1880 16592 2000 16624
rect 0 16552 2000 16592
rect 0 16520 120 16552
rect 152 16520 192 16552
rect 224 16520 264 16552
rect 296 16520 336 16552
rect 368 16520 408 16552
rect 440 16520 480 16552
rect 512 16520 552 16552
rect 584 16520 624 16552
rect 656 16520 696 16552
rect 728 16520 768 16552
rect 800 16520 840 16552
rect 872 16520 912 16552
rect 944 16520 984 16552
rect 1016 16520 1056 16552
rect 1088 16520 1128 16552
rect 1160 16520 1200 16552
rect 1232 16520 1272 16552
rect 1304 16520 1344 16552
rect 1376 16520 1416 16552
rect 1448 16520 1488 16552
rect 1520 16520 1560 16552
rect 1592 16520 1632 16552
rect 1664 16520 1704 16552
rect 1736 16520 1776 16552
rect 1808 16520 1848 16552
rect 1880 16520 2000 16552
rect 0 16480 2000 16520
rect 0 16448 120 16480
rect 152 16448 192 16480
rect 224 16448 264 16480
rect 296 16448 336 16480
rect 368 16448 408 16480
rect 440 16448 480 16480
rect 512 16448 552 16480
rect 584 16448 624 16480
rect 656 16448 696 16480
rect 728 16448 768 16480
rect 800 16448 840 16480
rect 872 16448 912 16480
rect 944 16448 984 16480
rect 1016 16448 1056 16480
rect 1088 16448 1128 16480
rect 1160 16448 1200 16480
rect 1232 16448 1272 16480
rect 1304 16448 1344 16480
rect 1376 16448 1416 16480
rect 1448 16448 1488 16480
rect 1520 16448 1560 16480
rect 1592 16448 1632 16480
rect 1664 16448 1704 16480
rect 1736 16448 1776 16480
rect 1808 16448 1848 16480
rect 1880 16448 2000 16480
rect 0 16408 2000 16448
rect 0 16376 120 16408
rect 152 16376 192 16408
rect 224 16376 264 16408
rect 296 16376 336 16408
rect 368 16376 408 16408
rect 440 16376 480 16408
rect 512 16376 552 16408
rect 584 16376 624 16408
rect 656 16376 696 16408
rect 728 16376 768 16408
rect 800 16376 840 16408
rect 872 16376 912 16408
rect 944 16376 984 16408
rect 1016 16376 1056 16408
rect 1088 16376 1128 16408
rect 1160 16376 1200 16408
rect 1232 16376 1272 16408
rect 1304 16376 1344 16408
rect 1376 16376 1416 16408
rect 1448 16376 1488 16408
rect 1520 16376 1560 16408
rect 1592 16376 1632 16408
rect 1664 16376 1704 16408
rect 1736 16376 1776 16408
rect 1808 16376 1848 16408
rect 1880 16376 2000 16408
rect 0 16336 2000 16376
rect 0 16304 120 16336
rect 152 16304 192 16336
rect 224 16304 264 16336
rect 296 16304 336 16336
rect 368 16304 408 16336
rect 440 16304 480 16336
rect 512 16304 552 16336
rect 584 16304 624 16336
rect 656 16304 696 16336
rect 728 16304 768 16336
rect 800 16304 840 16336
rect 872 16304 912 16336
rect 944 16304 984 16336
rect 1016 16304 1056 16336
rect 1088 16304 1128 16336
rect 1160 16304 1200 16336
rect 1232 16304 1272 16336
rect 1304 16304 1344 16336
rect 1376 16304 1416 16336
rect 1448 16304 1488 16336
rect 1520 16304 1560 16336
rect 1592 16304 1632 16336
rect 1664 16304 1704 16336
rect 1736 16304 1776 16336
rect 1808 16304 1848 16336
rect 1880 16304 2000 16336
rect 0 16264 2000 16304
rect 0 16232 120 16264
rect 152 16232 192 16264
rect 224 16232 264 16264
rect 296 16232 336 16264
rect 368 16232 408 16264
rect 440 16232 480 16264
rect 512 16232 552 16264
rect 584 16232 624 16264
rect 656 16232 696 16264
rect 728 16232 768 16264
rect 800 16232 840 16264
rect 872 16232 912 16264
rect 944 16232 984 16264
rect 1016 16232 1056 16264
rect 1088 16232 1128 16264
rect 1160 16232 1200 16264
rect 1232 16232 1272 16264
rect 1304 16232 1344 16264
rect 1376 16232 1416 16264
rect 1448 16232 1488 16264
rect 1520 16232 1560 16264
rect 1592 16232 1632 16264
rect 1664 16232 1704 16264
rect 1736 16232 1776 16264
rect 1808 16232 1848 16264
rect 1880 16232 2000 16264
rect 0 16192 2000 16232
rect 0 16160 120 16192
rect 152 16160 192 16192
rect 224 16160 264 16192
rect 296 16160 336 16192
rect 368 16160 408 16192
rect 440 16160 480 16192
rect 512 16160 552 16192
rect 584 16160 624 16192
rect 656 16160 696 16192
rect 728 16160 768 16192
rect 800 16160 840 16192
rect 872 16160 912 16192
rect 944 16160 984 16192
rect 1016 16160 1056 16192
rect 1088 16160 1128 16192
rect 1160 16160 1200 16192
rect 1232 16160 1272 16192
rect 1304 16160 1344 16192
rect 1376 16160 1416 16192
rect 1448 16160 1488 16192
rect 1520 16160 1560 16192
rect 1592 16160 1632 16192
rect 1664 16160 1704 16192
rect 1736 16160 1776 16192
rect 1808 16160 1848 16192
rect 1880 16160 2000 16192
rect 0 16120 2000 16160
rect 0 16088 120 16120
rect 152 16088 192 16120
rect 224 16088 264 16120
rect 296 16088 336 16120
rect 368 16088 408 16120
rect 440 16088 480 16120
rect 512 16088 552 16120
rect 584 16088 624 16120
rect 656 16088 696 16120
rect 728 16088 768 16120
rect 800 16088 840 16120
rect 872 16088 912 16120
rect 944 16088 984 16120
rect 1016 16088 1056 16120
rect 1088 16088 1128 16120
rect 1160 16088 1200 16120
rect 1232 16088 1272 16120
rect 1304 16088 1344 16120
rect 1376 16088 1416 16120
rect 1448 16088 1488 16120
rect 1520 16088 1560 16120
rect 1592 16088 1632 16120
rect 1664 16088 1704 16120
rect 1736 16088 1776 16120
rect 1808 16088 1848 16120
rect 1880 16088 2000 16120
rect 0 16048 2000 16088
rect 0 16016 120 16048
rect 152 16016 192 16048
rect 224 16016 264 16048
rect 296 16016 336 16048
rect 368 16016 408 16048
rect 440 16016 480 16048
rect 512 16016 552 16048
rect 584 16016 624 16048
rect 656 16016 696 16048
rect 728 16016 768 16048
rect 800 16016 840 16048
rect 872 16016 912 16048
rect 944 16016 984 16048
rect 1016 16016 1056 16048
rect 1088 16016 1128 16048
rect 1160 16016 1200 16048
rect 1232 16016 1272 16048
rect 1304 16016 1344 16048
rect 1376 16016 1416 16048
rect 1448 16016 1488 16048
rect 1520 16016 1560 16048
rect 1592 16016 1632 16048
rect 1664 16016 1704 16048
rect 1736 16016 1776 16048
rect 1808 16016 1848 16048
rect 1880 16016 2000 16048
rect 0 15976 2000 16016
rect 0 15944 120 15976
rect 152 15944 192 15976
rect 224 15944 264 15976
rect 296 15944 336 15976
rect 368 15944 408 15976
rect 440 15944 480 15976
rect 512 15944 552 15976
rect 584 15944 624 15976
rect 656 15944 696 15976
rect 728 15944 768 15976
rect 800 15944 840 15976
rect 872 15944 912 15976
rect 944 15944 984 15976
rect 1016 15944 1056 15976
rect 1088 15944 1128 15976
rect 1160 15944 1200 15976
rect 1232 15944 1272 15976
rect 1304 15944 1344 15976
rect 1376 15944 1416 15976
rect 1448 15944 1488 15976
rect 1520 15944 1560 15976
rect 1592 15944 1632 15976
rect 1664 15944 1704 15976
rect 1736 15944 1776 15976
rect 1808 15944 1848 15976
rect 1880 15944 2000 15976
rect 0 15904 2000 15944
rect 0 15872 120 15904
rect 152 15872 192 15904
rect 224 15872 264 15904
rect 296 15872 336 15904
rect 368 15872 408 15904
rect 440 15872 480 15904
rect 512 15872 552 15904
rect 584 15872 624 15904
rect 656 15872 696 15904
rect 728 15872 768 15904
rect 800 15872 840 15904
rect 872 15872 912 15904
rect 944 15872 984 15904
rect 1016 15872 1056 15904
rect 1088 15872 1128 15904
rect 1160 15872 1200 15904
rect 1232 15872 1272 15904
rect 1304 15872 1344 15904
rect 1376 15872 1416 15904
rect 1448 15872 1488 15904
rect 1520 15872 1560 15904
rect 1592 15872 1632 15904
rect 1664 15872 1704 15904
rect 1736 15872 1776 15904
rect 1808 15872 1848 15904
rect 1880 15872 2000 15904
rect 0 15832 2000 15872
rect 0 15800 120 15832
rect 152 15800 192 15832
rect 224 15800 264 15832
rect 296 15800 336 15832
rect 368 15800 408 15832
rect 440 15800 480 15832
rect 512 15800 552 15832
rect 584 15800 624 15832
rect 656 15800 696 15832
rect 728 15800 768 15832
rect 800 15800 840 15832
rect 872 15800 912 15832
rect 944 15800 984 15832
rect 1016 15800 1056 15832
rect 1088 15800 1128 15832
rect 1160 15800 1200 15832
rect 1232 15800 1272 15832
rect 1304 15800 1344 15832
rect 1376 15800 1416 15832
rect 1448 15800 1488 15832
rect 1520 15800 1560 15832
rect 1592 15800 1632 15832
rect 1664 15800 1704 15832
rect 1736 15800 1776 15832
rect 1808 15800 1848 15832
rect 1880 15800 2000 15832
rect 0 15760 2000 15800
rect 0 15728 120 15760
rect 152 15728 192 15760
rect 224 15728 264 15760
rect 296 15728 336 15760
rect 368 15728 408 15760
rect 440 15728 480 15760
rect 512 15728 552 15760
rect 584 15728 624 15760
rect 656 15728 696 15760
rect 728 15728 768 15760
rect 800 15728 840 15760
rect 872 15728 912 15760
rect 944 15728 984 15760
rect 1016 15728 1056 15760
rect 1088 15728 1128 15760
rect 1160 15728 1200 15760
rect 1232 15728 1272 15760
rect 1304 15728 1344 15760
rect 1376 15728 1416 15760
rect 1448 15728 1488 15760
rect 1520 15728 1560 15760
rect 1592 15728 1632 15760
rect 1664 15728 1704 15760
rect 1736 15728 1776 15760
rect 1808 15728 1848 15760
rect 1880 15728 2000 15760
rect 0 15688 2000 15728
rect 0 15656 120 15688
rect 152 15656 192 15688
rect 224 15656 264 15688
rect 296 15656 336 15688
rect 368 15656 408 15688
rect 440 15656 480 15688
rect 512 15656 552 15688
rect 584 15656 624 15688
rect 656 15656 696 15688
rect 728 15656 768 15688
rect 800 15656 840 15688
rect 872 15656 912 15688
rect 944 15656 984 15688
rect 1016 15656 1056 15688
rect 1088 15656 1128 15688
rect 1160 15656 1200 15688
rect 1232 15656 1272 15688
rect 1304 15656 1344 15688
rect 1376 15656 1416 15688
rect 1448 15656 1488 15688
rect 1520 15656 1560 15688
rect 1592 15656 1632 15688
rect 1664 15656 1704 15688
rect 1736 15656 1776 15688
rect 1808 15656 1848 15688
rect 1880 15656 2000 15688
rect 0 15616 2000 15656
rect 0 15584 120 15616
rect 152 15584 192 15616
rect 224 15584 264 15616
rect 296 15584 336 15616
rect 368 15584 408 15616
rect 440 15584 480 15616
rect 512 15584 552 15616
rect 584 15584 624 15616
rect 656 15584 696 15616
rect 728 15584 768 15616
rect 800 15584 840 15616
rect 872 15584 912 15616
rect 944 15584 984 15616
rect 1016 15584 1056 15616
rect 1088 15584 1128 15616
rect 1160 15584 1200 15616
rect 1232 15584 1272 15616
rect 1304 15584 1344 15616
rect 1376 15584 1416 15616
rect 1448 15584 1488 15616
rect 1520 15584 1560 15616
rect 1592 15584 1632 15616
rect 1664 15584 1704 15616
rect 1736 15584 1776 15616
rect 1808 15584 1848 15616
rect 1880 15584 2000 15616
rect 0 15544 2000 15584
rect 0 15512 120 15544
rect 152 15512 192 15544
rect 224 15512 264 15544
rect 296 15512 336 15544
rect 368 15512 408 15544
rect 440 15512 480 15544
rect 512 15512 552 15544
rect 584 15512 624 15544
rect 656 15512 696 15544
rect 728 15512 768 15544
rect 800 15512 840 15544
rect 872 15512 912 15544
rect 944 15512 984 15544
rect 1016 15512 1056 15544
rect 1088 15512 1128 15544
rect 1160 15512 1200 15544
rect 1232 15512 1272 15544
rect 1304 15512 1344 15544
rect 1376 15512 1416 15544
rect 1448 15512 1488 15544
rect 1520 15512 1560 15544
rect 1592 15512 1632 15544
rect 1664 15512 1704 15544
rect 1736 15512 1776 15544
rect 1808 15512 1848 15544
rect 1880 15512 2000 15544
rect 0 15472 2000 15512
rect 0 15440 120 15472
rect 152 15440 192 15472
rect 224 15440 264 15472
rect 296 15440 336 15472
rect 368 15440 408 15472
rect 440 15440 480 15472
rect 512 15440 552 15472
rect 584 15440 624 15472
rect 656 15440 696 15472
rect 728 15440 768 15472
rect 800 15440 840 15472
rect 872 15440 912 15472
rect 944 15440 984 15472
rect 1016 15440 1056 15472
rect 1088 15440 1128 15472
rect 1160 15440 1200 15472
rect 1232 15440 1272 15472
rect 1304 15440 1344 15472
rect 1376 15440 1416 15472
rect 1448 15440 1488 15472
rect 1520 15440 1560 15472
rect 1592 15440 1632 15472
rect 1664 15440 1704 15472
rect 1736 15440 1776 15472
rect 1808 15440 1848 15472
rect 1880 15440 2000 15472
rect 0 15400 2000 15440
rect 0 15368 120 15400
rect 152 15368 192 15400
rect 224 15368 264 15400
rect 296 15368 336 15400
rect 368 15368 408 15400
rect 440 15368 480 15400
rect 512 15368 552 15400
rect 584 15368 624 15400
rect 656 15368 696 15400
rect 728 15368 768 15400
rect 800 15368 840 15400
rect 872 15368 912 15400
rect 944 15368 984 15400
rect 1016 15368 1056 15400
rect 1088 15368 1128 15400
rect 1160 15368 1200 15400
rect 1232 15368 1272 15400
rect 1304 15368 1344 15400
rect 1376 15368 1416 15400
rect 1448 15368 1488 15400
rect 1520 15368 1560 15400
rect 1592 15368 1632 15400
rect 1664 15368 1704 15400
rect 1736 15368 1776 15400
rect 1808 15368 1848 15400
rect 1880 15368 2000 15400
rect 0 15328 2000 15368
rect 0 15296 120 15328
rect 152 15296 192 15328
rect 224 15296 264 15328
rect 296 15296 336 15328
rect 368 15296 408 15328
rect 440 15296 480 15328
rect 512 15296 552 15328
rect 584 15296 624 15328
rect 656 15296 696 15328
rect 728 15296 768 15328
rect 800 15296 840 15328
rect 872 15296 912 15328
rect 944 15296 984 15328
rect 1016 15296 1056 15328
rect 1088 15296 1128 15328
rect 1160 15296 1200 15328
rect 1232 15296 1272 15328
rect 1304 15296 1344 15328
rect 1376 15296 1416 15328
rect 1448 15296 1488 15328
rect 1520 15296 1560 15328
rect 1592 15296 1632 15328
rect 1664 15296 1704 15328
rect 1736 15296 1776 15328
rect 1808 15296 1848 15328
rect 1880 15296 2000 15328
rect 0 15256 2000 15296
rect 0 15224 120 15256
rect 152 15224 192 15256
rect 224 15224 264 15256
rect 296 15224 336 15256
rect 368 15224 408 15256
rect 440 15224 480 15256
rect 512 15224 552 15256
rect 584 15224 624 15256
rect 656 15224 696 15256
rect 728 15224 768 15256
rect 800 15224 840 15256
rect 872 15224 912 15256
rect 944 15224 984 15256
rect 1016 15224 1056 15256
rect 1088 15224 1128 15256
rect 1160 15224 1200 15256
rect 1232 15224 1272 15256
rect 1304 15224 1344 15256
rect 1376 15224 1416 15256
rect 1448 15224 1488 15256
rect 1520 15224 1560 15256
rect 1592 15224 1632 15256
rect 1664 15224 1704 15256
rect 1736 15224 1776 15256
rect 1808 15224 1848 15256
rect 1880 15224 2000 15256
rect 0 15184 2000 15224
rect 0 15152 120 15184
rect 152 15152 192 15184
rect 224 15152 264 15184
rect 296 15152 336 15184
rect 368 15152 408 15184
rect 440 15152 480 15184
rect 512 15152 552 15184
rect 584 15152 624 15184
rect 656 15152 696 15184
rect 728 15152 768 15184
rect 800 15152 840 15184
rect 872 15152 912 15184
rect 944 15152 984 15184
rect 1016 15152 1056 15184
rect 1088 15152 1128 15184
rect 1160 15152 1200 15184
rect 1232 15152 1272 15184
rect 1304 15152 1344 15184
rect 1376 15152 1416 15184
rect 1448 15152 1488 15184
rect 1520 15152 1560 15184
rect 1592 15152 1632 15184
rect 1664 15152 1704 15184
rect 1736 15152 1776 15184
rect 1808 15152 1848 15184
rect 1880 15152 2000 15184
rect 0 15112 2000 15152
rect 0 15080 120 15112
rect 152 15080 192 15112
rect 224 15080 264 15112
rect 296 15080 336 15112
rect 368 15080 408 15112
rect 440 15080 480 15112
rect 512 15080 552 15112
rect 584 15080 624 15112
rect 656 15080 696 15112
rect 728 15080 768 15112
rect 800 15080 840 15112
rect 872 15080 912 15112
rect 944 15080 984 15112
rect 1016 15080 1056 15112
rect 1088 15080 1128 15112
rect 1160 15080 1200 15112
rect 1232 15080 1272 15112
rect 1304 15080 1344 15112
rect 1376 15080 1416 15112
rect 1448 15080 1488 15112
rect 1520 15080 1560 15112
rect 1592 15080 1632 15112
rect 1664 15080 1704 15112
rect 1736 15080 1776 15112
rect 1808 15080 1848 15112
rect 1880 15080 2000 15112
rect 0 15040 2000 15080
rect 0 15008 120 15040
rect 152 15008 192 15040
rect 224 15008 264 15040
rect 296 15008 336 15040
rect 368 15008 408 15040
rect 440 15008 480 15040
rect 512 15008 552 15040
rect 584 15008 624 15040
rect 656 15008 696 15040
rect 728 15008 768 15040
rect 800 15008 840 15040
rect 872 15008 912 15040
rect 944 15008 984 15040
rect 1016 15008 1056 15040
rect 1088 15008 1128 15040
rect 1160 15008 1200 15040
rect 1232 15008 1272 15040
rect 1304 15008 1344 15040
rect 1376 15008 1416 15040
rect 1448 15008 1488 15040
rect 1520 15008 1560 15040
rect 1592 15008 1632 15040
rect 1664 15008 1704 15040
rect 1736 15008 1776 15040
rect 1808 15008 1848 15040
rect 1880 15008 2000 15040
rect 0 14968 2000 15008
rect 0 14936 120 14968
rect 152 14936 192 14968
rect 224 14936 264 14968
rect 296 14936 336 14968
rect 368 14936 408 14968
rect 440 14936 480 14968
rect 512 14936 552 14968
rect 584 14936 624 14968
rect 656 14936 696 14968
rect 728 14936 768 14968
rect 800 14936 840 14968
rect 872 14936 912 14968
rect 944 14936 984 14968
rect 1016 14936 1056 14968
rect 1088 14936 1128 14968
rect 1160 14936 1200 14968
rect 1232 14936 1272 14968
rect 1304 14936 1344 14968
rect 1376 14936 1416 14968
rect 1448 14936 1488 14968
rect 1520 14936 1560 14968
rect 1592 14936 1632 14968
rect 1664 14936 1704 14968
rect 1736 14936 1776 14968
rect 1808 14936 1848 14968
rect 1880 14936 2000 14968
rect 0 14896 2000 14936
rect 0 14864 120 14896
rect 152 14864 192 14896
rect 224 14864 264 14896
rect 296 14864 336 14896
rect 368 14864 408 14896
rect 440 14864 480 14896
rect 512 14864 552 14896
rect 584 14864 624 14896
rect 656 14864 696 14896
rect 728 14864 768 14896
rect 800 14864 840 14896
rect 872 14864 912 14896
rect 944 14864 984 14896
rect 1016 14864 1056 14896
rect 1088 14864 1128 14896
rect 1160 14864 1200 14896
rect 1232 14864 1272 14896
rect 1304 14864 1344 14896
rect 1376 14864 1416 14896
rect 1448 14864 1488 14896
rect 1520 14864 1560 14896
rect 1592 14864 1632 14896
rect 1664 14864 1704 14896
rect 1736 14864 1776 14896
rect 1808 14864 1848 14896
rect 1880 14864 2000 14896
rect 0 14824 2000 14864
rect 0 14792 120 14824
rect 152 14792 192 14824
rect 224 14792 264 14824
rect 296 14792 336 14824
rect 368 14792 408 14824
rect 440 14792 480 14824
rect 512 14792 552 14824
rect 584 14792 624 14824
rect 656 14792 696 14824
rect 728 14792 768 14824
rect 800 14792 840 14824
rect 872 14792 912 14824
rect 944 14792 984 14824
rect 1016 14792 1056 14824
rect 1088 14792 1128 14824
rect 1160 14792 1200 14824
rect 1232 14792 1272 14824
rect 1304 14792 1344 14824
rect 1376 14792 1416 14824
rect 1448 14792 1488 14824
rect 1520 14792 1560 14824
rect 1592 14792 1632 14824
rect 1664 14792 1704 14824
rect 1736 14792 1776 14824
rect 1808 14792 1848 14824
rect 1880 14792 2000 14824
rect 0 14752 2000 14792
rect 0 14720 120 14752
rect 152 14720 192 14752
rect 224 14720 264 14752
rect 296 14720 336 14752
rect 368 14720 408 14752
rect 440 14720 480 14752
rect 512 14720 552 14752
rect 584 14720 624 14752
rect 656 14720 696 14752
rect 728 14720 768 14752
rect 800 14720 840 14752
rect 872 14720 912 14752
rect 944 14720 984 14752
rect 1016 14720 1056 14752
rect 1088 14720 1128 14752
rect 1160 14720 1200 14752
rect 1232 14720 1272 14752
rect 1304 14720 1344 14752
rect 1376 14720 1416 14752
rect 1448 14720 1488 14752
rect 1520 14720 1560 14752
rect 1592 14720 1632 14752
rect 1664 14720 1704 14752
rect 1736 14720 1776 14752
rect 1808 14720 1848 14752
rect 1880 14720 2000 14752
rect 0 14680 2000 14720
rect 0 14648 120 14680
rect 152 14648 192 14680
rect 224 14648 264 14680
rect 296 14648 336 14680
rect 368 14648 408 14680
rect 440 14648 480 14680
rect 512 14648 552 14680
rect 584 14648 624 14680
rect 656 14648 696 14680
rect 728 14648 768 14680
rect 800 14648 840 14680
rect 872 14648 912 14680
rect 944 14648 984 14680
rect 1016 14648 1056 14680
rect 1088 14648 1128 14680
rect 1160 14648 1200 14680
rect 1232 14648 1272 14680
rect 1304 14648 1344 14680
rect 1376 14648 1416 14680
rect 1448 14648 1488 14680
rect 1520 14648 1560 14680
rect 1592 14648 1632 14680
rect 1664 14648 1704 14680
rect 1736 14648 1776 14680
rect 1808 14648 1848 14680
rect 1880 14648 2000 14680
rect 0 14608 2000 14648
rect 0 14576 120 14608
rect 152 14576 192 14608
rect 224 14576 264 14608
rect 296 14576 336 14608
rect 368 14576 408 14608
rect 440 14576 480 14608
rect 512 14576 552 14608
rect 584 14576 624 14608
rect 656 14576 696 14608
rect 728 14576 768 14608
rect 800 14576 840 14608
rect 872 14576 912 14608
rect 944 14576 984 14608
rect 1016 14576 1056 14608
rect 1088 14576 1128 14608
rect 1160 14576 1200 14608
rect 1232 14576 1272 14608
rect 1304 14576 1344 14608
rect 1376 14576 1416 14608
rect 1448 14576 1488 14608
rect 1520 14576 1560 14608
rect 1592 14576 1632 14608
rect 1664 14576 1704 14608
rect 1736 14576 1776 14608
rect 1808 14576 1848 14608
rect 1880 14576 2000 14608
rect 0 14536 2000 14576
rect 0 14504 120 14536
rect 152 14504 192 14536
rect 224 14504 264 14536
rect 296 14504 336 14536
rect 368 14504 408 14536
rect 440 14504 480 14536
rect 512 14504 552 14536
rect 584 14504 624 14536
rect 656 14504 696 14536
rect 728 14504 768 14536
rect 800 14504 840 14536
rect 872 14504 912 14536
rect 944 14504 984 14536
rect 1016 14504 1056 14536
rect 1088 14504 1128 14536
rect 1160 14504 1200 14536
rect 1232 14504 1272 14536
rect 1304 14504 1344 14536
rect 1376 14504 1416 14536
rect 1448 14504 1488 14536
rect 1520 14504 1560 14536
rect 1592 14504 1632 14536
rect 1664 14504 1704 14536
rect 1736 14504 1776 14536
rect 1808 14504 1848 14536
rect 1880 14504 2000 14536
rect 0 14464 2000 14504
rect 0 14432 120 14464
rect 152 14432 192 14464
rect 224 14432 264 14464
rect 296 14432 336 14464
rect 368 14432 408 14464
rect 440 14432 480 14464
rect 512 14432 552 14464
rect 584 14432 624 14464
rect 656 14432 696 14464
rect 728 14432 768 14464
rect 800 14432 840 14464
rect 872 14432 912 14464
rect 944 14432 984 14464
rect 1016 14432 1056 14464
rect 1088 14432 1128 14464
rect 1160 14432 1200 14464
rect 1232 14432 1272 14464
rect 1304 14432 1344 14464
rect 1376 14432 1416 14464
rect 1448 14432 1488 14464
rect 1520 14432 1560 14464
rect 1592 14432 1632 14464
rect 1664 14432 1704 14464
rect 1736 14432 1776 14464
rect 1808 14432 1848 14464
rect 1880 14432 2000 14464
rect 0 14392 2000 14432
rect 0 14360 120 14392
rect 152 14360 192 14392
rect 224 14360 264 14392
rect 296 14360 336 14392
rect 368 14360 408 14392
rect 440 14360 480 14392
rect 512 14360 552 14392
rect 584 14360 624 14392
rect 656 14360 696 14392
rect 728 14360 768 14392
rect 800 14360 840 14392
rect 872 14360 912 14392
rect 944 14360 984 14392
rect 1016 14360 1056 14392
rect 1088 14360 1128 14392
rect 1160 14360 1200 14392
rect 1232 14360 1272 14392
rect 1304 14360 1344 14392
rect 1376 14360 1416 14392
rect 1448 14360 1488 14392
rect 1520 14360 1560 14392
rect 1592 14360 1632 14392
rect 1664 14360 1704 14392
rect 1736 14360 1776 14392
rect 1808 14360 1848 14392
rect 1880 14360 2000 14392
rect 0 14320 2000 14360
rect 0 14288 120 14320
rect 152 14288 192 14320
rect 224 14288 264 14320
rect 296 14288 336 14320
rect 368 14288 408 14320
rect 440 14288 480 14320
rect 512 14288 552 14320
rect 584 14288 624 14320
rect 656 14288 696 14320
rect 728 14288 768 14320
rect 800 14288 840 14320
rect 872 14288 912 14320
rect 944 14288 984 14320
rect 1016 14288 1056 14320
rect 1088 14288 1128 14320
rect 1160 14288 1200 14320
rect 1232 14288 1272 14320
rect 1304 14288 1344 14320
rect 1376 14288 1416 14320
rect 1448 14288 1488 14320
rect 1520 14288 1560 14320
rect 1592 14288 1632 14320
rect 1664 14288 1704 14320
rect 1736 14288 1776 14320
rect 1808 14288 1848 14320
rect 1880 14288 2000 14320
rect 0 14248 2000 14288
rect 0 14216 120 14248
rect 152 14216 192 14248
rect 224 14216 264 14248
rect 296 14216 336 14248
rect 368 14216 408 14248
rect 440 14216 480 14248
rect 512 14216 552 14248
rect 584 14216 624 14248
rect 656 14216 696 14248
rect 728 14216 768 14248
rect 800 14216 840 14248
rect 872 14216 912 14248
rect 944 14216 984 14248
rect 1016 14216 1056 14248
rect 1088 14216 1128 14248
rect 1160 14216 1200 14248
rect 1232 14216 1272 14248
rect 1304 14216 1344 14248
rect 1376 14216 1416 14248
rect 1448 14216 1488 14248
rect 1520 14216 1560 14248
rect 1592 14216 1632 14248
rect 1664 14216 1704 14248
rect 1736 14216 1776 14248
rect 1808 14216 1848 14248
rect 1880 14216 2000 14248
rect 0 14176 2000 14216
rect 0 14144 120 14176
rect 152 14144 192 14176
rect 224 14144 264 14176
rect 296 14144 336 14176
rect 368 14144 408 14176
rect 440 14144 480 14176
rect 512 14144 552 14176
rect 584 14144 624 14176
rect 656 14144 696 14176
rect 728 14144 768 14176
rect 800 14144 840 14176
rect 872 14144 912 14176
rect 944 14144 984 14176
rect 1016 14144 1056 14176
rect 1088 14144 1128 14176
rect 1160 14144 1200 14176
rect 1232 14144 1272 14176
rect 1304 14144 1344 14176
rect 1376 14144 1416 14176
rect 1448 14144 1488 14176
rect 1520 14144 1560 14176
rect 1592 14144 1632 14176
rect 1664 14144 1704 14176
rect 1736 14144 1776 14176
rect 1808 14144 1848 14176
rect 1880 14144 2000 14176
rect 0 14104 2000 14144
rect 0 14072 120 14104
rect 152 14072 192 14104
rect 224 14072 264 14104
rect 296 14072 336 14104
rect 368 14072 408 14104
rect 440 14072 480 14104
rect 512 14072 552 14104
rect 584 14072 624 14104
rect 656 14072 696 14104
rect 728 14072 768 14104
rect 800 14072 840 14104
rect 872 14072 912 14104
rect 944 14072 984 14104
rect 1016 14072 1056 14104
rect 1088 14072 1128 14104
rect 1160 14072 1200 14104
rect 1232 14072 1272 14104
rect 1304 14072 1344 14104
rect 1376 14072 1416 14104
rect 1448 14072 1488 14104
rect 1520 14072 1560 14104
rect 1592 14072 1632 14104
rect 1664 14072 1704 14104
rect 1736 14072 1776 14104
rect 1808 14072 1848 14104
rect 1880 14072 2000 14104
rect 0 14032 2000 14072
rect 0 14000 120 14032
rect 152 14000 192 14032
rect 224 14000 264 14032
rect 296 14000 336 14032
rect 368 14000 408 14032
rect 440 14000 480 14032
rect 512 14000 552 14032
rect 584 14000 624 14032
rect 656 14000 696 14032
rect 728 14000 768 14032
rect 800 14000 840 14032
rect 872 14000 912 14032
rect 944 14000 984 14032
rect 1016 14000 1056 14032
rect 1088 14000 1128 14032
rect 1160 14000 1200 14032
rect 1232 14000 1272 14032
rect 1304 14000 1344 14032
rect 1376 14000 1416 14032
rect 1448 14000 1488 14032
rect 1520 14000 1560 14032
rect 1592 14000 1632 14032
rect 1664 14000 1704 14032
rect 1736 14000 1776 14032
rect 1808 14000 1848 14032
rect 1880 14000 2000 14032
rect 0 13960 2000 14000
rect 0 13928 120 13960
rect 152 13928 192 13960
rect 224 13928 264 13960
rect 296 13928 336 13960
rect 368 13928 408 13960
rect 440 13928 480 13960
rect 512 13928 552 13960
rect 584 13928 624 13960
rect 656 13928 696 13960
rect 728 13928 768 13960
rect 800 13928 840 13960
rect 872 13928 912 13960
rect 944 13928 984 13960
rect 1016 13928 1056 13960
rect 1088 13928 1128 13960
rect 1160 13928 1200 13960
rect 1232 13928 1272 13960
rect 1304 13928 1344 13960
rect 1376 13928 1416 13960
rect 1448 13928 1488 13960
rect 1520 13928 1560 13960
rect 1592 13928 1632 13960
rect 1664 13928 1704 13960
rect 1736 13928 1776 13960
rect 1808 13928 1848 13960
rect 1880 13928 2000 13960
rect 0 13888 2000 13928
rect 0 13856 120 13888
rect 152 13856 192 13888
rect 224 13856 264 13888
rect 296 13856 336 13888
rect 368 13856 408 13888
rect 440 13856 480 13888
rect 512 13856 552 13888
rect 584 13856 624 13888
rect 656 13856 696 13888
rect 728 13856 768 13888
rect 800 13856 840 13888
rect 872 13856 912 13888
rect 944 13856 984 13888
rect 1016 13856 1056 13888
rect 1088 13856 1128 13888
rect 1160 13856 1200 13888
rect 1232 13856 1272 13888
rect 1304 13856 1344 13888
rect 1376 13856 1416 13888
rect 1448 13856 1488 13888
rect 1520 13856 1560 13888
rect 1592 13856 1632 13888
rect 1664 13856 1704 13888
rect 1736 13856 1776 13888
rect 1808 13856 1848 13888
rect 1880 13856 2000 13888
rect 0 13816 2000 13856
rect 0 13784 120 13816
rect 152 13784 192 13816
rect 224 13784 264 13816
rect 296 13784 336 13816
rect 368 13784 408 13816
rect 440 13784 480 13816
rect 512 13784 552 13816
rect 584 13784 624 13816
rect 656 13784 696 13816
rect 728 13784 768 13816
rect 800 13784 840 13816
rect 872 13784 912 13816
rect 944 13784 984 13816
rect 1016 13784 1056 13816
rect 1088 13784 1128 13816
rect 1160 13784 1200 13816
rect 1232 13784 1272 13816
rect 1304 13784 1344 13816
rect 1376 13784 1416 13816
rect 1448 13784 1488 13816
rect 1520 13784 1560 13816
rect 1592 13784 1632 13816
rect 1664 13784 1704 13816
rect 1736 13784 1776 13816
rect 1808 13784 1848 13816
rect 1880 13784 2000 13816
rect 0 13744 2000 13784
rect 0 13712 120 13744
rect 152 13712 192 13744
rect 224 13712 264 13744
rect 296 13712 336 13744
rect 368 13712 408 13744
rect 440 13712 480 13744
rect 512 13712 552 13744
rect 584 13712 624 13744
rect 656 13712 696 13744
rect 728 13712 768 13744
rect 800 13712 840 13744
rect 872 13712 912 13744
rect 944 13712 984 13744
rect 1016 13712 1056 13744
rect 1088 13712 1128 13744
rect 1160 13712 1200 13744
rect 1232 13712 1272 13744
rect 1304 13712 1344 13744
rect 1376 13712 1416 13744
rect 1448 13712 1488 13744
rect 1520 13712 1560 13744
rect 1592 13712 1632 13744
rect 1664 13712 1704 13744
rect 1736 13712 1776 13744
rect 1808 13712 1848 13744
rect 1880 13712 2000 13744
rect 0 13672 2000 13712
rect 0 13640 120 13672
rect 152 13640 192 13672
rect 224 13640 264 13672
rect 296 13640 336 13672
rect 368 13640 408 13672
rect 440 13640 480 13672
rect 512 13640 552 13672
rect 584 13640 624 13672
rect 656 13640 696 13672
rect 728 13640 768 13672
rect 800 13640 840 13672
rect 872 13640 912 13672
rect 944 13640 984 13672
rect 1016 13640 1056 13672
rect 1088 13640 1128 13672
rect 1160 13640 1200 13672
rect 1232 13640 1272 13672
rect 1304 13640 1344 13672
rect 1376 13640 1416 13672
rect 1448 13640 1488 13672
rect 1520 13640 1560 13672
rect 1592 13640 1632 13672
rect 1664 13640 1704 13672
rect 1736 13640 1776 13672
rect 1808 13640 1848 13672
rect 1880 13640 2000 13672
rect 0 13600 2000 13640
rect 0 13568 120 13600
rect 152 13568 192 13600
rect 224 13568 264 13600
rect 296 13568 336 13600
rect 368 13568 408 13600
rect 440 13568 480 13600
rect 512 13568 552 13600
rect 584 13568 624 13600
rect 656 13568 696 13600
rect 728 13568 768 13600
rect 800 13568 840 13600
rect 872 13568 912 13600
rect 944 13568 984 13600
rect 1016 13568 1056 13600
rect 1088 13568 1128 13600
rect 1160 13568 1200 13600
rect 1232 13568 1272 13600
rect 1304 13568 1344 13600
rect 1376 13568 1416 13600
rect 1448 13568 1488 13600
rect 1520 13568 1560 13600
rect 1592 13568 1632 13600
rect 1664 13568 1704 13600
rect 1736 13568 1776 13600
rect 1808 13568 1848 13600
rect 1880 13568 2000 13600
rect 0 13528 2000 13568
rect 0 13496 120 13528
rect 152 13496 192 13528
rect 224 13496 264 13528
rect 296 13496 336 13528
rect 368 13496 408 13528
rect 440 13496 480 13528
rect 512 13496 552 13528
rect 584 13496 624 13528
rect 656 13496 696 13528
rect 728 13496 768 13528
rect 800 13496 840 13528
rect 872 13496 912 13528
rect 944 13496 984 13528
rect 1016 13496 1056 13528
rect 1088 13496 1128 13528
rect 1160 13496 1200 13528
rect 1232 13496 1272 13528
rect 1304 13496 1344 13528
rect 1376 13496 1416 13528
rect 1448 13496 1488 13528
rect 1520 13496 1560 13528
rect 1592 13496 1632 13528
rect 1664 13496 1704 13528
rect 1736 13496 1776 13528
rect 1808 13496 1848 13528
rect 1880 13496 2000 13528
rect 0 13456 2000 13496
rect 0 13424 120 13456
rect 152 13424 192 13456
rect 224 13424 264 13456
rect 296 13424 336 13456
rect 368 13424 408 13456
rect 440 13424 480 13456
rect 512 13424 552 13456
rect 584 13424 624 13456
rect 656 13424 696 13456
rect 728 13424 768 13456
rect 800 13424 840 13456
rect 872 13424 912 13456
rect 944 13424 984 13456
rect 1016 13424 1056 13456
rect 1088 13424 1128 13456
rect 1160 13424 1200 13456
rect 1232 13424 1272 13456
rect 1304 13424 1344 13456
rect 1376 13424 1416 13456
rect 1448 13424 1488 13456
rect 1520 13424 1560 13456
rect 1592 13424 1632 13456
rect 1664 13424 1704 13456
rect 1736 13424 1776 13456
rect 1808 13424 1848 13456
rect 1880 13424 2000 13456
rect 0 13384 2000 13424
rect 0 13352 120 13384
rect 152 13352 192 13384
rect 224 13352 264 13384
rect 296 13352 336 13384
rect 368 13352 408 13384
rect 440 13352 480 13384
rect 512 13352 552 13384
rect 584 13352 624 13384
rect 656 13352 696 13384
rect 728 13352 768 13384
rect 800 13352 840 13384
rect 872 13352 912 13384
rect 944 13352 984 13384
rect 1016 13352 1056 13384
rect 1088 13352 1128 13384
rect 1160 13352 1200 13384
rect 1232 13352 1272 13384
rect 1304 13352 1344 13384
rect 1376 13352 1416 13384
rect 1448 13352 1488 13384
rect 1520 13352 1560 13384
rect 1592 13352 1632 13384
rect 1664 13352 1704 13384
rect 1736 13352 1776 13384
rect 1808 13352 1848 13384
rect 1880 13352 2000 13384
rect 0 13312 2000 13352
rect 0 13280 120 13312
rect 152 13280 192 13312
rect 224 13280 264 13312
rect 296 13280 336 13312
rect 368 13280 408 13312
rect 440 13280 480 13312
rect 512 13280 552 13312
rect 584 13280 624 13312
rect 656 13280 696 13312
rect 728 13280 768 13312
rect 800 13280 840 13312
rect 872 13280 912 13312
rect 944 13280 984 13312
rect 1016 13280 1056 13312
rect 1088 13280 1128 13312
rect 1160 13280 1200 13312
rect 1232 13280 1272 13312
rect 1304 13280 1344 13312
rect 1376 13280 1416 13312
rect 1448 13280 1488 13312
rect 1520 13280 1560 13312
rect 1592 13280 1632 13312
rect 1664 13280 1704 13312
rect 1736 13280 1776 13312
rect 1808 13280 1848 13312
rect 1880 13280 2000 13312
rect 0 13240 2000 13280
rect 0 13208 120 13240
rect 152 13208 192 13240
rect 224 13208 264 13240
rect 296 13208 336 13240
rect 368 13208 408 13240
rect 440 13208 480 13240
rect 512 13208 552 13240
rect 584 13208 624 13240
rect 656 13208 696 13240
rect 728 13208 768 13240
rect 800 13208 840 13240
rect 872 13208 912 13240
rect 944 13208 984 13240
rect 1016 13208 1056 13240
rect 1088 13208 1128 13240
rect 1160 13208 1200 13240
rect 1232 13208 1272 13240
rect 1304 13208 1344 13240
rect 1376 13208 1416 13240
rect 1448 13208 1488 13240
rect 1520 13208 1560 13240
rect 1592 13208 1632 13240
rect 1664 13208 1704 13240
rect 1736 13208 1776 13240
rect 1808 13208 1848 13240
rect 1880 13208 2000 13240
rect 0 13168 2000 13208
rect 0 13136 120 13168
rect 152 13136 192 13168
rect 224 13136 264 13168
rect 296 13136 336 13168
rect 368 13136 408 13168
rect 440 13136 480 13168
rect 512 13136 552 13168
rect 584 13136 624 13168
rect 656 13136 696 13168
rect 728 13136 768 13168
rect 800 13136 840 13168
rect 872 13136 912 13168
rect 944 13136 984 13168
rect 1016 13136 1056 13168
rect 1088 13136 1128 13168
rect 1160 13136 1200 13168
rect 1232 13136 1272 13168
rect 1304 13136 1344 13168
rect 1376 13136 1416 13168
rect 1448 13136 1488 13168
rect 1520 13136 1560 13168
rect 1592 13136 1632 13168
rect 1664 13136 1704 13168
rect 1736 13136 1776 13168
rect 1808 13136 1848 13168
rect 1880 13136 2000 13168
rect 0 13096 2000 13136
rect 0 13064 120 13096
rect 152 13064 192 13096
rect 224 13064 264 13096
rect 296 13064 336 13096
rect 368 13064 408 13096
rect 440 13064 480 13096
rect 512 13064 552 13096
rect 584 13064 624 13096
rect 656 13064 696 13096
rect 728 13064 768 13096
rect 800 13064 840 13096
rect 872 13064 912 13096
rect 944 13064 984 13096
rect 1016 13064 1056 13096
rect 1088 13064 1128 13096
rect 1160 13064 1200 13096
rect 1232 13064 1272 13096
rect 1304 13064 1344 13096
rect 1376 13064 1416 13096
rect 1448 13064 1488 13096
rect 1520 13064 1560 13096
rect 1592 13064 1632 13096
rect 1664 13064 1704 13096
rect 1736 13064 1776 13096
rect 1808 13064 1848 13096
rect 1880 13064 2000 13096
rect 0 13000 2000 13064
rect 0 12144 2000 12200
rect 0 12112 48 12144
rect 80 12112 120 12144
rect 152 12112 192 12144
rect 224 12112 264 12144
rect 296 12112 336 12144
rect 368 12112 408 12144
rect 440 12112 480 12144
rect 512 12112 552 12144
rect 584 12112 624 12144
rect 656 12112 696 12144
rect 728 12112 768 12144
rect 800 12112 840 12144
rect 872 12112 912 12144
rect 944 12112 984 12144
rect 1016 12112 1056 12144
rect 1088 12112 1128 12144
rect 1160 12112 1200 12144
rect 1232 12112 1272 12144
rect 1304 12112 1344 12144
rect 1376 12112 1416 12144
rect 1448 12112 1488 12144
rect 1520 12112 1560 12144
rect 1592 12112 1632 12144
rect 1664 12112 1704 12144
rect 1736 12112 1776 12144
rect 1808 12112 1848 12144
rect 1880 12112 1920 12144
rect 1952 12112 2000 12144
rect 0 12072 2000 12112
rect 0 12040 48 12072
rect 80 12040 120 12072
rect 152 12040 192 12072
rect 224 12040 264 12072
rect 296 12040 336 12072
rect 368 12040 408 12072
rect 440 12040 480 12072
rect 512 12040 552 12072
rect 584 12040 624 12072
rect 656 12040 696 12072
rect 728 12040 768 12072
rect 800 12040 840 12072
rect 872 12040 912 12072
rect 944 12040 984 12072
rect 1016 12040 1056 12072
rect 1088 12040 1128 12072
rect 1160 12040 1200 12072
rect 1232 12040 1272 12072
rect 1304 12040 1344 12072
rect 1376 12040 1416 12072
rect 1448 12040 1488 12072
rect 1520 12040 1560 12072
rect 1592 12040 1632 12072
rect 1664 12040 1704 12072
rect 1736 12040 1776 12072
rect 1808 12040 1848 12072
rect 1880 12040 1920 12072
rect 1952 12040 2000 12072
rect 0 12000 2000 12040
rect 0 11968 48 12000
rect 80 11968 120 12000
rect 152 11968 192 12000
rect 224 11968 264 12000
rect 296 11968 336 12000
rect 368 11968 408 12000
rect 440 11968 480 12000
rect 512 11968 552 12000
rect 584 11968 624 12000
rect 656 11968 696 12000
rect 728 11968 768 12000
rect 800 11968 840 12000
rect 872 11968 912 12000
rect 944 11968 984 12000
rect 1016 11968 1056 12000
rect 1088 11968 1128 12000
rect 1160 11968 1200 12000
rect 1232 11968 1272 12000
rect 1304 11968 1344 12000
rect 1376 11968 1416 12000
rect 1448 11968 1488 12000
rect 1520 11968 1560 12000
rect 1592 11968 1632 12000
rect 1664 11968 1704 12000
rect 1736 11968 1776 12000
rect 1808 11968 1848 12000
rect 1880 11968 1920 12000
rect 1952 11968 2000 12000
rect 0 11928 2000 11968
rect 0 11896 48 11928
rect 80 11896 120 11928
rect 152 11896 192 11928
rect 224 11896 264 11928
rect 296 11896 336 11928
rect 368 11896 408 11928
rect 440 11896 480 11928
rect 512 11896 552 11928
rect 584 11896 624 11928
rect 656 11896 696 11928
rect 728 11896 768 11928
rect 800 11896 840 11928
rect 872 11896 912 11928
rect 944 11896 984 11928
rect 1016 11896 1056 11928
rect 1088 11896 1128 11928
rect 1160 11896 1200 11928
rect 1232 11896 1272 11928
rect 1304 11896 1344 11928
rect 1376 11896 1416 11928
rect 1448 11896 1488 11928
rect 1520 11896 1560 11928
rect 1592 11896 1632 11928
rect 1664 11896 1704 11928
rect 1736 11896 1776 11928
rect 1808 11896 1848 11928
rect 1880 11896 1920 11928
rect 1952 11896 2000 11928
rect 0 11856 2000 11896
rect 0 11824 48 11856
rect 80 11824 120 11856
rect 152 11824 192 11856
rect 224 11824 264 11856
rect 296 11824 336 11856
rect 368 11824 408 11856
rect 440 11824 480 11856
rect 512 11824 552 11856
rect 584 11824 624 11856
rect 656 11824 696 11856
rect 728 11824 768 11856
rect 800 11824 840 11856
rect 872 11824 912 11856
rect 944 11824 984 11856
rect 1016 11824 1056 11856
rect 1088 11824 1128 11856
rect 1160 11824 1200 11856
rect 1232 11824 1272 11856
rect 1304 11824 1344 11856
rect 1376 11824 1416 11856
rect 1448 11824 1488 11856
rect 1520 11824 1560 11856
rect 1592 11824 1632 11856
rect 1664 11824 1704 11856
rect 1736 11824 1776 11856
rect 1808 11824 1848 11856
rect 1880 11824 1920 11856
rect 1952 11824 2000 11856
rect 0 11784 2000 11824
rect 0 11752 48 11784
rect 80 11752 120 11784
rect 152 11752 192 11784
rect 224 11752 264 11784
rect 296 11752 336 11784
rect 368 11752 408 11784
rect 440 11752 480 11784
rect 512 11752 552 11784
rect 584 11752 624 11784
rect 656 11752 696 11784
rect 728 11752 768 11784
rect 800 11752 840 11784
rect 872 11752 912 11784
rect 944 11752 984 11784
rect 1016 11752 1056 11784
rect 1088 11752 1128 11784
rect 1160 11752 1200 11784
rect 1232 11752 1272 11784
rect 1304 11752 1344 11784
rect 1376 11752 1416 11784
rect 1448 11752 1488 11784
rect 1520 11752 1560 11784
rect 1592 11752 1632 11784
rect 1664 11752 1704 11784
rect 1736 11752 1776 11784
rect 1808 11752 1848 11784
rect 1880 11752 1920 11784
rect 1952 11752 2000 11784
rect 0 11712 2000 11752
rect 0 11680 48 11712
rect 80 11680 120 11712
rect 152 11680 192 11712
rect 224 11680 264 11712
rect 296 11680 336 11712
rect 368 11680 408 11712
rect 440 11680 480 11712
rect 512 11680 552 11712
rect 584 11680 624 11712
rect 656 11680 696 11712
rect 728 11680 768 11712
rect 800 11680 840 11712
rect 872 11680 912 11712
rect 944 11680 984 11712
rect 1016 11680 1056 11712
rect 1088 11680 1128 11712
rect 1160 11680 1200 11712
rect 1232 11680 1272 11712
rect 1304 11680 1344 11712
rect 1376 11680 1416 11712
rect 1448 11680 1488 11712
rect 1520 11680 1560 11712
rect 1592 11680 1632 11712
rect 1664 11680 1704 11712
rect 1736 11680 1776 11712
rect 1808 11680 1848 11712
rect 1880 11680 1920 11712
rect 1952 11680 2000 11712
rect 0 11640 2000 11680
rect 0 11608 48 11640
rect 80 11608 120 11640
rect 152 11608 192 11640
rect 224 11608 264 11640
rect 296 11608 336 11640
rect 368 11608 408 11640
rect 440 11608 480 11640
rect 512 11608 552 11640
rect 584 11608 624 11640
rect 656 11608 696 11640
rect 728 11608 768 11640
rect 800 11608 840 11640
rect 872 11608 912 11640
rect 944 11608 984 11640
rect 1016 11608 1056 11640
rect 1088 11608 1128 11640
rect 1160 11608 1200 11640
rect 1232 11608 1272 11640
rect 1304 11608 1344 11640
rect 1376 11608 1416 11640
rect 1448 11608 1488 11640
rect 1520 11608 1560 11640
rect 1592 11608 1632 11640
rect 1664 11608 1704 11640
rect 1736 11608 1776 11640
rect 1808 11608 1848 11640
rect 1880 11608 1920 11640
rect 1952 11608 2000 11640
rect 0 11568 2000 11608
rect 0 11536 48 11568
rect 80 11536 120 11568
rect 152 11536 192 11568
rect 224 11536 264 11568
rect 296 11536 336 11568
rect 368 11536 408 11568
rect 440 11536 480 11568
rect 512 11536 552 11568
rect 584 11536 624 11568
rect 656 11536 696 11568
rect 728 11536 768 11568
rect 800 11536 840 11568
rect 872 11536 912 11568
rect 944 11536 984 11568
rect 1016 11536 1056 11568
rect 1088 11536 1128 11568
rect 1160 11536 1200 11568
rect 1232 11536 1272 11568
rect 1304 11536 1344 11568
rect 1376 11536 1416 11568
rect 1448 11536 1488 11568
rect 1520 11536 1560 11568
rect 1592 11536 1632 11568
rect 1664 11536 1704 11568
rect 1736 11536 1776 11568
rect 1808 11536 1848 11568
rect 1880 11536 1920 11568
rect 1952 11536 2000 11568
rect 0 11496 2000 11536
rect 0 11464 48 11496
rect 80 11464 120 11496
rect 152 11464 192 11496
rect 224 11464 264 11496
rect 296 11464 336 11496
rect 368 11464 408 11496
rect 440 11464 480 11496
rect 512 11464 552 11496
rect 584 11464 624 11496
rect 656 11464 696 11496
rect 728 11464 768 11496
rect 800 11464 840 11496
rect 872 11464 912 11496
rect 944 11464 984 11496
rect 1016 11464 1056 11496
rect 1088 11464 1128 11496
rect 1160 11464 1200 11496
rect 1232 11464 1272 11496
rect 1304 11464 1344 11496
rect 1376 11464 1416 11496
rect 1448 11464 1488 11496
rect 1520 11464 1560 11496
rect 1592 11464 1632 11496
rect 1664 11464 1704 11496
rect 1736 11464 1776 11496
rect 1808 11464 1848 11496
rect 1880 11464 1920 11496
rect 1952 11464 2000 11496
rect 0 11424 2000 11464
rect 0 11392 48 11424
rect 80 11392 120 11424
rect 152 11392 192 11424
rect 224 11392 264 11424
rect 296 11392 336 11424
rect 368 11392 408 11424
rect 440 11392 480 11424
rect 512 11392 552 11424
rect 584 11392 624 11424
rect 656 11392 696 11424
rect 728 11392 768 11424
rect 800 11392 840 11424
rect 872 11392 912 11424
rect 944 11392 984 11424
rect 1016 11392 1056 11424
rect 1088 11392 1128 11424
rect 1160 11392 1200 11424
rect 1232 11392 1272 11424
rect 1304 11392 1344 11424
rect 1376 11392 1416 11424
rect 1448 11392 1488 11424
rect 1520 11392 1560 11424
rect 1592 11392 1632 11424
rect 1664 11392 1704 11424
rect 1736 11392 1776 11424
rect 1808 11392 1848 11424
rect 1880 11392 1920 11424
rect 1952 11392 2000 11424
rect 0 11352 2000 11392
rect 0 11320 48 11352
rect 80 11320 120 11352
rect 152 11320 192 11352
rect 224 11320 264 11352
rect 296 11320 336 11352
rect 368 11320 408 11352
rect 440 11320 480 11352
rect 512 11320 552 11352
rect 584 11320 624 11352
rect 656 11320 696 11352
rect 728 11320 768 11352
rect 800 11320 840 11352
rect 872 11320 912 11352
rect 944 11320 984 11352
rect 1016 11320 1056 11352
rect 1088 11320 1128 11352
rect 1160 11320 1200 11352
rect 1232 11320 1272 11352
rect 1304 11320 1344 11352
rect 1376 11320 1416 11352
rect 1448 11320 1488 11352
rect 1520 11320 1560 11352
rect 1592 11320 1632 11352
rect 1664 11320 1704 11352
rect 1736 11320 1776 11352
rect 1808 11320 1848 11352
rect 1880 11320 1920 11352
rect 1952 11320 2000 11352
rect 0 11280 2000 11320
rect 0 11248 48 11280
rect 80 11248 120 11280
rect 152 11248 192 11280
rect 224 11248 264 11280
rect 296 11248 336 11280
rect 368 11248 408 11280
rect 440 11248 480 11280
rect 512 11248 552 11280
rect 584 11248 624 11280
rect 656 11248 696 11280
rect 728 11248 768 11280
rect 800 11248 840 11280
rect 872 11248 912 11280
rect 944 11248 984 11280
rect 1016 11248 1056 11280
rect 1088 11248 1128 11280
rect 1160 11248 1200 11280
rect 1232 11248 1272 11280
rect 1304 11248 1344 11280
rect 1376 11248 1416 11280
rect 1448 11248 1488 11280
rect 1520 11248 1560 11280
rect 1592 11248 1632 11280
rect 1664 11248 1704 11280
rect 1736 11248 1776 11280
rect 1808 11248 1848 11280
rect 1880 11248 1920 11280
rect 1952 11248 2000 11280
rect 0 11208 2000 11248
rect 0 11176 48 11208
rect 80 11176 120 11208
rect 152 11176 192 11208
rect 224 11176 264 11208
rect 296 11176 336 11208
rect 368 11176 408 11208
rect 440 11176 480 11208
rect 512 11176 552 11208
rect 584 11176 624 11208
rect 656 11176 696 11208
rect 728 11176 768 11208
rect 800 11176 840 11208
rect 872 11176 912 11208
rect 944 11176 984 11208
rect 1016 11176 1056 11208
rect 1088 11176 1128 11208
rect 1160 11176 1200 11208
rect 1232 11176 1272 11208
rect 1304 11176 1344 11208
rect 1376 11176 1416 11208
rect 1448 11176 1488 11208
rect 1520 11176 1560 11208
rect 1592 11176 1632 11208
rect 1664 11176 1704 11208
rect 1736 11176 1776 11208
rect 1808 11176 1848 11208
rect 1880 11176 1920 11208
rect 1952 11176 2000 11208
rect 0 11136 2000 11176
rect 0 11104 48 11136
rect 80 11104 120 11136
rect 152 11104 192 11136
rect 224 11104 264 11136
rect 296 11104 336 11136
rect 368 11104 408 11136
rect 440 11104 480 11136
rect 512 11104 552 11136
rect 584 11104 624 11136
rect 656 11104 696 11136
rect 728 11104 768 11136
rect 800 11104 840 11136
rect 872 11104 912 11136
rect 944 11104 984 11136
rect 1016 11104 1056 11136
rect 1088 11104 1128 11136
rect 1160 11104 1200 11136
rect 1232 11104 1272 11136
rect 1304 11104 1344 11136
rect 1376 11104 1416 11136
rect 1448 11104 1488 11136
rect 1520 11104 1560 11136
rect 1592 11104 1632 11136
rect 1664 11104 1704 11136
rect 1736 11104 1776 11136
rect 1808 11104 1848 11136
rect 1880 11104 1920 11136
rect 1952 11104 2000 11136
rect 0 11064 2000 11104
rect 0 11032 48 11064
rect 80 11032 120 11064
rect 152 11032 192 11064
rect 224 11032 264 11064
rect 296 11032 336 11064
rect 368 11032 408 11064
rect 440 11032 480 11064
rect 512 11032 552 11064
rect 584 11032 624 11064
rect 656 11032 696 11064
rect 728 11032 768 11064
rect 800 11032 840 11064
rect 872 11032 912 11064
rect 944 11032 984 11064
rect 1016 11032 1056 11064
rect 1088 11032 1128 11064
rect 1160 11032 1200 11064
rect 1232 11032 1272 11064
rect 1304 11032 1344 11064
rect 1376 11032 1416 11064
rect 1448 11032 1488 11064
rect 1520 11032 1560 11064
rect 1592 11032 1632 11064
rect 1664 11032 1704 11064
rect 1736 11032 1776 11064
rect 1808 11032 1848 11064
rect 1880 11032 1920 11064
rect 1952 11032 2000 11064
rect 0 10992 2000 11032
rect 0 10960 48 10992
rect 80 10960 120 10992
rect 152 10960 192 10992
rect 224 10960 264 10992
rect 296 10960 336 10992
rect 368 10960 408 10992
rect 440 10960 480 10992
rect 512 10960 552 10992
rect 584 10960 624 10992
rect 656 10960 696 10992
rect 728 10960 768 10992
rect 800 10960 840 10992
rect 872 10960 912 10992
rect 944 10960 984 10992
rect 1016 10960 1056 10992
rect 1088 10960 1128 10992
rect 1160 10960 1200 10992
rect 1232 10960 1272 10992
rect 1304 10960 1344 10992
rect 1376 10960 1416 10992
rect 1448 10960 1488 10992
rect 1520 10960 1560 10992
rect 1592 10960 1632 10992
rect 1664 10960 1704 10992
rect 1736 10960 1776 10992
rect 1808 10960 1848 10992
rect 1880 10960 1920 10992
rect 1952 10960 2000 10992
rect 0 10920 2000 10960
rect 0 10888 48 10920
rect 80 10888 120 10920
rect 152 10888 192 10920
rect 224 10888 264 10920
rect 296 10888 336 10920
rect 368 10888 408 10920
rect 440 10888 480 10920
rect 512 10888 552 10920
rect 584 10888 624 10920
rect 656 10888 696 10920
rect 728 10888 768 10920
rect 800 10888 840 10920
rect 872 10888 912 10920
rect 944 10888 984 10920
rect 1016 10888 1056 10920
rect 1088 10888 1128 10920
rect 1160 10888 1200 10920
rect 1232 10888 1272 10920
rect 1304 10888 1344 10920
rect 1376 10888 1416 10920
rect 1448 10888 1488 10920
rect 1520 10888 1560 10920
rect 1592 10888 1632 10920
rect 1664 10888 1704 10920
rect 1736 10888 1776 10920
rect 1808 10888 1848 10920
rect 1880 10888 1920 10920
rect 1952 10888 2000 10920
rect 0 10848 2000 10888
rect 0 10816 48 10848
rect 80 10816 120 10848
rect 152 10816 192 10848
rect 224 10816 264 10848
rect 296 10816 336 10848
rect 368 10816 408 10848
rect 440 10816 480 10848
rect 512 10816 552 10848
rect 584 10816 624 10848
rect 656 10816 696 10848
rect 728 10816 768 10848
rect 800 10816 840 10848
rect 872 10816 912 10848
rect 944 10816 984 10848
rect 1016 10816 1056 10848
rect 1088 10816 1128 10848
rect 1160 10816 1200 10848
rect 1232 10816 1272 10848
rect 1304 10816 1344 10848
rect 1376 10816 1416 10848
rect 1448 10816 1488 10848
rect 1520 10816 1560 10848
rect 1592 10816 1632 10848
rect 1664 10816 1704 10848
rect 1736 10816 1776 10848
rect 1808 10816 1848 10848
rect 1880 10816 1920 10848
rect 1952 10816 2000 10848
rect 0 10776 2000 10816
rect 0 10744 48 10776
rect 80 10744 120 10776
rect 152 10744 192 10776
rect 224 10744 264 10776
rect 296 10744 336 10776
rect 368 10744 408 10776
rect 440 10744 480 10776
rect 512 10744 552 10776
rect 584 10744 624 10776
rect 656 10744 696 10776
rect 728 10744 768 10776
rect 800 10744 840 10776
rect 872 10744 912 10776
rect 944 10744 984 10776
rect 1016 10744 1056 10776
rect 1088 10744 1128 10776
rect 1160 10744 1200 10776
rect 1232 10744 1272 10776
rect 1304 10744 1344 10776
rect 1376 10744 1416 10776
rect 1448 10744 1488 10776
rect 1520 10744 1560 10776
rect 1592 10744 1632 10776
rect 1664 10744 1704 10776
rect 1736 10744 1776 10776
rect 1808 10744 1848 10776
rect 1880 10744 1920 10776
rect 1952 10744 2000 10776
rect 0 10704 2000 10744
rect 0 10672 48 10704
rect 80 10672 120 10704
rect 152 10672 192 10704
rect 224 10672 264 10704
rect 296 10672 336 10704
rect 368 10672 408 10704
rect 440 10672 480 10704
rect 512 10672 552 10704
rect 584 10672 624 10704
rect 656 10672 696 10704
rect 728 10672 768 10704
rect 800 10672 840 10704
rect 872 10672 912 10704
rect 944 10672 984 10704
rect 1016 10672 1056 10704
rect 1088 10672 1128 10704
rect 1160 10672 1200 10704
rect 1232 10672 1272 10704
rect 1304 10672 1344 10704
rect 1376 10672 1416 10704
rect 1448 10672 1488 10704
rect 1520 10672 1560 10704
rect 1592 10672 1632 10704
rect 1664 10672 1704 10704
rect 1736 10672 1776 10704
rect 1808 10672 1848 10704
rect 1880 10672 1920 10704
rect 1952 10672 2000 10704
rect 0 10632 2000 10672
rect 0 10600 48 10632
rect 80 10600 120 10632
rect 152 10600 192 10632
rect 224 10600 264 10632
rect 296 10600 336 10632
rect 368 10600 408 10632
rect 440 10600 480 10632
rect 512 10600 552 10632
rect 584 10600 624 10632
rect 656 10600 696 10632
rect 728 10600 768 10632
rect 800 10600 840 10632
rect 872 10600 912 10632
rect 944 10600 984 10632
rect 1016 10600 1056 10632
rect 1088 10600 1128 10632
rect 1160 10600 1200 10632
rect 1232 10600 1272 10632
rect 1304 10600 1344 10632
rect 1376 10600 1416 10632
rect 1448 10600 1488 10632
rect 1520 10600 1560 10632
rect 1592 10600 1632 10632
rect 1664 10600 1704 10632
rect 1736 10600 1776 10632
rect 1808 10600 1848 10632
rect 1880 10600 1920 10632
rect 1952 10600 2000 10632
rect 0 10560 2000 10600
rect 0 10528 48 10560
rect 80 10528 120 10560
rect 152 10528 192 10560
rect 224 10528 264 10560
rect 296 10528 336 10560
rect 368 10528 408 10560
rect 440 10528 480 10560
rect 512 10528 552 10560
rect 584 10528 624 10560
rect 656 10528 696 10560
rect 728 10528 768 10560
rect 800 10528 840 10560
rect 872 10528 912 10560
rect 944 10528 984 10560
rect 1016 10528 1056 10560
rect 1088 10528 1128 10560
rect 1160 10528 1200 10560
rect 1232 10528 1272 10560
rect 1304 10528 1344 10560
rect 1376 10528 1416 10560
rect 1448 10528 1488 10560
rect 1520 10528 1560 10560
rect 1592 10528 1632 10560
rect 1664 10528 1704 10560
rect 1736 10528 1776 10560
rect 1808 10528 1848 10560
rect 1880 10528 1920 10560
rect 1952 10528 2000 10560
rect 0 10488 2000 10528
rect 0 10456 48 10488
rect 80 10456 120 10488
rect 152 10456 192 10488
rect 224 10456 264 10488
rect 296 10456 336 10488
rect 368 10456 408 10488
rect 440 10456 480 10488
rect 512 10456 552 10488
rect 584 10456 624 10488
rect 656 10456 696 10488
rect 728 10456 768 10488
rect 800 10456 840 10488
rect 872 10456 912 10488
rect 944 10456 984 10488
rect 1016 10456 1056 10488
rect 1088 10456 1128 10488
rect 1160 10456 1200 10488
rect 1232 10456 1272 10488
rect 1304 10456 1344 10488
rect 1376 10456 1416 10488
rect 1448 10456 1488 10488
rect 1520 10456 1560 10488
rect 1592 10456 1632 10488
rect 1664 10456 1704 10488
rect 1736 10456 1776 10488
rect 1808 10456 1848 10488
rect 1880 10456 1920 10488
rect 1952 10456 2000 10488
rect 0 10416 2000 10456
rect 0 10384 48 10416
rect 80 10384 120 10416
rect 152 10384 192 10416
rect 224 10384 264 10416
rect 296 10384 336 10416
rect 368 10384 408 10416
rect 440 10384 480 10416
rect 512 10384 552 10416
rect 584 10384 624 10416
rect 656 10384 696 10416
rect 728 10384 768 10416
rect 800 10384 840 10416
rect 872 10384 912 10416
rect 944 10384 984 10416
rect 1016 10384 1056 10416
rect 1088 10384 1128 10416
rect 1160 10384 1200 10416
rect 1232 10384 1272 10416
rect 1304 10384 1344 10416
rect 1376 10384 1416 10416
rect 1448 10384 1488 10416
rect 1520 10384 1560 10416
rect 1592 10384 1632 10416
rect 1664 10384 1704 10416
rect 1736 10384 1776 10416
rect 1808 10384 1848 10416
rect 1880 10384 1920 10416
rect 1952 10384 2000 10416
rect 0 10344 2000 10384
rect 0 10312 48 10344
rect 80 10312 120 10344
rect 152 10312 192 10344
rect 224 10312 264 10344
rect 296 10312 336 10344
rect 368 10312 408 10344
rect 440 10312 480 10344
rect 512 10312 552 10344
rect 584 10312 624 10344
rect 656 10312 696 10344
rect 728 10312 768 10344
rect 800 10312 840 10344
rect 872 10312 912 10344
rect 944 10312 984 10344
rect 1016 10312 1056 10344
rect 1088 10312 1128 10344
rect 1160 10312 1200 10344
rect 1232 10312 1272 10344
rect 1304 10312 1344 10344
rect 1376 10312 1416 10344
rect 1448 10312 1488 10344
rect 1520 10312 1560 10344
rect 1592 10312 1632 10344
rect 1664 10312 1704 10344
rect 1736 10312 1776 10344
rect 1808 10312 1848 10344
rect 1880 10312 1920 10344
rect 1952 10312 2000 10344
rect 0 10272 2000 10312
rect 0 10240 48 10272
rect 80 10240 120 10272
rect 152 10240 192 10272
rect 224 10240 264 10272
rect 296 10240 336 10272
rect 368 10240 408 10272
rect 440 10240 480 10272
rect 512 10240 552 10272
rect 584 10240 624 10272
rect 656 10240 696 10272
rect 728 10240 768 10272
rect 800 10240 840 10272
rect 872 10240 912 10272
rect 944 10240 984 10272
rect 1016 10240 1056 10272
rect 1088 10240 1128 10272
rect 1160 10240 1200 10272
rect 1232 10240 1272 10272
rect 1304 10240 1344 10272
rect 1376 10240 1416 10272
rect 1448 10240 1488 10272
rect 1520 10240 1560 10272
rect 1592 10240 1632 10272
rect 1664 10240 1704 10272
rect 1736 10240 1776 10272
rect 1808 10240 1848 10272
rect 1880 10240 1920 10272
rect 1952 10240 2000 10272
rect 0 10200 2000 10240
rect 0 10168 48 10200
rect 80 10168 120 10200
rect 152 10168 192 10200
rect 224 10168 264 10200
rect 296 10168 336 10200
rect 368 10168 408 10200
rect 440 10168 480 10200
rect 512 10168 552 10200
rect 584 10168 624 10200
rect 656 10168 696 10200
rect 728 10168 768 10200
rect 800 10168 840 10200
rect 872 10168 912 10200
rect 944 10168 984 10200
rect 1016 10168 1056 10200
rect 1088 10168 1128 10200
rect 1160 10168 1200 10200
rect 1232 10168 1272 10200
rect 1304 10168 1344 10200
rect 1376 10168 1416 10200
rect 1448 10168 1488 10200
rect 1520 10168 1560 10200
rect 1592 10168 1632 10200
rect 1664 10168 1704 10200
rect 1736 10168 1776 10200
rect 1808 10168 1848 10200
rect 1880 10168 1920 10200
rect 1952 10168 2000 10200
rect 0 10128 2000 10168
rect 0 10096 48 10128
rect 80 10096 120 10128
rect 152 10096 192 10128
rect 224 10096 264 10128
rect 296 10096 336 10128
rect 368 10096 408 10128
rect 440 10096 480 10128
rect 512 10096 552 10128
rect 584 10096 624 10128
rect 656 10096 696 10128
rect 728 10096 768 10128
rect 800 10096 840 10128
rect 872 10096 912 10128
rect 944 10096 984 10128
rect 1016 10096 1056 10128
rect 1088 10096 1128 10128
rect 1160 10096 1200 10128
rect 1232 10096 1272 10128
rect 1304 10096 1344 10128
rect 1376 10096 1416 10128
rect 1448 10096 1488 10128
rect 1520 10096 1560 10128
rect 1592 10096 1632 10128
rect 1664 10096 1704 10128
rect 1736 10096 1776 10128
rect 1808 10096 1848 10128
rect 1880 10096 1920 10128
rect 1952 10096 2000 10128
rect 0 10056 2000 10096
rect 0 10024 48 10056
rect 80 10024 120 10056
rect 152 10024 192 10056
rect 224 10024 264 10056
rect 296 10024 336 10056
rect 368 10024 408 10056
rect 440 10024 480 10056
rect 512 10024 552 10056
rect 584 10024 624 10056
rect 656 10024 696 10056
rect 728 10024 768 10056
rect 800 10024 840 10056
rect 872 10024 912 10056
rect 944 10024 984 10056
rect 1016 10024 1056 10056
rect 1088 10024 1128 10056
rect 1160 10024 1200 10056
rect 1232 10024 1272 10056
rect 1304 10024 1344 10056
rect 1376 10024 1416 10056
rect 1448 10024 1488 10056
rect 1520 10024 1560 10056
rect 1592 10024 1632 10056
rect 1664 10024 1704 10056
rect 1736 10024 1776 10056
rect 1808 10024 1848 10056
rect 1880 10024 1920 10056
rect 1952 10024 2000 10056
rect 0 9984 2000 10024
rect 0 9952 48 9984
rect 80 9952 120 9984
rect 152 9952 192 9984
rect 224 9952 264 9984
rect 296 9952 336 9984
rect 368 9952 408 9984
rect 440 9952 480 9984
rect 512 9952 552 9984
rect 584 9952 624 9984
rect 656 9952 696 9984
rect 728 9952 768 9984
rect 800 9952 840 9984
rect 872 9952 912 9984
rect 944 9952 984 9984
rect 1016 9952 1056 9984
rect 1088 9952 1128 9984
rect 1160 9952 1200 9984
rect 1232 9952 1272 9984
rect 1304 9952 1344 9984
rect 1376 9952 1416 9984
rect 1448 9952 1488 9984
rect 1520 9952 1560 9984
rect 1592 9952 1632 9984
rect 1664 9952 1704 9984
rect 1736 9952 1776 9984
rect 1808 9952 1848 9984
rect 1880 9952 1920 9984
rect 1952 9952 2000 9984
rect 0 9912 2000 9952
rect 0 9880 48 9912
rect 80 9880 120 9912
rect 152 9880 192 9912
rect 224 9880 264 9912
rect 296 9880 336 9912
rect 368 9880 408 9912
rect 440 9880 480 9912
rect 512 9880 552 9912
rect 584 9880 624 9912
rect 656 9880 696 9912
rect 728 9880 768 9912
rect 800 9880 840 9912
rect 872 9880 912 9912
rect 944 9880 984 9912
rect 1016 9880 1056 9912
rect 1088 9880 1128 9912
rect 1160 9880 1200 9912
rect 1232 9880 1272 9912
rect 1304 9880 1344 9912
rect 1376 9880 1416 9912
rect 1448 9880 1488 9912
rect 1520 9880 1560 9912
rect 1592 9880 1632 9912
rect 1664 9880 1704 9912
rect 1736 9880 1776 9912
rect 1808 9880 1848 9912
rect 1880 9880 1920 9912
rect 1952 9880 2000 9912
rect 0 9840 2000 9880
rect 0 9808 48 9840
rect 80 9808 120 9840
rect 152 9808 192 9840
rect 224 9808 264 9840
rect 296 9808 336 9840
rect 368 9808 408 9840
rect 440 9808 480 9840
rect 512 9808 552 9840
rect 584 9808 624 9840
rect 656 9808 696 9840
rect 728 9808 768 9840
rect 800 9808 840 9840
rect 872 9808 912 9840
rect 944 9808 984 9840
rect 1016 9808 1056 9840
rect 1088 9808 1128 9840
rect 1160 9808 1200 9840
rect 1232 9808 1272 9840
rect 1304 9808 1344 9840
rect 1376 9808 1416 9840
rect 1448 9808 1488 9840
rect 1520 9808 1560 9840
rect 1592 9808 1632 9840
rect 1664 9808 1704 9840
rect 1736 9808 1776 9840
rect 1808 9808 1848 9840
rect 1880 9808 1920 9840
rect 1952 9808 2000 9840
rect 0 9768 2000 9808
rect 0 9736 48 9768
rect 80 9736 120 9768
rect 152 9736 192 9768
rect 224 9736 264 9768
rect 296 9736 336 9768
rect 368 9736 408 9768
rect 440 9736 480 9768
rect 512 9736 552 9768
rect 584 9736 624 9768
rect 656 9736 696 9768
rect 728 9736 768 9768
rect 800 9736 840 9768
rect 872 9736 912 9768
rect 944 9736 984 9768
rect 1016 9736 1056 9768
rect 1088 9736 1128 9768
rect 1160 9736 1200 9768
rect 1232 9736 1272 9768
rect 1304 9736 1344 9768
rect 1376 9736 1416 9768
rect 1448 9736 1488 9768
rect 1520 9736 1560 9768
rect 1592 9736 1632 9768
rect 1664 9736 1704 9768
rect 1736 9736 1776 9768
rect 1808 9736 1848 9768
rect 1880 9736 1920 9768
rect 1952 9736 2000 9768
rect 0 9696 2000 9736
rect 0 9664 48 9696
rect 80 9664 120 9696
rect 152 9664 192 9696
rect 224 9664 264 9696
rect 296 9664 336 9696
rect 368 9664 408 9696
rect 440 9664 480 9696
rect 512 9664 552 9696
rect 584 9664 624 9696
rect 656 9664 696 9696
rect 728 9664 768 9696
rect 800 9664 840 9696
rect 872 9664 912 9696
rect 944 9664 984 9696
rect 1016 9664 1056 9696
rect 1088 9664 1128 9696
rect 1160 9664 1200 9696
rect 1232 9664 1272 9696
rect 1304 9664 1344 9696
rect 1376 9664 1416 9696
rect 1448 9664 1488 9696
rect 1520 9664 1560 9696
rect 1592 9664 1632 9696
rect 1664 9664 1704 9696
rect 1736 9664 1776 9696
rect 1808 9664 1848 9696
rect 1880 9664 1920 9696
rect 1952 9664 2000 9696
rect 0 9624 2000 9664
rect 0 9592 48 9624
rect 80 9592 120 9624
rect 152 9592 192 9624
rect 224 9592 264 9624
rect 296 9592 336 9624
rect 368 9592 408 9624
rect 440 9592 480 9624
rect 512 9592 552 9624
rect 584 9592 624 9624
rect 656 9592 696 9624
rect 728 9592 768 9624
rect 800 9592 840 9624
rect 872 9592 912 9624
rect 944 9592 984 9624
rect 1016 9592 1056 9624
rect 1088 9592 1128 9624
rect 1160 9592 1200 9624
rect 1232 9592 1272 9624
rect 1304 9592 1344 9624
rect 1376 9592 1416 9624
rect 1448 9592 1488 9624
rect 1520 9592 1560 9624
rect 1592 9592 1632 9624
rect 1664 9592 1704 9624
rect 1736 9592 1776 9624
rect 1808 9592 1848 9624
rect 1880 9592 1920 9624
rect 1952 9592 2000 9624
rect 0 9552 2000 9592
rect 0 9520 48 9552
rect 80 9520 120 9552
rect 152 9520 192 9552
rect 224 9520 264 9552
rect 296 9520 336 9552
rect 368 9520 408 9552
rect 440 9520 480 9552
rect 512 9520 552 9552
rect 584 9520 624 9552
rect 656 9520 696 9552
rect 728 9520 768 9552
rect 800 9520 840 9552
rect 872 9520 912 9552
rect 944 9520 984 9552
rect 1016 9520 1056 9552
rect 1088 9520 1128 9552
rect 1160 9520 1200 9552
rect 1232 9520 1272 9552
rect 1304 9520 1344 9552
rect 1376 9520 1416 9552
rect 1448 9520 1488 9552
rect 1520 9520 1560 9552
rect 1592 9520 1632 9552
rect 1664 9520 1704 9552
rect 1736 9520 1776 9552
rect 1808 9520 1848 9552
rect 1880 9520 1920 9552
rect 1952 9520 2000 9552
rect 0 9480 2000 9520
rect 0 9448 48 9480
rect 80 9448 120 9480
rect 152 9448 192 9480
rect 224 9448 264 9480
rect 296 9448 336 9480
rect 368 9448 408 9480
rect 440 9448 480 9480
rect 512 9448 552 9480
rect 584 9448 624 9480
rect 656 9448 696 9480
rect 728 9448 768 9480
rect 800 9448 840 9480
rect 872 9448 912 9480
rect 944 9448 984 9480
rect 1016 9448 1056 9480
rect 1088 9448 1128 9480
rect 1160 9448 1200 9480
rect 1232 9448 1272 9480
rect 1304 9448 1344 9480
rect 1376 9448 1416 9480
rect 1448 9448 1488 9480
rect 1520 9448 1560 9480
rect 1592 9448 1632 9480
rect 1664 9448 1704 9480
rect 1736 9448 1776 9480
rect 1808 9448 1848 9480
rect 1880 9448 1920 9480
rect 1952 9448 2000 9480
rect 0 9408 2000 9448
rect 0 9376 48 9408
rect 80 9376 120 9408
rect 152 9376 192 9408
rect 224 9376 264 9408
rect 296 9376 336 9408
rect 368 9376 408 9408
rect 440 9376 480 9408
rect 512 9376 552 9408
rect 584 9376 624 9408
rect 656 9376 696 9408
rect 728 9376 768 9408
rect 800 9376 840 9408
rect 872 9376 912 9408
rect 944 9376 984 9408
rect 1016 9376 1056 9408
rect 1088 9376 1128 9408
rect 1160 9376 1200 9408
rect 1232 9376 1272 9408
rect 1304 9376 1344 9408
rect 1376 9376 1416 9408
rect 1448 9376 1488 9408
rect 1520 9376 1560 9408
rect 1592 9376 1632 9408
rect 1664 9376 1704 9408
rect 1736 9376 1776 9408
rect 1808 9376 1848 9408
rect 1880 9376 1920 9408
rect 1952 9376 2000 9408
rect 0 9336 2000 9376
rect 0 9304 48 9336
rect 80 9304 120 9336
rect 152 9304 192 9336
rect 224 9304 264 9336
rect 296 9304 336 9336
rect 368 9304 408 9336
rect 440 9304 480 9336
rect 512 9304 552 9336
rect 584 9304 624 9336
rect 656 9304 696 9336
rect 728 9304 768 9336
rect 800 9304 840 9336
rect 872 9304 912 9336
rect 944 9304 984 9336
rect 1016 9304 1056 9336
rect 1088 9304 1128 9336
rect 1160 9304 1200 9336
rect 1232 9304 1272 9336
rect 1304 9304 1344 9336
rect 1376 9304 1416 9336
rect 1448 9304 1488 9336
rect 1520 9304 1560 9336
rect 1592 9304 1632 9336
rect 1664 9304 1704 9336
rect 1736 9304 1776 9336
rect 1808 9304 1848 9336
rect 1880 9304 1920 9336
rect 1952 9304 2000 9336
rect 0 9264 2000 9304
rect 0 9232 48 9264
rect 80 9232 120 9264
rect 152 9232 192 9264
rect 224 9232 264 9264
rect 296 9232 336 9264
rect 368 9232 408 9264
rect 440 9232 480 9264
rect 512 9232 552 9264
rect 584 9232 624 9264
rect 656 9232 696 9264
rect 728 9232 768 9264
rect 800 9232 840 9264
rect 872 9232 912 9264
rect 944 9232 984 9264
rect 1016 9232 1056 9264
rect 1088 9232 1128 9264
rect 1160 9232 1200 9264
rect 1232 9232 1272 9264
rect 1304 9232 1344 9264
rect 1376 9232 1416 9264
rect 1448 9232 1488 9264
rect 1520 9232 1560 9264
rect 1592 9232 1632 9264
rect 1664 9232 1704 9264
rect 1736 9232 1776 9264
rect 1808 9232 1848 9264
rect 1880 9232 1920 9264
rect 1952 9232 2000 9264
rect 0 9192 2000 9232
rect 0 9160 48 9192
rect 80 9160 120 9192
rect 152 9160 192 9192
rect 224 9160 264 9192
rect 296 9160 336 9192
rect 368 9160 408 9192
rect 440 9160 480 9192
rect 512 9160 552 9192
rect 584 9160 624 9192
rect 656 9160 696 9192
rect 728 9160 768 9192
rect 800 9160 840 9192
rect 872 9160 912 9192
rect 944 9160 984 9192
rect 1016 9160 1056 9192
rect 1088 9160 1128 9192
rect 1160 9160 1200 9192
rect 1232 9160 1272 9192
rect 1304 9160 1344 9192
rect 1376 9160 1416 9192
rect 1448 9160 1488 9192
rect 1520 9160 1560 9192
rect 1592 9160 1632 9192
rect 1664 9160 1704 9192
rect 1736 9160 1776 9192
rect 1808 9160 1848 9192
rect 1880 9160 1920 9192
rect 1952 9160 2000 9192
rect 0 9120 2000 9160
rect 0 9088 48 9120
rect 80 9088 120 9120
rect 152 9088 192 9120
rect 224 9088 264 9120
rect 296 9088 336 9120
rect 368 9088 408 9120
rect 440 9088 480 9120
rect 512 9088 552 9120
rect 584 9088 624 9120
rect 656 9088 696 9120
rect 728 9088 768 9120
rect 800 9088 840 9120
rect 872 9088 912 9120
rect 944 9088 984 9120
rect 1016 9088 1056 9120
rect 1088 9088 1128 9120
rect 1160 9088 1200 9120
rect 1232 9088 1272 9120
rect 1304 9088 1344 9120
rect 1376 9088 1416 9120
rect 1448 9088 1488 9120
rect 1520 9088 1560 9120
rect 1592 9088 1632 9120
rect 1664 9088 1704 9120
rect 1736 9088 1776 9120
rect 1808 9088 1848 9120
rect 1880 9088 1920 9120
rect 1952 9088 2000 9120
rect 0 9048 2000 9088
rect 0 9016 48 9048
rect 80 9016 120 9048
rect 152 9016 192 9048
rect 224 9016 264 9048
rect 296 9016 336 9048
rect 368 9016 408 9048
rect 440 9016 480 9048
rect 512 9016 552 9048
rect 584 9016 624 9048
rect 656 9016 696 9048
rect 728 9016 768 9048
rect 800 9016 840 9048
rect 872 9016 912 9048
rect 944 9016 984 9048
rect 1016 9016 1056 9048
rect 1088 9016 1128 9048
rect 1160 9016 1200 9048
rect 1232 9016 1272 9048
rect 1304 9016 1344 9048
rect 1376 9016 1416 9048
rect 1448 9016 1488 9048
rect 1520 9016 1560 9048
rect 1592 9016 1632 9048
rect 1664 9016 1704 9048
rect 1736 9016 1776 9048
rect 1808 9016 1848 9048
rect 1880 9016 1920 9048
rect 1952 9016 2000 9048
rect 0 8976 2000 9016
rect 0 8944 48 8976
rect 80 8944 120 8976
rect 152 8944 192 8976
rect 224 8944 264 8976
rect 296 8944 336 8976
rect 368 8944 408 8976
rect 440 8944 480 8976
rect 512 8944 552 8976
rect 584 8944 624 8976
rect 656 8944 696 8976
rect 728 8944 768 8976
rect 800 8944 840 8976
rect 872 8944 912 8976
rect 944 8944 984 8976
rect 1016 8944 1056 8976
rect 1088 8944 1128 8976
rect 1160 8944 1200 8976
rect 1232 8944 1272 8976
rect 1304 8944 1344 8976
rect 1376 8944 1416 8976
rect 1448 8944 1488 8976
rect 1520 8944 1560 8976
rect 1592 8944 1632 8976
rect 1664 8944 1704 8976
rect 1736 8944 1776 8976
rect 1808 8944 1848 8976
rect 1880 8944 1920 8976
rect 1952 8944 2000 8976
rect 0 8904 2000 8944
rect 0 8872 48 8904
rect 80 8872 120 8904
rect 152 8872 192 8904
rect 224 8872 264 8904
rect 296 8872 336 8904
rect 368 8872 408 8904
rect 440 8872 480 8904
rect 512 8872 552 8904
rect 584 8872 624 8904
rect 656 8872 696 8904
rect 728 8872 768 8904
rect 800 8872 840 8904
rect 872 8872 912 8904
rect 944 8872 984 8904
rect 1016 8872 1056 8904
rect 1088 8872 1128 8904
rect 1160 8872 1200 8904
rect 1232 8872 1272 8904
rect 1304 8872 1344 8904
rect 1376 8872 1416 8904
rect 1448 8872 1488 8904
rect 1520 8872 1560 8904
rect 1592 8872 1632 8904
rect 1664 8872 1704 8904
rect 1736 8872 1776 8904
rect 1808 8872 1848 8904
rect 1880 8872 1920 8904
rect 1952 8872 2000 8904
rect 0 8832 2000 8872
rect 0 8800 48 8832
rect 80 8800 120 8832
rect 152 8800 192 8832
rect 224 8800 264 8832
rect 296 8800 336 8832
rect 368 8800 408 8832
rect 440 8800 480 8832
rect 512 8800 552 8832
rect 584 8800 624 8832
rect 656 8800 696 8832
rect 728 8800 768 8832
rect 800 8800 840 8832
rect 872 8800 912 8832
rect 944 8800 984 8832
rect 1016 8800 1056 8832
rect 1088 8800 1128 8832
rect 1160 8800 1200 8832
rect 1232 8800 1272 8832
rect 1304 8800 1344 8832
rect 1376 8800 1416 8832
rect 1448 8800 1488 8832
rect 1520 8800 1560 8832
rect 1592 8800 1632 8832
rect 1664 8800 1704 8832
rect 1736 8800 1776 8832
rect 1808 8800 1848 8832
rect 1880 8800 1920 8832
rect 1952 8800 2000 8832
rect 0 8760 2000 8800
rect 0 8728 48 8760
rect 80 8728 120 8760
rect 152 8728 192 8760
rect 224 8728 264 8760
rect 296 8728 336 8760
rect 368 8728 408 8760
rect 440 8728 480 8760
rect 512 8728 552 8760
rect 584 8728 624 8760
rect 656 8728 696 8760
rect 728 8728 768 8760
rect 800 8728 840 8760
rect 872 8728 912 8760
rect 944 8728 984 8760
rect 1016 8728 1056 8760
rect 1088 8728 1128 8760
rect 1160 8728 1200 8760
rect 1232 8728 1272 8760
rect 1304 8728 1344 8760
rect 1376 8728 1416 8760
rect 1448 8728 1488 8760
rect 1520 8728 1560 8760
rect 1592 8728 1632 8760
rect 1664 8728 1704 8760
rect 1736 8728 1776 8760
rect 1808 8728 1848 8760
rect 1880 8728 1920 8760
rect 1952 8728 2000 8760
rect 0 8688 2000 8728
rect 0 8656 48 8688
rect 80 8656 120 8688
rect 152 8656 192 8688
rect 224 8656 264 8688
rect 296 8656 336 8688
rect 368 8656 408 8688
rect 440 8656 480 8688
rect 512 8656 552 8688
rect 584 8656 624 8688
rect 656 8656 696 8688
rect 728 8656 768 8688
rect 800 8656 840 8688
rect 872 8656 912 8688
rect 944 8656 984 8688
rect 1016 8656 1056 8688
rect 1088 8656 1128 8688
rect 1160 8656 1200 8688
rect 1232 8656 1272 8688
rect 1304 8656 1344 8688
rect 1376 8656 1416 8688
rect 1448 8656 1488 8688
rect 1520 8656 1560 8688
rect 1592 8656 1632 8688
rect 1664 8656 1704 8688
rect 1736 8656 1776 8688
rect 1808 8656 1848 8688
rect 1880 8656 1920 8688
rect 1952 8656 2000 8688
rect 0 8616 2000 8656
rect 0 8584 48 8616
rect 80 8584 120 8616
rect 152 8584 192 8616
rect 224 8584 264 8616
rect 296 8584 336 8616
rect 368 8584 408 8616
rect 440 8584 480 8616
rect 512 8584 552 8616
rect 584 8584 624 8616
rect 656 8584 696 8616
rect 728 8584 768 8616
rect 800 8584 840 8616
rect 872 8584 912 8616
rect 944 8584 984 8616
rect 1016 8584 1056 8616
rect 1088 8584 1128 8616
rect 1160 8584 1200 8616
rect 1232 8584 1272 8616
rect 1304 8584 1344 8616
rect 1376 8584 1416 8616
rect 1448 8584 1488 8616
rect 1520 8584 1560 8616
rect 1592 8584 1632 8616
rect 1664 8584 1704 8616
rect 1736 8584 1776 8616
rect 1808 8584 1848 8616
rect 1880 8584 1920 8616
rect 1952 8584 2000 8616
rect 0 8544 2000 8584
rect 0 8512 48 8544
rect 80 8512 120 8544
rect 152 8512 192 8544
rect 224 8512 264 8544
rect 296 8512 336 8544
rect 368 8512 408 8544
rect 440 8512 480 8544
rect 512 8512 552 8544
rect 584 8512 624 8544
rect 656 8512 696 8544
rect 728 8512 768 8544
rect 800 8512 840 8544
rect 872 8512 912 8544
rect 944 8512 984 8544
rect 1016 8512 1056 8544
rect 1088 8512 1128 8544
rect 1160 8512 1200 8544
rect 1232 8512 1272 8544
rect 1304 8512 1344 8544
rect 1376 8512 1416 8544
rect 1448 8512 1488 8544
rect 1520 8512 1560 8544
rect 1592 8512 1632 8544
rect 1664 8512 1704 8544
rect 1736 8512 1776 8544
rect 1808 8512 1848 8544
rect 1880 8512 1920 8544
rect 1952 8512 2000 8544
rect 0 8472 2000 8512
rect 0 8440 48 8472
rect 80 8440 120 8472
rect 152 8440 192 8472
rect 224 8440 264 8472
rect 296 8440 336 8472
rect 368 8440 408 8472
rect 440 8440 480 8472
rect 512 8440 552 8472
rect 584 8440 624 8472
rect 656 8440 696 8472
rect 728 8440 768 8472
rect 800 8440 840 8472
rect 872 8440 912 8472
rect 944 8440 984 8472
rect 1016 8440 1056 8472
rect 1088 8440 1128 8472
rect 1160 8440 1200 8472
rect 1232 8440 1272 8472
rect 1304 8440 1344 8472
rect 1376 8440 1416 8472
rect 1448 8440 1488 8472
rect 1520 8440 1560 8472
rect 1592 8440 1632 8472
rect 1664 8440 1704 8472
rect 1736 8440 1776 8472
rect 1808 8440 1848 8472
rect 1880 8440 1920 8472
rect 1952 8440 2000 8472
rect 0 8400 2000 8440
rect 0 8368 48 8400
rect 80 8368 120 8400
rect 152 8368 192 8400
rect 224 8368 264 8400
rect 296 8368 336 8400
rect 368 8368 408 8400
rect 440 8368 480 8400
rect 512 8368 552 8400
rect 584 8368 624 8400
rect 656 8368 696 8400
rect 728 8368 768 8400
rect 800 8368 840 8400
rect 872 8368 912 8400
rect 944 8368 984 8400
rect 1016 8368 1056 8400
rect 1088 8368 1128 8400
rect 1160 8368 1200 8400
rect 1232 8368 1272 8400
rect 1304 8368 1344 8400
rect 1376 8368 1416 8400
rect 1448 8368 1488 8400
rect 1520 8368 1560 8400
rect 1592 8368 1632 8400
rect 1664 8368 1704 8400
rect 1736 8368 1776 8400
rect 1808 8368 1848 8400
rect 1880 8368 1920 8400
rect 1952 8368 2000 8400
rect 0 8328 2000 8368
rect 0 8296 48 8328
rect 80 8296 120 8328
rect 152 8296 192 8328
rect 224 8296 264 8328
rect 296 8296 336 8328
rect 368 8296 408 8328
rect 440 8296 480 8328
rect 512 8296 552 8328
rect 584 8296 624 8328
rect 656 8296 696 8328
rect 728 8296 768 8328
rect 800 8296 840 8328
rect 872 8296 912 8328
rect 944 8296 984 8328
rect 1016 8296 1056 8328
rect 1088 8296 1128 8328
rect 1160 8296 1200 8328
rect 1232 8296 1272 8328
rect 1304 8296 1344 8328
rect 1376 8296 1416 8328
rect 1448 8296 1488 8328
rect 1520 8296 1560 8328
rect 1592 8296 1632 8328
rect 1664 8296 1704 8328
rect 1736 8296 1776 8328
rect 1808 8296 1848 8328
rect 1880 8296 1920 8328
rect 1952 8296 2000 8328
rect 0 8256 2000 8296
rect 0 8224 48 8256
rect 80 8224 120 8256
rect 152 8224 192 8256
rect 224 8224 264 8256
rect 296 8224 336 8256
rect 368 8224 408 8256
rect 440 8224 480 8256
rect 512 8224 552 8256
rect 584 8224 624 8256
rect 656 8224 696 8256
rect 728 8224 768 8256
rect 800 8224 840 8256
rect 872 8224 912 8256
rect 944 8224 984 8256
rect 1016 8224 1056 8256
rect 1088 8224 1128 8256
rect 1160 8224 1200 8256
rect 1232 8224 1272 8256
rect 1304 8224 1344 8256
rect 1376 8224 1416 8256
rect 1448 8224 1488 8256
rect 1520 8224 1560 8256
rect 1592 8224 1632 8256
rect 1664 8224 1704 8256
rect 1736 8224 1776 8256
rect 1808 8224 1848 8256
rect 1880 8224 1920 8256
rect 1952 8224 2000 8256
rect 0 8184 2000 8224
rect 0 8152 48 8184
rect 80 8152 120 8184
rect 152 8152 192 8184
rect 224 8152 264 8184
rect 296 8152 336 8184
rect 368 8152 408 8184
rect 440 8152 480 8184
rect 512 8152 552 8184
rect 584 8152 624 8184
rect 656 8152 696 8184
rect 728 8152 768 8184
rect 800 8152 840 8184
rect 872 8152 912 8184
rect 944 8152 984 8184
rect 1016 8152 1056 8184
rect 1088 8152 1128 8184
rect 1160 8152 1200 8184
rect 1232 8152 1272 8184
rect 1304 8152 1344 8184
rect 1376 8152 1416 8184
rect 1448 8152 1488 8184
rect 1520 8152 1560 8184
rect 1592 8152 1632 8184
rect 1664 8152 1704 8184
rect 1736 8152 1776 8184
rect 1808 8152 1848 8184
rect 1880 8152 1920 8184
rect 1952 8152 2000 8184
rect 0 8112 2000 8152
rect 0 8080 48 8112
rect 80 8080 120 8112
rect 152 8080 192 8112
rect 224 8080 264 8112
rect 296 8080 336 8112
rect 368 8080 408 8112
rect 440 8080 480 8112
rect 512 8080 552 8112
rect 584 8080 624 8112
rect 656 8080 696 8112
rect 728 8080 768 8112
rect 800 8080 840 8112
rect 872 8080 912 8112
rect 944 8080 984 8112
rect 1016 8080 1056 8112
rect 1088 8080 1128 8112
rect 1160 8080 1200 8112
rect 1232 8080 1272 8112
rect 1304 8080 1344 8112
rect 1376 8080 1416 8112
rect 1448 8080 1488 8112
rect 1520 8080 1560 8112
rect 1592 8080 1632 8112
rect 1664 8080 1704 8112
rect 1736 8080 1776 8112
rect 1808 8080 1848 8112
rect 1880 8080 1920 8112
rect 1952 8080 2000 8112
rect 0 8040 2000 8080
rect 0 8008 48 8040
rect 80 8008 120 8040
rect 152 8008 192 8040
rect 224 8008 264 8040
rect 296 8008 336 8040
rect 368 8008 408 8040
rect 440 8008 480 8040
rect 512 8008 552 8040
rect 584 8008 624 8040
rect 656 8008 696 8040
rect 728 8008 768 8040
rect 800 8008 840 8040
rect 872 8008 912 8040
rect 944 8008 984 8040
rect 1016 8008 1056 8040
rect 1088 8008 1128 8040
rect 1160 8008 1200 8040
rect 1232 8008 1272 8040
rect 1304 8008 1344 8040
rect 1376 8008 1416 8040
rect 1448 8008 1488 8040
rect 1520 8008 1560 8040
rect 1592 8008 1632 8040
rect 1664 8008 1704 8040
rect 1736 8008 1776 8040
rect 1808 8008 1848 8040
rect 1880 8008 1920 8040
rect 1952 8008 2000 8040
rect 0 7968 2000 8008
rect 0 7936 48 7968
rect 80 7936 120 7968
rect 152 7936 192 7968
rect 224 7936 264 7968
rect 296 7936 336 7968
rect 368 7936 408 7968
rect 440 7936 480 7968
rect 512 7936 552 7968
rect 584 7936 624 7968
rect 656 7936 696 7968
rect 728 7936 768 7968
rect 800 7936 840 7968
rect 872 7936 912 7968
rect 944 7936 984 7968
rect 1016 7936 1056 7968
rect 1088 7936 1128 7968
rect 1160 7936 1200 7968
rect 1232 7936 1272 7968
rect 1304 7936 1344 7968
rect 1376 7936 1416 7968
rect 1448 7936 1488 7968
rect 1520 7936 1560 7968
rect 1592 7936 1632 7968
rect 1664 7936 1704 7968
rect 1736 7936 1776 7968
rect 1808 7936 1848 7968
rect 1880 7936 1920 7968
rect 1952 7936 2000 7968
rect 0 7896 2000 7936
rect 0 7864 48 7896
rect 80 7864 120 7896
rect 152 7864 192 7896
rect 224 7864 264 7896
rect 296 7864 336 7896
rect 368 7864 408 7896
rect 440 7864 480 7896
rect 512 7864 552 7896
rect 584 7864 624 7896
rect 656 7864 696 7896
rect 728 7864 768 7896
rect 800 7864 840 7896
rect 872 7864 912 7896
rect 944 7864 984 7896
rect 1016 7864 1056 7896
rect 1088 7864 1128 7896
rect 1160 7864 1200 7896
rect 1232 7864 1272 7896
rect 1304 7864 1344 7896
rect 1376 7864 1416 7896
rect 1448 7864 1488 7896
rect 1520 7864 1560 7896
rect 1592 7864 1632 7896
rect 1664 7864 1704 7896
rect 1736 7864 1776 7896
rect 1808 7864 1848 7896
rect 1880 7864 1920 7896
rect 1952 7864 2000 7896
rect 0 7824 2000 7864
rect 0 7792 48 7824
rect 80 7792 120 7824
rect 152 7792 192 7824
rect 224 7792 264 7824
rect 296 7792 336 7824
rect 368 7792 408 7824
rect 440 7792 480 7824
rect 512 7792 552 7824
rect 584 7792 624 7824
rect 656 7792 696 7824
rect 728 7792 768 7824
rect 800 7792 840 7824
rect 872 7792 912 7824
rect 944 7792 984 7824
rect 1016 7792 1056 7824
rect 1088 7792 1128 7824
rect 1160 7792 1200 7824
rect 1232 7792 1272 7824
rect 1304 7792 1344 7824
rect 1376 7792 1416 7824
rect 1448 7792 1488 7824
rect 1520 7792 1560 7824
rect 1592 7792 1632 7824
rect 1664 7792 1704 7824
rect 1736 7792 1776 7824
rect 1808 7792 1848 7824
rect 1880 7792 1920 7824
rect 1952 7792 2000 7824
rect 0 7752 2000 7792
rect 0 7720 48 7752
rect 80 7720 120 7752
rect 152 7720 192 7752
rect 224 7720 264 7752
rect 296 7720 336 7752
rect 368 7720 408 7752
rect 440 7720 480 7752
rect 512 7720 552 7752
rect 584 7720 624 7752
rect 656 7720 696 7752
rect 728 7720 768 7752
rect 800 7720 840 7752
rect 872 7720 912 7752
rect 944 7720 984 7752
rect 1016 7720 1056 7752
rect 1088 7720 1128 7752
rect 1160 7720 1200 7752
rect 1232 7720 1272 7752
rect 1304 7720 1344 7752
rect 1376 7720 1416 7752
rect 1448 7720 1488 7752
rect 1520 7720 1560 7752
rect 1592 7720 1632 7752
rect 1664 7720 1704 7752
rect 1736 7720 1776 7752
rect 1808 7720 1848 7752
rect 1880 7720 1920 7752
rect 1952 7720 2000 7752
rect 0 7680 2000 7720
rect 0 7648 48 7680
rect 80 7648 120 7680
rect 152 7648 192 7680
rect 224 7648 264 7680
rect 296 7648 336 7680
rect 368 7648 408 7680
rect 440 7648 480 7680
rect 512 7648 552 7680
rect 584 7648 624 7680
rect 656 7648 696 7680
rect 728 7648 768 7680
rect 800 7648 840 7680
rect 872 7648 912 7680
rect 944 7648 984 7680
rect 1016 7648 1056 7680
rect 1088 7648 1128 7680
rect 1160 7648 1200 7680
rect 1232 7648 1272 7680
rect 1304 7648 1344 7680
rect 1376 7648 1416 7680
rect 1448 7648 1488 7680
rect 1520 7648 1560 7680
rect 1592 7648 1632 7680
rect 1664 7648 1704 7680
rect 1736 7648 1776 7680
rect 1808 7648 1848 7680
rect 1880 7648 1920 7680
rect 1952 7648 2000 7680
rect 0 7608 2000 7648
rect 0 7576 48 7608
rect 80 7576 120 7608
rect 152 7576 192 7608
rect 224 7576 264 7608
rect 296 7576 336 7608
rect 368 7576 408 7608
rect 440 7576 480 7608
rect 512 7576 552 7608
rect 584 7576 624 7608
rect 656 7576 696 7608
rect 728 7576 768 7608
rect 800 7576 840 7608
rect 872 7576 912 7608
rect 944 7576 984 7608
rect 1016 7576 1056 7608
rect 1088 7576 1128 7608
rect 1160 7576 1200 7608
rect 1232 7576 1272 7608
rect 1304 7576 1344 7608
rect 1376 7576 1416 7608
rect 1448 7576 1488 7608
rect 1520 7576 1560 7608
rect 1592 7576 1632 7608
rect 1664 7576 1704 7608
rect 1736 7576 1776 7608
rect 1808 7576 1848 7608
rect 1880 7576 1920 7608
rect 1952 7576 2000 7608
rect 0 7536 2000 7576
rect 0 7504 48 7536
rect 80 7504 120 7536
rect 152 7504 192 7536
rect 224 7504 264 7536
rect 296 7504 336 7536
rect 368 7504 408 7536
rect 440 7504 480 7536
rect 512 7504 552 7536
rect 584 7504 624 7536
rect 656 7504 696 7536
rect 728 7504 768 7536
rect 800 7504 840 7536
rect 872 7504 912 7536
rect 944 7504 984 7536
rect 1016 7504 1056 7536
rect 1088 7504 1128 7536
rect 1160 7504 1200 7536
rect 1232 7504 1272 7536
rect 1304 7504 1344 7536
rect 1376 7504 1416 7536
rect 1448 7504 1488 7536
rect 1520 7504 1560 7536
rect 1592 7504 1632 7536
rect 1664 7504 1704 7536
rect 1736 7504 1776 7536
rect 1808 7504 1848 7536
rect 1880 7504 1920 7536
rect 1952 7504 2000 7536
rect 0 7464 2000 7504
rect 0 7432 48 7464
rect 80 7432 120 7464
rect 152 7432 192 7464
rect 224 7432 264 7464
rect 296 7432 336 7464
rect 368 7432 408 7464
rect 440 7432 480 7464
rect 512 7432 552 7464
rect 584 7432 624 7464
rect 656 7432 696 7464
rect 728 7432 768 7464
rect 800 7432 840 7464
rect 872 7432 912 7464
rect 944 7432 984 7464
rect 1016 7432 1056 7464
rect 1088 7432 1128 7464
rect 1160 7432 1200 7464
rect 1232 7432 1272 7464
rect 1304 7432 1344 7464
rect 1376 7432 1416 7464
rect 1448 7432 1488 7464
rect 1520 7432 1560 7464
rect 1592 7432 1632 7464
rect 1664 7432 1704 7464
rect 1736 7432 1776 7464
rect 1808 7432 1848 7464
rect 1880 7432 1920 7464
rect 1952 7432 2000 7464
rect 0 7392 2000 7432
rect 0 7360 48 7392
rect 80 7360 120 7392
rect 152 7360 192 7392
rect 224 7360 264 7392
rect 296 7360 336 7392
rect 368 7360 408 7392
rect 440 7360 480 7392
rect 512 7360 552 7392
rect 584 7360 624 7392
rect 656 7360 696 7392
rect 728 7360 768 7392
rect 800 7360 840 7392
rect 872 7360 912 7392
rect 944 7360 984 7392
rect 1016 7360 1056 7392
rect 1088 7360 1128 7392
rect 1160 7360 1200 7392
rect 1232 7360 1272 7392
rect 1304 7360 1344 7392
rect 1376 7360 1416 7392
rect 1448 7360 1488 7392
rect 1520 7360 1560 7392
rect 1592 7360 1632 7392
rect 1664 7360 1704 7392
rect 1736 7360 1776 7392
rect 1808 7360 1848 7392
rect 1880 7360 1920 7392
rect 1952 7360 2000 7392
rect 0 7320 2000 7360
rect 0 7288 48 7320
rect 80 7288 120 7320
rect 152 7288 192 7320
rect 224 7288 264 7320
rect 296 7288 336 7320
rect 368 7288 408 7320
rect 440 7288 480 7320
rect 512 7288 552 7320
rect 584 7288 624 7320
rect 656 7288 696 7320
rect 728 7288 768 7320
rect 800 7288 840 7320
rect 872 7288 912 7320
rect 944 7288 984 7320
rect 1016 7288 1056 7320
rect 1088 7288 1128 7320
rect 1160 7288 1200 7320
rect 1232 7288 1272 7320
rect 1304 7288 1344 7320
rect 1376 7288 1416 7320
rect 1448 7288 1488 7320
rect 1520 7288 1560 7320
rect 1592 7288 1632 7320
rect 1664 7288 1704 7320
rect 1736 7288 1776 7320
rect 1808 7288 1848 7320
rect 1880 7288 1920 7320
rect 1952 7288 2000 7320
rect 0 7248 2000 7288
rect 0 7216 48 7248
rect 80 7216 120 7248
rect 152 7216 192 7248
rect 224 7216 264 7248
rect 296 7216 336 7248
rect 368 7216 408 7248
rect 440 7216 480 7248
rect 512 7216 552 7248
rect 584 7216 624 7248
rect 656 7216 696 7248
rect 728 7216 768 7248
rect 800 7216 840 7248
rect 872 7216 912 7248
rect 944 7216 984 7248
rect 1016 7216 1056 7248
rect 1088 7216 1128 7248
rect 1160 7216 1200 7248
rect 1232 7216 1272 7248
rect 1304 7216 1344 7248
rect 1376 7216 1416 7248
rect 1448 7216 1488 7248
rect 1520 7216 1560 7248
rect 1592 7216 1632 7248
rect 1664 7216 1704 7248
rect 1736 7216 1776 7248
rect 1808 7216 1848 7248
rect 1880 7216 1920 7248
rect 1952 7216 2000 7248
rect 0 7176 2000 7216
rect 0 7144 48 7176
rect 80 7144 120 7176
rect 152 7144 192 7176
rect 224 7144 264 7176
rect 296 7144 336 7176
rect 368 7144 408 7176
rect 440 7144 480 7176
rect 512 7144 552 7176
rect 584 7144 624 7176
rect 656 7144 696 7176
rect 728 7144 768 7176
rect 800 7144 840 7176
rect 872 7144 912 7176
rect 944 7144 984 7176
rect 1016 7144 1056 7176
rect 1088 7144 1128 7176
rect 1160 7144 1200 7176
rect 1232 7144 1272 7176
rect 1304 7144 1344 7176
rect 1376 7144 1416 7176
rect 1448 7144 1488 7176
rect 1520 7144 1560 7176
rect 1592 7144 1632 7176
rect 1664 7144 1704 7176
rect 1736 7144 1776 7176
rect 1808 7144 1848 7176
rect 1880 7144 1920 7176
rect 1952 7144 2000 7176
rect 0 7104 2000 7144
rect 0 7072 48 7104
rect 80 7072 120 7104
rect 152 7072 192 7104
rect 224 7072 264 7104
rect 296 7072 336 7104
rect 368 7072 408 7104
rect 440 7072 480 7104
rect 512 7072 552 7104
rect 584 7072 624 7104
rect 656 7072 696 7104
rect 728 7072 768 7104
rect 800 7072 840 7104
rect 872 7072 912 7104
rect 944 7072 984 7104
rect 1016 7072 1056 7104
rect 1088 7072 1128 7104
rect 1160 7072 1200 7104
rect 1232 7072 1272 7104
rect 1304 7072 1344 7104
rect 1376 7072 1416 7104
rect 1448 7072 1488 7104
rect 1520 7072 1560 7104
rect 1592 7072 1632 7104
rect 1664 7072 1704 7104
rect 1736 7072 1776 7104
rect 1808 7072 1848 7104
rect 1880 7072 1920 7104
rect 1952 7072 2000 7104
rect 0 7032 2000 7072
rect 0 7000 48 7032
rect 80 7000 120 7032
rect 152 7000 192 7032
rect 224 7000 264 7032
rect 296 7000 336 7032
rect 368 7000 408 7032
rect 440 7000 480 7032
rect 512 7000 552 7032
rect 584 7000 624 7032
rect 656 7000 696 7032
rect 728 7000 768 7032
rect 800 7000 840 7032
rect 872 7000 912 7032
rect 944 7000 984 7032
rect 1016 7000 1056 7032
rect 1088 7000 1128 7032
rect 1160 7000 1200 7032
rect 1232 7000 1272 7032
rect 1304 7000 1344 7032
rect 1376 7000 1416 7032
rect 1448 7000 1488 7032
rect 1520 7000 1560 7032
rect 1592 7000 1632 7032
rect 1664 7000 1704 7032
rect 1736 7000 1776 7032
rect 1808 7000 1848 7032
rect 1880 7000 1920 7032
rect 1952 7000 2000 7032
rect 0 6960 2000 7000
rect 0 6928 48 6960
rect 80 6928 120 6960
rect 152 6928 192 6960
rect 224 6928 264 6960
rect 296 6928 336 6960
rect 368 6928 408 6960
rect 440 6928 480 6960
rect 512 6928 552 6960
rect 584 6928 624 6960
rect 656 6928 696 6960
rect 728 6928 768 6960
rect 800 6928 840 6960
rect 872 6928 912 6960
rect 944 6928 984 6960
rect 1016 6928 1056 6960
rect 1088 6928 1128 6960
rect 1160 6928 1200 6960
rect 1232 6928 1272 6960
rect 1304 6928 1344 6960
rect 1376 6928 1416 6960
rect 1448 6928 1488 6960
rect 1520 6928 1560 6960
rect 1592 6928 1632 6960
rect 1664 6928 1704 6960
rect 1736 6928 1776 6960
rect 1808 6928 1848 6960
rect 1880 6928 1920 6960
rect 1952 6928 2000 6960
rect 0 6888 2000 6928
rect 0 6856 48 6888
rect 80 6856 120 6888
rect 152 6856 192 6888
rect 224 6856 264 6888
rect 296 6856 336 6888
rect 368 6856 408 6888
rect 440 6856 480 6888
rect 512 6856 552 6888
rect 584 6856 624 6888
rect 656 6856 696 6888
rect 728 6856 768 6888
rect 800 6856 840 6888
rect 872 6856 912 6888
rect 944 6856 984 6888
rect 1016 6856 1056 6888
rect 1088 6856 1128 6888
rect 1160 6856 1200 6888
rect 1232 6856 1272 6888
rect 1304 6856 1344 6888
rect 1376 6856 1416 6888
rect 1448 6856 1488 6888
rect 1520 6856 1560 6888
rect 1592 6856 1632 6888
rect 1664 6856 1704 6888
rect 1736 6856 1776 6888
rect 1808 6856 1848 6888
rect 1880 6856 1920 6888
rect 1952 6856 2000 6888
rect 0 6800 2000 6856
rect 0 6544 2000 6600
rect 0 6512 48 6544
rect 80 6512 120 6544
rect 152 6512 192 6544
rect 224 6512 264 6544
rect 296 6512 336 6544
rect 368 6512 408 6544
rect 440 6512 480 6544
rect 512 6512 552 6544
rect 584 6512 624 6544
rect 656 6512 696 6544
rect 728 6512 768 6544
rect 800 6512 840 6544
rect 872 6512 912 6544
rect 944 6512 984 6544
rect 1016 6512 1056 6544
rect 1088 6512 1128 6544
rect 1160 6512 1200 6544
rect 1232 6512 1272 6544
rect 1304 6512 1344 6544
rect 1376 6512 1416 6544
rect 1448 6512 1488 6544
rect 1520 6512 1560 6544
rect 1592 6512 1632 6544
rect 1664 6512 1704 6544
rect 1736 6512 1776 6544
rect 1808 6512 1848 6544
rect 1880 6512 1920 6544
rect 1952 6512 2000 6544
rect 0 6472 2000 6512
rect 0 6440 48 6472
rect 80 6440 120 6472
rect 152 6440 192 6472
rect 224 6440 264 6472
rect 296 6440 336 6472
rect 368 6440 408 6472
rect 440 6440 480 6472
rect 512 6440 552 6472
rect 584 6440 624 6472
rect 656 6440 696 6472
rect 728 6440 768 6472
rect 800 6440 840 6472
rect 872 6440 912 6472
rect 944 6440 984 6472
rect 1016 6440 1056 6472
rect 1088 6440 1128 6472
rect 1160 6440 1200 6472
rect 1232 6440 1272 6472
rect 1304 6440 1344 6472
rect 1376 6440 1416 6472
rect 1448 6440 1488 6472
rect 1520 6440 1560 6472
rect 1592 6440 1632 6472
rect 1664 6440 1704 6472
rect 1736 6440 1776 6472
rect 1808 6440 1848 6472
rect 1880 6440 1920 6472
rect 1952 6440 2000 6472
rect 0 6400 2000 6440
rect 0 6368 48 6400
rect 80 6368 120 6400
rect 152 6368 192 6400
rect 224 6368 264 6400
rect 296 6368 336 6400
rect 368 6368 408 6400
rect 440 6368 480 6400
rect 512 6368 552 6400
rect 584 6368 624 6400
rect 656 6368 696 6400
rect 728 6368 768 6400
rect 800 6368 840 6400
rect 872 6368 912 6400
rect 944 6368 984 6400
rect 1016 6368 1056 6400
rect 1088 6368 1128 6400
rect 1160 6368 1200 6400
rect 1232 6368 1272 6400
rect 1304 6368 1344 6400
rect 1376 6368 1416 6400
rect 1448 6368 1488 6400
rect 1520 6368 1560 6400
rect 1592 6368 1632 6400
rect 1664 6368 1704 6400
rect 1736 6368 1776 6400
rect 1808 6368 1848 6400
rect 1880 6368 1920 6400
rect 1952 6368 2000 6400
rect 0 6328 2000 6368
rect 0 6296 48 6328
rect 80 6296 120 6328
rect 152 6296 192 6328
rect 224 6296 264 6328
rect 296 6296 336 6328
rect 368 6296 408 6328
rect 440 6296 480 6328
rect 512 6296 552 6328
rect 584 6296 624 6328
rect 656 6296 696 6328
rect 728 6296 768 6328
rect 800 6296 840 6328
rect 872 6296 912 6328
rect 944 6296 984 6328
rect 1016 6296 1056 6328
rect 1088 6296 1128 6328
rect 1160 6296 1200 6328
rect 1232 6296 1272 6328
rect 1304 6296 1344 6328
rect 1376 6296 1416 6328
rect 1448 6296 1488 6328
rect 1520 6296 1560 6328
rect 1592 6296 1632 6328
rect 1664 6296 1704 6328
rect 1736 6296 1776 6328
rect 1808 6296 1848 6328
rect 1880 6296 1920 6328
rect 1952 6296 2000 6328
rect 0 6256 2000 6296
rect 0 6224 48 6256
rect 80 6224 120 6256
rect 152 6224 192 6256
rect 224 6224 264 6256
rect 296 6224 336 6256
rect 368 6224 408 6256
rect 440 6224 480 6256
rect 512 6224 552 6256
rect 584 6224 624 6256
rect 656 6224 696 6256
rect 728 6224 768 6256
rect 800 6224 840 6256
rect 872 6224 912 6256
rect 944 6224 984 6256
rect 1016 6224 1056 6256
rect 1088 6224 1128 6256
rect 1160 6224 1200 6256
rect 1232 6224 1272 6256
rect 1304 6224 1344 6256
rect 1376 6224 1416 6256
rect 1448 6224 1488 6256
rect 1520 6224 1560 6256
rect 1592 6224 1632 6256
rect 1664 6224 1704 6256
rect 1736 6224 1776 6256
rect 1808 6224 1848 6256
rect 1880 6224 1920 6256
rect 1952 6224 2000 6256
rect 0 6184 2000 6224
rect 0 6152 48 6184
rect 80 6152 120 6184
rect 152 6152 192 6184
rect 224 6152 264 6184
rect 296 6152 336 6184
rect 368 6152 408 6184
rect 440 6152 480 6184
rect 512 6152 552 6184
rect 584 6152 624 6184
rect 656 6152 696 6184
rect 728 6152 768 6184
rect 800 6152 840 6184
rect 872 6152 912 6184
rect 944 6152 984 6184
rect 1016 6152 1056 6184
rect 1088 6152 1128 6184
rect 1160 6152 1200 6184
rect 1232 6152 1272 6184
rect 1304 6152 1344 6184
rect 1376 6152 1416 6184
rect 1448 6152 1488 6184
rect 1520 6152 1560 6184
rect 1592 6152 1632 6184
rect 1664 6152 1704 6184
rect 1736 6152 1776 6184
rect 1808 6152 1848 6184
rect 1880 6152 1920 6184
rect 1952 6152 2000 6184
rect 0 6112 2000 6152
rect 0 6080 48 6112
rect 80 6080 120 6112
rect 152 6080 192 6112
rect 224 6080 264 6112
rect 296 6080 336 6112
rect 368 6080 408 6112
rect 440 6080 480 6112
rect 512 6080 552 6112
rect 584 6080 624 6112
rect 656 6080 696 6112
rect 728 6080 768 6112
rect 800 6080 840 6112
rect 872 6080 912 6112
rect 944 6080 984 6112
rect 1016 6080 1056 6112
rect 1088 6080 1128 6112
rect 1160 6080 1200 6112
rect 1232 6080 1272 6112
rect 1304 6080 1344 6112
rect 1376 6080 1416 6112
rect 1448 6080 1488 6112
rect 1520 6080 1560 6112
rect 1592 6080 1632 6112
rect 1664 6080 1704 6112
rect 1736 6080 1776 6112
rect 1808 6080 1848 6112
rect 1880 6080 1920 6112
rect 1952 6080 2000 6112
rect 0 6040 2000 6080
rect 0 6008 48 6040
rect 80 6008 120 6040
rect 152 6008 192 6040
rect 224 6008 264 6040
rect 296 6008 336 6040
rect 368 6008 408 6040
rect 440 6008 480 6040
rect 512 6008 552 6040
rect 584 6008 624 6040
rect 656 6008 696 6040
rect 728 6008 768 6040
rect 800 6008 840 6040
rect 872 6008 912 6040
rect 944 6008 984 6040
rect 1016 6008 1056 6040
rect 1088 6008 1128 6040
rect 1160 6008 1200 6040
rect 1232 6008 1272 6040
rect 1304 6008 1344 6040
rect 1376 6008 1416 6040
rect 1448 6008 1488 6040
rect 1520 6008 1560 6040
rect 1592 6008 1632 6040
rect 1664 6008 1704 6040
rect 1736 6008 1776 6040
rect 1808 6008 1848 6040
rect 1880 6008 1920 6040
rect 1952 6008 2000 6040
rect 0 5968 2000 6008
rect 0 5936 48 5968
rect 80 5936 120 5968
rect 152 5936 192 5968
rect 224 5936 264 5968
rect 296 5936 336 5968
rect 368 5936 408 5968
rect 440 5936 480 5968
rect 512 5936 552 5968
rect 584 5936 624 5968
rect 656 5936 696 5968
rect 728 5936 768 5968
rect 800 5936 840 5968
rect 872 5936 912 5968
rect 944 5936 984 5968
rect 1016 5936 1056 5968
rect 1088 5936 1128 5968
rect 1160 5936 1200 5968
rect 1232 5936 1272 5968
rect 1304 5936 1344 5968
rect 1376 5936 1416 5968
rect 1448 5936 1488 5968
rect 1520 5936 1560 5968
rect 1592 5936 1632 5968
rect 1664 5936 1704 5968
rect 1736 5936 1776 5968
rect 1808 5936 1848 5968
rect 1880 5936 1920 5968
rect 1952 5936 2000 5968
rect 0 5896 2000 5936
rect 0 5864 48 5896
rect 80 5864 120 5896
rect 152 5864 192 5896
rect 224 5864 264 5896
rect 296 5864 336 5896
rect 368 5864 408 5896
rect 440 5864 480 5896
rect 512 5864 552 5896
rect 584 5864 624 5896
rect 656 5864 696 5896
rect 728 5864 768 5896
rect 800 5864 840 5896
rect 872 5864 912 5896
rect 944 5864 984 5896
rect 1016 5864 1056 5896
rect 1088 5864 1128 5896
rect 1160 5864 1200 5896
rect 1232 5864 1272 5896
rect 1304 5864 1344 5896
rect 1376 5864 1416 5896
rect 1448 5864 1488 5896
rect 1520 5864 1560 5896
rect 1592 5864 1632 5896
rect 1664 5864 1704 5896
rect 1736 5864 1776 5896
rect 1808 5864 1848 5896
rect 1880 5864 1920 5896
rect 1952 5864 2000 5896
rect 0 5824 2000 5864
rect 0 5792 48 5824
rect 80 5792 120 5824
rect 152 5792 192 5824
rect 224 5792 264 5824
rect 296 5792 336 5824
rect 368 5792 408 5824
rect 440 5792 480 5824
rect 512 5792 552 5824
rect 584 5792 624 5824
rect 656 5792 696 5824
rect 728 5792 768 5824
rect 800 5792 840 5824
rect 872 5792 912 5824
rect 944 5792 984 5824
rect 1016 5792 1056 5824
rect 1088 5792 1128 5824
rect 1160 5792 1200 5824
rect 1232 5792 1272 5824
rect 1304 5792 1344 5824
rect 1376 5792 1416 5824
rect 1448 5792 1488 5824
rect 1520 5792 1560 5824
rect 1592 5792 1632 5824
rect 1664 5792 1704 5824
rect 1736 5792 1776 5824
rect 1808 5792 1848 5824
rect 1880 5792 1920 5824
rect 1952 5792 2000 5824
rect 0 5752 2000 5792
rect 0 5720 48 5752
rect 80 5720 120 5752
rect 152 5720 192 5752
rect 224 5720 264 5752
rect 296 5720 336 5752
rect 368 5720 408 5752
rect 440 5720 480 5752
rect 512 5720 552 5752
rect 584 5720 624 5752
rect 656 5720 696 5752
rect 728 5720 768 5752
rect 800 5720 840 5752
rect 872 5720 912 5752
rect 944 5720 984 5752
rect 1016 5720 1056 5752
rect 1088 5720 1128 5752
rect 1160 5720 1200 5752
rect 1232 5720 1272 5752
rect 1304 5720 1344 5752
rect 1376 5720 1416 5752
rect 1448 5720 1488 5752
rect 1520 5720 1560 5752
rect 1592 5720 1632 5752
rect 1664 5720 1704 5752
rect 1736 5720 1776 5752
rect 1808 5720 1848 5752
rect 1880 5720 1920 5752
rect 1952 5720 2000 5752
rect 0 5680 2000 5720
rect 0 5648 48 5680
rect 80 5648 120 5680
rect 152 5648 192 5680
rect 224 5648 264 5680
rect 296 5648 336 5680
rect 368 5648 408 5680
rect 440 5648 480 5680
rect 512 5648 552 5680
rect 584 5648 624 5680
rect 656 5648 696 5680
rect 728 5648 768 5680
rect 800 5648 840 5680
rect 872 5648 912 5680
rect 944 5648 984 5680
rect 1016 5648 1056 5680
rect 1088 5648 1128 5680
rect 1160 5648 1200 5680
rect 1232 5648 1272 5680
rect 1304 5648 1344 5680
rect 1376 5648 1416 5680
rect 1448 5648 1488 5680
rect 1520 5648 1560 5680
rect 1592 5648 1632 5680
rect 1664 5648 1704 5680
rect 1736 5648 1776 5680
rect 1808 5648 1848 5680
rect 1880 5648 1920 5680
rect 1952 5648 2000 5680
rect 0 5608 2000 5648
rect 0 5576 48 5608
rect 80 5576 120 5608
rect 152 5576 192 5608
rect 224 5576 264 5608
rect 296 5576 336 5608
rect 368 5576 408 5608
rect 440 5576 480 5608
rect 512 5576 552 5608
rect 584 5576 624 5608
rect 656 5576 696 5608
rect 728 5576 768 5608
rect 800 5576 840 5608
rect 872 5576 912 5608
rect 944 5576 984 5608
rect 1016 5576 1056 5608
rect 1088 5576 1128 5608
rect 1160 5576 1200 5608
rect 1232 5576 1272 5608
rect 1304 5576 1344 5608
rect 1376 5576 1416 5608
rect 1448 5576 1488 5608
rect 1520 5576 1560 5608
rect 1592 5576 1632 5608
rect 1664 5576 1704 5608
rect 1736 5576 1776 5608
rect 1808 5576 1848 5608
rect 1880 5576 1920 5608
rect 1952 5576 2000 5608
rect 0 5536 2000 5576
rect 0 5504 48 5536
rect 80 5504 120 5536
rect 152 5504 192 5536
rect 224 5504 264 5536
rect 296 5504 336 5536
rect 368 5504 408 5536
rect 440 5504 480 5536
rect 512 5504 552 5536
rect 584 5504 624 5536
rect 656 5504 696 5536
rect 728 5504 768 5536
rect 800 5504 840 5536
rect 872 5504 912 5536
rect 944 5504 984 5536
rect 1016 5504 1056 5536
rect 1088 5504 1128 5536
rect 1160 5504 1200 5536
rect 1232 5504 1272 5536
rect 1304 5504 1344 5536
rect 1376 5504 1416 5536
rect 1448 5504 1488 5536
rect 1520 5504 1560 5536
rect 1592 5504 1632 5536
rect 1664 5504 1704 5536
rect 1736 5504 1776 5536
rect 1808 5504 1848 5536
rect 1880 5504 1920 5536
rect 1952 5504 2000 5536
rect 0 5464 2000 5504
rect 0 5432 48 5464
rect 80 5432 120 5464
rect 152 5432 192 5464
rect 224 5432 264 5464
rect 296 5432 336 5464
rect 368 5432 408 5464
rect 440 5432 480 5464
rect 512 5432 552 5464
rect 584 5432 624 5464
rect 656 5432 696 5464
rect 728 5432 768 5464
rect 800 5432 840 5464
rect 872 5432 912 5464
rect 944 5432 984 5464
rect 1016 5432 1056 5464
rect 1088 5432 1128 5464
rect 1160 5432 1200 5464
rect 1232 5432 1272 5464
rect 1304 5432 1344 5464
rect 1376 5432 1416 5464
rect 1448 5432 1488 5464
rect 1520 5432 1560 5464
rect 1592 5432 1632 5464
rect 1664 5432 1704 5464
rect 1736 5432 1776 5464
rect 1808 5432 1848 5464
rect 1880 5432 1920 5464
rect 1952 5432 2000 5464
rect 0 5392 2000 5432
rect 0 5360 48 5392
rect 80 5360 120 5392
rect 152 5360 192 5392
rect 224 5360 264 5392
rect 296 5360 336 5392
rect 368 5360 408 5392
rect 440 5360 480 5392
rect 512 5360 552 5392
rect 584 5360 624 5392
rect 656 5360 696 5392
rect 728 5360 768 5392
rect 800 5360 840 5392
rect 872 5360 912 5392
rect 944 5360 984 5392
rect 1016 5360 1056 5392
rect 1088 5360 1128 5392
rect 1160 5360 1200 5392
rect 1232 5360 1272 5392
rect 1304 5360 1344 5392
rect 1376 5360 1416 5392
rect 1448 5360 1488 5392
rect 1520 5360 1560 5392
rect 1592 5360 1632 5392
rect 1664 5360 1704 5392
rect 1736 5360 1776 5392
rect 1808 5360 1848 5392
rect 1880 5360 1920 5392
rect 1952 5360 2000 5392
rect 0 5320 2000 5360
rect 0 5288 48 5320
rect 80 5288 120 5320
rect 152 5288 192 5320
rect 224 5288 264 5320
rect 296 5288 336 5320
rect 368 5288 408 5320
rect 440 5288 480 5320
rect 512 5288 552 5320
rect 584 5288 624 5320
rect 656 5288 696 5320
rect 728 5288 768 5320
rect 800 5288 840 5320
rect 872 5288 912 5320
rect 944 5288 984 5320
rect 1016 5288 1056 5320
rect 1088 5288 1128 5320
rect 1160 5288 1200 5320
rect 1232 5288 1272 5320
rect 1304 5288 1344 5320
rect 1376 5288 1416 5320
rect 1448 5288 1488 5320
rect 1520 5288 1560 5320
rect 1592 5288 1632 5320
rect 1664 5288 1704 5320
rect 1736 5288 1776 5320
rect 1808 5288 1848 5320
rect 1880 5288 1920 5320
rect 1952 5288 2000 5320
rect 0 5248 2000 5288
rect 0 5216 48 5248
rect 80 5216 120 5248
rect 152 5216 192 5248
rect 224 5216 264 5248
rect 296 5216 336 5248
rect 368 5216 408 5248
rect 440 5216 480 5248
rect 512 5216 552 5248
rect 584 5216 624 5248
rect 656 5216 696 5248
rect 728 5216 768 5248
rect 800 5216 840 5248
rect 872 5216 912 5248
rect 944 5216 984 5248
rect 1016 5216 1056 5248
rect 1088 5216 1128 5248
rect 1160 5216 1200 5248
rect 1232 5216 1272 5248
rect 1304 5216 1344 5248
rect 1376 5216 1416 5248
rect 1448 5216 1488 5248
rect 1520 5216 1560 5248
rect 1592 5216 1632 5248
rect 1664 5216 1704 5248
rect 1736 5216 1776 5248
rect 1808 5216 1848 5248
rect 1880 5216 1920 5248
rect 1952 5216 2000 5248
rect 0 5176 2000 5216
rect 0 5144 48 5176
rect 80 5144 120 5176
rect 152 5144 192 5176
rect 224 5144 264 5176
rect 296 5144 336 5176
rect 368 5144 408 5176
rect 440 5144 480 5176
rect 512 5144 552 5176
rect 584 5144 624 5176
rect 656 5144 696 5176
rect 728 5144 768 5176
rect 800 5144 840 5176
rect 872 5144 912 5176
rect 944 5144 984 5176
rect 1016 5144 1056 5176
rect 1088 5144 1128 5176
rect 1160 5144 1200 5176
rect 1232 5144 1272 5176
rect 1304 5144 1344 5176
rect 1376 5144 1416 5176
rect 1448 5144 1488 5176
rect 1520 5144 1560 5176
rect 1592 5144 1632 5176
rect 1664 5144 1704 5176
rect 1736 5144 1776 5176
rect 1808 5144 1848 5176
rect 1880 5144 1920 5176
rect 1952 5144 2000 5176
rect 0 5104 2000 5144
rect 0 5072 48 5104
rect 80 5072 120 5104
rect 152 5072 192 5104
rect 224 5072 264 5104
rect 296 5072 336 5104
rect 368 5072 408 5104
rect 440 5072 480 5104
rect 512 5072 552 5104
rect 584 5072 624 5104
rect 656 5072 696 5104
rect 728 5072 768 5104
rect 800 5072 840 5104
rect 872 5072 912 5104
rect 944 5072 984 5104
rect 1016 5072 1056 5104
rect 1088 5072 1128 5104
rect 1160 5072 1200 5104
rect 1232 5072 1272 5104
rect 1304 5072 1344 5104
rect 1376 5072 1416 5104
rect 1448 5072 1488 5104
rect 1520 5072 1560 5104
rect 1592 5072 1632 5104
rect 1664 5072 1704 5104
rect 1736 5072 1776 5104
rect 1808 5072 1848 5104
rect 1880 5072 1920 5104
rect 1952 5072 2000 5104
rect 0 5032 2000 5072
rect 0 5000 48 5032
rect 80 5000 120 5032
rect 152 5000 192 5032
rect 224 5000 264 5032
rect 296 5000 336 5032
rect 368 5000 408 5032
rect 440 5000 480 5032
rect 512 5000 552 5032
rect 584 5000 624 5032
rect 656 5000 696 5032
rect 728 5000 768 5032
rect 800 5000 840 5032
rect 872 5000 912 5032
rect 944 5000 984 5032
rect 1016 5000 1056 5032
rect 1088 5000 1128 5032
rect 1160 5000 1200 5032
rect 1232 5000 1272 5032
rect 1304 5000 1344 5032
rect 1376 5000 1416 5032
rect 1448 5000 1488 5032
rect 1520 5000 1560 5032
rect 1592 5000 1632 5032
rect 1664 5000 1704 5032
rect 1736 5000 1776 5032
rect 1808 5000 1848 5032
rect 1880 5000 1920 5032
rect 1952 5000 2000 5032
rect 0 4960 2000 5000
rect 0 4928 48 4960
rect 80 4928 120 4960
rect 152 4928 192 4960
rect 224 4928 264 4960
rect 296 4928 336 4960
rect 368 4928 408 4960
rect 440 4928 480 4960
rect 512 4928 552 4960
rect 584 4928 624 4960
rect 656 4928 696 4960
rect 728 4928 768 4960
rect 800 4928 840 4960
rect 872 4928 912 4960
rect 944 4928 984 4960
rect 1016 4928 1056 4960
rect 1088 4928 1128 4960
rect 1160 4928 1200 4960
rect 1232 4928 1272 4960
rect 1304 4928 1344 4960
rect 1376 4928 1416 4960
rect 1448 4928 1488 4960
rect 1520 4928 1560 4960
rect 1592 4928 1632 4960
rect 1664 4928 1704 4960
rect 1736 4928 1776 4960
rect 1808 4928 1848 4960
rect 1880 4928 1920 4960
rect 1952 4928 2000 4960
rect 0 4888 2000 4928
rect 0 4856 48 4888
rect 80 4856 120 4888
rect 152 4856 192 4888
rect 224 4856 264 4888
rect 296 4856 336 4888
rect 368 4856 408 4888
rect 440 4856 480 4888
rect 512 4856 552 4888
rect 584 4856 624 4888
rect 656 4856 696 4888
rect 728 4856 768 4888
rect 800 4856 840 4888
rect 872 4856 912 4888
rect 944 4856 984 4888
rect 1016 4856 1056 4888
rect 1088 4856 1128 4888
rect 1160 4856 1200 4888
rect 1232 4856 1272 4888
rect 1304 4856 1344 4888
rect 1376 4856 1416 4888
rect 1448 4856 1488 4888
rect 1520 4856 1560 4888
rect 1592 4856 1632 4888
rect 1664 4856 1704 4888
rect 1736 4856 1776 4888
rect 1808 4856 1848 4888
rect 1880 4856 1920 4888
rect 1952 4856 2000 4888
rect 0 4816 2000 4856
rect 0 4784 48 4816
rect 80 4784 120 4816
rect 152 4784 192 4816
rect 224 4784 264 4816
rect 296 4784 336 4816
rect 368 4784 408 4816
rect 440 4784 480 4816
rect 512 4784 552 4816
rect 584 4784 624 4816
rect 656 4784 696 4816
rect 728 4784 768 4816
rect 800 4784 840 4816
rect 872 4784 912 4816
rect 944 4784 984 4816
rect 1016 4784 1056 4816
rect 1088 4784 1128 4816
rect 1160 4784 1200 4816
rect 1232 4784 1272 4816
rect 1304 4784 1344 4816
rect 1376 4784 1416 4816
rect 1448 4784 1488 4816
rect 1520 4784 1560 4816
rect 1592 4784 1632 4816
rect 1664 4784 1704 4816
rect 1736 4784 1776 4816
rect 1808 4784 1848 4816
rect 1880 4784 1920 4816
rect 1952 4784 2000 4816
rect 0 4744 2000 4784
rect 0 4712 48 4744
rect 80 4712 120 4744
rect 152 4712 192 4744
rect 224 4712 264 4744
rect 296 4712 336 4744
rect 368 4712 408 4744
rect 440 4712 480 4744
rect 512 4712 552 4744
rect 584 4712 624 4744
rect 656 4712 696 4744
rect 728 4712 768 4744
rect 800 4712 840 4744
rect 872 4712 912 4744
rect 944 4712 984 4744
rect 1016 4712 1056 4744
rect 1088 4712 1128 4744
rect 1160 4712 1200 4744
rect 1232 4712 1272 4744
rect 1304 4712 1344 4744
rect 1376 4712 1416 4744
rect 1448 4712 1488 4744
rect 1520 4712 1560 4744
rect 1592 4712 1632 4744
rect 1664 4712 1704 4744
rect 1736 4712 1776 4744
rect 1808 4712 1848 4744
rect 1880 4712 1920 4744
rect 1952 4712 2000 4744
rect 0 4672 2000 4712
rect 0 4640 48 4672
rect 80 4640 120 4672
rect 152 4640 192 4672
rect 224 4640 264 4672
rect 296 4640 336 4672
rect 368 4640 408 4672
rect 440 4640 480 4672
rect 512 4640 552 4672
rect 584 4640 624 4672
rect 656 4640 696 4672
rect 728 4640 768 4672
rect 800 4640 840 4672
rect 872 4640 912 4672
rect 944 4640 984 4672
rect 1016 4640 1056 4672
rect 1088 4640 1128 4672
rect 1160 4640 1200 4672
rect 1232 4640 1272 4672
rect 1304 4640 1344 4672
rect 1376 4640 1416 4672
rect 1448 4640 1488 4672
rect 1520 4640 1560 4672
rect 1592 4640 1632 4672
rect 1664 4640 1704 4672
rect 1736 4640 1776 4672
rect 1808 4640 1848 4672
rect 1880 4640 1920 4672
rect 1952 4640 2000 4672
rect 0 4600 2000 4640
rect 0 4568 48 4600
rect 80 4568 120 4600
rect 152 4568 192 4600
rect 224 4568 264 4600
rect 296 4568 336 4600
rect 368 4568 408 4600
rect 440 4568 480 4600
rect 512 4568 552 4600
rect 584 4568 624 4600
rect 656 4568 696 4600
rect 728 4568 768 4600
rect 800 4568 840 4600
rect 872 4568 912 4600
rect 944 4568 984 4600
rect 1016 4568 1056 4600
rect 1088 4568 1128 4600
rect 1160 4568 1200 4600
rect 1232 4568 1272 4600
rect 1304 4568 1344 4600
rect 1376 4568 1416 4600
rect 1448 4568 1488 4600
rect 1520 4568 1560 4600
rect 1592 4568 1632 4600
rect 1664 4568 1704 4600
rect 1736 4568 1776 4600
rect 1808 4568 1848 4600
rect 1880 4568 1920 4600
rect 1952 4568 2000 4600
rect 0 4528 2000 4568
rect 0 4496 48 4528
rect 80 4496 120 4528
rect 152 4496 192 4528
rect 224 4496 264 4528
rect 296 4496 336 4528
rect 368 4496 408 4528
rect 440 4496 480 4528
rect 512 4496 552 4528
rect 584 4496 624 4528
rect 656 4496 696 4528
rect 728 4496 768 4528
rect 800 4496 840 4528
rect 872 4496 912 4528
rect 944 4496 984 4528
rect 1016 4496 1056 4528
rect 1088 4496 1128 4528
rect 1160 4496 1200 4528
rect 1232 4496 1272 4528
rect 1304 4496 1344 4528
rect 1376 4496 1416 4528
rect 1448 4496 1488 4528
rect 1520 4496 1560 4528
rect 1592 4496 1632 4528
rect 1664 4496 1704 4528
rect 1736 4496 1776 4528
rect 1808 4496 1848 4528
rect 1880 4496 1920 4528
rect 1952 4496 2000 4528
rect 0 4456 2000 4496
rect 0 4424 48 4456
rect 80 4424 120 4456
rect 152 4424 192 4456
rect 224 4424 264 4456
rect 296 4424 336 4456
rect 368 4424 408 4456
rect 440 4424 480 4456
rect 512 4424 552 4456
rect 584 4424 624 4456
rect 656 4424 696 4456
rect 728 4424 768 4456
rect 800 4424 840 4456
rect 872 4424 912 4456
rect 944 4424 984 4456
rect 1016 4424 1056 4456
rect 1088 4424 1128 4456
rect 1160 4424 1200 4456
rect 1232 4424 1272 4456
rect 1304 4424 1344 4456
rect 1376 4424 1416 4456
rect 1448 4424 1488 4456
rect 1520 4424 1560 4456
rect 1592 4424 1632 4456
rect 1664 4424 1704 4456
rect 1736 4424 1776 4456
rect 1808 4424 1848 4456
rect 1880 4424 1920 4456
rect 1952 4424 2000 4456
rect 0 4384 2000 4424
rect 0 4352 48 4384
rect 80 4352 120 4384
rect 152 4352 192 4384
rect 224 4352 264 4384
rect 296 4352 336 4384
rect 368 4352 408 4384
rect 440 4352 480 4384
rect 512 4352 552 4384
rect 584 4352 624 4384
rect 656 4352 696 4384
rect 728 4352 768 4384
rect 800 4352 840 4384
rect 872 4352 912 4384
rect 944 4352 984 4384
rect 1016 4352 1056 4384
rect 1088 4352 1128 4384
rect 1160 4352 1200 4384
rect 1232 4352 1272 4384
rect 1304 4352 1344 4384
rect 1376 4352 1416 4384
rect 1448 4352 1488 4384
rect 1520 4352 1560 4384
rect 1592 4352 1632 4384
rect 1664 4352 1704 4384
rect 1736 4352 1776 4384
rect 1808 4352 1848 4384
rect 1880 4352 1920 4384
rect 1952 4352 2000 4384
rect 0 4312 2000 4352
rect 0 4280 48 4312
rect 80 4280 120 4312
rect 152 4280 192 4312
rect 224 4280 264 4312
rect 296 4280 336 4312
rect 368 4280 408 4312
rect 440 4280 480 4312
rect 512 4280 552 4312
rect 584 4280 624 4312
rect 656 4280 696 4312
rect 728 4280 768 4312
rect 800 4280 840 4312
rect 872 4280 912 4312
rect 944 4280 984 4312
rect 1016 4280 1056 4312
rect 1088 4280 1128 4312
rect 1160 4280 1200 4312
rect 1232 4280 1272 4312
rect 1304 4280 1344 4312
rect 1376 4280 1416 4312
rect 1448 4280 1488 4312
rect 1520 4280 1560 4312
rect 1592 4280 1632 4312
rect 1664 4280 1704 4312
rect 1736 4280 1776 4312
rect 1808 4280 1848 4312
rect 1880 4280 1920 4312
rect 1952 4280 2000 4312
rect 0 4240 2000 4280
rect 0 4208 48 4240
rect 80 4208 120 4240
rect 152 4208 192 4240
rect 224 4208 264 4240
rect 296 4208 336 4240
rect 368 4208 408 4240
rect 440 4208 480 4240
rect 512 4208 552 4240
rect 584 4208 624 4240
rect 656 4208 696 4240
rect 728 4208 768 4240
rect 800 4208 840 4240
rect 872 4208 912 4240
rect 944 4208 984 4240
rect 1016 4208 1056 4240
rect 1088 4208 1128 4240
rect 1160 4208 1200 4240
rect 1232 4208 1272 4240
rect 1304 4208 1344 4240
rect 1376 4208 1416 4240
rect 1448 4208 1488 4240
rect 1520 4208 1560 4240
rect 1592 4208 1632 4240
rect 1664 4208 1704 4240
rect 1736 4208 1776 4240
rect 1808 4208 1848 4240
rect 1880 4208 1920 4240
rect 1952 4208 2000 4240
rect 0 4168 2000 4208
rect 0 4136 48 4168
rect 80 4136 120 4168
rect 152 4136 192 4168
rect 224 4136 264 4168
rect 296 4136 336 4168
rect 368 4136 408 4168
rect 440 4136 480 4168
rect 512 4136 552 4168
rect 584 4136 624 4168
rect 656 4136 696 4168
rect 728 4136 768 4168
rect 800 4136 840 4168
rect 872 4136 912 4168
rect 944 4136 984 4168
rect 1016 4136 1056 4168
rect 1088 4136 1128 4168
rect 1160 4136 1200 4168
rect 1232 4136 1272 4168
rect 1304 4136 1344 4168
rect 1376 4136 1416 4168
rect 1448 4136 1488 4168
rect 1520 4136 1560 4168
rect 1592 4136 1632 4168
rect 1664 4136 1704 4168
rect 1736 4136 1776 4168
rect 1808 4136 1848 4168
rect 1880 4136 1920 4168
rect 1952 4136 2000 4168
rect 0 4096 2000 4136
rect 0 4064 48 4096
rect 80 4064 120 4096
rect 152 4064 192 4096
rect 224 4064 264 4096
rect 296 4064 336 4096
rect 368 4064 408 4096
rect 440 4064 480 4096
rect 512 4064 552 4096
rect 584 4064 624 4096
rect 656 4064 696 4096
rect 728 4064 768 4096
rect 800 4064 840 4096
rect 872 4064 912 4096
rect 944 4064 984 4096
rect 1016 4064 1056 4096
rect 1088 4064 1128 4096
rect 1160 4064 1200 4096
rect 1232 4064 1272 4096
rect 1304 4064 1344 4096
rect 1376 4064 1416 4096
rect 1448 4064 1488 4096
rect 1520 4064 1560 4096
rect 1592 4064 1632 4096
rect 1664 4064 1704 4096
rect 1736 4064 1776 4096
rect 1808 4064 1848 4096
rect 1880 4064 1920 4096
rect 1952 4064 2000 4096
rect 0 4024 2000 4064
rect 0 3992 48 4024
rect 80 3992 120 4024
rect 152 3992 192 4024
rect 224 3992 264 4024
rect 296 3992 336 4024
rect 368 3992 408 4024
rect 440 3992 480 4024
rect 512 3992 552 4024
rect 584 3992 624 4024
rect 656 3992 696 4024
rect 728 3992 768 4024
rect 800 3992 840 4024
rect 872 3992 912 4024
rect 944 3992 984 4024
rect 1016 3992 1056 4024
rect 1088 3992 1128 4024
rect 1160 3992 1200 4024
rect 1232 3992 1272 4024
rect 1304 3992 1344 4024
rect 1376 3992 1416 4024
rect 1448 3992 1488 4024
rect 1520 3992 1560 4024
rect 1592 3992 1632 4024
rect 1664 3992 1704 4024
rect 1736 3992 1776 4024
rect 1808 3992 1848 4024
rect 1880 3992 1920 4024
rect 1952 3992 2000 4024
rect 0 3952 2000 3992
rect 0 3920 48 3952
rect 80 3920 120 3952
rect 152 3920 192 3952
rect 224 3920 264 3952
rect 296 3920 336 3952
rect 368 3920 408 3952
rect 440 3920 480 3952
rect 512 3920 552 3952
rect 584 3920 624 3952
rect 656 3920 696 3952
rect 728 3920 768 3952
rect 800 3920 840 3952
rect 872 3920 912 3952
rect 944 3920 984 3952
rect 1016 3920 1056 3952
rect 1088 3920 1128 3952
rect 1160 3920 1200 3952
rect 1232 3920 1272 3952
rect 1304 3920 1344 3952
rect 1376 3920 1416 3952
rect 1448 3920 1488 3952
rect 1520 3920 1560 3952
rect 1592 3920 1632 3952
rect 1664 3920 1704 3952
rect 1736 3920 1776 3952
rect 1808 3920 1848 3952
rect 1880 3920 1920 3952
rect 1952 3920 2000 3952
rect 0 3880 2000 3920
rect 0 3848 48 3880
rect 80 3848 120 3880
rect 152 3848 192 3880
rect 224 3848 264 3880
rect 296 3848 336 3880
rect 368 3848 408 3880
rect 440 3848 480 3880
rect 512 3848 552 3880
rect 584 3848 624 3880
rect 656 3848 696 3880
rect 728 3848 768 3880
rect 800 3848 840 3880
rect 872 3848 912 3880
rect 944 3848 984 3880
rect 1016 3848 1056 3880
rect 1088 3848 1128 3880
rect 1160 3848 1200 3880
rect 1232 3848 1272 3880
rect 1304 3848 1344 3880
rect 1376 3848 1416 3880
rect 1448 3848 1488 3880
rect 1520 3848 1560 3880
rect 1592 3848 1632 3880
rect 1664 3848 1704 3880
rect 1736 3848 1776 3880
rect 1808 3848 1848 3880
rect 1880 3848 1920 3880
rect 1952 3848 2000 3880
rect 0 3808 2000 3848
rect 0 3776 48 3808
rect 80 3776 120 3808
rect 152 3776 192 3808
rect 224 3776 264 3808
rect 296 3776 336 3808
rect 368 3776 408 3808
rect 440 3776 480 3808
rect 512 3776 552 3808
rect 584 3776 624 3808
rect 656 3776 696 3808
rect 728 3776 768 3808
rect 800 3776 840 3808
rect 872 3776 912 3808
rect 944 3776 984 3808
rect 1016 3776 1056 3808
rect 1088 3776 1128 3808
rect 1160 3776 1200 3808
rect 1232 3776 1272 3808
rect 1304 3776 1344 3808
rect 1376 3776 1416 3808
rect 1448 3776 1488 3808
rect 1520 3776 1560 3808
rect 1592 3776 1632 3808
rect 1664 3776 1704 3808
rect 1736 3776 1776 3808
rect 1808 3776 1848 3808
rect 1880 3776 1920 3808
rect 1952 3776 2000 3808
rect 0 3736 2000 3776
rect 0 3704 48 3736
rect 80 3704 120 3736
rect 152 3704 192 3736
rect 224 3704 264 3736
rect 296 3704 336 3736
rect 368 3704 408 3736
rect 440 3704 480 3736
rect 512 3704 552 3736
rect 584 3704 624 3736
rect 656 3704 696 3736
rect 728 3704 768 3736
rect 800 3704 840 3736
rect 872 3704 912 3736
rect 944 3704 984 3736
rect 1016 3704 1056 3736
rect 1088 3704 1128 3736
rect 1160 3704 1200 3736
rect 1232 3704 1272 3736
rect 1304 3704 1344 3736
rect 1376 3704 1416 3736
rect 1448 3704 1488 3736
rect 1520 3704 1560 3736
rect 1592 3704 1632 3736
rect 1664 3704 1704 3736
rect 1736 3704 1776 3736
rect 1808 3704 1848 3736
rect 1880 3704 1920 3736
rect 1952 3704 2000 3736
rect 0 3664 2000 3704
rect 0 3632 48 3664
rect 80 3632 120 3664
rect 152 3632 192 3664
rect 224 3632 264 3664
rect 296 3632 336 3664
rect 368 3632 408 3664
rect 440 3632 480 3664
rect 512 3632 552 3664
rect 584 3632 624 3664
rect 656 3632 696 3664
rect 728 3632 768 3664
rect 800 3632 840 3664
rect 872 3632 912 3664
rect 944 3632 984 3664
rect 1016 3632 1056 3664
rect 1088 3632 1128 3664
rect 1160 3632 1200 3664
rect 1232 3632 1272 3664
rect 1304 3632 1344 3664
rect 1376 3632 1416 3664
rect 1448 3632 1488 3664
rect 1520 3632 1560 3664
rect 1592 3632 1632 3664
rect 1664 3632 1704 3664
rect 1736 3632 1776 3664
rect 1808 3632 1848 3664
rect 1880 3632 1920 3664
rect 1952 3632 2000 3664
rect 0 3592 2000 3632
rect 0 3560 48 3592
rect 80 3560 120 3592
rect 152 3560 192 3592
rect 224 3560 264 3592
rect 296 3560 336 3592
rect 368 3560 408 3592
rect 440 3560 480 3592
rect 512 3560 552 3592
rect 584 3560 624 3592
rect 656 3560 696 3592
rect 728 3560 768 3592
rect 800 3560 840 3592
rect 872 3560 912 3592
rect 944 3560 984 3592
rect 1016 3560 1056 3592
rect 1088 3560 1128 3592
rect 1160 3560 1200 3592
rect 1232 3560 1272 3592
rect 1304 3560 1344 3592
rect 1376 3560 1416 3592
rect 1448 3560 1488 3592
rect 1520 3560 1560 3592
rect 1592 3560 1632 3592
rect 1664 3560 1704 3592
rect 1736 3560 1776 3592
rect 1808 3560 1848 3592
rect 1880 3560 1920 3592
rect 1952 3560 2000 3592
rect 0 3520 2000 3560
rect 0 3488 48 3520
rect 80 3488 120 3520
rect 152 3488 192 3520
rect 224 3488 264 3520
rect 296 3488 336 3520
rect 368 3488 408 3520
rect 440 3488 480 3520
rect 512 3488 552 3520
rect 584 3488 624 3520
rect 656 3488 696 3520
rect 728 3488 768 3520
rect 800 3488 840 3520
rect 872 3488 912 3520
rect 944 3488 984 3520
rect 1016 3488 1056 3520
rect 1088 3488 1128 3520
rect 1160 3488 1200 3520
rect 1232 3488 1272 3520
rect 1304 3488 1344 3520
rect 1376 3488 1416 3520
rect 1448 3488 1488 3520
rect 1520 3488 1560 3520
rect 1592 3488 1632 3520
rect 1664 3488 1704 3520
rect 1736 3488 1776 3520
rect 1808 3488 1848 3520
rect 1880 3488 1920 3520
rect 1952 3488 2000 3520
rect 0 3448 2000 3488
rect 0 3416 48 3448
rect 80 3416 120 3448
rect 152 3416 192 3448
rect 224 3416 264 3448
rect 296 3416 336 3448
rect 368 3416 408 3448
rect 440 3416 480 3448
rect 512 3416 552 3448
rect 584 3416 624 3448
rect 656 3416 696 3448
rect 728 3416 768 3448
rect 800 3416 840 3448
rect 872 3416 912 3448
rect 944 3416 984 3448
rect 1016 3416 1056 3448
rect 1088 3416 1128 3448
rect 1160 3416 1200 3448
rect 1232 3416 1272 3448
rect 1304 3416 1344 3448
rect 1376 3416 1416 3448
rect 1448 3416 1488 3448
rect 1520 3416 1560 3448
rect 1592 3416 1632 3448
rect 1664 3416 1704 3448
rect 1736 3416 1776 3448
rect 1808 3416 1848 3448
rect 1880 3416 1920 3448
rect 1952 3416 2000 3448
rect 0 3376 2000 3416
rect 0 3344 48 3376
rect 80 3344 120 3376
rect 152 3344 192 3376
rect 224 3344 264 3376
rect 296 3344 336 3376
rect 368 3344 408 3376
rect 440 3344 480 3376
rect 512 3344 552 3376
rect 584 3344 624 3376
rect 656 3344 696 3376
rect 728 3344 768 3376
rect 800 3344 840 3376
rect 872 3344 912 3376
rect 944 3344 984 3376
rect 1016 3344 1056 3376
rect 1088 3344 1128 3376
rect 1160 3344 1200 3376
rect 1232 3344 1272 3376
rect 1304 3344 1344 3376
rect 1376 3344 1416 3376
rect 1448 3344 1488 3376
rect 1520 3344 1560 3376
rect 1592 3344 1632 3376
rect 1664 3344 1704 3376
rect 1736 3344 1776 3376
rect 1808 3344 1848 3376
rect 1880 3344 1920 3376
rect 1952 3344 2000 3376
rect 0 3304 2000 3344
rect 0 3272 48 3304
rect 80 3272 120 3304
rect 152 3272 192 3304
rect 224 3272 264 3304
rect 296 3272 336 3304
rect 368 3272 408 3304
rect 440 3272 480 3304
rect 512 3272 552 3304
rect 584 3272 624 3304
rect 656 3272 696 3304
rect 728 3272 768 3304
rect 800 3272 840 3304
rect 872 3272 912 3304
rect 944 3272 984 3304
rect 1016 3272 1056 3304
rect 1088 3272 1128 3304
rect 1160 3272 1200 3304
rect 1232 3272 1272 3304
rect 1304 3272 1344 3304
rect 1376 3272 1416 3304
rect 1448 3272 1488 3304
rect 1520 3272 1560 3304
rect 1592 3272 1632 3304
rect 1664 3272 1704 3304
rect 1736 3272 1776 3304
rect 1808 3272 1848 3304
rect 1880 3272 1920 3304
rect 1952 3272 2000 3304
rect 0 3232 2000 3272
rect 0 3200 48 3232
rect 80 3200 120 3232
rect 152 3200 192 3232
rect 224 3200 264 3232
rect 296 3200 336 3232
rect 368 3200 408 3232
rect 440 3200 480 3232
rect 512 3200 552 3232
rect 584 3200 624 3232
rect 656 3200 696 3232
rect 728 3200 768 3232
rect 800 3200 840 3232
rect 872 3200 912 3232
rect 944 3200 984 3232
rect 1016 3200 1056 3232
rect 1088 3200 1128 3232
rect 1160 3200 1200 3232
rect 1232 3200 1272 3232
rect 1304 3200 1344 3232
rect 1376 3200 1416 3232
rect 1448 3200 1488 3232
rect 1520 3200 1560 3232
rect 1592 3200 1632 3232
rect 1664 3200 1704 3232
rect 1736 3200 1776 3232
rect 1808 3200 1848 3232
rect 1880 3200 1920 3232
rect 1952 3200 2000 3232
rect 0 3160 2000 3200
rect 0 3128 48 3160
rect 80 3128 120 3160
rect 152 3128 192 3160
rect 224 3128 264 3160
rect 296 3128 336 3160
rect 368 3128 408 3160
rect 440 3128 480 3160
rect 512 3128 552 3160
rect 584 3128 624 3160
rect 656 3128 696 3160
rect 728 3128 768 3160
rect 800 3128 840 3160
rect 872 3128 912 3160
rect 944 3128 984 3160
rect 1016 3128 1056 3160
rect 1088 3128 1128 3160
rect 1160 3128 1200 3160
rect 1232 3128 1272 3160
rect 1304 3128 1344 3160
rect 1376 3128 1416 3160
rect 1448 3128 1488 3160
rect 1520 3128 1560 3160
rect 1592 3128 1632 3160
rect 1664 3128 1704 3160
rect 1736 3128 1776 3160
rect 1808 3128 1848 3160
rect 1880 3128 1920 3160
rect 1952 3128 2000 3160
rect 0 3088 2000 3128
rect 0 3056 48 3088
rect 80 3056 120 3088
rect 152 3056 192 3088
rect 224 3056 264 3088
rect 296 3056 336 3088
rect 368 3056 408 3088
rect 440 3056 480 3088
rect 512 3056 552 3088
rect 584 3056 624 3088
rect 656 3056 696 3088
rect 728 3056 768 3088
rect 800 3056 840 3088
rect 872 3056 912 3088
rect 944 3056 984 3088
rect 1016 3056 1056 3088
rect 1088 3056 1128 3088
rect 1160 3056 1200 3088
rect 1232 3056 1272 3088
rect 1304 3056 1344 3088
rect 1376 3056 1416 3088
rect 1448 3056 1488 3088
rect 1520 3056 1560 3088
rect 1592 3056 1632 3088
rect 1664 3056 1704 3088
rect 1736 3056 1776 3088
rect 1808 3056 1848 3088
rect 1880 3056 1920 3088
rect 1952 3056 2000 3088
rect 0 3016 2000 3056
rect 0 2984 48 3016
rect 80 2984 120 3016
rect 152 2984 192 3016
rect 224 2984 264 3016
rect 296 2984 336 3016
rect 368 2984 408 3016
rect 440 2984 480 3016
rect 512 2984 552 3016
rect 584 2984 624 3016
rect 656 2984 696 3016
rect 728 2984 768 3016
rect 800 2984 840 3016
rect 872 2984 912 3016
rect 944 2984 984 3016
rect 1016 2984 1056 3016
rect 1088 2984 1128 3016
rect 1160 2984 1200 3016
rect 1232 2984 1272 3016
rect 1304 2984 1344 3016
rect 1376 2984 1416 3016
rect 1448 2984 1488 3016
rect 1520 2984 1560 3016
rect 1592 2984 1632 3016
rect 1664 2984 1704 3016
rect 1736 2984 1776 3016
rect 1808 2984 1848 3016
rect 1880 2984 1920 3016
rect 1952 2984 2000 3016
rect 0 2944 2000 2984
rect 0 2912 48 2944
rect 80 2912 120 2944
rect 152 2912 192 2944
rect 224 2912 264 2944
rect 296 2912 336 2944
rect 368 2912 408 2944
rect 440 2912 480 2944
rect 512 2912 552 2944
rect 584 2912 624 2944
rect 656 2912 696 2944
rect 728 2912 768 2944
rect 800 2912 840 2944
rect 872 2912 912 2944
rect 944 2912 984 2944
rect 1016 2912 1056 2944
rect 1088 2912 1128 2944
rect 1160 2912 1200 2944
rect 1232 2912 1272 2944
rect 1304 2912 1344 2944
rect 1376 2912 1416 2944
rect 1448 2912 1488 2944
rect 1520 2912 1560 2944
rect 1592 2912 1632 2944
rect 1664 2912 1704 2944
rect 1736 2912 1776 2944
rect 1808 2912 1848 2944
rect 1880 2912 1920 2944
rect 1952 2912 2000 2944
rect 0 2872 2000 2912
rect 0 2840 48 2872
rect 80 2840 120 2872
rect 152 2840 192 2872
rect 224 2840 264 2872
rect 296 2840 336 2872
rect 368 2840 408 2872
rect 440 2840 480 2872
rect 512 2840 552 2872
rect 584 2840 624 2872
rect 656 2840 696 2872
rect 728 2840 768 2872
rect 800 2840 840 2872
rect 872 2840 912 2872
rect 944 2840 984 2872
rect 1016 2840 1056 2872
rect 1088 2840 1128 2872
rect 1160 2840 1200 2872
rect 1232 2840 1272 2872
rect 1304 2840 1344 2872
rect 1376 2840 1416 2872
rect 1448 2840 1488 2872
rect 1520 2840 1560 2872
rect 1592 2840 1632 2872
rect 1664 2840 1704 2872
rect 1736 2840 1776 2872
rect 1808 2840 1848 2872
rect 1880 2840 1920 2872
rect 1952 2840 2000 2872
rect 0 2800 2000 2840
rect 0 2768 48 2800
rect 80 2768 120 2800
rect 152 2768 192 2800
rect 224 2768 264 2800
rect 296 2768 336 2800
rect 368 2768 408 2800
rect 440 2768 480 2800
rect 512 2768 552 2800
rect 584 2768 624 2800
rect 656 2768 696 2800
rect 728 2768 768 2800
rect 800 2768 840 2800
rect 872 2768 912 2800
rect 944 2768 984 2800
rect 1016 2768 1056 2800
rect 1088 2768 1128 2800
rect 1160 2768 1200 2800
rect 1232 2768 1272 2800
rect 1304 2768 1344 2800
rect 1376 2768 1416 2800
rect 1448 2768 1488 2800
rect 1520 2768 1560 2800
rect 1592 2768 1632 2800
rect 1664 2768 1704 2800
rect 1736 2768 1776 2800
rect 1808 2768 1848 2800
rect 1880 2768 1920 2800
rect 1952 2768 2000 2800
rect 0 2728 2000 2768
rect 0 2696 48 2728
rect 80 2696 120 2728
rect 152 2696 192 2728
rect 224 2696 264 2728
rect 296 2696 336 2728
rect 368 2696 408 2728
rect 440 2696 480 2728
rect 512 2696 552 2728
rect 584 2696 624 2728
rect 656 2696 696 2728
rect 728 2696 768 2728
rect 800 2696 840 2728
rect 872 2696 912 2728
rect 944 2696 984 2728
rect 1016 2696 1056 2728
rect 1088 2696 1128 2728
rect 1160 2696 1200 2728
rect 1232 2696 1272 2728
rect 1304 2696 1344 2728
rect 1376 2696 1416 2728
rect 1448 2696 1488 2728
rect 1520 2696 1560 2728
rect 1592 2696 1632 2728
rect 1664 2696 1704 2728
rect 1736 2696 1776 2728
rect 1808 2696 1848 2728
rect 1880 2696 1920 2728
rect 1952 2696 2000 2728
rect 0 2656 2000 2696
rect 0 2624 48 2656
rect 80 2624 120 2656
rect 152 2624 192 2656
rect 224 2624 264 2656
rect 296 2624 336 2656
rect 368 2624 408 2656
rect 440 2624 480 2656
rect 512 2624 552 2656
rect 584 2624 624 2656
rect 656 2624 696 2656
rect 728 2624 768 2656
rect 800 2624 840 2656
rect 872 2624 912 2656
rect 944 2624 984 2656
rect 1016 2624 1056 2656
rect 1088 2624 1128 2656
rect 1160 2624 1200 2656
rect 1232 2624 1272 2656
rect 1304 2624 1344 2656
rect 1376 2624 1416 2656
rect 1448 2624 1488 2656
rect 1520 2624 1560 2656
rect 1592 2624 1632 2656
rect 1664 2624 1704 2656
rect 1736 2624 1776 2656
rect 1808 2624 1848 2656
rect 1880 2624 1920 2656
rect 1952 2624 2000 2656
rect 0 2584 2000 2624
rect 0 2552 48 2584
rect 80 2552 120 2584
rect 152 2552 192 2584
rect 224 2552 264 2584
rect 296 2552 336 2584
rect 368 2552 408 2584
rect 440 2552 480 2584
rect 512 2552 552 2584
rect 584 2552 624 2584
rect 656 2552 696 2584
rect 728 2552 768 2584
rect 800 2552 840 2584
rect 872 2552 912 2584
rect 944 2552 984 2584
rect 1016 2552 1056 2584
rect 1088 2552 1128 2584
rect 1160 2552 1200 2584
rect 1232 2552 1272 2584
rect 1304 2552 1344 2584
rect 1376 2552 1416 2584
rect 1448 2552 1488 2584
rect 1520 2552 1560 2584
rect 1592 2552 1632 2584
rect 1664 2552 1704 2584
rect 1736 2552 1776 2584
rect 1808 2552 1848 2584
rect 1880 2552 1920 2584
rect 1952 2552 2000 2584
rect 0 2512 2000 2552
rect 0 2480 48 2512
rect 80 2480 120 2512
rect 152 2480 192 2512
rect 224 2480 264 2512
rect 296 2480 336 2512
rect 368 2480 408 2512
rect 440 2480 480 2512
rect 512 2480 552 2512
rect 584 2480 624 2512
rect 656 2480 696 2512
rect 728 2480 768 2512
rect 800 2480 840 2512
rect 872 2480 912 2512
rect 944 2480 984 2512
rect 1016 2480 1056 2512
rect 1088 2480 1128 2512
rect 1160 2480 1200 2512
rect 1232 2480 1272 2512
rect 1304 2480 1344 2512
rect 1376 2480 1416 2512
rect 1448 2480 1488 2512
rect 1520 2480 1560 2512
rect 1592 2480 1632 2512
rect 1664 2480 1704 2512
rect 1736 2480 1776 2512
rect 1808 2480 1848 2512
rect 1880 2480 1920 2512
rect 1952 2480 2000 2512
rect 0 2440 2000 2480
rect 0 2408 48 2440
rect 80 2408 120 2440
rect 152 2408 192 2440
rect 224 2408 264 2440
rect 296 2408 336 2440
rect 368 2408 408 2440
rect 440 2408 480 2440
rect 512 2408 552 2440
rect 584 2408 624 2440
rect 656 2408 696 2440
rect 728 2408 768 2440
rect 800 2408 840 2440
rect 872 2408 912 2440
rect 944 2408 984 2440
rect 1016 2408 1056 2440
rect 1088 2408 1128 2440
rect 1160 2408 1200 2440
rect 1232 2408 1272 2440
rect 1304 2408 1344 2440
rect 1376 2408 1416 2440
rect 1448 2408 1488 2440
rect 1520 2408 1560 2440
rect 1592 2408 1632 2440
rect 1664 2408 1704 2440
rect 1736 2408 1776 2440
rect 1808 2408 1848 2440
rect 1880 2408 1920 2440
rect 1952 2408 2000 2440
rect 0 2368 2000 2408
rect 0 2336 48 2368
rect 80 2336 120 2368
rect 152 2336 192 2368
rect 224 2336 264 2368
rect 296 2336 336 2368
rect 368 2336 408 2368
rect 440 2336 480 2368
rect 512 2336 552 2368
rect 584 2336 624 2368
rect 656 2336 696 2368
rect 728 2336 768 2368
rect 800 2336 840 2368
rect 872 2336 912 2368
rect 944 2336 984 2368
rect 1016 2336 1056 2368
rect 1088 2336 1128 2368
rect 1160 2336 1200 2368
rect 1232 2336 1272 2368
rect 1304 2336 1344 2368
rect 1376 2336 1416 2368
rect 1448 2336 1488 2368
rect 1520 2336 1560 2368
rect 1592 2336 1632 2368
rect 1664 2336 1704 2368
rect 1736 2336 1776 2368
rect 1808 2336 1848 2368
rect 1880 2336 1920 2368
rect 1952 2336 2000 2368
rect 0 2296 2000 2336
rect 0 2264 48 2296
rect 80 2264 120 2296
rect 152 2264 192 2296
rect 224 2264 264 2296
rect 296 2264 336 2296
rect 368 2264 408 2296
rect 440 2264 480 2296
rect 512 2264 552 2296
rect 584 2264 624 2296
rect 656 2264 696 2296
rect 728 2264 768 2296
rect 800 2264 840 2296
rect 872 2264 912 2296
rect 944 2264 984 2296
rect 1016 2264 1056 2296
rect 1088 2264 1128 2296
rect 1160 2264 1200 2296
rect 1232 2264 1272 2296
rect 1304 2264 1344 2296
rect 1376 2264 1416 2296
rect 1448 2264 1488 2296
rect 1520 2264 1560 2296
rect 1592 2264 1632 2296
rect 1664 2264 1704 2296
rect 1736 2264 1776 2296
rect 1808 2264 1848 2296
rect 1880 2264 1920 2296
rect 1952 2264 2000 2296
rect 0 2224 2000 2264
rect 0 2192 48 2224
rect 80 2192 120 2224
rect 152 2192 192 2224
rect 224 2192 264 2224
rect 296 2192 336 2224
rect 368 2192 408 2224
rect 440 2192 480 2224
rect 512 2192 552 2224
rect 584 2192 624 2224
rect 656 2192 696 2224
rect 728 2192 768 2224
rect 800 2192 840 2224
rect 872 2192 912 2224
rect 944 2192 984 2224
rect 1016 2192 1056 2224
rect 1088 2192 1128 2224
rect 1160 2192 1200 2224
rect 1232 2192 1272 2224
rect 1304 2192 1344 2224
rect 1376 2192 1416 2224
rect 1448 2192 1488 2224
rect 1520 2192 1560 2224
rect 1592 2192 1632 2224
rect 1664 2192 1704 2224
rect 1736 2192 1776 2224
rect 1808 2192 1848 2224
rect 1880 2192 1920 2224
rect 1952 2192 2000 2224
rect 0 2152 2000 2192
rect 0 2120 48 2152
rect 80 2120 120 2152
rect 152 2120 192 2152
rect 224 2120 264 2152
rect 296 2120 336 2152
rect 368 2120 408 2152
rect 440 2120 480 2152
rect 512 2120 552 2152
rect 584 2120 624 2152
rect 656 2120 696 2152
rect 728 2120 768 2152
rect 800 2120 840 2152
rect 872 2120 912 2152
rect 944 2120 984 2152
rect 1016 2120 1056 2152
rect 1088 2120 1128 2152
rect 1160 2120 1200 2152
rect 1232 2120 1272 2152
rect 1304 2120 1344 2152
rect 1376 2120 1416 2152
rect 1448 2120 1488 2152
rect 1520 2120 1560 2152
rect 1592 2120 1632 2152
rect 1664 2120 1704 2152
rect 1736 2120 1776 2152
rect 1808 2120 1848 2152
rect 1880 2120 1920 2152
rect 1952 2120 2000 2152
rect 0 2080 2000 2120
rect 0 2048 48 2080
rect 80 2048 120 2080
rect 152 2048 192 2080
rect 224 2048 264 2080
rect 296 2048 336 2080
rect 368 2048 408 2080
rect 440 2048 480 2080
rect 512 2048 552 2080
rect 584 2048 624 2080
rect 656 2048 696 2080
rect 728 2048 768 2080
rect 800 2048 840 2080
rect 872 2048 912 2080
rect 944 2048 984 2080
rect 1016 2048 1056 2080
rect 1088 2048 1128 2080
rect 1160 2048 1200 2080
rect 1232 2048 1272 2080
rect 1304 2048 1344 2080
rect 1376 2048 1416 2080
rect 1448 2048 1488 2080
rect 1520 2048 1560 2080
rect 1592 2048 1632 2080
rect 1664 2048 1704 2080
rect 1736 2048 1776 2080
rect 1808 2048 1848 2080
rect 1880 2048 1920 2080
rect 1952 2048 2000 2080
rect 0 2008 2000 2048
rect 0 1976 48 2008
rect 80 1976 120 2008
rect 152 1976 192 2008
rect 224 1976 264 2008
rect 296 1976 336 2008
rect 368 1976 408 2008
rect 440 1976 480 2008
rect 512 1976 552 2008
rect 584 1976 624 2008
rect 656 1976 696 2008
rect 728 1976 768 2008
rect 800 1976 840 2008
rect 872 1976 912 2008
rect 944 1976 984 2008
rect 1016 1976 1056 2008
rect 1088 1976 1128 2008
rect 1160 1976 1200 2008
rect 1232 1976 1272 2008
rect 1304 1976 1344 2008
rect 1376 1976 1416 2008
rect 1448 1976 1488 2008
rect 1520 1976 1560 2008
rect 1592 1976 1632 2008
rect 1664 1976 1704 2008
rect 1736 1976 1776 2008
rect 1808 1976 1848 2008
rect 1880 1976 1920 2008
rect 1952 1976 2000 2008
rect 0 1936 2000 1976
rect 0 1904 48 1936
rect 80 1904 120 1936
rect 152 1904 192 1936
rect 224 1904 264 1936
rect 296 1904 336 1936
rect 368 1904 408 1936
rect 440 1904 480 1936
rect 512 1904 552 1936
rect 584 1904 624 1936
rect 656 1904 696 1936
rect 728 1904 768 1936
rect 800 1904 840 1936
rect 872 1904 912 1936
rect 944 1904 984 1936
rect 1016 1904 1056 1936
rect 1088 1904 1128 1936
rect 1160 1904 1200 1936
rect 1232 1904 1272 1936
rect 1304 1904 1344 1936
rect 1376 1904 1416 1936
rect 1448 1904 1488 1936
rect 1520 1904 1560 1936
rect 1592 1904 1632 1936
rect 1664 1904 1704 1936
rect 1736 1904 1776 1936
rect 1808 1904 1848 1936
rect 1880 1904 1920 1936
rect 1952 1904 2000 1936
rect 0 1864 2000 1904
rect 0 1832 48 1864
rect 80 1832 120 1864
rect 152 1832 192 1864
rect 224 1832 264 1864
rect 296 1832 336 1864
rect 368 1832 408 1864
rect 440 1832 480 1864
rect 512 1832 552 1864
rect 584 1832 624 1864
rect 656 1832 696 1864
rect 728 1832 768 1864
rect 800 1832 840 1864
rect 872 1832 912 1864
rect 944 1832 984 1864
rect 1016 1832 1056 1864
rect 1088 1832 1128 1864
rect 1160 1832 1200 1864
rect 1232 1832 1272 1864
rect 1304 1832 1344 1864
rect 1376 1832 1416 1864
rect 1448 1832 1488 1864
rect 1520 1832 1560 1864
rect 1592 1832 1632 1864
rect 1664 1832 1704 1864
rect 1736 1832 1776 1864
rect 1808 1832 1848 1864
rect 1880 1832 1920 1864
rect 1952 1832 2000 1864
rect 0 1792 2000 1832
rect 0 1760 48 1792
rect 80 1760 120 1792
rect 152 1760 192 1792
rect 224 1760 264 1792
rect 296 1760 336 1792
rect 368 1760 408 1792
rect 440 1760 480 1792
rect 512 1760 552 1792
rect 584 1760 624 1792
rect 656 1760 696 1792
rect 728 1760 768 1792
rect 800 1760 840 1792
rect 872 1760 912 1792
rect 944 1760 984 1792
rect 1016 1760 1056 1792
rect 1088 1760 1128 1792
rect 1160 1760 1200 1792
rect 1232 1760 1272 1792
rect 1304 1760 1344 1792
rect 1376 1760 1416 1792
rect 1448 1760 1488 1792
rect 1520 1760 1560 1792
rect 1592 1760 1632 1792
rect 1664 1760 1704 1792
rect 1736 1760 1776 1792
rect 1808 1760 1848 1792
rect 1880 1760 1920 1792
rect 1952 1760 2000 1792
rect 0 1720 2000 1760
rect 0 1688 48 1720
rect 80 1688 120 1720
rect 152 1688 192 1720
rect 224 1688 264 1720
rect 296 1688 336 1720
rect 368 1688 408 1720
rect 440 1688 480 1720
rect 512 1688 552 1720
rect 584 1688 624 1720
rect 656 1688 696 1720
rect 728 1688 768 1720
rect 800 1688 840 1720
rect 872 1688 912 1720
rect 944 1688 984 1720
rect 1016 1688 1056 1720
rect 1088 1688 1128 1720
rect 1160 1688 1200 1720
rect 1232 1688 1272 1720
rect 1304 1688 1344 1720
rect 1376 1688 1416 1720
rect 1448 1688 1488 1720
rect 1520 1688 1560 1720
rect 1592 1688 1632 1720
rect 1664 1688 1704 1720
rect 1736 1688 1776 1720
rect 1808 1688 1848 1720
rect 1880 1688 1920 1720
rect 1952 1688 2000 1720
rect 0 1648 2000 1688
rect 0 1616 48 1648
rect 80 1616 120 1648
rect 152 1616 192 1648
rect 224 1616 264 1648
rect 296 1616 336 1648
rect 368 1616 408 1648
rect 440 1616 480 1648
rect 512 1616 552 1648
rect 584 1616 624 1648
rect 656 1616 696 1648
rect 728 1616 768 1648
rect 800 1616 840 1648
rect 872 1616 912 1648
rect 944 1616 984 1648
rect 1016 1616 1056 1648
rect 1088 1616 1128 1648
rect 1160 1616 1200 1648
rect 1232 1616 1272 1648
rect 1304 1616 1344 1648
rect 1376 1616 1416 1648
rect 1448 1616 1488 1648
rect 1520 1616 1560 1648
rect 1592 1616 1632 1648
rect 1664 1616 1704 1648
rect 1736 1616 1776 1648
rect 1808 1616 1848 1648
rect 1880 1616 1920 1648
rect 1952 1616 2000 1648
rect 0 1576 2000 1616
rect 0 1544 48 1576
rect 80 1544 120 1576
rect 152 1544 192 1576
rect 224 1544 264 1576
rect 296 1544 336 1576
rect 368 1544 408 1576
rect 440 1544 480 1576
rect 512 1544 552 1576
rect 584 1544 624 1576
rect 656 1544 696 1576
rect 728 1544 768 1576
rect 800 1544 840 1576
rect 872 1544 912 1576
rect 944 1544 984 1576
rect 1016 1544 1056 1576
rect 1088 1544 1128 1576
rect 1160 1544 1200 1576
rect 1232 1544 1272 1576
rect 1304 1544 1344 1576
rect 1376 1544 1416 1576
rect 1448 1544 1488 1576
rect 1520 1544 1560 1576
rect 1592 1544 1632 1576
rect 1664 1544 1704 1576
rect 1736 1544 1776 1576
rect 1808 1544 1848 1576
rect 1880 1544 1920 1576
rect 1952 1544 2000 1576
rect 0 1504 2000 1544
rect 0 1472 48 1504
rect 80 1472 120 1504
rect 152 1472 192 1504
rect 224 1472 264 1504
rect 296 1472 336 1504
rect 368 1472 408 1504
rect 440 1472 480 1504
rect 512 1472 552 1504
rect 584 1472 624 1504
rect 656 1472 696 1504
rect 728 1472 768 1504
rect 800 1472 840 1504
rect 872 1472 912 1504
rect 944 1472 984 1504
rect 1016 1472 1056 1504
rect 1088 1472 1128 1504
rect 1160 1472 1200 1504
rect 1232 1472 1272 1504
rect 1304 1472 1344 1504
rect 1376 1472 1416 1504
rect 1448 1472 1488 1504
rect 1520 1472 1560 1504
rect 1592 1472 1632 1504
rect 1664 1472 1704 1504
rect 1736 1472 1776 1504
rect 1808 1472 1848 1504
rect 1880 1472 1920 1504
rect 1952 1472 2000 1504
rect 0 1432 2000 1472
rect 0 1400 48 1432
rect 80 1400 120 1432
rect 152 1400 192 1432
rect 224 1400 264 1432
rect 296 1400 336 1432
rect 368 1400 408 1432
rect 440 1400 480 1432
rect 512 1400 552 1432
rect 584 1400 624 1432
rect 656 1400 696 1432
rect 728 1400 768 1432
rect 800 1400 840 1432
rect 872 1400 912 1432
rect 944 1400 984 1432
rect 1016 1400 1056 1432
rect 1088 1400 1128 1432
rect 1160 1400 1200 1432
rect 1232 1400 1272 1432
rect 1304 1400 1344 1432
rect 1376 1400 1416 1432
rect 1448 1400 1488 1432
rect 1520 1400 1560 1432
rect 1592 1400 1632 1432
rect 1664 1400 1704 1432
rect 1736 1400 1776 1432
rect 1808 1400 1848 1432
rect 1880 1400 1920 1432
rect 1952 1400 2000 1432
rect 0 1360 2000 1400
rect 0 1328 48 1360
rect 80 1328 120 1360
rect 152 1328 192 1360
rect 224 1328 264 1360
rect 296 1328 336 1360
rect 368 1328 408 1360
rect 440 1328 480 1360
rect 512 1328 552 1360
rect 584 1328 624 1360
rect 656 1328 696 1360
rect 728 1328 768 1360
rect 800 1328 840 1360
rect 872 1328 912 1360
rect 944 1328 984 1360
rect 1016 1328 1056 1360
rect 1088 1328 1128 1360
rect 1160 1328 1200 1360
rect 1232 1328 1272 1360
rect 1304 1328 1344 1360
rect 1376 1328 1416 1360
rect 1448 1328 1488 1360
rect 1520 1328 1560 1360
rect 1592 1328 1632 1360
rect 1664 1328 1704 1360
rect 1736 1328 1776 1360
rect 1808 1328 1848 1360
rect 1880 1328 1920 1360
rect 1952 1328 2000 1360
rect 0 1288 2000 1328
rect 0 1256 48 1288
rect 80 1256 120 1288
rect 152 1256 192 1288
rect 224 1256 264 1288
rect 296 1256 336 1288
rect 368 1256 408 1288
rect 440 1256 480 1288
rect 512 1256 552 1288
rect 584 1256 624 1288
rect 656 1256 696 1288
rect 728 1256 768 1288
rect 800 1256 840 1288
rect 872 1256 912 1288
rect 944 1256 984 1288
rect 1016 1256 1056 1288
rect 1088 1256 1128 1288
rect 1160 1256 1200 1288
rect 1232 1256 1272 1288
rect 1304 1256 1344 1288
rect 1376 1256 1416 1288
rect 1448 1256 1488 1288
rect 1520 1256 1560 1288
rect 1592 1256 1632 1288
rect 1664 1256 1704 1288
rect 1736 1256 1776 1288
rect 1808 1256 1848 1288
rect 1880 1256 1920 1288
rect 1952 1256 2000 1288
rect 0 1200 2000 1256
<< metal3 >>
rect 0 32000 2000 35600
rect 0 28000 2000 31600
rect 0 25200 2000 26800
rect 0 18700 2000 23800
rect 0 13200 2000 18300
rect 0 6900 2000 12000
rect 0 1400 2000 6500
<< metal4 >>
rect 0 32440 2000 35600
rect 0 28000 2000 31160
rect 0 25200 2000 26800
rect 0 18700 2000 23800
rect 0 13200 2000 18300
rect 0 6900 2000 12000
rect 0 1400 2000 6500
<< metal5 >>
rect 0 32000 2000 35600
rect 0 28000 2000 31600
rect 0 25200 2000 26800
rect 0 18700 2000 23800
rect 0 13200 2000 18300
rect 0 6900 2000 12000
rect 0 1400 2000 6500
<< metal6 >>
rect 0 32000 2000 35600
rect 0 28000 2000 31600
rect 0 25200 2000 26800
rect 0 18700 2000 23800
rect 0 13200 2000 18300
rect 0 6900 2000 12000
rect 0 1400 2000 6500
<< metal7 >>
rect 0 25500 2000 26500
rect 0 19000 2000 23500
rect 0 13500 2000 18000
rect 0 7200 2000 11700
rect 0 1700 2000 6200
<< labels >>
rlabel metal3 s 0 32000 2000 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 2000 31600 4 vss
port 1 nsew
rlabel metal3 s 0 18700 2000 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 13200 2000 18300 4 iovdd
port 4 nsew
rlabel metal3 s 0 6900 2000 12000 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 2000 6500 4 iovss
port 3 nsew
rlabel metal3 s 0 25200 2000 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 2000 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 2000 35600 4 vss
port 1 nsew
rlabel metal4 s 0 18700 2000 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 13200 2000 18300 4 iovdd
port 4 nsew
rlabel metal4 s 0 6900 2000 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 2000 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 25200 2000 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 2000 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 2000 35600 4 vss
port 1 nsew
rlabel metal5 s 0 18700 2000 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 13200 2000 18300 4 iovdd
port 4 nsew
rlabel metal5 s 0 6900 2000 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 2000 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 25200 2000 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 2000 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 2000 35600 4 vss
port 1 nsew
rlabel metal6 s 0 18700 2000 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 13200 2000 18300 4 iovdd
port 4 nsew
rlabel metal6 s 0 6900 2000 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 2000 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 25200 2000 26800 4 iovss
port 3 nsew
rlabel metal7 s 0 19000 2000 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 13500 2000 18000 4 iovdd
port 4 nsew
rlabel metal7 s 0 25500 2000 26500 4 iovss
port 3 nsew
rlabel metal7 s 0 7200 2000 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 1700 2000 6200 4 iovss
port 3 nsew
flabel comment s 1010 31400 1010 31400 0 FreeSans 400 0 0 0 sub!
flabel comment s 359 17636 359 17636 0 FreeSans 400 0 0 0 sub!
flabel comment s 353 22637 353 22637 0 FreeSans 400 0 0 0 sub!
flabel comment s 408 27723 408 27723 0 FreeSans 400 0 0 0 sub!
flabel metal1 s 659 31384 749 31416 0 FreeSans 400 0 0 0 vss
port 1 nsew
flabel metal1 s 225 6176 485 6389 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 256 11768 501 11981 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 488 17550 728 17654 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 488 22532 728 22636 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 488 27795 728 27899 0 FreeSans 400 0 0 0 iovss
port 3 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 2000 36000
string GDS_END 64440556
string GDS_FILE sg13g2_io.gds
string GDS_START 63852652
<< end >>
