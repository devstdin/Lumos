magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -924 3124 37600
<< isosubstrate >>
rect 50 23124 950 28034
rect 50 18112 950 22924
rect 50 13000 950 17912
<< nwell >>
rect -124 33246 1124 33554
rect -124 29546 1124 29854
rect -124 1076 1124 12324
<< pwell >>
rect 18 31344 982 31456
rect 24 12974 976 28060
<< psubdiff >>
rect 292 31384 324 31416
rect 362 31384 394 31416
rect 431 31384 463 31416
rect 502 31384 534 31416
rect 572 31384 604 31416
rect 640 31384 672 31416
rect 710 31384 742 31416
rect 196 27939 228 27971
rect 268 27939 300 27971
rect 340 27939 372 27971
rect 412 27939 444 27971
rect 484 27939 516 27971
rect 556 27939 588 27971
rect 628 27939 660 27971
rect 700 27939 732 27971
rect 772 27939 804 27971
rect 844 27939 876 27971
rect 124 27867 156 27899
rect 196 27867 228 27899
rect 268 27867 300 27899
rect 340 27867 372 27899
rect 412 27867 444 27899
rect 484 27867 516 27899
rect 556 27867 588 27899
rect 628 27867 660 27899
rect 700 27867 732 27899
rect 772 27867 804 27899
rect 844 27867 876 27899
rect 124 27795 156 27827
rect 196 27795 228 27827
rect 268 27795 300 27827
rect 340 27795 372 27827
rect 412 27795 444 27827
rect 484 27795 516 27827
rect 556 27795 588 27827
rect 628 27795 660 27827
rect 700 27795 732 27827
rect 772 27795 804 27827
rect 844 27795 876 27827
rect 124 27723 156 27755
rect 196 27723 228 27755
rect 268 27723 300 27755
rect 340 27723 372 27755
rect 412 27723 444 27755
rect 484 27723 516 27755
rect 556 27723 588 27755
rect 628 27723 660 27755
rect 700 27723 732 27755
rect 772 27723 804 27755
rect 844 27723 876 27755
rect 124 27651 156 27683
rect 196 27651 228 27683
rect 268 27651 300 27683
rect 340 27651 372 27683
rect 412 27651 444 27683
rect 484 27651 516 27683
rect 556 27651 588 27683
rect 628 27651 660 27683
rect 700 27651 732 27683
rect 772 27651 804 27683
rect 844 27651 876 27683
rect 124 27579 156 27611
rect 196 27579 228 27611
rect 268 27579 300 27611
rect 340 27579 372 27611
rect 412 27579 444 27611
rect 484 27579 516 27611
rect 556 27579 588 27611
rect 628 27579 660 27611
rect 700 27579 732 27611
rect 772 27579 804 27611
rect 844 27579 876 27611
rect 124 27507 156 27539
rect 196 27507 228 27539
rect 268 27507 300 27539
rect 340 27507 372 27539
rect 412 27507 444 27539
rect 484 27507 516 27539
rect 556 27507 588 27539
rect 628 27507 660 27539
rect 700 27507 732 27539
rect 772 27507 804 27539
rect 844 27507 876 27539
rect 124 27435 156 27467
rect 196 27435 228 27467
rect 268 27435 300 27467
rect 340 27435 372 27467
rect 412 27435 444 27467
rect 484 27435 516 27467
rect 556 27435 588 27467
rect 628 27435 660 27467
rect 700 27435 732 27467
rect 772 27435 804 27467
rect 844 27435 876 27467
rect 124 27363 156 27395
rect 196 27363 228 27395
rect 268 27363 300 27395
rect 340 27363 372 27395
rect 412 27363 444 27395
rect 484 27363 516 27395
rect 556 27363 588 27395
rect 628 27363 660 27395
rect 700 27363 732 27395
rect 772 27363 804 27395
rect 844 27363 876 27395
rect 124 27291 156 27323
rect 196 27291 228 27323
rect 268 27291 300 27323
rect 340 27291 372 27323
rect 412 27291 444 27323
rect 484 27291 516 27323
rect 556 27291 588 27323
rect 628 27291 660 27323
rect 700 27291 732 27323
rect 772 27291 804 27323
rect 844 27291 876 27323
rect 124 27219 156 27251
rect 196 27219 228 27251
rect 268 27219 300 27251
rect 340 27219 372 27251
rect 412 27219 444 27251
rect 484 27219 516 27251
rect 556 27219 588 27251
rect 628 27219 660 27251
rect 700 27219 732 27251
rect 772 27219 804 27251
rect 844 27219 876 27251
rect 124 27147 156 27179
rect 196 27147 228 27179
rect 268 27147 300 27179
rect 340 27147 372 27179
rect 412 27147 444 27179
rect 484 27147 516 27179
rect 556 27147 588 27179
rect 628 27147 660 27179
rect 700 27147 732 27179
rect 772 27147 804 27179
rect 844 27147 876 27179
rect 124 27075 156 27107
rect 196 27075 228 27107
rect 268 27075 300 27107
rect 340 27075 372 27107
rect 412 27075 444 27107
rect 484 27075 516 27107
rect 556 27075 588 27107
rect 628 27075 660 27107
rect 700 27075 732 27107
rect 772 27075 804 27107
rect 844 27075 876 27107
rect 124 27003 156 27035
rect 196 27003 228 27035
rect 268 27003 300 27035
rect 340 27003 372 27035
rect 412 27003 444 27035
rect 484 27003 516 27035
rect 556 27003 588 27035
rect 628 27003 660 27035
rect 700 27003 732 27035
rect 772 27003 804 27035
rect 844 27003 876 27035
rect 124 26931 156 26963
rect 196 26931 228 26963
rect 268 26931 300 26963
rect 340 26931 372 26963
rect 412 26931 444 26963
rect 484 26931 516 26963
rect 556 26931 588 26963
rect 628 26931 660 26963
rect 700 26931 732 26963
rect 772 26931 804 26963
rect 844 26931 876 26963
rect 124 26859 156 26891
rect 196 26859 228 26891
rect 268 26859 300 26891
rect 340 26859 372 26891
rect 412 26859 444 26891
rect 484 26859 516 26891
rect 556 26859 588 26891
rect 628 26859 660 26891
rect 700 26859 732 26891
rect 772 26859 804 26891
rect 844 26859 876 26891
rect 124 26787 156 26819
rect 196 26787 228 26819
rect 268 26787 300 26819
rect 340 26787 372 26819
rect 412 26787 444 26819
rect 484 26787 516 26819
rect 556 26787 588 26819
rect 628 26787 660 26819
rect 700 26787 732 26819
rect 772 26787 804 26819
rect 844 26787 876 26819
rect 124 26715 156 26747
rect 196 26715 228 26747
rect 268 26715 300 26747
rect 340 26715 372 26747
rect 412 26715 444 26747
rect 484 26715 516 26747
rect 556 26715 588 26747
rect 628 26715 660 26747
rect 700 26715 732 26747
rect 772 26715 804 26747
rect 844 26715 876 26747
rect 124 26643 156 26675
rect 196 26643 228 26675
rect 268 26643 300 26675
rect 340 26643 372 26675
rect 412 26643 444 26675
rect 484 26643 516 26675
rect 556 26643 588 26675
rect 628 26643 660 26675
rect 700 26643 732 26675
rect 772 26643 804 26675
rect 844 26643 876 26675
rect 124 26571 156 26603
rect 196 26571 228 26603
rect 268 26571 300 26603
rect 340 26571 372 26603
rect 412 26571 444 26603
rect 484 26571 516 26603
rect 556 26571 588 26603
rect 628 26571 660 26603
rect 700 26571 732 26603
rect 772 26571 804 26603
rect 844 26571 876 26603
rect 124 26499 156 26531
rect 196 26499 228 26531
rect 268 26499 300 26531
rect 340 26499 372 26531
rect 412 26499 444 26531
rect 484 26499 516 26531
rect 556 26499 588 26531
rect 628 26499 660 26531
rect 700 26499 732 26531
rect 772 26499 804 26531
rect 844 26499 876 26531
rect 124 26427 156 26459
rect 196 26427 228 26459
rect 268 26427 300 26459
rect 340 26427 372 26459
rect 412 26427 444 26459
rect 484 26427 516 26459
rect 556 26427 588 26459
rect 628 26427 660 26459
rect 700 26427 732 26459
rect 772 26427 804 26459
rect 844 26427 876 26459
rect 124 26355 156 26387
rect 196 26355 228 26387
rect 268 26355 300 26387
rect 340 26355 372 26387
rect 412 26355 444 26387
rect 484 26355 516 26387
rect 556 26355 588 26387
rect 628 26355 660 26387
rect 700 26355 732 26387
rect 772 26355 804 26387
rect 844 26355 876 26387
rect 124 26283 156 26315
rect 196 26283 228 26315
rect 268 26283 300 26315
rect 340 26283 372 26315
rect 412 26283 444 26315
rect 484 26283 516 26315
rect 556 26283 588 26315
rect 628 26283 660 26315
rect 700 26283 732 26315
rect 772 26283 804 26315
rect 844 26283 876 26315
rect 124 26211 156 26243
rect 196 26211 228 26243
rect 268 26211 300 26243
rect 340 26211 372 26243
rect 412 26211 444 26243
rect 484 26211 516 26243
rect 556 26211 588 26243
rect 628 26211 660 26243
rect 700 26211 732 26243
rect 772 26211 804 26243
rect 844 26211 876 26243
rect 124 26139 156 26171
rect 196 26139 228 26171
rect 268 26139 300 26171
rect 340 26139 372 26171
rect 412 26139 444 26171
rect 484 26139 516 26171
rect 556 26139 588 26171
rect 628 26139 660 26171
rect 700 26139 732 26171
rect 772 26139 804 26171
rect 844 26139 876 26171
rect 124 26067 156 26099
rect 196 26067 228 26099
rect 268 26067 300 26099
rect 340 26067 372 26099
rect 412 26067 444 26099
rect 484 26067 516 26099
rect 556 26067 588 26099
rect 628 26067 660 26099
rect 700 26067 732 26099
rect 772 26067 804 26099
rect 844 26067 876 26099
rect 124 25995 156 26027
rect 196 25995 228 26027
rect 268 25995 300 26027
rect 340 25995 372 26027
rect 412 25995 444 26027
rect 484 25995 516 26027
rect 556 25995 588 26027
rect 628 25995 660 26027
rect 700 25995 732 26027
rect 772 25995 804 26027
rect 844 25995 876 26027
rect 124 25923 156 25955
rect 196 25923 228 25955
rect 268 25923 300 25955
rect 340 25923 372 25955
rect 412 25923 444 25955
rect 484 25923 516 25955
rect 556 25923 588 25955
rect 628 25923 660 25955
rect 700 25923 732 25955
rect 772 25923 804 25955
rect 844 25923 876 25955
rect 124 25851 156 25883
rect 196 25851 228 25883
rect 268 25851 300 25883
rect 340 25851 372 25883
rect 412 25851 444 25883
rect 484 25851 516 25883
rect 556 25851 588 25883
rect 628 25851 660 25883
rect 700 25851 732 25883
rect 772 25851 804 25883
rect 844 25851 876 25883
rect 124 25779 156 25811
rect 196 25779 228 25811
rect 268 25779 300 25811
rect 340 25779 372 25811
rect 412 25779 444 25811
rect 484 25779 516 25811
rect 556 25779 588 25811
rect 628 25779 660 25811
rect 700 25779 732 25811
rect 772 25779 804 25811
rect 844 25779 876 25811
rect 124 25707 156 25739
rect 196 25707 228 25739
rect 268 25707 300 25739
rect 340 25707 372 25739
rect 412 25707 444 25739
rect 484 25707 516 25739
rect 556 25707 588 25739
rect 628 25707 660 25739
rect 700 25707 732 25739
rect 772 25707 804 25739
rect 844 25707 876 25739
rect 124 25635 156 25667
rect 196 25635 228 25667
rect 268 25635 300 25667
rect 340 25635 372 25667
rect 412 25635 444 25667
rect 484 25635 516 25667
rect 556 25635 588 25667
rect 628 25635 660 25667
rect 700 25635 732 25667
rect 772 25635 804 25667
rect 844 25635 876 25667
rect 124 25563 156 25595
rect 196 25563 228 25595
rect 268 25563 300 25595
rect 340 25563 372 25595
rect 412 25563 444 25595
rect 484 25563 516 25595
rect 556 25563 588 25595
rect 628 25563 660 25595
rect 700 25563 732 25595
rect 772 25563 804 25595
rect 844 25563 876 25595
rect 124 25491 156 25523
rect 196 25491 228 25523
rect 268 25491 300 25523
rect 340 25491 372 25523
rect 412 25491 444 25523
rect 484 25491 516 25523
rect 556 25491 588 25523
rect 628 25491 660 25523
rect 700 25491 732 25523
rect 772 25491 804 25523
rect 844 25491 876 25523
rect 124 25419 156 25451
rect 196 25419 228 25451
rect 268 25419 300 25451
rect 340 25419 372 25451
rect 412 25419 444 25451
rect 484 25419 516 25451
rect 556 25419 588 25451
rect 628 25419 660 25451
rect 700 25419 732 25451
rect 772 25419 804 25451
rect 844 25419 876 25451
rect 124 25347 156 25379
rect 196 25347 228 25379
rect 268 25347 300 25379
rect 340 25347 372 25379
rect 412 25347 444 25379
rect 484 25347 516 25379
rect 556 25347 588 25379
rect 628 25347 660 25379
rect 700 25347 732 25379
rect 772 25347 804 25379
rect 844 25347 876 25379
rect 124 25275 156 25307
rect 196 25275 228 25307
rect 268 25275 300 25307
rect 340 25275 372 25307
rect 412 25275 444 25307
rect 484 25275 516 25307
rect 556 25275 588 25307
rect 628 25275 660 25307
rect 700 25275 732 25307
rect 772 25275 804 25307
rect 844 25275 876 25307
rect 124 25203 156 25235
rect 196 25203 228 25235
rect 268 25203 300 25235
rect 340 25203 372 25235
rect 412 25203 444 25235
rect 484 25203 516 25235
rect 556 25203 588 25235
rect 628 25203 660 25235
rect 700 25203 732 25235
rect 772 25203 804 25235
rect 844 25203 876 25235
rect 124 25131 156 25163
rect 196 25131 228 25163
rect 268 25131 300 25163
rect 340 25131 372 25163
rect 412 25131 444 25163
rect 484 25131 516 25163
rect 556 25131 588 25163
rect 628 25131 660 25163
rect 700 25131 732 25163
rect 772 25131 804 25163
rect 844 25131 876 25163
rect 124 25059 156 25091
rect 196 25059 228 25091
rect 268 25059 300 25091
rect 340 25059 372 25091
rect 412 25059 444 25091
rect 484 25059 516 25091
rect 556 25059 588 25091
rect 628 25059 660 25091
rect 700 25059 732 25091
rect 772 25059 804 25091
rect 844 25059 876 25091
rect 124 24987 156 25019
rect 196 24987 228 25019
rect 268 24987 300 25019
rect 340 24987 372 25019
rect 412 24987 444 25019
rect 484 24987 516 25019
rect 556 24987 588 25019
rect 628 24987 660 25019
rect 700 24987 732 25019
rect 772 24987 804 25019
rect 844 24987 876 25019
rect 124 24915 156 24947
rect 196 24915 228 24947
rect 268 24915 300 24947
rect 340 24915 372 24947
rect 412 24915 444 24947
rect 484 24915 516 24947
rect 556 24915 588 24947
rect 628 24915 660 24947
rect 700 24915 732 24947
rect 772 24915 804 24947
rect 844 24915 876 24947
rect 124 24843 156 24875
rect 196 24843 228 24875
rect 268 24843 300 24875
rect 340 24843 372 24875
rect 412 24843 444 24875
rect 484 24843 516 24875
rect 556 24843 588 24875
rect 628 24843 660 24875
rect 700 24843 732 24875
rect 772 24843 804 24875
rect 844 24843 876 24875
rect 124 24771 156 24803
rect 196 24771 228 24803
rect 268 24771 300 24803
rect 340 24771 372 24803
rect 412 24771 444 24803
rect 484 24771 516 24803
rect 556 24771 588 24803
rect 628 24771 660 24803
rect 700 24771 732 24803
rect 772 24771 804 24803
rect 844 24771 876 24803
rect 124 24699 156 24731
rect 196 24699 228 24731
rect 268 24699 300 24731
rect 340 24699 372 24731
rect 412 24699 444 24731
rect 484 24699 516 24731
rect 556 24699 588 24731
rect 628 24699 660 24731
rect 700 24699 732 24731
rect 772 24699 804 24731
rect 844 24699 876 24731
rect 124 24627 156 24659
rect 196 24627 228 24659
rect 268 24627 300 24659
rect 340 24627 372 24659
rect 412 24627 444 24659
rect 484 24627 516 24659
rect 556 24627 588 24659
rect 628 24627 660 24659
rect 700 24627 732 24659
rect 772 24627 804 24659
rect 844 24627 876 24659
rect 124 24555 156 24587
rect 196 24555 228 24587
rect 268 24555 300 24587
rect 340 24555 372 24587
rect 412 24555 444 24587
rect 484 24555 516 24587
rect 556 24555 588 24587
rect 628 24555 660 24587
rect 700 24555 732 24587
rect 772 24555 804 24587
rect 844 24555 876 24587
rect 124 24483 156 24515
rect 196 24483 228 24515
rect 268 24483 300 24515
rect 340 24483 372 24515
rect 412 24483 444 24515
rect 484 24483 516 24515
rect 556 24483 588 24515
rect 628 24483 660 24515
rect 700 24483 732 24515
rect 772 24483 804 24515
rect 844 24483 876 24515
rect 124 24411 156 24443
rect 196 24411 228 24443
rect 268 24411 300 24443
rect 340 24411 372 24443
rect 412 24411 444 24443
rect 484 24411 516 24443
rect 556 24411 588 24443
rect 628 24411 660 24443
rect 700 24411 732 24443
rect 772 24411 804 24443
rect 844 24411 876 24443
rect 124 24339 156 24371
rect 196 24339 228 24371
rect 268 24339 300 24371
rect 340 24339 372 24371
rect 412 24339 444 24371
rect 484 24339 516 24371
rect 556 24339 588 24371
rect 628 24339 660 24371
rect 700 24339 732 24371
rect 772 24339 804 24371
rect 844 24339 876 24371
rect 124 24267 156 24299
rect 196 24267 228 24299
rect 268 24267 300 24299
rect 340 24267 372 24299
rect 412 24267 444 24299
rect 484 24267 516 24299
rect 556 24267 588 24299
rect 628 24267 660 24299
rect 700 24267 732 24299
rect 772 24267 804 24299
rect 844 24267 876 24299
rect 124 24195 156 24227
rect 196 24195 228 24227
rect 268 24195 300 24227
rect 340 24195 372 24227
rect 412 24195 444 24227
rect 484 24195 516 24227
rect 556 24195 588 24227
rect 628 24195 660 24227
rect 700 24195 732 24227
rect 772 24195 804 24227
rect 844 24195 876 24227
rect 124 24123 156 24155
rect 196 24123 228 24155
rect 268 24123 300 24155
rect 340 24123 372 24155
rect 412 24123 444 24155
rect 484 24123 516 24155
rect 556 24123 588 24155
rect 628 24123 660 24155
rect 700 24123 732 24155
rect 772 24123 804 24155
rect 844 24123 876 24155
rect 124 24051 156 24083
rect 196 24051 228 24083
rect 268 24051 300 24083
rect 340 24051 372 24083
rect 412 24051 444 24083
rect 484 24051 516 24083
rect 556 24051 588 24083
rect 628 24051 660 24083
rect 700 24051 732 24083
rect 772 24051 804 24083
rect 844 24051 876 24083
rect 124 23979 156 24011
rect 196 23979 228 24011
rect 268 23979 300 24011
rect 340 23979 372 24011
rect 412 23979 444 24011
rect 484 23979 516 24011
rect 556 23979 588 24011
rect 628 23979 660 24011
rect 700 23979 732 24011
rect 772 23979 804 24011
rect 844 23979 876 24011
rect 124 23907 156 23939
rect 196 23907 228 23939
rect 268 23907 300 23939
rect 340 23907 372 23939
rect 412 23907 444 23939
rect 484 23907 516 23939
rect 556 23907 588 23939
rect 628 23907 660 23939
rect 700 23907 732 23939
rect 772 23907 804 23939
rect 844 23907 876 23939
rect 124 23835 156 23867
rect 196 23835 228 23867
rect 268 23835 300 23867
rect 340 23835 372 23867
rect 412 23835 444 23867
rect 484 23835 516 23867
rect 556 23835 588 23867
rect 628 23835 660 23867
rect 700 23835 732 23867
rect 772 23835 804 23867
rect 844 23835 876 23867
rect 124 23763 156 23795
rect 196 23763 228 23795
rect 268 23763 300 23795
rect 340 23763 372 23795
rect 412 23763 444 23795
rect 484 23763 516 23795
rect 556 23763 588 23795
rect 628 23763 660 23795
rect 700 23763 732 23795
rect 772 23763 804 23795
rect 844 23763 876 23795
rect 124 23691 156 23723
rect 196 23691 228 23723
rect 268 23691 300 23723
rect 340 23691 372 23723
rect 412 23691 444 23723
rect 484 23691 516 23723
rect 556 23691 588 23723
rect 628 23691 660 23723
rect 700 23691 732 23723
rect 772 23691 804 23723
rect 844 23691 876 23723
rect 124 23619 156 23651
rect 196 23619 228 23651
rect 268 23619 300 23651
rect 340 23619 372 23651
rect 412 23619 444 23651
rect 484 23619 516 23651
rect 556 23619 588 23651
rect 628 23619 660 23651
rect 700 23619 732 23651
rect 772 23619 804 23651
rect 844 23619 876 23651
rect 124 23547 156 23579
rect 196 23547 228 23579
rect 268 23547 300 23579
rect 340 23547 372 23579
rect 412 23547 444 23579
rect 484 23547 516 23579
rect 556 23547 588 23579
rect 628 23547 660 23579
rect 700 23547 732 23579
rect 772 23547 804 23579
rect 844 23547 876 23579
rect 124 23475 156 23507
rect 196 23475 228 23507
rect 268 23475 300 23507
rect 340 23475 372 23507
rect 412 23475 444 23507
rect 484 23475 516 23507
rect 556 23475 588 23507
rect 628 23475 660 23507
rect 700 23475 732 23507
rect 772 23475 804 23507
rect 844 23475 876 23507
rect 124 23403 156 23435
rect 196 23403 228 23435
rect 268 23403 300 23435
rect 340 23403 372 23435
rect 412 23403 444 23435
rect 484 23403 516 23435
rect 556 23403 588 23435
rect 628 23403 660 23435
rect 700 23403 732 23435
rect 772 23403 804 23435
rect 844 23403 876 23435
rect 124 23331 156 23363
rect 196 23331 228 23363
rect 268 23331 300 23363
rect 340 23331 372 23363
rect 412 23331 444 23363
rect 484 23331 516 23363
rect 556 23331 588 23363
rect 628 23331 660 23363
rect 700 23331 732 23363
rect 772 23331 804 23363
rect 844 23331 876 23363
rect 124 23259 156 23291
rect 196 23259 228 23291
rect 268 23259 300 23291
rect 340 23259 372 23291
rect 412 23259 444 23291
rect 484 23259 516 23291
rect 556 23259 588 23291
rect 628 23259 660 23291
rect 700 23259 732 23291
rect 772 23259 804 23291
rect 844 23259 876 23291
rect 124 23187 156 23219
rect 196 23187 228 23219
rect 268 23187 300 23219
rect 340 23187 372 23219
rect 412 23187 444 23219
rect 484 23187 516 23219
rect 556 23187 588 23219
rect 628 23187 660 23219
rect 700 23187 732 23219
rect 772 23187 804 23219
rect 844 23187 876 23219
rect 196 22842 228 22874
rect 268 22842 300 22874
rect 340 22842 372 22874
rect 412 22842 444 22874
rect 484 22842 516 22874
rect 556 22842 588 22874
rect 628 22842 660 22874
rect 700 22842 732 22874
rect 772 22842 804 22874
rect 844 22842 876 22874
rect 124 22770 156 22802
rect 196 22770 228 22802
rect 268 22770 300 22802
rect 340 22770 372 22802
rect 412 22770 444 22802
rect 484 22770 516 22802
rect 556 22770 588 22802
rect 628 22770 660 22802
rect 700 22770 732 22802
rect 772 22770 804 22802
rect 844 22770 876 22802
rect 124 22698 156 22730
rect 196 22698 228 22730
rect 268 22698 300 22730
rect 340 22698 372 22730
rect 412 22698 444 22730
rect 484 22698 516 22730
rect 556 22698 588 22730
rect 628 22698 660 22730
rect 700 22698 732 22730
rect 772 22698 804 22730
rect 844 22698 876 22730
rect 124 22626 156 22658
rect 196 22626 228 22658
rect 268 22626 300 22658
rect 340 22626 372 22658
rect 412 22626 444 22658
rect 484 22626 516 22658
rect 556 22626 588 22658
rect 628 22626 660 22658
rect 700 22626 732 22658
rect 772 22626 804 22658
rect 844 22626 876 22658
rect 124 22554 156 22586
rect 196 22554 228 22586
rect 268 22554 300 22586
rect 340 22554 372 22586
rect 412 22554 444 22586
rect 484 22554 516 22586
rect 556 22554 588 22586
rect 628 22554 660 22586
rect 700 22554 732 22586
rect 772 22554 804 22586
rect 844 22554 876 22586
rect 124 22482 156 22514
rect 196 22482 228 22514
rect 268 22482 300 22514
rect 340 22482 372 22514
rect 412 22482 444 22514
rect 484 22482 516 22514
rect 556 22482 588 22514
rect 628 22482 660 22514
rect 700 22482 732 22514
rect 772 22482 804 22514
rect 844 22482 876 22514
rect 124 22410 156 22442
rect 196 22410 228 22442
rect 268 22410 300 22442
rect 340 22410 372 22442
rect 412 22410 444 22442
rect 484 22410 516 22442
rect 556 22410 588 22442
rect 628 22410 660 22442
rect 700 22410 732 22442
rect 772 22410 804 22442
rect 844 22410 876 22442
rect 124 22338 156 22370
rect 196 22338 228 22370
rect 268 22338 300 22370
rect 340 22338 372 22370
rect 412 22338 444 22370
rect 484 22338 516 22370
rect 556 22338 588 22370
rect 628 22338 660 22370
rect 700 22338 732 22370
rect 772 22338 804 22370
rect 844 22338 876 22370
rect 124 22266 156 22298
rect 196 22266 228 22298
rect 268 22266 300 22298
rect 340 22266 372 22298
rect 412 22266 444 22298
rect 484 22266 516 22298
rect 556 22266 588 22298
rect 628 22266 660 22298
rect 700 22266 732 22298
rect 772 22266 804 22298
rect 844 22266 876 22298
rect 124 22194 156 22226
rect 196 22194 228 22226
rect 268 22194 300 22226
rect 340 22194 372 22226
rect 412 22194 444 22226
rect 484 22194 516 22226
rect 556 22194 588 22226
rect 628 22194 660 22226
rect 700 22194 732 22226
rect 772 22194 804 22226
rect 844 22194 876 22226
rect 124 22122 156 22154
rect 196 22122 228 22154
rect 268 22122 300 22154
rect 340 22122 372 22154
rect 412 22122 444 22154
rect 484 22122 516 22154
rect 556 22122 588 22154
rect 628 22122 660 22154
rect 700 22122 732 22154
rect 772 22122 804 22154
rect 844 22122 876 22154
rect 124 22050 156 22082
rect 196 22050 228 22082
rect 268 22050 300 22082
rect 340 22050 372 22082
rect 412 22050 444 22082
rect 484 22050 516 22082
rect 556 22050 588 22082
rect 628 22050 660 22082
rect 700 22050 732 22082
rect 772 22050 804 22082
rect 844 22050 876 22082
rect 124 21978 156 22010
rect 196 21978 228 22010
rect 268 21978 300 22010
rect 340 21978 372 22010
rect 412 21978 444 22010
rect 484 21978 516 22010
rect 556 21978 588 22010
rect 628 21978 660 22010
rect 700 21978 732 22010
rect 772 21978 804 22010
rect 844 21978 876 22010
rect 124 21906 156 21938
rect 196 21906 228 21938
rect 268 21906 300 21938
rect 340 21906 372 21938
rect 412 21906 444 21938
rect 484 21906 516 21938
rect 556 21906 588 21938
rect 628 21906 660 21938
rect 700 21906 732 21938
rect 772 21906 804 21938
rect 844 21906 876 21938
rect 124 21834 156 21866
rect 196 21834 228 21866
rect 268 21834 300 21866
rect 340 21834 372 21866
rect 412 21834 444 21866
rect 484 21834 516 21866
rect 556 21834 588 21866
rect 628 21834 660 21866
rect 700 21834 732 21866
rect 772 21834 804 21866
rect 844 21834 876 21866
rect 124 21762 156 21794
rect 196 21762 228 21794
rect 268 21762 300 21794
rect 340 21762 372 21794
rect 412 21762 444 21794
rect 484 21762 516 21794
rect 556 21762 588 21794
rect 628 21762 660 21794
rect 700 21762 732 21794
rect 772 21762 804 21794
rect 844 21762 876 21794
rect 124 21690 156 21722
rect 196 21690 228 21722
rect 268 21690 300 21722
rect 340 21690 372 21722
rect 412 21690 444 21722
rect 484 21690 516 21722
rect 556 21690 588 21722
rect 628 21690 660 21722
rect 700 21690 732 21722
rect 772 21690 804 21722
rect 844 21690 876 21722
rect 124 21618 156 21650
rect 196 21618 228 21650
rect 268 21618 300 21650
rect 340 21618 372 21650
rect 412 21618 444 21650
rect 484 21618 516 21650
rect 556 21618 588 21650
rect 628 21618 660 21650
rect 700 21618 732 21650
rect 772 21618 804 21650
rect 844 21618 876 21650
rect 124 21546 156 21578
rect 196 21546 228 21578
rect 268 21546 300 21578
rect 340 21546 372 21578
rect 412 21546 444 21578
rect 484 21546 516 21578
rect 556 21546 588 21578
rect 628 21546 660 21578
rect 700 21546 732 21578
rect 772 21546 804 21578
rect 844 21546 876 21578
rect 124 21474 156 21506
rect 196 21474 228 21506
rect 268 21474 300 21506
rect 340 21474 372 21506
rect 412 21474 444 21506
rect 484 21474 516 21506
rect 556 21474 588 21506
rect 628 21474 660 21506
rect 700 21474 732 21506
rect 772 21474 804 21506
rect 844 21474 876 21506
rect 124 21402 156 21434
rect 196 21402 228 21434
rect 268 21402 300 21434
rect 340 21402 372 21434
rect 412 21402 444 21434
rect 484 21402 516 21434
rect 556 21402 588 21434
rect 628 21402 660 21434
rect 700 21402 732 21434
rect 772 21402 804 21434
rect 844 21402 876 21434
rect 124 21330 156 21362
rect 196 21330 228 21362
rect 268 21330 300 21362
rect 340 21330 372 21362
rect 412 21330 444 21362
rect 484 21330 516 21362
rect 556 21330 588 21362
rect 628 21330 660 21362
rect 700 21330 732 21362
rect 772 21330 804 21362
rect 844 21330 876 21362
rect 124 21258 156 21290
rect 196 21258 228 21290
rect 268 21258 300 21290
rect 340 21258 372 21290
rect 412 21258 444 21290
rect 484 21258 516 21290
rect 556 21258 588 21290
rect 628 21258 660 21290
rect 700 21258 732 21290
rect 772 21258 804 21290
rect 844 21258 876 21290
rect 124 21186 156 21218
rect 196 21186 228 21218
rect 268 21186 300 21218
rect 340 21186 372 21218
rect 412 21186 444 21218
rect 484 21186 516 21218
rect 556 21186 588 21218
rect 628 21186 660 21218
rect 700 21186 732 21218
rect 772 21186 804 21218
rect 844 21186 876 21218
rect 124 21114 156 21146
rect 196 21114 228 21146
rect 268 21114 300 21146
rect 340 21114 372 21146
rect 412 21114 444 21146
rect 484 21114 516 21146
rect 556 21114 588 21146
rect 628 21114 660 21146
rect 700 21114 732 21146
rect 772 21114 804 21146
rect 844 21114 876 21146
rect 124 21042 156 21074
rect 196 21042 228 21074
rect 268 21042 300 21074
rect 340 21042 372 21074
rect 412 21042 444 21074
rect 484 21042 516 21074
rect 556 21042 588 21074
rect 628 21042 660 21074
rect 700 21042 732 21074
rect 772 21042 804 21074
rect 844 21042 876 21074
rect 124 20970 156 21002
rect 196 20970 228 21002
rect 268 20970 300 21002
rect 340 20970 372 21002
rect 412 20970 444 21002
rect 484 20970 516 21002
rect 556 20970 588 21002
rect 628 20970 660 21002
rect 700 20970 732 21002
rect 772 20970 804 21002
rect 844 20970 876 21002
rect 124 20898 156 20930
rect 196 20898 228 20930
rect 268 20898 300 20930
rect 340 20898 372 20930
rect 412 20898 444 20930
rect 484 20898 516 20930
rect 556 20898 588 20930
rect 628 20898 660 20930
rect 700 20898 732 20930
rect 772 20898 804 20930
rect 844 20898 876 20930
rect 124 20826 156 20858
rect 196 20826 228 20858
rect 268 20826 300 20858
rect 340 20826 372 20858
rect 412 20826 444 20858
rect 484 20826 516 20858
rect 556 20826 588 20858
rect 628 20826 660 20858
rect 700 20826 732 20858
rect 772 20826 804 20858
rect 844 20826 876 20858
rect 124 20754 156 20786
rect 196 20754 228 20786
rect 268 20754 300 20786
rect 340 20754 372 20786
rect 412 20754 444 20786
rect 484 20754 516 20786
rect 556 20754 588 20786
rect 628 20754 660 20786
rect 700 20754 732 20786
rect 772 20754 804 20786
rect 844 20754 876 20786
rect 124 20682 156 20714
rect 196 20682 228 20714
rect 268 20682 300 20714
rect 340 20682 372 20714
rect 412 20682 444 20714
rect 484 20682 516 20714
rect 556 20682 588 20714
rect 628 20682 660 20714
rect 700 20682 732 20714
rect 772 20682 804 20714
rect 844 20682 876 20714
rect 124 20610 156 20642
rect 196 20610 228 20642
rect 268 20610 300 20642
rect 340 20610 372 20642
rect 412 20610 444 20642
rect 484 20610 516 20642
rect 556 20610 588 20642
rect 628 20610 660 20642
rect 700 20610 732 20642
rect 772 20610 804 20642
rect 844 20610 876 20642
rect 124 20538 156 20570
rect 196 20538 228 20570
rect 268 20538 300 20570
rect 340 20538 372 20570
rect 412 20538 444 20570
rect 484 20538 516 20570
rect 556 20538 588 20570
rect 628 20538 660 20570
rect 700 20538 732 20570
rect 772 20538 804 20570
rect 844 20538 876 20570
rect 124 20466 156 20498
rect 196 20466 228 20498
rect 268 20466 300 20498
rect 340 20466 372 20498
rect 412 20466 444 20498
rect 484 20466 516 20498
rect 556 20466 588 20498
rect 628 20466 660 20498
rect 700 20466 732 20498
rect 772 20466 804 20498
rect 844 20466 876 20498
rect 124 20394 156 20426
rect 196 20394 228 20426
rect 268 20394 300 20426
rect 340 20394 372 20426
rect 412 20394 444 20426
rect 484 20394 516 20426
rect 556 20394 588 20426
rect 628 20394 660 20426
rect 700 20394 732 20426
rect 772 20394 804 20426
rect 844 20394 876 20426
rect 124 20322 156 20354
rect 196 20322 228 20354
rect 268 20322 300 20354
rect 340 20322 372 20354
rect 412 20322 444 20354
rect 484 20322 516 20354
rect 556 20322 588 20354
rect 628 20322 660 20354
rect 700 20322 732 20354
rect 772 20322 804 20354
rect 844 20322 876 20354
rect 124 20250 156 20282
rect 196 20250 228 20282
rect 268 20250 300 20282
rect 340 20250 372 20282
rect 412 20250 444 20282
rect 484 20250 516 20282
rect 556 20250 588 20282
rect 628 20250 660 20282
rect 700 20250 732 20282
rect 772 20250 804 20282
rect 844 20250 876 20282
rect 124 20178 156 20210
rect 196 20178 228 20210
rect 268 20178 300 20210
rect 340 20178 372 20210
rect 412 20178 444 20210
rect 484 20178 516 20210
rect 556 20178 588 20210
rect 628 20178 660 20210
rect 700 20178 732 20210
rect 772 20178 804 20210
rect 844 20178 876 20210
rect 124 20106 156 20138
rect 196 20106 228 20138
rect 268 20106 300 20138
rect 340 20106 372 20138
rect 412 20106 444 20138
rect 484 20106 516 20138
rect 556 20106 588 20138
rect 628 20106 660 20138
rect 700 20106 732 20138
rect 772 20106 804 20138
rect 844 20106 876 20138
rect 124 20034 156 20066
rect 196 20034 228 20066
rect 268 20034 300 20066
rect 340 20034 372 20066
rect 412 20034 444 20066
rect 484 20034 516 20066
rect 556 20034 588 20066
rect 628 20034 660 20066
rect 700 20034 732 20066
rect 772 20034 804 20066
rect 844 20034 876 20066
rect 124 19962 156 19994
rect 196 19962 228 19994
rect 268 19962 300 19994
rect 340 19962 372 19994
rect 412 19962 444 19994
rect 484 19962 516 19994
rect 556 19962 588 19994
rect 628 19962 660 19994
rect 700 19962 732 19994
rect 772 19962 804 19994
rect 844 19962 876 19994
rect 124 19890 156 19922
rect 196 19890 228 19922
rect 268 19890 300 19922
rect 340 19890 372 19922
rect 412 19890 444 19922
rect 484 19890 516 19922
rect 556 19890 588 19922
rect 628 19890 660 19922
rect 700 19890 732 19922
rect 772 19890 804 19922
rect 844 19890 876 19922
rect 124 19818 156 19850
rect 196 19818 228 19850
rect 268 19818 300 19850
rect 340 19818 372 19850
rect 412 19818 444 19850
rect 484 19818 516 19850
rect 556 19818 588 19850
rect 628 19818 660 19850
rect 700 19818 732 19850
rect 772 19818 804 19850
rect 844 19818 876 19850
rect 124 19746 156 19778
rect 196 19746 228 19778
rect 268 19746 300 19778
rect 340 19746 372 19778
rect 412 19746 444 19778
rect 484 19746 516 19778
rect 556 19746 588 19778
rect 628 19746 660 19778
rect 700 19746 732 19778
rect 772 19746 804 19778
rect 844 19746 876 19778
rect 124 19674 156 19706
rect 196 19674 228 19706
rect 268 19674 300 19706
rect 340 19674 372 19706
rect 412 19674 444 19706
rect 484 19674 516 19706
rect 556 19674 588 19706
rect 628 19674 660 19706
rect 700 19674 732 19706
rect 772 19674 804 19706
rect 844 19674 876 19706
rect 124 19602 156 19634
rect 196 19602 228 19634
rect 268 19602 300 19634
rect 340 19602 372 19634
rect 412 19602 444 19634
rect 484 19602 516 19634
rect 556 19602 588 19634
rect 628 19602 660 19634
rect 700 19602 732 19634
rect 772 19602 804 19634
rect 844 19602 876 19634
rect 124 19530 156 19562
rect 196 19530 228 19562
rect 268 19530 300 19562
rect 340 19530 372 19562
rect 412 19530 444 19562
rect 484 19530 516 19562
rect 556 19530 588 19562
rect 628 19530 660 19562
rect 700 19530 732 19562
rect 772 19530 804 19562
rect 844 19530 876 19562
rect 124 19458 156 19490
rect 196 19458 228 19490
rect 268 19458 300 19490
rect 340 19458 372 19490
rect 412 19458 444 19490
rect 484 19458 516 19490
rect 556 19458 588 19490
rect 628 19458 660 19490
rect 700 19458 732 19490
rect 772 19458 804 19490
rect 844 19458 876 19490
rect 124 19386 156 19418
rect 196 19386 228 19418
rect 268 19386 300 19418
rect 340 19386 372 19418
rect 412 19386 444 19418
rect 484 19386 516 19418
rect 556 19386 588 19418
rect 628 19386 660 19418
rect 700 19386 732 19418
rect 772 19386 804 19418
rect 844 19386 876 19418
rect 124 19314 156 19346
rect 196 19314 228 19346
rect 268 19314 300 19346
rect 340 19314 372 19346
rect 412 19314 444 19346
rect 484 19314 516 19346
rect 556 19314 588 19346
rect 628 19314 660 19346
rect 700 19314 732 19346
rect 772 19314 804 19346
rect 844 19314 876 19346
rect 124 19242 156 19274
rect 196 19242 228 19274
rect 268 19242 300 19274
rect 340 19242 372 19274
rect 412 19242 444 19274
rect 484 19242 516 19274
rect 556 19242 588 19274
rect 628 19242 660 19274
rect 700 19242 732 19274
rect 772 19242 804 19274
rect 844 19242 876 19274
rect 124 19170 156 19202
rect 196 19170 228 19202
rect 268 19170 300 19202
rect 340 19170 372 19202
rect 412 19170 444 19202
rect 484 19170 516 19202
rect 556 19170 588 19202
rect 628 19170 660 19202
rect 700 19170 732 19202
rect 772 19170 804 19202
rect 844 19170 876 19202
rect 124 19098 156 19130
rect 196 19098 228 19130
rect 268 19098 300 19130
rect 340 19098 372 19130
rect 412 19098 444 19130
rect 484 19098 516 19130
rect 556 19098 588 19130
rect 628 19098 660 19130
rect 700 19098 732 19130
rect 772 19098 804 19130
rect 844 19098 876 19130
rect 124 19026 156 19058
rect 196 19026 228 19058
rect 268 19026 300 19058
rect 340 19026 372 19058
rect 412 19026 444 19058
rect 484 19026 516 19058
rect 556 19026 588 19058
rect 628 19026 660 19058
rect 700 19026 732 19058
rect 772 19026 804 19058
rect 844 19026 876 19058
rect 124 18954 156 18986
rect 196 18954 228 18986
rect 268 18954 300 18986
rect 340 18954 372 18986
rect 412 18954 444 18986
rect 484 18954 516 18986
rect 556 18954 588 18986
rect 628 18954 660 18986
rect 700 18954 732 18986
rect 772 18954 804 18986
rect 844 18954 876 18986
rect 124 18882 156 18914
rect 196 18882 228 18914
rect 268 18882 300 18914
rect 340 18882 372 18914
rect 412 18882 444 18914
rect 484 18882 516 18914
rect 556 18882 588 18914
rect 628 18882 660 18914
rect 700 18882 732 18914
rect 772 18882 804 18914
rect 844 18882 876 18914
rect 124 18810 156 18842
rect 196 18810 228 18842
rect 268 18810 300 18842
rect 340 18810 372 18842
rect 412 18810 444 18842
rect 484 18810 516 18842
rect 556 18810 588 18842
rect 628 18810 660 18842
rect 700 18810 732 18842
rect 772 18810 804 18842
rect 844 18810 876 18842
rect 124 18738 156 18770
rect 196 18738 228 18770
rect 268 18738 300 18770
rect 340 18738 372 18770
rect 412 18738 444 18770
rect 484 18738 516 18770
rect 556 18738 588 18770
rect 628 18738 660 18770
rect 700 18738 732 18770
rect 772 18738 804 18770
rect 844 18738 876 18770
rect 124 18666 156 18698
rect 196 18666 228 18698
rect 268 18666 300 18698
rect 340 18666 372 18698
rect 412 18666 444 18698
rect 484 18666 516 18698
rect 556 18666 588 18698
rect 628 18666 660 18698
rect 700 18666 732 18698
rect 772 18666 804 18698
rect 844 18666 876 18698
rect 124 18594 156 18626
rect 196 18594 228 18626
rect 268 18594 300 18626
rect 340 18594 372 18626
rect 412 18594 444 18626
rect 484 18594 516 18626
rect 556 18594 588 18626
rect 628 18594 660 18626
rect 700 18594 732 18626
rect 772 18594 804 18626
rect 844 18594 876 18626
rect 124 18522 156 18554
rect 196 18522 228 18554
rect 268 18522 300 18554
rect 340 18522 372 18554
rect 412 18522 444 18554
rect 484 18522 516 18554
rect 556 18522 588 18554
rect 628 18522 660 18554
rect 700 18522 732 18554
rect 772 18522 804 18554
rect 844 18522 876 18554
rect 124 18450 156 18482
rect 196 18450 228 18482
rect 268 18450 300 18482
rect 340 18450 372 18482
rect 412 18450 444 18482
rect 484 18450 516 18482
rect 556 18450 588 18482
rect 628 18450 660 18482
rect 700 18450 732 18482
rect 772 18450 804 18482
rect 844 18450 876 18482
rect 124 18378 156 18410
rect 196 18378 228 18410
rect 268 18378 300 18410
rect 340 18378 372 18410
rect 412 18378 444 18410
rect 484 18378 516 18410
rect 556 18378 588 18410
rect 628 18378 660 18410
rect 700 18378 732 18410
rect 772 18378 804 18410
rect 844 18378 876 18410
rect 124 18306 156 18338
rect 196 18306 228 18338
rect 268 18306 300 18338
rect 340 18306 372 18338
rect 412 18306 444 18338
rect 484 18306 516 18338
rect 556 18306 588 18338
rect 628 18306 660 18338
rect 700 18306 732 18338
rect 772 18306 804 18338
rect 844 18306 876 18338
rect 124 18234 156 18266
rect 196 18234 228 18266
rect 268 18234 300 18266
rect 340 18234 372 18266
rect 412 18234 444 18266
rect 484 18234 516 18266
rect 556 18234 588 18266
rect 628 18234 660 18266
rect 700 18234 732 18266
rect 772 18234 804 18266
rect 844 18234 876 18266
rect 124 18162 156 18194
rect 196 18162 228 18194
rect 268 18162 300 18194
rect 340 18162 372 18194
rect 412 18162 444 18194
rect 484 18162 516 18194
rect 556 18162 588 18194
rect 628 18162 660 18194
rect 700 18162 732 18194
rect 772 18162 804 18194
rect 844 18162 876 18194
rect 196 17816 228 17848
rect 268 17816 300 17848
rect 340 17816 372 17848
rect 412 17816 444 17848
rect 484 17816 516 17848
rect 556 17816 588 17848
rect 628 17816 660 17848
rect 700 17816 732 17848
rect 772 17816 804 17848
rect 844 17816 876 17848
rect 124 17744 156 17776
rect 196 17744 228 17776
rect 268 17744 300 17776
rect 340 17744 372 17776
rect 412 17744 444 17776
rect 484 17744 516 17776
rect 556 17744 588 17776
rect 628 17744 660 17776
rect 700 17744 732 17776
rect 772 17744 804 17776
rect 844 17744 876 17776
rect 124 17672 156 17704
rect 196 17672 228 17704
rect 268 17672 300 17704
rect 340 17672 372 17704
rect 412 17672 444 17704
rect 484 17672 516 17704
rect 556 17672 588 17704
rect 628 17672 660 17704
rect 700 17672 732 17704
rect 772 17672 804 17704
rect 844 17672 876 17704
rect 124 17600 156 17632
rect 196 17600 228 17632
rect 268 17600 300 17632
rect 340 17600 372 17632
rect 412 17600 444 17632
rect 484 17600 516 17632
rect 556 17600 588 17632
rect 628 17600 660 17632
rect 700 17600 732 17632
rect 772 17600 804 17632
rect 844 17600 876 17632
rect 124 17528 156 17560
rect 196 17528 228 17560
rect 268 17528 300 17560
rect 340 17528 372 17560
rect 412 17528 444 17560
rect 484 17528 516 17560
rect 556 17528 588 17560
rect 628 17528 660 17560
rect 700 17528 732 17560
rect 772 17528 804 17560
rect 844 17528 876 17560
rect 124 17456 156 17488
rect 196 17456 228 17488
rect 268 17456 300 17488
rect 340 17456 372 17488
rect 412 17456 444 17488
rect 484 17456 516 17488
rect 556 17456 588 17488
rect 628 17456 660 17488
rect 700 17456 732 17488
rect 772 17456 804 17488
rect 844 17456 876 17488
rect 124 17384 156 17416
rect 196 17384 228 17416
rect 268 17384 300 17416
rect 340 17384 372 17416
rect 412 17384 444 17416
rect 484 17384 516 17416
rect 556 17384 588 17416
rect 628 17384 660 17416
rect 700 17384 732 17416
rect 772 17384 804 17416
rect 844 17384 876 17416
rect 124 17312 156 17344
rect 196 17312 228 17344
rect 268 17312 300 17344
rect 340 17312 372 17344
rect 412 17312 444 17344
rect 484 17312 516 17344
rect 556 17312 588 17344
rect 628 17312 660 17344
rect 700 17312 732 17344
rect 772 17312 804 17344
rect 844 17312 876 17344
rect 124 17240 156 17272
rect 196 17240 228 17272
rect 268 17240 300 17272
rect 340 17240 372 17272
rect 412 17240 444 17272
rect 484 17240 516 17272
rect 556 17240 588 17272
rect 628 17240 660 17272
rect 700 17240 732 17272
rect 772 17240 804 17272
rect 844 17240 876 17272
rect 124 17168 156 17200
rect 196 17168 228 17200
rect 268 17168 300 17200
rect 340 17168 372 17200
rect 412 17168 444 17200
rect 484 17168 516 17200
rect 556 17168 588 17200
rect 628 17168 660 17200
rect 700 17168 732 17200
rect 772 17168 804 17200
rect 844 17168 876 17200
rect 124 17096 156 17128
rect 196 17096 228 17128
rect 268 17096 300 17128
rect 340 17096 372 17128
rect 412 17096 444 17128
rect 484 17096 516 17128
rect 556 17096 588 17128
rect 628 17096 660 17128
rect 700 17096 732 17128
rect 772 17096 804 17128
rect 844 17096 876 17128
rect 124 17024 156 17056
rect 196 17024 228 17056
rect 268 17024 300 17056
rect 340 17024 372 17056
rect 412 17024 444 17056
rect 484 17024 516 17056
rect 556 17024 588 17056
rect 628 17024 660 17056
rect 700 17024 732 17056
rect 772 17024 804 17056
rect 844 17024 876 17056
rect 124 16952 156 16984
rect 196 16952 228 16984
rect 268 16952 300 16984
rect 340 16952 372 16984
rect 412 16952 444 16984
rect 484 16952 516 16984
rect 556 16952 588 16984
rect 628 16952 660 16984
rect 700 16952 732 16984
rect 772 16952 804 16984
rect 844 16952 876 16984
rect 124 16880 156 16912
rect 196 16880 228 16912
rect 268 16880 300 16912
rect 340 16880 372 16912
rect 412 16880 444 16912
rect 484 16880 516 16912
rect 556 16880 588 16912
rect 628 16880 660 16912
rect 700 16880 732 16912
rect 772 16880 804 16912
rect 844 16880 876 16912
rect 124 16808 156 16840
rect 196 16808 228 16840
rect 268 16808 300 16840
rect 340 16808 372 16840
rect 412 16808 444 16840
rect 484 16808 516 16840
rect 556 16808 588 16840
rect 628 16808 660 16840
rect 700 16808 732 16840
rect 772 16808 804 16840
rect 844 16808 876 16840
rect 124 16736 156 16768
rect 196 16736 228 16768
rect 268 16736 300 16768
rect 340 16736 372 16768
rect 412 16736 444 16768
rect 484 16736 516 16768
rect 556 16736 588 16768
rect 628 16736 660 16768
rect 700 16736 732 16768
rect 772 16736 804 16768
rect 844 16736 876 16768
rect 124 16664 156 16696
rect 196 16664 228 16696
rect 268 16664 300 16696
rect 340 16664 372 16696
rect 412 16664 444 16696
rect 484 16664 516 16696
rect 556 16664 588 16696
rect 628 16664 660 16696
rect 700 16664 732 16696
rect 772 16664 804 16696
rect 844 16664 876 16696
rect 124 16592 156 16624
rect 196 16592 228 16624
rect 268 16592 300 16624
rect 340 16592 372 16624
rect 412 16592 444 16624
rect 484 16592 516 16624
rect 556 16592 588 16624
rect 628 16592 660 16624
rect 700 16592 732 16624
rect 772 16592 804 16624
rect 844 16592 876 16624
rect 124 16520 156 16552
rect 196 16520 228 16552
rect 268 16520 300 16552
rect 340 16520 372 16552
rect 412 16520 444 16552
rect 484 16520 516 16552
rect 556 16520 588 16552
rect 628 16520 660 16552
rect 700 16520 732 16552
rect 772 16520 804 16552
rect 844 16520 876 16552
rect 124 16448 156 16480
rect 196 16448 228 16480
rect 268 16448 300 16480
rect 340 16448 372 16480
rect 412 16448 444 16480
rect 484 16448 516 16480
rect 556 16448 588 16480
rect 628 16448 660 16480
rect 700 16448 732 16480
rect 772 16448 804 16480
rect 844 16448 876 16480
rect 124 16376 156 16408
rect 196 16376 228 16408
rect 268 16376 300 16408
rect 340 16376 372 16408
rect 412 16376 444 16408
rect 484 16376 516 16408
rect 556 16376 588 16408
rect 628 16376 660 16408
rect 700 16376 732 16408
rect 772 16376 804 16408
rect 844 16376 876 16408
rect 124 16304 156 16336
rect 196 16304 228 16336
rect 268 16304 300 16336
rect 340 16304 372 16336
rect 412 16304 444 16336
rect 484 16304 516 16336
rect 556 16304 588 16336
rect 628 16304 660 16336
rect 700 16304 732 16336
rect 772 16304 804 16336
rect 844 16304 876 16336
rect 124 16232 156 16264
rect 196 16232 228 16264
rect 268 16232 300 16264
rect 340 16232 372 16264
rect 412 16232 444 16264
rect 484 16232 516 16264
rect 556 16232 588 16264
rect 628 16232 660 16264
rect 700 16232 732 16264
rect 772 16232 804 16264
rect 844 16232 876 16264
rect 124 16160 156 16192
rect 196 16160 228 16192
rect 268 16160 300 16192
rect 340 16160 372 16192
rect 412 16160 444 16192
rect 484 16160 516 16192
rect 556 16160 588 16192
rect 628 16160 660 16192
rect 700 16160 732 16192
rect 772 16160 804 16192
rect 844 16160 876 16192
rect 124 16088 156 16120
rect 196 16088 228 16120
rect 268 16088 300 16120
rect 340 16088 372 16120
rect 412 16088 444 16120
rect 484 16088 516 16120
rect 556 16088 588 16120
rect 628 16088 660 16120
rect 700 16088 732 16120
rect 772 16088 804 16120
rect 844 16088 876 16120
rect 124 16016 156 16048
rect 196 16016 228 16048
rect 268 16016 300 16048
rect 340 16016 372 16048
rect 412 16016 444 16048
rect 484 16016 516 16048
rect 556 16016 588 16048
rect 628 16016 660 16048
rect 700 16016 732 16048
rect 772 16016 804 16048
rect 844 16016 876 16048
rect 124 15944 156 15976
rect 196 15944 228 15976
rect 268 15944 300 15976
rect 340 15944 372 15976
rect 412 15944 444 15976
rect 484 15944 516 15976
rect 556 15944 588 15976
rect 628 15944 660 15976
rect 700 15944 732 15976
rect 772 15944 804 15976
rect 844 15944 876 15976
rect 124 15872 156 15904
rect 196 15872 228 15904
rect 268 15872 300 15904
rect 340 15872 372 15904
rect 412 15872 444 15904
rect 484 15872 516 15904
rect 556 15872 588 15904
rect 628 15872 660 15904
rect 700 15872 732 15904
rect 772 15872 804 15904
rect 844 15872 876 15904
rect 124 15800 156 15832
rect 196 15800 228 15832
rect 268 15800 300 15832
rect 340 15800 372 15832
rect 412 15800 444 15832
rect 484 15800 516 15832
rect 556 15800 588 15832
rect 628 15800 660 15832
rect 700 15800 732 15832
rect 772 15800 804 15832
rect 844 15800 876 15832
rect 124 15728 156 15760
rect 196 15728 228 15760
rect 268 15728 300 15760
rect 340 15728 372 15760
rect 412 15728 444 15760
rect 484 15728 516 15760
rect 556 15728 588 15760
rect 628 15728 660 15760
rect 700 15728 732 15760
rect 772 15728 804 15760
rect 844 15728 876 15760
rect 124 15656 156 15688
rect 196 15656 228 15688
rect 268 15656 300 15688
rect 340 15656 372 15688
rect 412 15656 444 15688
rect 484 15656 516 15688
rect 556 15656 588 15688
rect 628 15656 660 15688
rect 700 15656 732 15688
rect 772 15656 804 15688
rect 844 15656 876 15688
rect 124 15584 156 15616
rect 196 15584 228 15616
rect 268 15584 300 15616
rect 340 15584 372 15616
rect 412 15584 444 15616
rect 484 15584 516 15616
rect 556 15584 588 15616
rect 628 15584 660 15616
rect 700 15584 732 15616
rect 772 15584 804 15616
rect 844 15584 876 15616
rect 124 15512 156 15544
rect 196 15512 228 15544
rect 268 15512 300 15544
rect 340 15512 372 15544
rect 412 15512 444 15544
rect 484 15512 516 15544
rect 556 15512 588 15544
rect 628 15512 660 15544
rect 700 15512 732 15544
rect 772 15512 804 15544
rect 844 15512 876 15544
rect 124 15440 156 15472
rect 196 15440 228 15472
rect 268 15440 300 15472
rect 340 15440 372 15472
rect 412 15440 444 15472
rect 484 15440 516 15472
rect 556 15440 588 15472
rect 628 15440 660 15472
rect 700 15440 732 15472
rect 772 15440 804 15472
rect 844 15440 876 15472
rect 124 15368 156 15400
rect 196 15368 228 15400
rect 268 15368 300 15400
rect 340 15368 372 15400
rect 412 15368 444 15400
rect 484 15368 516 15400
rect 556 15368 588 15400
rect 628 15368 660 15400
rect 700 15368 732 15400
rect 772 15368 804 15400
rect 844 15368 876 15400
rect 124 15296 156 15328
rect 196 15296 228 15328
rect 268 15296 300 15328
rect 340 15296 372 15328
rect 412 15296 444 15328
rect 484 15296 516 15328
rect 556 15296 588 15328
rect 628 15296 660 15328
rect 700 15296 732 15328
rect 772 15296 804 15328
rect 844 15296 876 15328
rect 124 15224 156 15256
rect 196 15224 228 15256
rect 268 15224 300 15256
rect 340 15224 372 15256
rect 412 15224 444 15256
rect 484 15224 516 15256
rect 556 15224 588 15256
rect 628 15224 660 15256
rect 700 15224 732 15256
rect 772 15224 804 15256
rect 844 15224 876 15256
rect 124 15152 156 15184
rect 196 15152 228 15184
rect 268 15152 300 15184
rect 340 15152 372 15184
rect 412 15152 444 15184
rect 484 15152 516 15184
rect 556 15152 588 15184
rect 628 15152 660 15184
rect 700 15152 732 15184
rect 772 15152 804 15184
rect 844 15152 876 15184
rect 124 15080 156 15112
rect 196 15080 228 15112
rect 268 15080 300 15112
rect 340 15080 372 15112
rect 412 15080 444 15112
rect 484 15080 516 15112
rect 556 15080 588 15112
rect 628 15080 660 15112
rect 700 15080 732 15112
rect 772 15080 804 15112
rect 844 15080 876 15112
rect 124 15008 156 15040
rect 196 15008 228 15040
rect 268 15008 300 15040
rect 340 15008 372 15040
rect 412 15008 444 15040
rect 484 15008 516 15040
rect 556 15008 588 15040
rect 628 15008 660 15040
rect 700 15008 732 15040
rect 772 15008 804 15040
rect 844 15008 876 15040
rect 124 14936 156 14968
rect 196 14936 228 14968
rect 268 14936 300 14968
rect 340 14936 372 14968
rect 412 14936 444 14968
rect 484 14936 516 14968
rect 556 14936 588 14968
rect 628 14936 660 14968
rect 700 14936 732 14968
rect 772 14936 804 14968
rect 844 14936 876 14968
rect 124 14864 156 14896
rect 196 14864 228 14896
rect 268 14864 300 14896
rect 340 14864 372 14896
rect 412 14864 444 14896
rect 484 14864 516 14896
rect 556 14864 588 14896
rect 628 14864 660 14896
rect 700 14864 732 14896
rect 772 14864 804 14896
rect 844 14864 876 14896
rect 124 14792 156 14824
rect 196 14792 228 14824
rect 268 14792 300 14824
rect 340 14792 372 14824
rect 412 14792 444 14824
rect 484 14792 516 14824
rect 556 14792 588 14824
rect 628 14792 660 14824
rect 700 14792 732 14824
rect 772 14792 804 14824
rect 844 14792 876 14824
rect 124 14720 156 14752
rect 196 14720 228 14752
rect 268 14720 300 14752
rect 340 14720 372 14752
rect 412 14720 444 14752
rect 484 14720 516 14752
rect 556 14720 588 14752
rect 628 14720 660 14752
rect 700 14720 732 14752
rect 772 14720 804 14752
rect 844 14720 876 14752
rect 124 14648 156 14680
rect 196 14648 228 14680
rect 268 14648 300 14680
rect 340 14648 372 14680
rect 412 14648 444 14680
rect 484 14648 516 14680
rect 556 14648 588 14680
rect 628 14648 660 14680
rect 700 14648 732 14680
rect 772 14648 804 14680
rect 844 14648 876 14680
rect 124 14576 156 14608
rect 196 14576 228 14608
rect 268 14576 300 14608
rect 340 14576 372 14608
rect 412 14576 444 14608
rect 484 14576 516 14608
rect 556 14576 588 14608
rect 628 14576 660 14608
rect 700 14576 732 14608
rect 772 14576 804 14608
rect 844 14576 876 14608
rect 124 14504 156 14536
rect 196 14504 228 14536
rect 268 14504 300 14536
rect 340 14504 372 14536
rect 412 14504 444 14536
rect 484 14504 516 14536
rect 556 14504 588 14536
rect 628 14504 660 14536
rect 700 14504 732 14536
rect 772 14504 804 14536
rect 844 14504 876 14536
rect 124 14432 156 14464
rect 196 14432 228 14464
rect 268 14432 300 14464
rect 340 14432 372 14464
rect 412 14432 444 14464
rect 484 14432 516 14464
rect 556 14432 588 14464
rect 628 14432 660 14464
rect 700 14432 732 14464
rect 772 14432 804 14464
rect 844 14432 876 14464
rect 124 14360 156 14392
rect 196 14360 228 14392
rect 268 14360 300 14392
rect 340 14360 372 14392
rect 412 14360 444 14392
rect 484 14360 516 14392
rect 556 14360 588 14392
rect 628 14360 660 14392
rect 700 14360 732 14392
rect 772 14360 804 14392
rect 844 14360 876 14392
rect 124 14288 156 14320
rect 196 14288 228 14320
rect 268 14288 300 14320
rect 340 14288 372 14320
rect 412 14288 444 14320
rect 484 14288 516 14320
rect 556 14288 588 14320
rect 628 14288 660 14320
rect 700 14288 732 14320
rect 772 14288 804 14320
rect 844 14288 876 14320
rect 124 14216 156 14248
rect 196 14216 228 14248
rect 268 14216 300 14248
rect 340 14216 372 14248
rect 412 14216 444 14248
rect 484 14216 516 14248
rect 556 14216 588 14248
rect 628 14216 660 14248
rect 700 14216 732 14248
rect 772 14216 804 14248
rect 844 14216 876 14248
rect 124 14144 156 14176
rect 196 14144 228 14176
rect 268 14144 300 14176
rect 340 14144 372 14176
rect 412 14144 444 14176
rect 484 14144 516 14176
rect 556 14144 588 14176
rect 628 14144 660 14176
rect 700 14144 732 14176
rect 772 14144 804 14176
rect 844 14144 876 14176
rect 124 14072 156 14104
rect 196 14072 228 14104
rect 268 14072 300 14104
rect 340 14072 372 14104
rect 412 14072 444 14104
rect 484 14072 516 14104
rect 556 14072 588 14104
rect 628 14072 660 14104
rect 700 14072 732 14104
rect 772 14072 804 14104
rect 844 14072 876 14104
rect 124 14000 156 14032
rect 196 14000 228 14032
rect 268 14000 300 14032
rect 340 14000 372 14032
rect 412 14000 444 14032
rect 484 14000 516 14032
rect 556 14000 588 14032
rect 628 14000 660 14032
rect 700 14000 732 14032
rect 772 14000 804 14032
rect 844 14000 876 14032
rect 124 13928 156 13960
rect 196 13928 228 13960
rect 268 13928 300 13960
rect 340 13928 372 13960
rect 412 13928 444 13960
rect 484 13928 516 13960
rect 556 13928 588 13960
rect 628 13928 660 13960
rect 700 13928 732 13960
rect 772 13928 804 13960
rect 844 13928 876 13960
rect 124 13856 156 13888
rect 196 13856 228 13888
rect 268 13856 300 13888
rect 340 13856 372 13888
rect 412 13856 444 13888
rect 484 13856 516 13888
rect 556 13856 588 13888
rect 628 13856 660 13888
rect 700 13856 732 13888
rect 772 13856 804 13888
rect 844 13856 876 13888
rect 124 13784 156 13816
rect 196 13784 228 13816
rect 268 13784 300 13816
rect 340 13784 372 13816
rect 412 13784 444 13816
rect 484 13784 516 13816
rect 556 13784 588 13816
rect 628 13784 660 13816
rect 700 13784 732 13816
rect 772 13784 804 13816
rect 844 13784 876 13816
rect 124 13712 156 13744
rect 196 13712 228 13744
rect 268 13712 300 13744
rect 340 13712 372 13744
rect 412 13712 444 13744
rect 484 13712 516 13744
rect 556 13712 588 13744
rect 628 13712 660 13744
rect 700 13712 732 13744
rect 772 13712 804 13744
rect 844 13712 876 13744
rect 124 13640 156 13672
rect 196 13640 228 13672
rect 268 13640 300 13672
rect 340 13640 372 13672
rect 412 13640 444 13672
rect 484 13640 516 13672
rect 556 13640 588 13672
rect 628 13640 660 13672
rect 700 13640 732 13672
rect 772 13640 804 13672
rect 844 13640 876 13672
rect 124 13568 156 13600
rect 196 13568 228 13600
rect 268 13568 300 13600
rect 340 13568 372 13600
rect 412 13568 444 13600
rect 484 13568 516 13600
rect 556 13568 588 13600
rect 628 13568 660 13600
rect 700 13568 732 13600
rect 772 13568 804 13600
rect 844 13568 876 13600
rect 124 13496 156 13528
rect 196 13496 228 13528
rect 268 13496 300 13528
rect 340 13496 372 13528
rect 412 13496 444 13528
rect 484 13496 516 13528
rect 556 13496 588 13528
rect 628 13496 660 13528
rect 700 13496 732 13528
rect 772 13496 804 13528
rect 844 13496 876 13528
rect 124 13424 156 13456
rect 196 13424 228 13456
rect 268 13424 300 13456
rect 340 13424 372 13456
rect 412 13424 444 13456
rect 484 13424 516 13456
rect 556 13424 588 13456
rect 628 13424 660 13456
rect 700 13424 732 13456
rect 772 13424 804 13456
rect 844 13424 876 13456
rect 124 13352 156 13384
rect 196 13352 228 13384
rect 268 13352 300 13384
rect 340 13352 372 13384
rect 412 13352 444 13384
rect 484 13352 516 13384
rect 556 13352 588 13384
rect 628 13352 660 13384
rect 700 13352 732 13384
rect 772 13352 804 13384
rect 844 13352 876 13384
rect 124 13280 156 13312
rect 196 13280 228 13312
rect 268 13280 300 13312
rect 340 13280 372 13312
rect 412 13280 444 13312
rect 484 13280 516 13312
rect 556 13280 588 13312
rect 628 13280 660 13312
rect 700 13280 732 13312
rect 772 13280 804 13312
rect 844 13280 876 13312
rect 124 13208 156 13240
rect 196 13208 228 13240
rect 268 13208 300 13240
rect 340 13208 372 13240
rect 412 13208 444 13240
rect 484 13208 516 13240
rect 556 13208 588 13240
rect 628 13208 660 13240
rect 700 13208 732 13240
rect 772 13208 804 13240
rect 844 13208 876 13240
rect 124 13136 156 13168
rect 196 13136 228 13168
rect 268 13136 300 13168
rect 340 13136 372 13168
rect 412 13136 444 13168
rect 484 13136 516 13168
rect 556 13136 588 13168
rect 628 13136 660 13168
rect 700 13136 732 13168
rect 772 13136 804 13168
rect 844 13136 876 13168
rect 124 13064 156 13096
rect 196 13064 228 13096
rect 268 13064 300 13096
rect 340 13064 372 13096
rect 412 13064 444 13096
rect 484 13064 516 13096
rect 556 13064 588 13096
rect 628 13064 660 13096
rect 700 13064 732 13096
rect 772 13064 804 13096
rect 844 13064 876 13096
rect 44 31416 956 31430
rect 44 31384 223 31416
rect 255 31384 292 31416
rect 324 31384 362 31416
rect 394 31384 431 31416
rect 463 31384 502 31416
rect 534 31384 572 31416
rect 604 31384 640 31416
rect 672 31384 710 31416
rect 742 31384 956 31416
rect 44 31370 956 31384
rect 50 27971 950 28034
rect 50 27939 124 27971
rect 156 27939 196 27971
rect 228 27939 268 27971
rect 300 27939 340 27971
rect 372 27939 412 27971
rect 444 27939 484 27971
rect 516 27939 556 27971
rect 588 27939 628 27971
rect 660 27939 700 27971
rect 732 27939 772 27971
rect 804 27939 844 27971
rect 876 27939 950 27971
rect 50 27899 950 27939
rect 50 27867 124 27899
rect 156 27867 196 27899
rect 228 27867 268 27899
rect 300 27867 340 27899
rect 372 27867 412 27899
rect 444 27867 484 27899
rect 516 27867 556 27899
rect 588 27867 628 27899
rect 660 27867 700 27899
rect 732 27867 772 27899
rect 804 27867 844 27899
rect 876 27867 950 27899
rect 50 27827 950 27867
rect 50 27795 124 27827
rect 156 27795 196 27827
rect 228 27795 268 27827
rect 300 27795 340 27827
rect 372 27795 412 27827
rect 444 27795 484 27827
rect 516 27795 556 27827
rect 588 27795 628 27827
rect 660 27795 700 27827
rect 732 27795 772 27827
rect 804 27795 844 27827
rect 876 27795 950 27827
rect 50 27755 950 27795
rect 50 27723 124 27755
rect 156 27723 196 27755
rect 228 27723 268 27755
rect 300 27723 340 27755
rect 372 27723 412 27755
rect 444 27723 484 27755
rect 516 27723 556 27755
rect 588 27723 628 27755
rect 660 27723 700 27755
rect 732 27723 772 27755
rect 804 27723 844 27755
rect 876 27723 950 27755
rect 50 27683 950 27723
rect 50 27651 124 27683
rect 156 27651 196 27683
rect 228 27651 268 27683
rect 300 27651 340 27683
rect 372 27651 412 27683
rect 444 27651 484 27683
rect 516 27651 556 27683
rect 588 27651 628 27683
rect 660 27651 700 27683
rect 732 27651 772 27683
rect 804 27651 844 27683
rect 876 27651 950 27683
rect 50 27611 950 27651
rect 50 27579 124 27611
rect 156 27579 196 27611
rect 228 27579 268 27611
rect 300 27579 340 27611
rect 372 27579 412 27611
rect 444 27579 484 27611
rect 516 27579 556 27611
rect 588 27579 628 27611
rect 660 27579 700 27611
rect 732 27579 772 27611
rect 804 27579 844 27611
rect 876 27579 950 27611
rect 50 27539 950 27579
rect 50 27507 124 27539
rect 156 27507 196 27539
rect 228 27507 268 27539
rect 300 27507 340 27539
rect 372 27507 412 27539
rect 444 27507 484 27539
rect 516 27507 556 27539
rect 588 27507 628 27539
rect 660 27507 700 27539
rect 732 27507 772 27539
rect 804 27507 844 27539
rect 876 27507 950 27539
rect 50 27467 950 27507
rect 50 27435 124 27467
rect 156 27435 196 27467
rect 228 27435 268 27467
rect 300 27435 340 27467
rect 372 27435 412 27467
rect 444 27435 484 27467
rect 516 27435 556 27467
rect 588 27435 628 27467
rect 660 27435 700 27467
rect 732 27435 772 27467
rect 804 27435 844 27467
rect 876 27435 950 27467
rect 50 27395 950 27435
rect 50 27363 124 27395
rect 156 27363 196 27395
rect 228 27363 268 27395
rect 300 27363 340 27395
rect 372 27363 412 27395
rect 444 27363 484 27395
rect 516 27363 556 27395
rect 588 27363 628 27395
rect 660 27363 700 27395
rect 732 27363 772 27395
rect 804 27363 844 27395
rect 876 27363 950 27395
rect 50 27323 950 27363
rect 50 27291 124 27323
rect 156 27291 196 27323
rect 228 27291 268 27323
rect 300 27291 340 27323
rect 372 27291 412 27323
rect 444 27291 484 27323
rect 516 27291 556 27323
rect 588 27291 628 27323
rect 660 27291 700 27323
rect 732 27291 772 27323
rect 804 27291 844 27323
rect 876 27291 950 27323
rect 50 27251 950 27291
rect 50 27219 124 27251
rect 156 27219 196 27251
rect 228 27219 268 27251
rect 300 27219 340 27251
rect 372 27219 412 27251
rect 444 27219 484 27251
rect 516 27219 556 27251
rect 588 27219 628 27251
rect 660 27219 700 27251
rect 732 27219 772 27251
rect 804 27219 844 27251
rect 876 27219 950 27251
rect 50 27179 950 27219
rect 50 27147 124 27179
rect 156 27147 196 27179
rect 228 27147 268 27179
rect 300 27147 340 27179
rect 372 27147 412 27179
rect 444 27147 484 27179
rect 516 27147 556 27179
rect 588 27147 628 27179
rect 660 27147 700 27179
rect 732 27147 772 27179
rect 804 27147 844 27179
rect 876 27147 950 27179
rect 50 27107 950 27147
rect 50 27075 124 27107
rect 156 27075 196 27107
rect 228 27075 268 27107
rect 300 27075 340 27107
rect 372 27075 412 27107
rect 444 27075 484 27107
rect 516 27075 556 27107
rect 588 27075 628 27107
rect 660 27075 700 27107
rect 732 27075 772 27107
rect 804 27075 844 27107
rect 876 27075 950 27107
rect 50 27035 950 27075
rect 50 27003 124 27035
rect 156 27003 196 27035
rect 228 27003 268 27035
rect 300 27003 340 27035
rect 372 27003 412 27035
rect 444 27003 484 27035
rect 516 27003 556 27035
rect 588 27003 628 27035
rect 660 27003 700 27035
rect 732 27003 772 27035
rect 804 27003 844 27035
rect 876 27003 950 27035
rect 50 26963 950 27003
rect 50 26931 124 26963
rect 156 26931 196 26963
rect 228 26931 268 26963
rect 300 26931 340 26963
rect 372 26931 412 26963
rect 444 26931 484 26963
rect 516 26931 556 26963
rect 588 26931 628 26963
rect 660 26931 700 26963
rect 732 26931 772 26963
rect 804 26931 844 26963
rect 876 26931 950 26963
rect 50 26891 950 26931
rect 50 26859 124 26891
rect 156 26859 196 26891
rect 228 26859 268 26891
rect 300 26859 340 26891
rect 372 26859 412 26891
rect 444 26859 484 26891
rect 516 26859 556 26891
rect 588 26859 628 26891
rect 660 26859 700 26891
rect 732 26859 772 26891
rect 804 26859 844 26891
rect 876 26859 950 26891
rect 50 26819 950 26859
rect 50 26787 124 26819
rect 156 26787 196 26819
rect 228 26787 268 26819
rect 300 26787 340 26819
rect 372 26787 412 26819
rect 444 26787 484 26819
rect 516 26787 556 26819
rect 588 26787 628 26819
rect 660 26787 700 26819
rect 732 26787 772 26819
rect 804 26787 844 26819
rect 876 26787 950 26819
rect 50 26747 950 26787
rect 50 26715 124 26747
rect 156 26715 196 26747
rect 228 26715 268 26747
rect 300 26715 340 26747
rect 372 26715 412 26747
rect 444 26715 484 26747
rect 516 26715 556 26747
rect 588 26715 628 26747
rect 660 26715 700 26747
rect 732 26715 772 26747
rect 804 26715 844 26747
rect 876 26715 950 26747
rect 50 26675 950 26715
rect 50 26643 124 26675
rect 156 26643 196 26675
rect 228 26643 268 26675
rect 300 26643 340 26675
rect 372 26643 412 26675
rect 444 26643 484 26675
rect 516 26643 556 26675
rect 588 26643 628 26675
rect 660 26643 700 26675
rect 732 26643 772 26675
rect 804 26643 844 26675
rect 876 26643 950 26675
rect 50 26603 950 26643
rect 50 26571 124 26603
rect 156 26571 196 26603
rect 228 26571 268 26603
rect 300 26571 340 26603
rect 372 26571 412 26603
rect 444 26571 484 26603
rect 516 26571 556 26603
rect 588 26571 628 26603
rect 660 26571 700 26603
rect 732 26571 772 26603
rect 804 26571 844 26603
rect 876 26571 950 26603
rect 50 26531 950 26571
rect 50 26499 124 26531
rect 156 26499 196 26531
rect 228 26499 268 26531
rect 300 26499 340 26531
rect 372 26499 412 26531
rect 444 26499 484 26531
rect 516 26499 556 26531
rect 588 26499 628 26531
rect 660 26499 700 26531
rect 732 26499 772 26531
rect 804 26499 844 26531
rect 876 26499 950 26531
rect 50 26459 950 26499
rect 50 26427 124 26459
rect 156 26427 196 26459
rect 228 26427 268 26459
rect 300 26427 340 26459
rect 372 26427 412 26459
rect 444 26427 484 26459
rect 516 26427 556 26459
rect 588 26427 628 26459
rect 660 26427 700 26459
rect 732 26427 772 26459
rect 804 26427 844 26459
rect 876 26427 950 26459
rect 50 26387 950 26427
rect 50 26355 124 26387
rect 156 26355 196 26387
rect 228 26355 268 26387
rect 300 26355 340 26387
rect 372 26355 412 26387
rect 444 26355 484 26387
rect 516 26355 556 26387
rect 588 26355 628 26387
rect 660 26355 700 26387
rect 732 26355 772 26387
rect 804 26355 844 26387
rect 876 26355 950 26387
rect 50 26315 950 26355
rect 50 26283 124 26315
rect 156 26283 196 26315
rect 228 26283 268 26315
rect 300 26283 340 26315
rect 372 26283 412 26315
rect 444 26283 484 26315
rect 516 26283 556 26315
rect 588 26283 628 26315
rect 660 26283 700 26315
rect 732 26283 772 26315
rect 804 26283 844 26315
rect 876 26283 950 26315
rect 50 26243 950 26283
rect 50 26211 124 26243
rect 156 26211 196 26243
rect 228 26211 268 26243
rect 300 26211 340 26243
rect 372 26211 412 26243
rect 444 26211 484 26243
rect 516 26211 556 26243
rect 588 26211 628 26243
rect 660 26211 700 26243
rect 732 26211 772 26243
rect 804 26211 844 26243
rect 876 26211 950 26243
rect 50 26171 950 26211
rect 50 26139 124 26171
rect 156 26139 196 26171
rect 228 26139 268 26171
rect 300 26139 340 26171
rect 372 26139 412 26171
rect 444 26139 484 26171
rect 516 26139 556 26171
rect 588 26139 628 26171
rect 660 26139 700 26171
rect 732 26139 772 26171
rect 804 26139 844 26171
rect 876 26139 950 26171
rect 50 26099 950 26139
rect 50 26067 124 26099
rect 156 26067 196 26099
rect 228 26067 268 26099
rect 300 26067 340 26099
rect 372 26067 412 26099
rect 444 26067 484 26099
rect 516 26067 556 26099
rect 588 26067 628 26099
rect 660 26067 700 26099
rect 732 26067 772 26099
rect 804 26067 844 26099
rect 876 26067 950 26099
rect 50 26027 950 26067
rect 50 25995 124 26027
rect 156 25995 196 26027
rect 228 25995 268 26027
rect 300 25995 340 26027
rect 372 25995 412 26027
rect 444 25995 484 26027
rect 516 25995 556 26027
rect 588 25995 628 26027
rect 660 25995 700 26027
rect 732 25995 772 26027
rect 804 25995 844 26027
rect 876 25995 950 26027
rect 50 25955 950 25995
rect 50 25923 124 25955
rect 156 25923 196 25955
rect 228 25923 268 25955
rect 300 25923 340 25955
rect 372 25923 412 25955
rect 444 25923 484 25955
rect 516 25923 556 25955
rect 588 25923 628 25955
rect 660 25923 700 25955
rect 732 25923 772 25955
rect 804 25923 844 25955
rect 876 25923 950 25955
rect 50 25883 950 25923
rect 50 25851 124 25883
rect 156 25851 196 25883
rect 228 25851 268 25883
rect 300 25851 340 25883
rect 372 25851 412 25883
rect 444 25851 484 25883
rect 516 25851 556 25883
rect 588 25851 628 25883
rect 660 25851 700 25883
rect 732 25851 772 25883
rect 804 25851 844 25883
rect 876 25851 950 25883
rect 50 25811 950 25851
rect 50 25779 124 25811
rect 156 25779 196 25811
rect 228 25779 268 25811
rect 300 25779 340 25811
rect 372 25779 412 25811
rect 444 25779 484 25811
rect 516 25779 556 25811
rect 588 25779 628 25811
rect 660 25779 700 25811
rect 732 25779 772 25811
rect 804 25779 844 25811
rect 876 25779 950 25811
rect 50 25739 950 25779
rect 50 25707 124 25739
rect 156 25707 196 25739
rect 228 25707 268 25739
rect 300 25707 340 25739
rect 372 25707 412 25739
rect 444 25707 484 25739
rect 516 25707 556 25739
rect 588 25707 628 25739
rect 660 25707 700 25739
rect 732 25707 772 25739
rect 804 25707 844 25739
rect 876 25707 950 25739
rect 50 25667 950 25707
rect 50 25635 124 25667
rect 156 25635 196 25667
rect 228 25635 268 25667
rect 300 25635 340 25667
rect 372 25635 412 25667
rect 444 25635 484 25667
rect 516 25635 556 25667
rect 588 25635 628 25667
rect 660 25635 700 25667
rect 732 25635 772 25667
rect 804 25635 844 25667
rect 876 25635 950 25667
rect 50 25595 950 25635
rect 50 25563 124 25595
rect 156 25563 196 25595
rect 228 25563 268 25595
rect 300 25563 340 25595
rect 372 25563 412 25595
rect 444 25563 484 25595
rect 516 25563 556 25595
rect 588 25563 628 25595
rect 660 25563 700 25595
rect 732 25563 772 25595
rect 804 25563 844 25595
rect 876 25563 950 25595
rect 50 25523 950 25563
rect 50 25491 124 25523
rect 156 25491 196 25523
rect 228 25491 268 25523
rect 300 25491 340 25523
rect 372 25491 412 25523
rect 444 25491 484 25523
rect 516 25491 556 25523
rect 588 25491 628 25523
rect 660 25491 700 25523
rect 732 25491 772 25523
rect 804 25491 844 25523
rect 876 25491 950 25523
rect 50 25451 950 25491
rect 50 25419 124 25451
rect 156 25419 196 25451
rect 228 25419 268 25451
rect 300 25419 340 25451
rect 372 25419 412 25451
rect 444 25419 484 25451
rect 516 25419 556 25451
rect 588 25419 628 25451
rect 660 25419 700 25451
rect 732 25419 772 25451
rect 804 25419 844 25451
rect 876 25419 950 25451
rect 50 25379 950 25419
rect 50 25347 124 25379
rect 156 25347 196 25379
rect 228 25347 268 25379
rect 300 25347 340 25379
rect 372 25347 412 25379
rect 444 25347 484 25379
rect 516 25347 556 25379
rect 588 25347 628 25379
rect 660 25347 700 25379
rect 732 25347 772 25379
rect 804 25347 844 25379
rect 876 25347 950 25379
rect 50 25307 950 25347
rect 50 25275 124 25307
rect 156 25275 196 25307
rect 228 25275 268 25307
rect 300 25275 340 25307
rect 372 25275 412 25307
rect 444 25275 484 25307
rect 516 25275 556 25307
rect 588 25275 628 25307
rect 660 25275 700 25307
rect 732 25275 772 25307
rect 804 25275 844 25307
rect 876 25275 950 25307
rect 50 25235 950 25275
rect 50 25203 124 25235
rect 156 25203 196 25235
rect 228 25203 268 25235
rect 300 25203 340 25235
rect 372 25203 412 25235
rect 444 25203 484 25235
rect 516 25203 556 25235
rect 588 25203 628 25235
rect 660 25203 700 25235
rect 732 25203 772 25235
rect 804 25203 844 25235
rect 876 25203 950 25235
rect 50 25163 950 25203
rect 50 25131 124 25163
rect 156 25131 196 25163
rect 228 25131 268 25163
rect 300 25131 340 25163
rect 372 25131 412 25163
rect 444 25131 484 25163
rect 516 25131 556 25163
rect 588 25131 628 25163
rect 660 25131 700 25163
rect 732 25131 772 25163
rect 804 25131 844 25163
rect 876 25131 950 25163
rect 50 25091 950 25131
rect 50 25059 124 25091
rect 156 25059 196 25091
rect 228 25059 268 25091
rect 300 25059 340 25091
rect 372 25059 412 25091
rect 444 25059 484 25091
rect 516 25059 556 25091
rect 588 25059 628 25091
rect 660 25059 700 25091
rect 732 25059 772 25091
rect 804 25059 844 25091
rect 876 25059 950 25091
rect 50 25019 950 25059
rect 50 24987 124 25019
rect 156 24987 196 25019
rect 228 24987 268 25019
rect 300 24987 340 25019
rect 372 24987 412 25019
rect 444 24987 484 25019
rect 516 24987 556 25019
rect 588 24987 628 25019
rect 660 24987 700 25019
rect 732 24987 772 25019
rect 804 24987 844 25019
rect 876 24987 950 25019
rect 50 24947 950 24987
rect 50 24915 124 24947
rect 156 24915 196 24947
rect 228 24915 268 24947
rect 300 24915 340 24947
rect 372 24915 412 24947
rect 444 24915 484 24947
rect 516 24915 556 24947
rect 588 24915 628 24947
rect 660 24915 700 24947
rect 732 24915 772 24947
rect 804 24915 844 24947
rect 876 24915 950 24947
rect 50 24875 950 24915
rect 50 24843 124 24875
rect 156 24843 196 24875
rect 228 24843 268 24875
rect 300 24843 340 24875
rect 372 24843 412 24875
rect 444 24843 484 24875
rect 516 24843 556 24875
rect 588 24843 628 24875
rect 660 24843 700 24875
rect 732 24843 772 24875
rect 804 24843 844 24875
rect 876 24843 950 24875
rect 50 24803 950 24843
rect 50 24771 124 24803
rect 156 24771 196 24803
rect 228 24771 268 24803
rect 300 24771 340 24803
rect 372 24771 412 24803
rect 444 24771 484 24803
rect 516 24771 556 24803
rect 588 24771 628 24803
rect 660 24771 700 24803
rect 732 24771 772 24803
rect 804 24771 844 24803
rect 876 24771 950 24803
rect 50 24731 950 24771
rect 50 24699 124 24731
rect 156 24699 196 24731
rect 228 24699 268 24731
rect 300 24699 340 24731
rect 372 24699 412 24731
rect 444 24699 484 24731
rect 516 24699 556 24731
rect 588 24699 628 24731
rect 660 24699 700 24731
rect 732 24699 772 24731
rect 804 24699 844 24731
rect 876 24699 950 24731
rect 50 24659 950 24699
rect 50 24627 124 24659
rect 156 24627 196 24659
rect 228 24627 268 24659
rect 300 24627 340 24659
rect 372 24627 412 24659
rect 444 24627 484 24659
rect 516 24627 556 24659
rect 588 24627 628 24659
rect 660 24627 700 24659
rect 732 24627 772 24659
rect 804 24627 844 24659
rect 876 24627 950 24659
rect 50 24587 950 24627
rect 50 24555 124 24587
rect 156 24555 196 24587
rect 228 24555 268 24587
rect 300 24555 340 24587
rect 372 24555 412 24587
rect 444 24555 484 24587
rect 516 24555 556 24587
rect 588 24555 628 24587
rect 660 24555 700 24587
rect 732 24555 772 24587
rect 804 24555 844 24587
rect 876 24555 950 24587
rect 50 24515 950 24555
rect 50 24483 124 24515
rect 156 24483 196 24515
rect 228 24483 268 24515
rect 300 24483 340 24515
rect 372 24483 412 24515
rect 444 24483 484 24515
rect 516 24483 556 24515
rect 588 24483 628 24515
rect 660 24483 700 24515
rect 732 24483 772 24515
rect 804 24483 844 24515
rect 876 24483 950 24515
rect 50 24443 950 24483
rect 50 24411 124 24443
rect 156 24411 196 24443
rect 228 24411 268 24443
rect 300 24411 340 24443
rect 372 24411 412 24443
rect 444 24411 484 24443
rect 516 24411 556 24443
rect 588 24411 628 24443
rect 660 24411 700 24443
rect 732 24411 772 24443
rect 804 24411 844 24443
rect 876 24411 950 24443
rect 50 24371 950 24411
rect 50 24339 124 24371
rect 156 24339 196 24371
rect 228 24339 268 24371
rect 300 24339 340 24371
rect 372 24339 412 24371
rect 444 24339 484 24371
rect 516 24339 556 24371
rect 588 24339 628 24371
rect 660 24339 700 24371
rect 732 24339 772 24371
rect 804 24339 844 24371
rect 876 24339 950 24371
rect 50 24299 950 24339
rect 50 24267 124 24299
rect 156 24267 196 24299
rect 228 24267 268 24299
rect 300 24267 340 24299
rect 372 24267 412 24299
rect 444 24267 484 24299
rect 516 24267 556 24299
rect 588 24267 628 24299
rect 660 24267 700 24299
rect 732 24267 772 24299
rect 804 24267 844 24299
rect 876 24267 950 24299
rect 50 24227 950 24267
rect 50 24195 124 24227
rect 156 24195 196 24227
rect 228 24195 268 24227
rect 300 24195 340 24227
rect 372 24195 412 24227
rect 444 24195 484 24227
rect 516 24195 556 24227
rect 588 24195 628 24227
rect 660 24195 700 24227
rect 732 24195 772 24227
rect 804 24195 844 24227
rect 876 24195 950 24227
rect 50 24155 950 24195
rect 50 24123 124 24155
rect 156 24123 196 24155
rect 228 24123 268 24155
rect 300 24123 340 24155
rect 372 24123 412 24155
rect 444 24123 484 24155
rect 516 24123 556 24155
rect 588 24123 628 24155
rect 660 24123 700 24155
rect 732 24123 772 24155
rect 804 24123 844 24155
rect 876 24123 950 24155
rect 50 24083 950 24123
rect 50 24051 124 24083
rect 156 24051 196 24083
rect 228 24051 268 24083
rect 300 24051 340 24083
rect 372 24051 412 24083
rect 444 24051 484 24083
rect 516 24051 556 24083
rect 588 24051 628 24083
rect 660 24051 700 24083
rect 732 24051 772 24083
rect 804 24051 844 24083
rect 876 24051 950 24083
rect 50 24011 950 24051
rect 50 23979 124 24011
rect 156 23979 196 24011
rect 228 23979 268 24011
rect 300 23979 340 24011
rect 372 23979 412 24011
rect 444 23979 484 24011
rect 516 23979 556 24011
rect 588 23979 628 24011
rect 660 23979 700 24011
rect 732 23979 772 24011
rect 804 23979 844 24011
rect 876 23979 950 24011
rect 50 23939 950 23979
rect 50 23907 124 23939
rect 156 23907 196 23939
rect 228 23907 268 23939
rect 300 23907 340 23939
rect 372 23907 412 23939
rect 444 23907 484 23939
rect 516 23907 556 23939
rect 588 23907 628 23939
rect 660 23907 700 23939
rect 732 23907 772 23939
rect 804 23907 844 23939
rect 876 23907 950 23939
rect 50 23867 950 23907
rect 50 23835 124 23867
rect 156 23835 196 23867
rect 228 23835 268 23867
rect 300 23835 340 23867
rect 372 23835 412 23867
rect 444 23835 484 23867
rect 516 23835 556 23867
rect 588 23835 628 23867
rect 660 23835 700 23867
rect 732 23835 772 23867
rect 804 23835 844 23867
rect 876 23835 950 23867
rect 50 23795 950 23835
rect 50 23763 124 23795
rect 156 23763 196 23795
rect 228 23763 268 23795
rect 300 23763 340 23795
rect 372 23763 412 23795
rect 444 23763 484 23795
rect 516 23763 556 23795
rect 588 23763 628 23795
rect 660 23763 700 23795
rect 732 23763 772 23795
rect 804 23763 844 23795
rect 876 23763 950 23795
rect 50 23723 950 23763
rect 50 23691 124 23723
rect 156 23691 196 23723
rect 228 23691 268 23723
rect 300 23691 340 23723
rect 372 23691 412 23723
rect 444 23691 484 23723
rect 516 23691 556 23723
rect 588 23691 628 23723
rect 660 23691 700 23723
rect 732 23691 772 23723
rect 804 23691 844 23723
rect 876 23691 950 23723
rect 50 23651 950 23691
rect 50 23619 124 23651
rect 156 23619 196 23651
rect 228 23619 268 23651
rect 300 23619 340 23651
rect 372 23619 412 23651
rect 444 23619 484 23651
rect 516 23619 556 23651
rect 588 23619 628 23651
rect 660 23619 700 23651
rect 732 23619 772 23651
rect 804 23619 844 23651
rect 876 23619 950 23651
rect 50 23579 950 23619
rect 50 23547 124 23579
rect 156 23547 196 23579
rect 228 23547 268 23579
rect 300 23547 340 23579
rect 372 23547 412 23579
rect 444 23547 484 23579
rect 516 23547 556 23579
rect 588 23547 628 23579
rect 660 23547 700 23579
rect 732 23547 772 23579
rect 804 23547 844 23579
rect 876 23547 950 23579
rect 50 23507 950 23547
rect 50 23475 124 23507
rect 156 23475 196 23507
rect 228 23475 268 23507
rect 300 23475 340 23507
rect 372 23475 412 23507
rect 444 23475 484 23507
rect 516 23475 556 23507
rect 588 23475 628 23507
rect 660 23475 700 23507
rect 732 23475 772 23507
rect 804 23475 844 23507
rect 876 23475 950 23507
rect 50 23435 950 23475
rect 50 23403 124 23435
rect 156 23403 196 23435
rect 228 23403 268 23435
rect 300 23403 340 23435
rect 372 23403 412 23435
rect 444 23403 484 23435
rect 516 23403 556 23435
rect 588 23403 628 23435
rect 660 23403 700 23435
rect 732 23403 772 23435
rect 804 23403 844 23435
rect 876 23403 950 23435
rect 50 23363 950 23403
rect 50 23331 124 23363
rect 156 23331 196 23363
rect 228 23331 268 23363
rect 300 23331 340 23363
rect 372 23331 412 23363
rect 444 23331 484 23363
rect 516 23331 556 23363
rect 588 23331 628 23363
rect 660 23331 700 23363
rect 732 23331 772 23363
rect 804 23331 844 23363
rect 876 23331 950 23363
rect 50 23291 950 23331
rect 50 23259 124 23291
rect 156 23259 196 23291
rect 228 23259 268 23291
rect 300 23259 340 23291
rect 372 23259 412 23291
rect 444 23259 484 23291
rect 516 23259 556 23291
rect 588 23259 628 23291
rect 660 23259 700 23291
rect 732 23259 772 23291
rect 804 23259 844 23291
rect 876 23259 950 23291
rect 50 23219 950 23259
rect 50 23187 124 23219
rect 156 23187 196 23219
rect 228 23187 268 23219
rect 300 23187 340 23219
rect 372 23187 412 23219
rect 444 23187 484 23219
rect 516 23187 556 23219
rect 588 23187 628 23219
rect 660 23187 700 23219
rect 732 23187 772 23219
rect 804 23187 844 23219
rect 876 23187 950 23219
rect 50 23124 950 23187
rect 50 22874 950 22924
rect 50 22842 124 22874
rect 156 22842 196 22874
rect 228 22842 268 22874
rect 300 22842 340 22874
rect 372 22842 412 22874
rect 444 22842 484 22874
rect 516 22842 556 22874
rect 588 22842 628 22874
rect 660 22842 700 22874
rect 732 22842 772 22874
rect 804 22842 844 22874
rect 876 22842 950 22874
rect 50 22802 950 22842
rect 50 22770 124 22802
rect 156 22770 196 22802
rect 228 22770 268 22802
rect 300 22770 340 22802
rect 372 22770 412 22802
rect 444 22770 484 22802
rect 516 22770 556 22802
rect 588 22770 628 22802
rect 660 22770 700 22802
rect 732 22770 772 22802
rect 804 22770 844 22802
rect 876 22770 950 22802
rect 50 22730 950 22770
rect 50 22698 124 22730
rect 156 22698 196 22730
rect 228 22698 268 22730
rect 300 22698 340 22730
rect 372 22698 412 22730
rect 444 22698 484 22730
rect 516 22698 556 22730
rect 588 22698 628 22730
rect 660 22698 700 22730
rect 732 22698 772 22730
rect 804 22698 844 22730
rect 876 22698 950 22730
rect 50 22658 950 22698
rect 50 22626 124 22658
rect 156 22626 196 22658
rect 228 22626 268 22658
rect 300 22626 340 22658
rect 372 22626 412 22658
rect 444 22626 484 22658
rect 516 22626 556 22658
rect 588 22626 628 22658
rect 660 22626 700 22658
rect 732 22626 772 22658
rect 804 22626 844 22658
rect 876 22626 950 22658
rect 50 22586 950 22626
rect 50 22554 124 22586
rect 156 22554 196 22586
rect 228 22554 268 22586
rect 300 22554 340 22586
rect 372 22554 412 22586
rect 444 22554 484 22586
rect 516 22554 556 22586
rect 588 22554 628 22586
rect 660 22554 700 22586
rect 732 22554 772 22586
rect 804 22554 844 22586
rect 876 22554 950 22586
rect 50 22514 950 22554
rect 50 22482 124 22514
rect 156 22482 196 22514
rect 228 22482 268 22514
rect 300 22482 340 22514
rect 372 22482 412 22514
rect 444 22482 484 22514
rect 516 22482 556 22514
rect 588 22482 628 22514
rect 660 22482 700 22514
rect 732 22482 772 22514
rect 804 22482 844 22514
rect 876 22482 950 22514
rect 50 22442 950 22482
rect 50 22410 124 22442
rect 156 22410 196 22442
rect 228 22410 268 22442
rect 300 22410 340 22442
rect 372 22410 412 22442
rect 444 22410 484 22442
rect 516 22410 556 22442
rect 588 22410 628 22442
rect 660 22410 700 22442
rect 732 22410 772 22442
rect 804 22410 844 22442
rect 876 22410 950 22442
rect 50 22370 950 22410
rect 50 22338 124 22370
rect 156 22338 196 22370
rect 228 22338 268 22370
rect 300 22338 340 22370
rect 372 22338 412 22370
rect 444 22338 484 22370
rect 516 22338 556 22370
rect 588 22338 628 22370
rect 660 22338 700 22370
rect 732 22338 772 22370
rect 804 22338 844 22370
rect 876 22338 950 22370
rect 50 22298 950 22338
rect 50 22266 124 22298
rect 156 22266 196 22298
rect 228 22266 268 22298
rect 300 22266 340 22298
rect 372 22266 412 22298
rect 444 22266 484 22298
rect 516 22266 556 22298
rect 588 22266 628 22298
rect 660 22266 700 22298
rect 732 22266 772 22298
rect 804 22266 844 22298
rect 876 22266 950 22298
rect 50 22226 950 22266
rect 50 22194 124 22226
rect 156 22194 196 22226
rect 228 22194 268 22226
rect 300 22194 340 22226
rect 372 22194 412 22226
rect 444 22194 484 22226
rect 516 22194 556 22226
rect 588 22194 628 22226
rect 660 22194 700 22226
rect 732 22194 772 22226
rect 804 22194 844 22226
rect 876 22194 950 22226
rect 50 22154 950 22194
rect 50 22122 124 22154
rect 156 22122 196 22154
rect 228 22122 268 22154
rect 300 22122 340 22154
rect 372 22122 412 22154
rect 444 22122 484 22154
rect 516 22122 556 22154
rect 588 22122 628 22154
rect 660 22122 700 22154
rect 732 22122 772 22154
rect 804 22122 844 22154
rect 876 22122 950 22154
rect 50 22082 950 22122
rect 50 22050 124 22082
rect 156 22050 196 22082
rect 228 22050 268 22082
rect 300 22050 340 22082
rect 372 22050 412 22082
rect 444 22050 484 22082
rect 516 22050 556 22082
rect 588 22050 628 22082
rect 660 22050 700 22082
rect 732 22050 772 22082
rect 804 22050 844 22082
rect 876 22050 950 22082
rect 50 22010 950 22050
rect 50 21978 124 22010
rect 156 21978 196 22010
rect 228 21978 268 22010
rect 300 21978 340 22010
rect 372 21978 412 22010
rect 444 21978 484 22010
rect 516 21978 556 22010
rect 588 21978 628 22010
rect 660 21978 700 22010
rect 732 21978 772 22010
rect 804 21978 844 22010
rect 876 21978 950 22010
rect 50 21938 950 21978
rect 50 21906 124 21938
rect 156 21906 196 21938
rect 228 21906 268 21938
rect 300 21906 340 21938
rect 372 21906 412 21938
rect 444 21906 484 21938
rect 516 21906 556 21938
rect 588 21906 628 21938
rect 660 21906 700 21938
rect 732 21906 772 21938
rect 804 21906 844 21938
rect 876 21906 950 21938
rect 50 21866 950 21906
rect 50 21834 124 21866
rect 156 21834 196 21866
rect 228 21834 268 21866
rect 300 21834 340 21866
rect 372 21834 412 21866
rect 444 21834 484 21866
rect 516 21834 556 21866
rect 588 21834 628 21866
rect 660 21834 700 21866
rect 732 21834 772 21866
rect 804 21834 844 21866
rect 876 21834 950 21866
rect 50 21794 950 21834
rect 50 21762 124 21794
rect 156 21762 196 21794
rect 228 21762 268 21794
rect 300 21762 340 21794
rect 372 21762 412 21794
rect 444 21762 484 21794
rect 516 21762 556 21794
rect 588 21762 628 21794
rect 660 21762 700 21794
rect 732 21762 772 21794
rect 804 21762 844 21794
rect 876 21762 950 21794
rect 50 21722 950 21762
rect 50 21690 124 21722
rect 156 21690 196 21722
rect 228 21690 268 21722
rect 300 21690 340 21722
rect 372 21690 412 21722
rect 444 21690 484 21722
rect 516 21690 556 21722
rect 588 21690 628 21722
rect 660 21690 700 21722
rect 732 21690 772 21722
rect 804 21690 844 21722
rect 876 21690 950 21722
rect 50 21650 950 21690
rect 50 21618 124 21650
rect 156 21618 196 21650
rect 228 21618 268 21650
rect 300 21618 340 21650
rect 372 21618 412 21650
rect 444 21618 484 21650
rect 516 21618 556 21650
rect 588 21618 628 21650
rect 660 21618 700 21650
rect 732 21618 772 21650
rect 804 21618 844 21650
rect 876 21618 950 21650
rect 50 21578 950 21618
rect 50 21546 124 21578
rect 156 21546 196 21578
rect 228 21546 268 21578
rect 300 21546 340 21578
rect 372 21546 412 21578
rect 444 21546 484 21578
rect 516 21546 556 21578
rect 588 21546 628 21578
rect 660 21546 700 21578
rect 732 21546 772 21578
rect 804 21546 844 21578
rect 876 21546 950 21578
rect 50 21506 950 21546
rect 50 21474 124 21506
rect 156 21474 196 21506
rect 228 21474 268 21506
rect 300 21474 340 21506
rect 372 21474 412 21506
rect 444 21474 484 21506
rect 516 21474 556 21506
rect 588 21474 628 21506
rect 660 21474 700 21506
rect 732 21474 772 21506
rect 804 21474 844 21506
rect 876 21474 950 21506
rect 50 21434 950 21474
rect 50 21402 124 21434
rect 156 21402 196 21434
rect 228 21402 268 21434
rect 300 21402 340 21434
rect 372 21402 412 21434
rect 444 21402 484 21434
rect 516 21402 556 21434
rect 588 21402 628 21434
rect 660 21402 700 21434
rect 732 21402 772 21434
rect 804 21402 844 21434
rect 876 21402 950 21434
rect 50 21362 950 21402
rect 50 21330 124 21362
rect 156 21330 196 21362
rect 228 21330 268 21362
rect 300 21330 340 21362
rect 372 21330 412 21362
rect 444 21330 484 21362
rect 516 21330 556 21362
rect 588 21330 628 21362
rect 660 21330 700 21362
rect 732 21330 772 21362
rect 804 21330 844 21362
rect 876 21330 950 21362
rect 50 21290 950 21330
rect 50 21258 124 21290
rect 156 21258 196 21290
rect 228 21258 268 21290
rect 300 21258 340 21290
rect 372 21258 412 21290
rect 444 21258 484 21290
rect 516 21258 556 21290
rect 588 21258 628 21290
rect 660 21258 700 21290
rect 732 21258 772 21290
rect 804 21258 844 21290
rect 876 21258 950 21290
rect 50 21218 950 21258
rect 50 21186 124 21218
rect 156 21186 196 21218
rect 228 21186 268 21218
rect 300 21186 340 21218
rect 372 21186 412 21218
rect 444 21186 484 21218
rect 516 21186 556 21218
rect 588 21186 628 21218
rect 660 21186 700 21218
rect 732 21186 772 21218
rect 804 21186 844 21218
rect 876 21186 950 21218
rect 50 21146 950 21186
rect 50 21114 124 21146
rect 156 21114 196 21146
rect 228 21114 268 21146
rect 300 21114 340 21146
rect 372 21114 412 21146
rect 444 21114 484 21146
rect 516 21114 556 21146
rect 588 21114 628 21146
rect 660 21114 700 21146
rect 732 21114 772 21146
rect 804 21114 844 21146
rect 876 21114 950 21146
rect 50 21074 950 21114
rect 50 21042 124 21074
rect 156 21042 196 21074
rect 228 21042 268 21074
rect 300 21042 340 21074
rect 372 21042 412 21074
rect 444 21042 484 21074
rect 516 21042 556 21074
rect 588 21042 628 21074
rect 660 21042 700 21074
rect 732 21042 772 21074
rect 804 21042 844 21074
rect 876 21042 950 21074
rect 50 21002 950 21042
rect 50 20970 124 21002
rect 156 20970 196 21002
rect 228 20970 268 21002
rect 300 20970 340 21002
rect 372 20970 412 21002
rect 444 20970 484 21002
rect 516 20970 556 21002
rect 588 20970 628 21002
rect 660 20970 700 21002
rect 732 20970 772 21002
rect 804 20970 844 21002
rect 876 20970 950 21002
rect 50 20930 950 20970
rect 50 20898 124 20930
rect 156 20898 196 20930
rect 228 20898 268 20930
rect 300 20898 340 20930
rect 372 20898 412 20930
rect 444 20898 484 20930
rect 516 20898 556 20930
rect 588 20898 628 20930
rect 660 20898 700 20930
rect 732 20898 772 20930
rect 804 20898 844 20930
rect 876 20898 950 20930
rect 50 20858 950 20898
rect 50 20826 124 20858
rect 156 20826 196 20858
rect 228 20826 268 20858
rect 300 20826 340 20858
rect 372 20826 412 20858
rect 444 20826 484 20858
rect 516 20826 556 20858
rect 588 20826 628 20858
rect 660 20826 700 20858
rect 732 20826 772 20858
rect 804 20826 844 20858
rect 876 20826 950 20858
rect 50 20786 950 20826
rect 50 20754 124 20786
rect 156 20754 196 20786
rect 228 20754 268 20786
rect 300 20754 340 20786
rect 372 20754 412 20786
rect 444 20754 484 20786
rect 516 20754 556 20786
rect 588 20754 628 20786
rect 660 20754 700 20786
rect 732 20754 772 20786
rect 804 20754 844 20786
rect 876 20754 950 20786
rect 50 20714 950 20754
rect 50 20682 124 20714
rect 156 20682 196 20714
rect 228 20682 268 20714
rect 300 20682 340 20714
rect 372 20682 412 20714
rect 444 20682 484 20714
rect 516 20682 556 20714
rect 588 20682 628 20714
rect 660 20682 700 20714
rect 732 20682 772 20714
rect 804 20682 844 20714
rect 876 20682 950 20714
rect 50 20642 950 20682
rect 50 20610 124 20642
rect 156 20610 196 20642
rect 228 20610 268 20642
rect 300 20610 340 20642
rect 372 20610 412 20642
rect 444 20610 484 20642
rect 516 20610 556 20642
rect 588 20610 628 20642
rect 660 20610 700 20642
rect 732 20610 772 20642
rect 804 20610 844 20642
rect 876 20610 950 20642
rect 50 20570 950 20610
rect 50 20538 124 20570
rect 156 20538 196 20570
rect 228 20538 268 20570
rect 300 20538 340 20570
rect 372 20538 412 20570
rect 444 20538 484 20570
rect 516 20538 556 20570
rect 588 20538 628 20570
rect 660 20538 700 20570
rect 732 20538 772 20570
rect 804 20538 844 20570
rect 876 20538 950 20570
rect 50 20498 950 20538
rect 50 20466 124 20498
rect 156 20466 196 20498
rect 228 20466 268 20498
rect 300 20466 340 20498
rect 372 20466 412 20498
rect 444 20466 484 20498
rect 516 20466 556 20498
rect 588 20466 628 20498
rect 660 20466 700 20498
rect 732 20466 772 20498
rect 804 20466 844 20498
rect 876 20466 950 20498
rect 50 20426 950 20466
rect 50 20394 124 20426
rect 156 20394 196 20426
rect 228 20394 268 20426
rect 300 20394 340 20426
rect 372 20394 412 20426
rect 444 20394 484 20426
rect 516 20394 556 20426
rect 588 20394 628 20426
rect 660 20394 700 20426
rect 732 20394 772 20426
rect 804 20394 844 20426
rect 876 20394 950 20426
rect 50 20354 950 20394
rect 50 20322 124 20354
rect 156 20322 196 20354
rect 228 20322 268 20354
rect 300 20322 340 20354
rect 372 20322 412 20354
rect 444 20322 484 20354
rect 516 20322 556 20354
rect 588 20322 628 20354
rect 660 20322 700 20354
rect 732 20322 772 20354
rect 804 20322 844 20354
rect 876 20322 950 20354
rect 50 20282 950 20322
rect 50 20250 124 20282
rect 156 20250 196 20282
rect 228 20250 268 20282
rect 300 20250 340 20282
rect 372 20250 412 20282
rect 444 20250 484 20282
rect 516 20250 556 20282
rect 588 20250 628 20282
rect 660 20250 700 20282
rect 732 20250 772 20282
rect 804 20250 844 20282
rect 876 20250 950 20282
rect 50 20210 950 20250
rect 50 20178 124 20210
rect 156 20178 196 20210
rect 228 20178 268 20210
rect 300 20178 340 20210
rect 372 20178 412 20210
rect 444 20178 484 20210
rect 516 20178 556 20210
rect 588 20178 628 20210
rect 660 20178 700 20210
rect 732 20178 772 20210
rect 804 20178 844 20210
rect 876 20178 950 20210
rect 50 20138 950 20178
rect 50 20106 124 20138
rect 156 20106 196 20138
rect 228 20106 268 20138
rect 300 20106 340 20138
rect 372 20106 412 20138
rect 444 20106 484 20138
rect 516 20106 556 20138
rect 588 20106 628 20138
rect 660 20106 700 20138
rect 732 20106 772 20138
rect 804 20106 844 20138
rect 876 20106 950 20138
rect 50 20066 950 20106
rect 50 20034 124 20066
rect 156 20034 196 20066
rect 228 20034 268 20066
rect 300 20034 340 20066
rect 372 20034 412 20066
rect 444 20034 484 20066
rect 516 20034 556 20066
rect 588 20034 628 20066
rect 660 20034 700 20066
rect 732 20034 772 20066
rect 804 20034 844 20066
rect 876 20034 950 20066
rect 50 19994 950 20034
rect 50 19962 124 19994
rect 156 19962 196 19994
rect 228 19962 268 19994
rect 300 19962 340 19994
rect 372 19962 412 19994
rect 444 19962 484 19994
rect 516 19962 556 19994
rect 588 19962 628 19994
rect 660 19962 700 19994
rect 732 19962 772 19994
rect 804 19962 844 19994
rect 876 19962 950 19994
rect 50 19922 950 19962
rect 50 19890 124 19922
rect 156 19890 196 19922
rect 228 19890 268 19922
rect 300 19890 340 19922
rect 372 19890 412 19922
rect 444 19890 484 19922
rect 516 19890 556 19922
rect 588 19890 628 19922
rect 660 19890 700 19922
rect 732 19890 772 19922
rect 804 19890 844 19922
rect 876 19890 950 19922
rect 50 19850 950 19890
rect 50 19818 124 19850
rect 156 19818 196 19850
rect 228 19818 268 19850
rect 300 19818 340 19850
rect 372 19818 412 19850
rect 444 19818 484 19850
rect 516 19818 556 19850
rect 588 19818 628 19850
rect 660 19818 700 19850
rect 732 19818 772 19850
rect 804 19818 844 19850
rect 876 19818 950 19850
rect 50 19778 950 19818
rect 50 19746 124 19778
rect 156 19746 196 19778
rect 228 19746 268 19778
rect 300 19746 340 19778
rect 372 19746 412 19778
rect 444 19746 484 19778
rect 516 19746 556 19778
rect 588 19746 628 19778
rect 660 19746 700 19778
rect 732 19746 772 19778
rect 804 19746 844 19778
rect 876 19746 950 19778
rect 50 19706 950 19746
rect 50 19674 124 19706
rect 156 19674 196 19706
rect 228 19674 268 19706
rect 300 19674 340 19706
rect 372 19674 412 19706
rect 444 19674 484 19706
rect 516 19674 556 19706
rect 588 19674 628 19706
rect 660 19674 700 19706
rect 732 19674 772 19706
rect 804 19674 844 19706
rect 876 19674 950 19706
rect 50 19634 950 19674
rect 50 19602 124 19634
rect 156 19602 196 19634
rect 228 19602 268 19634
rect 300 19602 340 19634
rect 372 19602 412 19634
rect 444 19602 484 19634
rect 516 19602 556 19634
rect 588 19602 628 19634
rect 660 19602 700 19634
rect 732 19602 772 19634
rect 804 19602 844 19634
rect 876 19602 950 19634
rect 50 19562 950 19602
rect 50 19530 124 19562
rect 156 19530 196 19562
rect 228 19530 268 19562
rect 300 19530 340 19562
rect 372 19530 412 19562
rect 444 19530 484 19562
rect 516 19530 556 19562
rect 588 19530 628 19562
rect 660 19530 700 19562
rect 732 19530 772 19562
rect 804 19530 844 19562
rect 876 19530 950 19562
rect 50 19490 950 19530
rect 50 19458 124 19490
rect 156 19458 196 19490
rect 228 19458 268 19490
rect 300 19458 340 19490
rect 372 19458 412 19490
rect 444 19458 484 19490
rect 516 19458 556 19490
rect 588 19458 628 19490
rect 660 19458 700 19490
rect 732 19458 772 19490
rect 804 19458 844 19490
rect 876 19458 950 19490
rect 50 19418 950 19458
rect 50 19386 124 19418
rect 156 19386 196 19418
rect 228 19386 268 19418
rect 300 19386 340 19418
rect 372 19386 412 19418
rect 444 19386 484 19418
rect 516 19386 556 19418
rect 588 19386 628 19418
rect 660 19386 700 19418
rect 732 19386 772 19418
rect 804 19386 844 19418
rect 876 19386 950 19418
rect 50 19346 950 19386
rect 50 19314 124 19346
rect 156 19314 196 19346
rect 228 19314 268 19346
rect 300 19314 340 19346
rect 372 19314 412 19346
rect 444 19314 484 19346
rect 516 19314 556 19346
rect 588 19314 628 19346
rect 660 19314 700 19346
rect 732 19314 772 19346
rect 804 19314 844 19346
rect 876 19314 950 19346
rect 50 19274 950 19314
rect 50 19242 124 19274
rect 156 19242 196 19274
rect 228 19242 268 19274
rect 300 19242 340 19274
rect 372 19242 412 19274
rect 444 19242 484 19274
rect 516 19242 556 19274
rect 588 19242 628 19274
rect 660 19242 700 19274
rect 732 19242 772 19274
rect 804 19242 844 19274
rect 876 19242 950 19274
rect 50 19202 950 19242
rect 50 19170 124 19202
rect 156 19170 196 19202
rect 228 19170 268 19202
rect 300 19170 340 19202
rect 372 19170 412 19202
rect 444 19170 484 19202
rect 516 19170 556 19202
rect 588 19170 628 19202
rect 660 19170 700 19202
rect 732 19170 772 19202
rect 804 19170 844 19202
rect 876 19170 950 19202
rect 50 19130 950 19170
rect 50 19098 124 19130
rect 156 19098 196 19130
rect 228 19098 268 19130
rect 300 19098 340 19130
rect 372 19098 412 19130
rect 444 19098 484 19130
rect 516 19098 556 19130
rect 588 19098 628 19130
rect 660 19098 700 19130
rect 732 19098 772 19130
rect 804 19098 844 19130
rect 876 19098 950 19130
rect 50 19058 950 19098
rect 50 19026 124 19058
rect 156 19026 196 19058
rect 228 19026 268 19058
rect 300 19026 340 19058
rect 372 19026 412 19058
rect 444 19026 484 19058
rect 516 19026 556 19058
rect 588 19026 628 19058
rect 660 19026 700 19058
rect 732 19026 772 19058
rect 804 19026 844 19058
rect 876 19026 950 19058
rect 50 18986 950 19026
rect 50 18954 124 18986
rect 156 18954 196 18986
rect 228 18954 268 18986
rect 300 18954 340 18986
rect 372 18954 412 18986
rect 444 18954 484 18986
rect 516 18954 556 18986
rect 588 18954 628 18986
rect 660 18954 700 18986
rect 732 18954 772 18986
rect 804 18954 844 18986
rect 876 18954 950 18986
rect 50 18914 950 18954
rect 50 18882 124 18914
rect 156 18882 196 18914
rect 228 18882 268 18914
rect 300 18882 340 18914
rect 372 18882 412 18914
rect 444 18882 484 18914
rect 516 18882 556 18914
rect 588 18882 628 18914
rect 660 18882 700 18914
rect 732 18882 772 18914
rect 804 18882 844 18914
rect 876 18882 950 18914
rect 50 18842 950 18882
rect 50 18810 124 18842
rect 156 18810 196 18842
rect 228 18810 268 18842
rect 300 18810 340 18842
rect 372 18810 412 18842
rect 444 18810 484 18842
rect 516 18810 556 18842
rect 588 18810 628 18842
rect 660 18810 700 18842
rect 732 18810 772 18842
rect 804 18810 844 18842
rect 876 18810 950 18842
rect 50 18770 950 18810
rect 50 18738 124 18770
rect 156 18738 196 18770
rect 228 18738 268 18770
rect 300 18738 340 18770
rect 372 18738 412 18770
rect 444 18738 484 18770
rect 516 18738 556 18770
rect 588 18738 628 18770
rect 660 18738 700 18770
rect 732 18738 772 18770
rect 804 18738 844 18770
rect 876 18738 950 18770
rect 50 18698 950 18738
rect 50 18666 124 18698
rect 156 18666 196 18698
rect 228 18666 268 18698
rect 300 18666 340 18698
rect 372 18666 412 18698
rect 444 18666 484 18698
rect 516 18666 556 18698
rect 588 18666 628 18698
rect 660 18666 700 18698
rect 732 18666 772 18698
rect 804 18666 844 18698
rect 876 18666 950 18698
rect 50 18626 950 18666
rect 50 18594 124 18626
rect 156 18594 196 18626
rect 228 18594 268 18626
rect 300 18594 340 18626
rect 372 18594 412 18626
rect 444 18594 484 18626
rect 516 18594 556 18626
rect 588 18594 628 18626
rect 660 18594 700 18626
rect 732 18594 772 18626
rect 804 18594 844 18626
rect 876 18594 950 18626
rect 50 18554 950 18594
rect 50 18522 124 18554
rect 156 18522 196 18554
rect 228 18522 268 18554
rect 300 18522 340 18554
rect 372 18522 412 18554
rect 444 18522 484 18554
rect 516 18522 556 18554
rect 588 18522 628 18554
rect 660 18522 700 18554
rect 732 18522 772 18554
rect 804 18522 844 18554
rect 876 18522 950 18554
rect 50 18482 950 18522
rect 50 18450 124 18482
rect 156 18450 196 18482
rect 228 18450 268 18482
rect 300 18450 340 18482
rect 372 18450 412 18482
rect 444 18450 484 18482
rect 516 18450 556 18482
rect 588 18450 628 18482
rect 660 18450 700 18482
rect 732 18450 772 18482
rect 804 18450 844 18482
rect 876 18450 950 18482
rect 50 18410 950 18450
rect 50 18378 124 18410
rect 156 18378 196 18410
rect 228 18378 268 18410
rect 300 18378 340 18410
rect 372 18378 412 18410
rect 444 18378 484 18410
rect 516 18378 556 18410
rect 588 18378 628 18410
rect 660 18378 700 18410
rect 732 18378 772 18410
rect 804 18378 844 18410
rect 876 18378 950 18410
rect 50 18338 950 18378
rect 50 18306 124 18338
rect 156 18306 196 18338
rect 228 18306 268 18338
rect 300 18306 340 18338
rect 372 18306 412 18338
rect 444 18306 484 18338
rect 516 18306 556 18338
rect 588 18306 628 18338
rect 660 18306 700 18338
rect 732 18306 772 18338
rect 804 18306 844 18338
rect 876 18306 950 18338
rect 50 18266 950 18306
rect 50 18234 124 18266
rect 156 18234 196 18266
rect 228 18234 268 18266
rect 300 18234 340 18266
rect 372 18234 412 18266
rect 444 18234 484 18266
rect 516 18234 556 18266
rect 588 18234 628 18266
rect 660 18234 700 18266
rect 732 18234 772 18266
rect 804 18234 844 18266
rect 876 18234 950 18266
rect 50 18194 950 18234
rect 50 18162 124 18194
rect 156 18162 196 18194
rect 228 18162 268 18194
rect 300 18162 340 18194
rect 372 18162 412 18194
rect 444 18162 484 18194
rect 516 18162 556 18194
rect 588 18162 628 18194
rect 660 18162 700 18194
rect 732 18162 772 18194
rect 804 18162 844 18194
rect 876 18162 950 18194
rect 50 18112 950 18162
rect 50 17848 950 17912
rect 50 17816 124 17848
rect 156 17816 196 17848
rect 228 17816 268 17848
rect 300 17816 340 17848
rect 372 17816 412 17848
rect 444 17816 484 17848
rect 516 17816 556 17848
rect 588 17816 628 17848
rect 660 17816 700 17848
rect 732 17816 772 17848
rect 804 17816 844 17848
rect 876 17816 950 17848
rect 50 17776 950 17816
rect 50 17744 124 17776
rect 156 17744 196 17776
rect 228 17744 268 17776
rect 300 17744 340 17776
rect 372 17744 412 17776
rect 444 17744 484 17776
rect 516 17744 556 17776
rect 588 17744 628 17776
rect 660 17744 700 17776
rect 732 17744 772 17776
rect 804 17744 844 17776
rect 876 17744 950 17776
rect 50 17704 950 17744
rect 50 17672 124 17704
rect 156 17672 196 17704
rect 228 17672 268 17704
rect 300 17672 340 17704
rect 372 17672 412 17704
rect 444 17672 484 17704
rect 516 17672 556 17704
rect 588 17672 628 17704
rect 660 17672 700 17704
rect 732 17672 772 17704
rect 804 17672 844 17704
rect 876 17672 950 17704
rect 50 17632 950 17672
rect 50 17600 124 17632
rect 156 17600 196 17632
rect 228 17600 268 17632
rect 300 17600 340 17632
rect 372 17600 412 17632
rect 444 17600 484 17632
rect 516 17600 556 17632
rect 588 17600 628 17632
rect 660 17600 700 17632
rect 732 17600 772 17632
rect 804 17600 844 17632
rect 876 17600 950 17632
rect 50 17560 950 17600
rect 50 17528 124 17560
rect 156 17528 196 17560
rect 228 17528 268 17560
rect 300 17528 340 17560
rect 372 17528 412 17560
rect 444 17528 484 17560
rect 516 17528 556 17560
rect 588 17528 628 17560
rect 660 17528 700 17560
rect 732 17528 772 17560
rect 804 17528 844 17560
rect 876 17528 950 17560
rect 50 17488 950 17528
rect 50 17456 124 17488
rect 156 17456 196 17488
rect 228 17456 268 17488
rect 300 17456 340 17488
rect 372 17456 412 17488
rect 444 17456 484 17488
rect 516 17456 556 17488
rect 588 17456 628 17488
rect 660 17456 700 17488
rect 732 17456 772 17488
rect 804 17456 844 17488
rect 876 17456 950 17488
rect 50 17416 950 17456
rect 50 17384 124 17416
rect 156 17384 196 17416
rect 228 17384 268 17416
rect 300 17384 340 17416
rect 372 17384 412 17416
rect 444 17384 484 17416
rect 516 17384 556 17416
rect 588 17384 628 17416
rect 660 17384 700 17416
rect 732 17384 772 17416
rect 804 17384 844 17416
rect 876 17384 950 17416
rect 50 17344 950 17384
rect 50 17312 124 17344
rect 156 17312 196 17344
rect 228 17312 268 17344
rect 300 17312 340 17344
rect 372 17312 412 17344
rect 444 17312 484 17344
rect 516 17312 556 17344
rect 588 17312 628 17344
rect 660 17312 700 17344
rect 732 17312 772 17344
rect 804 17312 844 17344
rect 876 17312 950 17344
rect 50 17272 950 17312
rect 50 17240 124 17272
rect 156 17240 196 17272
rect 228 17240 268 17272
rect 300 17240 340 17272
rect 372 17240 412 17272
rect 444 17240 484 17272
rect 516 17240 556 17272
rect 588 17240 628 17272
rect 660 17240 700 17272
rect 732 17240 772 17272
rect 804 17240 844 17272
rect 876 17240 950 17272
rect 50 17200 950 17240
rect 50 17168 124 17200
rect 156 17168 196 17200
rect 228 17168 268 17200
rect 300 17168 340 17200
rect 372 17168 412 17200
rect 444 17168 484 17200
rect 516 17168 556 17200
rect 588 17168 628 17200
rect 660 17168 700 17200
rect 732 17168 772 17200
rect 804 17168 844 17200
rect 876 17168 950 17200
rect 50 17128 950 17168
rect 50 17096 124 17128
rect 156 17096 196 17128
rect 228 17096 268 17128
rect 300 17096 340 17128
rect 372 17096 412 17128
rect 444 17096 484 17128
rect 516 17096 556 17128
rect 588 17096 628 17128
rect 660 17096 700 17128
rect 732 17096 772 17128
rect 804 17096 844 17128
rect 876 17096 950 17128
rect 50 17056 950 17096
rect 50 17024 124 17056
rect 156 17024 196 17056
rect 228 17024 268 17056
rect 300 17024 340 17056
rect 372 17024 412 17056
rect 444 17024 484 17056
rect 516 17024 556 17056
rect 588 17024 628 17056
rect 660 17024 700 17056
rect 732 17024 772 17056
rect 804 17024 844 17056
rect 876 17024 950 17056
rect 50 16984 950 17024
rect 50 16952 124 16984
rect 156 16952 196 16984
rect 228 16952 268 16984
rect 300 16952 340 16984
rect 372 16952 412 16984
rect 444 16952 484 16984
rect 516 16952 556 16984
rect 588 16952 628 16984
rect 660 16952 700 16984
rect 732 16952 772 16984
rect 804 16952 844 16984
rect 876 16952 950 16984
rect 50 16912 950 16952
rect 50 16880 124 16912
rect 156 16880 196 16912
rect 228 16880 268 16912
rect 300 16880 340 16912
rect 372 16880 412 16912
rect 444 16880 484 16912
rect 516 16880 556 16912
rect 588 16880 628 16912
rect 660 16880 700 16912
rect 732 16880 772 16912
rect 804 16880 844 16912
rect 876 16880 950 16912
rect 50 16840 950 16880
rect 50 16808 124 16840
rect 156 16808 196 16840
rect 228 16808 268 16840
rect 300 16808 340 16840
rect 372 16808 412 16840
rect 444 16808 484 16840
rect 516 16808 556 16840
rect 588 16808 628 16840
rect 660 16808 700 16840
rect 732 16808 772 16840
rect 804 16808 844 16840
rect 876 16808 950 16840
rect 50 16768 950 16808
rect 50 16736 124 16768
rect 156 16736 196 16768
rect 228 16736 268 16768
rect 300 16736 340 16768
rect 372 16736 412 16768
rect 444 16736 484 16768
rect 516 16736 556 16768
rect 588 16736 628 16768
rect 660 16736 700 16768
rect 732 16736 772 16768
rect 804 16736 844 16768
rect 876 16736 950 16768
rect 50 16696 950 16736
rect 50 16664 124 16696
rect 156 16664 196 16696
rect 228 16664 268 16696
rect 300 16664 340 16696
rect 372 16664 412 16696
rect 444 16664 484 16696
rect 516 16664 556 16696
rect 588 16664 628 16696
rect 660 16664 700 16696
rect 732 16664 772 16696
rect 804 16664 844 16696
rect 876 16664 950 16696
rect 50 16624 950 16664
rect 50 16592 124 16624
rect 156 16592 196 16624
rect 228 16592 268 16624
rect 300 16592 340 16624
rect 372 16592 412 16624
rect 444 16592 484 16624
rect 516 16592 556 16624
rect 588 16592 628 16624
rect 660 16592 700 16624
rect 732 16592 772 16624
rect 804 16592 844 16624
rect 876 16592 950 16624
rect 50 16552 950 16592
rect 50 16520 124 16552
rect 156 16520 196 16552
rect 228 16520 268 16552
rect 300 16520 340 16552
rect 372 16520 412 16552
rect 444 16520 484 16552
rect 516 16520 556 16552
rect 588 16520 628 16552
rect 660 16520 700 16552
rect 732 16520 772 16552
rect 804 16520 844 16552
rect 876 16520 950 16552
rect 50 16480 950 16520
rect 50 16448 124 16480
rect 156 16448 196 16480
rect 228 16448 268 16480
rect 300 16448 340 16480
rect 372 16448 412 16480
rect 444 16448 484 16480
rect 516 16448 556 16480
rect 588 16448 628 16480
rect 660 16448 700 16480
rect 732 16448 772 16480
rect 804 16448 844 16480
rect 876 16448 950 16480
rect 50 16408 950 16448
rect 50 16376 124 16408
rect 156 16376 196 16408
rect 228 16376 268 16408
rect 300 16376 340 16408
rect 372 16376 412 16408
rect 444 16376 484 16408
rect 516 16376 556 16408
rect 588 16376 628 16408
rect 660 16376 700 16408
rect 732 16376 772 16408
rect 804 16376 844 16408
rect 876 16376 950 16408
rect 50 16336 950 16376
rect 50 16304 124 16336
rect 156 16304 196 16336
rect 228 16304 268 16336
rect 300 16304 340 16336
rect 372 16304 412 16336
rect 444 16304 484 16336
rect 516 16304 556 16336
rect 588 16304 628 16336
rect 660 16304 700 16336
rect 732 16304 772 16336
rect 804 16304 844 16336
rect 876 16304 950 16336
rect 50 16264 950 16304
rect 50 16232 124 16264
rect 156 16232 196 16264
rect 228 16232 268 16264
rect 300 16232 340 16264
rect 372 16232 412 16264
rect 444 16232 484 16264
rect 516 16232 556 16264
rect 588 16232 628 16264
rect 660 16232 700 16264
rect 732 16232 772 16264
rect 804 16232 844 16264
rect 876 16232 950 16264
rect 50 16192 950 16232
rect 50 16160 124 16192
rect 156 16160 196 16192
rect 228 16160 268 16192
rect 300 16160 340 16192
rect 372 16160 412 16192
rect 444 16160 484 16192
rect 516 16160 556 16192
rect 588 16160 628 16192
rect 660 16160 700 16192
rect 732 16160 772 16192
rect 804 16160 844 16192
rect 876 16160 950 16192
rect 50 16120 950 16160
rect 50 16088 124 16120
rect 156 16088 196 16120
rect 228 16088 268 16120
rect 300 16088 340 16120
rect 372 16088 412 16120
rect 444 16088 484 16120
rect 516 16088 556 16120
rect 588 16088 628 16120
rect 660 16088 700 16120
rect 732 16088 772 16120
rect 804 16088 844 16120
rect 876 16088 950 16120
rect 50 16048 950 16088
rect 50 16016 124 16048
rect 156 16016 196 16048
rect 228 16016 268 16048
rect 300 16016 340 16048
rect 372 16016 412 16048
rect 444 16016 484 16048
rect 516 16016 556 16048
rect 588 16016 628 16048
rect 660 16016 700 16048
rect 732 16016 772 16048
rect 804 16016 844 16048
rect 876 16016 950 16048
rect 50 15976 950 16016
rect 50 15944 124 15976
rect 156 15944 196 15976
rect 228 15944 268 15976
rect 300 15944 340 15976
rect 372 15944 412 15976
rect 444 15944 484 15976
rect 516 15944 556 15976
rect 588 15944 628 15976
rect 660 15944 700 15976
rect 732 15944 772 15976
rect 804 15944 844 15976
rect 876 15944 950 15976
rect 50 15904 950 15944
rect 50 15872 124 15904
rect 156 15872 196 15904
rect 228 15872 268 15904
rect 300 15872 340 15904
rect 372 15872 412 15904
rect 444 15872 484 15904
rect 516 15872 556 15904
rect 588 15872 628 15904
rect 660 15872 700 15904
rect 732 15872 772 15904
rect 804 15872 844 15904
rect 876 15872 950 15904
rect 50 15832 950 15872
rect 50 15800 124 15832
rect 156 15800 196 15832
rect 228 15800 268 15832
rect 300 15800 340 15832
rect 372 15800 412 15832
rect 444 15800 484 15832
rect 516 15800 556 15832
rect 588 15800 628 15832
rect 660 15800 700 15832
rect 732 15800 772 15832
rect 804 15800 844 15832
rect 876 15800 950 15832
rect 50 15760 950 15800
rect 50 15728 124 15760
rect 156 15728 196 15760
rect 228 15728 268 15760
rect 300 15728 340 15760
rect 372 15728 412 15760
rect 444 15728 484 15760
rect 516 15728 556 15760
rect 588 15728 628 15760
rect 660 15728 700 15760
rect 732 15728 772 15760
rect 804 15728 844 15760
rect 876 15728 950 15760
rect 50 15688 950 15728
rect 50 15656 124 15688
rect 156 15656 196 15688
rect 228 15656 268 15688
rect 300 15656 340 15688
rect 372 15656 412 15688
rect 444 15656 484 15688
rect 516 15656 556 15688
rect 588 15656 628 15688
rect 660 15656 700 15688
rect 732 15656 772 15688
rect 804 15656 844 15688
rect 876 15656 950 15688
rect 50 15616 950 15656
rect 50 15584 124 15616
rect 156 15584 196 15616
rect 228 15584 268 15616
rect 300 15584 340 15616
rect 372 15584 412 15616
rect 444 15584 484 15616
rect 516 15584 556 15616
rect 588 15584 628 15616
rect 660 15584 700 15616
rect 732 15584 772 15616
rect 804 15584 844 15616
rect 876 15584 950 15616
rect 50 15544 950 15584
rect 50 15512 124 15544
rect 156 15512 196 15544
rect 228 15512 268 15544
rect 300 15512 340 15544
rect 372 15512 412 15544
rect 444 15512 484 15544
rect 516 15512 556 15544
rect 588 15512 628 15544
rect 660 15512 700 15544
rect 732 15512 772 15544
rect 804 15512 844 15544
rect 876 15512 950 15544
rect 50 15472 950 15512
rect 50 15440 124 15472
rect 156 15440 196 15472
rect 228 15440 268 15472
rect 300 15440 340 15472
rect 372 15440 412 15472
rect 444 15440 484 15472
rect 516 15440 556 15472
rect 588 15440 628 15472
rect 660 15440 700 15472
rect 732 15440 772 15472
rect 804 15440 844 15472
rect 876 15440 950 15472
rect 50 15400 950 15440
rect 50 15368 124 15400
rect 156 15368 196 15400
rect 228 15368 268 15400
rect 300 15368 340 15400
rect 372 15368 412 15400
rect 444 15368 484 15400
rect 516 15368 556 15400
rect 588 15368 628 15400
rect 660 15368 700 15400
rect 732 15368 772 15400
rect 804 15368 844 15400
rect 876 15368 950 15400
rect 50 15328 950 15368
rect 50 15296 124 15328
rect 156 15296 196 15328
rect 228 15296 268 15328
rect 300 15296 340 15328
rect 372 15296 412 15328
rect 444 15296 484 15328
rect 516 15296 556 15328
rect 588 15296 628 15328
rect 660 15296 700 15328
rect 732 15296 772 15328
rect 804 15296 844 15328
rect 876 15296 950 15328
rect 50 15256 950 15296
rect 50 15224 124 15256
rect 156 15224 196 15256
rect 228 15224 268 15256
rect 300 15224 340 15256
rect 372 15224 412 15256
rect 444 15224 484 15256
rect 516 15224 556 15256
rect 588 15224 628 15256
rect 660 15224 700 15256
rect 732 15224 772 15256
rect 804 15224 844 15256
rect 876 15224 950 15256
rect 50 15184 950 15224
rect 50 15152 124 15184
rect 156 15152 196 15184
rect 228 15152 268 15184
rect 300 15152 340 15184
rect 372 15152 412 15184
rect 444 15152 484 15184
rect 516 15152 556 15184
rect 588 15152 628 15184
rect 660 15152 700 15184
rect 732 15152 772 15184
rect 804 15152 844 15184
rect 876 15152 950 15184
rect 50 15112 950 15152
rect 50 15080 124 15112
rect 156 15080 196 15112
rect 228 15080 268 15112
rect 300 15080 340 15112
rect 372 15080 412 15112
rect 444 15080 484 15112
rect 516 15080 556 15112
rect 588 15080 628 15112
rect 660 15080 700 15112
rect 732 15080 772 15112
rect 804 15080 844 15112
rect 876 15080 950 15112
rect 50 15040 950 15080
rect 50 15008 124 15040
rect 156 15008 196 15040
rect 228 15008 268 15040
rect 300 15008 340 15040
rect 372 15008 412 15040
rect 444 15008 484 15040
rect 516 15008 556 15040
rect 588 15008 628 15040
rect 660 15008 700 15040
rect 732 15008 772 15040
rect 804 15008 844 15040
rect 876 15008 950 15040
rect 50 14968 950 15008
rect 50 14936 124 14968
rect 156 14936 196 14968
rect 228 14936 268 14968
rect 300 14936 340 14968
rect 372 14936 412 14968
rect 444 14936 484 14968
rect 516 14936 556 14968
rect 588 14936 628 14968
rect 660 14936 700 14968
rect 732 14936 772 14968
rect 804 14936 844 14968
rect 876 14936 950 14968
rect 50 14896 950 14936
rect 50 14864 124 14896
rect 156 14864 196 14896
rect 228 14864 268 14896
rect 300 14864 340 14896
rect 372 14864 412 14896
rect 444 14864 484 14896
rect 516 14864 556 14896
rect 588 14864 628 14896
rect 660 14864 700 14896
rect 732 14864 772 14896
rect 804 14864 844 14896
rect 876 14864 950 14896
rect 50 14824 950 14864
rect 50 14792 124 14824
rect 156 14792 196 14824
rect 228 14792 268 14824
rect 300 14792 340 14824
rect 372 14792 412 14824
rect 444 14792 484 14824
rect 516 14792 556 14824
rect 588 14792 628 14824
rect 660 14792 700 14824
rect 732 14792 772 14824
rect 804 14792 844 14824
rect 876 14792 950 14824
rect 50 14752 950 14792
rect 50 14720 124 14752
rect 156 14720 196 14752
rect 228 14720 268 14752
rect 300 14720 340 14752
rect 372 14720 412 14752
rect 444 14720 484 14752
rect 516 14720 556 14752
rect 588 14720 628 14752
rect 660 14720 700 14752
rect 732 14720 772 14752
rect 804 14720 844 14752
rect 876 14720 950 14752
rect 50 14680 950 14720
rect 50 14648 124 14680
rect 156 14648 196 14680
rect 228 14648 268 14680
rect 300 14648 340 14680
rect 372 14648 412 14680
rect 444 14648 484 14680
rect 516 14648 556 14680
rect 588 14648 628 14680
rect 660 14648 700 14680
rect 732 14648 772 14680
rect 804 14648 844 14680
rect 876 14648 950 14680
rect 50 14608 950 14648
rect 50 14576 124 14608
rect 156 14576 196 14608
rect 228 14576 268 14608
rect 300 14576 340 14608
rect 372 14576 412 14608
rect 444 14576 484 14608
rect 516 14576 556 14608
rect 588 14576 628 14608
rect 660 14576 700 14608
rect 732 14576 772 14608
rect 804 14576 844 14608
rect 876 14576 950 14608
rect 50 14536 950 14576
rect 50 14504 124 14536
rect 156 14504 196 14536
rect 228 14504 268 14536
rect 300 14504 340 14536
rect 372 14504 412 14536
rect 444 14504 484 14536
rect 516 14504 556 14536
rect 588 14504 628 14536
rect 660 14504 700 14536
rect 732 14504 772 14536
rect 804 14504 844 14536
rect 876 14504 950 14536
rect 50 14464 950 14504
rect 50 14432 124 14464
rect 156 14432 196 14464
rect 228 14432 268 14464
rect 300 14432 340 14464
rect 372 14432 412 14464
rect 444 14432 484 14464
rect 516 14432 556 14464
rect 588 14432 628 14464
rect 660 14432 700 14464
rect 732 14432 772 14464
rect 804 14432 844 14464
rect 876 14432 950 14464
rect 50 14392 950 14432
rect 50 14360 124 14392
rect 156 14360 196 14392
rect 228 14360 268 14392
rect 300 14360 340 14392
rect 372 14360 412 14392
rect 444 14360 484 14392
rect 516 14360 556 14392
rect 588 14360 628 14392
rect 660 14360 700 14392
rect 732 14360 772 14392
rect 804 14360 844 14392
rect 876 14360 950 14392
rect 50 14320 950 14360
rect 50 14288 124 14320
rect 156 14288 196 14320
rect 228 14288 268 14320
rect 300 14288 340 14320
rect 372 14288 412 14320
rect 444 14288 484 14320
rect 516 14288 556 14320
rect 588 14288 628 14320
rect 660 14288 700 14320
rect 732 14288 772 14320
rect 804 14288 844 14320
rect 876 14288 950 14320
rect 50 14248 950 14288
rect 50 14216 124 14248
rect 156 14216 196 14248
rect 228 14216 268 14248
rect 300 14216 340 14248
rect 372 14216 412 14248
rect 444 14216 484 14248
rect 516 14216 556 14248
rect 588 14216 628 14248
rect 660 14216 700 14248
rect 732 14216 772 14248
rect 804 14216 844 14248
rect 876 14216 950 14248
rect 50 14176 950 14216
rect 50 14144 124 14176
rect 156 14144 196 14176
rect 228 14144 268 14176
rect 300 14144 340 14176
rect 372 14144 412 14176
rect 444 14144 484 14176
rect 516 14144 556 14176
rect 588 14144 628 14176
rect 660 14144 700 14176
rect 732 14144 772 14176
rect 804 14144 844 14176
rect 876 14144 950 14176
rect 50 14104 950 14144
rect 50 14072 124 14104
rect 156 14072 196 14104
rect 228 14072 268 14104
rect 300 14072 340 14104
rect 372 14072 412 14104
rect 444 14072 484 14104
rect 516 14072 556 14104
rect 588 14072 628 14104
rect 660 14072 700 14104
rect 732 14072 772 14104
rect 804 14072 844 14104
rect 876 14072 950 14104
rect 50 14032 950 14072
rect 50 14000 124 14032
rect 156 14000 196 14032
rect 228 14000 268 14032
rect 300 14000 340 14032
rect 372 14000 412 14032
rect 444 14000 484 14032
rect 516 14000 556 14032
rect 588 14000 628 14032
rect 660 14000 700 14032
rect 732 14000 772 14032
rect 804 14000 844 14032
rect 876 14000 950 14032
rect 50 13960 950 14000
rect 50 13928 124 13960
rect 156 13928 196 13960
rect 228 13928 268 13960
rect 300 13928 340 13960
rect 372 13928 412 13960
rect 444 13928 484 13960
rect 516 13928 556 13960
rect 588 13928 628 13960
rect 660 13928 700 13960
rect 732 13928 772 13960
rect 804 13928 844 13960
rect 876 13928 950 13960
rect 50 13888 950 13928
rect 50 13856 124 13888
rect 156 13856 196 13888
rect 228 13856 268 13888
rect 300 13856 340 13888
rect 372 13856 412 13888
rect 444 13856 484 13888
rect 516 13856 556 13888
rect 588 13856 628 13888
rect 660 13856 700 13888
rect 732 13856 772 13888
rect 804 13856 844 13888
rect 876 13856 950 13888
rect 50 13816 950 13856
rect 50 13784 124 13816
rect 156 13784 196 13816
rect 228 13784 268 13816
rect 300 13784 340 13816
rect 372 13784 412 13816
rect 444 13784 484 13816
rect 516 13784 556 13816
rect 588 13784 628 13816
rect 660 13784 700 13816
rect 732 13784 772 13816
rect 804 13784 844 13816
rect 876 13784 950 13816
rect 50 13744 950 13784
rect 50 13712 124 13744
rect 156 13712 196 13744
rect 228 13712 268 13744
rect 300 13712 340 13744
rect 372 13712 412 13744
rect 444 13712 484 13744
rect 516 13712 556 13744
rect 588 13712 628 13744
rect 660 13712 700 13744
rect 732 13712 772 13744
rect 804 13712 844 13744
rect 876 13712 950 13744
rect 50 13672 950 13712
rect 50 13640 124 13672
rect 156 13640 196 13672
rect 228 13640 268 13672
rect 300 13640 340 13672
rect 372 13640 412 13672
rect 444 13640 484 13672
rect 516 13640 556 13672
rect 588 13640 628 13672
rect 660 13640 700 13672
rect 732 13640 772 13672
rect 804 13640 844 13672
rect 876 13640 950 13672
rect 50 13600 950 13640
rect 50 13568 124 13600
rect 156 13568 196 13600
rect 228 13568 268 13600
rect 300 13568 340 13600
rect 372 13568 412 13600
rect 444 13568 484 13600
rect 516 13568 556 13600
rect 588 13568 628 13600
rect 660 13568 700 13600
rect 732 13568 772 13600
rect 804 13568 844 13600
rect 876 13568 950 13600
rect 50 13528 950 13568
rect 50 13496 124 13528
rect 156 13496 196 13528
rect 228 13496 268 13528
rect 300 13496 340 13528
rect 372 13496 412 13528
rect 444 13496 484 13528
rect 516 13496 556 13528
rect 588 13496 628 13528
rect 660 13496 700 13528
rect 732 13496 772 13528
rect 804 13496 844 13528
rect 876 13496 950 13528
rect 50 13456 950 13496
rect 50 13424 124 13456
rect 156 13424 196 13456
rect 228 13424 268 13456
rect 300 13424 340 13456
rect 372 13424 412 13456
rect 444 13424 484 13456
rect 516 13424 556 13456
rect 588 13424 628 13456
rect 660 13424 700 13456
rect 732 13424 772 13456
rect 804 13424 844 13456
rect 876 13424 950 13456
rect 50 13384 950 13424
rect 50 13352 124 13384
rect 156 13352 196 13384
rect 228 13352 268 13384
rect 300 13352 340 13384
rect 372 13352 412 13384
rect 444 13352 484 13384
rect 516 13352 556 13384
rect 588 13352 628 13384
rect 660 13352 700 13384
rect 732 13352 772 13384
rect 804 13352 844 13384
rect 876 13352 950 13384
rect 50 13312 950 13352
rect 50 13280 124 13312
rect 156 13280 196 13312
rect 228 13280 268 13312
rect 300 13280 340 13312
rect 372 13280 412 13312
rect 444 13280 484 13312
rect 516 13280 556 13312
rect 588 13280 628 13312
rect 660 13280 700 13312
rect 732 13280 772 13312
rect 804 13280 844 13312
rect 876 13280 950 13312
rect 50 13240 950 13280
rect 50 13208 124 13240
rect 156 13208 196 13240
rect 228 13208 268 13240
rect 300 13208 340 13240
rect 372 13208 412 13240
rect 444 13208 484 13240
rect 516 13208 556 13240
rect 588 13208 628 13240
rect 660 13208 700 13240
rect 732 13208 772 13240
rect 804 13208 844 13240
rect 876 13208 950 13240
rect 50 13168 950 13208
rect 50 13136 124 13168
rect 156 13136 196 13168
rect 228 13136 268 13168
rect 300 13136 340 13168
rect 372 13136 412 13168
rect 444 13136 484 13168
rect 516 13136 556 13168
rect 588 13136 628 13168
rect 660 13136 700 13168
rect 732 13136 772 13168
rect 804 13136 844 13168
rect 876 13136 950 13168
rect 50 13096 950 13136
rect 50 13064 124 13096
rect 156 13064 196 13096
rect 228 13064 268 13096
rect 300 13064 340 13096
rect 372 13064 412 13096
rect 444 13064 484 13096
rect 516 13064 556 13096
rect 588 13064 628 13096
rect 660 13064 700 13096
rect 732 13064 772 13096
rect 804 13064 844 13096
rect 876 13064 950 13096
rect 50 13000 950 13064
<< nsubdiff >>
rect 196 33384 228 33416
rect 268 33384 300 33416
rect 340 33384 372 33416
rect 412 33384 444 33416
rect 484 33384 516 33416
rect 556 33384 588 33416
rect 628 33384 660 33416
rect 700 33384 732 33416
rect 772 33384 804 33416
rect 844 33384 876 33416
rect 196 29684 228 29716
rect 268 29684 300 29716
rect 340 29684 372 29716
rect 412 29684 444 29716
rect 484 29684 516 29716
rect 556 29684 588 29716
rect 628 29684 660 29716
rect 700 29684 732 29716
rect 772 29684 804 29716
rect 844 29684 876 29716
rect 124 12112 156 12144
rect 196 12112 228 12144
rect 268 12112 300 12144
rect 340 12112 372 12144
rect 412 12112 444 12144
rect 484 12112 516 12144
rect 556 12112 588 12144
rect 628 12112 660 12144
rect 700 12112 732 12144
rect 772 12112 804 12144
rect 844 12112 876 12144
rect 916 12112 948 12144
rect 52 12040 84 12072
rect 124 12040 156 12072
rect 196 12040 228 12072
rect 268 12040 300 12072
rect 340 12040 372 12072
rect 412 12040 444 12072
rect 484 12040 516 12072
rect 556 12040 588 12072
rect 628 12040 660 12072
rect 700 12040 732 12072
rect 772 12040 804 12072
rect 844 12040 876 12072
rect 916 12040 948 12072
rect 52 11968 84 12000
rect 124 11968 156 12000
rect 196 11968 228 12000
rect 268 11968 300 12000
rect 340 11968 372 12000
rect 412 11968 444 12000
rect 484 11968 516 12000
rect 556 11968 588 12000
rect 628 11968 660 12000
rect 700 11968 732 12000
rect 772 11968 804 12000
rect 844 11968 876 12000
rect 916 11968 948 12000
rect 52 11896 84 11928
rect 124 11896 156 11928
rect 196 11896 228 11928
rect 268 11896 300 11928
rect 340 11896 372 11928
rect 412 11896 444 11928
rect 484 11896 516 11928
rect 556 11896 588 11928
rect 628 11896 660 11928
rect 700 11896 732 11928
rect 772 11896 804 11928
rect 844 11896 876 11928
rect 916 11896 948 11928
rect 52 11824 84 11856
rect 124 11824 156 11856
rect 196 11824 228 11856
rect 268 11824 300 11856
rect 340 11824 372 11856
rect 412 11824 444 11856
rect 484 11824 516 11856
rect 556 11824 588 11856
rect 628 11824 660 11856
rect 700 11824 732 11856
rect 772 11824 804 11856
rect 844 11824 876 11856
rect 916 11824 948 11856
rect 52 11752 84 11784
rect 124 11752 156 11784
rect 196 11752 228 11784
rect 268 11752 300 11784
rect 340 11752 372 11784
rect 412 11752 444 11784
rect 484 11752 516 11784
rect 556 11752 588 11784
rect 628 11752 660 11784
rect 700 11752 732 11784
rect 772 11752 804 11784
rect 844 11752 876 11784
rect 916 11752 948 11784
rect 52 11680 84 11712
rect 124 11680 156 11712
rect 196 11680 228 11712
rect 268 11680 300 11712
rect 340 11680 372 11712
rect 412 11680 444 11712
rect 484 11680 516 11712
rect 556 11680 588 11712
rect 628 11680 660 11712
rect 700 11680 732 11712
rect 772 11680 804 11712
rect 844 11680 876 11712
rect 916 11680 948 11712
rect 52 11608 84 11640
rect 124 11608 156 11640
rect 196 11608 228 11640
rect 268 11608 300 11640
rect 340 11608 372 11640
rect 412 11608 444 11640
rect 484 11608 516 11640
rect 556 11608 588 11640
rect 628 11608 660 11640
rect 700 11608 732 11640
rect 772 11608 804 11640
rect 844 11608 876 11640
rect 916 11608 948 11640
rect 52 11536 84 11568
rect 124 11536 156 11568
rect 196 11536 228 11568
rect 268 11536 300 11568
rect 340 11536 372 11568
rect 412 11536 444 11568
rect 484 11536 516 11568
rect 556 11536 588 11568
rect 628 11536 660 11568
rect 700 11536 732 11568
rect 772 11536 804 11568
rect 844 11536 876 11568
rect 916 11536 948 11568
rect 52 11464 84 11496
rect 124 11464 156 11496
rect 196 11464 228 11496
rect 268 11464 300 11496
rect 340 11464 372 11496
rect 412 11464 444 11496
rect 484 11464 516 11496
rect 556 11464 588 11496
rect 628 11464 660 11496
rect 700 11464 732 11496
rect 772 11464 804 11496
rect 844 11464 876 11496
rect 916 11464 948 11496
rect 52 11392 84 11424
rect 124 11392 156 11424
rect 196 11392 228 11424
rect 268 11392 300 11424
rect 340 11392 372 11424
rect 412 11392 444 11424
rect 484 11392 516 11424
rect 556 11392 588 11424
rect 628 11392 660 11424
rect 700 11392 732 11424
rect 772 11392 804 11424
rect 844 11392 876 11424
rect 916 11392 948 11424
rect 52 11320 84 11352
rect 124 11320 156 11352
rect 196 11320 228 11352
rect 268 11320 300 11352
rect 340 11320 372 11352
rect 412 11320 444 11352
rect 484 11320 516 11352
rect 556 11320 588 11352
rect 628 11320 660 11352
rect 700 11320 732 11352
rect 772 11320 804 11352
rect 844 11320 876 11352
rect 916 11320 948 11352
rect 52 11248 84 11280
rect 124 11248 156 11280
rect 196 11248 228 11280
rect 268 11248 300 11280
rect 340 11248 372 11280
rect 412 11248 444 11280
rect 484 11248 516 11280
rect 556 11248 588 11280
rect 628 11248 660 11280
rect 700 11248 732 11280
rect 772 11248 804 11280
rect 844 11248 876 11280
rect 916 11248 948 11280
rect 52 11176 84 11208
rect 124 11176 156 11208
rect 196 11176 228 11208
rect 268 11176 300 11208
rect 340 11176 372 11208
rect 412 11176 444 11208
rect 484 11176 516 11208
rect 556 11176 588 11208
rect 628 11176 660 11208
rect 700 11176 732 11208
rect 772 11176 804 11208
rect 844 11176 876 11208
rect 916 11176 948 11208
rect 52 11104 84 11136
rect 124 11104 156 11136
rect 196 11104 228 11136
rect 268 11104 300 11136
rect 340 11104 372 11136
rect 412 11104 444 11136
rect 484 11104 516 11136
rect 556 11104 588 11136
rect 628 11104 660 11136
rect 700 11104 732 11136
rect 772 11104 804 11136
rect 844 11104 876 11136
rect 916 11104 948 11136
rect 52 11032 84 11064
rect 124 11032 156 11064
rect 196 11032 228 11064
rect 268 11032 300 11064
rect 340 11032 372 11064
rect 412 11032 444 11064
rect 484 11032 516 11064
rect 556 11032 588 11064
rect 628 11032 660 11064
rect 700 11032 732 11064
rect 772 11032 804 11064
rect 844 11032 876 11064
rect 916 11032 948 11064
rect 52 10960 84 10992
rect 124 10960 156 10992
rect 196 10960 228 10992
rect 268 10960 300 10992
rect 340 10960 372 10992
rect 412 10960 444 10992
rect 484 10960 516 10992
rect 556 10960 588 10992
rect 628 10960 660 10992
rect 700 10960 732 10992
rect 772 10960 804 10992
rect 844 10960 876 10992
rect 916 10960 948 10992
rect 52 10888 84 10920
rect 124 10888 156 10920
rect 196 10888 228 10920
rect 268 10888 300 10920
rect 340 10888 372 10920
rect 412 10888 444 10920
rect 484 10888 516 10920
rect 556 10888 588 10920
rect 628 10888 660 10920
rect 700 10888 732 10920
rect 772 10888 804 10920
rect 844 10888 876 10920
rect 916 10888 948 10920
rect 52 10816 84 10848
rect 124 10816 156 10848
rect 196 10816 228 10848
rect 268 10816 300 10848
rect 340 10816 372 10848
rect 412 10816 444 10848
rect 484 10816 516 10848
rect 556 10816 588 10848
rect 628 10816 660 10848
rect 700 10816 732 10848
rect 772 10816 804 10848
rect 844 10816 876 10848
rect 916 10816 948 10848
rect 52 10744 84 10776
rect 124 10744 156 10776
rect 196 10744 228 10776
rect 268 10744 300 10776
rect 340 10744 372 10776
rect 412 10744 444 10776
rect 484 10744 516 10776
rect 556 10744 588 10776
rect 628 10744 660 10776
rect 700 10744 732 10776
rect 772 10744 804 10776
rect 844 10744 876 10776
rect 916 10744 948 10776
rect 52 10672 84 10704
rect 124 10672 156 10704
rect 196 10672 228 10704
rect 268 10672 300 10704
rect 340 10672 372 10704
rect 412 10672 444 10704
rect 484 10672 516 10704
rect 556 10672 588 10704
rect 628 10672 660 10704
rect 700 10672 732 10704
rect 772 10672 804 10704
rect 844 10672 876 10704
rect 916 10672 948 10704
rect 52 10600 84 10632
rect 124 10600 156 10632
rect 196 10600 228 10632
rect 268 10600 300 10632
rect 340 10600 372 10632
rect 412 10600 444 10632
rect 484 10600 516 10632
rect 556 10600 588 10632
rect 628 10600 660 10632
rect 700 10600 732 10632
rect 772 10600 804 10632
rect 844 10600 876 10632
rect 916 10600 948 10632
rect 52 10528 84 10560
rect 124 10528 156 10560
rect 196 10528 228 10560
rect 268 10528 300 10560
rect 340 10528 372 10560
rect 412 10528 444 10560
rect 484 10528 516 10560
rect 556 10528 588 10560
rect 628 10528 660 10560
rect 700 10528 732 10560
rect 772 10528 804 10560
rect 844 10528 876 10560
rect 916 10528 948 10560
rect 52 10456 84 10488
rect 124 10456 156 10488
rect 196 10456 228 10488
rect 268 10456 300 10488
rect 340 10456 372 10488
rect 412 10456 444 10488
rect 484 10456 516 10488
rect 556 10456 588 10488
rect 628 10456 660 10488
rect 700 10456 732 10488
rect 772 10456 804 10488
rect 844 10456 876 10488
rect 916 10456 948 10488
rect 52 10384 84 10416
rect 124 10384 156 10416
rect 196 10384 228 10416
rect 268 10384 300 10416
rect 340 10384 372 10416
rect 412 10384 444 10416
rect 484 10384 516 10416
rect 556 10384 588 10416
rect 628 10384 660 10416
rect 700 10384 732 10416
rect 772 10384 804 10416
rect 844 10384 876 10416
rect 916 10384 948 10416
rect 52 10312 84 10344
rect 124 10312 156 10344
rect 196 10312 228 10344
rect 268 10312 300 10344
rect 340 10312 372 10344
rect 412 10312 444 10344
rect 484 10312 516 10344
rect 556 10312 588 10344
rect 628 10312 660 10344
rect 700 10312 732 10344
rect 772 10312 804 10344
rect 844 10312 876 10344
rect 916 10312 948 10344
rect 52 10240 84 10272
rect 124 10240 156 10272
rect 196 10240 228 10272
rect 268 10240 300 10272
rect 340 10240 372 10272
rect 412 10240 444 10272
rect 484 10240 516 10272
rect 556 10240 588 10272
rect 628 10240 660 10272
rect 700 10240 732 10272
rect 772 10240 804 10272
rect 844 10240 876 10272
rect 916 10240 948 10272
rect 52 10168 84 10200
rect 124 10168 156 10200
rect 196 10168 228 10200
rect 268 10168 300 10200
rect 340 10168 372 10200
rect 412 10168 444 10200
rect 484 10168 516 10200
rect 556 10168 588 10200
rect 628 10168 660 10200
rect 700 10168 732 10200
rect 772 10168 804 10200
rect 844 10168 876 10200
rect 916 10168 948 10200
rect 52 10096 84 10128
rect 124 10096 156 10128
rect 196 10096 228 10128
rect 268 10096 300 10128
rect 340 10096 372 10128
rect 412 10096 444 10128
rect 484 10096 516 10128
rect 556 10096 588 10128
rect 628 10096 660 10128
rect 700 10096 732 10128
rect 772 10096 804 10128
rect 844 10096 876 10128
rect 916 10096 948 10128
rect 52 10024 84 10056
rect 124 10024 156 10056
rect 196 10024 228 10056
rect 268 10024 300 10056
rect 340 10024 372 10056
rect 412 10024 444 10056
rect 484 10024 516 10056
rect 556 10024 588 10056
rect 628 10024 660 10056
rect 700 10024 732 10056
rect 772 10024 804 10056
rect 844 10024 876 10056
rect 916 10024 948 10056
rect 52 9952 84 9984
rect 124 9952 156 9984
rect 196 9952 228 9984
rect 268 9952 300 9984
rect 340 9952 372 9984
rect 412 9952 444 9984
rect 484 9952 516 9984
rect 556 9952 588 9984
rect 628 9952 660 9984
rect 700 9952 732 9984
rect 772 9952 804 9984
rect 844 9952 876 9984
rect 916 9952 948 9984
rect 52 9880 84 9912
rect 124 9880 156 9912
rect 196 9880 228 9912
rect 268 9880 300 9912
rect 340 9880 372 9912
rect 412 9880 444 9912
rect 484 9880 516 9912
rect 556 9880 588 9912
rect 628 9880 660 9912
rect 700 9880 732 9912
rect 772 9880 804 9912
rect 844 9880 876 9912
rect 916 9880 948 9912
rect 52 9808 84 9840
rect 124 9808 156 9840
rect 196 9808 228 9840
rect 268 9808 300 9840
rect 340 9808 372 9840
rect 412 9808 444 9840
rect 484 9808 516 9840
rect 556 9808 588 9840
rect 628 9808 660 9840
rect 700 9808 732 9840
rect 772 9808 804 9840
rect 844 9808 876 9840
rect 916 9808 948 9840
rect 52 9736 84 9768
rect 124 9736 156 9768
rect 196 9736 228 9768
rect 268 9736 300 9768
rect 340 9736 372 9768
rect 412 9736 444 9768
rect 484 9736 516 9768
rect 556 9736 588 9768
rect 628 9736 660 9768
rect 700 9736 732 9768
rect 772 9736 804 9768
rect 844 9736 876 9768
rect 916 9736 948 9768
rect 52 9664 84 9696
rect 124 9664 156 9696
rect 196 9664 228 9696
rect 268 9664 300 9696
rect 340 9664 372 9696
rect 412 9664 444 9696
rect 484 9664 516 9696
rect 556 9664 588 9696
rect 628 9664 660 9696
rect 700 9664 732 9696
rect 772 9664 804 9696
rect 844 9664 876 9696
rect 916 9664 948 9696
rect 52 9592 84 9624
rect 124 9592 156 9624
rect 196 9592 228 9624
rect 268 9592 300 9624
rect 340 9592 372 9624
rect 412 9592 444 9624
rect 484 9592 516 9624
rect 556 9592 588 9624
rect 628 9592 660 9624
rect 700 9592 732 9624
rect 772 9592 804 9624
rect 844 9592 876 9624
rect 916 9592 948 9624
rect 52 9520 84 9552
rect 124 9520 156 9552
rect 196 9520 228 9552
rect 268 9520 300 9552
rect 340 9520 372 9552
rect 412 9520 444 9552
rect 484 9520 516 9552
rect 556 9520 588 9552
rect 628 9520 660 9552
rect 700 9520 732 9552
rect 772 9520 804 9552
rect 844 9520 876 9552
rect 916 9520 948 9552
rect 52 9448 84 9480
rect 124 9448 156 9480
rect 196 9448 228 9480
rect 268 9448 300 9480
rect 340 9448 372 9480
rect 412 9448 444 9480
rect 484 9448 516 9480
rect 556 9448 588 9480
rect 628 9448 660 9480
rect 700 9448 732 9480
rect 772 9448 804 9480
rect 844 9448 876 9480
rect 916 9448 948 9480
rect 52 9376 84 9408
rect 124 9376 156 9408
rect 196 9376 228 9408
rect 268 9376 300 9408
rect 340 9376 372 9408
rect 412 9376 444 9408
rect 484 9376 516 9408
rect 556 9376 588 9408
rect 628 9376 660 9408
rect 700 9376 732 9408
rect 772 9376 804 9408
rect 844 9376 876 9408
rect 916 9376 948 9408
rect 52 9304 84 9336
rect 124 9304 156 9336
rect 196 9304 228 9336
rect 268 9304 300 9336
rect 340 9304 372 9336
rect 412 9304 444 9336
rect 484 9304 516 9336
rect 556 9304 588 9336
rect 628 9304 660 9336
rect 700 9304 732 9336
rect 772 9304 804 9336
rect 844 9304 876 9336
rect 916 9304 948 9336
rect 52 9232 84 9264
rect 124 9232 156 9264
rect 196 9232 228 9264
rect 268 9232 300 9264
rect 340 9232 372 9264
rect 412 9232 444 9264
rect 484 9232 516 9264
rect 556 9232 588 9264
rect 628 9232 660 9264
rect 700 9232 732 9264
rect 772 9232 804 9264
rect 844 9232 876 9264
rect 916 9232 948 9264
rect 52 9160 84 9192
rect 124 9160 156 9192
rect 196 9160 228 9192
rect 268 9160 300 9192
rect 340 9160 372 9192
rect 412 9160 444 9192
rect 484 9160 516 9192
rect 556 9160 588 9192
rect 628 9160 660 9192
rect 700 9160 732 9192
rect 772 9160 804 9192
rect 844 9160 876 9192
rect 916 9160 948 9192
rect 52 9088 84 9120
rect 124 9088 156 9120
rect 196 9088 228 9120
rect 268 9088 300 9120
rect 340 9088 372 9120
rect 412 9088 444 9120
rect 484 9088 516 9120
rect 556 9088 588 9120
rect 628 9088 660 9120
rect 700 9088 732 9120
rect 772 9088 804 9120
rect 844 9088 876 9120
rect 916 9088 948 9120
rect 52 9016 84 9048
rect 124 9016 156 9048
rect 196 9016 228 9048
rect 268 9016 300 9048
rect 340 9016 372 9048
rect 412 9016 444 9048
rect 484 9016 516 9048
rect 556 9016 588 9048
rect 628 9016 660 9048
rect 700 9016 732 9048
rect 772 9016 804 9048
rect 844 9016 876 9048
rect 916 9016 948 9048
rect 52 8944 84 8976
rect 124 8944 156 8976
rect 196 8944 228 8976
rect 268 8944 300 8976
rect 340 8944 372 8976
rect 412 8944 444 8976
rect 484 8944 516 8976
rect 556 8944 588 8976
rect 628 8944 660 8976
rect 700 8944 732 8976
rect 772 8944 804 8976
rect 844 8944 876 8976
rect 916 8944 948 8976
rect 52 8872 84 8904
rect 124 8872 156 8904
rect 196 8872 228 8904
rect 268 8872 300 8904
rect 340 8872 372 8904
rect 412 8872 444 8904
rect 484 8872 516 8904
rect 556 8872 588 8904
rect 628 8872 660 8904
rect 700 8872 732 8904
rect 772 8872 804 8904
rect 844 8872 876 8904
rect 916 8872 948 8904
rect 52 8800 84 8832
rect 124 8800 156 8832
rect 196 8800 228 8832
rect 268 8800 300 8832
rect 340 8800 372 8832
rect 412 8800 444 8832
rect 484 8800 516 8832
rect 556 8800 588 8832
rect 628 8800 660 8832
rect 700 8800 732 8832
rect 772 8800 804 8832
rect 844 8800 876 8832
rect 916 8800 948 8832
rect 52 8728 84 8760
rect 124 8728 156 8760
rect 196 8728 228 8760
rect 268 8728 300 8760
rect 340 8728 372 8760
rect 412 8728 444 8760
rect 484 8728 516 8760
rect 556 8728 588 8760
rect 628 8728 660 8760
rect 700 8728 732 8760
rect 772 8728 804 8760
rect 844 8728 876 8760
rect 916 8728 948 8760
rect 52 8656 84 8688
rect 124 8656 156 8688
rect 196 8656 228 8688
rect 268 8656 300 8688
rect 340 8656 372 8688
rect 412 8656 444 8688
rect 484 8656 516 8688
rect 556 8656 588 8688
rect 628 8656 660 8688
rect 700 8656 732 8688
rect 772 8656 804 8688
rect 844 8656 876 8688
rect 916 8656 948 8688
rect 52 8584 84 8616
rect 124 8584 156 8616
rect 196 8584 228 8616
rect 268 8584 300 8616
rect 340 8584 372 8616
rect 412 8584 444 8616
rect 484 8584 516 8616
rect 556 8584 588 8616
rect 628 8584 660 8616
rect 700 8584 732 8616
rect 772 8584 804 8616
rect 844 8584 876 8616
rect 916 8584 948 8616
rect 52 8512 84 8544
rect 124 8512 156 8544
rect 196 8512 228 8544
rect 268 8512 300 8544
rect 340 8512 372 8544
rect 412 8512 444 8544
rect 484 8512 516 8544
rect 556 8512 588 8544
rect 628 8512 660 8544
rect 700 8512 732 8544
rect 772 8512 804 8544
rect 844 8512 876 8544
rect 916 8512 948 8544
rect 52 8440 84 8472
rect 124 8440 156 8472
rect 196 8440 228 8472
rect 268 8440 300 8472
rect 340 8440 372 8472
rect 412 8440 444 8472
rect 484 8440 516 8472
rect 556 8440 588 8472
rect 628 8440 660 8472
rect 700 8440 732 8472
rect 772 8440 804 8472
rect 844 8440 876 8472
rect 916 8440 948 8472
rect 52 8368 84 8400
rect 124 8368 156 8400
rect 196 8368 228 8400
rect 268 8368 300 8400
rect 340 8368 372 8400
rect 412 8368 444 8400
rect 484 8368 516 8400
rect 556 8368 588 8400
rect 628 8368 660 8400
rect 700 8368 732 8400
rect 772 8368 804 8400
rect 844 8368 876 8400
rect 916 8368 948 8400
rect 52 8296 84 8328
rect 124 8296 156 8328
rect 196 8296 228 8328
rect 268 8296 300 8328
rect 340 8296 372 8328
rect 412 8296 444 8328
rect 484 8296 516 8328
rect 556 8296 588 8328
rect 628 8296 660 8328
rect 700 8296 732 8328
rect 772 8296 804 8328
rect 844 8296 876 8328
rect 916 8296 948 8328
rect 52 8224 84 8256
rect 124 8224 156 8256
rect 196 8224 228 8256
rect 268 8224 300 8256
rect 340 8224 372 8256
rect 412 8224 444 8256
rect 484 8224 516 8256
rect 556 8224 588 8256
rect 628 8224 660 8256
rect 700 8224 732 8256
rect 772 8224 804 8256
rect 844 8224 876 8256
rect 916 8224 948 8256
rect 52 8152 84 8184
rect 124 8152 156 8184
rect 196 8152 228 8184
rect 268 8152 300 8184
rect 340 8152 372 8184
rect 412 8152 444 8184
rect 484 8152 516 8184
rect 556 8152 588 8184
rect 628 8152 660 8184
rect 700 8152 732 8184
rect 772 8152 804 8184
rect 844 8152 876 8184
rect 916 8152 948 8184
rect 52 8080 84 8112
rect 124 8080 156 8112
rect 196 8080 228 8112
rect 268 8080 300 8112
rect 340 8080 372 8112
rect 412 8080 444 8112
rect 484 8080 516 8112
rect 556 8080 588 8112
rect 628 8080 660 8112
rect 700 8080 732 8112
rect 772 8080 804 8112
rect 844 8080 876 8112
rect 916 8080 948 8112
rect 52 8008 84 8040
rect 124 8008 156 8040
rect 196 8008 228 8040
rect 268 8008 300 8040
rect 340 8008 372 8040
rect 412 8008 444 8040
rect 484 8008 516 8040
rect 556 8008 588 8040
rect 628 8008 660 8040
rect 700 8008 732 8040
rect 772 8008 804 8040
rect 844 8008 876 8040
rect 916 8008 948 8040
rect 52 7936 84 7968
rect 124 7936 156 7968
rect 196 7936 228 7968
rect 268 7936 300 7968
rect 340 7936 372 7968
rect 412 7936 444 7968
rect 484 7936 516 7968
rect 556 7936 588 7968
rect 628 7936 660 7968
rect 700 7936 732 7968
rect 772 7936 804 7968
rect 844 7936 876 7968
rect 916 7936 948 7968
rect 52 7864 84 7896
rect 124 7864 156 7896
rect 196 7864 228 7896
rect 268 7864 300 7896
rect 340 7864 372 7896
rect 412 7864 444 7896
rect 484 7864 516 7896
rect 556 7864 588 7896
rect 628 7864 660 7896
rect 700 7864 732 7896
rect 772 7864 804 7896
rect 844 7864 876 7896
rect 916 7864 948 7896
rect 52 7792 84 7824
rect 124 7792 156 7824
rect 196 7792 228 7824
rect 268 7792 300 7824
rect 340 7792 372 7824
rect 412 7792 444 7824
rect 484 7792 516 7824
rect 556 7792 588 7824
rect 628 7792 660 7824
rect 700 7792 732 7824
rect 772 7792 804 7824
rect 844 7792 876 7824
rect 916 7792 948 7824
rect 52 7720 84 7752
rect 124 7720 156 7752
rect 196 7720 228 7752
rect 268 7720 300 7752
rect 340 7720 372 7752
rect 412 7720 444 7752
rect 484 7720 516 7752
rect 556 7720 588 7752
rect 628 7720 660 7752
rect 700 7720 732 7752
rect 772 7720 804 7752
rect 844 7720 876 7752
rect 916 7720 948 7752
rect 52 7648 84 7680
rect 124 7648 156 7680
rect 196 7648 228 7680
rect 268 7648 300 7680
rect 340 7648 372 7680
rect 412 7648 444 7680
rect 484 7648 516 7680
rect 556 7648 588 7680
rect 628 7648 660 7680
rect 700 7648 732 7680
rect 772 7648 804 7680
rect 844 7648 876 7680
rect 916 7648 948 7680
rect 52 7576 84 7608
rect 124 7576 156 7608
rect 196 7576 228 7608
rect 268 7576 300 7608
rect 340 7576 372 7608
rect 412 7576 444 7608
rect 484 7576 516 7608
rect 556 7576 588 7608
rect 628 7576 660 7608
rect 700 7576 732 7608
rect 772 7576 804 7608
rect 844 7576 876 7608
rect 916 7576 948 7608
rect 52 7504 84 7536
rect 124 7504 156 7536
rect 196 7504 228 7536
rect 268 7504 300 7536
rect 340 7504 372 7536
rect 412 7504 444 7536
rect 484 7504 516 7536
rect 556 7504 588 7536
rect 628 7504 660 7536
rect 700 7504 732 7536
rect 772 7504 804 7536
rect 844 7504 876 7536
rect 916 7504 948 7536
rect 52 7432 84 7464
rect 124 7432 156 7464
rect 196 7432 228 7464
rect 268 7432 300 7464
rect 340 7432 372 7464
rect 412 7432 444 7464
rect 484 7432 516 7464
rect 556 7432 588 7464
rect 628 7432 660 7464
rect 700 7432 732 7464
rect 772 7432 804 7464
rect 844 7432 876 7464
rect 916 7432 948 7464
rect 52 7360 84 7392
rect 124 7360 156 7392
rect 196 7360 228 7392
rect 268 7360 300 7392
rect 340 7360 372 7392
rect 412 7360 444 7392
rect 484 7360 516 7392
rect 556 7360 588 7392
rect 628 7360 660 7392
rect 700 7360 732 7392
rect 772 7360 804 7392
rect 844 7360 876 7392
rect 916 7360 948 7392
rect 52 7288 84 7320
rect 124 7288 156 7320
rect 196 7288 228 7320
rect 268 7288 300 7320
rect 340 7288 372 7320
rect 412 7288 444 7320
rect 484 7288 516 7320
rect 556 7288 588 7320
rect 628 7288 660 7320
rect 700 7288 732 7320
rect 772 7288 804 7320
rect 844 7288 876 7320
rect 916 7288 948 7320
rect 52 7216 84 7248
rect 124 7216 156 7248
rect 196 7216 228 7248
rect 268 7216 300 7248
rect 340 7216 372 7248
rect 412 7216 444 7248
rect 484 7216 516 7248
rect 556 7216 588 7248
rect 628 7216 660 7248
rect 700 7216 732 7248
rect 772 7216 804 7248
rect 844 7216 876 7248
rect 916 7216 948 7248
rect 52 7144 84 7176
rect 124 7144 156 7176
rect 196 7144 228 7176
rect 268 7144 300 7176
rect 340 7144 372 7176
rect 412 7144 444 7176
rect 484 7144 516 7176
rect 556 7144 588 7176
rect 628 7144 660 7176
rect 700 7144 732 7176
rect 772 7144 804 7176
rect 844 7144 876 7176
rect 916 7144 948 7176
rect 52 7072 84 7104
rect 124 7072 156 7104
rect 196 7072 228 7104
rect 268 7072 300 7104
rect 340 7072 372 7104
rect 412 7072 444 7104
rect 484 7072 516 7104
rect 556 7072 588 7104
rect 628 7072 660 7104
rect 700 7072 732 7104
rect 772 7072 804 7104
rect 844 7072 876 7104
rect 916 7072 948 7104
rect 52 7000 84 7032
rect 124 7000 156 7032
rect 196 7000 228 7032
rect 268 7000 300 7032
rect 340 7000 372 7032
rect 412 7000 444 7032
rect 484 7000 516 7032
rect 556 7000 588 7032
rect 628 7000 660 7032
rect 700 7000 732 7032
rect 772 7000 804 7032
rect 844 7000 876 7032
rect 916 7000 948 7032
rect 52 6928 84 6960
rect 124 6928 156 6960
rect 196 6928 228 6960
rect 268 6928 300 6960
rect 340 6928 372 6960
rect 412 6928 444 6960
rect 484 6928 516 6960
rect 556 6928 588 6960
rect 628 6928 660 6960
rect 700 6928 732 6960
rect 772 6928 804 6960
rect 844 6928 876 6960
rect 916 6928 948 6960
rect 52 6856 84 6888
rect 124 6856 156 6888
rect 196 6856 228 6888
rect 268 6856 300 6888
rect 340 6856 372 6888
rect 412 6856 444 6888
rect 484 6856 516 6888
rect 556 6856 588 6888
rect 628 6856 660 6888
rect 700 6856 732 6888
rect 772 6856 804 6888
rect 844 6856 876 6888
rect 916 6856 948 6888
rect 124 6512 156 6544
rect 196 6512 228 6544
rect 268 6512 300 6544
rect 340 6512 372 6544
rect 412 6512 444 6544
rect 484 6512 516 6544
rect 556 6512 588 6544
rect 628 6512 660 6544
rect 700 6512 732 6544
rect 772 6512 804 6544
rect 844 6512 876 6544
rect 916 6512 948 6544
rect 52 6440 84 6472
rect 124 6440 156 6472
rect 196 6440 228 6472
rect 268 6440 300 6472
rect 340 6440 372 6472
rect 412 6440 444 6472
rect 484 6440 516 6472
rect 556 6440 588 6472
rect 628 6440 660 6472
rect 700 6440 732 6472
rect 772 6440 804 6472
rect 844 6440 876 6472
rect 916 6440 948 6472
rect 52 6368 84 6400
rect 124 6368 156 6400
rect 196 6368 228 6400
rect 268 6368 300 6400
rect 340 6368 372 6400
rect 412 6368 444 6400
rect 484 6368 516 6400
rect 556 6368 588 6400
rect 628 6368 660 6400
rect 700 6368 732 6400
rect 772 6368 804 6400
rect 844 6368 876 6400
rect 916 6368 948 6400
rect 52 6296 84 6328
rect 124 6296 156 6328
rect 196 6296 228 6328
rect 268 6296 300 6328
rect 340 6296 372 6328
rect 412 6296 444 6328
rect 484 6296 516 6328
rect 556 6296 588 6328
rect 628 6296 660 6328
rect 700 6296 732 6328
rect 772 6296 804 6328
rect 844 6296 876 6328
rect 916 6296 948 6328
rect 52 6224 84 6256
rect 124 6224 156 6256
rect 196 6224 228 6256
rect 268 6224 300 6256
rect 340 6224 372 6256
rect 412 6224 444 6256
rect 484 6224 516 6256
rect 556 6224 588 6256
rect 628 6224 660 6256
rect 700 6224 732 6256
rect 772 6224 804 6256
rect 844 6224 876 6256
rect 916 6224 948 6256
rect 52 6152 84 6184
rect 124 6152 156 6184
rect 196 6152 228 6184
rect 268 6152 300 6184
rect 340 6152 372 6184
rect 412 6152 444 6184
rect 484 6152 516 6184
rect 556 6152 588 6184
rect 628 6152 660 6184
rect 700 6152 732 6184
rect 772 6152 804 6184
rect 844 6152 876 6184
rect 916 6152 948 6184
rect 52 6080 84 6112
rect 124 6080 156 6112
rect 196 6080 228 6112
rect 268 6080 300 6112
rect 340 6080 372 6112
rect 412 6080 444 6112
rect 484 6080 516 6112
rect 556 6080 588 6112
rect 628 6080 660 6112
rect 700 6080 732 6112
rect 772 6080 804 6112
rect 844 6080 876 6112
rect 916 6080 948 6112
rect 52 6008 84 6040
rect 124 6008 156 6040
rect 196 6008 228 6040
rect 268 6008 300 6040
rect 340 6008 372 6040
rect 412 6008 444 6040
rect 484 6008 516 6040
rect 556 6008 588 6040
rect 628 6008 660 6040
rect 700 6008 732 6040
rect 772 6008 804 6040
rect 844 6008 876 6040
rect 916 6008 948 6040
rect 52 5936 84 5968
rect 124 5936 156 5968
rect 196 5936 228 5968
rect 268 5936 300 5968
rect 340 5936 372 5968
rect 412 5936 444 5968
rect 484 5936 516 5968
rect 556 5936 588 5968
rect 628 5936 660 5968
rect 700 5936 732 5968
rect 772 5936 804 5968
rect 844 5936 876 5968
rect 916 5936 948 5968
rect 52 5864 84 5896
rect 124 5864 156 5896
rect 196 5864 228 5896
rect 268 5864 300 5896
rect 340 5864 372 5896
rect 412 5864 444 5896
rect 484 5864 516 5896
rect 556 5864 588 5896
rect 628 5864 660 5896
rect 700 5864 732 5896
rect 772 5864 804 5896
rect 844 5864 876 5896
rect 916 5864 948 5896
rect 52 5792 84 5824
rect 124 5792 156 5824
rect 196 5792 228 5824
rect 268 5792 300 5824
rect 340 5792 372 5824
rect 412 5792 444 5824
rect 484 5792 516 5824
rect 556 5792 588 5824
rect 628 5792 660 5824
rect 700 5792 732 5824
rect 772 5792 804 5824
rect 844 5792 876 5824
rect 916 5792 948 5824
rect 52 5720 84 5752
rect 124 5720 156 5752
rect 196 5720 228 5752
rect 268 5720 300 5752
rect 340 5720 372 5752
rect 412 5720 444 5752
rect 484 5720 516 5752
rect 556 5720 588 5752
rect 628 5720 660 5752
rect 700 5720 732 5752
rect 772 5720 804 5752
rect 844 5720 876 5752
rect 916 5720 948 5752
rect 52 5648 84 5680
rect 124 5648 156 5680
rect 196 5648 228 5680
rect 268 5648 300 5680
rect 340 5648 372 5680
rect 412 5648 444 5680
rect 484 5648 516 5680
rect 556 5648 588 5680
rect 628 5648 660 5680
rect 700 5648 732 5680
rect 772 5648 804 5680
rect 844 5648 876 5680
rect 916 5648 948 5680
rect 52 5576 84 5608
rect 124 5576 156 5608
rect 196 5576 228 5608
rect 268 5576 300 5608
rect 340 5576 372 5608
rect 412 5576 444 5608
rect 484 5576 516 5608
rect 556 5576 588 5608
rect 628 5576 660 5608
rect 700 5576 732 5608
rect 772 5576 804 5608
rect 844 5576 876 5608
rect 916 5576 948 5608
rect 52 5504 84 5536
rect 124 5504 156 5536
rect 196 5504 228 5536
rect 268 5504 300 5536
rect 340 5504 372 5536
rect 412 5504 444 5536
rect 484 5504 516 5536
rect 556 5504 588 5536
rect 628 5504 660 5536
rect 700 5504 732 5536
rect 772 5504 804 5536
rect 844 5504 876 5536
rect 916 5504 948 5536
rect 52 5432 84 5464
rect 124 5432 156 5464
rect 196 5432 228 5464
rect 268 5432 300 5464
rect 340 5432 372 5464
rect 412 5432 444 5464
rect 484 5432 516 5464
rect 556 5432 588 5464
rect 628 5432 660 5464
rect 700 5432 732 5464
rect 772 5432 804 5464
rect 844 5432 876 5464
rect 916 5432 948 5464
rect 52 5360 84 5392
rect 124 5360 156 5392
rect 196 5360 228 5392
rect 268 5360 300 5392
rect 340 5360 372 5392
rect 412 5360 444 5392
rect 484 5360 516 5392
rect 556 5360 588 5392
rect 628 5360 660 5392
rect 700 5360 732 5392
rect 772 5360 804 5392
rect 844 5360 876 5392
rect 916 5360 948 5392
rect 52 5288 84 5320
rect 124 5288 156 5320
rect 196 5288 228 5320
rect 268 5288 300 5320
rect 340 5288 372 5320
rect 412 5288 444 5320
rect 484 5288 516 5320
rect 556 5288 588 5320
rect 628 5288 660 5320
rect 700 5288 732 5320
rect 772 5288 804 5320
rect 844 5288 876 5320
rect 916 5288 948 5320
rect 52 5216 84 5248
rect 124 5216 156 5248
rect 196 5216 228 5248
rect 268 5216 300 5248
rect 340 5216 372 5248
rect 412 5216 444 5248
rect 484 5216 516 5248
rect 556 5216 588 5248
rect 628 5216 660 5248
rect 700 5216 732 5248
rect 772 5216 804 5248
rect 844 5216 876 5248
rect 916 5216 948 5248
rect 52 5144 84 5176
rect 124 5144 156 5176
rect 196 5144 228 5176
rect 268 5144 300 5176
rect 340 5144 372 5176
rect 412 5144 444 5176
rect 484 5144 516 5176
rect 556 5144 588 5176
rect 628 5144 660 5176
rect 700 5144 732 5176
rect 772 5144 804 5176
rect 844 5144 876 5176
rect 916 5144 948 5176
rect 52 5072 84 5104
rect 124 5072 156 5104
rect 196 5072 228 5104
rect 268 5072 300 5104
rect 340 5072 372 5104
rect 412 5072 444 5104
rect 484 5072 516 5104
rect 556 5072 588 5104
rect 628 5072 660 5104
rect 700 5072 732 5104
rect 772 5072 804 5104
rect 844 5072 876 5104
rect 916 5072 948 5104
rect 52 5000 84 5032
rect 124 5000 156 5032
rect 196 5000 228 5032
rect 268 5000 300 5032
rect 340 5000 372 5032
rect 412 5000 444 5032
rect 484 5000 516 5032
rect 556 5000 588 5032
rect 628 5000 660 5032
rect 700 5000 732 5032
rect 772 5000 804 5032
rect 844 5000 876 5032
rect 916 5000 948 5032
rect 52 4928 84 4960
rect 124 4928 156 4960
rect 196 4928 228 4960
rect 268 4928 300 4960
rect 340 4928 372 4960
rect 412 4928 444 4960
rect 484 4928 516 4960
rect 556 4928 588 4960
rect 628 4928 660 4960
rect 700 4928 732 4960
rect 772 4928 804 4960
rect 844 4928 876 4960
rect 916 4928 948 4960
rect 52 4856 84 4888
rect 124 4856 156 4888
rect 196 4856 228 4888
rect 268 4856 300 4888
rect 340 4856 372 4888
rect 412 4856 444 4888
rect 484 4856 516 4888
rect 556 4856 588 4888
rect 628 4856 660 4888
rect 700 4856 732 4888
rect 772 4856 804 4888
rect 844 4856 876 4888
rect 916 4856 948 4888
rect 52 4784 84 4816
rect 124 4784 156 4816
rect 196 4784 228 4816
rect 268 4784 300 4816
rect 340 4784 372 4816
rect 412 4784 444 4816
rect 484 4784 516 4816
rect 556 4784 588 4816
rect 628 4784 660 4816
rect 700 4784 732 4816
rect 772 4784 804 4816
rect 844 4784 876 4816
rect 916 4784 948 4816
rect 52 4712 84 4744
rect 124 4712 156 4744
rect 196 4712 228 4744
rect 268 4712 300 4744
rect 340 4712 372 4744
rect 412 4712 444 4744
rect 484 4712 516 4744
rect 556 4712 588 4744
rect 628 4712 660 4744
rect 700 4712 732 4744
rect 772 4712 804 4744
rect 844 4712 876 4744
rect 916 4712 948 4744
rect 52 4640 84 4672
rect 124 4640 156 4672
rect 196 4640 228 4672
rect 268 4640 300 4672
rect 340 4640 372 4672
rect 412 4640 444 4672
rect 484 4640 516 4672
rect 556 4640 588 4672
rect 628 4640 660 4672
rect 700 4640 732 4672
rect 772 4640 804 4672
rect 844 4640 876 4672
rect 916 4640 948 4672
rect 52 4568 84 4600
rect 124 4568 156 4600
rect 196 4568 228 4600
rect 268 4568 300 4600
rect 340 4568 372 4600
rect 412 4568 444 4600
rect 484 4568 516 4600
rect 556 4568 588 4600
rect 628 4568 660 4600
rect 700 4568 732 4600
rect 772 4568 804 4600
rect 844 4568 876 4600
rect 916 4568 948 4600
rect 52 4496 84 4528
rect 124 4496 156 4528
rect 196 4496 228 4528
rect 268 4496 300 4528
rect 340 4496 372 4528
rect 412 4496 444 4528
rect 484 4496 516 4528
rect 556 4496 588 4528
rect 628 4496 660 4528
rect 700 4496 732 4528
rect 772 4496 804 4528
rect 844 4496 876 4528
rect 916 4496 948 4528
rect 52 4424 84 4456
rect 124 4424 156 4456
rect 196 4424 228 4456
rect 268 4424 300 4456
rect 340 4424 372 4456
rect 412 4424 444 4456
rect 484 4424 516 4456
rect 556 4424 588 4456
rect 628 4424 660 4456
rect 700 4424 732 4456
rect 772 4424 804 4456
rect 844 4424 876 4456
rect 916 4424 948 4456
rect 52 4352 84 4384
rect 124 4352 156 4384
rect 196 4352 228 4384
rect 268 4352 300 4384
rect 340 4352 372 4384
rect 412 4352 444 4384
rect 484 4352 516 4384
rect 556 4352 588 4384
rect 628 4352 660 4384
rect 700 4352 732 4384
rect 772 4352 804 4384
rect 844 4352 876 4384
rect 916 4352 948 4384
rect 52 4280 84 4312
rect 124 4280 156 4312
rect 196 4280 228 4312
rect 268 4280 300 4312
rect 340 4280 372 4312
rect 412 4280 444 4312
rect 484 4280 516 4312
rect 556 4280 588 4312
rect 628 4280 660 4312
rect 700 4280 732 4312
rect 772 4280 804 4312
rect 844 4280 876 4312
rect 916 4280 948 4312
rect 52 4208 84 4240
rect 124 4208 156 4240
rect 196 4208 228 4240
rect 268 4208 300 4240
rect 340 4208 372 4240
rect 412 4208 444 4240
rect 484 4208 516 4240
rect 556 4208 588 4240
rect 628 4208 660 4240
rect 700 4208 732 4240
rect 772 4208 804 4240
rect 844 4208 876 4240
rect 916 4208 948 4240
rect 52 4136 84 4168
rect 124 4136 156 4168
rect 196 4136 228 4168
rect 268 4136 300 4168
rect 340 4136 372 4168
rect 412 4136 444 4168
rect 484 4136 516 4168
rect 556 4136 588 4168
rect 628 4136 660 4168
rect 700 4136 732 4168
rect 772 4136 804 4168
rect 844 4136 876 4168
rect 916 4136 948 4168
rect 52 4064 84 4096
rect 124 4064 156 4096
rect 196 4064 228 4096
rect 268 4064 300 4096
rect 340 4064 372 4096
rect 412 4064 444 4096
rect 484 4064 516 4096
rect 556 4064 588 4096
rect 628 4064 660 4096
rect 700 4064 732 4096
rect 772 4064 804 4096
rect 844 4064 876 4096
rect 916 4064 948 4096
rect 52 3992 84 4024
rect 124 3992 156 4024
rect 196 3992 228 4024
rect 268 3992 300 4024
rect 340 3992 372 4024
rect 412 3992 444 4024
rect 484 3992 516 4024
rect 556 3992 588 4024
rect 628 3992 660 4024
rect 700 3992 732 4024
rect 772 3992 804 4024
rect 844 3992 876 4024
rect 916 3992 948 4024
rect 52 3920 84 3952
rect 124 3920 156 3952
rect 196 3920 228 3952
rect 268 3920 300 3952
rect 340 3920 372 3952
rect 412 3920 444 3952
rect 484 3920 516 3952
rect 556 3920 588 3952
rect 628 3920 660 3952
rect 700 3920 732 3952
rect 772 3920 804 3952
rect 844 3920 876 3952
rect 916 3920 948 3952
rect 52 3848 84 3880
rect 124 3848 156 3880
rect 196 3848 228 3880
rect 268 3848 300 3880
rect 340 3848 372 3880
rect 412 3848 444 3880
rect 484 3848 516 3880
rect 556 3848 588 3880
rect 628 3848 660 3880
rect 700 3848 732 3880
rect 772 3848 804 3880
rect 844 3848 876 3880
rect 916 3848 948 3880
rect 52 3776 84 3808
rect 124 3776 156 3808
rect 196 3776 228 3808
rect 268 3776 300 3808
rect 340 3776 372 3808
rect 412 3776 444 3808
rect 484 3776 516 3808
rect 556 3776 588 3808
rect 628 3776 660 3808
rect 700 3776 732 3808
rect 772 3776 804 3808
rect 844 3776 876 3808
rect 916 3776 948 3808
rect 52 3704 84 3736
rect 124 3704 156 3736
rect 196 3704 228 3736
rect 268 3704 300 3736
rect 340 3704 372 3736
rect 412 3704 444 3736
rect 484 3704 516 3736
rect 556 3704 588 3736
rect 628 3704 660 3736
rect 700 3704 732 3736
rect 772 3704 804 3736
rect 844 3704 876 3736
rect 916 3704 948 3736
rect 52 3632 84 3664
rect 124 3632 156 3664
rect 196 3632 228 3664
rect 268 3632 300 3664
rect 340 3632 372 3664
rect 412 3632 444 3664
rect 484 3632 516 3664
rect 556 3632 588 3664
rect 628 3632 660 3664
rect 700 3632 732 3664
rect 772 3632 804 3664
rect 844 3632 876 3664
rect 916 3632 948 3664
rect 52 3560 84 3592
rect 124 3560 156 3592
rect 196 3560 228 3592
rect 268 3560 300 3592
rect 340 3560 372 3592
rect 412 3560 444 3592
rect 484 3560 516 3592
rect 556 3560 588 3592
rect 628 3560 660 3592
rect 700 3560 732 3592
rect 772 3560 804 3592
rect 844 3560 876 3592
rect 916 3560 948 3592
rect 52 3488 84 3520
rect 124 3488 156 3520
rect 196 3488 228 3520
rect 268 3488 300 3520
rect 340 3488 372 3520
rect 412 3488 444 3520
rect 484 3488 516 3520
rect 556 3488 588 3520
rect 628 3488 660 3520
rect 700 3488 732 3520
rect 772 3488 804 3520
rect 844 3488 876 3520
rect 916 3488 948 3520
rect 52 3416 84 3448
rect 124 3416 156 3448
rect 196 3416 228 3448
rect 268 3416 300 3448
rect 340 3416 372 3448
rect 412 3416 444 3448
rect 484 3416 516 3448
rect 556 3416 588 3448
rect 628 3416 660 3448
rect 700 3416 732 3448
rect 772 3416 804 3448
rect 844 3416 876 3448
rect 916 3416 948 3448
rect 52 3344 84 3376
rect 124 3344 156 3376
rect 196 3344 228 3376
rect 268 3344 300 3376
rect 340 3344 372 3376
rect 412 3344 444 3376
rect 484 3344 516 3376
rect 556 3344 588 3376
rect 628 3344 660 3376
rect 700 3344 732 3376
rect 772 3344 804 3376
rect 844 3344 876 3376
rect 916 3344 948 3376
rect 52 3272 84 3304
rect 124 3272 156 3304
rect 196 3272 228 3304
rect 268 3272 300 3304
rect 340 3272 372 3304
rect 412 3272 444 3304
rect 484 3272 516 3304
rect 556 3272 588 3304
rect 628 3272 660 3304
rect 700 3272 732 3304
rect 772 3272 804 3304
rect 844 3272 876 3304
rect 916 3272 948 3304
rect 52 3200 84 3232
rect 124 3200 156 3232
rect 196 3200 228 3232
rect 268 3200 300 3232
rect 340 3200 372 3232
rect 412 3200 444 3232
rect 484 3200 516 3232
rect 556 3200 588 3232
rect 628 3200 660 3232
rect 700 3200 732 3232
rect 772 3200 804 3232
rect 844 3200 876 3232
rect 916 3200 948 3232
rect 52 3128 84 3160
rect 124 3128 156 3160
rect 196 3128 228 3160
rect 268 3128 300 3160
rect 340 3128 372 3160
rect 412 3128 444 3160
rect 484 3128 516 3160
rect 556 3128 588 3160
rect 628 3128 660 3160
rect 700 3128 732 3160
rect 772 3128 804 3160
rect 844 3128 876 3160
rect 916 3128 948 3160
rect 52 3056 84 3088
rect 124 3056 156 3088
rect 196 3056 228 3088
rect 268 3056 300 3088
rect 340 3056 372 3088
rect 412 3056 444 3088
rect 484 3056 516 3088
rect 556 3056 588 3088
rect 628 3056 660 3088
rect 700 3056 732 3088
rect 772 3056 804 3088
rect 844 3056 876 3088
rect 916 3056 948 3088
rect 52 2984 84 3016
rect 124 2984 156 3016
rect 196 2984 228 3016
rect 268 2984 300 3016
rect 340 2984 372 3016
rect 412 2984 444 3016
rect 484 2984 516 3016
rect 556 2984 588 3016
rect 628 2984 660 3016
rect 700 2984 732 3016
rect 772 2984 804 3016
rect 844 2984 876 3016
rect 916 2984 948 3016
rect 52 2912 84 2944
rect 124 2912 156 2944
rect 196 2912 228 2944
rect 268 2912 300 2944
rect 340 2912 372 2944
rect 412 2912 444 2944
rect 484 2912 516 2944
rect 556 2912 588 2944
rect 628 2912 660 2944
rect 700 2912 732 2944
rect 772 2912 804 2944
rect 844 2912 876 2944
rect 916 2912 948 2944
rect 52 2840 84 2872
rect 124 2840 156 2872
rect 196 2840 228 2872
rect 268 2840 300 2872
rect 340 2840 372 2872
rect 412 2840 444 2872
rect 484 2840 516 2872
rect 556 2840 588 2872
rect 628 2840 660 2872
rect 700 2840 732 2872
rect 772 2840 804 2872
rect 844 2840 876 2872
rect 916 2840 948 2872
rect 52 2768 84 2800
rect 124 2768 156 2800
rect 196 2768 228 2800
rect 268 2768 300 2800
rect 340 2768 372 2800
rect 412 2768 444 2800
rect 484 2768 516 2800
rect 556 2768 588 2800
rect 628 2768 660 2800
rect 700 2768 732 2800
rect 772 2768 804 2800
rect 844 2768 876 2800
rect 916 2768 948 2800
rect 52 2696 84 2728
rect 124 2696 156 2728
rect 196 2696 228 2728
rect 268 2696 300 2728
rect 340 2696 372 2728
rect 412 2696 444 2728
rect 484 2696 516 2728
rect 556 2696 588 2728
rect 628 2696 660 2728
rect 700 2696 732 2728
rect 772 2696 804 2728
rect 844 2696 876 2728
rect 916 2696 948 2728
rect 52 2624 84 2656
rect 124 2624 156 2656
rect 196 2624 228 2656
rect 268 2624 300 2656
rect 340 2624 372 2656
rect 412 2624 444 2656
rect 484 2624 516 2656
rect 556 2624 588 2656
rect 628 2624 660 2656
rect 700 2624 732 2656
rect 772 2624 804 2656
rect 844 2624 876 2656
rect 916 2624 948 2656
rect 52 2552 84 2584
rect 124 2552 156 2584
rect 196 2552 228 2584
rect 268 2552 300 2584
rect 340 2552 372 2584
rect 412 2552 444 2584
rect 484 2552 516 2584
rect 556 2552 588 2584
rect 628 2552 660 2584
rect 700 2552 732 2584
rect 772 2552 804 2584
rect 844 2552 876 2584
rect 916 2552 948 2584
rect 52 2480 84 2512
rect 124 2480 156 2512
rect 196 2480 228 2512
rect 268 2480 300 2512
rect 340 2480 372 2512
rect 412 2480 444 2512
rect 484 2480 516 2512
rect 556 2480 588 2512
rect 628 2480 660 2512
rect 700 2480 732 2512
rect 772 2480 804 2512
rect 844 2480 876 2512
rect 916 2480 948 2512
rect 52 2408 84 2440
rect 124 2408 156 2440
rect 196 2408 228 2440
rect 268 2408 300 2440
rect 340 2408 372 2440
rect 412 2408 444 2440
rect 484 2408 516 2440
rect 556 2408 588 2440
rect 628 2408 660 2440
rect 700 2408 732 2440
rect 772 2408 804 2440
rect 844 2408 876 2440
rect 916 2408 948 2440
rect 52 2336 84 2368
rect 124 2336 156 2368
rect 196 2336 228 2368
rect 268 2336 300 2368
rect 340 2336 372 2368
rect 412 2336 444 2368
rect 484 2336 516 2368
rect 556 2336 588 2368
rect 628 2336 660 2368
rect 700 2336 732 2368
rect 772 2336 804 2368
rect 844 2336 876 2368
rect 916 2336 948 2368
rect 52 2264 84 2296
rect 124 2264 156 2296
rect 196 2264 228 2296
rect 268 2264 300 2296
rect 340 2264 372 2296
rect 412 2264 444 2296
rect 484 2264 516 2296
rect 556 2264 588 2296
rect 628 2264 660 2296
rect 700 2264 732 2296
rect 772 2264 804 2296
rect 844 2264 876 2296
rect 916 2264 948 2296
rect 52 2192 84 2224
rect 124 2192 156 2224
rect 196 2192 228 2224
rect 268 2192 300 2224
rect 340 2192 372 2224
rect 412 2192 444 2224
rect 484 2192 516 2224
rect 556 2192 588 2224
rect 628 2192 660 2224
rect 700 2192 732 2224
rect 772 2192 804 2224
rect 844 2192 876 2224
rect 916 2192 948 2224
rect 52 2120 84 2152
rect 124 2120 156 2152
rect 196 2120 228 2152
rect 268 2120 300 2152
rect 340 2120 372 2152
rect 412 2120 444 2152
rect 484 2120 516 2152
rect 556 2120 588 2152
rect 628 2120 660 2152
rect 700 2120 732 2152
rect 772 2120 804 2152
rect 844 2120 876 2152
rect 916 2120 948 2152
rect 52 2048 84 2080
rect 124 2048 156 2080
rect 196 2048 228 2080
rect 268 2048 300 2080
rect 340 2048 372 2080
rect 412 2048 444 2080
rect 484 2048 516 2080
rect 556 2048 588 2080
rect 628 2048 660 2080
rect 700 2048 732 2080
rect 772 2048 804 2080
rect 844 2048 876 2080
rect 916 2048 948 2080
rect 52 1976 84 2008
rect 124 1976 156 2008
rect 196 1976 228 2008
rect 268 1976 300 2008
rect 340 1976 372 2008
rect 412 1976 444 2008
rect 484 1976 516 2008
rect 556 1976 588 2008
rect 628 1976 660 2008
rect 700 1976 732 2008
rect 772 1976 804 2008
rect 844 1976 876 2008
rect 916 1976 948 2008
rect 52 1904 84 1936
rect 124 1904 156 1936
rect 196 1904 228 1936
rect 268 1904 300 1936
rect 340 1904 372 1936
rect 412 1904 444 1936
rect 484 1904 516 1936
rect 556 1904 588 1936
rect 628 1904 660 1936
rect 700 1904 732 1936
rect 772 1904 804 1936
rect 844 1904 876 1936
rect 916 1904 948 1936
rect 52 1832 84 1864
rect 124 1832 156 1864
rect 196 1832 228 1864
rect 268 1832 300 1864
rect 340 1832 372 1864
rect 412 1832 444 1864
rect 484 1832 516 1864
rect 556 1832 588 1864
rect 628 1832 660 1864
rect 700 1832 732 1864
rect 772 1832 804 1864
rect 844 1832 876 1864
rect 916 1832 948 1864
rect 52 1760 84 1792
rect 124 1760 156 1792
rect 196 1760 228 1792
rect 268 1760 300 1792
rect 340 1760 372 1792
rect 412 1760 444 1792
rect 484 1760 516 1792
rect 556 1760 588 1792
rect 628 1760 660 1792
rect 700 1760 732 1792
rect 772 1760 804 1792
rect 844 1760 876 1792
rect 916 1760 948 1792
rect 52 1688 84 1720
rect 124 1688 156 1720
rect 196 1688 228 1720
rect 268 1688 300 1720
rect 340 1688 372 1720
rect 412 1688 444 1720
rect 484 1688 516 1720
rect 556 1688 588 1720
rect 628 1688 660 1720
rect 700 1688 732 1720
rect 772 1688 804 1720
rect 844 1688 876 1720
rect 916 1688 948 1720
rect 52 1616 84 1648
rect 124 1616 156 1648
rect 196 1616 228 1648
rect 268 1616 300 1648
rect 340 1616 372 1648
rect 412 1616 444 1648
rect 484 1616 516 1648
rect 556 1616 588 1648
rect 628 1616 660 1648
rect 700 1616 732 1648
rect 772 1616 804 1648
rect 844 1616 876 1648
rect 916 1616 948 1648
rect 52 1544 84 1576
rect 124 1544 156 1576
rect 196 1544 228 1576
rect 268 1544 300 1576
rect 340 1544 372 1576
rect 412 1544 444 1576
rect 484 1544 516 1576
rect 556 1544 588 1576
rect 628 1544 660 1576
rect 700 1544 732 1576
rect 772 1544 804 1576
rect 844 1544 876 1576
rect 916 1544 948 1576
rect 52 1472 84 1504
rect 124 1472 156 1504
rect 196 1472 228 1504
rect 268 1472 300 1504
rect 340 1472 372 1504
rect 412 1472 444 1504
rect 484 1472 516 1504
rect 556 1472 588 1504
rect 628 1472 660 1504
rect 700 1472 732 1504
rect 772 1472 804 1504
rect 844 1472 876 1504
rect 916 1472 948 1504
rect 52 1400 84 1432
rect 124 1400 156 1432
rect 196 1400 228 1432
rect 268 1400 300 1432
rect 340 1400 372 1432
rect 412 1400 444 1432
rect 484 1400 516 1432
rect 556 1400 588 1432
rect 628 1400 660 1432
rect 700 1400 732 1432
rect 772 1400 804 1432
rect 844 1400 876 1432
rect 916 1400 948 1432
rect 52 1328 84 1360
rect 124 1328 156 1360
rect 196 1328 228 1360
rect 268 1328 300 1360
rect 340 1328 372 1360
rect 412 1328 444 1360
rect 484 1328 516 1360
rect 556 1328 588 1360
rect 628 1328 660 1360
rect 700 1328 732 1360
rect 772 1328 804 1360
rect 844 1328 876 1360
rect 916 1328 948 1360
rect 52 1256 84 1288
rect 124 1256 156 1288
rect 196 1256 228 1288
rect 268 1256 300 1288
rect 340 1256 372 1288
rect 412 1256 444 1288
rect 484 1256 516 1288
rect 556 1256 588 1288
rect 628 1256 660 1288
rect 700 1256 732 1288
rect 772 1256 804 1288
rect 844 1256 876 1288
rect 916 1256 948 1288
rect 0 33416 1000 33430
rect 0 33384 124 33416
rect 156 33384 196 33416
rect 228 33384 268 33416
rect 300 33384 340 33416
rect 372 33384 412 33416
rect 444 33384 484 33416
rect 516 33384 556 33416
rect 588 33384 628 33416
rect 660 33384 700 33416
rect 732 33384 772 33416
rect 804 33384 844 33416
rect 876 33384 1000 33416
rect 0 33370 1000 33384
rect 0 29716 1000 29730
rect 0 29684 124 29716
rect 156 29684 196 29716
rect 228 29684 268 29716
rect 300 29684 340 29716
rect 372 29684 412 29716
rect 444 29684 484 29716
rect 516 29684 556 29716
rect 588 29684 628 29716
rect 660 29684 700 29716
rect 732 29684 772 29716
rect 804 29684 844 29716
rect 876 29684 1000 29716
rect 0 29670 1000 29684
rect 0 12144 1000 12200
rect 0 12112 52 12144
rect 84 12112 124 12144
rect 156 12112 196 12144
rect 228 12112 268 12144
rect 300 12112 340 12144
rect 372 12112 412 12144
rect 444 12112 484 12144
rect 516 12112 556 12144
rect 588 12112 628 12144
rect 660 12112 700 12144
rect 732 12112 772 12144
rect 804 12112 844 12144
rect 876 12112 916 12144
rect 948 12112 1000 12144
rect 0 12072 1000 12112
rect 0 12040 52 12072
rect 84 12040 124 12072
rect 156 12040 196 12072
rect 228 12040 268 12072
rect 300 12040 340 12072
rect 372 12040 412 12072
rect 444 12040 484 12072
rect 516 12040 556 12072
rect 588 12040 628 12072
rect 660 12040 700 12072
rect 732 12040 772 12072
rect 804 12040 844 12072
rect 876 12040 916 12072
rect 948 12040 1000 12072
rect 0 12000 1000 12040
rect 0 11968 52 12000
rect 84 11968 124 12000
rect 156 11968 196 12000
rect 228 11968 268 12000
rect 300 11968 340 12000
rect 372 11968 412 12000
rect 444 11968 484 12000
rect 516 11968 556 12000
rect 588 11968 628 12000
rect 660 11968 700 12000
rect 732 11968 772 12000
rect 804 11968 844 12000
rect 876 11968 916 12000
rect 948 11968 1000 12000
rect 0 11928 1000 11968
rect 0 11896 52 11928
rect 84 11896 124 11928
rect 156 11896 196 11928
rect 228 11896 268 11928
rect 300 11896 340 11928
rect 372 11896 412 11928
rect 444 11896 484 11928
rect 516 11896 556 11928
rect 588 11896 628 11928
rect 660 11896 700 11928
rect 732 11896 772 11928
rect 804 11896 844 11928
rect 876 11896 916 11928
rect 948 11896 1000 11928
rect 0 11856 1000 11896
rect 0 11824 52 11856
rect 84 11824 124 11856
rect 156 11824 196 11856
rect 228 11824 268 11856
rect 300 11824 340 11856
rect 372 11824 412 11856
rect 444 11824 484 11856
rect 516 11824 556 11856
rect 588 11824 628 11856
rect 660 11824 700 11856
rect 732 11824 772 11856
rect 804 11824 844 11856
rect 876 11824 916 11856
rect 948 11824 1000 11856
rect 0 11784 1000 11824
rect 0 11752 52 11784
rect 84 11752 124 11784
rect 156 11752 196 11784
rect 228 11752 268 11784
rect 300 11752 340 11784
rect 372 11752 412 11784
rect 444 11752 484 11784
rect 516 11752 556 11784
rect 588 11752 628 11784
rect 660 11752 700 11784
rect 732 11752 772 11784
rect 804 11752 844 11784
rect 876 11752 916 11784
rect 948 11752 1000 11784
rect 0 11712 1000 11752
rect 0 11680 52 11712
rect 84 11680 124 11712
rect 156 11680 196 11712
rect 228 11680 268 11712
rect 300 11680 340 11712
rect 372 11680 412 11712
rect 444 11680 484 11712
rect 516 11680 556 11712
rect 588 11680 628 11712
rect 660 11680 700 11712
rect 732 11680 772 11712
rect 804 11680 844 11712
rect 876 11680 916 11712
rect 948 11680 1000 11712
rect 0 11640 1000 11680
rect 0 11608 52 11640
rect 84 11608 124 11640
rect 156 11608 196 11640
rect 228 11608 268 11640
rect 300 11608 340 11640
rect 372 11608 412 11640
rect 444 11608 484 11640
rect 516 11608 556 11640
rect 588 11608 628 11640
rect 660 11608 700 11640
rect 732 11608 772 11640
rect 804 11608 844 11640
rect 876 11608 916 11640
rect 948 11608 1000 11640
rect 0 11568 1000 11608
rect 0 11536 52 11568
rect 84 11536 124 11568
rect 156 11536 196 11568
rect 228 11536 268 11568
rect 300 11536 340 11568
rect 372 11536 412 11568
rect 444 11536 484 11568
rect 516 11536 556 11568
rect 588 11536 628 11568
rect 660 11536 700 11568
rect 732 11536 772 11568
rect 804 11536 844 11568
rect 876 11536 916 11568
rect 948 11536 1000 11568
rect 0 11496 1000 11536
rect 0 11464 52 11496
rect 84 11464 124 11496
rect 156 11464 196 11496
rect 228 11464 268 11496
rect 300 11464 340 11496
rect 372 11464 412 11496
rect 444 11464 484 11496
rect 516 11464 556 11496
rect 588 11464 628 11496
rect 660 11464 700 11496
rect 732 11464 772 11496
rect 804 11464 844 11496
rect 876 11464 916 11496
rect 948 11464 1000 11496
rect 0 11424 1000 11464
rect 0 11392 52 11424
rect 84 11392 124 11424
rect 156 11392 196 11424
rect 228 11392 268 11424
rect 300 11392 340 11424
rect 372 11392 412 11424
rect 444 11392 484 11424
rect 516 11392 556 11424
rect 588 11392 628 11424
rect 660 11392 700 11424
rect 732 11392 772 11424
rect 804 11392 844 11424
rect 876 11392 916 11424
rect 948 11392 1000 11424
rect 0 11352 1000 11392
rect 0 11320 52 11352
rect 84 11320 124 11352
rect 156 11320 196 11352
rect 228 11320 268 11352
rect 300 11320 340 11352
rect 372 11320 412 11352
rect 444 11320 484 11352
rect 516 11320 556 11352
rect 588 11320 628 11352
rect 660 11320 700 11352
rect 732 11320 772 11352
rect 804 11320 844 11352
rect 876 11320 916 11352
rect 948 11320 1000 11352
rect 0 11280 1000 11320
rect 0 11248 52 11280
rect 84 11248 124 11280
rect 156 11248 196 11280
rect 228 11248 268 11280
rect 300 11248 340 11280
rect 372 11248 412 11280
rect 444 11248 484 11280
rect 516 11248 556 11280
rect 588 11248 628 11280
rect 660 11248 700 11280
rect 732 11248 772 11280
rect 804 11248 844 11280
rect 876 11248 916 11280
rect 948 11248 1000 11280
rect 0 11208 1000 11248
rect 0 11176 52 11208
rect 84 11176 124 11208
rect 156 11176 196 11208
rect 228 11176 268 11208
rect 300 11176 340 11208
rect 372 11176 412 11208
rect 444 11176 484 11208
rect 516 11176 556 11208
rect 588 11176 628 11208
rect 660 11176 700 11208
rect 732 11176 772 11208
rect 804 11176 844 11208
rect 876 11176 916 11208
rect 948 11176 1000 11208
rect 0 11136 1000 11176
rect 0 11104 52 11136
rect 84 11104 124 11136
rect 156 11104 196 11136
rect 228 11104 268 11136
rect 300 11104 340 11136
rect 372 11104 412 11136
rect 444 11104 484 11136
rect 516 11104 556 11136
rect 588 11104 628 11136
rect 660 11104 700 11136
rect 732 11104 772 11136
rect 804 11104 844 11136
rect 876 11104 916 11136
rect 948 11104 1000 11136
rect 0 11064 1000 11104
rect 0 11032 52 11064
rect 84 11032 124 11064
rect 156 11032 196 11064
rect 228 11032 268 11064
rect 300 11032 340 11064
rect 372 11032 412 11064
rect 444 11032 484 11064
rect 516 11032 556 11064
rect 588 11032 628 11064
rect 660 11032 700 11064
rect 732 11032 772 11064
rect 804 11032 844 11064
rect 876 11032 916 11064
rect 948 11032 1000 11064
rect 0 10992 1000 11032
rect 0 10960 52 10992
rect 84 10960 124 10992
rect 156 10960 196 10992
rect 228 10960 268 10992
rect 300 10960 340 10992
rect 372 10960 412 10992
rect 444 10960 484 10992
rect 516 10960 556 10992
rect 588 10960 628 10992
rect 660 10960 700 10992
rect 732 10960 772 10992
rect 804 10960 844 10992
rect 876 10960 916 10992
rect 948 10960 1000 10992
rect 0 10920 1000 10960
rect 0 10888 52 10920
rect 84 10888 124 10920
rect 156 10888 196 10920
rect 228 10888 268 10920
rect 300 10888 340 10920
rect 372 10888 412 10920
rect 444 10888 484 10920
rect 516 10888 556 10920
rect 588 10888 628 10920
rect 660 10888 700 10920
rect 732 10888 772 10920
rect 804 10888 844 10920
rect 876 10888 916 10920
rect 948 10888 1000 10920
rect 0 10848 1000 10888
rect 0 10816 52 10848
rect 84 10816 124 10848
rect 156 10816 196 10848
rect 228 10816 268 10848
rect 300 10816 340 10848
rect 372 10816 412 10848
rect 444 10816 484 10848
rect 516 10816 556 10848
rect 588 10816 628 10848
rect 660 10816 700 10848
rect 732 10816 772 10848
rect 804 10816 844 10848
rect 876 10816 916 10848
rect 948 10816 1000 10848
rect 0 10776 1000 10816
rect 0 10744 52 10776
rect 84 10744 124 10776
rect 156 10744 196 10776
rect 228 10744 268 10776
rect 300 10744 340 10776
rect 372 10744 412 10776
rect 444 10744 484 10776
rect 516 10744 556 10776
rect 588 10744 628 10776
rect 660 10744 700 10776
rect 732 10744 772 10776
rect 804 10744 844 10776
rect 876 10744 916 10776
rect 948 10744 1000 10776
rect 0 10704 1000 10744
rect 0 10672 52 10704
rect 84 10672 124 10704
rect 156 10672 196 10704
rect 228 10672 268 10704
rect 300 10672 340 10704
rect 372 10672 412 10704
rect 444 10672 484 10704
rect 516 10672 556 10704
rect 588 10672 628 10704
rect 660 10672 700 10704
rect 732 10672 772 10704
rect 804 10672 844 10704
rect 876 10672 916 10704
rect 948 10672 1000 10704
rect 0 10632 1000 10672
rect 0 10600 52 10632
rect 84 10600 124 10632
rect 156 10600 196 10632
rect 228 10600 268 10632
rect 300 10600 340 10632
rect 372 10600 412 10632
rect 444 10600 484 10632
rect 516 10600 556 10632
rect 588 10600 628 10632
rect 660 10600 700 10632
rect 732 10600 772 10632
rect 804 10600 844 10632
rect 876 10600 916 10632
rect 948 10600 1000 10632
rect 0 10560 1000 10600
rect 0 10528 52 10560
rect 84 10528 124 10560
rect 156 10528 196 10560
rect 228 10528 268 10560
rect 300 10528 340 10560
rect 372 10528 412 10560
rect 444 10528 484 10560
rect 516 10528 556 10560
rect 588 10528 628 10560
rect 660 10528 700 10560
rect 732 10528 772 10560
rect 804 10528 844 10560
rect 876 10528 916 10560
rect 948 10528 1000 10560
rect 0 10488 1000 10528
rect 0 10456 52 10488
rect 84 10456 124 10488
rect 156 10456 196 10488
rect 228 10456 268 10488
rect 300 10456 340 10488
rect 372 10456 412 10488
rect 444 10456 484 10488
rect 516 10456 556 10488
rect 588 10456 628 10488
rect 660 10456 700 10488
rect 732 10456 772 10488
rect 804 10456 844 10488
rect 876 10456 916 10488
rect 948 10456 1000 10488
rect 0 10416 1000 10456
rect 0 10384 52 10416
rect 84 10384 124 10416
rect 156 10384 196 10416
rect 228 10384 268 10416
rect 300 10384 340 10416
rect 372 10384 412 10416
rect 444 10384 484 10416
rect 516 10384 556 10416
rect 588 10384 628 10416
rect 660 10384 700 10416
rect 732 10384 772 10416
rect 804 10384 844 10416
rect 876 10384 916 10416
rect 948 10384 1000 10416
rect 0 10344 1000 10384
rect 0 10312 52 10344
rect 84 10312 124 10344
rect 156 10312 196 10344
rect 228 10312 268 10344
rect 300 10312 340 10344
rect 372 10312 412 10344
rect 444 10312 484 10344
rect 516 10312 556 10344
rect 588 10312 628 10344
rect 660 10312 700 10344
rect 732 10312 772 10344
rect 804 10312 844 10344
rect 876 10312 916 10344
rect 948 10312 1000 10344
rect 0 10272 1000 10312
rect 0 10240 52 10272
rect 84 10240 124 10272
rect 156 10240 196 10272
rect 228 10240 268 10272
rect 300 10240 340 10272
rect 372 10240 412 10272
rect 444 10240 484 10272
rect 516 10240 556 10272
rect 588 10240 628 10272
rect 660 10240 700 10272
rect 732 10240 772 10272
rect 804 10240 844 10272
rect 876 10240 916 10272
rect 948 10240 1000 10272
rect 0 10200 1000 10240
rect 0 10168 52 10200
rect 84 10168 124 10200
rect 156 10168 196 10200
rect 228 10168 268 10200
rect 300 10168 340 10200
rect 372 10168 412 10200
rect 444 10168 484 10200
rect 516 10168 556 10200
rect 588 10168 628 10200
rect 660 10168 700 10200
rect 732 10168 772 10200
rect 804 10168 844 10200
rect 876 10168 916 10200
rect 948 10168 1000 10200
rect 0 10128 1000 10168
rect 0 10096 52 10128
rect 84 10096 124 10128
rect 156 10096 196 10128
rect 228 10096 268 10128
rect 300 10096 340 10128
rect 372 10096 412 10128
rect 444 10096 484 10128
rect 516 10096 556 10128
rect 588 10096 628 10128
rect 660 10096 700 10128
rect 732 10096 772 10128
rect 804 10096 844 10128
rect 876 10096 916 10128
rect 948 10096 1000 10128
rect 0 10056 1000 10096
rect 0 10024 52 10056
rect 84 10024 124 10056
rect 156 10024 196 10056
rect 228 10024 268 10056
rect 300 10024 340 10056
rect 372 10024 412 10056
rect 444 10024 484 10056
rect 516 10024 556 10056
rect 588 10024 628 10056
rect 660 10024 700 10056
rect 732 10024 772 10056
rect 804 10024 844 10056
rect 876 10024 916 10056
rect 948 10024 1000 10056
rect 0 9984 1000 10024
rect 0 9952 52 9984
rect 84 9952 124 9984
rect 156 9952 196 9984
rect 228 9952 268 9984
rect 300 9952 340 9984
rect 372 9952 412 9984
rect 444 9952 484 9984
rect 516 9952 556 9984
rect 588 9952 628 9984
rect 660 9952 700 9984
rect 732 9952 772 9984
rect 804 9952 844 9984
rect 876 9952 916 9984
rect 948 9952 1000 9984
rect 0 9912 1000 9952
rect 0 9880 52 9912
rect 84 9880 124 9912
rect 156 9880 196 9912
rect 228 9880 268 9912
rect 300 9880 340 9912
rect 372 9880 412 9912
rect 444 9880 484 9912
rect 516 9880 556 9912
rect 588 9880 628 9912
rect 660 9880 700 9912
rect 732 9880 772 9912
rect 804 9880 844 9912
rect 876 9880 916 9912
rect 948 9880 1000 9912
rect 0 9840 1000 9880
rect 0 9808 52 9840
rect 84 9808 124 9840
rect 156 9808 196 9840
rect 228 9808 268 9840
rect 300 9808 340 9840
rect 372 9808 412 9840
rect 444 9808 484 9840
rect 516 9808 556 9840
rect 588 9808 628 9840
rect 660 9808 700 9840
rect 732 9808 772 9840
rect 804 9808 844 9840
rect 876 9808 916 9840
rect 948 9808 1000 9840
rect 0 9768 1000 9808
rect 0 9736 52 9768
rect 84 9736 124 9768
rect 156 9736 196 9768
rect 228 9736 268 9768
rect 300 9736 340 9768
rect 372 9736 412 9768
rect 444 9736 484 9768
rect 516 9736 556 9768
rect 588 9736 628 9768
rect 660 9736 700 9768
rect 732 9736 772 9768
rect 804 9736 844 9768
rect 876 9736 916 9768
rect 948 9736 1000 9768
rect 0 9696 1000 9736
rect 0 9664 52 9696
rect 84 9664 124 9696
rect 156 9664 196 9696
rect 228 9664 268 9696
rect 300 9664 340 9696
rect 372 9664 412 9696
rect 444 9664 484 9696
rect 516 9664 556 9696
rect 588 9664 628 9696
rect 660 9664 700 9696
rect 732 9664 772 9696
rect 804 9664 844 9696
rect 876 9664 916 9696
rect 948 9664 1000 9696
rect 0 9624 1000 9664
rect 0 9592 52 9624
rect 84 9592 124 9624
rect 156 9592 196 9624
rect 228 9592 268 9624
rect 300 9592 340 9624
rect 372 9592 412 9624
rect 444 9592 484 9624
rect 516 9592 556 9624
rect 588 9592 628 9624
rect 660 9592 700 9624
rect 732 9592 772 9624
rect 804 9592 844 9624
rect 876 9592 916 9624
rect 948 9592 1000 9624
rect 0 9552 1000 9592
rect 0 9520 52 9552
rect 84 9520 124 9552
rect 156 9520 196 9552
rect 228 9520 268 9552
rect 300 9520 340 9552
rect 372 9520 412 9552
rect 444 9520 484 9552
rect 516 9520 556 9552
rect 588 9520 628 9552
rect 660 9520 700 9552
rect 732 9520 772 9552
rect 804 9520 844 9552
rect 876 9520 916 9552
rect 948 9520 1000 9552
rect 0 9480 1000 9520
rect 0 9448 52 9480
rect 84 9448 124 9480
rect 156 9448 196 9480
rect 228 9448 268 9480
rect 300 9448 340 9480
rect 372 9448 412 9480
rect 444 9448 484 9480
rect 516 9448 556 9480
rect 588 9448 628 9480
rect 660 9448 700 9480
rect 732 9448 772 9480
rect 804 9448 844 9480
rect 876 9448 916 9480
rect 948 9448 1000 9480
rect 0 9408 1000 9448
rect 0 9376 52 9408
rect 84 9376 124 9408
rect 156 9376 196 9408
rect 228 9376 268 9408
rect 300 9376 340 9408
rect 372 9376 412 9408
rect 444 9376 484 9408
rect 516 9376 556 9408
rect 588 9376 628 9408
rect 660 9376 700 9408
rect 732 9376 772 9408
rect 804 9376 844 9408
rect 876 9376 916 9408
rect 948 9376 1000 9408
rect 0 9336 1000 9376
rect 0 9304 52 9336
rect 84 9304 124 9336
rect 156 9304 196 9336
rect 228 9304 268 9336
rect 300 9304 340 9336
rect 372 9304 412 9336
rect 444 9304 484 9336
rect 516 9304 556 9336
rect 588 9304 628 9336
rect 660 9304 700 9336
rect 732 9304 772 9336
rect 804 9304 844 9336
rect 876 9304 916 9336
rect 948 9304 1000 9336
rect 0 9264 1000 9304
rect 0 9232 52 9264
rect 84 9232 124 9264
rect 156 9232 196 9264
rect 228 9232 268 9264
rect 300 9232 340 9264
rect 372 9232 412 9264
rect 444 9232 484 9264
rect 516 9232 556 9264
rect 588 9232 628 9264
rect 660 9232 700 9264
rect 732 9232 772 9264
rect 804 9232 844 9264
rect 876 9232 916 9264
rect 948 9232 1000 9264
rect 0 9192 1000 9232
rect 0 9160 52 9192
rect 84 9160 124 9192
rect 156 9160 196 9192
rect 228 9160 268 9192
rect 300 9160 340 9192
rect 372 9160 412 9192
rect 444 9160 484 9192
rect 516 9160 556 9192
rect 588 9160 628 9192
rect 660 9160 700 9192
rect 732 9160 772 9192
rect 804 9160 844 9192
rect 876 9160 916 9192
rect 948 9160 1000 9192
rect 0 9120 1000 9160
rect 0 9088 52 9120
rect 84 9088 124 9120
rect 156 9088 196 9120
rect 228 9088 268 9120
rect 300 9088 340 9120
rect 372 9088 412 9120
rect 444 9088 484 9120
rect 516 9088 556 9120
rect 588 9088 628 9120
rect 660 9088 700 9120
rect 732 9088 772 9120
rect 804 9088 844 9120
rect 876 9088 916 9120
rect 948 9088 1000 9120
rect 0 9048 1000 9088
rect 0 9016 52 9048
rect 84 9016 124 9048
rect 156 9016 196 9048
rect 228 9016 268 9048
rect 300 9016 340 9048
rect 372 9016 412 9048
rect 444 9016 484 9048
rect 516 9016 556 9048
rect 588 9016 628 9048
rect 660 9016 700 9048
rect 732 9016 772 9048
rect 804 9016 844 9048
rect 876 9016 916 9048
rect 948 9016 1000 9048
rect 0 8976 1000 9016
rect 0 8944 52 8976
rect 84 8944 124 8976
rect 156 8944 196 8976
rect 228 8944 268 8976
rect 300 8944 340 8976
rect 372 8944 412 8976
rect 444 8944 484 8976
rect 516 8944 556 8976
rect 588 8944 628 8976
rect 660 8944 700 8976
rect 732 8944 772 8976
rect 804 8944 844 8976
rect 876 8944 916 8976
rect 948 8944 1000 8976
rect 0 8904 1000 8944
rect 0 8872 52 8904
rect 84 8872 124 8904
rect 156 8872 196 8904
rect 228 8872 268 8904
rect 300 8872 340 8904
rect 372 8872 412 8904
rect 444 8872 484 8904
rect 516 8872 556 8904
rect 588 8872 628 8904
rect 660 8872 700 8904
rect 732 8872 772 8904
rect 804 8872 844 8904
rect 876 8872 916 8904
rect 948 8872 1000 8904
rect 0 8832 1000 8872
rect 0 8800 52 8832
rect 84 8800 124 8832
rect 156 8800 196 8832
rect 228 8800 268 8832
rect 300 8800 340 8832
rect 372 8800 412 8832
rect 444 8800 484 8832
rect 516 8800 556 8832
rect 588 8800 628 8832
rect 660 8800 700 8832
rect 732 8800 772 8832
rect 804 8800 844 8832
rect 876 8800 916 8832
rect 948 8800 1000 8832
rect 0 8760 1000 8800
rect 0 8728 52 8760
rect 84 8728 124 8760
rect 156 8728 196 8760
rect 228 8728 268 8760
rect 300 8728 340 8760
rect 372 8728 412 8760
rect 444 8728 484 8760
rect 516 8728 556 8760
rect 588 8728 628 8760
rect 660 8728 700 8760
rect 732 8728 772 8760
rect 804 8728 844 8760
rect 876 8728 916 8760
rect 948 8728 1000 8760
rect 0 8688 1000 8728
rect 0 8656 52 8688
rect 84 8656 124 8688
rect 156 8656 196 8688
rect 228 8656 268 8688
rect 300 8656 340 8688
rect 372 8656 412 8688
rect 444 8656 484 8688
rect 516 8656 556 8688
rect 588 8656 628 8688
rect 660 8656 700 8688
rect 732 8656 772 8688
rect 804 8656 844 8688
rect 876 8656 916 8688
rect 948 8656 1000 8688
rect 0 8616 1000 8656
rect 0 8584 52 8616
rect 84 8584 124 8616
rect 156 8584 196 8616
rect 228 8584 268 8616
rect 300 8584 340 8616
rect 372 8584 412 8616
rect 444 8584 484 8616
rect 516 8584 556 8616
rect 588 8584 628 8616
rect 660 8584 700 8616
rect 732 8584 772 8616
rect 804 8584 844 8616
rect 876 8584 916 8616
rect 948 8584 1000 8616
rect 0 8544 1000 8584
rect 0 8512 52 8544
rect 84 8512 124 8544
rect 156 8512 196 8544
rect 228 8512 268 8544
rect 300 8512 340 8544
rect 372 8512 412 8544
rect 444 8512 484 8544
rect 516 8512 556 8544
rect 588 8512 628 8544
rect 660 8512 700 8544
rect 732 8512 772 8544
rect 804 8512 844 8544
rect 876 8512 916 8544
rect 948 8512 1000 8544
rect 0 8472 1000 8512
rect 0 8440 52 8472
rect 84 8440 124 8472
rect 156 8440 196 8472
rect 228 8440 268 8472
rect 300 8440 340 8472
rect 372 8440 412 8472
rect 444 8440 484 8472
rect 516 8440 556 8472
rect 588 8440 628 8472
rect 660 8440 700 8472
rect 732 8440 772 8472
rect 804 8440 844 8472
rect 876 8440 916 8472
rect 948 8440 1000 8472
rect 0 8400 1000 8440
rect 0 8368 52 8400
rect 84 8368 124 8400
rect 156 8368 196 8400
rect 228 8368 268 8400
rect 300 8368 340 8400
rect 372 8368 412 8400
rect 444 8368 484 8400
rect 516 8368 556 8400
rect 588 8368 628 8400
rect 660 8368 700 8400
rect 732 8368 772 8400
rect 804 8368 844 8400
rect 876 8368 916 8400
rect 948 8368 1000 8400
rect 0 8328 1000 8368
rect 0 8296 52 8328
rect 84 8296 124 8328
rect 156 8296 196 8328
rect 228 8296 268 8328
rect 300 8296 340 8328
rect 372 8296 412 8328
rect 444 8296 484 8328
rect 516 8296 556 8328
rect 588 8296 628 8328
rect 660 8296 700 8328
rect 732 8296 772 8328
rect 804 8296 844 8328
rect 876 8296 916 8328
rect 948 8296 1000 8328
rect 0 8256 1000 8296
rect 0 8224 52 8256
rect 84 8224 124 8256
rect 156 8224 196 8256
rect 228 8224 268 8256
rect 300 8224 340 8256
rect 372 8224 412 8256
rect 444 8224 484 8256
rect 516 8224 556 8256
rect 588 8224 628 8256
rect 660 8224 700 8256
rect 732 8224 772 8256
rect 804 8224 844 8256
rect 876 8224 916 8256
rect 948 8224 1000 8256
rect 0 8184 1000 8224
rect 0 8152 52 8184
rect 84 8152 124 8184
rect 156 8152 196 8184
rect 228 8152 268 8184
rect 300 8152 340 8184
rect 372 8152 412 8184
rect 444 8152 484 8184
rect 516 8152 556 8184
rect 588 8152 628 8184
rect 660 8152 700 8184
rect 732 8152 772 8184
rect 804 8152 844 8184
rect 876 8152 916 8184
rect 948 8152 1000 8184
rect 0 8112 1000 8152
rect 0 8080 52 8112
rect 84 8080 124 8112
rect 156 8080 196 8112
rect 228 8080 268 8112
rect 300 8080 340 8112
rect 372 8080 412 8112
rect 444 8080 484 8112
rect 516 8080 556 8112
rect 588 8080 628 8112
rect 660 8080 700 8112
rect 732 8080 772 8112
rect 804 8080 844 8112
rect 876 8080 916 8112
rect 948 8080 1000 8112
rect 0 8040 1000 8080
rect 0 8008 52 8040
rect 84 8008 124 8040
rect 156 8008 196 8040
rect 228 8008 268 8040
rect 300 8008 340 8040
rect 372 8008 412 8040
rect 444 8008 484 8040
rect 516 8008 556 8040
rect 588 8008 628 8040
rect 660 8008 700 8040
rect 732 8008 772 8040
rect 804 8008 844 8040
rect 876 8008 916 8040
rect 948 8008 1000 8040
rect 0 7968 1000 8008
rect 0 7936 52 7968
rect 84 7936 124 7968
rect 156 7936 196 7968
rect 228 7936 268 7968
rect 300 7936 340 7968
rect 372 7936 412 7968
rect 444 7936 484 7968
rect 516 7936 556 7968
rect 588 7936 628 7968
rect 660 7936 700 7968
rect 732 7936 772 7968
rect 804 7936 844 7968
rect 876 7936 916 7968
rect 948 7936 1000 7968
rect 0 7896 1000 7936
rect 0 7864 52 7896
rect 84 7864 124 7896
rect 156 7864 196 7896
rect 228 7864 268 7896
rect 300 7864 340 7896
rect 372 7864 412 7896
rect 444 7864 484 7896
rect 516 7864 556 7896
rect 588 7864 628 7896
rect 660 7864 700 7896
rect 732 7864 772 7896
rect 804 7864 844 7896
rect 876 7864 916 7896
rect 948 7864 1000 7896
rect 0 7824 1000 7864
rect 0 7792 52 7824
rect 84 7792 124 7824
rect 156 7792 196 7824
rect 228 7792 268 7824
rect 300 7792 340 7824
rect 372 7792 412 7824
rect 444 7792 484 7824
rect 516 7792 556 7824
rect 588 7792 628 7824
rect 660 7792 700 7824
rect 732 7792 772 7824
rect 804 7792 844 7824
rect 876 7792 916 7824
rect 948 7792 1000 7824
rect 0 7752 1000 7792
rect 0 7720 52 7752
rect 84 7720 124 7752
rect 156 7720 196 7752
rect 228 7720 268 7752
rect 300 7720 340 7752
rect 372 7720 412 7752
rect 444 7720 484 7752
rect 516 7720 556 7752
rect 588 7720 628 7752
rect 660 7720 700 7752
rect 732 7720 772 7752
rect 804 7720 844 7752
rect 876 7720 916 7752
rect 948 7720 1000 7752
rect 0 7680 1000 7720
rect 0 7648 52 7680
rect 84 7648 124 7680
rect 156 7648 196 7680
rect 228 7648 268 7680
rect 300 7648 340 7680
rect 372 7648 412 7680
rect 444 7648 484 7680
rect 516 7648 556 7680
rect 588 7648 628 7680
rect 660 7648 700 7680
rect 732 7648 772 7680
rect 804 7648 844 7680
rect 876 7648 916 7680
rect 948 7648 1000 7680
rect 0 7608 1000 7648
rect 0 7576 52 7608
rect 84 7576 124 7608
rect 156 7576 196 7608
rect 228 7576 268 7608
rect 300 7576 340 7608
rect 372 7576 412 7608
rect 444 7576 484 7608
rect 516 7576 556 7608
rect 588 7576 628 7608
rect 660 7576 700 7608
rect 732 7576 772 7608
rect 804 7576 844 7608
rect 876 7576 916 7608
rect 948 7576 1000 7608
rect 0 7536 1000 7576
rect 0 7504 52 7536
rect 84 7504 124 7536
rect 156 7504 196 7536
rect 228 7504 268 7536
rect 300 7504 340 7536
rect 372 7504 412 7536
rect 444 7504 484 7536
rect 516 7504 556 7536
rect 588 7504 628 7536
rect 660 7504 700 7536
rect 732 7504 772 7536
rect 804 7504 844 7536
rect 876 7504 916 7536
rect 948 7504 1000 7536
rect 0 7464 1000 7504
rect 0 7432 52 7464
rect 84 7432 124 7464
rect 156 7432 196 7464
rect 228 7432 268 7464
rect 300 7432 340 7464
rect 372 7432 412 7464
rect 444 7432 484 7464
rect 516 7432 556 7464
rect 588 7432 628 7464
rect 660 7432 700 7464
rect 732 7432 772 7464
rect 804 7432 844 7464
rect 876 7432 916 7464
rect 948 7432 1000 7464
rect 0 7392 1000 7432
rect 0 7360 52 7392
rect 84 7360 124 7392
rect 156 7360 196 7392
rect 228 7360 268 7392
rect 300 7360 340 7392
rect 372 7360 412 7392
rect 444 7360 484 7392
rect 516 7360 556 7392
rect 588 7360 628 7392
rect 660 7360 700 7392
rect 732 7360 772 7392
rect 804 7360 844 7392
rect 876 7360 916 7392
rect 948 7360 1000 7392
rect 0 7320 1000 7360
rect 0 7288 52 7320
rect 84 7288 124 7320
rect 156 7288 196 7320
rect 228 7288 268 7320
rect 300 7288 340 7320
rect 372 7288 412 7320
rect 444 7288 484 7320
rect 516 7288 556 7320
rect 588 7288 628 7320
rect 660 7288 700 7320
rect 732 7288 772 7320
rect 804 7288 844 7320
rect 876 7288 916 7320
rect 948 7288 1000 7320
rect 0 7248 1000 7288
rect 0 7216 52 7248
rect 84 7216 124 7248
rect 156 7216 196 7248
rect 228 7216 268 7248
rect 300 7216 340 7248
rect 372 7216 412 7248
rect 444 7216 484 7248
rect 516 7216 556 7248
rect 588 7216 628 7248
rect 660 7216 700 7248
rect 732 7216 772 7248
rect 804 7216 844 7248
rect 876 7216 916 7248
rect 948 7216 1000 7248
rect 0 7176 1000 7216
rect 0 7144 52 7176
rect 84 7144 124 7176
rect 156 7144 196 7176
rect 228 7144 268 7176
rect 300 7144 340 7176
rect 372 7144 412 7176
rect 444 7144 484 7176
rect 516 7144 556 7176
rect 588 7144 628 7176
rect 660 7144 700 7176
rect 732 7144 772 7176
rect 804 7144 844 7176
rect 876 7144 916 7176
rect 948 7144 1000 7176
rect 0 7104 1000 7144
rect 0 7072 52 7104
rect 84 7072 124 7104
rect 156 7072 196 7104
rect 228 7072 268 7104
rect 300 7072 340 7104
rect 372 7072 412 7104
rect 444 7072 484 7104
rect 516 7072 556 7104
rect 588 7072 628 7104
rect 660 7072 700 7104
rect 732 7072 772 7104
rect 804 7072 844 7104
rect 876 7072 916 7104
rect 948 7072 1000 7104
rect 0 7032 1000 7072
rect 0 7000 52 7032
rect 84 7000 124 7032
rect 156 7000 196 7032
rect 228 7000 268 7032
rect 300 7000 340 7032
rect 372 7000 412 7032
rect 444 7000 484 7032
rect 516 7000 556 7032
rect 588 7000 628 7032
rect 660 7000 700 7032
rect 732 7000 772 7032
rect 804 7000 844 7032
rect 876 7000 916 7032
rect 948 7000 1000 7032
rect 0 6960 1000 7000
rect 0 6928 52 6960
rect 84 6928 124 6960
rect 156 6928 196 6960
rect 228 6928 268 6960
rect 300 6928 340 6960
rect 372 6928 412 6960
rect 444 6928 484 6960
rect 516 6928 556 6960
rect 588 6928 628 6960
rect 660 6928 700 6960
rect 732 6928 772 6960
rect 804 6928 844 6960
rect 876 6928 916 6960
rect 948 6928 1000 6960
rect 0 6888 1000 6928
rect 0 6856 52 6888
rect 84 6856 124 6888
rect 156 6856 196 6888
rect 228 6856 268 6888
rect 300 6856 340 6888
rect 372 6856 412 6888
rect 444 6856 484 6888
rect 516 6856 556 6888
rect 588 6856 628 6888
rect 660 6856 700 6888
rect 732 6856 772 6888
rect 804 6856 844 6888
rect 876 6856 916 6888
rect 948 6856 1000 6888
rect 0 6800 1000 6856
rect 0 6544 1000 6600
rect 0 6512 52 6544
rect 84 6512 124 6544
rect 156 6512 196 6544
rect 228 6512 268 6544
rect 300 6512 340 6544
rect 372 6512 412 6544
rect 444 6512 484 6544
rect 516 6512 556 6544
rect 588 6512 628 6544
rect 660 6512 700 6544
rect 732 6512 772 6544
rect 804 6512 844 6544
rect 876 6512 916 6544
rect 948 6512 1000 6544
rect 0 6472 1000 6512
rect 0 6440 52 6472
rect 84 6440 124 6472
rect 156 6440 196 6472
rect 228 6440 268 6472
rect 300 6440 340 6472
rect 372 6440 412 6472
rect 444 6440 484 6472
rect 516 6440 556 6472
rect 588 6440 628 6472
rect 660 6440 700 6472
rect 732 6440 772 6472
rect 804 6440 844 6472
rect 876 6440 916 6472
rect 948 6440 1000 6472
rect 0 6400 1000 6440
rect 0 6368 52 6400
rect 84 6368 124 6400
rect 156 6368 196 6400
rect 228 6368 268 6400
rect 300 6368 340 6400
rect 372 6368 412 6400
rect 444 6368 484 6400
rect 516 6368 556 6400
rect 588 6368 628 6400
rect 660 6368 700 6400
rect 732 6368 772 6400
rect 804 6368 844 6400
rect 876 6368 916 6400
rect 948 6368 1000 6400
rect 0 6328 1000 6368
rect 0 6296 52 6328
rect 84 6296 124 6328
rect 156 6296 196 6328
rect 228 6296 268 6328
rect 300 6296 340 6328
rect 372 6296 412 6328
rect 444 6296 484 6328
rect 516 6296 556 6328
rect 588 6296 628 6328
rect 660 6296 700 6328
rect 732 6296 772 6328
rect 804 6296 844 6328
rect 876 6296 916 6328
rect 948 6296 1000 6328
rect 0 6256 1000 6296
rect 0 6224 52 6256
rect 84 6224 124 6256
rect 156 6224 196 6256
rect 228 6224 268 6256
rect 300 6224 340 6256
rect 372 6224 412 6256
rect 444 6224 484 6256
rect 516 6224 556 6256
rect 588 6224 628 6256
rect 660 6224 700 6256
rect 732 6224 772 6256
rect 804 6224 844 6256
rect 876 6224 916 6256
rect 948 6224 1000 6256
rect 0 6184 1000 6224
rect 0 6152 52 6184
rect 84 6152 124 6184
rect 156 6152 196 6184
rect 228 6152 268 6184
rect 300 6152 340 6184
rect 372 6152 412 6184
rect 444 6152 484 6184
rect 516 6152 556 6184
rect 588 6152 628 6184
rect 660 6152 700 6184
rect 732 6152 772 6184
rect 804 6152 844 6184
rect 876 6152 916 6184
rect 948 6152 1000 6184
rect 0 6112 1000 6152
rect 0 6080 52 6112
rect 84 6080 124 6112
rect 156 6080 196 6112
rect 228 6080 268 6112
rect 300 6080 340 6112
rect 372 6080 412 6112
rect 444 6080 484 6112
rect 516 6080 556 6112
rect 588 6080 628 6112
rect 660 6080 700 6112
rect 732 6080 772 6112
rect 804 6080 844 6112
rect 876 6080 916 6112
rect 948 6080 1000 6112
rect 0 6040 1000 6080
rect 0 6008 52 6040
rect 84 6008 124 6040
rect 156 6008 196 6040
rect 228 6008 268 6040
rect 300 6008 340 6040
rect 372 6008 412 6040
rect 444 6008 484 6040
rect 516 6008 556 6040
rect 588 6008 628 6040
rect 660 6008 700 6040
rect 732 6008 772 6040
rect 804 6008 844 6040
rect 876 6008 916 6040
rect 948 6008 1000 6040
rect 0 5968 1000 6008
rect 0 5936 52 5968
rect 84 5936 124 5968
rect 156 5936 196 5968
rect 228 5936 268 5968
rect 300 5936 340 5968
rect 372 5936 412 5968
rect 444 5936 484 5968
rect 516 5936 556 5968
rect 588 5936 628 5968
rect 660 5936 700 5968
rect 732 5936 772 5968
rect 804 5936 844 5968
rect 876 5936 916 5968
rect 948 5936 1000 5968
rect 0 5896 1000 5936
rect 0 5864 52 5896
rect 84 5864 124 5896
rect 156 5864 196 5896
rect 228 5864 268 5896
rect 300 5864 340 5896
rect 372 5864 412 5896
rect 444 5864 484 5896
rect 516 5864 556 5896
rect 588 5864 628 5896
rect 660 5864 700 5896
rect 732 5864 772 5896
rect 804 5864 844 5896
rect 876 5864 916 5896
rect 948 5864 1000 5896
rect 0 5824 1000 5864
rect 0 5792 52 5824
rect 84 5792 124 5824
rect 156 5792 196 5824
rect 228 5792 268 5824
rect 300 5792 340 5824
rect 372 5792 412 5824
rect 444 5792 484 5824
rect 516 5792 556 5824
rect 588 5792 628 5824
rect 660 5792 700 5824
rect 732 5792 772 5824
rect 804 5792 844 5824
rect 876 5792 916 5824
rect 948 5792 1000 5824
rect 0 5752 1000 5792
rect 0 5720 52 5752
rect 84 5720 124 5752
rect 156 5720 196 5752
rect 228 5720 268 5752
rect 300 5720 340 5752
rect 372 5720 412 5752
rect 444 5720 484 5752
rect 516 5720 556 5752
rect 588 5720 628 5752
rect 660 5720 700 5752
rect 732 5720 772 5752
rect 804 5720 844 5752
rect 876 5720 916 5752
rect 948 5720 1000 5752
rect 0 5680 1000 5720
rect 0 5648 52 5680
rect 84 5648 124 5680
rect 156 5648 196 5680
rect 228 5648 268 5680
rect 300 5648 340 5680
rect 372 5648 412 5680
rect 444 5648 484 5680
rect 516 5648 556 5680
rect 588 5648 628 5680
rect 660 5648 700 5680
rect 732 5648 772 5680
rect 804 5648 844 5680
rect 876 5648 916 5680
rect 948 5648 1000 5680
rect 0 5608 1000 5648
rect 0 5576 52 5608
rect 84 5576 124 5608
rect 156 5576 196 5608
rect 228 5576 268 5608
rect 300 5576 340 5608
rect 372 5576 412 5608
rect 444 5576 484 5608
rect 516 5576 556 5608
rect 588 5576 628 5608
rect 660 5576 700 5608
rect 732 5576 772 5608
rect 804 5576 844 5608
rect 876 5576 916 5608
rect 948 5576 1000 5608
rect 0 5536 1000 5576
rect 0 5504 52 5536
rect 84 5504 124 5536
rect 156 5504 196 5536
rect 228 5504 268 5536
rect 300 5504 340 5536
rect 372 5504 412 5536
rect 444 5504 484 5536
rect 516 5504 556 5536
rect 588 5504 628 5536
rect 660 5504 700 5536
rect 732 5504 772 5536
rect 804 5504 844 5536
rect 876 5504 916 5536
rect 948 5504 1000 5536
rect 0 5464 1000 5504
rect 0 5432 52 5464
rect 84 5432 124 5464
rect 156 5432 196 5464
rect 228 5432 268 5464
rect 300 5432 340 5464
rect 372 5432 412 5464
rect 444 5432 484 5464
rect 516 5432 556 5464
rect 588 5432 628 5464
rect 660 5432 700 5464
rect 732 5432 772 5464
rect 804 5432 844 5464
rect 876 5432 916 5464
rect 948 5432 1000 5464
rect 0 5392 1000 5432
rect 0 5360 52 5392
rect 84 5360 124 5392
rect 156 5360 196 5392
rect 228 5360 268 5392
rect 300 5360 340 5392
rect 372 5360 412 5392
rect 444 5360 484 5392
rect 516 5360 556 5392
rect 588 5360 628 5392
rect 660 5360 700 5392
rect 732 5360 772 5392
rect 804 5360 844 5392
rect 876 5360 916 5392
rect 948 5360 1000 5392
rect 0 5320 1000 5360
rect 0 5288 52 5320
rect 84 5288 124 5320
rect 156 5288 196 5320
rect 228 5288 268 5320
rect 300 5288 340 5320
rect 372 5288 412 5320
rect 444 5288 484 5320
rect 516 5288 556 5320
rect 588 5288 628 5320
rect 660 5288 700 5320
rect 732 5288 772 5320
rect 804 5288 844 5320
rect 876 5288 916 5320
rect 948 5288 1000 5320
rect 0 5248 1000 5288
rect 0 5216 52 5248
rect 84 5216 124 5248
rect 156 5216 196 5248
rect 228 5216 268 5248
rect 300 5216 340 5248
rect 372 5216 412 5248
rect 444 5216 484 5248
rect 516 5216 556 5248
rect 588 5216 628 5248
rect 660 5216 700 5248
rect 732 5216 772 5248
rect 804 5216 844 5248
rect 876 5216 916 5248
rect 948 5216 1000 5248
rect 0 5176 1000 5216
rect 0 5144 52 5176
rect 84 5144 124 5176
rect 156 5144 196 5176
rect 228 5144 268 5176
rect 300 5144 340 5176
rect 372 5144 412 5176
rect 444 5144 484 5176
rect 516 5144 556 5176
rect 588 5144 628 5176
rect 660 5144 700 5176
rect 732 5144 772 5176
rect 804 5144 844 5176
rect 876 5144 916 5176
rect 948 5144 1000 5176
rect 0 5104 1000 5144
rect 0 5072 52 5104
rect 84 5072 124 5104
rect 156 5072 196 5104
rect 228 5072 268 5104
rect 300 5072 340 5104
rect 372 5072 412 5104
rect 444 5072 484 5104
rect 516 5072 556 5104
rect 588 5072 628 5104
rect 660 5072 700 5104
rect 732 5072 772 5104
rect 804 5072 844 5104
rect 876 5072 916 5104
rect 948 5072 1000 5104
rect 0 5032 1000 5072
rect 0 5000 52 5032
rect 84 5000 124 5032
rect 156 5000 196 5032
rect 228 5000 268 5032
rect 300 5000 340 5032
rect 372 5000 412 5032
rect 444 5000 484 5032
rect 516 5000 556 5032
rect 588 5000 628 5032
rect 660 5000 700 5032
rect 732 5000 772 5032
rect 804 5000 844 5032
rect 876 5000 916 5032
rect 948 5000 1000 5032
rect 0 4960 1000 5000
rect 0 4928 52 4960
rect 84 4928 124 4960
rect 156 4928 196 4960
rect 228 4928 268 4960
rect 300 4928 340 4960
rect 372 4928 412 4960
rect 444 4928 484 4960
rect 516 4928 556 4960
rect 588 4928 628 4960
rect 660 4928 700 4960
rect 732 4928 772 4960
rect 804 4928 844 4960
rect 876 4928 916 4960
rect 948 4928 1000 4960
rect 0 4888 1000 4928
rect 0 4856 52 4888
rect 84 4856 124 4888
rect 156 4856 196 4888
rect 228 4856 268 4888
rect 300 4856 340 4888
rect 372 4856 412 4888
rect 444 4856 484 4888
rect 516 4856 556 4888
rect 588 4856 628 4888
rect 660 4856 700 4888
rect 732 4856 772 4888
rect 804 4856 844 4888
rect 876 4856 916 4888
rect 948 4856 1000 4888
rect 0 4816 1000 4856
rect 0 4784 52 4816
rect 84 4784 124 4816
rect 156 4784 196 4816
rect 228 4784 268 4816
rect 300 4784 340 4816
rect 372 4784 412 4816
rect 444 4784 484 4816
rect 516 4784 556 4816
rect 588 4784 628 4816
rect 660 4784 700 4816
rect 732 4784 772 4816
rect 804 4784 844 4816
rect 876 4784 916 4816
rect 948 4784 1000 4816
rect 0 4744 1000 4784
rect 0 4712 52 4744
rect 84 4712 124 4744
rect 156 4712 196 4744
rect 228 4712 268 4744
rect 300 4712 340 4744
rect 372 4712 412 4744
rect 444 4712 484 4744
rect 516 4712 556 4744
rect 588 4712 628 4744
rect 660 4712 700 4744
rect 732 4712 772 4744
rect 804 4712 844 4744
rect 876 4712 916 4744
rect 948 4712 1000 4744
rect 0 4672 1000 4712
rect 0 4640 52 4672
rect 84 4640 124 4672
rect 156 4640 196 4672
rect 228 4640 268 4672
rect 300 4640 340 4672
rect 372 4640 412 4672
rect 444 4640 484 4672
rect 516 4640 556 4672
rect 588 4640 628 4672
rect 660 4640 700 4672
rect 732 4640 772 4672
rect 804 4640 844 4672
rect 876 4640 916 4672
rect 948 4640 1000 4672
rect 0 4600 1000 4640
rect 0 4568 52 4600
rect 84 4568 124 4600
rect 156 4568 196 4600
rect 228 4568 268 4600
rect 300 4568 340 4600
rect 372 4568 412 4600
rect 444 4568 484 4600
rect 516 4568 556 4600
rect 588 4568 628 4600
rect 660 4568 700 4600
rect 732 4568 772 4600
rect 804 4568 844 4600
rect 876 4568 916 4600
rect 948 4568 1000 4600
rect 0 4528 1000 4568
rect 0 4496 52 4528
rect 84 4496 124 4528
rect 156 4496 196 4528
rect 228 4496 268 4528
rect 300 4496 340 4528
rect 372 4496 412 4528
rect 444 4496 484 4528
rect 516 4496 556 4528
rect 588 4496 628 4528
rect 660 4496 700 4528
rect 732 4496 772 4528
rect 804 4496 844 4528
rect 876 4496 916 4528
rect 948 4496 1000 4528
rect 0 4456 1000 4496
rect 0 4424 52 4456
rect 84 4424 124 4456
rect 156 4424 196 4456
rect 228 4424 268 4456
rect 300 4424 340 4456
rect 372 4424 412 4456
rect 444 4424 484 4456
rect 516 4424 556 4456
rect 588 4424 628 4456
rect 660 4424 700 4456
rect 732 4424 772 4456
rect 804 4424 844 4456
rect 876 4424 916 4456
rect 948 4424 1000 4456
rect 0 4384 1000 4424
rect 0 4352 52 4384
rect 84 4352 124 4384
rect 156 4352 196 4384
rect 228 4352 268 4384
rect 300 4352 340 4384
rect 372 4352 412 4384
rect 444 4352 484 4384
rect 516 4352 556 4384
rect 588 4352 628 4384
rect 660 4352 700 4384
rect 732 4352 772 4384
rect 804 4352 844 4384
rect 876 4352 916 4384
rect 948 4352 1000 4384
rect 0 4312 1000 4352
rect 0 4280 52 4312
rect 84 4280 124 4312
rect 156 4280 196 4312
rect 228 4280 268 4312
rect 300 4280 340 4312
rect 372 4280 412 4312
rect 444 4280 484 4312
rect 516 4280 556 4312
rect 588 4280 628 4312
rect 660 4280 700 4312
rect 732 4280 772 4312
rect 804 4280 844 4312
rect 876 4280 916 4312
rect 948 4280 1000 4312
rect 0 4240 1000 4280
rect 0 4208 52 4240
rect 84 4208 124 4240
rect 156 4208 196 4240
rect 228 4208 268 4240
rect 300 4208 340 4240
rect 372 4208 412 4240
rect 444 4208 484 4240
rect 516 4208 556 4240
rect 588 4208 628 4240
rect 660 4208 700 4240
rect 732 4208 772 4240
rect 804 4208 844 4240
rect 876 4208 916 4240
rect 948 4208 1000 4240
rect 0 4168 1000 4208
rect 0 4136 52 4168
rect 84 4136 124 4168
rect 156 4136 196 4168
rect 228 4136 268 4168
rect 300 4136 340 4168
rect 372 4136 412 4168
rect 444 4136 484 4168
rect 516 4136 556 4168
rect 588 4136 628 4168
rect 660 4136 700 4168
rect 732 4136 772 4168
rect 804 4136 844 4168
rect 876 4136 916 4168
rect 948 4136 1000 4168
rect 0 4096 1000 4136
rect 0 4064 52 4096
rect 84 4064 124 4096
rect 156 4064 196 4096
rect 228 4064 268 4096
rect 300 4064 340 4096
rect 372 4064 412 4096
rect 444 4064 484 4096
rect 516 4064 556 4096
rect 588 4064 628 4096
rect 660 4064 700 4096
rect 732 4064 772 4096
rect 804 4064 844 4096
rect 876 4064 916 4096
rect 948 4064 1000 4096
rect 0 4024 1000 4064
rect 0 3992 52 4024
rect 84 3992 124 4024
rect 156 3992 196 4024
rect 228 3992 268 4024
rect 300 3992 340 4024
rect 372 3992 412 4024
rect 444 3992 484 4024
rect 516 3992 556 4024
rect 588 3992 628 4024
rect 660 3992 700 4024
rect 732 3992 772 4024
rect 804 3992 844 4024
rect 876 3992 916 4024
rect 948 3992 1000 4024
rect 0 3952 1000 3992
rect 0 3920 52 3952
rect 84 3920 124 3952
rect 156 3920 196 3952
rect 228 3920 268 3952
rect 300 3920 340 3952
rect 372 3920 412 3952
rect 444 3920 484 3952
rect 516 3920 556 3952
rect 588 3920 628 3952
rect 660 3920 700 3952
rect 732 3920 772 3952
rect 804 3920 844 3952
rect 876 3920 916 3952
rect 948 3920 1000 3952
rect 0 3880 1000 3920
rect 0 3848 52 3880
rect 84 3848 124 3880
rect 156 3848 196 3880
rect 228 3848 268 3880
rect 300 3848 340 3880
rect 372 3848 412 3880
rect 444 3848 484 3880
rect 516 3848 556 3880
rect 588 3848 628 3880
rect 660 3848 700 3880
rect 732 3848 772 3880
rect 804 3848 844 3880
rect 876 3848 916 3880
rect 948 3848 1000 3880
rect 0 3808 1000 3848
rect 0 3776 52 3808
rect 84 3776 124 3808
rect 156 3776 196 3808
rect 228 3776 268 3808
rect 300 3776 340 3808
rect 372 3776 412 3808
rect 444 3776 484 3808
rect 516 3776 556 3808
rect 588 3776 628 3808
rect 660 3776 700 3808
rect 732 3776 772 3808
rect 804 3776 844 3808
rect 876 3776 916 3808
rect 948 3776 1000 3808
rect 0 3736 1000 3776
rect 0 3704 52 3736
rect 84 3704 124 3736
rect 156 3704 196 3736
rect 228 3704 268 3736
rect 300 3704 340 3736
rect 372 3704 412 3736
rect 444 3704 484 3736
rect 516 3704 556 3736
rect 588 3704 628 3736
rect 660 3704 700 3736
rect 732 3704 772 3736
rect 804 3704 844 3736
rect 876 3704 916 3736
rect 948 3704 1000 3736
rect 0 3664 1000 3704
rect 0 3632 52 3664
rect 84 3632 124 3664
rect 156 3632 196 3664
rect 228 3632 268 3664
rect 300 3632 340 3664
rect 372 3632 412 3664
rect 444 3632 484 3664
rect 516 3632 556 3664
rect 588 3632 628 3664
rect 660 3632 700 3664
rect 732 3632 772 3664
rect 804 3632 844 3664
rect 876 3632 916 3664
rect 948 3632 1000 3664
rect 0 3592 1000 3632
rect 0 3560 52 3592
rect 84 3560 124 3592
rect 156 3560 196 3592
rect 228 3560 268 3592
rect 300 3560 340 3592
rect 372 3560 412 3592
rect 444 3560 484 3592
rect 516 3560 556 3592
rect 588 3560 628 3592
rect 660 3560 700 3592
rect 732 3560 772 3592
rect 804 3560 844 3592
rect 876 3560 916 3592
rect 948 3560 1000 3592
rect 0 3520 1000 3560
rect 0 3488 52 3520
rect 84 3488 124 3520
rect 156 3488 196 3520
rect 228 3488 268 3520
rect 300 3488 340 3520
rect 372 3488 412 3520
rect 444 3488 484 3520
rect 516 3488 556 3520
rect 588 3488 628 3520
rect 660 3488 700 3520
rect 732 3488 772 3520
rect 804 3488 844 3520
rect 876 3488 916 3520
rect 948 3488 1000 3520
rect 0 3448 1000 3488
rect 0 3416 52 3448
rect 84 3416 124 3448
rect 156 3416 196 3448
rect 228 3416 268 3448
rect 300 3416 340 3448
rect 372 3416 412 3448
rect 444 3416 484 3448
rect 516 3416 556 3448
rect 588 3416 628 3448
rect 660 3416 700 3448
rect 732 3416 772 3448
rect 804 3416 844 3448
rect 876 3416 916 3448
rect 948 3416 1000 3448
rect 0 3376 1000 3416
rect 0 3344 52 3376
rect 84 3344 124 3376
rect 156 3344 196 3376
rect 228 3344 268 3376
rect 300 3344 340 3376
rect 372 3344 412 3376
rect 444 3344 484 3376
rect 516 3344 556 3376
rect 588 3344 628 3376
rect 660 3344 700 3376
rect 732 3344 772 3376
rect 804 3344 844 3376
rect 876 3344 916 3376
rect 948 3344 1000 3376
rect 0 3304 1000 3344
rect 0 3272 52 3304
rect 84 3272 124 3304
rect 156 3272 196 3304
rect 228 3272 268 3304
rect 300 3272 340 3304
rect 372 3272 412 3304
rect 444 3272 484 3304
rect 516 3272 556 3304
rect 588 3272 628 3304
rect 660 3272 700 3304
rect 732 3272 772 3304
rect 804 3272 844 3304
rect 876 3272 916 3304
rect 948 3272 1000 3304
rect 0 3232 1000 3272
rect 0 3200 52 3232
rect 84 3200 124 3232
rect 156 3200 196 3232
rect 228 3200 268 3232
rect 300 3200 340 3232
rect 372 3200 412 3232
rect 444 3200 484 3232
rect 516 3200 556 3232
rect 588 3200 628 3232
rect 660 3200 700 3232
rect 732 3200 772 3232
rect 804 3200 844 3232
rect 876 3200 916 3232
rect 948 3200 1000 3232
rect 0 3160 1000 3200
rect 0 3128 52 3160
rect 84 3128 124 3160
rect 156 3128 196 3160
rect 228 3128 268 3160
rect 300 3128 340 3160
rect 372 3128 412 3160
rect 444 3128 484 3160
rect 516 3128 556 3160
rect 588 3128 628 3160
rect 660 3128 700 3160
rect 732 3128 772 3160
rect 804 3128 844 3160
rect 876 3128 916 3160
rect 948 3128 1000 3160
rect 0 3088 1000 3128
rect 0 3056 52 3088
rect 84 3056 124 3088
rect 156 3056 196 3088
rect 228 3056 268 3088
rect 300 3056 340 3088
rect 372 3056 412 3088
rect 444 3056 484 3088
rect 516 3056 556 3088
rect 588 3056 628 3088
rect 660 3056 700 3088
rect 732 3056 772 3088
rect 804 3056 844 3088
rect 876 3056 916 3088
rect 948 3056 1000 3088
rect 0 3016 1000 3056
rect 0 2984 52 3016
rect 84 2984 124 3016
rect 156 2984 196 3016
rect 228 2984 268 3016
rect 300 2984 340 3016
rect 372 2984 412 3016
rect 444 2984 484 3016
rect 516 2984 556 3016
rect 588 2984 628 3016
rect 660 2984 700 3016
rect 732 2984 772 3016
rect 804 2984 844 3016
rect 876 2984 916 3016
rect 948 2984 1000 3016
rect 0 2944 1000 2984
rect 0 2912 52 2944
rect 84 2912 124 2944
rect 156 2912 196 2944
rect 228 2912 268 2944
rect 300 2912 340 2944
rect 372 2912 412 2944
rect 444 2912 484 2944
rect 516 2912 556 2944
rect 588 2912 628 2944
rect 660 2912 700 2944
rect 732 2912 772 2944
rect 804 2912 844 2944
rect 876 2912 916 2944
rect 948 2912 1000 2944
rect 0 2872 1000 2912
rect 0 2840 52 2872
rect 84 2840 124 2872
rect 156 2840 196 2872
rect 228 2840 268 2872
rect 300 2840 340 2872
rect 372 2840 412 2872
rect 444 2840 484 2872
rect 516 2840 556 2872
rect 588 2840 628 2872
rect 660 2840 700 2872
rect 732 2840 772 2872
rect 804 2840 844 2872
rect 876 2840 916 2872
rect 948 2840 1000 2872
rect 0 2800 1000 2840
rect 0 2768 52 2800
rect 84 2768 124 2800
rect 156 2768 196 2800
rect 228 2768 268 2800
rect 300 2768 340 2800
rect 372 2768 412 2800
rect 444 2768 484 2800
rect 516 2768 556 2800
rect 588 2768 628 2800
rect 660 2768 700 2800
rect 732 2768 772 2800
rect 804 2768 844 2800
rect 876 2768 916 2800
rect 948 2768 1000 2800
rect 0 2728 1000 2768
rect 0 2696 52 2728
rect 84 2696 124 2728
rect 156 2696 196 2728
rect 228 2696 268 2728
rect 300 2696 340 2728
rect 372 2696 412 2728
rect 444 2696 484 2728
rect 516 2696 556 2728
rect 588 2696 628 2728
rect 660 2696 700 2728
rect 732 2696 772 2728
rect 804 2696 844 2728
rect 876 2696 916 2728
rect 948 2696 1000 2728
rect 0 2656 1000 2696
rect 0 2624 52 2656
rect 84 2624 124 2656
rect 156 2624 196 2656
rect 228 2624 268 2656
rect 300 2624 340 2656
rect 372 2624 412 2656
rect 444 2624 484 2656
rect 516 2624 556 2656
rect 588 2624 628 2656
rect 660 2624 700 2656
rect 732 2624 772 2656
rect 804 2624 844 2656
rect 876 2624 916 2656
rect 948 2624 1000 2656
rect 0 2584 1000 2624
rect 0 2552 52 2584
rect 84 2552 124 2584
rect 156 2552 196 2584
rect 228 2552 268 2584
rect 300 2552 340 2584
rect 372 2552 412 2584
rect 444 2552 484 2584
rect 516 2552 556 2584
rect 588 2552 628 2584
rect 660 2552 700 2584
rect 732 2552 772 2584
rect 804 2552 844 2584
rect 876 2552 916 2584
rect 948 2552 1000 2584
rect 0 2512 1000 2552
rect 0 2480 52 2512
rect 84 2480 124 2512
rect 156 2480 196 2512
rect 228 2480 268 2512
rect 300 2480 340 2512
rect 372 2480 412 2512
rect 444 2480 484 2512
rect 516 2480 556 2512
rect 588 2480 628 2512
rect 660 2480 700 2512
rect 732 2480 772 2512
rect 804 2480 844 2512
rect 876 2480 916 2512
rect 948 2480 1000 2512
rect 0 2440 1000 2480
rect 0 2408 52 2440
rect 84 2408 124 2440
rect 156 2408 196 2440
rect 228 2408 268 2440
rect 300 2408 340 2440
rect 372 2408 412 2440
rect 444 2408 484 2440
rect 516 2408 556 2440
rect 588 2408 628 2440
rect 660 2408 700 2440
rect 732 2408 772 2440
rect 804 2408 844 2440
rect 876 2408 916 2440
rect 948 2408 1000 2440
rect 0 2368 1000 2408
rect 0 2336 52 2368
rect 84 2336 124 2368
rect 156 2336 196 2368
rect 228 2336 268 2368
rect 300 2336 340 2368
rect 372 2336 412 2368
rect 444 2336 484 2368
rect 516 2336 556 2368
rect 588 2336 628 2368
rect 660 2336 700 2368
rect 732 2336 772 2368
rect 804 2336 844 2368
rect 876 2336 916 2368
rect 948 2336 1000 2368
rect 0 2296 1000 2336
rect 0 2264 52 2296
rect 84 2264 124 2296
rect 156 2264 196 2296
rect 228 2264 268 2296
rect 300 2264 340 2296
rect 372 2264 412 2296
rect 444 2264 484 2296
rect 516 2264 556 2296
rect 588 2264 628 2296
rect 660 2264 700 2296
rect 732 2264 772 2296
rect 804 2264 844 2296
rect 876 2264 916 2296
rect 948 2264 1000 2296
rect 0 2224 1000 2264
rect 0 2192 52 2224
rect 84 2192 124 2224
rect 156 2192 196 2224
rect 228 2192 268 2224
rect 300 2192 340 2224
rect 372 2192 412 2224
rect 444 2192 484 2224
rect 516 2192 556 2224
rect 588 2192 628 2224
rect 660 2192 700 2224
rect 732 2192 772 2224
rect 804 2192 844 2224
rect 876 2192 916 2224
rect 948 2192 1000 2224
rect 0 2152 1000 2192
rect 0 2120 52 2152
rect 84 2120 124 2152
rect 156 2120 196 2152
rect 228 2120 268 2152
rect 300 2120 340 2152
rect 372 2120 412 2152
rect 444 2120 484 2152
rect 516 2120 556 2152
rect 588 2120 628 2152
rect 660 2120 700 2152
rect 732 2120 772 2152
rect 804 2120 844 2152
rect 876 2120 916 2152
rect 948 2120 1000 2152
rect 0 2080 1000 2120
rect 0 2048 52 2080
rect 84 2048 124 2080
rect 156 2048 196 2080
rect 228 2048 268 2080
rect 300 2048 340 2080
rect 372 2048 412 2080
rect 444 2048 484 2080
rect 516 2048 556 2080
rect 588 2048 628 2080
rect 660 2048 700 2080
rect 732 2048 772 2080
rect 804 2048 844 2080
rect 876 2048 916 2080
rect 948 2048 1000 2080
rect 0 2008 1000 2048
rect 0 1976 52 2008
rect 84 1976 124 2008
rect 156 1976 196 2008
rect 228 1976 268 2008
rect 300 1976 340 2008
rect 372 1976 412 2008
rect 444 1976 484 2008
rect 516 1976 556 2008
rect 588 1976 628 2008
rect 660 1976 700 2008
rect 732 1976 772 2008
rect 804 1976 844 2008
rect 876 1976 916 2008
rect 948 1976 1000 2008
rect 0 1936 1000 1976
rect 0 1904 52 1936
rect 84 1904 124 1936
rect 156 1904 196 1936
rect 228 1904 268 1936
rect 300 1904 340 1936
rect 372 1904 412 1936
rect 444 1904 484 1936
rect 516 1904 556 1936
rect 588 1904 628 1936
rect 660 1904 700 1936
rect 732 1904 772 1936
rect 804 1904 844 1936
rect 876 1904 916 1936
rect 948 1904 1000 1936
rect 0 1864 1000 1904
rect 0 1832 52 1864
rect 84 1832 124 1864
rect 156 1832 196 1864
rect 228 1832 268 1864
rect 300 1832 340 1864
rect 372 1832 412 1864
rect 444 1832 484 1864
rect 516 1832 556 1864
rect 588 1832 628 1864
rect 660 1832 700 1864
rect 732 1832 772 1864
rect 804 1832 844 1864
rect 876 1832 916 1864
rect 948 1832 1000 1864
rect 0 1792 1000 1832
rect 0 1760 52 1792
rect 84 1760 124 1792
rect 156 1760 196 1792
rect 228 1760 268 1792
rect 300 1760 340 1792
rect 372 1760 412 1792
rect 444 1760 484 1792
rect 516 1760 556 1792
rect 588 1760 628 1792
rect 660 1760 700 1792
rect 732 1760 772 1792
rect 804 1760 844 1792
rect 876 1760 916 1792
rect 948 1760 1000 1792
rect 0 1720 1000 1760
rect 0 1688 52 1720
rect 84 1688 124 1720
rect 156 1688 196 1720
rect 228 1688 268 1720
rect 300 1688 340 1720
rect 372 1688 412 1720
rect 444 1688 484 1720
rect 516 1688 556 1720
rect 588 1688 628 1720
rect 660 1688 700 1720
rect 732 1688 772 1720
rect 804 1688 844 1720
rect 876 1688 916 1720
rect 948 1688 1000 1720
rect 0 1648 1000 1688
rect 0 1616 52 1648
rect 84 1616 124 1648
rect 156 1616 196 1648
rect 228 1616 268 1648
rect 300 1616 340 1648
rect 372 1616 412 1648
rect 444 1616 484 1648
rect 516 1616 556 1648
rect 588 1616 628 1648
rect 660 1616 700 1648
rect 732 1616 772 1648
rect 804 1616 844 1648
rect 876 1616 916 1648
rect 948 1616 1000 1648
rect 0 1576 1000 1616
rect 0 1544 52 1576
rect 84 1544 124 1576
rect 156 1544 196 1576
rect 228 1544 268 1576
rect 300 1544 340 1576
rect 372 1544 412 1576
rect 444 1544 484 1576
rect 516 1544 556 1576
rect 588 1544 628 1576
rect 660 1544 700 1576
rect 732 1544 772 1576
rect 804 1544 844 1576
rect 876 1544 916 1576
rect 948 1544 1000 1576
rect 0 1504 1000 1544
rect 0 1472 52 1504
rect 84 1472 124 1504
rect 156 1472 196 1504
rect 228 1472 268 1504
rect 300 1472 340 1504
rect 372 1472 412 1504
rect 444 1472 484 1504
rect 516 1472 556 1504
rect 588 1472 628 1504
rect 660 1472 700 1504
rect 732 1472 772 1504
rect 804 1472 844 1504
rect 876 1472 916 1504
rect 948 1472 1000 1504
rect 0 1432 1000 1472
rect 0 1400 52 1432
rect 84 1400 124 1432
rect 156 1400 196 1432
rect 228 1400 268 1432
rect 300 1400 340 1432
rect 372 1400 412 1432
rect 444 1400 484 1432
rect 516 1400 556 1432
rect 588 1400 628 1432
rect 660 1400 700 1432
rect 732 1400 772 1432
rect 804 1400 844 1432
rect 876 1400 916 1432
rect 948 1400 1000 1432
rect 0 1360 1000 1400
rect 0 1328 52 1360
rect 84 1328 124 1360
rect 156 1328 196 1360
rect 228 1328 268 1360
rect 300 1328 340 1360
rect 372 1328 412 1360
rect 444 1328 484 1360
rect 516 1328 556 1360
rect 588 1328 628 1360
rect 660 1328 700 1360
rect 732 1328 772 1360
rect 804 1328 844 1360
rect 876 1328 916 1360
rect 948 1328 1000 1360
rect 0 1288 1000 1328
rect 0 1256 52 1288
rect 84 1256 124 1288
rect 156 1256 196 1288
rect 228 1256 268 1288
rect 300 1256 340 1288
rect 372 1256 412 1288
rect 444 1256 484 1288
rect 516 1256 556 1288
rect 588 1256 628 1288
rect 660 1256 700 1288
rect 732 1256 772 1288
rect 804 1256 844 1288
rect 876 1256 916 1288
rect 948 1256 1000 1288
rect 0 1200 1000 1256
<< psubdiffcont >>
rect 223 31384 255 31416
rect 124 27939 156 27971
rect 124 22842 156 22874
rect 124 17816 156 17848
<< nsubdiffcont >>
rect 124 33384 156 33416
rect 124 29684 156 29716
rect 52 12112 84 12144
rect 52 6512 84 6544
<< metal1 >>
rect 196 33384 228 33416
rect 268 33384 300 33416
rect 340 33384 372 33416
rect 412 33384 444 33416
rect 484 33384 516 33416
rect 556 33384 588 33416
rect 628 33384 660 33416
rect 700 33384 732 33416
rect 772 33384 804 33416
rect 844 33384 876 33416
rect 196 29684 228 29716
rect 268 29684 300 29716
rect 340 29684 372 29716
rect 412 29684 444 29716
rect 484 29684 516 29716
rect 556 29684 588 29716
rect 628 29684 660 29716
rect 700 29684 732 29716
rect 772 29684 804 29716
rect 844 29684 876 29716
rect 124 12112 156 12144
rect 196 12112 228 12144
rect 268 12112 300 12144
rect 340 12112 372 12144
rect 412 12112 444 12144
rect 484 12112 516 12144
rect 556 12112 588 12144
rect 628 12112 660 12144
rect 700 12112 732 12144
rect 772 12112 804 12144
rect 844 12112 876 12144
rect 916 12112 948 12144
rect 52 12040 84 12072
rect 124 12040 156 12072
rect 196 12040 228 12072
rect 268 12040 300 12072
rect 340 12040 372 12072
rect 412 12040 444 12072
rect 484 12040 516 12072
rect 556 12040 588 12072
rect 628 12040 660 12072
rect 700 12040 732 12072
rect 772 12040 804 12072
rect 844 12040 876 12072
rect 916 12040 948 12072
rect 52 11968 84 12000
rect 124 11968 156 12000
rect 196 11968 228 12000
rect 268 11968 300 12000
rect 340 11968 372 12000
rect 412 11968 444 12000
rect 484 11968 516 12000
rect 556 11968 588 12000
rect 628 11968 660 12000
rect 700 11968 732 12000
rect 772 11968 804 12000
rect 844 11968 876 12000
rect 916 11968 948 12000
rect 52 11896 84 11928
rect 124 11896 156 11928
rect 196 11896 228 11928
rect 268 11896 300 11928
rect 340 11896 372 11928
rect 412 11896 444 11928
rect 484 11896 516 11928
rect 556 11896 588 11928
rect 628 11896 660 11928
rect 700 11896 732 11928
rect 772 11896 804 11928
rect 844 11896 876 11928
rect 916 11896 948 11928
rect 52 11824 84 11856
rect 124 11824 156 11856
rect 196 11824 228 11856
rect 268 11824 300 11856
rect 340 11824 372 11856
rect 412 11824 444 11856
rect 484 11824 516 11856
rect 556 11824 588 11856
rect 628 11824 660 11856
rect 700 11824 732 11856
rect 772 11824 804 11856
rect 844 11824 876 11856
rect 916 11824 948 11856
rect 52 11752 84 11784
rect 124 11752 156 11784
rect 196 11752 228 11784
rect 268 11752 300 11784
rect 340 11752 372 11784
rect 412 11752 444 11784
rect 484 11752 516 11784
rect 556 11752 588 11784
rect 628 11752 660 11784
rect 700 11752 732 11784
rect 772 11752 804 11784
rect 844 11752 876 11784
rect 916 11752 948 11784
rect 52 11680 84 11712
rect 124 11680 156 11712
rect 196 11680 228 11712
rect 268 11680 300 11712
rect 340 11680 372 11712
rect 412 11680 444 11712
rect 484 11680 516 11712
rect 556 11680 588 11712
rect 628 11680 660 11712
rect 700 11680 732 11712
rect 772 11680 804 11712
rect 844 11680 876 11712
rect 916 11680 948 11712
rect 52 11608 84 11640
rect 124 11608 156 11640
rect 196 11608 228 11640
rect 268 11608 300 11640
rect 340 11608 372 11640
rect 412 11608 444 11640
rect 484 11608 516 11640
rect 556 11608 588 11640
rect 628 11608 660 11640
rect 700 11608 732 11640
rect 772 11608 804 11640
rect 844 11608 876 11640
rect 916 11608 948 11640
rect 52 11536 84 11568
rect 124 11536 156 11568
rect 196 11536 228 11568
rect 268 11536 300 11568
rect 340 11536 372 11568
rect 412 11536 444 11568
rect 484 11536 516 11568
rect 556 11536 588 11568
rect 628 11536 660 11568
rect 700 11536 732 11568
rect 772 11536 804 11568
rect 844 11536 876 11568
rect 916 11536 948 11568
rect 52 11464 84 11496
rect 124 11464 156 11496
rect 196 11464 228 11496
rect 268 11464 300 11496
rect 340 11464 372 11496
rect 412 11464 444 11496
rect 484 11464 516 11496
rect 556 11464 588 11496
rect 628 11464 660 11496
rect 700 11464 732 11496
rect 772 11464 804 11496
rect 844 11464 876 11496
rect 916 11464 948 11496
rect 52 11392 84 11424
rect 124 11392 156 11424
rect 196 11392 228 11424
rect 268 11392 300 11424
rect 340 11392 372 11424
rect 412 11392 444 11424
rect 484 11392 516 11424
rect 556 11392 588 11424
rect 628 11392 660 11424
rect 700 11392 732 11424
rect 772 11392 804 11424
rect 844 11392 876 11424
rect 916 11392 948 11424
rect 52 11320 84 11352
rect 124 11320 156 11352
rect 196 11320 228 11352
rect 268 11320 300 11352
rect 340 11320 372 11352
rect 412 11320 444 11352
rect 484 11320 516 11352
rect 556 11320 588 11352
rect 628 11320 660 11352
rect 700 11320 732 11352
rect 772 11320 804 11352
rect 844 11320 876 11352
rect 916 11320 948 11352
rect 52 11248 84 11280
rect 124 11248 156 11280
rect 196 11248 228 11280
rect 268 11248 300 11280
rect 340 11248 372 11280
rect 412 11248 444 11280
rect 484 11248 516 11280
rect 556 11248 588 11280
rect 628 11248 660 11280
rect 700 11248 732 11280
rect 772 11248 804 11280
rect 844 11248 876 11280
rect 916 11248 948 11280
rect 52 11176 84 11208
rect 124 11176 156 11208
rect 196 11176 228 11208
rect 268 11176 300 11208
rect 340 11176 372 11208
rect 412 11176 444 11208
rect 484 11176 516 11208
rect 556 11176 588 11208
rect 628 11176 660 11208
rect 700 11176 732 11208
rect 772 11176 804 11208
rect 844 11176 876 11208
rect 916 11176 948 11208
rect 52 11104 84 11136
rect 124 11104 156 11136
rect 196 11104 228 11136
rect 268 11104 300 11136
rect 340 11104 372 11136
rect 412 11104 444 11136
rect 484 11104 516 11136
rect 556 11104 588 11136
rect 628 11104 660 11136
rect 700 11104 732 11136
rect 772 11104 804 11136
rect 844 11104 876 11136
rect 916 11104 948 11136
rect 52 11032 84 11064
rect 124 11032 156 11064
rect 196 11032 228 11064
rect 268 11032 300 11064
rect 340 11032 372 11064
rect 412 11032 444 11064
rect 484 11032 516 11064
rect 556 11032 588 11064
rect 628 11032 660 11064
rect 700 11032 732 11064
rect 772 11032 804 11064
rect 844 11032 876 11064
rect 916 11032 948 11064
rect 52 10960 84 10992
rect 124 10960 156 10992
rect 196 10960 228 10992
rect 268 10960 300 10992
rect 340 10960 372 10992
rect 412 10960 444 10992
rect 484 10960 516 10992
rect 556 10960 588 10992
rect 628 10960 660 10992
rect 700 10960 732 10992
rect 772 10960 804 10992
rect 844 10960 876 10992
rect 916 10960 948 10992
rect 52 10888 84 10920
rect 124 10888 156 10920
rect 196 10888 228 10920
rect 268 10888 300 10920
rect 340 10888 372 10920
rect 412 10888 444 10920
rect 484 10888 516 10920
rect 556 10888 588 10920
rect 628 10888 660 10920
rect 700 10888 732 10920
rect 772 10888 804 10920
rect 844 10888 876 10920
rect 916 10888 948 10920
rect 52 10816 84 10848
rect 124 10816 156 10848
rect 196 10816 228 10848
rect 268 10816 300 10848
rect 340 10816 372 10848
rect 412 10816 444 10848
rect 484 10816 516 10848
rect 556 10816 588 10848
rect 628 10816 660 10848
rect 700 10816 732 10848
rect 772 10816 804 10848
rect 844 10816 876 10848
rect 916 10816 948 10848
rect 52 10744 84 10776
rect 124 10744 156 10776
rect 196 10744 228 10776
rect 268 10744 300 10776
rect 340 10744 372 10776
rect 412 10744 444 10776
rect 484 10744 516 10776
rect 556 10744 588 10776
rect 628 10744 660 10776
rect 700 10744 732 10776
rect 772 10744 804 10776
rect 844 10744 876 10776
rect 916 10744 948 10776
rect 52 10672 84 10704
rect 124 10672 156 10704
rect 196 10672 228 10704
rect 268 10672 300 10704
rect 340 10672 372 10704
rect 412 10672 444 10704
rect 484 10672 516 10704
rect 556 10672 588 10704
rect 628 10672 660 10704
rect 700 10672 732 10704
rect 772 10672 804 10704
rect 844 10672 876 10704
rect 916 10672 948 10704
rect 52 10600 84 10632
rect 124 10600 156 10632
rect 196 10600 228 10632
rect 268 10600 300 10632
rect 340 10600 372 10632
rect 412 10600 444 10632
rect 484 10600 516 10632
rect 556 10600 588 10632
rect 628 10600 660 10632
rect 700 10600 732 10632
rect 772 10600 804 10632
rect 844 10600 876 10632
rect 916 10600 948 10632
rect 52 10528 84 10560
rect 124 10528 156 10560
rect 196 10528 228 10560
rect 268 10528 300 10560
rect 340 10528 372 10560
rect 412 10528 444 10560
rect 484 10528 516 10560
rect 556 10528 588 10560
rect 628 10528 660 10560
rect 700 10528 732 10560
rect 772 10528 804 10560
rect 844 10528 876 10560
rect 916 10528 948 10560
rect 52 10456 84 10488
rect 124 10456 156 10488
rect 196 10456 228 10488
rect 268 10456 300 10488
rect 340 10456 372 10488
rect 412 10456 444 10488
rect 484 10456 516 10488
rect 556 10456 588 10488
rect 628 10456 660 10488
rect 700 10456 732 10488
rect 772 10456 804 10488
rect 844 10456 876 10488
rect 916 10456 948 10488
rect 52 10384 84 10416
rect 124 10384 156 10416
rect 196 10384 228 10416
rect 268 10384 300 10416
rect 340 10384 372 10416
rect 412 10384 444 10416
rect 484 10384 516 10416
rect 556 10384 588 10416
rect 628 10384 660 10416
rect 700 10384 732 10416
rect 772 10384 804 10416
rect 844 10384 876 10416
rect 916 10384 948 10416
rect 52 10312 84 10344
rect 124 10312 156 10344
rect 196 10312 228 10344
rect 268 10312 300 10344
rect 340 10312 372 10344
rect 412 10312 444 10344
rect 484 10312 516 10344
rect 556 10312 588 10344
rect 628 10312 660 10344
rect 700 10312 732 10344
rect 772 10312 804 10344
rect 844 10312 876 10344
rect 916 10312 948 10344
rect 52 10240 84 10272
rect 124 10240 156 10272
rect 196 10240 228 10272
rect 268 10240 300 10272
rect 340 10240 372 10272
rect 412 10240 444 10272
rect 484 10240 516 10272
rect 556 10240 588 10272
rect 628 10240 660 10272
rect 700 10240 732 10272
rect 772 10240 804 10272
rect 844 10240 876 10272
rect 916 10240 948 10272
rect 52 10168 84 10200
rect 124 10168 156 10200
rect 196 10168 228 10200
rect 268 10168 300 10200
rect 340 10168 372 10200
rect 412 10168 444 10200
rect 484 10168 516 10200
rect 556 10168 588 10200
rect 628 10168 660 10200
rect 700 10168 732 10200
rect 772 10168 804 10200
rect 844 10168 876 10200
rect 916 10168 948 10200
rect 52 10096 84 10128
rect 124 10096 156 10128
rect 196 10096 228 10128
rect 268 10096 300 10128
rect 340 10096 372 10128
rect 412 10096 444 10128
rect 484 10096 516 10128
rect 556 10096 588 10128
rect 628 10096 660 10128
rect 700 10096 732 10128
rect 772 10096 804 10128
rect 844 10096 876 10128
rect 916 10096 948 10128
rect 52 10024 84 10056
rect 124 10024 156 10056
rect 196 10024 228 10056
rect 268 10024 300 10056
rect 340 10024 372 10056
rect 412 10024 444 10056
rect 484 10024 516 10056
rect 556 10024 588 10056
rect 628 10024 660 10056
rect 700 10024 732 10056
rect 772 10024 804 10056
rect 844 10024 876 10056
rect 916 10024 948 10056
rect 52 9952 84 9984
rect 124 9952 156 9984
rect 196 9952 228 9984
rect 268 9952 300 9984
rect 340 9952 372 9984
rect 412 9952 444 9984
rect 484 9952 516 9984
rect 556 9952 588 9984
rect 628 9952 660 9984
rect 700 9952 732 9984
rect 772 9952 804 9984
rect 844 9952 876 9984
rect 916 9952 948 9984
rect 52 9880 84 9912
rect 124 9880 156 9912
rect 196 9880 228 9912
rect 268 9880 300 9912
rect 340 9880 372 9912
rect 412 9880 444 9912
rect 484 9880 516 9912
rect 556 9880 588 9912
rect 628 9880 660 9912
rect 700 9880 732 9912
rect 772 9880 804 9912
rect 844 9880 876 9912
rect 916 9880 948 9912
rect 52 9808 84 9840
rect 124 9808 156 9840
rect 196 9808 228 9840
rect 268 9808 300 9840
rect 340 9808 372 9840
rect 412 9808 444 9840
rect 484 9808 516 9840
rect 556 9808 588 9840
rect 628 9808 660 9840
rect 700 9808 732 9840
rect 772 9808 804 9840
rect 844 9808 876 9840
rect 916 9808 948 9840
rect 52 9736 84 9768
rect 124 9736 156 9768
rect 196 9736 228 9768
rect 268 9736 300 9768
rect 340 9736 372 9768
rect 412 9736 444 9768
rect 484 9736 516 9768
rect 556 9736 588 9768
rect 628 9736 660 9768
rect 700 9736 732 9768
rect 772 9736 804 9768
rect 844 9736 876 9768
rect 916 9736 948 9768
rect 52 9664 84 9696
rect 124 9664 156 9696
rect 196 9664 228 9696
rect 268 9664 300 9696
rect 340 9664 372 9696
rect 412 9664 444 9696
rect 484 9664 516 9696
rect 556 9664 588 9696
rect 628 9664 660 9696
rect 700 9664 732 9696
rect 772 9664 804 9696
rect 844 9664 876 9696
rect 916 9664 948 9696
rect 52 9592 84 9624
rect 124 9592 156 9624
rect 196 9592 228 9624
rect 268 9592 300 9624
rect 340 9592 372 9624
rect 412 9592 444 9624
rect 484 9592 516 9624
rect 556 9592 588 9624
rect 628 9592 660 9624
rect 700 9592 732 9624
rect 772 9592 804 9624
rect 844 9592 876 9624
rect 916 9592 948 9624
rect 52 9520 84 9552
rect 124 9520 156 9552
rect 196 9520 228 9552
rect 268 9520 300 9552
rect 340 9520 372 9552
rect 412 9520 444 9552
rect 484 9520 516 9552
rect 556 9520 588 9552
rect 628 9520 660 9552
rect 700 9520 732 9552
rect 772 9520 804 9552
rect 844 9520 876 9552
rect 916 9520 948 9552
rect 52 9448 84 9480
rect 124 9448 156 9480
rect 196 9448 228 9480
rect 268 9448 300 9480
rect 340 9448 372 9480
rect 412 9448 444 9480
rect 484 9448 516 9480
rect 556 9448 588 9480
rect 628 9448 660 9480
rect 700 9448 732 9480
rect 772 9448 804 9480
rect 844 9448 876 9480
rect 916 9448 948 9480
rect 52 9376 84 9408
rect 124 9376 156 9408
rect 196 9376 228 9408
rect 268 9376 300 9408
rect 340 9376 372 9408
rect 412 9376 444 9408
rect 484 9376 516 9408
rect 556 9376 588 9408
rect 628 9376 660 9408
rect 700 9376 732 9408
rect 772 9376 804 9408
rect 844 9376 876 9408
rect 916 9376 948 9408
rect 52 9304 84 9336
rect 124 9304 156 9336
rect 196 9304 228 9336
rect 268 9304 300 9336
rect 340 9304 372 9336
rect 412 9304 444 9336
rect 484 9304 516 9336
rect 556 9304 588 9336
rect 628 9304 660 9336
rect 700 9304 732 9336
rect 772 9304 804 9336
rect 844 9304 876 9336
rect 916 9304 948 9336
rect 52 9232 84 9264
rect 124 9232 156 9264
rect 196 9232 228 9264
rect 268 9232 300 9264
rect 340 9232 372 9264
rect 412 9232 444 9264
rect 484 9232 516 9264
rect 556 9232 588 9264
rect 628 9232 660 9264
rect 700 9232 732 9264
rect 772 9232 804 9264
rect 844 9232 876 9264
rect 916 9232 948 9264
rect 52 9160 84 9192
rect 124 9160 156 9192
rect 196 9160 228 9192
rect 268 9160 300 9192
rect 340 9160 372 9192
rect 412 9160 444 9192
rect 484 9160 516 9192
rect 556 9160 588 9192
rect 628 9160 660 9192
rect 700 9160 732 9192
rect 772 9160 804 9192
rect 844 9160 876 9192
rect 916 9160 948 9192
rect 52 9088 84 9120
rect 124 9088 156 9120
rect 196 9088 228 9120
rect 268 9088 300 9120
rect 340 9088 372 9120
rect 412 9088 444 9120
rect 484 9088 516 9120
rect 556 9088 588 9120
rect 628 9088 660 9120
rect 700 9088 732 9120
rect 772 9088 804 9120
rect 844 9088 876 9120
rect 916 9088 948 9120
rect 52 9016 84 9048
rect 124 9016 156 9048
rect 196 9016 228 9048
rect 268 9016 300 9048
rect 340 9016 372 9048
rect 412 9016 444 9048
rect 484 9016 516 9048
rect 556 9016 588 9048
rect 628 9016 660 9048
rect 700 9016 732 9048
rect 772 9016 804 9048
rect 844 9016 876 9048
rect 916 9016 948 9048
rect 52 8944 84 8976
rect 124 8944 156 8976
rect 196 8944 228 8976
rect 268 8944 300 8976
rect 340 8944 372 8976
rect 412 8944 444 8976
rect 484 8944 516 8976
rect 556 8944 588 8976
rect 628 8944 660 8976
rect 700 8944 732 8976
rect 772 8944 804 8976
rect 844 8944 876 8976
rect 916 8944 948 8976
rect 52 8872 84 8904
rect 124 8872 156 8904
rect 196 8872 228 8904
rect 268 8872 300 8904
rect 340 8872 372 8904
rect 412 8872 444 8904
rect 484 8872 516 8904
rect 556 8872 588 8904
rect 628 8872 660 8904
rect 700 8872 732 8904
rect 772 8872 804 8904
rect 844 8872 876 8904
rect 916 8872 948 8904
rect 52 8800 84 8832
rect 124 8800 156 8832
rect 196 8800 228 8832
rect 268 8800 300 8832
rect 340 8800 372 8832
rect 412 8800 444 8832
rect 484 8800 516 8832
rect 556 8800 588 8832
rect 628 8800 660 8832
rect 700 8800 732 8832
rect 772 8800 804 8832
rect 844 8800 876 8832
rect 916 8800 948 8832
rect 52 8728 84 8760
rect 124 8728 156 8760
rect 196 8728 228 8760
rect 268 8728 300 8760
rect 340 8728 372 8760
rect 412 8728 444 8760
rect 484 8728 516 8760
rect 556 8728 588 8760
rect 628 8728 660 8760
rect 700 8728 732 8760
rect 772 8728 804 8760
rect 844 8728 876 8760
rect 916 8728 948 8760
rect 52 8656 84 8688
rect 124 8656 156 8688
rect 196 8656 228 8688
rect 268 8656 300 8688
rect 340 8656 372 8688
rect 412 8656 444 8688
rect 484 8656 516 8688
rect 556 8656 588 8688
rect 628 8656 660 8688
rect 700 8656 732 8688
rect 772 8656 804 8688
rect 844 8656 876 8688
rect 916 8656 948 8688
rect 52 8584 84 8616
rect 124 8584 156 8616
rect 196 8584 228 8616
rect 268 8584 300 8616
rect 340 8584 372 8616
rect 412 8584 444 8616
rect 484 8584 516 8616
rect 556 8584 588 8616
rect 628 8584 660 8616
rect 700 8584 732 8616
rect 772 8584 804 8616
rect 844 8584 876 8616
rect 916 8584 948 8616
rect 52 8512 84 8544
rect 124 8512 156 8544
rect 196 8512 228 8544
rect 268 8512 300 8544
rect 340 8512 372 8544
rect 412 8512 444 8544
rect 484 8512 516 8544
rect 556 8512 588 8544
rect 628 8512 660 8544
rect 700 8512 732 8544
rect 772 8512 804 8544
rect 844 8512 876 8544
rect 916 8512 948 8544
rect 52 8440 84 8472
rect 124 8440 156 8472
rect 196 8440 228 8472
rect 268 8440 300 8472
rect 340 8440 372 8472
rect 412 8440 444 8472
rect 484 8440 516 8472
rect 556 8440 588 8472
rect 628 8440 660 8472
rect 700 8440 732 8472
rect 772 8440 804 8472
rect 844 8440 876 8472
rect 916 8440 948 8472
rect 52 8368 84 8400
rect 124 8368 156 8400
rect 196 8368 228 8400
rect 268 8368 300 8400
rect 340 8368 372 8400
rect 412 8368 444 8400
rect 484 8368 516 8400
rect 556 8368 588 8400
rect 628 8368 660 8400
rect 700 8368 732 8400
rect 772 8368 804 8400
rect 844 8368 876 8400
rect 916 8368 948 8400
rect 52 8296 84 8328
rect 124 8296 156 8328
rect 196 8296 228 8328
rect 268 8296 300 8328
rect 340 8296 372 8328
rect 412 8296 444 8328
rect 484 8296 516 8328
rect 556 8296 588 8328
rect 628 8296 660 8328
rect 700 8296 732 8328
rect 772 8296 804 8328
rect 844 8296 876 8328
rect 916 8296 948 8328
rect 52 8224 84 8256
rect 124 8224 156 8256
rect 196 8224 228 8256
rect 268 8224 300 8256
rect 340 8224 372 8256
rect 412 8224 444 8256
rect 484 8224 516 8256
rect 556 8224 588 8256
rect 628 8224 660 8256
rect 700 8224 732 8256
rect 772 8224 804 8256
rect 844 8224 876 8256
rect 916 8224 948 8256
rect 52 8152 84 8184
rect 124 8152 156 8184
rect 196 8152 228 8184
rect 268 8152 300 8184
rect 340 8152 372 8184
rect 412 8152 444 8184
rect 484 8152 516 8184
rect 556 8152 588 8184
rect 628 8152 660 8184
rect 700 8152 732 8184
rect 772 8152 804 8184
rect 844 8152 876 8184
rect 916 8152 948 8184
rect 52 8080 84 8112
rect 124 8080 156 8112
rect 196 8080 228 8112
rect 268 8080 300 8112
rect 340 8080 372 8112
rect 412 8080 444 8112
rect 484 8080 516 8112
rect 556 8080 588 8112
rect 628 8080 660 8112
rect 700 8080 732 8112
rect 772 8080 804 8112
rect 844 8080 876 8112
rect 916 8080 948 8112
rect 52 8008 84 8040
rect 124 8008 156 8040
rect 196 8008 228 8040
rect 268 8008 300 8040
rect 340 8008 372 8040
rect 412 8008 444 8040
rect 484 8008 516 8040
rect 556 8008 588 8040
rect 628 8008 660 8040
rect 700 8008 732 8040
rect 772 8008 804 8040
rect 844 8008 876 8040
rect 916 8008 948 8040
rect 52 7936 84 7968
rect 124 7936 156 7968
rect 196 7936 228 7968
rect 268 7936 300 7968
rect 340 7936 372 7968
rect 412 7936 444 7968
rect 484 7936 516 7968
rect 556 7936 588 7968
rect 628 7936 660 7968
rect 700 7936 732 7968
rect 772 7936 804 7968
rect 844 7936 876 7968
rect 916 7936 948 7968
rect 52 7864 84 7896
rect 124 7864 156 7896
rect 196 7864 228 7896
rect 268 7864 300 7896
rect 340 7864 372 7896
rect 412 7864 444 7896
rect 484 7864 516 7896
rect 556 7864 588 7896
rect 628 7864 660 7896
rect 700 7864 732 7896
rect 772 7864 804 7896
rect 844 7864 876 7896
rect 916 7864 948 7896
rect 52 7792 84 7824
rect 124 7792 156 7824
rect 196 7792 228 7824
rect 268 7792 300 7824
rect 340 7792 372 7824
rect 412 7792 444 7824
rect 484 7792 516 7824
rect 556 7792 588 7824
rect 628 7792 660 7824
rect 700 7792 732 7824
rect 772 7792 804 7824
rect 844 7792 876 7824
rect 916 7792 948 7824
rect 52 7720 84 7752
rect 124 7720 156 7752
rect 196 7720 228 7752
rect 268 7720 300 7752
rect 340 7720 372 7752
rect 412 7720 444 7752
rect 484 7720 516 7752
rect 556 7720 588 7752
rect 628 7720 660 7752
rect 700 7720 732 7752
rect 772 7720 804 7752
rect 844 7720 876 7752
rect 916 7720 948 7752
rect 52 7648 84 7680
rect 124 7648 156 7680
rect 196 7648 228 7680
rect 268 7648 300 7680
rect 340 7648 372 7680
rect 412 7648 444 7680
rect 484 7648 516 7680
rect 556 7648 588 7680
rect 628 7648 660 7680
rect 700 7648 732 7680
rect 772 7648 804 7680
rect 844 7648 876 7680
rect 916 7648 948 7680
rect 52 7576 84 7608
rect 124 7576 156 7608
rect 196 7576 228 7608
rect 268 7576 300 7608
rect 340 7576 372 7608
rect 412 7576 444 7608
rect 484 7576 516 7608
rect 556 7576 588 7608
rect 628 7576 660 7608
rect 700 7576 732 7608
rect 772 7576 804 7608
rect 844 7576 876 7608
rect 916 7576 948 7608
rect 52 7504 84 7536
rect 124 7504 156 7536
rect 196 7504 228 7536
rect 268 7504 300 7536
rect 340 7504 372 7536
rect 412 7504 444 7536
rect 484 7504 516 7536
rect 556 7504 588 7536
rect 628 7504 660 7536
rect 700 7504 732 7536
rect 772 7504 804 7536
rect 844 7504 876 7536
rect 916 7504 948 7536
rect 52 7432 84 7464
rect 124 7432 156 7464
rect 196 7432 228 7464
rect 268 7432 300 7464
rect 340 7432 372 7464
rect 412 7432 444 7464
rect 484 7432 516 7464
rect 556 7432 588 7464
rect 628 7432 660 7464
rect 700 7432 732 7464
rect 772 7432 804 7464
rect 844 7432 876 7464
rect 916 7432 948 7464
rect 52 7360 84 7392
rect 124 7360 156 7392
rect 196 7360 228 7392
rect 268 7360 300 7392
rect 340 7360 372 7392
rect 412 7360 444 7392
rect 484 7360 516 7392
rect 556 7360 588 7392
rect 628 7360 660 7392
rect 700 7360 732 7392
rect 772 7360 804 7392
rect 844 7360 876 7392
rect 916 7360 948 7392
rect 52 7288 84 7320
rect 124 7288 156 7320
rect 196 7288 228 7320
rect 268 7288 300 7320
rect 340 7288 372 7320
rect 412 7288 444 7320
rect 484 7288 516 7320
rect 556 7288 588 7320
rect 628 7288 660 7320
rect 700 7288 732 7320
rect 772 7288 804 7320
rect 844 7288 876 7320
rect 916 7288 948 7320
rect 52 7216 84 7248
rect 124 7216 156 7248
rect 196 7216 228 7248
rect 268 7216 300 7248
rect 340 7216 372 7248
rect 412 7216 444 7248
rect 484 7216 516 7248
rect 556 7216 588 7248
rect 628 7216 660 7248
rect 700 7216 732 7248
rect 772 7216 804 7248
rect 844 7216 876 7248
rect 916 7216 948 7248
rect 52 7144 84 7176
rect 124 7144 156 7176
rect 196 7144 228 7176
rect 268 7144 300 7176
rect 340 7144 372 7176
rect 412 7144 444 7176
rect 484 7144 516 7176
rect 556 7144 588 7176
rect 628 7144 660 7176
rect 700 7144 732 7176
rect 772 7144 804 7176
rect 844 7144 876 7176
rect 916 7144 948 7176
rect 52 7072 84 7104
rect 124 7072 156 7104
rect 196 7072 228 7104
rect 268 7072 300 7104
rect 340 7072 372 7104
rect 412 7072 444 7104
rect 484 7072 516 7104
rect 556 7072 588 7104
rect 628 7072 660 7104
rect 700 7072 732 7104
rect 772 7072 804 7104
rect 844 7072 876 7104
rect 916 7072 948 7104
rect 52 7000 84 7032
rect 124 7000 156 7032
rect 196 7000 228 7032
rect 268 7000 300 7032
rect 340 7000 372 7032
rect 412 7000 444 7032
rect 484 7000 516 7032
rect 556 7000 588 7032
rect 628 7000 660 7032
rect 700 7000 732 7032
rect 772 7000 804 7032
rect 844 7000 876 7032
rect 916 7000 948 7032
rect 52 6928 84 6960
rect 124 6928 156 6960
rect 196 6928 228 6960
rect 268 6928 300 6960
rect 340 6928 372 6960
rect 412 6928 444 6960
rect 484 6928 516 6960
rect 556 6928 588 6960
rect 628 6928 660 6960
rect 700 6928 732 6960
rect 772 6928 804 6960
rect 844 6928 876 6960
rect 916 6928 948 6960
rect 52 6856 84 6888
rect 124 6856 156 6888
rect 196 6856 228 6888
rect 268 6856 300 6888
rect 340 6856 372 6888
rect 412 6856 444 6888
rect 484 6856 516 6888
rect 556 6856 588 6888
rect 628 6856 660 6888
rect 700 6856 732 6888
rect 772 6856 804 6888
rect 844 6856 876 6888
rect 916 6856 948 6888
rect 124 6512 156 6544
rect 196 6512 228 6544
rect 268 6512 300 6544
rect 340 6512 372 6544
rect 412 6512 444 6544
rect 484 6512 516 6544
rect 556 6512 588 6544
rect 628 6512 660 6544
rect 700 6512 732 6544
rect 772 6512 804 6544
rect 844 6512 876 6544
rect 916 6512 948 6544
rect 52 6440 84 6472
rect 124 6440 156 6472
rect 196 6440 228 6472
rect 268 6440 300 6472
rect 340 6440 372 6472
rect 412 6440 444 6472
rect 484 6440 516 6472
rect 556 6440 588 6472
rect 628 6440 660 6472
rect 700 6440 732 6472
rect 772 6440 804 6472
rect 844 6440 876 6472
rect 916 6440 948 6472
rect 52 6368 84 6400
rect 124 6368 156 6400
rect 196 6368 228 6400
rect 268 6368 300 6400
rect 340 6368 372 6400
rect 412 6368 444 6400
rect 484 6368 516 6400
rect 556 6368 588 6400
rect 628 6368 660 6400
rect 700 6368 732 6400
rect 772 6368 804 6400
rect 844 6368 876 6400
rect 916 6368 948 6400
rect 52 6296 84 6328
rect 124 6296 156 6328
rect 196 6296 228 6328
rect 268 6296 300 6328
rect 340 6296 372 6328
rect 412 6296 444 6328
rect 484 6296 516 6328
rect 556 6296 588 6328
rect 628 6296 660 6328
rect 700 6296 732 6328
rect 772 6296 804 6328
rect 844 6296 876 6328
rect 916 6296 948 6328
rect 52 6224 84 6256
rect 124 6224 156 6256
rect 196 6224 228 6256
rect 268 6224 300 6256
rect 340 6224 372 6256
rect 412 6224 444 6256
rect 484 6224 516 6256
rect 556 6224 588 6256
rect 628 6224 660 6256
rect 700 6224 732 6256
rect 772 6224 804 6256
rect 844 6224 876 6256
rect 916 6224 948 6256
rect 52 6152 84 6184
rect 124 6152 156 6184
rect 196 6152 228 6184
rect 268 6152 300 6184
rect 340 6152 372 6184
rect 412 6152 444 6184
rect 484 6152 516 6184
rect 556 6152 588 6184
rect 628 6152 660 6184
rect 700 6152 732 6184
rect 772 6152 804 6184
rect 844 6152 876 6184
rect 916 6152 948 6184
rect 52 6080 84 6112
rect 124 6080 156 6112
rect 196 6080 228 6112
rect 268 6080 300 6112
rect 340 6080 372 6112
rect 412 6080 444 6112
rect 484 6080 516 6112
rect 556 6080 588 6112
rect 628 6080 660 6112
rect 700 6080 732 6112
rect 772 6080 804 6112
rect 844 6080 876 6112
rect 916 6080 948 6112
rect 52 6008 84 6040
rect 124 6008 156 6040
rect 196 6008 228 6040
rect 268 6008 300 6040
rect 340 6008 372 6040
rect 412 6008 444 6040
rect 484 6008 516 6040
rect 556 6008 588 6040
rect 628 6008 660 6040
rect 700 6008 732 6040
rect 772 6008 804 6040
rect 844 6008 876 6040
rect 916 6008 948 6040
rect 52 5936 84 5968
rect 124 5936 156 5968
rect 196 5936 228 5968
rect 268 5936 300 5968
rect 340 5936 372 5968
rect 412 5936 444 5968
rect 484 5936 516 5968
rect 556 5936 588 5968
rect 628 5936 660 5968
rect 700 5936 732 5968
rect 772 5936 804 5968
rect 844 5936 876 5968
rect 916 5936 948 5968
rect 52 5864 84 5896
rect 124 5864 156 5896
rect 196 5864 228 5896
rect 268 5864 300 5896
rect 340 5864 372 5896
rect 412 5864 444 5896
rect 484 5864 516 5896
rect 556 5864 588 5896
rect 628 5864 660 5896
rect 700 5864 732 5896
rect 772 5864 804 5896
rect 844 5864 876 5896
rect 916 5864 948 5896
rect 52 5792 84 5824
rect 124 5792 156 5824
rect 196 5792 228 5824
rect 268 5792 300 5824
rect 340 5792 372 5824
rect 412 5792 444 5824
rect 484 5792 516 5824
rect 556 5792 588 5824
rect 628 5792 660 5824
rect 700 5792 732 5824
rect 772 5792 804 5824
rect 844 5792 876 5824
rect 916 5792 948 5824
rect 52 5720 84 5752
rect 124 5720 156 5752
rect 196 5720 228 5752
rect 268 5720 300 5752
rect 340 5720 372 5752
rect 412 5720 444 5752
rect 484 5720 516 5752
rect 556 5720 588 5752
rect 628 5720 660 5752
rect 700 5720 732 5752
rect 772 5720 804 5752
rect 844 5720 876 5752
rect 916 5720 948 5752
rect 52 5648 84 5680
rect 124 5648 156 5680
rect 196 5648 228 5680
rect 268 5648 300 5680
rect 340 5648 372 5680
rect 412 5648 444 5680
rect 484 5648 516 5680
rect 556 5648 588 5680
rect 628 5648 660 5680
rect 700 5648 732 5680
rect 772 5648 804 5680
rect 844 5648 876 5680
rect 916 5648 948 5680
rect 52 5576 84 5608
rect 124 5576 156 5608
rect 196 5576 228 5608
rect 268 5576 300 5608
rect 340 5576 372 5608
rect 412 5576 444 5608
rect 484 5576 516 5608
rect 556 5576 588 5608
rect 628 5576 660 5608
rect 700 5576 732 5608
rect 772 5576 804 5608
rect 844 5576 876 5608
rect 916 5576 948 5608
rect 52 5504 84 5536
rect 124 5504 156 5536
rect 196 5504 228 5536
rect 268 5504 300 5536
rect 340 5504 372 5536
rect 412 5504 444 5536
rect 484 5504 516 5536
rect 556 5504 588 5536
rect 628 5504 660 5536
rect 700 5504 732 5536
rect 772 5504 804 5536
rect 844 5504 876 5536
rect 916 5504 948 5536
rect 52 5432 84 5464
rect 124 5432 156 5464
rect 196 5432 228 5464
rect 268 5432 300 5464
rect 340 5432 372 5464
rect 412 5432 444 5464
rect 484 5432 516 5464
rect 556 5432 588 5464
rect 628 5432 660 5464
rect 700 5432 732 5464
rect 772 5432 804 5464
rect 844 5432 876 5464
rect 916 5432 948 5464
rect 52 5360 84 5392
rect 124 5360 156 5392
rect 196 5360 228 5392
rect 268 5360 300 5392
rect 340 5360 372 5392
rect 412 5360 444 5392
rect 484 5360 516 5392
rect 556 5360 588 5392
rect 628 5360 660 5392
rect 700 5360 732 5392
rect 772 5360 804 5392
rect 844 5360 876 5392
rect 916 5360 948 5392
rect 52 5288 84 5320
rect 124 5288 156 5320
rect 196 5288 228 5320
rect 268 5288 300 5320
rect 340 5288 372 5320
rect 412 5288 444 5320
rect 484 5288 516 5320
rect 556 5288 588 5320
rect 628 5288 660 5320
rect 700 5288 732 5320
rect 772 5288 804 5320
rect 844 5288 876 5320
rect 916 5288 948 5320
rect 52 5216 84 5248
rect 124 5216 156 5248
rect 196 5216 228 5248
rect 268 5216 300 5248
rect 340 5216 372 5248
rect 412 5216 444 5248
rect 484 5216 516 5248
rect 556 5216 588 5248
rect 628 5216 660 5248
rect 700 5216 732 5248
rect 772 5216 804 5248
rect 844 5216 876 5248
rect 916 5216 948 5248
rect 52 5144 84 5176
rect 124 5144 156 5176
rect 196 5144 228 5176
rect 268 5144 300 5176
rect 340 5144 372 5176
rect 412 5144 444 5176
rect 484 5144 516 5176
rect 556 5144 588 5176
rect 628 5144 660 5176
rect 700 5144 732 5176
rect 772 5144 804 5176
rect 844 5144 876 5176
rect 916 5144 948 5176
rect 52 5072 84 5104
rect 124 5072 156 5104
rect 196 5072 228 5104
rect 268 5072 300 5104
rect 340 5072 372 5104
rect 412 5072 444 5104
rect 484 5072 516 5104
rect 556 5072 588 5104
rect 628 5072 660 5104
rect 700 5072 732 5104
rect 772 5072 804 5104
rect 844 5072 876 5104
rect 916 5072 948 5104
rect 52 5000 84 5032
rect 124 5000 156 5032
rect 196 5000 228 5032
rect 268 5000 300 5032
rect 340 5000 372 5032
rect 412 5000 444 5032
rect 484 5000 516 5032
rect 556 5000 588 5032
rect 628 5000 660 5032
rect 700 5000 732 5032
rect 772 5000 804 5032
rect 844 5000 876 5032
rect 916 5000 948 5032
rect 52 4928 84 4960
rect 124 4928 156 4960
rect 196 4928 228 4960
rect 268 4928 300 4960
rect 340 4928 372 4960
rect 412 4928 444 4960
rect 484 4928 516 4960
rect 556 4928 588 4960
rect 628 4928 660 4960
rect 700 4928 732 4960
rect 772 4928 804 4960
rect 844 4928 876 4960
rect 916 4928 948 4960
rect 52 4856 84 4888
rect 124 4856 156 4888
rect 196 4856 228 4888
rect 268 4856 300 4888
rect 340 4856 372 4888
rect 412 4856 444 4888
rect 484 4856 516 4888
rect 556 4856 588 4888
rect 628 4856 660 4888
rect 700 4856 732 4888
rect 772 4856 804 4888
rect 844 4856 876 4888
rect 916 4856 948 4888
rect 52 4784 84 4816
rect 124 4784 156 4816
rect 196 4784 228 4816
rect 268 4784 300 4816
rect 340 4784 372 4816
rect 412 4784 444 4816
rect 484 4784 516 4816
rect 556 4784 588 4816
rect 628 4784 660 4816
rect 700 4784 732 4816
rect 772 4784 804 4816
rect 844 4784 876 4816
rect 916 4784 948 4816
rect 52 4712 84 4744
rect 124 4712 156 4744
rect 196 4712 228 4744
rect 268 4712 300 4744
rect 340 4712 372 4744
rect 412 4712 444 4744
rect 484 4712 516 4744
rect 556 4712 588 4744
rect 628 4712 660 4744
rect 700 4712 732 4744
rect 772 4712 804 4744
rect 844 4712 876 4744
rect 916 4712 948 4744
rect 52 4640 84 4672
rect 124 4640 156 4672
rect 196 4640 228 4672
rect 268 4640 300 4672
rect 340 4640 372 4672
rect 412 4640 444 4672
rect 484 4640 516 4672
rect 556 4640 588 4672
rect 628 4640 660 4672
rect 700 4640 732 4672
rect 772 4640 804 4672
rect 844 4640 876 4672
rect 916 4640 948 4672
rect 52 4568 84 4600
rect 124 4568 156 4600
rect 196 4568 228 4600
rect 268 4568 300 4600
rect 340 4568 372 4600
rect 412 4568 444 4600
rect 484 4568 516 4600
rect 556 4568 588 4600
rect 628 4568 660 4600
rect 700 4568 732 4600
rect 772 4568 804 4600
rect 844 4568 876 4600
rect 916 4568 948 4600
rect 52 4496 84 4528
rect 124 4496 156 4528
rect 196 4496 228 4528
rect 268 4496 300 4528
rect 340 4496 372 4528
rect 412 4496 444 4528
rect 484 4496 516 4528
rect 556 4496 588 4528
rect 628 4496 660 4528
rect 700 4496 732 4528
rect 772 4496 804 4528
rect 844 4496 876 4528
rect 916 4496 948 4528
rect 52 4424 84 4456
rect 124 4424 156 4456
rect 196 4424 228 4456
rect 268 4424 300 4456
rect 340 4424 372 4456
rect 412 4424 444 4456
rect 484 4424 516 4456
rect 556 4424 588 4456
rect 628 4424 660 4456
rect 700 4424 732 4456
rect 772 4424 804 4456
rect 844 4424 876 4456
rect 916 4424 948 4456
rect 52 4352 84 4384
rect 124 4352 156 4384
rect 196 4352 228 4384
rect 268 4352 300 4384
rect 340 4352 372 4384
rect 412 4352 444 4384
rect 484 4352 516 4384
rect 556 4352 588 4384
rect 628 4352 660 4384
rect 700 4352 732 4384
rect 772 4352 804 4384
rect 844 4352 876 4384
rect 916 4352 948 4384
rect 52 4280 84 4312
rect 124 4280 156 4312
rect 196 4280 228 4312
rect 268 4280 300 4312
rect 340 4280 372 4312
rect 412 4280 444 4312
rect 484 4280 516 4312
rect 556 4280 588 4312
rect 628 4280 660 4312
rect 700 4280 732 4312
rect 772 4280 804 4312
rect 844 4280 876 4312
rect 916 4280 948 4312
rect 52 4208 84 4240
rect 124 4208 156 4240
rect 196 4208 228 4240
rect 268 4208 300 4240
rect 340 4208 372 4240
rect 412 4208 444 4240
rect 484 4208 516 4240
rect 556 4208 588 4240
rect 628 4208 660 4240
rect 700 4208 732 4240
rect 772 4208 804 4240
rect 844 4208 876 4240
rect 916 4208 948 4240
rect 52 4136 84 4168
rect 124 4136 156 4168
rect 196 4136 228 4168
rect 268 4136 300 4168
rect 340 4136 372 4168
rect 412 4136 444 4168
rect 484 4136 516 4168
rect 556 4136 588 4168
rect 628 4136 660 4168
rect 700 4136 732 4168
rect 772 4136 804 4168
rect 844 4136 876 4168
rect 916 4136 948 4168
rect 52 4064 84 4096
rect 124 4064 156 4096
rect 196 4064 228 4096
rect 268 4064 300 4096
rect 340 4064 372 4096
rect 412 4064 444 4096
rect 484 4064 516 4096
rect 556 4064 588 4096
rect 628 4064 660 4096
rect 700 4064 732 4096
rect 772 4064 804 4096
rect 844 4064 876 4096
rect 916 4064 948 4096
rect 52 3992 84 4024
rect 124 3992 156 4024
rect 196 3992 228 4024
rect 268 3992 300 4024
rect 340 3992 372 4024
rect 412 3992 444 4024
rect 484 3992 516 4024
rect 556 3992 588 4024
rect 628 3992 660 4024
rect 700 3992 732 4024
rect 772 3992 804 4024
rect 844 3992 876 4024
rect 916 3992 948 4024
rect 52 3920 84 3952
rect 124 3920 156 3952
rect 196 3920 228 3952
rect 268 3920 300 3952
rect 340 3920 372 3952
rect 412 3920 444 3952
rect 484 3920 516 3952
rect 556 3920 588 3952
rect 628 3920 660 3952
rect 700 3920 732 3952
rect 772 3920 804 3952
rect 844 3920 876 3952
rect 916 3920 948 3952
rect 52 3848 84 3880
rect 124 3848 156 3880
rect 196 3848 228 3880
rect 268 3848 300 3880
rect 340 3848 372 3880
rect 412 3848 444 3880
rect 484 3848 516 3880
rect 556 3848 588 3880
rect 628 3848 660 3880
rect 700 3848 732 3880
rect 772 3848 804 3880
rect 844 3848 876 3880
rect 916 3848 948 3880
rect 52 3776 84 3808
rect 124 3776 156 3808
rect 196 3776 228 3808
rect 268 3776 300 3808
rect 340 3776 372 3808
rect 412 3776 444 3808
rect 484 3776 516 3808
rect 556 3776 588 3808
rect 628 3776 660 3808
rect 700 3776 732 3808
rect 772 3776 804 3808
rect 844 3776 876 3808
rect 916 3776 948 3808
rect 52 3704 84 3736
rect 124 3704 156 3736
rect 196 3704 228 3736
rect 268 3704 300 3736
rect 340 3704 372 3736
rect 412 3704 444 3736
rect 484 3704 516 3736
rect 556 3704 588 3736
rect 628 3704 660 3736
rect 700 3704 732 3736
rect 772 3704 804 3736
rect 844 3704 876 3736
rect 916 3704 948 3736
rect 52 3632 84 3664
rect 124 3632 156 3664
rect 196 3632 228 3664
rect 268 3632 300 3664
rect 340 3632 372 3664
rect 412 3632 444 3664
rect 484 3632 516 3664
rect 556 3632 588 3664
rect 628 3632 660 3664
rect 700 3632 732 3664
rect 772 3632 804 3664
rect 844 3632 876 3664
rect 916 3632 948 3664
rect 52 3560 84 3592
rect 124 3560 156 3592
rect 196 3560 228 3592
rect 268 3560 300 3592
rect 340 3560 372 3592
rect 412 3560 444 3592
rect 484 3560 516 3592
rect 556 3560 588 3592
rect 628 3560 660 3592
rect 700 3560 732 3592
rect 772 3560 804 3592
rect 844 3560 876 3592
rect 916 3560 948 3592
rect 52 3488 84 3520
rect 124 3488 156 3520
rect 196 3488 228 3520
rect 268 3488 300 3520
rect 340 3488 372 3520
rect 412 3488 444 3520
rect 484 3488 516 3520
rect 556 3488 588 3520
rect 628 3488 660 3520
rect 700 3488 732 3520
rect 772 3488 804 3520
rect 844 3488 876 3520
rect 916 3488 948 3520
rect 52 3416 84 3448
rect 124 3416 156 3448
rect 196 3416 228 3448
rect 268 3416 300 3448
rect 340 3416 372 3448
rect 412 3416 444 3448
rect 484 3416 516 3448
rect 556 3416 588 3448
rect 628 3416 660 3448
rect 700 3416 732 3448
rect 772 3416 804 3448
rect 844 3416 876 3448
rect 916 3416 948 3448
rect 52 3344 84 3376
rect 124 3344 156 3376
rect 196 3344 228 3376
rect 268 3344 300 3376
rect 340 3344 372 3376
rect 412 3344 444 3376
rect 484 3344 516 3376
rect 556 3344 588 3376
rect 628 3344 660 3376
rect 700 3344 732 3376
rect 772 3344 804 3376
rect 844 3344 876 3376
rect 916 3344 948 3376
rect 52 3272 84 3304
rect 124 3272 156 3304
rect 196 3272 228 3304
rect 268 3272 300 3304
rect 340 3272 372 3304
rect 412 3272 444 3304
rect 484 3272 516 3304
rect 556 3272 588 3304
rect 628 3272 660 3304
rect 700 3272 732 3304
rect 772 3272 804 3304
rect 844 3272 876 3304
rect 916 3272 948 3304
rect 52 3200 84 3232
rect 124 3200 156 3232
rect 196 3200 228 3232
rect 268 3200 300 3232
rect 340 3200 372 3232
rect 412 3200 444 3232
rect 484 3200 516 3232
rect 556 3200 588 3232
rect 628 3200 660 3232
rect 700 3200 732 3232
rect 772 3200 804 3232
rect 844 3200 876 3232
rect 916 3200 948 3232
rect 52 3128 84 3160
rect 124 3128 156 3160
rect 196 3128 228 3160
rect 268 3128 300 3160
rect 340 3128 372 3160
rect 412 3128 444 3160
rect 484 3128 516 3160
rect 556 3128 588 3160
rect 628 3128 660 3160
rect 700 3128 732 3160
rect 772 3128 804 3160
rect 844 3128 876 3160
rect 916 3128 948 3160
rect 52 3056 84 3088
rect 124 3056 156 3088
rect 196 3056 228 3088
rect 268 3056 300 3088
rect 340 3056 372 3088
rect 412 3056 444 3088
rect 484 3056 516 3088
rect 556 3056 588 3088
rect 628 3056 660 3088
rect 700 3056 732 3088
rect 772 3056 804 3088
rect 844 3056 876 3088
rect 916 3056 948 3088
rect 52 2984 84 3016
rect 124 2984 156 3016
rect 196 2984 228 3016
rect 268 2984 300 3016
rect 340 2984 372 3016
rect 412 2984 444 3016
rect 484 2984 516 3016
rect 556 2984 588 3016
rect 628 2984 660 3016
rect 700 2984 732 3016
rect 772 2984 804 3016
rect 844 2984 876 3016
rect 916 2984 948 3016
rect 52 2912 84 2944
rect 124 2912 156 2944
rect 196 2912 228 2944
rect 268 2912 300 2944
rect 340 2912 372 2944
rect 412 2912 444 2944
rect 484 2912 516 2944
rect 556 2912 588 2944
rect 628 2912 660 2944
rect 700 2912 732 2944
rect 772 2912 804 2944
rect 844 2912 876 2944
rect 916 2912 948 2944
rect 52 2840 84 2872
rect 124 2840 156 2872
rect 196 2840 228 2872
rect 268 2840 300 2872
rect 340 2840 372 2872
rect 412 2840 444 2872
rect 484 2840 516 2872
rect 556 2840 588 2872
rect 628 2840 660 2872
rect 700 2840 732 2872
rect 772 2840 804 2872
rect 844 2840 876 2872
rect 916 2840 948 2872
rect 52 2768 84 2800
rect 124 2768 156 2800
rect 196 2768 228 2800
rect 268 2768 300 2800
rect 340 2768 372 2800
rect 412 2768 444 2800
rect 484 2768 516 2800
rect 556 2768 588 2800
rect 628 2768 660 2800
rect 700 2768 732 2800
rect 772 2768 804 2800
rect 844 2768 876 2800
rect 916 2768 948 2800
rect 52 2696 84 2728
rect 124 2696 156 2728
rect 196 2696 228 2728
rect 268 2696 300 2728
rect 340 2696 372 2728
rect 412 2696 444 2728
rect 484 2696 516 2728
rect 556 2696 588 2728
rect 628 2696 660 2728
rect 700 2696 732 2728
rect 772 2696 804 2728
rect 844 2696 876 2728
rect 916 2696 948 2728
rect 52 2624 84 2656
rect 124 2624 156 2656
rect 196 2624 228 2656
rect 268 2624 300 2656
rect 340 2624 372 2656
rect 412 2624 444 2656
rect 484 2624 516 2656
rect 556 2624 588 2656
rect 628 2624 660 2656
rect 700 2624 732 2656
rect 772 2624 804 2656
rect 844 2624 876 2656
rect 916 2624 948 2656
rect 52 2552 84 2584
rect 124 2552 156 2584
rect 196 2552 228 2584
rect 268 2552 300 2584
rect 340 2552 372 2584
rect 412 2552 444 2584
rect 484 2552 516 2584
rect 556 2552 588 2584
rect 628 2552 660 2584
rect 700 2552 732 2584
rect 772 2552 804 2584
rect 844 2552 876 2584
rect 916 2552 948 2584
rect 52 2480 84 2512
rect 124 2480 156 2512
rect 196 2480 228 2512
rect 268 2480 300 2512
rect 340 2480 372 2512
rect 412 2480 444 2512
rect 484 2480 516 2512
rect 556 2480 588 2512
rect 628 2480 660 2512
rect 700 2480 732 2512
rect 772 2480 804 2512
rect 844 2480 876 2512
rect 916 2480 948 2512
rect 52 2408 84 2440
rect 124 2408 156 2440
rect 196 2408 228 2440
rect 268 2408 300 2440
rect 340 2408 372 2440
rect 412 2408 444 2440
rect 484 2408 516 2440
rect 556 2408 588 2440
rect 628 2408 660 2440
rect 700 2408 732 2440
rect 772 2408 804 2440
rect 844 2408 876 2440
rect 916 2408 948 2440
rect 52 2336 84 2368
rect 124 2336 156 2368
rect 196 2336 228 2368
rect 268 2336 300 2368
rect 340 2336 372 2368
rect 412 2336 444 2368
rect 484 2336 516 2368
rect 556 2336 588 2368
rect 628 2336 660 2368
rect 700 2336 732 2368
rect 772 2336 804 2368
rect 844 2336 876 2368
rect 916 2336 948 2368
rect 52 2264 84 2296
rect 124 2264 156 2296
rect 196 2264 228 2296
rect 268 2264 300 2296
rect 340 2264 372 2296
rect 412 2264 444 2296
rect 484 2264 516 2296
rect 556 2264 588 2296
rect 628 2264 660 2296
rect 700 2264 732 2296
rect 772 2264 804 2296
rect 844 2264 876 2296
rect 916 2264 948 2296
rect 52 2192 84 2224
rect 124 2192 156 2224
rect 196 2192 228 2224
rect 268 2192 300 2224
rect 340 2192 372 2224
rect 412 2192 444 2224
rect 484 2192 516 2224
rect 556 2192 588 2224
rect 628 2192 660 2224
rect 700 2192 732 2224
rect 772 2192 804 2224
rect 844 2192 876 2224
rect 916 2192 948 2224
rect 52 2120 84 2152
rect 124 2120 156 2152
rect 196 2120 228 2152
rect 268 2120 300 2152
rect 340 2120 372 2152
rect 412 2120 444 2152
rect 484 2120 516 2152
rect 556 2120 588 2152
rect 628 2120 660 2152
rect 700 2120 732 2152
rect 772 2120 804 2152
rect 844 2120 876 2152
rect 916 2120 948 2152
rect 52 2048 84 2080
rect 124 2048 156 2080
rect 196 2048 228 2080
rect 268 2048 300 2080
rect 340 2048 372 2080
rect 412 2048 444 2080
rect 484 2048 516 2080
rect 556 2048 588 2080
rect 628 2048 660 2080
rect 700 2048 732 2080
rect 772 2048 804 2080
rect 844 2048 876 2080
rect 916 2048 948 2080
rect 52 1976 84 2008
rect 124 1976 156 2008
rect 196 1976 228 2008
rect 268 1976 300 2008
rect 340 1976 372 2008
rect 412 1976 444 2008
rect 484 1976 516 2008
rect 556 1976 588 2008
rect 628 1976 660 2008
rect 700 1976 732 2008
rect 772 1976 804 2008
rect 844 1976 876 2008
rect 916 1976 948 2008
rect 52 1904 84 1936
rect 124 1904 156 1936
rect 196 1904 228 1936
rect 268 1904 300 1936
rect 340 1904 372 1936
rect 412 1904 444 1936
rect 484 1904 516 1936
rect 556 1904 588 1936
rect 628 1904 660 1936
rect 700 1904 732 1936
rect 772 1904 804 1936
rect 844 1904 876 1936
rect 916 1904 948 1936
rect 52 1832 84 1864
rect 124 1832 156 1864
rect 196 1832 228 1864
rect 268 1832 300 1864
rect 340 1832 372 1864
rect 412 1832 444 1864
rect 484 1832 516 1864
rect 556 1832 588 1864
rect 628 1832 660 1864
rect 700 1832 732 1864
rect 772 1832 804 1864
rect 844 1832 876 1864
rect 916 1832 948 1864
rect 52 1760 84 1792
rect 124 1760 156 1792
rect 196 1760 228 1792
rect 268 1760 300 1792
rect 340 1760 372 1792
rect 412 1760 444 1792
rect 484 1760 516 1792
rect 556 1760 588 1792
rect 628 1760 660 1792
rect 700 1760 732 1792
rect 772 1760 804 1792
rect 844 1760 876 1792
rect 916 1760 948 1792
rect 52 1688 84 1720
rect 124 1688 156 1720
rect 196 1688 228 1720
rect 268 1688 300 1720
rect 340 1688 372 1720
rect 412 1688 444 1720
rect 484 1688 516 1720
rect 556 1688 588 1720
rect 628 1688 660 1720
rect 700 1688 732 1720
rect 772 1688 804 1720
rect 844 1688 876 1720
rect 916 1688 948 1720
rect 52 1616 84 1648
rect 124 1616 156 1648
rect 196 1616 228 1648
rect 268 1616 300 1648
rect 340 1616 372 1648
rect 412 1616 444 1648
rect 484 1616 516 1648
rect 556 1616 588 1648
rect 628 1616 660 1648
rect 700 1616 732 1648
rect 772 1616 804 1648
rect 844 1616 876 1648
rect 916 1616 948 1648
rect 52 1544 84 1576
rect 124 1544 156 1576
rect 196 1544 228 1576
rect 268 1544 300 1576
rect 340 1544 372 1576
rect 412 1544 444 1576
rect 484 1544 516 1576
rect 556 1544 588 1576
rect 628 1544 660 1576
rect 700 1544 732 1576
rect 772 1544 804 1576
rect 844 1544 876 1576
rect 916 1544 948 1576
rect 52 1472 84 1504
rect 124 1472 156 1504
rect 196 1472 228 1504
rect 268 1472 300 1504
rect 340 1472 372 1504
rect 412 1472 444 1504
rect 484 1472 516 1504
rect 556 1472 588 1504
rect 628 1472 660 1504
rect 700 1472 732 1504
rect 772 1472 804 1504
rect 844 1472 876 1504
rect 916 1472 948 1504
rect 52 1400 84 1432
rect 124 1400 156 1432
rect 196 1400 228 1432
rect 268 1400 300 1432
rect 340 1400 372 1432
rect 412 1400 444 1432
rect 484 1400 516 1432
rect 556 1400 588 1432
rect 628 1400 660 1432
rect 700 1400 732 1432
rect 772 1400 804 1432
rect 844 1400 876 1432
rect 916 1400 948 1432
rect 52 1328 84 1360
rect 124 1328 156 1360
rect 196 1328 228 1360
rect 268 1328 300 1360
rect 340 1328 372 1360
rect 412 1328 444 1360
rect 484 1328 516 1360
rect 556 1328 588 1360
rect 628 1328 660 1360
rect 700 1328 732 1360
rect 772 1328 804 1360
rect 844 1328 876 1360
rect 916 1328 948 1360
rect 52 1256 84 1288
rect 124 1256 156 1288
rect 196 1256 228 1288
rect 268 1256 300 1288
rect 340 1256 372 1288
rect 412 1256 444 1288
rect 484 1256 516 1288
rect 556 1256 588 1288
rect 628 1256 660 1288
rect 700 1256 732 1288
rect 772 1256 804 1288
rect 844 1256 876 1288
rect 916 1256 948 1288
rect 292 31384 324 31416
rect 362 31384 394 31416
rect 431 31384 463 31416
rect 502 31384 534 31416
rect 572 31384 604 31416
rect 640 31384 672 31416
rect 710 31384 742 31416
rect 196 27939 228 27971
rect 268 27939 300 27971
rect 340 27939 372 27971
rect 412 27939 444 27971
rect 484 27939 516 27971
rect 556 27939 588 27971
rect 628 27939 660 27971
rect 700 27939 732 27971
rect 772 27939 804 27971
rect 844 27939 876 27971
rect 124 27867 156 27899
rect 196 27867 228 27899
rect 268 27867 300 27899
rect 340 27867 372 27899
rect 412 27867 444 27899
rect 484 27867 516 27899
rect 556 27867 588 27899
rect 628 27867 660 27899
rect 700 27867 732 27899
rect 772 27867 804 27899
rect 844 27867 876 27899
rect 124 27795 156 27827
rect 196 27795 228 27827
rect 268 27795 300 27827
rect 340 27795 372 27827
rect 412 27795 444 27827
rect 484 27795 516 27827
rect 556 27795 588 27827
rect 628 27795 660 27827
rect 700 27795 732 27827
rect 772 27795 804 27827
rect 844 27795 876 27827
rect 124 27723 156 27755
rect 196 27723 228 27755
rect 268 27723 300 27755
rect 340 27723 372 27755
rect 412 27723 444 27755
rect 484 27723 516 27755
rect 556 27723 588 27755
rect 628 27723 660 27755
rect 700 27723 732 27755
rect 772 27723 804 27755
rect 844 27723 876 27755
rect 124 27651 156 27683
rect 196 27651 228 27683
rect 268 27651 300 27683
rect 340 27651 372 27683
rect 412 27651 444 27683
rect 484 27651 516 27683
rect 556 27651 588 27683
rect 628 27651 660 27683
rect 700 27651 732 27683
rect 772 27651 804 27683
rect 844 27651 876 27683
rect 124 27579 156 27611
rect 196 27579 228 27611
rect 268 27579 300 27611
rect 340 27579 372 27611
rect 412 27579 444 27611
rect 484 27579 516 27611
rect 556 27579 588 27611
rect 628 27579 660 27611
rect 700 27579 732 27611
rect 772 27579 804 27611
rect 844 27579 876 27611
rect 124 27507 156 27539
rect 196 27507 228 27539
rect 268 27507 300 27539
rect 340 27507 372 27539
rect 412 27507 444 27539
rect 484 27507 516 27539
rect 556 27507 588 27539
rect 628 27507 660 27539
rect 700 27507 732 27539
rect 772 27507 804 27539
rect 844 27507 876 27539
rect 124 27435 156 27467
rect 196 27435 228 27467
rect 268 27435 300 27467
rect 340 27435 372 27467
rect 412 27435 444 27467
rect 484 27435 516 27467
rect 556 27435 588 27467
rect 628 27435 660 27467
rect 700 27435 732 27467
rect 772 27435 804 27467
rect 844 27435 876 27467
rect 124 27363 156 27395
rect 196 27363 228 27395
rect 268 27363 300 27395
rect 340 27363 372 27395
rect 412 27363 444 27395
rect 484 27363 516 27395
rect 556 27363 588 27395
rect 628 27363 660 27395
rect 700 27363 732 27395
rect 772 27363 804 27395
rect 844 27363 876 27395
rect 124 27291 156 27323
rect 196 27291 228 27323
rect 268 27291 300 27323
rect 340 27291 372 27323
rect 412 27291 444 27323
rect 484 27291 516 27323
rect 556 27291 588 27323
rect 628 27291 660 27323
rect 700 27291 732 27323
rect 772 27291 804 27323
rect 844 27291 876 27323
rect 124 27219 156 27251
rect 196 27219 228 27251
rect 268 27219 300 27251
rect 340 27219 372 27251
rect 412 27219 444 27251
rect 484 27219 516 27251
rect 556 27219 588 27251
rect 628 27219 660 27251
rect 700 27219 732 27251
rect 772 27219 804 27251
rect 844 27219 876 27251
rect 124 27147 156 27179
rect 196 27147 228 27179
rect 268 27147 300 27179
rect 340 27147 372 27179
rect 412 27147 444 27179
rect 484 27147 516 27179
rect 556 27147 588 27179
rect 628 27147 660 27179
rect 700 27147 732 27179
rect 772 27147 804 27179
rect 844 27147 876 27179
rect 124 27075 156 27107
rect 196 27075 228 27107
rect 268 27075 300 27107
rect 340 27075 372 27107
rect 412 27075 444 27107
rect 484 27075 516 27107
rect 556 27075 588 27107
rect 628 27075 660 27107
rect 700 27075 732 27107
rect 772 27075 804 27107
rect 844 27075 876 27107
rect 124 27003 156 27035
rect 196 27003 228 27035
rect 268 27003 300 27035
rect 340 27003 372 27035
rect 412 27003 444 27035
rect 484 27003 516 27035
rect 556 27003 588 27035
rect 628 27003 660 27035
rect 700 27003 732 27035
rect 772 27003 804 27035
rect 844 27003 876 27035
rect 124 26931 156 26963
rect 196 26931 228 26963
rect 268 26931 300 26963
rect 340 26931 372 26963
rect 412 26931 444 26963
rect 484 26931 516 26963
rect 556 26931 588 26963
rect 628 26931 660 26963
rect 700 26931 732 26963
rect 772 26931 804 26963
rect 844 26931 876 26963
rect 124 26859 156 26891
rect 196 26859 228 26891
rect 268 26859 300 26891
rect 340 26859 372 26891
rect 412 26859 444 26891
rect 484 26859 516 26891
rect 556 26859 588 26891
rect 628 26859 660 26891
rect 700 26859 732 26891
rect 772 26859 804 26891
rect 844 26859 876 26891
rect 124 26787 156 26819
rect 196 26787 228 26819
rect 268 26787 300 26819
rect 340 26787 372 26819
rect 412 26787 444 26819
rect 484 26787 516 26819
rect 556 26787 588 26819
rect 628 26787 660 26819
rect 700 26787 732 26819
rect 772 26787 804 26819
rect 844 26787 876 26819
rect 124 26715 156 26747
rect 196 26715 228 26747
rect 268 26715 300 26747
rect 340 26715 372 26747
rect 412 26715 444 26747
rect 484 26715 516 26747
rect 556 26715 588 26747
rect 628 26715 660 26747
rect 700 26715 732 26747
rect 772 26715 804 26747
rect 844 26715 876 26747
rect 124 26643 156 26675
rect 196 26643 228 26675
rect 268 26643 300 26675
rect 340 26643 372 26675
rect 412 26643 444 26675
rect 484 26643 516 26675
rect 556 26643 588 26675
rect 628 26643 660 26675
rect 700 26643 732 26675
rect 772 26643 804 26675
rect 844 26643 876 26675
rect 124 26571 156 26603
rect 196 26571 228 26603
rect 268 26571 300 26603
rect 340 26571 372 26603
rect 412 26571 444 26603
rect 484 26571 516 26603
rect 556 26571 588 26603
rect 628 26571 660 26603
rect 700 26571 732 26603
rect 772 26571 804 26603
rect 844 26571 876 26603
rect 124 26499 156 26531
rect 196 26499 228 26531
rect 268 26499 300 26531
rect 340 26499 372 26531
rect 412 26499 444 26531
rect 484 26499 516 26531
rect 556 26499 588 26531
rect 628 26499 660 26531
rect 700 26499 732 26531
rect 772 26499 804 26531
rect 844 26499 876 26531
rect 124 26427 156 26459
rect 196 26427 228 26459
rect 268 26427 300 26459
rect 340 26427 372 26459
rect 412 26427 444 26459
rect 484 26427 516 26459
rect 556 26427 588 26459
rect 628 26427 660 26459
rect 700 26427 732 26459
rect 772 26427 804 26459
rect 844 26427 876 26459
rect 124 26355 156 26387
rect 196 26355 228 26387
rect 268 26355 300 26387
rect 340 26355 372 26387
rect 412 26355 444 26387
rect 484 26355 516 26387
rect 556 26355 588 26387
rect 628 26355 660 26387
rect 700 26355 732 26387
rect 772 26355 804 26387
rect 844 26355 876 26387
rect 124 26283 156 26315
rect 196 26283 228 26315
rect 268 26283 300 26315
rect 340 26283 372 26315
rect 412 26283 444 26315
rect 484 26283 516 26315
rect 556 26283 588 26315
rect 628 26283 660 26315
rect 700 26283 732 26315
rect 772 26283 804 26315
rect 844 26283 876 26315
rect 124 26211 156 26243
rect 196 26211 228 26243
rect 268 26211 300 26243
rect 340 26211 372 26243
rect 412 26211 444 26243
rect 484 26211 516 26243
rect 556 26211 588 26243
rect 628 26211 660 26243
rect 700 26211 732 26243
rect 772 26211 804 26243
rect 844 26211 876 26243
rect 124 26139 156 26171
rect 196 26139 228 26171
rect 268 26139 300 26171
rect 340 26139 372 26171
rect 412 26139 444 26171
rect 484 26139 516 26171
rect 556 26139 588 26171
rect 628 26139 660 26171
rect 700 26139 732 26171
rect 772 26139 804 26171
rect 844 26139 876 26171
rect 124 26067 156 26099
rect 196 26067 228 26099
rect 268 26067 300 26099
rect 340 26067 372 26099
rect 412 26067 444 26099
rect 484 26067 516 26099
rect 556 26067 588 26099
rect 628 26067 660 26099
rect 700 26067 732 26099
rect 772 26067 804 26099
rect 844 26067 876 26099
rect 124 25995 156 26027
rect 196 25995 228 26027
rect 268 25995 300 26027
rect 340 25995 372 26027
rect 412 25995 444 26027
rect 484 25995 516 26027
rect 556 25995 588 26027
rect 628 25995 660 26027
rect 700 25995 732 26027
rect 772 25995 804 26027
rect 844 25995 876 26027
rect 124 25923 156 25955
rect 196 25923 228 25955
rect 268 25923 300 25955
rect 340 25923 372 25955
rect 412 25923 444 25955
rect 484 25923 516 25955
rect 556 25923 588 25955
rect 628 25923 660 25955
rect 700 25923 732 25955
rect 772 25923 804 25955
rect 844 25923 876 25955
rect 124 25851 156 25883
rect 196 25851 228 25883
rect 268 25851 300 25883
rect 340 25851 372 25883
rect 412 25851 444 25883
rect 484 25851 516 25883
rect 556 25851 588 25883
rect 628 25851 660 25883
rect 700 25851 732 25883
rect 772 25851 804 25883
rect 844 25851 876 25883
rect 124 25779 156 25811
rect 196 25779 228 25811
rect 268 25779 300 25811
rect 340 25779 372 25811
rect 412 25779 444 25811
rect 484 25779 516 25811
rect 556 25779 588 25811
rect 628 25779 660 25811
rect 700 25779 732 25811
rect 772 25779 804 25811
rect 844 25779 876 25811
rect 124 25707 156 25739
rect 196 25707 228 25739
rect 268 25707 300 25739
rect 340 25707 372 25739
rect 412 25707 444 25739
rect 484 25707 516 25739
rect 556 25707 588 25739
rect 628 25707 660 25739
rect 700 25707 732 25739
rect 772 25707 804 25739
rect 844 25707 876 25739
rect 124 25635 156 25667
rect 196 25635 228 25667
rect 268 25635 300 25667
rect 340 25635 372 25667
rect 412 25635 444 25667
rect 484 25635 516 25667
rect 556 25635 588 25667
rect 628 25635 660 25667
rect 700 25635 732 25667
rect 772 25635 804 25667
rect 844 25635 876 25667
rect 124 25563 156 25595
rect 196 25563 228 25595
rect 268 25563 300 25595
rect 340 25563 372 25595
rect 412 25563 444 25595
rect 484 25563 516 25595
rect 556 25563 588 25595
rect 628 25563 660 25595
rect 700 25563 732 25595
rect 772 25563 804 25595
rect 844 25563 876 25595
rect 124 25491 156 25523
rect 196 25491 228 25523
rect 268 25491 300 25523
rect 340 25491 372 25523
rect 412 25491 444 25523
rect 484 25491 516 25523
rect 556 25491 588 25523
rect 628 25491 660 25523
rect 700 25491 732 25523
rect 772 25491 804 25523
rect 844 25491 876 25523
rect 124 25419 156 25451
rect 196 25419 228 25451
rect 268 25419 300 25451
rect 340 25419 372 25451
rect 412 25419 444 25451
rect 484 25419 516 25451
rect 556 25419 588 25451
rect 628 25419 660 25451
rect 700 25419 732 25451
rect 772 25419 804 25451
rect 844 25419 876 25451
rect 124 25347 156 25379
rect 196 25347 228 25379
rect 268 25347 300 25379
rect 340 25347 372 25379
rect 412 25347 444 25379
rect 484 25347 516 25379
rect 556 25347 588 25379
rect 628 25347 660 25379
rect 700 25347 732 25379
rect 772 25347 804 25379
rect 844 25347 876 25379
rect 124 25275 156 25307
rect 196 25275 228 25307
rect 268 25275 300 25307
rect 340 25275 372 25307
rect 412 25275 444 25307
rect 484 25275 516 25307
rect 556 25275 588 25307
rect 628 25275 660 25307
rect 700 25275 732 25307
rect 772 25275 804 25307
rect 844 25275 876 25307
rect 124 25203 156 25235
rect 196 25203 228 25235
rect 268 25203 300 25235
rect 340 25203 372 25235
rect 412 25203 444 25235
rect 484 25203 516 25235
rect 556 25203 588 25235
rect 628 25203 660 25235
rect 700 25203 732 25235
rect 772 25203 804 25235
rect 844 25203 876 25235
rect 124 25131 156 25163
rect 196 25131 228 25163
rect 268 25131 300 25163
rect 340 25131 372 25163
rect 412 25131 444 25163
rect 484 25131 516 25163
rect 556 25131 588 25163
rect 628 25131 660 25163
rect 700 25131 732 25163
rect 772 25131 804 25163
rect 844 25131 876 25163
rect 124 25059 156 25091
rect 196 25059 228 25091
rect 268 25059 300 25091
rect 340 25059 372 25091
rect 412 25059 444 25091
rect 484 25059 516 25091
rect 556 25059 588 25091
rect 628 25059 660 25091
rect 700 25059 732 25091
rect 772 25059 804 25091
rect 844 25059 876 25091
rect 124 24987 156 25019
rect 196 24987 228 25019
rect 268 24987 300 25019
rect 340 24987 372 25019
rect 412 24987 444 25019
rect 484 24987 516 25019
rect 556 24987 588 25019
rect 628 24987 660 25019
rect 700 24987 732 25019
rect 772 24987 804 25019
rect 844 24987 876 25019
rect 124 24915 156 24947
rect 196 24915 228 24947
rect 268 24915 300 24947
rect 340 24915 372 24947
rect 412 24915 444 24947
rect 484 24915 516 24947
rect 556 24915 588 24947
rect 628 24915 660 24947
rect 700 24915 732 24947
rect 772 24915 804 24947
rect 844 24915 876 24947
rect 124 24843 156 24875
rect 196 24843 228 24875
rect 268 24843 300 24875
rect 340 24843 372 24875
rect 412 24843 444 24875
rect 484 24843 516 24875
rect 556 24843 588 24875
rect 628 24843 660 24875
rect 700 24843 732 24875
rect 772 24843 804 24875
rect 844 24843 876 24875
rect 124 24771 156 24803
rect 196 24771 228 24803
rect 268 24771 300 24803
rect 340 24771 372 24803
rect 412 24771 444 24803
rect 484 24771 516 24803
rect 556 24771 588 24803
rect 628 24771 660 24803
rect 700 24771 732 24803
rect 772 24771 804 24803
rect 844 24771 876 24803
rect 124 24699 156 24731
rect 196 24699 228 24731
rect 268 24699 300 24731
rect 340 24699 372 24731
rect 412 24699 444 24731
rect 484 24699 516 24731
rect 556 24699 588 24731
rect 628 24699 660 24731
rect 700 24699 732 24731
rect 772 24699 804 24731
rect 844 24699 876 24731
rect 124 24627 156 24659
rect 196 24627 228 24659
rect 268 24627 300 24659
rect 340 24627 372 24659
rect 412 24627 444 24659
rect 484 24627 516 24659
rect 556 24627 588 24659
rect 628 24627 660 24659
rect 700 24627 732 24659
rect 772 24627 804 24659
rect 844 24627 876 24659
rect 124 24555 156 24587
rect 196 24555 228 24587
rect 268 24555 300 24587
rect 340 24555 372 24587
rect 412 24555 444 24587
rect 484 24555 516 24587
rect 556 24555 588 24587
rect 628 24555 660 24587
rect 700 24555 732 24587
rect 772 24555 804 24587
rect 844 24555 876 24587
rect 124 24483 156 24515
rect 196 24483 228 24515
rect 268 24483 300 24515
rect 340 24483 372 24515
rect 412 24483 444 24515
rect 484 24483 516 24515
rect 556 24483 588 24515
rect 628 24483 660 24515
rect 700 24483 732 24515
rect 772 24483 804 24515
rect 844 24483 876 24515
rect 124 24411 156 24443
rect 196 24411 228 24443
rect 268 24411 300 24443
rect 340 24411 372 24443
rect 412 24411 444 24443
rect 484 24411 516 24443
rect 556 24411 588 24443
rect 628 24411 660 24443
rect 700 24411 732 24443
rect 772 24411 804 24443
rect 844 24411 876 24443
rect 124 24339 156 24371
rect 196 24339 228 24371
rect 268 24339 300 24371
rect 340 24339 372 24371
rect 412 24339 444 24371
rect 484 24339 516 24371
rect 556 24339 588 24371
rect 628 24339 660 24371
rect 700 24339 732 24371
rect 772 24339 804 24371
rect 844 24339 876 24371
rect 124 24267 156 24299
rect 196 24267 228 24299
rect 268 24267 300 24299
rect 340 24267 372 24299
rect 412 24267 444 24299
rect 484 24267 516 24299
rect 556 24267 588 24299
rect 628 24267 660 24299
rect 700 24267 732 24299
rect 772 24267 804 24299
rect 844 24267 876 24299
rect 124 24195 156 24227
rect 196 24195 228 24227
rect 268 24195 300 24227
rect 340 24195 372 24227
rect 412 24195 444 24227
rect 484 24195 516 24227
rect 556 24195 588 24227
rect 628 24195 660 24227
rect 700 24195 732 24227
rect 772 24195 804 24227
rect 844 24195 876 24227
rect 124 24123 156 24155
rect 196 24123 228 24155
rect 268 24123 300 24155
rect 340 24123 372 24155
rect 412 24123 444 24155
rect 484 24123 516 24155
rect 556 24123 588 24155
rect 628 24123 660 24155
rect 700 24123 732 24155
rect 772 24123 804 24155
rect 844 24123 876 24155
rect 124 24051 156 24083
rect 196 24051 228 24083
rect 268 24051 300 24083
rect 340 24051 372 24083
rect 412 24051 444 24083
rect 484 24051 516 24083
rect 556 24051 588 24083
rect 628 24051 660 24083
rect 700 24051 732 24083
rect 772 24051 804 24083
rect 844 24051 876 24083
rect 124 23979 156 24011
rect 196 23979 228 24011
rect 268 23979 300 24011
rect 340 23979 372 24011
rect 412 23979 444 24011
rect 484 23979 516 24011
rect 556 23979 588 24011
rect 628 23979 660 24011
rect 700 23979 732 24011
rect 772 23979 804 24011
rect 844 23979 876 24011
rect 124 23907 156 23939
rect 196 23907 228 23939
rect 268 23907 300 23939
rect 340 23907 372 23939
rect 412 23907 444 23939
rect 484 23907 516 23939
rect 556 23907 588 23939
rect 628 23907 660 23939
rect 700 23907 732 23939
rect 772 23907 804 23939
rect 844 23907 876 23939
rect 124 23835 156 23867
rect 196 23835 228 23867
rect 268 23835 300 23867
rect 340 23835 372 23867
rect 412 23835 444 23867
rect 484 23835 516 23867
rect 556 23835 588 23867
rect 628 23835 660 23867
rect 700 23835 732 23867
rect 772 23835 804 23867
rect 844 23835 876 23867
rect 124 23763 156 23795
rect 196 23763 228 23795
rect 268 23763 300 23795
rect 340 23763 372 23795
rect 412 23763 444 23795
rect 484 23763 516 23795
rect 556 23763 588 23795
rect 628 23763 660 23795
rect 700 23763 732 23795
rect 772 23763 804 23795
rect 844 23763 876 23795
rect 124 23691 156 23723
rect 196 23691 228 23723
rect 268 23691 300 23723
rect 340 23691 372 23723
rect 412 23691 444 23723
rect 484 23691 516 23723
rect 556 23691 588 23723
rect 628 23691 660 23723
rect 700 23691 732 23723
rect 772 23691 804 23723
rect 844 23691 876 23723
rect 124 23619 156 23651
rect 196 23619 228 23651
rect 268 23619 300 23651
rect 340 23619 372 23651
rect 412 23619 444 23651
rect 484 23619 516 23651
rect 556 23619 588 23651
rect 628 23619 660 23651
rect 700 23619 732 23651
rect 772 23619 804 23651
rect 844 23619 876 23651
rect 124 23547 156 23579
rect 196 23547 228 23579
rect 268 23547 300 23579
rect 340 23547 372 23579
rect 412 23547 444 23579
rect 484 23547 516 23579
rect 556 23547 588 23579
rect 628 23547 660 23579
rect 700 23547 732 23579
rect 772 23547 804 23579
rect 844 23547 876 23579
rect 124 23475 156 23507
rect 196 23475 228 23507
rect 268 23475 300 23507
rect 340 23475 372 23507
rect 412 23475 444 23507
rect 484 23475 516 23507
rect 556 23475 588 23507
rect 628 23475 660 23507
rect 700 23475 732 23507
rect 772 23475 804 23507
rect 844 23475 876 23507
rect 124 23403 156 23435
rect 196 23403 228 23435
rect 268 23403 300 23435
rect 340 23403 372 23435
rect 412 23403 444 23435
rect 484 23403 516 23435
rect 556 23403 588 23435
rect 628 23403 660 23435
rect 700 23403 732 23435
rect 772 23403 804 23435
rect 844 23403 876 23435
rect 124 23331 156 23363
rect 196 23331 228 23363
rect 268 23331 300 23363
rect 340 23331 372 23363
rect 412 23331 444 23363
rect 484 23331 516 23363
rect 556 23331 588 23363
rect 628 23331 660 23363
rect 700 23331 732 23363
rect 772 23331 804 23363
rect 844 23331 876 23363
rect 124 23259 156 23291
rect 196 23259 228 23291
rect 268 23259 300 23291
rect 340 23259 372 23291
rect 412 23259 444 23291
rect 484 23259 516 23291
rect 556 23259 588 23291
rect 628 23259 660 23291
rect 700 23259 732 23291
rect 772 23259 804 23291
rect 844 23259 876 23291
rect 124 23187 156 23219
rect 196 23187 228 23219
rect 268 23187 300 23219
rect 340 23187 372 23219
rect 412 23187 444 23219
rect 484 23187 516 23219
rect 556 23187 588 23219
rect 628 23187 660 23219
rect 700 23187 732 23219
rect 772 23187 804 23219
rect 844 23187 876 23219
rect 196 22842 228 22874
rect 268 22842 300 22874
rect 340 22842 372 22874
rect 412 22842 444 22874
rect 484 22842 516 22874
rect 556 22842 588 22874
rect 628 22842 660 22874
rect 700 22842 732 22874
rect 772 22842 804 22874
rect 844 22842 876 22874
rect 124 22770 156 22802
rect 196 22770 228 22802
rect 268 22770 300 22802
rect 340 22770 372 22802
rect 412 22770 444 22802
rect 484 22770 516 22802
rect 556 22770 588 22802
rect 628 22770 660 22802
rect 700 22770 732 22802
rect 772 22770 804 22802
rect 844 22770 876 22802
rect 124 22698 156 22730
rect 196 22698 228 22730
rect 268 22698 300 22730
rect 340 22698 372 22730
rect 412 22698 444 22730
rect 484 22698 516 22730
rect 556 22698 588 22730
rect 628 22698 660 22730
rect 700 22698 732 22730
rect 772 22698 804 22730
rect 844 22698 876 22730
rect 124 22626 156 22658
rect 196 22626 228 22658
rect 268 22626 300 22658
rect 340 22626 372 22658
rect 412 22626 444 22658
rect 484 22626 516 22658
rect 556 22626 588 22658
rect 628 22626 660 22658
rect 700 22626 732 22658
rect 772 22626 804 22658
rect 844 22626 876 22658
rect 124 22554 156 22586
rect 196 22554 228 22586
rect 268 22554 300 22586
rect 340 22554 372 22586
rect 412 22554 444 22586
rect 484 22554 516 22586
rect 556 22554 588 22586
rect 628 22554 660 22586
rect 700 22554 732 22586
rect 772 22554 804 22586
rect 844 22554 876 22586
rect 124 22482 156 22514
rect 196 22482 228 22514
rect 268 22482 300 22514
rect 340 22482 372 22514
rect 412 22482 444 22514
rect 484 22482 516 22514
rect 556 22482 588 22514
rect 628 22482 660 22514
rect 700 22482 732 22514
rect 772 22482 804 22514
rect 844 22482 876 22514
rect 124 22410 156 22442
rect 196 22410 228 22442
rect 268 22410 300 22442
rect 340 22410 372 22442
rect 412 22410 444 22442
rect 484 22410 516 22442
rect 556 22410 588 22442
rect 628 22410 660 22442
rect 700 22410 732 22442
rect 772 22410 804 22442
rect 844 22410 876 22442
rect 124 22338 156 22370
rect 196 22338 228 22370
rect 268 22338 300 22370
rect 340 22338 372 22370
rect 412 22338 444 22370
rect 484 22338 516 22370
rect 556 22338 588 22370
rect 628 22338 660 22370
rect 700 22338 732 22370
rect 772 22338 804 22370
rect 844 22338 876 22370
rect 124 22266 156 22298
rect 196 22266 228 22298
rect 268 22266 300 22298
rect 340 22266 372 22298
rect 412 22266 444 22298
rect 484 22266 516 22298
rect 556 22266 588 22298
rect 628 22266 660 22298
rect 700 22266 732 22298
rect 772 22266 804 22298
rect 844 22266 876 22298
rect 124 22194 156 22226
rect 196 22194 228 22226
rect 268 22194 300 22226
rect 340 22194 372 22226
rect 412 22194 444 22226
rect 484 22194 516 22226
rect 556 22194 588 22226
rect 628 22194 660 22226
rect 700 22194 732 22226
rect 772 22194 804 22226
rect 844 22194 876 22226
rect 124 22122 156 22154
rect 196 22122 228 22154
rect 268 22122 300 22154
rect 340 22122 372 22154
rect 412 22122 444 22154
rect 484 22122 516 22154
rect 556 22122 588 22154
rect 628 22122 660 22154
rect 700 22122 732 22154
rect 772 22122 804 22154
rect 844 22122 876 22154
rect 124 22050 156 22082
rect 196 22050 228 22082
rect 268 22050 300 22082
rect 340 22050 372 22082
rect 412 22050 444 22082
rect 484 22050 516 22082
rect 556 22050 588 22082
rect 628 22050 660 22082
rect 700 22050 732 22082
rect 772 22050 804 22082
rect 844 22050 876 22082
rect 124 21978 156 22010
rect 196 21978 228 22010
rect 268 21978 300 22010
rect 340 21978 372 22010
rect 412 21978 444 22010
rect 484 21978 516 22010
rect 556 21978 588 22010
rect 628 21978 660 22010
rect 700 21978 732 22010
rect 772 21978 804 22010
rect 844 21978 876 22010
rect 124 21906 156 21938
rect 196 21906 228 21938
rect 268 21906 300 21938
rect 340 21906 372 21938
rect 412 21906 444 21938
rect 484 21906 516 21938
rect 556 21906 588 21938
rect 628 21906 660 21938
rect 700 21906 732 21938
rect 772 21906 804 21938
rect 844 21906 876 21938
rect 124 21834 156 21866
rect 196 21834 228 21866
rect 268 21834 300 21866
rect 340 21834 372 21866
rect 412 21834 444 21866
rect 484 21834 516 21866
rect 556 21834 588 21866
rect 628 21834 660 21866
rect 700 21834 732 21866
rect 772 21834 804 21866
rect 844 21834 876 21866
rect 124 21762 156 21794
rect 196 21762 228 21794
rect 268 21762 300 21794
rect 340 21762 372 21794
rect 412 21762 444 21794
rect 484 21762 516 21794
rect 556 21762 588 21794
rect 628 21762 660 21794
rect 700 21762 732 21794
rect 772 21762 804 21794
rect 844 21762 876 21794
rect 124 21690 156 21722
rect 196 21690 228 21722
rect 268 21690 300 21722
rect 340 21690 372 21722
rect 412 21690 444 21722
rect 484 21690 516 21722
rect 556 21690 588 21722
rect 628 21690 660 21722
rect 700 21690 732 21722
rect 772 21690 804 21722
rect 844 21690 876 21722
rect 124 21618 156 21650
rect 196 21618 228 21650
rect 268 21618 300 21650
rect 340 21618 372 21650
rect 412 21618 444 21650
rect 484 21618 516 21650
rect 556 21618 588 21650
rect 628 21618 660 21650
rect 700 21618 732 21650
rect 772 21618 804 21650
rect 844 21618 876 21650
rect 124 21546 156 21578
rect 196 21546 228 21578
rect 268 21546 300 21578
rect 340 21546 372 21578
rect 412 21546 444 21578
rect 484 21546 516 21578
rect 556 21546 588 21578
rect 628 21546 660 21578
rect 700 21546 732 21578
rect 772 21546 804 21578
rect 844 21546 876 21578
rect 124 21474 156 21506
rect 196 21474 228 21506
rect 268 21474 300 21506
rect 340 21474 372 21506
rect 412 21474 444 21506
rect 484 21474 516 21506
rect 556 21474 588 21506
rect 628 21474 660 21506
rect 700 21474 732 21506
rect 772 21474 804 21506
rect 844 21474 876 21506
rect 124 21402 156 21434
rect 196 21402 228 21434
rect 268 21402 300 21434
rect 340 21402 372 21434
rect 412 21402 444 21434
rect 484 21402 516 21434
rect 556 21402 588 21434
rect 628 21402 660 21434
rect 700 21402 732 21434
rect 772 21402 804 21434
rect 844 21402 876 21434
rect 124 21330 156 21362
rect 196 21330 228 21362
rect 268 21330 300 21362
rect 340 21330 372 21362
rect 412 21330 444 21362
rect 484 21330 516 21362
rect 556 21330 588 21362
rect 628 21330 660 21362
rect 700 21330 732 21362
rect 772 21330 804 21362
rect 844 21330 876 21362
rect 124 21258 156 21290
rect 196 21258 228 21290
rect 268 21258 300 21290
rect 340 21258 372 21290
rect 412 21258 444 21290
rect 484 21258 516 21290
rect 556 21258 588 21290
rect 628 21258 660 21290
rect 700 21258 732 21290
rect 772 21258 804 21290
rect 844 21258 876 21290
rect 124 21186 156 21218
rect 196 21186 228 21218
rect 268 21186 300 21218
rect 340 21186 372 21218
rect 412 21186 444 21218
rect 484 21186 516 21218
rect 556 21186 588 21218
rect 628 21186 660 21218
rect 700 21186 732 21218
rect 772 21186 804 21218
rect 844 21186 876 21218
rect 124 21114 156 21146
rect 196 21114 228 21146
rect 268 21114 300 21146
rect 340 21114 372 21146
rect 412 21114 444 21146
rect 484 21114 516 21146
rect 556 21114 588 21146
rect 628 21114 660 21146
rect 700 21114 732 21146
rect 772 21114 804 21146
rect 844 21114 876 21146
rect 124 21042 156 21074
rect 196 21042 228 21074
rect 268 21042 300 21074
rect 340 21042 372 21074
rect 412 21042 444 21074
rect 484 21042 516 21074
rect 556 21042 588 21074
rect 628 21042 660 21074
rect 700 21042 732 21074
rect 772 21042 804 21074
rect 844 21042 876 21074
rect 124 20970 156 21002
rect 196 20970 228 21002
rect 268 20970 300 21002
rect 340 20970 372 21002
rect 412 20970 444 21002
rect 484 20970 516 21002
rect 556 20970 588 21002
rect 628 20970 660 21002
rect 700 20970 732 21002
rect 772 20970 804 21002
rect 844 20970 876 21002
rect 124 20898 156 20930
rect 196 20898 228 20930
rect 268 20898 300 20930
rect 340 20898 372 20930
rect 412 20898 444 20930
rect 484 20898 516 20930
rect 556 20898 588 20930
rect 628 20898 660 20930
rect 700 20898 732 20930
rect 772 20898 804 20930
rect 844 20898 876 20930
rect 124 20826 156 20858
rect 196 20826 228 20858
rect 268 20826 300 20858
rect 340 20826 372 20858
rect 412 20826 444 20858
rect 484 20826 516 20858
rect 556 20826 588 20858
rect 628 20826 660 20858
rect 700 20826 732 20858
rect 772 20826 804 20858
rect 844 20826 876 20858
rect 124 20754 156 20786
rect 196 20754 228 20786
rect 268 20754 300 20786
rect 340 20754 372 20786
rect 412 20754 444 20786
rect 484 20754 516 20786
rect 556 20754 588 20786
rect 628 20754 660 20786
rect 700 20754 732 20786
rect 772 20754 804 20786
rect 844 20754 876 20786
rect 124 20682 156 20714
rect 196 20682 228 20714
rect 268 20682 300 20714
rect 340 20682 372 20714
rect 412 20682 444 20714
rect 484 20682 516 20714
rect 556 20682 588 20714
rect 628 20682 660 20714
rect 700 20682 732 20714
rect 772 20682 804 20714
rect 844 20682 876 20714
rect 124 20610 156 20642
rect 196 20610 228 20642
rect 268 20610 300 20642
rect 340 20610 372 20642
rect 412 20610 444 20642
rect 484 20610 516 20642
rect 556 20610 588 20642
rect 628 20610 660 20642
rect 700 20610 732 20642
rect 772 20610 804 20642
rect 844 20610 876 20642
rect 124 20538 156 20570
rect 196 20538 228 20570
rect 268 20538 300 20570
rect 340 20538 372 20570
rect 412 20538 444 20570
rect 484 20538 516 20570
rect 556 20538 588 20570
rect 628 20538 660 20570
rect 700 20538 732 20570
rect 772 20538 804 20570
rect 844 20538 876 20570
rect 124 20466 156 20498
rect 196 20466 228 20498
rect 268 20466 300 20498
rect 340 20466 372 20498
rect 412 20466 444 20498
rect 484 20466 516 20498
rect 556 20466 588 20498
rect 628 20466 660 20498
rect 700 20466 732 20498
rect 772 20466 804 20498
rect 844 20466 876 20498
rect 124 20394 156 20426
rect 196 20394 228 20426
rect 268 20394 300 20426
rect 340 20394 372 20426
rect 412 20394 444 20426
rect 484 20394 516 20426
rect 556 20394 588 20426
rect 628 20394 660 20426
rect 700 20394 732 20426
rect 772 20394 804 20426
rect 844 20394 876 20426
rect 124 20322 156 20354
rect 196 20322 228 20354
rect 268 20322 300 20354
rect 340 20322 372 20354
rect 412 20322 444 20354
rect 484 20322 516 20354
rect 556 20322 588 20354
rect 628 20322 660 20354
rect 700 20322 732 20354
rect 772 20322 804 20354
rect 844 20322 876 20354
rect 124 20250 156 20282
rect 196 20250 228 20282
rect 268 20250 300 20282
rect 340 20250 372 20282
rect 412 20250 444 20282
rect 484 20250 516 20282
rect 556 20250 588 20282
rect 628 20250 660 20282
rect 700 20250 732 20282
rect 772 20250 804 20282
rect 844 20250 876 20282
rect 124 20178 156 20210
rect 196 20178 228 20210
rect 268 20178 300 20210
rect 340 20178 372 20210
rect 412 20178 444 20210
rect 484 20178 516 20210
rect 556 20178 588 20210
rect 628 20178 660 20210
rect 700 20178 732 20210
rect 772 20178 804 20210
rect 844 20178 876 20210
rect 124 20106 156 20138
rect 196 20106 228 20138
rect 268 20106 300 20138
rect 340 20106 372 20138
rect 412 20106 444 20138
rect 484 20106 516 20138
rect 556 20106 588 20138
rect 628 20106 660 20138
rect 700 20106 732 20138
rect 772 20106 804 20138
rect 844 20106 876 20138
rect 124 20034 156 20066
rect 196 20034 228 20066
rect 268 20034 300 20066
rect 340 20034 372 20066
rect 412 20034 444 20066
rect 484 20034 516 20066
rect 556 20034 588 20066
rect 628 20034 660 20066
rect 700 20034 732 20066
rect 772 20034 804 20066
rect 844 20034 876 20066
rect 124 19962 156 19994
rect 196 19962 228 19994
rect 268 19962 300 19994
rect 340 19962 372 19994
rect 412 19962 444 19994
rect 484 19962 516 19994
rect 556 19962 588 19994
rect 628 19962 660 19994
rect 700 19962 732 19994
rect 772 19962 804 19994
rect 844 19962 876 19994
rect 124 19890 156 19922
rect 196 19890 228 19922
rect 268 19890 300 19922
rect 340 19890 372 19922
rect 412 19890 444 19922
rect 484 19890 516 19922
rect 556 19890 588 19922
rect 628 19890 660 19922
rect 700 19890 732 19922
rect 772 19890 804 19922
rect 844 19890 876 19922
rect 124 19818 156 19850
rect 196 19818 228 19850
rect 268 19818 300 19850
rect 340 19818 372 19850
rect 412 19818 444 19850
rect 484 19818 516 19850
rect 556 19818 588 19850
rect 628 19818 660 19850
rect 700 19818 732 19850
rect 772 19818 804 19850
rect 844 19818 876 19850
rect 124 19746 156 19778
rect 196 19746 228 19778
rect 268 19746 300 19778
rect 340 19746 372 19778
rect 412 19746 444 19778
rect 484 19746 516 19778
rect 556 19746 588 19778
rect 628 19746 660 19778
rect 700 19746 732 19778
rect 772 19746 804 19778
rect 844 19746 876 19778
rect 124 19674 156 19706
rect 196 19674 228 19706
rect 268 19674 300 19706
rect 340 19674 372 19706
rect 412 19674 444 19706
rect 484 19674 516 19706
rect 556 19674 588 19706
rect 628 19674 660 19706
rect 700 19674 732 19706
rect 772 19674 804 19706
rect 844 19674 876 19706
rect 124 19602 156 19634
rect 196 19602 228 19634
rect 268 19602 300 19634
rect 340 19602 372 19634
rect 412 19602 444 19634
rect 484 19602 516 19634
rect 556 19602 588 19634
rect 628 19602 660 19634
rect 700 19602 732 19634
rect 772 19602 804 19634
rect 844 19602 876 19634
rect 124 19530 156 19562
rect 196 19530 228 19562
rect 268 19530 300 19562
rect 340 19530 372 19562
rect 412 19530 444 19562
rect 484 19530 516 19562
rect 556 19530 588 19562
rect 628 19530 660 19562
rect 700 19530 732 19562
rect 772 19530 804 19562
rect 844 19530 876 19562
rect 124 19458 156 19490
rect 196 19458 228 19490
rect 268 19458 300 19490
rect 340 19458 372 19490
rect 412 19458 444 19490
rect 484 19458 516 19490
rect 556 19458 588 19490
rect 628 19458 660 19490
rect 700 19458 732 19490
rect 772 19458 804 19490
rect 844 19458 876 19490
rect 124 19386 156 19418
rect 196 19386 228 19418
rect 268 19386 300 19418
rect 340 19386 372 19418
rect 412 19386 444 19418
rect 484 19386 516 19418
rect 556 19386 588 19418
rect 628 19386 660 19418
rect 700 19386 732 19418
rect 772 19386 804 19418
rect 844 19386 876 19418
rect 124 19314 156 19346
rect 196 19314 228 19346
rect 268 19314 300 19346
rect 340 19314 372 19346
rect 412 19314 444 19346
rect 484 19314 516 19346
rect 556 19314 588 19346
rect 628 19314 660 19346
rect 700 19314 732 19346
rect 772 19314 804 19346
rect 844 19314 876 19346
rect 124 19242 156 19274
rect 196 19242 228 19274
rect 268 19242 300 19274
rect 340 19242 372 19274
rect 412 19242 444 19274
rect 484 19242 516 19274
rect 556 19242 588 19274
rect 628 19242 660 19274
rect 700 19242 732 19274
rect 772 19242 804 19274
rect 844 19242 876 19274
rect 124 19170 156 19202
rect 196 19170 228 19202
rect 268 19170 300 19202
rect 340 19170 372 19202
rect 412 19170 444 19202
rect 484 19170 516 19202
rect 556 19170 588 19202
rect 628 19170 660 19202
rect 700 19170 732 19202
rect 772 19170 804 19202
rect 844 19170 876 19202
rect 124 19098 156 19130
rect 196 19098 228 19130
rect 268 19098 300 19130
rect 340 19098 372 19130
rect 412 19098 444 19130
rect 484 19098 516 19130
rect 556 19098 588 19130
rect 628 19098 660 19130
rect 700 19098 732 19130
rect 772 19098 804 19130
rect 844 19098 876 19130
rect 124 19026 156 19058
rect 196 19026 228 19058
rect 268 19026 300 19058
rect 340 19026 372 19058
rect 412 19026 444 19058
rect 484 19026 516 19058
rect 556 19026 588 19058
rect 628 19026 660 19058
rect 700 19026 732 19058
rect 772 19026 804 19058
rect 844 19026 876 19058
rect 124 18954 156 18986
rect 196 18954 228 18986
rect 268 18954 300 18986
rect 340 18954 372 18986
rect 412 18954 444 18986
rect 484 18954 516 18986
rect 556 18954 588 18986
rect 628 18954 660 18986
rect 700 18954 732 18986
rect 772 18954 804 18986
rect 844 18954 876 18986
rect 124 18882 156 18914
rect 196 18882 228 18914
rect 268 18882 300 18914
rect 340 18882 372 18914
rect 412 18882 444 18914
rect 484 18882 516 18914
rect 556 18882 588 18914
rect 628 18882 660 18914
rect 700 18882 732 18914
rect 772 18882 804 18914
rect 844 18882 876 18914
rect 124 18810 156 18842
rect 196 18810 228 18842
rect 268 18810 300 18842
rect 340 18810 372 18842
rect 412 18810 444 18842
rect 484 18810 516 18842
rect 556 18810 588 18842
rect 628 18810 660 18842
rect 700 18810 732 18842
rect 772 18810 804 18842
rect 844 18810 876 18842
rect 124 18738 156 18770
rect 196 18738 228 18770
rect 268 18738 300 18770
rect 340 18738 372 18770
rect 412 18738 444 18770
rect 484 18738 516 18770
rect 556 18738 588 18770
rect 628 18738 660 18770
rect 700 18738 732 18770
rect 772 18738 804 18770
rect 844 18738 876 18770
rect 124 18666 156 18698
rect 196 18666 228 18698
rect 268 18666 300 18698
rect 340 18666 372 18698
rect 412 18666 444 18698
rect 484 18666 516 18698
rect 556 18666 588 18698
rect 628 18666 660 18698
rect 700 18666 732 18698
rect 772 18666 804 18698
rect 844 18666 876 18698
rect 124 18594 156 18626
rect 196 18594 228 18626
rect 268 18594 300 18626
rect 340 18594 372 18626
rect 412 18594 444 18626
rect 484 18594 516 18626
rect 556 18594 588 18626
rect 628 18594 660 18626
rect 700 18594 732 18626
rect 772 18594 804 18626
rect 844 18594 876 18626
rect 124 18522 156 18554
rect 196 18522 228 18554
rect 268 18522 300 18554
rect 340 18522 372 18554
rect 412 18522 444 18554
rect 484 18522 516 18554
rect 556 18522 588 18554
rect 628 18522 660 18554
rect 700 18522 732 18554
rect 772 18522 804 18554
rect 844 18522 876 18554
rect 124 18450 156 18482
rect 196 18450 228 18482
rect 268 18450 300 18482
rect 340 18450 372 18482
rect 412 18450 444 18482
rect 484 18450 516 18482
rect 556 18450 588 18482
rect 628 18450 660 18482
rect 700 18450 732 18482
rect 772 18450 804 18482
rect 844 18450 876 18482
rect 124 18378 156 18410
rect 196 18378 228 18410
rect 268 18378 300 18410
rect 340 18378 372 18410
rect 412 18378 444 18410
rect 484 18378 516 18410
rect 556 18378 588 18410
rect 628 18378 660 18410
rect 700 18378 732 18410
rect 772 18378 804 18410
rect 844 18378 876 18410
rect 124 18306 156 18338
rect 196 18306 228 18338
rect 268 18306 300 18338
rect 340 18306 372 18338
rect 412 18306 444 18338
rect 484 18306 516 18338
rect 556 18306 588 18338
rect 628 18306 660 18338
rect 700 18306 732 18338
rect 772 18306 804 18338
rect 844 18306 876 18338
rect 124 18234 156 18266
rect 196 18234 228 18266
rect 268 18234 300 18266
rect 340 18234 372 18266
rect 412 18234 444 18266
rect 484 18234 516 18266
rect 556 18234 588 18266
rect 628 18234 660 18266
rect 700 18234 732 18266
rect 772 18234 804 18266
rect 844 18234 876 18266
rect 124 18162 156 18194
rect 196 18162 228 18194
rect 268 18162 300 18194
rect 340 18162 372 18194
rect 412 18162 444 18194
rect 484 18162 516 18194
rect 556 18162 588 18194
rect 628 18162 660 18194
rect 700 18162 732 18194
rect 772 18162 804 18194
rect 844 18162 876 18194
rect 196 17816 228 17848
rect 268 17816 300 17848
rect 340 17816 372 17848
rect 412 17816 444 17848
rect 484 17816 516 17848
rect 556 17816 588 17848
rect 628 17816 660 17848
rect 700 17816 732 17848
rect 772 17816 804 17848
rect 844 17816 876 17848
rect 124 17744 156 17776
rect 196 17744 228 17776
rect 268 17744 300 17776
rect 340 17744 372 17776
rect 412 17744 444 17776
rect 484 17744 516 17776
rect 556 17744 588 17776
rect 628 17744 660 17776
rect 700 17744 732 17776
rect 772 17744 804 17776
rect 844 17744 876 17776
rect 124 17672 156 17704
rect 196 17672 228 17704
rect 268 17672 300 17704
rect 340 17672 372 17704
rect 412 17672 444 17704
rect 484 17672 516 17704
rect 556 17672 588 17704
rect 628 17672 660 17704
rect 700 17672 732 17704
rect 772 17672 804 17704
rect 844 17672 876 17704
rect 124 17600 156 17632
rect 196 17600 228 17632
rect 268 17600 300 17632
rect 340 17600 372 17632
rect 412 17600 444 17632
rect 484 17600 516 17632
rect 556 17600 588 17632
rect 628 17600 660 17632
rect 700 17600 732 17632
rect 772 17600 804 17632
rect 844 17600 876 17632
rect 124 17528 156 17560
rect 196 17528 228 17560
rect 268 17528 300 17560
rect 340 17528 372 17560
rect 412 17528 444 17560
rect 484 17528 516 17560
rect 556 17528 588 17560
rect 628 17528 660 17560
rect 700 17528 732 17560
rect 772 17528 804 17560
rect 844 17528 876 17560
rect 124 17456 156 17488
rect 196 17456 228 17488
rect 268 17456 300 17488
rect 340 17456 372 17488
rect 412 17456 444 17488
rect 484 17456 516 17488
rect 556 17456 588 17488
rect 628 17456 660 17488
rect 700 17456 732 17488
rect 772 17456 804 17488
rect 844 17456 876 17488
rect 124 17384 156 17416
rect 196 17384 228 17416
rect 268 17384 300 17416
rect 340 17384 372 17416
rect 412 17384 444 17416
rect 484 17384 516 17416
rect 556 17384 588 17416
rect 628 17384 660 17416
rect 700 17384 732 17416
rect 772 17384 804 17416
rect 844 17384 876 17416
rect 124 17312 156 17344
rect 196 17312 228 17344
rect 268 17312 300 17344
rect 340 17312 372 17344
rect 412 17312 444 17344
rect 484 17312 516 17344
rect 556 17312 588 17344
rect 628 17312 660 17344
rect 700 17312 732 17344
rect 772 17312 804 17344
rect 844 17312 876 17344
rect 124 17240 156 17272
rect 196 17240 228 17272
rect 268 17240 300 17272
rect 340 17240 372 17272
rect 412 17240 444 17272
rect 484 17240 516 17272
rect 556 17240 588 17272
rect 628 17240 660 17272
rect 700 17240 732 17272
rect 772 17240 804 17272
rect 844 17240 876 17272
rect 124 17168 156 17200
rect 196 17168 228 17200
rect 268 17168 300 17200
rect 340 17168 372 17200
rect 412 17168 444 17200
rect 484 17168 516 17200
rect 556 17168 588 17200
rect 628 17168 660 17200
rect 700 17168 732 17200
rect 772 17168 804 17200
rect 844 17168 876 17200
rect 124 17096 156 17128
rect 196 17096 228 17128
rect 268 17096 300 17128
rect 340 17096 372 17128
rect 412 17096 444 17128
rect 484 17096 516 17128
rect 556 17096 588 17128
rect 628 17096 660 17128
rect 700 17096 732 17128
rect 772 17096 804 17128
rect 844 17096 876 17128
rect 124 17024 156 17056
rect 196 17024 228 17056
rect 268 17024 300 17056
rect 340 17024 372 17056
rect 412 17024 444 17056
rect 484 17024 516 17056
rect 556 17024 588 17056
rect 628 17024 660 17056
rect 700 17024 732 17056
rect 772 17024 804 17056
rect 844 17024 876 17056
rect 124 16952 156 16984
rect 196 16952 228 16984
rect 268 16952 300 16984
rect 340 16952 372 16984
rect 412 16952 444 16984
rect 484 16952 516 16984
rect 556 16952 588 16984
rect 628 16952 660 16984
rect 700 16952 732 16984
rect 772 16952 804 16984
rect 844 16952 876 16984
rect 124 16880 156 16912
rect 196 16880 228 16912
rect 268 16880 300 16912
rect 340 16880 372 16912
rect 412 16880 444 16912
rect 484 16880 516 16912
rect 556 16880 588 16912
rect 628 16880 660 16912
rect 700 16880 732 16912
rect 772 16880 804 16912
rect 844 16880 876 16912
rect 124 16808 156 16840
rect 196 16808 228 16840
rect 268 16808 300 16840
rect 340 16808 372 16840
rect 412 16808 444 16840
rect 484 16808 516 16840
rect 556 16808 588 16840
rect 628 16808 660 16840
rect 700 16808 732 16840
rect 772 16808 804 16840
rect 844 16808 876 16840
rect 124 16736 156 16768
rect 196 16736 228 16768
rect 268 16736 300 16768
rect 340 16736 372 16768
rect 412 16736 444 16768
rect 484 16736 516 16768
rect 556 16736 588 16768
rect 628 16736 660 16768
rect 700 16736 732 16768
rect 772 16736 804 16768
rect 844 16736 876 16768
rect 124 16664 156 16696
rect 196 16664 228 16696
rect 268 16664 300 16696
rect 340 16664 372 16696
rect 412 16664 444 16696
rect 484 16664 516 16696
rect 556 16664 588 16696
rect 628 16664 660 16696
rect 700 16664 732 16696
rect 772 16664 804 16696
rect 844 16664 876 16696
rect 124 16592 156 16624
rect 196 16592 228 16624
rect 268 16592 300 16624
rect 340 16592 372 16624
rect 412 16592 444 16624
rect 484 16592 516 16624
rect 556 16592 588 16624
rect 628 16592 660 16624
rect 700 16592 732 16624
rect 772 16592 804 16624
rect 844 16592 876 16624
rect 124 16520 156 16552
rect 196 16520 228 16552
rect 268 16520 300 16552
rect 340 16520 372 16552
rect 412 16520 444 16552
rect 484 16520 516 16552
rect 556 16520 588 16552
rect 628 16520 660 16552
rect 700 16520 732 16552
rect 772 16520 804 16552
rect 844 16520 876 16552
rect 124 16448 156 16480
rect 196 16448 228 16480
rect 268 16448 300 16480
rect 340 16448 372 16480
rect 412 16448 444 16480
rect 484 16448 516 16480
rect 556 16448 588 16480
rect 628 16448 660 16480
rect 700 16448 732 16480
rect 772 16448 804 16480
rect 844 16448 876 16480
rect 124 16376 156 16408
rect 196 16376 228 16408
rect 268 16376 300 16408
rect 340 16376 372 16408
rect 412 16376 444 16408
rect 484 16376 516 16408
rect 556 16376 588 16408
rect 628 16376 660 16408
rect 700 16376 732 16408
rect 772 16376 804 16408
rect 844 16376 876 16408
rect 124 16304 156 16336
rect 196 16304 228 16336
rect 268 16304 300 16336
rect 340 16304 372 16336
rect 412 16304 444 16336
rect 484 16304 516 16336
rect 556 16304 588 16336
rect 628 16304 660 16336
rect 700 16304 732 16336
rect 772 16304 804 16336
rect 844 16304 876 16336
rect 124 16232 156 16264
rect 196 16232 228 16264
rect 268 16232 300 16264
rect 340 16232 372 16264
rect 412 16232 444 16264
rect 484 16232 516 16264
rect 556 16232 588 16264
rect 628 16232 660 16264
rect 700 16232 732 16264
rect 772 16232 804 16264
rect 844 16232 876 16264
rect 124 16160 156 16192
rect 196 16160 228 16192
rect 268 16160 300 16192
rect 340 16160 372 16192
rect 412 16160 444 16192
rect 484 16160 516 16192
rect 556 16160 588 16192
rect 628 16160 660 16192
rect 700 16160 732 16192
rect 772 16160 804 16192
rect 844 16160 876 16192
rect 124 16088 156 16120
rect 196 16088 228 16120
rect 268 16088 300 16120
rect 340 16088 372 16120
rect 412 16088 444 16120
rect 484 16088 516 16120
rect 556 16088 588 16120
rect 628 16088 660 16120
rect 700 16088 732 16120
rect 772 16088 804 16120
rect 844 16088 876 16120
rect 124 16016 156 16048
rect 196 16016 228 16048
rect 268 16016 300 16048
rect 340 16016 372 16048
rect 412 16016 444 16048
rect 484 16016 516 16048
rect 556 16016 588 16048
rect 628 16016 660 16048
rect 700 16016 732 16048
rect 772 16016 804 16048
rect 844 16016 876 16048
rect 124 15944 156 15976
rect 196 15944 228 15976
rect 268 15944 300 15976
rect 340 15944 372 15976
rect 412 15944 444 15976
rect 484 15944 516 15976
rect 556 15944 588 15976
rect 628 15944 660 15976
rect 700 15944 732 15976
rect 772 15944 804 15976
rect 844 15944 876 15976
rect 124 15872 156 15904
rect 196 15872 228 15904
rect 268 15872 300 15904
rect 340 15872 372 15904
rect 412 15872 444 15904
rect 484 15872 516 15904
rect 556 15872 588 15904
rect 628 15872 660 15904
rect 700 15872 732 15904
rect 772 15872 804 15904
rect 844 15872 876 15904
rect 124 15800 156 15832
rect 196 15800 228 15832
rect 268 15800 300 15832
rect 340 15800 372 15832
rect 412 15800 444 15832
rect 484 15800 516 15832
rect 556 15800 588 15832
rect 628 15800 660 15832
rect 700 15800 732 15832
rect 772 15800 804 15832
rect 844 15800 876 15832
rect 124 15728 156 15760
rect 196 15728 228 15760
rect 268 15728 300 15760
rect 340 15728 372 15760
rect 412 15728 444 15760
rect 484 15728 516 15760
rect 556 15728 588 15760
rect 628 15728 660 15760
rect 700 15728 732 15760
rect 772 15728 804 15760
rect 844 15728 876 15760
rect 124 15656 156 15688
rect 196 15656 228 15688
rect 268 15656 300 15688
rect 340 15656 372 15688
rect 412 15656 444 15688
rect 484 15656 516 15688
rect 556 15656 588 15688
rect 628 15656 660 15688
rect 700 15656 732 15688
rect 772 15656 804 15688
rect 844 15656 876 15688
rect 124 15584 156 15616
rect 196 15584 228 15616
rect 268 15584 300 15616
rect 340 15584 372 15616
rect 412 15584 444 15616
rect 484 15584 516 15616
rect 556 15584 588 15616
rect 628 15584 660 15616
rect 700 15584 732 15616
rect 772 15584 804 15616
rect 844 15584 876 15616
rect 124 15512 156 15544
rect 196 15512 228 15544
rect 268 15512 300 15544
rect 340 15512 372 15544
rect 412 15512 444 15544
rect 484 15512 516 15544
rect 556 15512 588 15544
rect 628 15512 660 15544
rect 700 15512 732 15544
rect 772 15512 804 15544
rect 844 15512 876 15544
rect 124 15440 156 15472
rect 196 15440 228 15472
rect 268 15440 300 15472
rect 340 15440 372 15472
rect 412 15440 444 15472
rect 484 15440 516 15472
rect 556 15440 588 15472
rect 628 15440 660 15472
rect 700 15440 732 15472
rect 772 15440 804 15472
rect 844 15440 876 15472
rect 124 15368 156 15400
rect 196 15368 228 15400
rect 268 15368 300 15400
rect 340 15368 372 15400
rect 412 15368 444 15400
rect 484 15368 516 15400
rect 556 15368 588 15400
rect 628 15368 660 15400
rect 700 15368 732 15400
rect 772 15368 804 15400
rect 844 15368 876 15400
rect 124 15296 156 15328
rect 196 15296 228 15328
rect 268 15296 300 15328
rect 340 15296 372 15328
rect 412 15296 444 15328
rect 484 15296 516 15328
rect 556 15296 588 15328
rect 628 15296 660 15328
rect 700 15296 732 15328
rect 772 15296 804 15328
rect 844 15296 876 15328
rect 124 15224 156 15256
rect 196 15224 228 15256
rect 268 15224 300 15256
rect 340 15224 372 15256
rect 412 15224 444 15256
rect 484 15224 516 15256
rect 556 15224 588 15256
rect 628 15224 660 15256
rect 700 15224 732 15256
rect 772 15224 804 15256
rect 844 15224 876 15256
rect 124 15152 156 15184
rect 196 15152 228 15184
rect 268 15152 300 15184
rect 340 15152 372 15184
rect 412 15152 444 15184
rect 484 15152 516 15184
rect 556 15152 588 15184
rect 628 15152 660 15184
rect 700 15152 732 15184
rect 772 15152 804 15184
rect 844 15152 876 15184
rect 124 15080 156 15112
rect 196 15080 228 15112
rect 268 15080 300 15112
rect 340 15080 372 15112
rect 412 15080 444 15112
rect 484 15080 516 15112
rect 556 15080 588 15112
rect 628 15080 660 15112
rect 700 15080 732 15112
rect 772 15080 804 15112
rect 844 15080 876 15112
rect 124 15008 156 15040
rect 196 15008 228 15040
rect 268 15008 300 15040
rect 340 15008 372 15040
rect 412 15008 444 15040
rect 484 15008 516 15040
rect 556 15008 588 15040
rect 628 15008 660 15040
rect 700 15008 732 15040
rect 772 15008 804 15040
rect 844 15008 876 15040
rect 124 14936 156 14968
rect 196 14936 228 14968
rect 268 14936 300 14968
rect 340 14936 372 14968
rect 412 14936 444 14968
rect 484 14936 516 14968
rect 556 14936 588 14968
rect 628 14936 660 14968
rect 700 14936 732 14968
rect 772 14936 804 14968
rect 844 14936 876 14968
rect 124 14864 156 14896
rect 196 14864 228 14896
rect 268 14864 300 14896
rect 340 14864 372 14896
rect 412 14864 444 14896
rect 484 14864 516 14896
rect 556 14864 588 14896
rect 628 14864 660 14896
rect 700 14864 732 14896
rect 772 14864 804 14896
rect 844 14864 876 14896
rect 124 14792 156 14824
rect 196 14792 228 14824
rect 268 14792 300 14824
rect 340 14792 372 14824
rect 412 14792 444 14824
rect 484 14792 516 14824
rect 556 14792 588 14824
rect 628 14792 660 14824
rect 700 14792 732 14824
rect 772 14792 804 14824
rect 844 14792 876 14824
rect 124 14720 156 14752
rect 196 14720 228 14752
rect 268 14720 300 14752
rect 340 14720 372 14752
rect 412 14720 444 14752
rect 484 14720 516 14752
rect 556 14720 588 14752
rect 628 14720 660 14752
rect 700 14720 732 14752
rect 772 14720 804 14752
rect 844 14720 876 14752
rect 124 14648 156 14680
rect 196 14648 228 14680
rect 268 14648 300 14680
rect 340 14648 372 14680
rect 412 14648 444 14680
rect 484 14648 516 14680
rect 556 14648 588 14680
rect 628 14648 660 14680
rect 700 14648 732 14680
rect 772 14648 804 14680
rect 844 14648 876 14680
rect 124 14576 156 14608
rect 196 14576 228 14608
rect 268 14576 300 14608
rect 340 14576 372 14608
rect 412 14576 444 14608
rect 484 14576 516 14608
rect 556 14576 588 14608
rect 628 14576 660 14608
rect 700 14576 732 14608
rect 772 14576 804 14608
rect 844 14576 876 14608
rect 124 14504 156 14536
rect 196 14504 228 14536
rect 268 14504 300 14536
rect 340 14504 372 14536
rect 412 14504 444 14536
rect 484 14504 516 14536
rect 556 14504 588 14536
rect 628 14504 660 14536
rect 700 14504 732 14536
rect 772 14504 804 14536
rect 844 14504 876 14536
rect 124 14432 156 14464
rect 196 14432 228 14464
rect 268 14432 300 14464
rect 340 14432 372 14464
rect 412 14432 444 14464
rect 484 14432 516 14464
rect 556 14432 588 14464
rect 628 14432 660 14464
rect 700 14432 732 14464
rect 772 14432 804 14464
rect 844 14432 876 14464
rect 124 14360 156 14392
rect 196 14360 228 14392
rect 268 14360 300 14392
rect 340 14360 372 14392
rect 412 14360 444 14392
rect 484 14360 516 14392
rect 556 14360 588 14392
rect 628 14360 660 14392
rect 700 14360 732 14392
rect 772 14360 804 14392
rect 844 14360 876 14392
rect 124 14288 156 14320
rect 196 14288 228 14320
rect 268 14288 300 14320
rect 340 14288 372 14320
rect 412 14288 444 14320
rect 484 14288 516 14320
rect 556 14288 588 14320
rect 628 14288 660 14320
rect 700 14288 732 14320
rect 772 14288 804 14320
rect 844 14288 876 14320
rect 124 14216 156 14248
rect 196 14216 228 14248
rect 268 14216 300 14248
rect 340 14216 372 14248
rect 412 14216 444 14248
rect 484 14216 516 14248
rect 556 14216 588 14248
rect 628 14216 660 14248
rect 700 14216 732 14248
rect 772 14216 804 14248
rect 844 14216 876 14248
rect 124 14144 156 14176
rect 196 14144 228 14176
rect 268 14144 300 14176
rect 340 14144 372 14176
rect 412 14144 444 14176
rect 484 14144 516 14176
rect 556 14144 588 14176
rect 628 14144 660 14176
rect 700 14144 732 14176
rect 772 14144 804 14176
rect 844 14144 876 14176
rect 124 14072 156 14104
rect 196 14072 228 14104
rect 268 14072 300 14104
rect 340 14072 372 14104
rect 412 14072 444 14104
rect 484 14072 516 14104
rect 556 14072 588 14104
rect 628 14072 660 14104
rect 700 14072 732 14104
rect 772 14072 804 14104
rect 844 14072 876 14104
rect 124 14000 156 14032
rect 196 14000 228 14032
rect 268 14000 300 14032
rect 340 14000 372 14032
rect 412 14000 444 14032
rect 484 14000 516 14032
rect 556 14000 588 14032
rect 628 14000 660 14032
rect 700 14000 732 14032
rect 772 14000 804 14032
rect 844 14000 876 14032
rect 124 13928 156 13960
rect 196 13928 228 13960
rect 268 13928 300 13960
rect 340 13928 372 13960
rect 412 13928 444 13960
rect 484 13928 516 13960
rect 556 13928 588 13960
rect 628 13928 660 13960
rect 700 13928 732 13960
rect 772 13928 804 13960
rect 844 13928 876 13960
rect 124 13856 156 13888
rect 196 13856 228 13888
rect 268 13856 300 13888
rect 340 13856 372 13888
rect 412 13856 444 13888
rect 484 13856 516 13888
rect 556 13856 588 13888
rect 628 13856 660 13888
rect 700 13856 732 13888
rect 772 13856 804 13888
rect 844 13856 876 13888
rect 124 13784 156 13816
rect 196 13784 228 13816
rect 268 13784 300 13816
rect 340 13784 372 13816
rect 412 13784 444 13816
rect 484 13784 516 13816
rect 556 13784 588 13816
rect 628 13784 660 13816
rect 700 13784 732 13816
rect 772 13784 804 13816
rect 844 13784 876 13816
rect 124 13712 156 13744
rect 196 13712 228 13744
rect 268 13712 300 13744
rect 340 13712 372 13744
rect 412 13712 444 13744
rect 484 13712 516 13744
rect 556 13712 588 13744
rect 628 13712 660 13744
rect 700 13712 732 13744
rect 772 13712 804 13744
rect 844 13712 876 13744
rect 124 13640 156 13672
rect 196 13640 228 13672
rect 268 13640 300 13672
rect 340 13640 372 13672
rect 412 13640 444 13672
rect 484 13640 516 13672
rect 556 13640 588 13672
rect 628 13640 660 13672
rect 700 13640 732 13672
rect 772 13640 804 13672
rect 844 13640 876 13672
rect 124 13568 156 13600
rect 196 13568 228 13600
rect 268 13568 300 13600
rect 340 13568 372 13600
rect 412 13568 444 13600
rect 484 13568 516 13600
rect 556 13568 588 13600
rect 628 13568 660 13600
rect 700 13568 732 13600
rect 772 13568 804 13600
rect 844 13568 876 13600
rect 124 13496 156 13528
rect 196 13496 228 13528
rect 268 13496 300 13528
rect 340 13496 372 13528
rect 412 13496 444 13528
rect 484 13496 516 13528
rect 556 13496 588 13528
rect 628 13496 660 13528
rect 700 13496 732 13528
rect 772 13496 804 13528
rect 844 13496 876 13528
rect 124 13424 156 13456
rect 196 13424 228 13456
rect 268 13424 300 13456
rect 340 13424 372 13456
rect 412 13424 444 13456
rect 484 13424 516 13456
rect 556 13424 588 13456
rect 628 13424 660 13456
rect 700 13424 732 13456
rect 772 13424 804 13456
rect 844 13424 876 13456
rect 124 13352 156 13384
rect 196 13352 228 13384
rect 268 13352 300 13384
rect 340 13352 372 13384
rect 412 13352 444 13384
rect 484 13352 516 13384
rect 556 13352 588 13384
rect 628 13352 660 13384
rect 700 13352 732 13384
rect 772 13352 804 13384
rect 844 13352 876 13384
rect 124 13280 156 13312
rect 196 13280 228 13312
rect 268 13280 300 13312
rect 340 13280 372 13312
rect 412 13280 444 13312
rect 484 13280 516 13312
rect 556 13280 588 13312
rect 628 13280 660 13312
rect 700 13280 732 13312
rect 772 13280 804 13312
rect 844 13280 876 13312
rect 124 13208 156 13240
rect 196 13208 228 13240
rect 268 13208 300 13240
rect 340 13208 372 13240
rect 412 13208 444 13240
rect 484 13208 516 13240
rect 556 13208 588 13240
rect 628 13208 660 13240
rect 700 13208 732 13240
rect 772 13208 804 13240
rect 844 13208 876 13240
rect 124 13136 156 13168
rect 196 13136 228 13168
rect 268 13136 300 13168
rect 340 13136 372 13168
rect 412 13136 444 13168
rect 484 13136 516 13168
rect 556 13136 588 13168
rect 628 13136 660 13168
rect 700 13136 732 13168
rect 772 13136 804 13168
rect 844 13136 876 13168
rect 124 13064 156 13096
rect 196 13064 228 13096
rect 268 13064 300 13096
rect 340 13064 372 13096
rect 412 13064 444 13096
rect 484 13064 516 13096
rect 556 13064 588 13096
rect 628 13064 660 13096
rect 700 13064 732 13096
rect 772 13064 804 13096
rect 844 13064 876 13096
rect 0 33384 124 33416
rect 156 33384 196 33416
rect 228 33384 268 33416
rect 300 33384 340 33416
rect 372 33384 412 33416
rect 444 33384 484 33416
rect 516 33384 556 33416
rect 588 33384 628 33416
rect 660 33384 700 33416
rect 732 33384 772 33416
rect 804 33384 844 33416
rect 876 33384 1000 33416
rect 0 31384 223 31416
rect 255 31384 292 31416
rect 324 31384 362 31416
rect 394 31384 431 31416
rect 463 31384 502 31416
rect 534 31384 572 31416
rect 604 31384 640 31416
rect 672 31384 710 31416
rect 742 31384 1000 31416
rect 0 29684 124 29716
rect 156 29684 196 29716
rect 228 29684 268 29716
rect 300 29684 340 29716
rect 372 29684 412 29716
rect 444 29684 484 29716
rect 516 29684 556 29716
rect 588 29684 628 29716
rect 660 29684 700 29716
rect 732 29684 772 29716
rect 804 29684 844 29716
rect 876 29684 1000 29716
rect 0 27971 1000 28034
rect 0 27939 124 27971
rect 156 27939 196 27971
rect 228 27939 268 27971
rect 300 27939 340 27971
rect 372 27939 412 27971
rect 444 27939 484 27971
rect 516 27939 556 27971
rect 588 27939 628 27971
rect 660 27939 700 27971
rect 732 27939 772 27971
rect 804 27939 844 27971
rect 876 27939 1000 27971
rect 0 27899 1000 27939
rect 0 27867 124 27899
rect 156 27867 196 27899
rect 228 27867 268 27899
rect 300 27867 340 27899
rect 372 27867 412 27899
rect 444 27867 484 27899
rect 516 27867 556 27899
rect 588 27867 628 27899
rect 660 27867 700 27899
rect 732 27867 772 27899
rect 804 27867 844 27899
rect 876 27867 1000 27899
rect 0 27827 1000 27867
rect 0 27795 124 27827
rect 156 27795 196 27827
rect 228 27795 268 27827
rect 300 27795 340 27827
rect 372 27795 412 27827
rect 444 27795 484 27827
rect 516 27795 556 27827
rect 588 27795 628 27827
rect 660 27795 700 27827
rect 732 27795 772 27827
rect 804 27795 844 27827
rect 876 27795 1000 27827
rect 0 27755 1000 27795
rect 0 27723 124 27755
rect 156 27723 196 27755
rect 228 27723 268 27755
rect 300 27723 340 27755
rect 372 27723 412 27755
rect 444 27723 484 27755
rect 516 27723 556 27755
rect 588 27723 628 27755
rect 660 27723 700 27755
rect 732 27723 772 27755
rect 804 27723 844 27755
rect 876 27723 1000 27755
rect 0 27683 1000 27723
rect 0 27651 124 27683
rect 156 27651 196 27683
rect 228 27651 268 27683
rect 300 27651 340 27683
rect 372 27651 412 27683
rect 444 27651 484 27683
rect 516 27651 556 27683
rect 588 27651 628 27683
rect 660 27651 700 27683
rect 732 27651 772 27683
rect 804 27651 844 27683
rect 876 27651 1000 27683
rect 0 27611 1000 27651
rect 0 27579 124 27611
rect 156 27579 196 27611
rect 228 27579 268 27611
rect 300 27579 340 27611
rect 372 27579 412 27611
rect 444 27579 484 27611
rect 516 27579 556 27611
rect 588 27579 628 27611
rect 660 27579 700 27611
rect 732 27579 772 27611
rect 804 27579 844 27611
rect 876 27579 1000 27611
rect 0 27539 1000 27579
rect 0 27507 124 27539
rect 156 27507 196 27539
rect 228 27507 268 27539
rect 300 27507 340 27539
rect 372 27507 412 27539
rect 444 27507 484 27539
rect 516 27507 556 27539
rect 588 27507 628 27539
rect 660 27507 700 27539
rect 732 27507 772 27539
rect 804 27507 844 27539
rect 876 27507 1000 27539
rect 0 27467 1000 27507
rect 0 27435 124 27467
rect 156 27435 196 27467
rect 228 27435 268 27467
rect 300 27435 340 27467
rect 372 27435 412 27467
rect 444 27435 484 27467
rect 516 27435 556 27467
rect 588 27435 628 27467
rect 660 27435 700 27467
rect 732 27435 772 27467
rect 804 27435 844 27467
rect 876 27435 1000 27467
rect 0 27395 1000 27435
rect 0 27363 124 27395
rect 156 27363 196 27395
rect 228 27363 268 27395
rect 300 27363 340 27395
rect 372 27363 412 27395
rect 444 27363 484 27395
rect 516 27363 556 27395
rect 588 27363 628 27395
rect 660 27363 700 27395
rect 732 27363 772 27395
rect 804 27363 844 27395
rect 876 27363 1000 27395
rect 0 27323 1000 27363
rect 0 27291 124 27323
rect 156 27291 196 27323
rect 228 27291 268 27323
rect 300 27291 340 27323
rect 372 27291 412 27323
rect 444 27291 484 27323
rect 516 27291 556 27323
rect 588 27291 628 27323
rect 660 27291 700 27323
rect 732 27291 772 27323
rect 804 27291 844 27323
rect 876 27291 1000 27323
rect 0 27251 1000 27291
rect 0 27219 124 27251
rect 156 27219 196 27251
rect 228 27219 268 27251
rect 300 27219 340 27251
rect 372 27219 412 27251
rect 444 27219 484 27251
rect 516 27219 556 27251
rect 588 27219 628 27251
rect 660 27219 700 27251
rect 732 27219 772 27251
rect 804 27219 844 27251
rect 876 27219 1000 27251
rect 0 27179 1000 27219
rect 0 27147 124 27179
rect 156 27147 196 27179
rect 228 27147 268 27179
rect 300 27147 340 27179
rect 372 27147 412 27179
rect 444 27147 484 27179
rect 516 27147 556 27179
rect 588 27147 628 27179
rect 660 27147 700 27179
rect 732 27147 772 27179
rect 804 27147 844 27179
rect 876 27147 1000 27179
rect 0 27107 1000 27147
rect 0 27075 124 27107
rect 156 27075 196 27107
rect 228 27075 268 27107
rect 300 27075 340 27107
rect 372 27075 412 27107
rect 444 27075 484 27107
rect 516 27075 556 27107
rect 588 27075 628 27107
rect 660 27075 700 27107
rect 732 27075 772 27107
rect 804 27075 844 27107
rect 876 27075 1000 27107
rect 0 27035 1000 27075
rect 0 27003 124 27035
rect 156 27003 196 27035
rect 228 27003 268 27035
rect 300 27003 340 27035
rect 372 27003 412 27035
rect 444 27003 484 27035
rect 516 27003 556 27035
rect 588 27003 628 27035
rect 660 27003 700 27035
rect 732 27003 772 27035
rect 804 27003 844 27035
rect 876 27003 1000 27035
rect 0 26963 1000 27003
rect 0 26931 124 26963
rect 156 26931 196 26963
rect 228 26931 268 26963
rect 300 26931 340 26963
rect 372 26931 412 26963
rect 444 26931 484 26963
rect 516 26931 556 26963
rect 588 26931 628 26963
rect 660 26931 700 26963
rect 732 26931 772 26963
rect 804 26931 844 26963
rect 876 26931 1000 26963
rect 0 26891 1000 26931
rect 0 26859 124 26891
rect 156 26859 196 26891
rect 228 26859 268 26891
rect 300 26859 340 26891
rect 372 26859 412 26891
rect 444 26859 484 26891
rect 516 26859 556 26891
rect 588 26859 628 26891
rect 660 26859 700 26891
rect 732 26859 772 26891
rect 804 26859 844 26891
rect 876 26859 1000 26891
rect 0 26819 1000 26859
rect 0 26787 124 26819
rect 156 26787 196 26819
rect 228 26787 268 26819
rect 300 26787 340 26819
rect 372 26787 412 26819
rect 444 26787 484 26819
rect 516 26787 556 26819
rect 588 26787 628 26819
rect 660 26787 700 26819
rect 732 26787 772 26819
rect 804 26787 844 26819
rect 876 26787 1000 26819
rect 0 26747 1000 26787
rect 0 26715 124 26747
rect 156 26715 196 26747
rect 228 26715 268 26747
rect 300 26715 340 26747
rect 372 26715 412 26747
rect 444 26715 484 26747
rect 516 26715 556 26747
rect 588 26715 628 26747
rect 660 26715 700 26747
rect 732 26715 772 26747
rect 804 26715 844 26747
rect 876 26715 1000 26747
rect 0 26675 1000 26715
rect 0 26643 124 26675
rect 156 26643 196 26675
rect 228 26643 268 26675
rect 300 26643 340 26675
rect 372 26643 412 26675
rect 444 26643 484 26675
rect 516 26643 556 26675
rect 588 26643 628 26675
rect 660 26643 700 26675
rect 732 26643 772 26675
rect 804 26643 844 26675
rect 876 26643 1000 26675
rect 0 26603 1000 26643
rect 0 26571 124 26603
rect 156 26571 196 26603
rect 228 26571 268 26603
rect 300 26571 340 26603
rect 372 26571 412 26603
rect 444 26571 484 26603
rect 516 26571 556 26603
rect 588 26571 628 26603
rect 660 26571 700 26603
rect 732 26571 772 26603
rect 804 26571 844 26603
rect 876 26571 1000 26603
rect 0 26531 1000 26571
rect 0 26499 124 26531
rect 156 26499 196 26531
rect 228 26499 268 26531
rect 300 26499 340 26531
rect 372 26499 412 26531
rect 444 26499 484 26531
rect 516 26499 556 26531
rect 588 26499 628 26531
rect 660 26499 700 26531
rect 732 26499 772 26531
rect 804 26499 844 26531
rect 876 26499 1000 26531
rect 0 26459 1000 26499
rect 0 26427 124 26459
rect 156 26427 196 26459
rect 228 26427 268 26459
rect 300 26427 340 26459
rect 372 26427 412 26459
rect 444 26427 484 26459
rect 516 26427 556 26459
rect 588 26427 628 26459
rect 660 26427 700 26459
rect 732 26427 772 26459
rect 804 26427 844 26459
rect 876 26427 1000 26459
rect 0 26387 1000 26427
rect 0 26355 124 26387
rect 156 26355 196 26387
rect 228 26355 268 26387
rect 300 26355 340 26387
rect 372 26355 412 26387
rect 444 26355 484 26387
rect 516 26355 556 26387
rect 588 26355 628 26387
rect 660 26355 700 26387
rect 732 26355 772 26387
rect 804 26355 844 26387
rect 876 26355 1000 26387
rect 0 26315 1000 26355
rect 0 26283 124 26315
rect 156 26283 196 26315
rect 228 26283 268 26315
rect 300 26283 340 26315
rect 372 26283 412 26315
rect 444 26283 484 26315
rect 516 26283 556 26315
rect 588 26283 628 26315
rect 660 26283 700 26315
rect 732 26283 772 26315
rect 804 26283 844 26315
rect 876 26283 1000 26315
rect 0 26243 1000 26283
rect 0 26211 124 26243
rect 156 26211 196 26243
rect 228 26211 268 26243
rect 300 26211 340 26243
rect 372 26211 412 26243
rect 444 26211 484 26243
rect 516 26211 556 26243
rect 588 26211 628 26243
rect 660 26211 700 26243
rect 732 26211 772 26243
rect 804 26211 844 26243
rect 876 26211 1000 26243
rect 0 26171 1000 26211
rect 0 26139 124 26171
rect 156 26139 196 26171
rect 228 26139 268 26171
rect 300 26139 340 26171
rect 372 26139 412 26171
rect 444 26139 484 26171
rect 516 26139 556 26171
rect 588 26139 628 26171
rect 660 26139 700 26171
rect 732 26139 772 26171
rect 804 26139 844 26171
rect 876 26139 1000 26171
rect 0 26099 1000 26139
rect 0 26067 124 26099
rect 156 26067 196 26099
rect 228 26067 268 26099
rect 300 26067 340 26099
rect 372 26067 412 26099
rect 444 26067 484 26099
rect 516 26067 556 26099
rect 588 26067 628 26099
rect 660 26067 700 26099
rect 732 26067 772 26099
rect 804 26067 844 26099
rect 876 26067 1000 26099
rect 0 26027 1000 26067
rect 0 25995 124 26027
rect 156 25995 196 26027
rect 228 25995 268 26027
rect 300 25995 340 26027
rect 372 25995 412 26027
rect 444 25995 484 26027
rect 516 25995 556 26027
rect 588 25995 628 26027
rect 660 25995 700 26027
rect 732 25995 772 26027
rect 804 25995 844 26027
rect 876 25995 1000 26027
rect 0 25955 1000 25995
rect 0 25923 124 25955
rect 156 25923 196 25955
rect 228 25923 268 25955
rect 300 25923 340 25955
rect 372 25923 412 25955
rect 444 25923 484 25955
rect 516 25923 556 25955
rect 588 25923 628 25955
rect 660 25923 700 25955
rect 732 25923 772 25955
rect 804 25923 844 25955
rect 876 25923 1000 25955
rect 0 25883 1000 25923
rect 0 25851 124 25883
rect 156 25851 196 25883
rect 228 25851 268 25883
rect 300 25851 340 25883
rect 372 25851 412 25883
rect 444 25851 484 25883
rect 516 25851 556 25883
rect 588 25851 628 25883
rect 660 25851 700 25883
rect 732 25851 772 25883
rect 804 25851 844 25883
rect 876 25851 1000 25883
rect 0 25811 1000 25851
rect 0 25779 124 25811
rect 156 25779 196 25811
rect 228 25779 268 25811
rect 300 25779 340 25811
rect 372 25779 412 25811
rect 444 25779 484 25811
rect 516 25779 556 25811
rect 588 25779 628 25811
rect 660 25779 700 25811
rect 732 25779 772 25811
rect 804 25779 844 25811
rect 876 25779 1000 25811
rect 0 25739 1000 25779
rect 0 25707 124 25739
rect 156 25707 196 25739
rect 228 25707 268 25739
rect 300 25707 340 25739
rect 372 25707 412 25739
rect 444 25707 484 25739
rect 516 25707 556 25739
rect 588 25707 628 25739
rect 660 25707 700 25739
rect 732 25707 772 25739
rect 804 25707 844 25739
rect 876 25707 1000 25739
rect 0 25667 1000 25707
rect 0 25635 124 25667
rect 156 25635 196 25667
rect 228 25635 268 25667
rect 300 25635 340 25667
rect 372 25635 412 25667
rect 444 25635 484 25667
rect 516 25635 556 25667
rect 588 25635 628 25667
rect 660 25635 700 25667
rect 732 25635 772 25667
rect 804 25635 844 25667
rect 876 25635 1000 25667
rect 0 25595 1000 25635
rect 0 25563 124 25595
rect 156 25563 196 25595
rect 228 25563 268 25595
rect 300 25563 340 25595
rect 372 25563 412 25595
rect 444 25563 484 25595
rect 516 25563 556 25595
rect 588 25563 628 25595
rect 660 25563 700 25595
rect 732 25563 772 25595
rect 804 25563 844 25595
rect 876 25563 1000 25595
rect 0 25523 1000 25563
rect 0 25491 124 25523
rect 156 25491 196 25523
rect 228 25491 268 25523
rect 300 25491 340 25523
rect 372 25491 412 25523
rect 444 25491 484 25523
rect 516 25491 556 25523
rect 588 25491 628 25523
rect 660 25491 700 25523
rect 732 25491 772 25523
rect 804 25491 844 25523
rect 876 25491 1000 25523
rect 0 25451 1000 25491
rect 0 25419 124 25451
rect 156 25419 196 25451
rect 228 25419 268 25451
rect 300 25419 340 25451
rect 372 25419 412 25451
rect 444 25419 484 25451
rect 516 25419 556 25451
rect 588 25419 628 25451
rect 660 25419 700 25451
rect 732 25419 772 25451
rect 804 25419 844 25451
rect 876 25419 1000 25451
rect 0 25379 1000 25419
rect 0 25347 124 25379
rect 156 25347 196 25379
rect 228 25347 268 25379
rect 300 25347 340 25379
rect 372 25347 412 25379
rect 444 25347 484 25379
rect 516 25347 556 25379
rect 588 25347 628 25379
rect 660 25347 700 25379
rect 732 25347 772 25379
rect 804 25347 844 25379
rect 876 25347 1000 25379
rect 0 25307 1000 25347
rect 0 25275 124 25307
rect 156 25275 196 25307
rect 228 25275 268 25307
rect 300 25275 340 25307
rect 372 25275 412 25307
rect 444 25275 484 25307
rect 516 25275 556 25307
rect 588 25275 628 25307
rect 660 25275 700 25307
rect 732 25275 772 25307
rect 804 25275 844 25307
rect 876 25275 1000 25307
rect 0 25235 1000 25275
rect 0 25203 124 25235
rect 156 25203 196 25235
rect 228 25203 268 25235
rect 300 25203 340 25235
rect 372 25203 412 25235
rect 444 25203 484 25235
rect 516 25203 556 25235
rect 588 25203 628 25235
rect 660 25203 700 25235
rect 732 25203 772 25235
rect 804 25203 844 25235
rect 876 25203 1000 25235
rect 0 25163 1000 25203
rect 0 25131 124 25163
rect 156 25131 196 25163
rect 228 25131 268 25163
rect 300 25131 340 25163
rect 372 25131 412 25163
rect 444 25131 484 25163
rect 516 25131 556 25163
rect 588 25131 628 25163
rect 660 25131 700 25163
rect 732 25131 772 25163
rect 804 25131 844 25163
rect 876 25131 1000 25163
rect 0 25091 1000 25131
rect 0 25059 124 25091
rect 156 25059 196 25091
rect 228 25059 268 25091
rect 300 25059 340 25091
rect 372 25059 412 25091
rect 444 25059 484 25091
rect 516 25059 556 25091
rect 588 25059 628 25091
rect 660 25059 700 25091
rect 732 25059 772 25091
rect 804 25059 844 25091
rect 876 25059 1000 25091
rect 0 25019 1000 25059
rect 0 24987 124 25019
rect 156 24987 196 25019
rect 228 24987 268 25019
rect 300 24987 340 25019
rect 372 24987 412 25019
rect 444 24987 484 25019
rect 516 24987 556 25019
rect 588 24987 628 25019
rect 660 24987 700 25019
rect 732 24987 772 25019
rect 804 24987 844 25019
rect 876 24987 1000 25019
rect 0 24947 1000 24987
rect 0 24915 124 24947
rect 156 24915 196 24947
rect 228 24915 268 24947
rect 300 24915 340 24947
rect 372 24915 412 24947
rect 444 24915 484 24947
rect 516 24915 556 24947
rect 588 24915 628 24947
rect 660 24915 700 24947
rect 732 24915 772 24947
rect 804 24915 844 24947
rect 876 24915 1000 24947
rect 0 24875 1000 24915
rect 0 24843 124 24875
rect 156 24843 196 24875
rect 228 24843 268 24875
rect 300 24843 340 24875
rect 372 24843 412 24875
rect 444 24843 484 24875
rect 516 24843 556 24875
rect 588 24843 628 24875
rect 660 24843 700 24875
rect 732 24843 772 24875
rect 804 24843 844 24875
rect 876 24843 1000 24875
rect 0 24803 1000 24843
rect 0 24771 124 24803
rect 156 24771 196 24803
rect 228 24771 268 24803
rect 300 24771 340 24803
rect 372 24771 412 24803
rect 444 24771 484 24803
rect 516 24771 556 24803
rect 588 24771 628 24803
rect 660 24771 700 24803
rect 732 24771 772 24803
rect 804 24771 844 24803
rect 876 24771 1000 24803
rect 0 24731 1000 24771
rect 0 24699 124 24731
rect 156 24699 196 24731
rect 228 24699 268 24731
rect 300 24699 340 24731
rect 372 24699 412 24731
rect 444 24699 484 24731
rect 516 24699 556 24731
rect 588 24699 628 24731
rect 660 24699 700 24731
rect 732 24699 772 24731
rect 804 24699 844 24731
rect 876 24699 1000 24731
rect 0 24659 1000 24699
rect 0 24627 124 24659
rect 156 24627 196 24659
rect 228 24627 268 24659
rect 300 24627 340 24659
rect 372 24627 412 24659
rect 444 24627 484 24659
rect 516 24627 556 24659
rect 588 24627 628 24659
rect 660 24627 700 24659
rect 732 24627 772 24659
rect 804 24627 844 24659
rect 876 24627 1000 24659
rect 0 24587 1000 24627
rect 0 24555 124 24587
rect 156 24555 196 24587
rect 228 24555 268 24587
rect 300 24555 340 24587
rect 372 24555 412 24587
rect 444 24555 484 24587
rect 516 24555 556 24587
rect 588 24555 628 24587
rect 660 24555 700 24587
rect 732 24555 772 24587
rect 804 24555 844 24587
rect 876 24555 1000 24587
rect 0 24515 1000 24555
rect 0 24483 124 24515
rect 156 24483 196 24515
rect 228 24483 268 24515
rect 300 24483 340 24515
rect 372 24483 412 24515
rect 444 24483 484 24515
rect 516 24483 556 24515
rect 588 24483 628 24515
rect 660 24483 700 24515
rect 732 24483 772 24515
rect 804 24483 844 24515
rect 876 24483 1000 24515
rect 0 24443 1000 24483
rect 0 24411 124 24443
rect 156 24411 196 24443
rect 228 24411 268 24443
rect 300 24411 340 24443
rect 372 24411 412 24443
rect 444 24411 484 24443
rect 516 24411 556 24443
rect 588 24411 628 24443
rect 660 24411 700 24443
rect 732 24411 772 24443
rect 804 24411 844 24443
rect 876 24411 1000 24443
rect 0 24371 1000 24411
rect 0 24339 124 24371
rect 156 24339 196 24371
rect 228 24339 268 24371
rect 300 24339 340 24371
rect 372 24339 412 24371
rect 444 24339 484 24371
rect 516 24339 556 24371
rect 588 24339 628 24371
rect 660 24339 700 24371
rect 732 24339 772 24371
rect 804 24339 844 24371
rect 876 24339 1000 24371
rect 0 24299 1000 24339
rect 0 24267 124 24299
rect 156 24267 196 24299
rect 228 24267 268 24299
rect 300 24267 340 24299
rect 372 24267 412 24299
rect 444 24267 484 24299
rect 516 24267 556 24299
rect 588 24267 628 24299
rect 660 24267 700 24299
rect 732 24267 772 24299
rect 804 24267 844 24299
rect 876 24267 1000 24299
rect 0 24227 1000 24267
rect 0 24195 124 24227
rect 156 24195 196 24227
rect 228 24195 268 24227
rect 300 24195 340 24227
rect 372 24195 412 24227
rect 444 24195 484 24227
rect 516 24195 556 24227
rect 588 24195 628 24227
rect 660 24195 700 24227
rect 732 24195 772 24227
rect 804 24195 844 24227
rect 876 24195 1000 24227
rect 0 24155 1000 24195
rect 0 24123 124 24155
rect 156 24123 196 24155
rect 228 24123 268 24155
rect 300 24123 340 24155
rect 372 24123 412 24155
rect 444 24123 484 24155
rect 516 24123 556 24155
rect 588 24123 628 24155
rect 660 24123 700 24155
rect 732 24123 772 24155
rect 804 24123 844 24155
rect 876 24123 1000 24155
rect 0 24083 1000 24123
rect 0 24051 124 24083
rect 156 24051 196 24083
rect 228 24051 268 24083
rect 300 24051 340 24083
rect 372 24051 412 24083
rect 444 24051 484 24083
rect 516 24051 556 24083
rect 588 24051 628 24083
rect 660 24051 700 24083
rect 732 24051 772 24083
rect 804 24051 844 24083
rect 876 24051 1000 24083
rect 0 24011 1000 24051
rect 0 23979 124 24011
rect 156 23979 196 24011
rect 228 23979 268 24011
rect 300 23979 340 24011
rect 372 23979 412 24011
rect 444 23979 484 24011
rect 516 23979 556 24011
rect 588 23979 628 24011
rect 660 23979 700 24011
rect 732 23979 772 24011
rect 804 23979 844 24011
rect 876 23979 1000 24011
rect 0 23939 1000 23979
rect 0 23907 124 23939
rect 156 23907 196 23939
rect 228 23907 268 23939
rect 300 23907 340 23939
rect 372 23907 412 23939
rect 444 23907 484 23939
rect 516 23907 556 23939
rect 588 23907 628 23939
rect 660 23907 700 23939
rect 732 23907 772 23939
rect 804 23907 844 23939
rect 876 23907 1000 23939
rect 0 23867 1000 23907
rect 0 23835 124 23867
rect 156 23835 196 23867
rect 228 23835 268 23867
rect 300 23835 340 23867
rect 372 23835 412 23867
rect 444 23835 484 23867
rect 516 23835 556 23867
rect 588 23835 628 23867
rect 660 23835 700 23867
rect 732 23835 772 23867
rect 804 23835 844 23867
rect 876 23835 1000 23867
rect 0 23795 1000 23835
rect 0 23763 124 23795
rect 156 23763 196 23795
rect 228 23763 268 23795
rect 300 23763 340 23795
rect 372 23763 412 23795
rect 444 23763 484 23795
rect 516 23763 556 23795
rect 588 23763 628 23795
rect 660 23763 700 23795
rect 732 23763 772 23795
rect 804 23763 844 23795
rect 876 23763 1000 23795
rect 0 23723 1000 23763
rect 0 23691 124 23723
rect 156 23691 196 23723
rect 228 23691 268 23723
rect 300 23691 340 23723
rect 372 23691 412 23723
rect 444 23691 484 23723
rect 516 23691 556 23723
rect 588 23691 628 23723
rect 660 23691 700 23723
rect 732 23691 772 23723
rect 804 23691 844 23723
rect 876 23691 1000 23723
rect 0 23651 1000 23691
rect 0 23619 124 23651
rect 156 23619 196 23651
rect 228 23619 268 23651
rect 300 23619 340 23651
rect 372 23619 412 23651
rect 444 23619 484 23651
rect 516 23619 556 23651
rect 588 23619 628 23651
rect 660 23619 700 23651
rect 732 23619 772 23651
rect 804 23619 844 23651
rect 876 23619 1000 23651
rect 0 23579 1000 23619
rect 0 23547 124 23579
rect 156 23547 196 23579
rect 228 23547 268 23579
rect 300 23547 340 23579
rect 372 23547 412 23579
rect 444 23547 484 23579
rect 516 23547 556 23579
rect 588 23547 628 23579
rect 660 23547 700 23579
rect 732 23547 772 23579
rect 804 23547 844 23579
rect 876 23547 1000 23579
rect 0 23507 1000 23547
rect 0 23475 124 23507
rect 156 23475 196 23507
rect 228 23475 268 23507
rect 300 23475 340 23507
rect 372 23475 412 23507
rect 444 23475 484 23507
rect 516 23475 556 23507
rect 588 23475 628 23507
rect 660 23475 700 23507
rect 732 23475 772 23507
rect 804 23475 844 23507
rect 876 23475 1000 23507
rect 0 23435 1000 23475
rect 0 23403 124 23435
rect 156 23403 196 23435
rect 228 23403 268 23435
rect 300 23403 340 23435
rect 372 23403 412 23435
rect 444 23403 484 23435
rect 516 23403 556 23435
rect 588 23403 628 23435
rect 660 23403 700 23435
rect 732 23403 772 23435
rect 804 23403 844 23435
rect 876 23403 1000 23435
rect 0 23363 1000 23403
rect 0 23331 124 23363
rect 156 23331 196 23363
rect 228 23331 268 23363
rect 300 23331 340 23363
rect 372 23331 412 23363
rect 444 23331 484 23363
rect 516 23331 556 23363
rect 588 23331 628 23363
rect 660 23331 700 23363
rect 732 23331 772 23363
rect 804 23331 844 23363
rect 876 23331 1000 23363
rect 0 23291 1000 23331
rect 0 23259 124 23291
rect 156 23259 196 23291
rect 228 23259 268 23291
rect 300 23259 340 23291
rect 372 23259 412 23291
rect 444 23259 484 23291
rect 516 23259 556 23291
rect 588 23259 628 23291
rect 660 23259 700 23291
rect 732 23259 772 23291
rect 804 23259 844 23291
rect 876 23259 1000 23291
rect 0 23219 1000 23259
rect 0 23187 124 23219
rect 156 23187 196 23219
rect 228 23187 268 23219
rect 300 23187 340 23219
rect 372 23187 412 23219
rect 444 23187 484 23219
rect 516 23187 556 23219
rect 588 23187 628 23219
rect 660 23187 700 23219
rect 732 23187 772 23219
rect 804 23187 844 23219
rect 876 23187 1000 23219
rect 0 23124 1000 23187
rect 0 22874 1000 22924
rect 0 22842 124 22874
rect 156 22842 196 22874
rect 228 22842 268 22874
rect 300 22842 340 22874
rect 372 22842 412 22874
rect 444 22842 484 22874
rect 516 22842 556 22874
rect 588 22842 628 22874
rect 660 22842 700 22874
rect 732 22842 772 22874
rect 804 22842 844 22874
rect 876 22842 1000 22874
rect 0 22802 1000 22842
rect 0 22770 124 22802
rect 156 22770 196 22802
rect 228 22770 268 22802
rect 300 22770 340 22802
rect 372 22770 412 22802
rect 444 22770 484 22802
rect 516 22770 556 22802
rect 588 22770 628 22802
rect 660 22770 700 22802
rect 732 22770 772 22802
rect 804 22770 844 22802
rect 876 22770 1000 22802
rect 0 22730 1000 22770
rect 0 22698 124 22730
rect 156 22698 196 22730
rect 228 22698 268 22730
rect 300 22698 340 22730
rect 372 22698 412 22730
rect 444 22698 484 22730
rect 516 22698 556 22730
rect 588 22698 628 22730
rect 660 22698 700 22730
rect 732 22698 772 22730
rect 804 22698 844 22730
rect 876 22698 1000 22730
rect 0 22658 1000 22698
rect 0 22626 124 22658
rect 156 22626 196 22658
rect 228 22626 268 22658
rect 300 22626 340 22658
rect 372 22626 412 22658
rect 444 22626 484 22658
rect 516 22626 556 22658
rect 588 22626 628 22658
rect 660 22626 700 22658
rect 732 22626 772 22658
rect 804 22626 844 22658
rect 876 22626 1000 22658
rect 0 22586 1000 22626
rect 0 22554 124 22586
rect 156 22554 196 22586
rect 228 22554 268 22586
rect 300 22554 340 22586
rect 372 22554 412 22586
rect 444 22554 484 22586
rect 516 22554 556 22586
rect 588 22554 628 22586
rect 660 22554 700 22586
rect 732 22554 772 22586
rect 804 22554 844 22586
rect 876 22554 1000 22586
rect 0 22514 1000 22554
rect 0 22482 124 22514
rect 156 22482 196 22514
rect 228 22482 268 22514
rect 300 22482 340 22514
rect 372 22482 412 22514
rect 444 22482 484 22514
rect 516 22482 556 22514
rect 588 22482 628 22514
rect 660 22482 700 22514
rect 732 22482 772 22514
rect 804 22482 844 22514
rect 876 22482 1000 22514
rect 0 22442 1000 22482
rect 0 22410 124 22442
rect 156 22410 196 22442
rect 228 22410 268 22442
rect 300 22410 340 22442
rect 372 22410 412 22442
rect 444 22410 484 22442
rect 516 22410 556 22442
rect 588 22410 628 22442
rect 660 22410 700 22442
rect 732 22410 772 22442
rect 804 22410 844 22442
rect 876 22410 1000 22442
rect 0 22370 1000 22410
rect 0 22338 124 22370
rect 156 22338 196 22370
rect 228 22338 268 22370
rect 300 22338 340 22370
rect 372 22338 412 22370
rect 444 22338 484 22370
rect 516 22338 556 22370
rect 588 22338 628 22370
rect 660 22338 700 22370
rect 732 22338 772 22370
rect 804 22338 844 22370
rect 876 22338 1000 22370
rect 0 22298 1000 22338
rect 0 22266 124 22298
rect 156 22266 196 22298
rect 228 22266 268 22298
rect 300 22266 340 22298
rect 372 22266 412 22298
rect 444 22266 484 22298
rect 516 22266 556 22298
rect 588 22266 628 22298
rect 660 22266 700 22298
rect 732 22266 772 22298
rect 804 22266 844 22298
rect 876 22266 1000 22298
rect 0 22226 1000 22266
rect 0 22194 124 22226
rect 156 22194 196 22226
rect 228 22194 268 22226
rect 300 22194 340 22226
rect 372 22194 412 22226
rect 444 22194 484 22226
rect 516 22194 556 22226
rect 588 22194 628 22226
rect 660 22194 700 22226
rect 732 22194 772 22226
rect 804 22194 844 22226
rect 876 22194 1000 22226
rect 0 22154 1000 22194
rect 0 22122 124 22154
rect 156 22122 196 22154
rect 228 22122 268 22154
rect 300 22122 340 22154
rect 372 22122 412 22154
rect 444 22122 484 22154
rect 516 22122 556 22154
rect 588 22122 628 22154
rect 660 22122 700 22154
rect 732 22122 772 22154
rect 804 22122 844 22154
rect 876 22122 1000 22154
rect 0 22082 1000 22122
rect 0 22050 124 22082
rect 156 22050 196 22082
rect 228 22050 268 22082
rect 300 22050 340 22082
rect 372 22050 412 22082
rect 444 22050 484 22082
rect 516 22050 556 22082
rect 588 22050 628 22082
rect 660 22050 700 22082
rect 732 22050 772 22082
rect 804 22050 844 22082
rect 876 22050 1000 22082
rect 0 22010 1000 22050
rect 0 21978 124 22010
rect 156 21978 196 22010
rect 228 21978 268 22010
rect 300 21978 340 22010
rect 372 21978 412 22010
rect 444 21978 484 22010
rect 516 21978 556 22010
rect 588 21978 628 22010
rect 660 21978 700 22010
rect 732 21978 772 22010
rect 804 21978 844 22010
rect 876 21978 1000 22010
rect 0 21938 1000 21978
rect 0 21906 124 21938
rect 156 21906 196 21938
rect 228 21906 268 21938
rect 300 21906 340 21938
rect 372 21906 412 21938
rect 444 21906 484 21938
rect 516 21906 556 21938
rect 588 21906 628 21938
rect 660 21906 700 21938
rect 732 21906 772 21938
rect 804 21906 844 21938
rect 876 21906 1000 21938
rect 0 21866 1000 21906
rect 0 21834 124 21866
rect 156 21834 196 21866
rect 228 21834 268 21866
rect 300 21834 340 21866
rect 372 21834 412 21866
rect 444 21834 484 21866
rect 516 21834 556 21866
rect 588 21834 628 21866
rect 660 21834 700 21866
rect 732 21834 772 21866
rect 804 21834 844 21866
rect 876 21834 1000 21866
rect 0 21794 1000 21834
rect 0 21762 124 21794
rect 156 21762 196 21794
rect 228 21762 268 21794
rect 300 21762 340 21794
rect 372 21762 412 21794
rect 444 21762 484 21794
rect 516 21762 556 21794
rect 588 21762 628 21794
rect 660 21762 700 21794
rect 732 21762 772 21794
rect 804 21762 844 21794
rect 876 21762 1000 21794
rect 0 21722 1000 21762
rect 0 21690 124 21722
rect 156 21690 196 21722
rect 228 21690 268 21722
rect 300 21690 340 21722
rect 372 21690 412 21722
rect 444 21690 484 21722
rect 516 21690 556 21722
rect 588 21690 628 21722
rect 660 21690 700 21722
rect 732 21690 772 21722
rect 804 21690 844 21722
rect 876 21690 1000 21722
rect 0 21650 1000 21690
rect 0 21618 124 21650
rect 156 21618 196 21650
rect 228 21618 268 21650
rect 300 21618 340 21650
rect 372 21618 412 21650
rect 444 21618 484 21650
rect 516 21618 556 21650
rect 588 21618 628 21650
rect 660 21618 700 21650
rect 732 21618 772 21650
rect 804 21618 844 21650
rect 876 21618 1000 21650
rect 0 21578 1000 21618
rect 0 21546 124 21578
rect 156 21546 196 21578
rect 228 21546 268 21578
rect 300 21546 340 21578
rect 372 21546 412 21578
rect 444 21546 484 21578
rect 516 21546 556 21578
rect 588 21546 628 21578
rect 660 21546 700 21578
rect 732 21546 772 21578
rect 804 21546 844 21578
rect 876 21546 1000 21578
rect 0 21506 1000 21546
rect 0 21474 124 21506
rect 156 21474 196 21506
rect 228 21474 268 21506
rect 300 21474 340 21506
rect 372 21474 412 21506
rect 444 21474 484 21506
rect 516 21474 556 21506
rect 588 21474 628 21506
rect 660 21474 700 21506
rect 732 21474 772 21506
rect 804 21474 844 21506
rect 876 21474 1000 21506
rect 0 21434 1000 21474
rect 0 21402 124 21434
rect 156 21402 196 21434
rect 228 21402 268 21434
rect 300 21402 340 21434
rect 372 21402 412 21434
rect 444 21402 484 21434
rect 516 21402 556 21434
rect 588 21402 628 21434
rect 660 21402 700 21434
rect 732 21402 772 21434
rect 804 21402 844 21434
rect 876 21402 1000 21434
rect 0 21362 1000 21402
rect 0 21330 124 21362
rect 156 21330 196 21362
rect 228 21330 268 21362
rect 300 21330 340 21362
rect 372 21330 412 21362
rect 444 21330 484 21362
rect 516 21330 556 21362
rect 588 21330 628 21362
rect 660 21330 700 21362
rect 732 21330 772 21362
rect 804 21330 844 21362
rect 876 21330 1000 21362
rect 0 21290 1000 21330
rect 0 21258 124 21290
rect 156 21258 196 21290
rect 228 21258 268 21290
rect 300 21258 340 21290
rect 372 21258 412 21290
rect 444 21258 484 21290
rect 516 21258 556 21290
rect 588 21258 628 21290
rect 660 21258 700 21290
rect 732 21258 772 21290
rect 804 21258 844 21290
rect 876 21258 1000 21290
rect 0 21218 1000 21258
rect 0 21186 124 21218
rect 156 21186 196 21218
rect 228 21186 268 21218
rect 300 21186 340 21218
rect 372 21186 412 21218
rect 444 21186 484 21218
rect 516 21186 556 21218
rect 588 21186 628 21218
rect 660 21186 700 21218
rect 732 21186 772 21218
rect 804 21186 844 21218
rect 876 21186 1000 21218
rect 0 21146 1000 21186
rect 0 21114 124 21146
rect 156 21114 196 21146
rect 228 21114 268 21146
rect 300 21114 340 21146
rect 372 21114 412 21146
rect 444 21114 484 21146
rect 516 21114 556 21146
rect 588 21114 628 21146
rect 660 21114 700 21146
rect 732 21114 772 21146
rect 804 21114 844 21146
rect 876 21114 1000 21146
rect 0 21074 1000 21114
rect 0 21042 124 21074
rect 156 21042 196 21074
rect 228 21042 268 21074
rect 300 21042 340 21074
rect 372 21042 412 21074
rect 444 21042 484 21074
rect 516 21042 556 21074
rect 588 21042 628 21074
rect 660 21042 700 21074
rect 732 21042 772 21074
rect 804 21042 844 21074
rect 876 21042 1000 21074
rect 0 21002 1000 21042
rect 0 20970 124 21002
rect 156 20970 196 21002
rect 228 20970 268 21002
rect 300 20970 340 21002
rect 372 20970 412 21002
rect 444 20970 484 21002
rect 516 20970 556 21002
rect 588 20970 628 21002
rect 660 20970 700 21002
rect 732 20970 772 21002
rect 804 20970 844 21002
rect 876 20970 1000 21002
rect 0 20930 1000 20970
rect 0 20898 124 20930
rect 156 20898 196 20930
rect 228 20898 268 20930
rect 300 20898 340 20930
rect 372 20898 412 20930
rect 444 20898 484 20930
rect 516 20898 556 20930
rect 588 20898 628 20930
rect 660 20898 700 20930
rect 732 20898 772 20930
rect 804 20898 844 20930
rect 876 20898 1000 20930
rect 0 20858 1000 20898
rect 0 20826 124 20858
rect 156 20826 196 20858
rect 228 20826 268 20858
rect 300 20826 340 20858
rect 372 20826 412 20858
rect 444 20826 484 20858
rect 516 20826 556 20858
rect 588 20826 628 20858
rect 660 20826 700 20858
rect 732 20826 772 20858
rect 804 20826 844 20858
rect 876 20826 1000 20858
rect 0 20786 1000 20826
rect 0 20754 124 20786
rect 156 20754 196 20786
rect 228 20754 268 20786
rect 300 20754 340 20786
rect 372 20754 412 20786
rect 444 20754 484 20786
rect 516 20754 556 20786
rect 588 20754 628 20786
rect 660 20754 700 20786
rect 732 20754 772 20786
rect 804 20754 844 20786
rect 876 20754 1000 20786
rect 0 20714 1000 20754
rect 0 20682 124 20714
rect 156 20682 196 20714
rect 228 20682 268 20714
rect 300 20682 340 20714
rect 372 20682 412 20714
rect 444 20682 484 20714
rect 516 20682 556 20714
rect 588 20682 628 20714
rect 660 20682 700 20714
rect 732 20682 772 20714
rect 804 20682 844 20714
rect 876 20682 1000 20714
rect 0 20642 1000 20682
rect 0 20610 124 20642
rect 156 20610 196 20642
rect 228 20610 268 20642
rect 300 20610 340 20642
rect 372 20610 412 20642
rect 444 20610 484 20642
rect 516 20610 556 20642
rect 588 20610 628 20642
rect 660 20610 700 20642
rect 732 20610 772 20642
rect 804 20610 844 20642
rect 876 20610 1000 20642
rect 0 20570 1000 20610
rect 0 20538 124 20570
rect 156 20538 196 20570
rect 228 20538 268 20570
rect 300 20538 340 20570
rect 372 20538 412 20570
rect 444 20538 484 20570
rect 516 20538 556 20570
rect 588 20538 628 20570
rect 660 20538 700 20570
rect 732 20538 772 20570
rect 804 20538 844 20570
rect 876 20538 1000 20570
rect 0 20498 1000 20538
rect 0 20466 124 20498
rect 156 20466 196 20498
rect 228 20466 268 20498
rect 300 20466 340 20498
rect 372 20466 412 20498
rect 444 20466 484 20498
rect 516 20466 556 20498
rect 588 20466 628 20498
rect 660 20466 700 20498
rect 732 20466 772 20498
rect 804 20466 844 20498
rect 876 20466 1000 20498
rect 0 20426 1000 20466
rect 0 20394 124 20426
rect 156 20394 196 20426
rect 228 20394 268 20426
rect 300 20394 340 20426
rect 372 20394 412 20426
rect 444 20394 484 20426
rect 516 20394 556 20426
rect 588 20394 628 20426
rect 660 20394 700 20426
rect 732 20394 772 20426
rect 804 20394 844 20426
rect 876 20394 1000 20426
rect 0 20354 1000 20394
rect 0 20322 124 20354
rect 156 20322 196 20354
rect 228 20322 268 20354
rect 300 20322 340 20354
rect 372 20322 412 20354
rect 444 20322 484 20354
rect 516 20322 556 20354
rect 588 20322 628 20354
rect 660 20322 700 20354
rect 732 20322 772 20354
rect 804 20322 844 20354
rect 876 20322 1000 20354
rect 0 20282 1000 20322
rect 0 20250 124 20282
rect 156 20250 196 20282
rect 228 20250 268 20282
rect 300 20250 340 20282
rect 372 20250 412 20282
rect 444 20250 484 20282
rect 516 20250 556 20282
rect 588 20250 628 20282
rect 660 20250 700 20282
rect 732 20250 772 20282
rect 804 20250 844 20282
rect 876 20250 1000 20282
rect 0 20210 1000 20250
rect 0 20178 124 20210
rect 156 20178 196 20210
rect 228 20178 268 20210
rect 300 20178 340 20210
rect 372 20178 412 20210
rect 444 20178 484 20210
rect 516 20178 556 20210
rect 588 20178 628 20210
rect 660 20178 700 20210
rect 732 20178 772 20210
rect 804 20178 844 20210
rect 876 20178 1000 20210
rect 0 20138 1000 20178
rect 0 20106 124 20138
rect 156 20106 196 20138
rect 228 20106 268 20138
rect 300 20106 340 20138
rect 372 20106 412 20138
rect 444 20106 484 20138
rect 516 20106 556 20138
rect 588 20106 628 20138
rect 660 20106 700 20138
rect 732 20106 772 20138
rect 804 20106 844 20138
rect 876 20106 1000 20138
rect 0 20066 1000 20106
rect 0 20034 124 20066
rect 156 20034 196 20066
rect 228 20034 268 20066
rect 300 20034 340 20066
rect 372 20034 412 20066
rect 444 20034 484 20066
rect 516 20034 556 20066
rect 588 20034 628 20066
rect 660 20034 700 20066
rect 732 20034 772 20066
rect 804 20034 844 20066
rect 876 20034 1000 20066
rect 0 19994 1000 20034
rect 0 19962 124 19994
rect 156 19962 196 19994
rect 228 19962 268 19994
rect 300 19962 340 19994
rect 372 19962 412 19994
rect 444 19962 484 19994
rect 516 19962 556 19994
rect 588 19962 628 19994
rect 660 19962 700 19994
rect 732 19962 772 19994
rect 804 19962 844 19994
rect 876 19962 1000 19994
rect 0 19922 1000 19962
rect 0 19890 124 19922
rect 156 19890 196 19922
rect 228 19890 268 19922
rect 300 19890 340 19922
rect 372 19890 412 19922
rect 444 19890 484 19922
rect 516 19890 556 19922
rect 588 19890 628 19922
rect 660 19890 700 19922
rect 732 19890 772 19922
rect 804 19890 844 19922
rect 876 19890 1000 19922
rect 0 19850 1000 19890
rect 0 19818 124 19850
rect 156 19818 196 19850
rect 228 19818 268 19850
rect 300 19818 340 19850
rect 372 19818 412 19850
rect 444 19818 484 19850
rect 516 19818 556 19850
rect 588 19818 628 19850
rect 660 19818 700 19850
rect 732 19818 772 19850
rect 804 19818 844 19850
rect 876 19818 1000 19850
rect 0 19778 1000 19818
rect 0 19746 124 19778
rect 156 19746 196 19778
rect 228 19746 268 19778
rect 300 19746 340 19778
rect 372 19746 412 19778
rect 444 19746 484 19778
rect 516 19746 556 19778
rect 588 19746 628 19778
rect 660 19746 700 19778
rect 732 19746 772 19778
rect 804 19746 844 19778
rect 876 19746 1000 19778
rect 0 19706 1000 19746
rect 0 19674 124 19706
rect 156 19674 196 19706
rect 228 19674 268 19706
rect 300 19674 340 19706
rect 372 19674 412 19706
rect 444 19674 484 19706
rect 516 19674 556 19706
rect 588 19674 628 19706
rect 660 19674 700 19706
rect 732 19674 772 19706
rect 804 19674 844 19706
rect 876 19674 1000 19706
rect 0 19634 1000 19674
rect 0 19602 124 19634
rect 156 19602 196 19634
rect 228 19602 268 19634
rect 300 19602 340 19634
rect 372 19602 412 19634
rect 444 19602 484 19634
rect 516 19602 556 19634
rect 588 19602 628 19634
rect 660 19602 700 19634
rect 732 19602 772 19634
rect 804 19602 844 19634
rect 876 19602 1000 19634
rect 0 19562 1000 19602
rect 0 19530 124 19562
rect 156 19530 196 19562
rect 228 19530 268 19562
rect 300 19530 340 19562
rect 372 19530 412 19562
rect 444 19530 484 19562
rect 516 19530 556 19562
rect 588 19530 628 19562
rect 660 19530 700 19562
rect 732 19530 772 19562
rect 804 19530 844 19562
rect 876 19530 1000 19562
rect 0 19490 1000 19530
rect 0 19458 124 19490
rect 156 19458 196 19490
rect 228 19458 268 19490
rect 300 19458 340 19490
rect 372 19458 412 19490
rect 444 19458 484 19490
rect 516 19458 556 19490
rect 588 19458 628 19490
rect 660 19458 700 19490
rect 732 19458 772 19490
rect 804 19458 844 19490
rect 876 19458 1000 19490
rect 0 19418 1000 19458
rect 0 19386 124 19418
rect 156 19386 196 19418
rect 228 19386 268 19418
rect 300 19386 340 19418
rect 372 19386 412 19418
rect 444 19386 484 19418
rect 516 19386 556 19418
rect 588 19386 628 19418
rect 660 19386 700 19418
rect 732 19386 772 19418
rect 804 19386 844 19418
rect 876 19386 1000 19418
rect 0 19346 1000 19386
rect 0 19314 124 19346
rect 156 19314 196 19346
rect 228 19314 268 19346
rect 300 19314 340 19346
rect 372 19314 412 19346
rect 444 19314 484 19346
rect 516 19314 556 19346
rect 588 19314 628 19346
rect 660 19314 700 19346
rect 732 19314 772 19346
rect 804 19314 844 19346
rect 876 19314 1000 19346
rect 0 19274 1000 19314
rect 0 19242 124 19274
rect 156 19242 196 19274
rect 228 19242 268 19274
rect 300 19242 340 19274
rect 372 19242 412 19274
rect 444 19242 484 19274
rect 516 19242 556 19274
rect 588 19242 628 19274
rect 660 19242 700 19274
rect 732 19242 772 19274
rect 804 19242 844 19274
rect 876 19242 1000 19274
rect 0 19202 1000 19242
rect 0 19170 124 19202
rect 156 19170 196 19202
rect 228 19170 268 19202
rect 300 19170 340 19202
rect 372 19170 412 19202
rect 444 19170 484 19202
rect 516 19170 556 19202
rect 588 19170 628 19202
rect 660 19170 700 19202
rect 732 19170 772 19202
rect 804 19170 844 19202
rect 876 19170 1000 19202
rect 0 19130 1000 19170
rect 0 19098 124 19130
rect 156 19098 196 19130
rect 228 19098 268 19130
rect 300 19098 340 19130
rect 372 19098 412 19130
rect 444 19098 484 19130
rect 516 19098 556 19130
rect 588 19098 628 19130
rect 660 19098 700 19130
rect 732 19098 772 19130
rect 804 19098 844 19130
rect 876 19098 1000 19130
rect 0 19058 1000 19098
rect 0 19026 124 19058
rect 156 19026 196 19058
rect 228 19026 268 19058
rect 300 19026 340 19058
rect 372 19026 412 19058
rect 444 19026 484 19058
rect 516 19026 556 19058
rect 588 19026 628 19058
rect 660 19026 700 19058
rect 732 19026 772 19058
rect 804 19026 844 19058
rect 876 19026 1000 19058
rect 0 18986 1000 19026
rect 0 18954 124 18986
rect 156 18954 196 18986
rect 228 18954 268 18986
rect 300 18954 340 18986
rect 372 18954 412 18986
rect 444 18954 484 18986
rect 516 18954 556 18986
rect 588 18954 628 18986
rect 660 18954 700 18986
rect 732 18954 772 18986
rect 804 18954 844 18986
rect 876 18954 1000 18986
rect 0 18914 1000 18954
rect 0 18882 124 18914
rect 156 18882 196 18914
rect 228 18882 268 18914
rect 300 18882 340 18914
rect 372 18882 412 18914
rect 444 18882 484 18914
rect 516 18882 556 18914
rect 588 18882 628 18914
rect 660 18882 700 18914
rect 732 18882 772 18914
rect 804 18882 844 18914
rect 876 18882 1000 18914
rect 0 18842 1000 18882
rect 0 18810 124 18842
rect 156 18810 196 18842
rect 228 18810 268 18842
rect 300 18810 340 18842
rect 372 18810 412 18842
rect 444 18810 484 18842
rect 516 18810 556 18842
rect 588 18810 628 18842
rect 660 18810 700 18842
rect 732 18810 772 18842
rect 804 18810 844 18842
rect 876 18810 1000 18842
rect 0 18770 1000 18810
rect 0 18738 124 18770
rect 156 18738 196 18770
rect 228 18738 268 18770
rect 300 18738 340 18770
rect 372 18738 412 18770
rect 444 18738 484 18770
rect 516 18738 556 18770
rect 588 18738 628 18770
rect 660 18738 700 18770
rect 732 18738 772 18770
rect 804 18738 844 18770
rect 876 18738 1000 18770
rect 0 18698 1000 18738
rect 0 18666 124 18698
rect 156 18666 196 18698
rect 228 18666 268 18698
rect 300 18666 340 18698
rect 372 18666 412 18698
rect 444 18666 484 18698
rect 516 18666 556 18698
rect 588 18666 628 18698
rect 660 18666 700 18698
rect 732 18666 772 18698
rect 804 18666 844 18698
rect 876 18666 1000 18698
rect 0 18626 1000 18666
rect 0 18594 124 18626
rect 156 18594 196 18626
rect 228 18594 268 18626
rect 300 18594 340 18626
rect 372 18594 412 18626
rect 444 18594 484 18626
rect 516 18594 556 18626
rect 588 18594 628 18626
rect 660 18594 700 18626
rect 732 18594 772 18626
rect 804 18594 844 18626
rect 876 18594 1000 18626
rect 0 18554 1000 18594
rect 0 18522 124 18554
rect 156 18522 196 18554
rect 228 18522 268 18554
rect 300 18522 340 18554
rect 372 18522 412 18554
rect 444 18522 484 18554
rect 516 18522 556 18554
rect 588 18522 628 18554
rect 660 18522 700 18554
rect 732 18522 772 18554
rect 804 18522 844 18554
rect 876 18522 1000 18554
rect 0 18482 1000 18522
rect 0 18450 124 18482
rect 156 18450 196 18482
rect 228 18450 268 18482
rect 300 18450 340 18482
rect 372 18450 412 18482
rect 444 18450 484 18482
rect 516 18450 556 18482
rect 588 18450 628 18482
rect 660 18450 700 18482
rect 732 18450 772 18482
rect 804 18450 844 18482
rect 876 18450 1000 18482
rect 0 18410 1000 18450
rect 0 18378 124 18410
rect 156 18378 196 18410
rect 228 18378 268 18410
rect 300 18378 340 18410
rect 372 18378 412 18410
rect 444 18378 484 18410
rect 516 18378 556 18410
rect 588 18378 628 18410
rect 660 18378 700 18410
rect 732 18378 772 18410
rect 804 18378 844 18410
rect 876 18378 1000 18410
rect 0 18338 1000 18378
rect 0 18306 124 18338
rect 156 18306 196 18338
rect 228 18306 268 18338
rect 300 18306 340 18338
rect 372 18306 412 18338
rect 444 18306 484 18338
rect 516 18306 556 18338
rect 588 18306 628 18338
rect 660 18306 700 18338
rect 732 18306 772 18338
rect 804 18306 844 18338
rect 876 18306 1000 18338
rect 0 18266 1000 18306
rect 0 18234 124 18266
rect 156 18234 196 18266
rect 228 18234 268 18266
rect 300 18234 340 18266
rect 372 18234 412 18266
rect 444 18234 484 18266
rect 516 18234 556 18266
rect 588 18234 628 18266
rect 660 18234 700 18266
rect 732 18234 772 18266
rect 804 18234 844 18266
rect 876 18234 1000 18266
rect 0 18194 1000 18234
rect 0 18162 124 18194
rect 156 18162 196 18194
rect 228 18162 268 18194
rect 300 18162 340 18194
rect 372 18162 412 18194
rect 444 18162 484 18194
rect 516 18162 556 18194
rect 588 18162 628 18194
rect 660 18162 700 18194
rect 732 18162 772 18194
rect 804 18162 844 18194
rect 876 18162 1000 18194
rect 0 18112 1000 18162
rect 0 17848 1000 17912
rect 0 17816 124 17848
rect 156 17816 196 17848
rect 228 17816 268 17848
rect 300 17816 340 17848
rect 372 17816 412 17848
rect 444 17816 484 17848
rect 516 17816 556 17848
rect 588 17816 628 17848
rect 660 17816 700 17848
rect 732 17816 772 17848
rect 804 17816 844 17848
rect 876 17816 1000 17848
rect 0 17776 1000 17816
rect 0 17744 124 17776
rect 156 17744 196 17776
rect 228 17744 268 17776
rect 300 17744 340 17776
rect 372 17744 412 17776
rect 444 17744 484 17776
rect 516 17744 556 17776
rect 588 17744 628 17776
rect 660 17744 700 17776
rect 732 17744 772 17776
rect 804 17744 844 17776
rect 876 17744 1000 17776
rect 0 17704 1000 17744
rect 0 17672 124 17704
rect 156 17672 196 17704
rect 228 17672 268 17704
rect 300 17672 340 17704
rect 372 17672 412 17704
rect 444 17672 484 17704
rect 516 17672 556 17704
rect 588 17672 628 17704
rect 660 17672 700 17704
rect 732 17672 772 17704
rect 804 17672 844 17704
rect 876 17672 1000 17704
rect 0 17632 1000 17672
rect 0 17600 124 17632
rect 156 17600 196 17632
rect 228 17600 268 17632
rect 300 17600 340 17632
rect 372 17600 412 17632
rect 444 17600 484 17632
rect 516 17600 556 17632
rect 588 17600 628 17632
rect 660 17600 700 17632
rect 732 17600 772 17632
rect 804 17600 844 17632
rect 876 17600 1000 17632
rect 0 17560 1000 17600
rect 0 17528 124 17560
rect 156 17528 196 17560
rect 228 17528 268 17560
rect 300 17528 340 17560
rect 372 17528 412 17560
rect 444 17528 484 17560
rect 516 17528 556 17560
rect 588 17528 628 17560
rect 660 17528 700 17560
rect 732 17528 772 17560
rect 804 17528 844 17560
rect 876 17528 1000 17560
rect 0 17488 1000 17528
rect 0 17456 124 17488
rect 156 17456 196 17488
rect 228 17456 268 17488
rect 300 17456 340 17488
rect 372 17456 412 17488
rect 444 17456 484 17488
rect 516 17456 556 17488
rect 588 17456 628 17488
rect 660 17456 700 17488
rect 732 17456 772 17488
rect 804 17456 844 17488
rect 876 17456 1000 17488
rect 0 17416 1000 17456
rect 0 17384 124 17416
rect 156 17384 196 17416
rect 228 17384 268 17416
rect 300 17384 340 17416
rect 372 17384 412 17416
rect 444 17384 484 17416
rect 516 17384 556 17416
rect 588 17384 628 17416
rect 660 17384 700 17416
rect 732 17384 772 17416
rect 804 17384 844 17416
rect 876 17384 1000 17416
rect 0 17344 1000 17384
rect 0 17312 124 17344
rect 156 17312 196 17344
rect 228 17312 268 17344
rect 300 17312 340 17344
rect 372 17312 412 17344
rect 444 17312 484 17344
rect 516 17312 556 17344
rect 588 17312 628 17344
rect 660 17312 700 17344
rect 732 17312 772 17344
rect 804 17312 844 17344
rect 876 17312 1000 17344
rect 0 17272 1000 17312
rect 0 17240 124 17272
rect 156 17240 196 17272
rect 228 17240 268 17272
rect 300 17240 340 17272
rect 372 17240 412 17272
rect 444 17240 484 17272
rect 516 17240 556 17272
rect 588 17240 628 17272
rect 660 17240 700 17272
rect 732 17240 772 17272
rect 804 17240 844 17272
rect 876 17240 1000 17272
rect 0 17200 1000 17240
rect 0 17168 124 17200
rect 156 17168 196 17200
rect 228 17168 268 17200
rect 300 17168 340 17200
rect 372 17168 412 17200
rect 444 17168 484 17200
rect 516 17168 556 17200
rect 588 17168 628 17200
rect 660 17168 700 17200
rect 732 17168 772 17200
rect 804 17168 844 17200
rect 876 17168 1000 17200
rect 0 17128 1000 17168
rect 0 17096 124 17128
rect 156 17096 196 17128
rect 228 17096 268 17128
rect 300 17096 340 17128
rect 372 17096 412 17128
rect 444 17096 484 17128
rect 516 17096 556 17128
rect 588 17096 628 17128
rect 660 17096 700 17128
rect 732 17096 772 17128
rect 804 17096 844 17128
rect 876 17096 1000 17128
rect 0 17056 1000 17096
rect 0 17024 124 17056
rect 156 17024 196 17056
rect 228 17024 268 17056
rect 300 17024 340 17056
rect 372 17024 412 17056
rect 444 17024 484 17056
rect 516 17024 556 17056
rect 588 17024 628 17056
rect 660 17024 700 17056
rect 732 17024 772 17056
rect 804 17024 844 17056
rect 876 17024 1000 17056
rect 0 16984 1000 17024
rect 0 16952 124 16984
rect 156 16952 196 16984
rect 228 16952 268 16984
rect 300 16952 340 16984
rect 372 16952 412 16984
rect 444 16952 484 16984
rect 516 16952 556 16984
rect 588 16952 628 16984
rect 660 16952 700 16984
rect 732 16952 772 16984
rect 804 16952 844 16984
rect 876 16952 1000 16984
rect 0 16912 1000 16952
rect 0 16880 124 16912
rect 156 16880 196 16912
rect 228 16880 268 16912
rect 300 16880 340 16912
rect 372 16880 412 16912
rect 444 16880 484 16912
rect 516 16880 556 16912
rect 588 16880 628 16912
rect 660 16880 700 16912
rect 732 16880 772 16912
rect 804 16880 844 16912
rect 876 16880 1000 16912
rect 0 16840 1000 16880
rect 0 16808 124 16840
rect 156 16808 196 16840
rect 228 16808 268 16840
rect 300 16808 340 16840
rect 372 16808 412 16840
rect 444 16808 484 16840
rect 516 16808 556 16840
rect 588 16808 628 16840
rect 660 16808 700 16840
rect 732 16808 772 16840
rect 804 16808 844 16840
rect 876 16808 1000 16840
rect 0 16768 1000 16808
rect 0 16736 124 16768
rect 156 16736 196 16768
rect 228 16736 268 16768
rect 300 16736 340 16768
rect 372 16736 412 16768
rect 444 16736 484 16768
rect 516 16736 556 16768
rect 588 16736 628 16768
rect 660 16736 700 16768
rect 732 16736 772 16768
rect 804 16736 844 16768
rect 876 16736 1000 16768
rect 0 16696 1000 16736
rect 0 16664 124 16696
rect 156 16664 196 16696
rect 228 16664 268 16696
rect 300 16664 340 16696
rect 372 16664 412 16696
rect 444 16664 484 16696
rect 516 16664 556 16696
rect 588 16664 628 16696
rect 660 16664 700 16696
rect 732 16664 772 16696
rect 804 16664 844 16696
rect 876 16664 1000 16696
rect 0 16624 1000 16664
rect 0 16592 124 16624
rect 156 16592 196 16624
rect 228 16592 268 16624
rect 300 16592 340 16624
rect 372 16592 412 16624
rect 444 16592 484 16624
rect 516 16592 556 16624
rect 588 16592 628 16624
rect 660 16592 700 16624
rect 732 16592 772 16624
rect 804 16592 844 16624
rect 876 16592 1000 16624
rect 0 16552 1000 16592
rect 0 16520 124 16552
rect 156 16520 196 16552
rect 228 16520 268 16552
rect 300 16520 340 16552
rect 372 16520 412 16552
rect 444 16520 484 16552
rect 516 16520 556 16552
rect 588 16520 628 16552
rect 660 16520 700 16552
rect 732 16520 772 16552
rect 804 16520 844 16552
rect 876 16520 1000 16552
rect 0 16480 1000 16520
rect 0 16448 124 16480
rect 156 16448 196 16480
rect 228 16448 268 16480
rect 300 16448 340 16480
rect 372 16448 412 16480
rect 444 16448 484 16480
rect 516 16448 556 16480
rect 588 16448 628 16480
rect 660 16448 700 16480
rect 732 16448 772 16480
rect 804 16448 844 16480
rect 876 16448 1000 16480
rect 0 16408 1000 16448
rect 0 16376 124 16408
rect 156 16376 196 16408
rect 228 16376 268 16408
rect 300 16376 340 16408
rect 372 16376 412 16408
rect 444 16376 484 16408
rect 516 16376 556 16408
rect 588 16376 628 16408
rect 660 16376 700 16408
rect 732 16376 772 16408
rect 804 16376 844 16408
rect 876 16376 1000 16408
rect 0 16336 1000 16376
rect 0 16304 124 16336
rect 156 16304 196 16336
rect 228 16304 268 16336
rect 300 16304 340 16336
rect 372 16304 412 16336
rect 444 16304 484 16336
rect 516 16304 556 16336
rect 588 16304 628 16336
rect 660 16304 700 16336
rect 732 16304 772 16336
rect 804 16304 844 16336
rect 876 16304 1000 16336
rect 0 16264 1000 16304
rect 0 16232 124 16264
rect 156 16232 196 16264
rect 228 16232 268 16264
rect 300 16232 340 16264
rect 372 16232 412 16264
rect 444 16232 484 16264
rect 516 16232 556 16264
rect 588 16232 628 16264
rect 660 16232 700 16264
rect 732 16232 772 16264
rect 804 16232 844 16264
rect 876 16232 1000 16264
rect 0 16192 1000 16232
rect 0 16160 124 16192
rect 156 16160 196 16192
rect 228 16160 268 16192
rect 300 16160 340 16192
rect 372 16160 412 16192
rect 444 16160 484 16192
rect 516 16160 556 16192
rect 588 16160 628 16192
rect 660 16160 700 16192
rect 732 16160 772 16192
rect 804 16160 844 16192
rect 876 16160 1000 16192
rect 0 16120 1000 16160
rect 0 16088 124 16120
rect 156 16088 196 16120
rect 228 16088 268 16120
rect 300 16088 340 16120
rect 372 16088 412 16120
rect 444 16088 484 16120
rect 516 16088 556 16120
rect 588 16088 628 16120
rect 660 16088 700 16120
rect 732 16088 772 16120
rect 804 16088 844 16120
rect 876 16088 1000 16120
rect 0 16048 1000 16088
rect 0 16016 124 16048
rect 156 16016 196 16048
rect 228 16016 268 16048
rect 300 16016 340 16048
rect 372 16016 412 16048
rect 444 16016 484 16048
rect 516 16016 556 16048
rect 588 16016 628 16048
rect 660 16016 700 16048
rect 732 16016 772 16048
rect 804 16016 844 16048
rect 876 16016 1000 16048
rect 0 15976 1000 16016
rect 0 15944 124 15976
rect 156 15944 196 15976
rect 228 15944 268 15976
rect 300 15944 340 15976
rect 372 15944 412 15976
rect 444 15944 484 15976
rect 516 15944 556 15976
rect 588 15944 628 15976
rect 660 15944 700 15976
rect 732 15944 772 15976
rect 804 15944 844 15976
rect 876 15944 1000 15976
rect 0 15904 1000 15944
rect 0 15872 124 15904
rect 156 15872 196 15904
rect 228 15872 268 15904
rect 300 15872 340 15904
rect 372 15872 412 15904
rect 444 15872 484 15904
rect 516 15872 556 15904
rect 588 15872 628 15904
rect 660 15872 700 15904
rect 732 15872 772 15904
rect 804 15872 844 15904
rect 876 15872 1000 15904
rect 0 15832 1000 15872
rect 0 15800 124 15832
rect 156 15800 196 15832
rect 228 15800 268 15832
rect 300 15800 340 15832
rect 372 15800 412 15832
rect 444 15800 484 15832
rect 516 15800 556 15832
rect 588 15800 628 15832
rect 660 15800 700 15832
rect 732 15800 772 15832
rect 804 15800 844 15832
rect 876 15800 1000 15832
rect 0 15760 1000 15800
rect 0 15728 124 15760
rect 156 15728 196 15760
rect 228 15728 268 15760
rect 300 15728 340 15760
rect 372 15728 412 15760
rect 444 15728 484 15760
rect 516 15728 556 15760
rect 588 15728 628 15760
rect 660 15728 700 15760
rect 732 15728 772 15760
rect 804 15728 844 15760
rect 876 15728 1000 15760
rect 0 15688 1000 15728
rect 0 15656 124 15688
rect 156 15656 196 15688
rect 228 15656 268 15688
rect 300 15656 340 15688
rect 372 15656 412 15688
rect 444 15656 484 15688
rect 516 15656 556 15688
rect 588 15656 628 15688
rect 660 15656 700 15688
rect 732 15656 772 15688
rect 804 15656 844 15688
rect 876 15656 1000 15688
rect 0 15616 1000 15656
rect 0 15584 124 15616
rect 156 15584 196 15616
rect 228 15584 268 15616
rect 300 15584 340 15616
rect 372 15584 412 15616
rect 444 15584 484 15616
rect 516 15584 556 15616
rect 588 15584 628 15616
rect 660 15584 700 15616
rect 732 15584 772 15616
rect 804 15584 844 15616
rect 876 15584 1000 15616
rect 0 15544 1000 15584
rect 0 15512 124 15544
rect 156 15512 196 15544
rect 228 15512 268 15544
rect 300 15512 340 15544
rect 372 15512 412 15544
rect 444 15512 484 15544
rect 516 15512 556 15544
rect 588 15512 628 15544
rect 660 15512 700 15544
rect 732 15512 772 15544
rect 804 15512 844 15544
rect 876 15512 1000 15544
rect 0 15472 1000 15512
rect 0 15440 124 15472
rect 156 15440 196 15472
rect 228 15440 268 15472
rect 300 15440 340 15472
rect 372 15440 412 15472
rect 444 15440 484 15472
rect 516 15440 556 15472
rect 588 15440 628 15472
rect 660 15440 700 15472
rect 732 15440 772 15472
rect 804 15440 844 15472
rect 876 15440 1000 15472
rect 0 15400 1000 15440
rect 0 15368 124 15400
rect 156 15368 196 15400
rect 228 15368 268 15400
rect 300 15368 340 15400
rect 372 15368 412 15400
rect 444 15368 484 15400
rect 516 15368 556 15400
rect 588 15368 628 15400
rect 660 15368 700 15400
rect 732 15368 772 15400
rect 804 15368 844 15400
rect 876 15368 1000 15400
rect 0 15328 1000 15368
rect 0 15296 124 15328
rect 156 15296 196 15328
rect 228 15296 268 15328
rect 300 15296 340 15328
rect 372 15296 412 15328
rect 444 15296 484 15328
rect 516 15296 556 15328
rect 588 15296 628 15328
rect 660 15296 700 15328
rect 732 15296 772 15328
rect 804 15296 844 15328
rect 876 15296 1000 15328
rect 0 15256 1000 15296
rect 0 15224 124 15256
rect 156 15224 196 15256
rect 228 15224 268 15256
rect 300 15224 340 15256
rect 372 15224 412 15256
rect 444 15224 484 15256
rect 516 15224 556 15256
rect 588 15224 628 15256
rect 660 15224 700 15256
rect 732 15224 772 15256
rect 804 15224 844 15256
rect 876 15224 1000 15256
rect 0 15184 1000 15224
rect 0 15152 124 15184
rect 156 15152 196 15184
rect 228 15152 268 15184
rect 300 15152 340 15184
rect 372 15152 412 15184
rect 444 15152 484 15184
rect 516 15152 556 15184
rect 588 15152 628 15184
rect 660 15152 700 15184
rect 732 15152 772 15184
rect 804 15152 844 15184
rect 876 15152 1000 15184
rect 0 15112 1000 15152
rect 0 15080 124 15112
rect 156 15080 196 15112
rect 228 15080 268 15112
rect 300 15080 340 15112
rect 372 15080 412 15112
rect 444 15080 484 15112
rect 516 15080 556 15112
rect 588 15080 628 15112
rect 660 15080 700 15112
rect 732 15080 772 15112
rect 804 15080 844 15112
rect 876 15080 1000 15112
rect 0 15040 1000 15080
rect 0 15008 124 15040
rect 156 15008 196 15040
rect 228 15008 268 15040
rect 300 15008 340 15040
rect 372 15008 412 15040
rect 444 15008 484 15040
rect 516 15008 556 15040
rect 588 15008 628 15040
rect 660 15008 700 15040
rect 732 15008 772 15040
rect 804 15008 844 15040
rect 876 15008 1000 15040
rect 0 14968 1000 15008
rect 0 14936 124 14968
rect 156 14936 196 14968
rect 228 14936 268 14968
rect 300 14936 340 14968
rect 372 14936 412 14968
rect 444 14936 484 14968
rect 516 14936 556 14968
rect 588 14936 628 14968
rect 660 14936 700 14968
rect 732 14936 772 14968
rect 804 14936 844 14968
rect 876 14936 1000 14968
rect 0 14896 1000 14936
rect 0 14864 124 14896
rect 156 14864 196 14896
rect 228 14864 268 14896
rect 300 14864 340 14896
rect 372 14864 412 14896
rect 444 14864 484 14896
rect 516 14864 556 14896
rect 588 14864 628 14896
rect 660 14864 700 14896
rect 732 14864 772 14896
rect 804 14864 844 14896
rect 876 14864 1000 14896
rect 0 14824 1000 14864
rect 0 14792 124 14824
rect 156 14792 196 14824
rect 228 14792 268 14824
rect 300 14792 340 14824
rect 372 14792 412 14824
rect 444 14792 484 14824
rect 516 14792 556 14824
rect 588 14792 628 14824
rect 660 14792 700 14824
rect 732 14792 772 14824
rect 804 14792 844 14824
rect 876 14792 1000 14824
rect 0 14752 1000 14792
rect 0 14720 124 14752
rect 156 14720 196 14752
rect 228 14720 268 14752
rect 300 14720 340 14752
rect 372 14720 412 14752
rect 444 14720 484 14752
rect 516 14720 556 14752
rect 588 14720 628 14752
rect 660 14720 700 14752
rect 732 14720 772 14752
rect 804 14720 844 14752
rect 876 14720 1000 14752
rect 0 14680 1000 14720
rect 0 14648 124 14680
rect 156 14648 196 14680
rect 228 14648 268 14680
rect 300 14648 340 14680
rect 372 14648 412 14680
rect 444 14648 484 14680
rect 516 14648 556 14680
rect 588 14648 628 14680
rect 660 14648 700 14680
rect 732 14648 772 14680
rect 804 14648 844 14680
rect 876 14648 1000 14680
rect 0 14608 1000 14648
rect 0 14576 124 14608
rect 156 14576 196 14608
rect 228 14576 268 14608
rect 300 14576 340 14608
rect 372 14576 412 14608
rect 444 14576 484 14608
rect 516 14576 556 14608
rect 588 14576 628 14608
rect 660 14576 700 14608
rect 732 14576 772 14608
rect 804 14576 844 14608
rect 876 14576 1000 14608
rect 0 14536 1000 14576
rect 0 14504 124 14536
rect 156 14504 196 14536
rect 228 14504 268 14536
rect 300 14504 340 14536
rect 372 14504 412 14536
rect 444 14504 484 14536
rect 516 14504 556 14536
rect 588 14504 628 14536
rect 660 14504 700 14536
rect 732 14504 772 14536
rect 804 14504 844 14536
rect 876 14504 1000 14536
rect 0 14464 1000 14504
rect 0 14432 124 14464
rect 156 14432 196 14464
rect 228 14432 268 14464
rect 300 14432 340 14464
rect 372 14432 412 14464
rect 444 14432 484 14464
rect 516 14432 556 14464
rect 588 14432 628 14464
rect 660 14432 700 14464
rect 732 14432 772 14464
rect 804 14432 844 14464
rect 876 14432 1000 14464
rect 0 14392 1000 14432
rect 0 14360 124 14392
rect 156 14360 196 14392
rect 228 14360 268 14392
rect 300 14360 340 14392
rect 372 14360 412 14392
rect 444 14360 484 14392
rect 516 14360 556 14392
rect 588 14360 628 14392
rect 660 14360 700 14392
rect 732 14360 772 14392
rect 804 14360 844 14392
rect 876 14360 1000 14392
rect 0 14320 1000 14360
rect 0 14288 124 14320
rect 156 14288 196 14320
rect 228 14288 268 14320
rect 300 14288 340 14320
rect 372 14288 412 14320
rect 444 14288 484 14320
rect 516 14288 556 14320
rect 588 14288 628 14320
rect 660 14288 700 14320
rect 732 14288 772 14320
rect 804 14288 844 14320
rect 876 14288 1000 14320
rect 0 14248 1000 14288
rect 0 14216 124 14248
rect 156 14216 196 14248
rect 228 14216 268 14248
rect 300 14216 340 14248
rect 372 14216 412 14248
rect 444 14216 484 14248
rect 516 14216 556 14248
rect 588 14216 628 14248
rect 660 14216 700 14248
rect 732 14216 772 14248
rect 804 14216 844 14248
rect 876 14216 1000 14248
rect 0 14176 1000 14216
rect 0 14144 124 14176
rect 156 14144 196 14176
rect 228 14144 268 14176
rect 300 14144 340 14176
rect 372 14144 412 14176
rect 444 14144 484 14176
rect 516 14144 556 14176
rect 588 14144 628 14176
rect 660 14144 700 14176
rect 732 14144 772 14176
rect 804 14144 844 14176
rect 876 14144 1000 14176
rect 0 14104 1000 14144
rect 0 14072 124 14104
rect 156 14072 196 14104
rect 228 14072 268 14104
rect 300 14072 340 14104
rect 372 14072 412 14104
rect 444 14072 484 14104
rect 516 14072 556 14104
rect 588 14072 628 14104
rect 660 14072 700 14104
rect 732 14072 772 14104
rect 804 14072 844 14104
rect 876 14072 1000 14104
rect 0 14032 1000 14072
rect 0 14000 124 14032
rect 156 14000 196 14032
rect 228 14000 268 14032
rect 300 14000 340 14032
rect 372 14000 412 14032
rect 444 14000 484 14032
rect 516 14000 556 14032
rect 588 14000 628 14032
rect 660 14000 700 14032
rect 732 14000 772 14032
rect 804 14000 844 14032
rect 876 14000 1000 14032
rect 0 13960 1000 14000
rect 0 13928 124 13960
rect 156 13928 196 13960
rect 228 13928 268 13960
rect 300 13928 340 13960
rect 372 13928 412 13960
rect 444 13928 484 13960
rect 516 13928 556 13960
rect 588 13928 628 13960
rect 660 13928 700 13960
rect 732 13928 772 13960
rect 804 13928 844 13960
rect 876 13928 1000 13960
rect 0 13888 1000 13928
rect 0 13856 124 13888
rect 156 13856 196 13888
rect 228 13856 268 13888
rect 300 13856 340 13888
rect 372 13856 412 13888
rect 444 13856 484 13888
rect 516 13856 556 13888
rect 588 13856 628 13888
rect 660 13856 700 13888
rect 732 13856 772 13888
rect 804 13856 844 13888
rect 876 13856 1000 13888
rect 0 13816 1000 13856
rect 0 13784 124 13816
rect 156 13784 196 13816
rect 228 13784 268 13816
rect 300 13784 340 13816
rect 372 13784 412 13816
rect 444 13784 484 13816
rect 516 13784 556 13816
rect 588 13784 628 13816
rect 660 13784 700 13816
rect 732 13784 772 13816
rect 804 13784 844 13816
rect 876 13784 1000 13816
rect 0 13744 1000 13784
rect 0 13712 124 13744
rect 156 13712 196 13744
rect 228 13712 268 13744
rect 300 13712 340 13744
rect 372 13712 412 13744
rect 444 13712 484 13744
rect 516 13712 556 13744
rect 588 13712 628 13744
rect 660 13712 700 13744
rect 732 13712 772 13744
rect 804 13712 844 13744
rect 876 13712 1000 13744
rect 0 13672 1000 13712
rect 0 13640 124 13672
rect 156 13640 196 13672
rect 228 13640 268 13672
rect 300 13640 340 13672
rect 372 13640 412 13672
rect 444 13640 484 13672
rect 516 13640 556 13672
rect 588 13640 628 13672
rect 660 13640 700 13672
rect 732 13640 772 13672
rect 804 13640 844 13672
rect 876 13640 1000 13672
rect 0 13600 1000 13640
rect 0 13568 124 13600
rect 156 13568 196 13600
rect 228 13568 268 13600
rect 300 13568 340 13600
rect 372 13568 412 13600
rect 444 13568 484 13600
rect 516 13568 556 13600
rect 588 13568 628 13600
rect 660 13568 700 13600
rect 732 13568 772 13600
rect 804 13568 844 13600
rect 876 13568 1000 13600
rect 0 13528 1000 13568
rect 0 13496 124 13528
rect 156 13496 196 13528
rect 228 13496 268 13528
rect 300 13496 340 13528
rect 372 13496 412 13528
rect 444 13496 484 13528
rect 516 13496 556 13528
rect 588 13496 628 13528
rect 660 13496 700 13528
rect 732 13496 772 13528
rect 804 13496 844 13528
rect 876 13496 1000 13528
rect 0 13456 1000 13496
rect 0 13424 124 13456
rect 156 13424 196 13456
rect 228 13424 268 13456
rect 300 13424 340 13456
rect 372 13424 412 13456
rect 444 13424 484 13456
rect 516 13424 556 13456
rect 588 13424 628 13456
rect 660 13424 700 13456
rect 732 13424 772 13456
rect 804 13424 844 13456
rect 876 13424 1000 13456
rect 0 13384 1000 13424
rect 0 13352 124 13384
rect 156 13352 196 13384
rect 228 13352 268 13384
rect 300 13352 340 13384
rect 372 13352 412 13384
rect 444 13352 484 13384
rect 516 13352 556 13384
rect 588 13352 628 13384
rect 660 13352 700 13384
rect 732 13352 772 13384
rect 804 13352 844 13384
rect 876 13352 1000 13384
rect 0 13312 1000 13352
rect 0 13280 124 13312
rect 156 13280 196 13312
rect 228 13280 268 13312
rect 300 13280 340 13312
rect 372 13280 412 13312
rect 444 13280 484 13312
rect 516 13280 556 13312
rect 588 13280 628 13312
rect 660 13280 700 13312
rect 732 13280 772 13312
rect 804 13280 844 13312
rect 876 13280 1000 13312
rect 0 13240 1000 13280
rect 0 13208 124 13240
rect 156 13208 196 13240
rect 228 13208 268 13240
rect 300 13208 340 13240
rect 372 13208 412 13240
rect 444 13208 484 13240
rect 516 13208 556 13240
rect 588 13208 628 13240
rect 660 13208 700 13240
rect 732 13208 772 13240
rect 804 13208 844 13240
rect 876 13208 1000 13240
rect 0 13168 1000 13208
rect 0 13136 124 13168
rect 156 13136 196 13168
rect 228 13136 268 13168
rect 300 13136 340 13168
rect 372 13136 412 13168
rect 444 13136 484 13168
rect 516 13136 556 13168
rect 588 13136 628 13168
rect 660 13136 700 13168
rect 732 13136 772 13168
rect 804 13136 844 13168
rect 876 13136 1000 13168
rect 0 13096 1000 13136
rect 0 13064 124 13096
rect 156 13064 196 13096
rect 228 13064 268 13096
rect 300 13064 340 13096
rect 372 13064 412 13096
rect 444 13064 484 13096
rect 516 13064 556 13096
rect 588 13064 628 13096
rect 660 13064 700 13096
rect 732 13064 772 13096
rect 804 13064 844 13096
rect 876 13064 1000 13096
rect 0 13000 1000 13064
rect 0 12144 1000 12200
rect 0 12112 52 12144
rect 84 12112 124 12144
rect 156 12112 196 12144
rect 228 12112 268 12144
rect 300 12112 340 12144
rect 372 12112 412 12144
rect 444 12112 484 12144
rect 516 12112 556 12144
rect 588 12112 628 12144
rect 660 12112 700 12144
rect 732 12112 772 12144
rect 804 12112 844 12144
rect 876 12112 916 12144
rect 948 12112 1000 12144
rect 0 12072 1000 12112
rect 0 12040 52 12072
rect 84 12040 124 12072
rect 156 12040 196 12072
rect 228 12040 268 12072
rect 300 12040 340 12072
rect 372 12040 412 12072
rect 444 12040 484 12072
rect 516 12040 556 12072
rect 588 12040 628 12072
rect 660 12040 700 12072
rect 732 12040 772 12072
rect 804 12040 844 12072
rect 876 12040 916 12072
rect 948 12040 1000 12072
rect 0 12000 1000 12040
rect 0 11968 52 12000
rect 84 11968 124 12000
rect 156 11968 196 12000
rect 228 11968 268 12000
rect 300 11968 340 12000
rect 372 11968 412 12000
rect 444 11968 484 12000
rect 516 11968 556 12000
rect 588 11968 628 12000
rect 660 11968 700 12000
rect 732 11968 772 12000
rect 804 11968 844 12000
rect 876 11968 916 12000
rect 948 11968 1000 12000
rect 0 11928 1000 11968
rect 0 11896 52 11928
rect 84 11896 124 11928
rect 156 11896 196 11928
rect 228 11896 268 11928
rect 300 11896 340 11928
rect 372 11896 412 11928
rect 444 11896 484 11928
rect 516 11896 556 11928
rect 588 11896 628 11928
rect 660 11896 700 11928
rect 732 11896 772 11928
rect 804 11896 844 11928
rect 876 11896 916 11928
rect 948 11896 1000 11928
rect 0 11856 1000 11896
rect 0 11824 52 11856
rect 84 11824 124 11856
rect 156 11824 196 11856
rect 228 11824 268 11856
rect 300 11824 340 11856
rect 372 11824 412 11856
rect 444 11824 484 11856
rect 516 11824 556 11856
rect 588 11824 628 11856
rect 660 11824 700 11856
rect 732 11824 772 11856
rect 804 11824 844 11856
rect 876 11824 916 11856
rect 948 11824 1000 11856
rect 0 11784 1000 11824
rect 0 11752 52 11784
rect 84 11752 124 11784
rect 156 11752 196 11784
rect 228 11752 268 11784
rect 300 11752 340 11784
rect 372 11752 412 11784
rect 444 11752 484 11784
rect 516 11752 556 11784
rect 588 11752 628 11784
rect 660 11752 700 11784
rect 732 11752 772 11784
rect 804 11752 844 11784
rect 876 11752 916 11784
rect 948 11752 1000 11784
rect 0 11712 1000 11752
rect 0 11680 52 11712
rect 84 11680 124 11712
rect 156 11680 196 11712
rect 228 11680 268 11712
rect 300 11680 340 11712
rect 372 11680 412 11712
rect 444 11680 484 11712
rect 516 11680 556 11712
rect 588 11680 628 11712
rect 660 11680 700 11712
rect 732 11680 772 11712
rect 804 11680 844 11712
rect 876 11680 916 11712
rect 948 11680 1000 11712
rect 0 11640 1000 11680
rect 0 11608 52 11640
rect 84 11608 124 11640
rect 156 11608 196 11640
rect 228 11608 268 11640
rect 300 11608 340 11640
rect 372 11608 412 11640
rect 444 11608 484 11640
rect 516 11608 556 11640
rect 588 11608 628 11640
rect 660 11608 700 11640
rect 732 11608 772 11640
rect 804 11608 844 11640
rect 876 11608 916 11640
rect 948 11608 1000 11640
rect 0 11568 1000 11608
rect 0 11536 52 11568
rect 84 11536 124 11568
rect 156 11536 196 11568
rect 228 11536 268 11568
rect 300 11536 340 11568
rect 372 11536 412 11568
rect 444 11536 484 11568
rect 516 11536 556 11568
rect 588 11536 628 11568
rect 660 11536 700 11568
rect 732 11536 772 11568
rect 804 11536 844 11568
rect 876 11536 916 11568
rect 948 11536 1000 11568
rect 0 11496 1000 11536
rect 0 11464 52 11496
rect 84 11464 124 11496
rect 156 11464 196 11496
rect 228 11464 268 11496
rect 300 11464 340 11496
rect 372 11464 412 11496
rect 444 11464 484 11496
rect 516 11464 556 11496
rect 588 11464 628 11496
rect 660 11464 700 11496
rect 732 11464 772 11496
rect 804 11464 844 11496
rect 876 11464 916 11496
rect 948 11464 1000 11496
rect 0 11424 1000 11464
rect 0 11392 52 11424
rect 84 11392 124 11424
rect 156 11392 196 11424
rect 228 11392 268 11424
rect 300 11392 340 11424
rect 372 11392 412 11424
rect 444 11392 484 11424
rect 516 11392 556 11424
rect 588 11392 628 11424
rect 660 11392 700 11424
rect 732 11392 772 11424
rect 804 11392 844 11424
rect 876 11392 916 11424
rect 948 11392 1000 11424
rect 0 11352 1000 11392
rect 0 11320 52 11352
rect 84 11320 124 11352
rect 156 11320 196 11352
rect 228 11320 268 11352
rect 300 11320 340 11352
rect 372 11320 412 11352
rect 444 11320 484 11352
rect 516 11320 556 11352
rect 588 11320 628 11352
rect 660 11320 700 11352
rect 732 11320 772 11352
rect 804 11320 844 11352
rect 876 11320 916 11352
rect 948 11320 1000 11352
rect 0 11280 1000 11320
rect 0 11248 52 11280
rect 84 11248 124 11280
rect 156 11248 196 11280
rect 228 11248 268 11280
rect 300 11248 340 11280
rect 372 11248 412 11280
rect 444 11248 484 11280
rect 516 11248 556 11280
rect 588 11248 628 11280
rect 660 11248 700 11280
rect 732 11248 772 11280
rect 804 11248 844 11280
rect 876 11248 916 11280
rect 948 11248 1000 11280
rect 0 11208 1000 11248
rect 0 11176 52 11208
rect 84 11176 124 11208
rect 156 11176 196 11208
rect 228 11176 268 11208
rect 300 11176 340 11208
rect 372 11176 412 11208
rect 444 11176 484 11208
rect 516 11176 556 11208
rect 588 11176 628 11208
rect 660 11176 700 11208
rect 732 11176 772 11208
rect 804 11176 844 11208
rect 876 11176 916 11208
rect 948 11176 1000 11208
rect 0 11136 1000 11176
rect 0 11104 52 11136
rect 84 11104 124 11136
rect 156 11104 196 11136
rect 228 11104 268 11136
rect 300 11104 340 11136
rect 372 11104 412 11136
rect 444 11104 484 11136
rect 516 11104 556 11136
rect 588 11104 628 11136
rect 660 11104 700 11136
rect 732 11104 772 11136
rect 804 11104 844 11136
rect 876 11104 916 11136
rect 948 11104 1000 11136
rect 0 11064 1000 11104
rect 0 11032 52 11064
rect 84 11032 124 11064
rect 156 11032 196 11064
rect 228 11032 268 11064
rect 300 11032 340 11064
rect 372 11032 412 11064
rect 444 11032 484 11064
rect 516 11032 556 11064
rect 588 11032 628 11064
rect 660 11032 700 11064
rect 732 11032 772 11064
rect 804 11032 844 11064
rect 876 11032 916 11064
rect 948 11032 1000 11064
rect 0 10992 1000 11032
rect 0 10960 52 10992
rect 84 10960 124 10992
rect 156 10960 196 10992
rect 228 10960 268 10992
rect 300 10960 340 10992
rect 372 10960 412 10992
rect 444 10960 484 10992
rect 516 10960 556 10992
rect 588 10960 628 10992
rect 660 10960 700 10992
rect 732 10960 772 10992
rect 804 10960 844 10992
rect 876 10960 916 10992
rect 948 10960 1000 10992
rect 0 10920 1000 10960
rect 0 10888 52 10920
rect 84 10888 124 10920
rect 156 10888 196 10920
rect 228 10888 268 10920
rect 300 10888 340 10920
rect 372 10888 412 10920
rect 444 10888 484 10920
rect 516 10888 556 10920
rect 588 10888 628 10920
rect 660 10888 700 10920
rect 732 10888 772 10920
rect 804 10888 844 10920
rect 876 10888 916 10920
rect 948 10888 1000 10920
rect 0 10848 1000 10888
rect 0 10816 52 10848
rect 84 10816 124 10848
rect 156 10816 196 10848
rect 228 10816 268 10848
rect 300 10816 340 10848
rect 372 10816 412 10848
rect 444 10816 484 10848
rect 516 10816 556 10848
rect 588 10816 628 10848
rect 660 10816 700 10848
rect 732 10816 772 10848
rect 804 10816 844 10848
rect 876 10816 916 10848
rect 948 10816 1000 10848
rect 0 10776 1000 10816
rect 0 10744 52 10776
rect 84 10744 124 10776
rect 156 10744 196 10776
rect 228 10744 268 10776
rect 300 10744 340 10776
rect 372 10744 412 10776
rect 444 10744 484 10776
rect 516 10744 556 10776
rect 588 10744 628 10776
rect 660 10744 700 10776
rect 732 10744 772 10776
rect 804 10744 844 10776
rect 876 10744 916 10776
rect 948 10744 1000 10776
rect 0 10704 1000 10744
rect 0 10672 52 10704
rect 84 10672 124 10704
rect 156 10672 196 10704
rect 228 10672 268 10704
rect 300 10672 340 10704
rect 372 10672 412 10704
rect 444 10672 484 10704
rect 516 10672 556 10704
rect 588 10672 628 10704
rect 660 10672 700 10704
rect 732 10672 772 10704
rect 804 10672 844 10704
rect 876 10672 916 10704
rect 948 10672 1000 10704
rect 0 10632 1000 10672
rect 0 10600 52 10632
rect 84 10600 124 10632
rect 156 10600 196 10632
rect 228 10600 268 10632
rect 300 10600 340 10632
rect 372 10600 412 10632
rect 444 10600 484 10632
rect 516 10600 556 10632
rect 588 10600 628 10632
rect 660 10600 700 10632
rect 732 10600 772 10632
rect 804 10600 844 10632
rect 876 10600 916 10632
rect 948 10600 1000 10632
rect 0 10560 1000 10600
rect 0 10528 52 10560
rect 84 10528 124 10560
rect 156 10528 196 10560
rect 228 10528 268 10560
rect 300 10528 340 10560
rect 372 10528 412 10560
rect 444 10528 484 10560
rect 516 10528 556 10560
rect 588 10528 628 10560
rect 660 10528 700 10560
rect 732 10528 772 10560
rect 804 10528 844 10560
rect 876 10528 916 10560
rect 948 10528 1000 10560
rect 0 10488 1000 10528
rect 0 10456 52 10488
rect 84 10456 124 10488
rect 156 10456 196 10488
rect 228 10456 268 10488
rect 300 10456 340 10488
rect 372 10456 412 10488
rect 444 10456 484 10488
rect 516 10456 556 10488
rect 588 10456 628 10488
rect 660 10456 700 10488
rect 732 10456 772 10488
rect 804 10456 844 10488
rect 876 10456 916 10488
rect 948 10456 1000 10488
rect 0 10416 1000 10456
rect 0 10384 52 10416
rect 84 10384 124 10416
rect 156 10384 196 10416
rect 228 10384 268 10416
rect 300 10384 340 10416
rect 372 10384 412 10416
rect 444 10384 484 10416
rect 516 10384 556 10416
rect 588 10384 628 10416
rect 660 10384 700 10416
rect 732 10384 772 10416
rect 804 10384 844 10416
rect 876 10384 916 10416
rect 948 10384 1000 10416
rect 0 10344 1000 10384
rect 0 10312 52 10344
rect 84 10312 124 10344
rect 156 10312 196 10344
rect 228 10312 268 10344
rect 300 10312 340 10344
rect 372 10312 412 10344
rect 444 10312 484 10344
rect 516 10312 556 10344
rect 588 10312 628 10344
rect 660 10312 700 10344
rect 732 10312 772 10344
rect 804 10312 844 10344
rect 876 10312 916 10344
rect 948 10312 1000 10344
rect 0 10272 1000 10312
rect 0 10240 52 10272
rect 84 10240 124 10272
rect 156 10240 196 10272
rect 228 10240 268 10272
rect 300 10240 340 10272
rect 372 10240 412 10272
rect 444 10240 484 10272
rect 516 10240 556 10272
rect 588 10240 628 10272
rect 660 10240 700 10272
rect 732 10240 772 10272
rect 804 10240 844 10272
rect 876 10240 916 10272
rect 948 10240 1000 10272
rect 0 10200 1000 10240
rect 0 10168 52 10200
rect 84 10168 124 10200
rect 156 10168 196 10200
rect 228 10168 268 10200
rect 300 10168 340 10200
rect 372 10168 412 10200
rect 444 10168 484 10200
rect 516 10168 556 10200
rect 588 10168 628 10200
rect 660 10168 700 10200
rect 732 10168 772 10200
rect 804 10168 844 10200
rect 876 10168 916 10200
rect 948 10168 1000 10200
rect 0 10128 1000 10168
rect 0 10096 52 10128
rect 84 10096 124 10128
rect 156 10096 196 10128
rect 228 10096 268 10128
rect 300 10096 340 10128
rect 372 10096 412 10128
rect 444 10096 484 10128
rect 516 10096 556 10128
rect 588 10096 628 10128
rect 660 10096 700 10128
rect 732 10096 772 10128
rect 804 10096 844 10128
rect 876 10096 916 10128
rect 948 10096 1000 10128
rect 0 10056 1000 10096
rect 0 10024 52 10056
rect 84 10024 124 10056
rect 156 10024 196 10056
rect 228 10024 268 10056
rect 300 10024 340 10056
rect 372 10024 412 10056
rect 444 10024 484 10056
rect 516 10024 556 10056
rect 588 10024 628 10056
rect 660 10024 700 10056
rect 732 10024 772 10056
rect 804 10024 844 10056
rect 876 10024 916 10056
rect 948 10024 1000 10056
rect 0 9984 1000 10024
rect 0 9952 52 9984
rect 84 9952 124 9984
rect 156 9952 196 9984
rect 228 9952 268 9984
rect 300 9952 340 9984
rect 372 9952 412 9984
rect 444 9952 484 9984
rect 516 9952 556 9984
rect 588 9952 628 9984
rect 660 9952 700 9984
rect 732 9952 772 9984
rect 804 9952 844 9984
rect 876 9952 916 9984
rect 948 9952 1000 9984
rect 0 9912 1000 9952
rect 0 9880 52 9912
rect 84 9880 124 9912
rect 156 9880 196 9912
rect 228 9880 268 9912
rect 300 9880 340 9912
rect 372 9880 412 9912
rect 444 9880 484 9912
rect 516 9880 556 9912
rect 588 9880 628 9912
rect 660 9880 700 9912
rect 732 9880 772 9912
rect 804 9880 844 9912
rect 876 9880 916 9912
rect 948 9880 1000 9912
rect 0 9840 1000 9880
rect 0 9808 52 9840
rect 84 9808 124 9840
rect 156 9808 196 9840
rect 228 9808 268 9840
rect 300 9808 340 9840
rect 372 9808 412 9840
rect 444 9808 484 9840
rect 516 9808 556 9840
rect 588 9808 628 9840
rect 660 9808 700 9840
rect 732 9808 772 9840
rect 804 9808 844 9840
rect 876 9808 916 9840
rect 948 9808 1000 9840
rect 0 9768 1000 9808
rect 0 9736 52 9768
rect 84 9736 124 9768
rect 156 9736 196 9768
rect 228 9736 268 9768
rect 300 9736 340 9768
rect 372 9736 412 9768
rect 444 9736 484 9768
rect 516 9736 556 9768
rect 588 9736 628 9768
rect 660 9736 700 9768
rect 732 9736 772 9768
rect 804 9736 844 9768
rect 876 9736 916 9768
rect 948 9736 1000 9768
rect 0 9696 1000 9736
rect 0 9664 52 9696
rect 84 9664 124 9696
rect 156 9664 196 9696
rect 228 9664 268 9696
rect 300 9664 340 9696
rect 372 9664 412 9696
rect 444 9664 484 9696
rect 516 9664 556 9696
rect 588 9664 628 9696
rect 660 9664 700 9696
rect 732 9664 772 9696
rect 804 9664 844 9696
rect 876 9664 916 9696
rect 948 9664 1000 9696
rect 0 9624 1000 9664
rect 0 9592 52 9624
rect 84 9592 124 9624
rect 156 9592 196 9624
rect 228 9592 268 9624
rect 300 9592 340 9624
rect 372 9592 412 9624
rect 444 9592 484 9624
rect 516 9592 556 9624
rect 588 9592 628 9624
rect 660 9592 700 9624
rect 732 9592 772 9624
rect 804 9592 844 9624
rect 876 9592 916 9624
rect 948 9592 1000 9624
rect 0 9552 1000 9592
rect 0 9520 52 9552
rect 84 9520 124 9552
rect 156 9520 196 9552
rect 228 9520 268 9552
rect 300 9520 340 9552
rect 372 9520 412 9552
rect 444 9520 484 9552
rect 516 9520 556 9552
rect 588 9520 628 9552
rect 660 9520 700 9552
rect 732 9520 772 9552
rect 804 9520 844 9552
rect 876 9520 916 9552
rect 948 9520 1000 9552
rect 0 9480 1000 9520
rect 0 9448 52 9480
rect 84 9448 124 9480
rect 156 9448 196 9480
rect 228 9448 268 9480
rect 300 9448 340 9480
rect 372 9448 412 9480
rect 444 9448 484 9480
rect 516 9448 556 9480
rect 588 9448 628 9480
rect 660 9448 700 9480
rect 732 9448 772 9480
rect 804 9448 844 9480
rect 876 9448 916 9480
rect 948 9448 1000 9480
rect 0 9408 1000 9448
rect 0 9376 52 9408
rect 84 9376 124 9408
rect 156 9376 196 9408
rect 228 9376 268 9408
rect 300 9376 340 9408
rect 372 9376 412 9408
rect 444 9376 484 9408
rect 516 9376 556 9408
rect 588 9376 628 9408
rect 660 9376 700 9408
rect 732 9376 772 9408
rect 804 9376 844 9408
rect 876 9376 916 9408
rect 948 9376 1000 9408
rect 0 9336 1000 9376
rect 0 9304 52 9336
rect 84 9304 124 9336
rect 156 9304 196 9336
rect 228 9304 268 9336
rect 300 9304 340 9336
rect 372 9304 412 9336
rect 444 9304 484 9336
rect 516 9304 556 9336
rect 588 9304 628 9336
rect 660 9304 700 9336
rect 732 9304 772 9336
rect 804 9304 844 9336
rect 876 9304 916 9336
rect 948 9304 1000 9336
rect 0 9264 1000 9304
rect 0 9232 52 9264
rect 84 9232 124 9264
rect 156 9232 196 9264
rect 228 9232 268 9264
rect 300 9232 340 9264
rect 372 9232 412 9264
rect 444 9232 484 9264
rect 516 9232 556 9264
rect 588 9232 628 9264
rect 660 9232 700 9264
rect 732 9232 772 9264
rect 804 9232 844 9264
rect 876 9232 916 9264
rect 948 9232 1000 9264
rect 0 9192 1000 9232
rect 0 9160 52 9192
rect 84 9160 124 9192
rect 156 9160 196 9192
rect 228 9160 268 9192
rect 300 9160 340 9192
rect 372 9160 412 9192
rect 444 9160 484 9192
rect 516 9160 556 9192
rect 588 9160 628 9192
rect 660 9160 700 9192
rect 732 9160 772 9192
rect 804 9160 844 9192
rect 876 9160 916 9192
rect 948 9160 1000 9192
rect 0 9120 1000 9160
rect 0 9088 52 9120
rect 84 9088 124 9120
rect 156 9088 196 9120
rect 228 9088 268 9120
rect 300 9088 340 9120
rect 372 9088 412 9120
rect 444 9088 484 9120
rect 516 9088 556 9120
rect 588 9088 628 9120
rect 660 9088 700 9120
rect 732 9088 772 9120
rect 804 9088 844 9120
rect 876 9088 916 9120
rect 948 9088 1000 9120
rect 0 9048 1000 9088
rect 0 9016 52 9048
rect 84 9016 124 9048
rect 156 9016 196 9048
rect 228 9016 268 9048
rect 300 9016 340 9048
rect 372 9016 412 9048
rect 444 9016 484 9048
rect 516 9016 556 9048
rect 588 9016 628 9048
rect 660 9016 700 9048
rect 732 9016 772 9048
rect 804 9016 844 9048
rect 876 9016 916 9048
rect 948 9016 1000 9048
rect 0 8976 1000 9016
rect 0 8944 52 8976
rect 84 8944 124 8976
rect 156 8944 196 8976
rect 228 8944 268 8976
rect 300 8944 340 8976
rect 372 8944 412 8976
rect 444 8944 484 8976
rect 516 8944 556 8976
rect 588 8944 628 8976
rect 660 8944 700 8976
rect 732 8944 772 8976
rect 804 8944 844 8976
rect 876 8944 916 8976
rect 948 8944 1000 8976
rect 0 8904 1000 8944
rect 0 8872 52 8904
rect 84 8872 124 8904
rect 156 8872 196 8904
rect 228 8872 268 8904
rect 300 8872 340 8904
rect 372 8872 412 8904
rect 444 8872 484 8904
rect 516 8872 556 8904
rect 588 8872 628 8904
rect 660 8872 700 8904
rect 732 8872 772 8904
rect 804 8872 844 8904
rect 876 8872 916 8904
rect 948 8872 1000 8904
rect 0 8832 1000 8872
rect 0 8800 52 8832
rect 84 8800 124 8832
rect 156 8800 196 8832
rect 228 8800 268 8832
rect 300 8800 340 8832
rect 372 8800 412 8832
rect 444 8800 484 8832
rect 516 8800 556 8832
rect 588 8800 628 8832
rect 660 8800 700 8832
rect 732 8800 772 8832
rect 804 8800 844 8832
rect 876 8800 916 8832
rect 948 8800 1000 8832
rect 0 8760 1000 8800
rect 0 8728 52 8760
rect 84 8728 124 8760
rect 156 8728 196 8760
rect 228 8728 268 8760
rect 300 8728 340 8760
rect 372 8728 412 8760
rect 444 8728 484 8760
rect 516 8728 556 8760
rect 588 8728 628 8760
rect 660 8728 700 8760
rect 732 8728 772 8760
rect 804 8728 844 8760
rect 876 8728 916 8760
rect 948 8728 1000 8760
rect 0 8688 1000 8728
rect 0 8656 52 8688
rect 84 8656 124 8688
rect 156 8656 196 8688
rect 228 8656 268 8688
rect 300 8656 340 8688
rect 372 8656 412 8688
rect 444 8656 484 8688
rect 516 8656 556 8688
rect 588 8656 628 8688
rect 660 8656 700 8688
rect 732 8656 772 8688
rect 804 8656 844 8688
rect 876 8656 916 8688
rect 948 8656 1000 8688
rect 0 8616 1000 8656
rect 0 8584 52 8616
rect 84 8584 124 8616
rect 156 8584 196 8616
rect 228 8584 268 8616
rect 300 8584 340 8616
rect 372 8584 412 8616
rect 444 8584 484 8616
rect 516 8584 556 8616
rect 588 8584 628 8616
rect 660 8584 700 8616
rect 732 8584 772 8616
rect 804 8584 844 8616
rect 876 8584 916 8616
rect 948 8584 1000 8616
rect 0 8544 1000 8584
rect 0 8512 52 8544
rect 84 8512 124 8544
rect 156 8512 196 8544
rect 228 8512 268 8544
rect 300 8512 340 8544
rect 372 8512 412 8544
rect 444 8512 484 8544
rect 516 8512 556 8544
rect 588 8512 628 8544
rect 660 8512 700 8544
rect 732 8512 772 8544
rect 804 8512 844 8544
rect 876 8512 916 8544
rect 948 8512 1000 8544
rect 0 8472 1000 8512
rect 0 8440 52 8472
rect 84 8440 124 8472
rect 156 8440 196 8472
rect 228 8440 268 8472
rect 300 8440 340 8472
rect 372 8440 412 8472
rect 444 8440 484 8472
rect 516 8440 556 8472
rect 588 8440 628 8472
rect 660 8440 700 8472
rect 732 8440 772 8472
rect 804 8440 844 8472
rect 876 8440 916 8472
rect 948 8440 1000 8472
rect 0 8400 1000 8440
rect 0 8368 52 8400
rect 84 8368 124 8400
rect 156 8368 196 8400
rect 228 8368 268 8400
rect 300 8368 340 8400
rect 372 8368 412 8400
rect 444 8368 484 8400
rect 516 8368 556 8400
rect 588 8368 628 8400
rect 660 8368 700 8400
rect 732 8368 772 8400
rect 804 8368 844 8400
rect 876 8368 916 8400
rect 948 8368 1000 8400
rect 0 8328 1000 8368
rect 0 8296 52 8328
rect 84 8296 124 8328
rect 156 8296 196 8328
rect 228 8296 268 8328
rect 300 8296 340 8328
rect 372 8296 412 8328
rect 444 8296 484 8328
rect 516 8296 556 8328
rect 588 8296 628 8328
rect 660 8296 700 8328
rect 732 8296 772 8328
rect 804 8296 844 8328
rect 876 8296 916 8328
rect 948 8296 1000 8328
rect 0 8256 1000 8296
rect 0 8224 52 8256
rect 84 8224 124 8256
rect 156 8224 196 8256
rect 228 8224 268 8256
rect 300 8224 340 8256
rect 372 8224 412 8256
rect 444 8224 484 8256
rect 516 8224 556 8256
rect 588 8224 628 8256
rect 660 8224 700 8256
rect 732 8224 772 8256
rect 804 8224 844 8256
rect 876 8224 916 8256
rect 948 8224 1000 8256
rect 0 8184 1000 8224
rect 0 8152 52 8184
rect 84 8152 124 8184
rect 156 8152 196 8184
rect 228 8152 268 8184
rect 300 8152 340 8184
rect 372 8152 412 8184
rect 444 8152 484 8184
rect 516 8152 556 8184
rect 588 8152 628 8184
rect 660 8152 700 8184
rect 732 8152 772 8184
rect 804 8152 844 8184
rect 876 8152 916 8184
rect 948 8152 1000 8184
rect 0 8112 1000 8152
rect 0 8080 52 8112
rect 84 8080 124 8112
rect 156 8080 196 8112
rect 228 8080 268 8112
rect 300 8080 340 8112
rect 372 8080 412 8112
rect 444 8080 484 8112
rect 516 8080 556 8112
rect 588 8080 628 8112
rect 660 8080 700 8112
rect 732 8080 772 8112
rect 804 8080 844 8112
rect 876 8080 916 8112
rect 948 8080 1000 8112
rect 0 8040 1000 8080
rect 0 8008 52 8040
rect 84 8008 124 8040
rect 156 8008 196 8040
rect 228 8008 268 8040
rect 300 8008 340 8040
rect 372 8008 412 8040
rect 444 8008 484 8040
rect 516 8008 556 8040
rect 588 8008 628 8040
rect 660 8008 700 8040
rect 732 8008 772 8040
rect 804 8008 844 8040
rect 876 8008 916 8040
rect 948 8008 1000 8040
rect 0 7968 1000 8008
rect 0 7936 52 7968
rect 84 7936 124 7968
rect 156 7936 196 7968
rect 228 7936 268 7968
rect 300 7936 340 7968
rect 372 7936 412 7968
rect 444 7936 484 7968
rect 516 7936 556 7968
rect 588 7936 628 7968
rect 660 7936 700 7968
rect 732 7936 772 7968
rect 804 7936 844 7968
rect 876 7936 916 7968
rect 948 7936 1000 7968
rect 0 7896 1000 7936
rect 0 7864 52 7896
rect 84 7864 124 7896
rect 156 7864 196 7896
rect 228 7864 268 7896
rect 300 7864 340 7896
rect 372 7864 412 7896
rect 444 7864 484 7896
rect 516 7864 556 7896
rect 588 7864 628 7896
rect 660 7864 700 7896
rect 732 7864 772 7896
rect 804 7864 844 7896
rect 876 7864 916 7896
rect 948 7864 1000 7896
rect 0 7824 1000 7864
rect 0 7792 52 7824
rect 84 7792 124 7824
rect 156 7792 196 7824
rect 228 7792 268 7824
rect 300 7792 340 7824
rect 372 7792 412 7824
rect 444 7792 484 7824
rect 516 7792 556 7824
rect 588 7792 628 7824
rect 660 7792 700 7824
rect 732 7792 772 7824
rect 804 7792 844 7824
rect 876 7792 916 7824
rect 948 7792 1000 7824
rect 0 7752 1000 7792
rect 0 7720 52 7752
rect 84 7720 124 7752
rect 156 7720 196 7752
rect 228 7720 268 7752
rect 300 7720 340 7752
rect 372 7720 412 7752
rect 444 7720 484 7752
rect 516 7720 556 7752
rect 588 7720 628 7752
rect 660 7720 700 7752
rect 732 7720 772 7752
rect 804 7720 844 7752
rect 876 7720 916 7752
rect 948 7720 1000 7752
rect 0 7680 1000 7720
rect 0 7648 52 7680
rect 84 7648 124 7680
rect 156 7648 196 7680
rect 228 7648 268 7680
rect 300 7648 340 7680
rect 372 7648 412 7680
rect 444 7648 484 7680
rect 516 7648 556 7680
rect 588 7648 628 7680
rect 660 7648 700 7680
rect 732 7648 772 7680
rect 804 7648 844 7680
rect 876 7648 916 7680
rect 948 7648 1000 7680
rect 0 7608 1000 7648
rect 0 7576 52 7608
rect 84 7576 124 7608
rect 156 7576 196 7608
rect 228 7576 268 7608
rect 300 7576 340 7608
rect 372 7576 412 7608
rect 444 7576 484 7608
rect 516 7576 556 7608
rect 588 7576 628 7608
rect 660 7576 700 7608
rect 732 7576 772 7608
rect 804 7576 844 7608
rect 876 7576 916 7608
rect 948 7576 1000 7608
rect 0 7536 1000 7576
rect 0 7504 52 7536
rect 84 7504 124 7536
rect 156 7504 196 7536
rect 228 7504 268 7536
rect 300 7504 340 7536
rect 372 7504 412 7536
rect 444 7504 484 7536
rect 516 7504 556 7536
rect 588 7504 628 7536
rect 660 7504 700 7536
rect 732 7504 772 7536
rect 804 7504 844 7536
rect 876 7504 916 7536
rect 948 7504 1000 7536
rect 0 7464 1000 7504
rect 0 7432 52 7464
rect 84 7432 124 7464
rect 156 7432 196 7464
rect 228 7432 268 7464
rect 300 7432 340 7464
rect 372 7432 412 7464
rect 444 7432 484 7464
rect 516 7432 556 7464
rect 588 7432 628 7464
rect 660 7432 700 7464
rect 732 7432 772 7464
rect 804 7432 844 7464
rect 876 7432 916 7464
rect 948 7432 1000 7464
rect 0 7392 1000 7432
rect 0 7360 52 7392
rect 84 7360 124 7392
rect 156 7360 196 7392
rect 228 7360 268 7392
rect 300 7360 340 7392
rect 372 7360 412 7392
rect 444 7360 484 7392
rect 516 7360 556 7392
rect 588 7360 628 7392
rect 660 7360 700 7392
rect 732 7360 772 7392
rect 804 7360 844 7392
rect 876 7360 916 7392
rect 948 7360 1000 7392
rect 0 7320 1000 7360
rect 0 7288 52 7320
rect 84 7288 124 7320
rect 156 7288 196 7320
rect 228 7288 268 7320
rect 300 7288 340 7320
rect 372 7288 412 7320
rect 444 7288 484 7320
rect 516 7288 556 7320
rect 588 7288 628 7320
rect 660 7288 700 7320
rect 732 7288 772 7320
rect 804 7288 844 7320
rect 876 7288 916 7320
rect 948 7288 1000 7320
rect 0 7248 1000 7288
rect 0 7216 52 7248
rect 84 7216 124 7248
rect 156 7216 196 7248
rect 228 7216 268 7248
rect 300 7216 340 7248
rect 372 7216 412 7248
rect 444 7216 484 7248
rect 516 7216 556 7248
rect 588 7216 628 7248
rect 660 7216 700 7248
rect 732 7216 772 7248
rect 804 7216 844 7248
rect 876 7216 916 7248
rect 948 7216 1000 7248
rect 0 7176 1000 7216
rect 0 7144 52 7176
rect 84 7144 124 7176
rect 156 7144 196 7176
rect 228 7144 268 7176
rect 300 7144 340 7176
rect 372 7144 412 7176
rect 444 7144 484 7176
rect 516 7144 556 7176
rect 588 7144 628 7176
rect 660 7144 700 7176
rect 732 7144 772 7176
rect 804 7144 844 7176
rect 876 7144 916 7176
rect 948 7144 1000 7176
rect 0 7104 1000 7144
rect 0 7072 52 7104
rect 84 7072 124 7104
rect 156 7072 196 7104
rect 228 7072 268 7104
rect 300 7072 340 7104
rect 372 7072 412 7104
rect 444 7072 484 7104
rect 516 7072 556 7104
rect 588 7072 628 7104
rect 660 7072 700 7104
rect 732 7072 772 7104
rect 804 7072 844 7104
rect 876 7072 916 7104
rect 948 7072 1000 7104
rect 0 7032 1000 7072
rect 0 7000 52 7032
rect 84 7000 124 7032
rect 156 7000 196 7032
rect 228 7000 268 7032
rect 300 7000 340 7032
rect 372 7000 412 7032
rect 444 7000 484 7032
rect 516 7000 556 7032
rect 588 7000 628 7032
rect 660 7000 700 7032
rect 732 7000 772 7032
rect 804 7000 844 7032
rect 876 7000 916 7032
rect 948 7000 1000 7032
rect 0 6960 1000 7000
rect 0 6928 52 6960
rect 84 6928 124 6960
rect 156 6928 196 6960
rect 228 6928 268 6960
rect 300 6928 340 6960
rect 372 6928 412 6960
rect 444 6928 484 6960
rect 516 6928 556 6960
rect 588 6928 628 6960
rect 660 6928 700 6960
rect 732 6928 772 6960
rect 804 6928 844 6960
rect 876 6928 916 6960
rect 948 6928 1000 6960
rect 0 6888 1000 6928
rect 0 6856 52 6888
rect 84 6856 124 6888
rect 156 6856 196 6888
rect 228 6856 268 6888
rect 300 6856 340 6888
rect 372 6856 412 6888
rect 444 6856 484 6888
rect 516 6856 556 6888
rect 588 6856 628 6888
rect 660 6856 700 6888
rect 732 6856 772 6888
rect 804 6856 844 6888
rect 876 6856 916 6888
rect 948 6856 1000 6888
rect 0 6800 1000 6856
rect 0 6544 1000 6600
rect 0 6512 52 6544
rect 84 6512 124 6544
rect 156 6512 196 6544
rect 228 6512 268 6544
rect 300 6512 340 6544
rect 372 6512 412 6544
rect 444 6512 484 6544
rect 516 6512 556 6544
rect 588 6512 628 6544
rect 660 6512 700 6544
rect 732 6512 772 6544
rect 804 6512 844 6544
rect 876 6512 916 6544
rect 948 6512 1000 6544
rect 0 6472 1000 6512
rect 0 6440 52 6472
rect 84 6440 124 6472
rect 156 6440 196 6472
rect 228 6440 268 6472
rect 300 6440 340 6472
rect 372 6440 412 6472
rect 444 6440 484 6472
rect 516 6440 556 6472
rect 588 6440 628 6472
rect 660 6440 700 6472
rect 732 6440 772 6472
rect 804 6440 844 6472
rect 876 6440 916 6472
rect 948 6440 1000 6472
rect 0 6400 1000 6440
rect 0 6368 52 6400
rect 84 6368 124 6400
rect 156 6368 196 6400
rect 228 6368 268 6400
rect 300 6368 340 6400
rect 372 6368 412 6400
rect 444 6368 484 6400
rect 516 6368 556 6400
rect 588 6368 628 6400
rect 660 6368 700 6400
rect 732 6368 772 6400
rect 804 6368 844 6400
rect 876 6368 916 6400
rect 948 6368 1000 6400
rect 0 6328 1000 6368
rect 0 6296 52 6328
rect 84 6296 124 6328
rect 156 6296 196 6328
rect 228 6296 268 6328
rect 300 6296 340 6328
rect 372 6296 412 6328
rect 444 6296 484 6328
rect 516 6296 556 6328
rect 588 6296 628 6328
rect 660 6296 700 6328
rect 732 6296 772 6328
rect 804 6296 844 6328
rect 876 6296 916 6328
rect 948 6296 1000 6328
rect 0 6256 1000 6296
rect 0 6224 52 6256
rect 84 6224 124 6256
rect 156 6224 196 6256
rect 228 6224 268 6256
rect 300 6224 340 6256
rect 372 6224 412 6256
rect 444 6224 484 6256
rect 516 6224 556 6256
rect 588 6224 628 6256
rect 660 6224 700 6256
rect 732 6224 772 6256
rect 804 6224 844 6256
rect 876 6224 916 6256
rect 948 6224 1000 6256
rect 0 6184 1000 6224
rect 0 6152 52 6184
rect 84 6152 124 6184
rect 156 6152 196 6184
rect 228 6152 268 6184
rect 300 6152 340 6184
rect 372 6152 412 6184
rect 444 6152 484 6184
rect 516 6152 556 6184
rect 588 6152 628 6184
rect 660 6152 700 6184
rect 732 6152 772 6184
rect 804 6152 844 6184
rect 876 6152 916 6184
rect 948 6152 1000 6184
rect 0 6112 1000 6152
rect 0 6080 52 6112
rect 84 6080 124 6112
rect 156 6080 196 6112
rect 228 6080 268 6112
rect 300 6080 340 6112
rect 372 6080 412 6112
rect 444 6080 484 6112
rect 516 6080 556 6112
rect 588 6080 628 6112
rect 660 6080 700 6112
rect 732 6080 772 6112
rect 804 6080 844 6112
rect 876 6080 916 6112
rect 948 6080 1000 6112
rect 0 6040 1000 6080
rect 0 6008 52 6040
rect 84 6008 124 6040
rect 156 6008 196 6040
rect 228 6008 268 6040
rect 300 6008 340 6040
rect 372 6008 412 6040
rect 444 6008 484 6040
rect 516 6008 556 6040
rect 588 6008 628 6040
rect 660 6008 700 6040
rect 732 6008 772 6040
rect 804 6008 844 6040
rect 876 6008 916 6040
rect 948 6008 1000 6040
rect 0 5968 1000 6008
rect 0 5936 52 5968
rect 84 5936 124 5968
rect 156 5936 196 5968
rect 228 5936 268 5968
rect 300 5936 340 5968
rect 372 5936 412 5968
rect 444 5936 484 5968
rect 516 5936 556 5968
rect 588 5936 628 5968
rect 660 5936 700 5968
rect 732 5936 772 5968
rect 804 5936 844 5968
rect 876 5936 916 5968
rect 948 5936 1000 5968
rect 0 5896 1000 5936
rect 0 5864 52 5896
rect 84 5864 124 5896
rect 156 5864 196 5896
rect 228 5864 268 5896
rect 300 5864 340 5896
rect 372 5864 412 5896
rect 444 5864 484 5896
rect 516 5864 556 5896
rect 588 5864 628 5896
rect 660 5864 700 5896
rect 732 5864 772 5896
rect 804 5864 844 5896
rect 876 5864 916 5896
rect 948 5864 1000 5896
rect 0 5824 1000 5864
rect 0 5792 52 5824
rect 84 5792 124 5824
rect 156 5792 196 5824
rect 228 5792 268 5824
rect 300 5792 340 5824
rect 372 5792 412 5824
rect 444 5792 484 5824
rect 516 5792 556 5824
rect 588 5792 628 5824
rect 660 5792 700 5824
rect 732 5792 772 5824
rect 804 5792 844 5824
rect 876 5792 916 5824
rect 948 5792 1000 5824
rect 0 5752 1000 5792
rect 0 5720 52 5752
rect 84 5720 124 5752
rect 156 5720 196 5752
rect 228 5720 268 5752
rect 300 5720 340 5752
rect 372 5720 412 5752
rect 444 5720 484 5752
rect 516 5720 556 5752
rect 588 5720 628 5752
rect 660 5720 700 5752
rect 732 5720 772 5752
rect 804 5720 844 5752
rect 876 5720 916 5752
rect 948 5720 1000 5752
rect 0 5680 1000 5720
rect 0 5648 52 5680
rect 84 5648 124 5680
rect 156 5648 196 5680
rect 228 5648 268 5680
rect 300 5648 340 5680
rect 372 5648 412 5680
rect 444 5648 484 5680
rect 516 5648 556 5680
rect 588 5648 628 5680
rect 660 5648 700 5680
rect 732 5648 772 5680
rect 804 5648 844 5680
rect 876 5648 916 5680
rect 948 5648 1000 5680
rect 0 5608 1000 5648
rect 0 5576 52 5608
rect 84 5576 124 5608
rect 156 5576 196 5608
rect 228 5576 268 5608
rect 300 5576 340 5608
rect 372 5576 412 5608
rect 444 5576 484 5608
rect 516 5576 556 5608
rect 588 5576 628 5608
rect 660 5576 700 5608
rect 732 5576 772 5608
rect 804 5576 844 5608
rect 876 5576 916 5608
rect 948 5576 1000 5608
rect 0 5536 1000 5576
rect 0 5504 52 5536
rect 84 5504 124 5536
rect 156 5504 196 5536
rect 228 5504 268 5536
rect 300 5504 340 5536
rect 372 5504 412 5536
rect 444 5504 484 5536
rect 516 5504 556 5536
rect 588 5504 628 5536
rect 660 5504 700 5536
rect 732 5504 772 5536
rect 804 5504 844 5536
rect 876 5504 916 5536
rect 948 5504 1000 5536
rect 0 5464 1000 5504
rect 0 5432 52 5464
rect 84 5432 124 5464
rect 156 5432 196 5464
rect 228 5432 268 5464
rect 300 5432 340 5464
rect 372 5432 412 5464
rect 444 5432 484 5464
rect 516 5432 556 5464
rect 588 5432 628 5464
rect 660 5432 700 5464
rect 732 5432 772 5464
rect 804 5432 844 5464
rect 876 5432 916 5464
rect 948 5432 1000 5464
rect 0 5392 1000 5432
rect 0 5360 52 5392
rect 84 5360 124 5392
rect 156 5360 196 5392
rect 228 5360 268 5392
rect 300 5360 340 5392
rect 372 5360 412 5392
rect 444 5360 484 5392
rect 516 5360 556 5392
rect 588 5360 628 5392
rect 660 5360 700 5392
rect 732 5360 772 5392
rect 804 5360 844 5392
rect 876 5360 916 5392
rect 948 5360 1000 5392
rect 0 5320 1000 5360
rect 0 5288 52 5320
rect 84 5288 124 5320
rect 156 5288 196 5320
rect 228 5288 268 5320
rect 300 5288 340 5320
rect 372 5288 412 5320
rect 444 5288 484 5320
rect 516 5288 556 5320
rect 588 5288 628 5320
rect 660 5288 700 5320
rect 732 5288 772 5320
rect 804 5288 844 5320
rect 876 5288 916 5320
rect 948 5288 1000 5320
rect 0 5248 1000 5288
rect 0 5216 52 5248
rect 84 5216 124 5248
rect 156 5216 196 5248
rect 228 5216 268 5248
rect 300 5216 340 5248
rect 372 5216 412 5248
rect 444 5216 484 5248
rect 516 5216 556 5248
rect 588 5216 628 5248
rect 660 5216 700 5248
rect 732 5216 772 5248
rect 804 5216 844 5248
rect 876 5216 916 5248
rect 948 5216 1000 5248
rect 0 5176 1000 5216
rect 0 5144 52 5176
rect 84 5144 124 5176
rect 156 5144 196 5176
rect 228 5144 268 5176
rect 300 5144 340 5176
rect 372 5144 412 5176
rect 444 5144 484 5176
rect 516 5144 556 5176
rect 588 5144 628 5176
rect 660 5144 700 5176
rect 732 5144 772 5176
rect 804 5144 844 5176
rect 876 5144 916 5176
rect 948 5144 1000 5176
rect 0 5104 1000 5144
rect 0 5072 52 5104
rect 84 5072 124 5104
rect 156 5072 196 5104
rect 228 5072 268 5104
rect 300 5072 340 5104
rect 372 5072 412 5104
rect 444 5072 484 5104
rect 516 5072 556 5104
rect 588 5072 628 5104
rect 660 5072 700 5104
rect 732 5072 772 5104
rect 804 5072 844 5104
rect 876 5072 916 5104
rect 948 5072 1000 5104
rect 0 5032 1000 5072
rect 0 5000 52 5032
rect 84 5000 124 5032
rect 156 5000 196 5032
rect 228 5000 268 5032
rect 300 5000 340 5032
rect 372 5000 412 5032
rect 444 5000 484 5032
rect 516 5000 556 5032
rect 588 5000 628 5032
rect 660 5000 700 5032
rect 732 5000 772 5032
rect 804 5000 844 5032
rect 876 5000 916 5032
rect 948 5000 1000 5032
rect 0 4960 1000 5000
rect 0 4928 52 4960
rect 84 4928 124 4960
rect 156 4928 196 4960
rect 228 4928 268 4960
rect 300 4928 340 4960
rect 372 4928 412 4960
rect 444 4928 484 4960
rect 516 4928 556 4960
rect 588 4928 628 4960
rect 660 4928 700 4960
rect 732 4928 772 4960
rect 804 4928 844 4960
rect 876 4928 916 4960
rect 948 4928 1000 4960
rect 0 4888 1000 4928
rect 0 4856 52 4888
rect 84 4856 124 4888
rect 156 4856 196 4888
rect 228 4856 268 4888
rect 300 4856 340 4888
rect 372 4856 412 4888
rect 444 4856 484 4888
rect 516 4856 556 4888
rect 588 4856 628 4888
rect 660 4856 700 4888
rect 732 4856 772 4888
rect 804 4856 844 4888
rect 876 4856 916 4888
rect 948 4856 1000 4888
rect 0 4816 1000 4856
rect 0 4784 52 4816
rect 84 4784 124 4816
rect 156 4784 196 4816
rect 228 4784 268 4816
rect 300 4784 340 4816
rect 372 4784 412 4816
rect 444 4784 484 4816
rect 516 4784 556 4816
rect 588 4784 628 4816
rect 660 4784 700 4816
rect 732 4784 772 4816
rect 804 4784 844 4816
rect 876 4784 916 4816
rect 948 4784 1000 4816
rect 0 4744 1000 4784
rect 0 4712 52 4744
rect 84 4712 124 4744
rect 156 4712 196 4744
rect 228 4712 268 4744
rect 300 4712 340 4744
rect 372 4712 412 4744
rect 444 4712 484 4744
rect 516 4712 556 4744
rect 588 4712 628 4744
rect 660 4712 700 4744
rect 732 4712 772 4744
rect 804 4712 844 4744
rect 876 4712 916 4744
rect 948 4712 1000 4744
rect 0 4672 1000 4712
rect 0 4640 52 4672
rect 84 4640 124 4672
rect 156 4640 196 4672
rect 228 4640 268 4672
rect 300 4640 340 4672
rect 372 4640 412 4672
rect 444 4640 484 4672
rect 516 4640 556 4672
rect 588 4640 628 4672
rect 660 4640 700 4672
rect 732 4640 772 4672
rect 804 4640 844 4672
rect 876 4640 916 4672
rect 948 4640 1000 4672
rect 0 4600 1000 4640
rect 0 4568 52 4600
rect 84 4568 124 4600
rect 156 4568 196 4600
rect 228 4568 268 4600
rect 300 4568 340 4600
rect 372 4568 412 4600
rect 444 4568 484 4600
rect 516 4568 556 4600
rect 588 4568 628 4600
rect 660 4568 700 4600
rect 732 4568 772 4600
rect 804 4568 844 4600
rect 876 4568 916 4600
rect 948 4568 1000 4600
rect 0 4528 1000 4568
rect 0 4496 52 4528
rect 84 4496 124 4528
rect 156 4496 196 4528
rect 228 4496 268 4528
rect 300 4496 340 4528
rect 372 4496 412 4528
rect 444 4496 484 4528
rect 516 4496 556 4528
rect 588 4496 628 4528
rect 660 4496 700 4528
rect 732 4496 772 4528
rect 804 4496 844 4528
rect 876 4496 916 4528
rect 948 4496 1000 4528
rect 0 4456 1000 4496
rect 0 4424 52 4456
rect 84 4424 124 4456
rect 156 4424 196 4456
rect 228 4424 268 4456
rect 300 4424 340 4456
rect 372 4424 412 4456
rect 444 4424 484 4456
rect 516 4424 556 4456
rect 588 4424 628 4456
rect 660 4424 700 4456
rect 732 4424 772 4456
rect 804 4424 844 4456
rect 876 4424 916 4456
rect 948 4424 1000 4456
rect 0 4384 1000 4424
rect 0 4352 52 4384
rect 84 4352 124 4384
rect 156 4352 196 4384
rect 228 4352 268 4384
rect 300 4352 340 4384
rect 372 4352 412 4384
rect 444 4352 484 4384
rect 516 4352 556 4384
rect 588 4352 628 4384
rect 660 4352 700 4384
rect 732 4352 772 4384
rect 804 4352 844 4384
rect 876 4352 916 4384
rect 948 4352 1000 4384
rect 0 4312 1000 4352
rect 0 4280 52 4312
rect 84 4280 124 4312
rect 156 4280 196 4312
rect 228 4280 268 4312
rect 300 4280 340 4312
rect 372 4280 412 4312
rect 444 4280 484 4312
rect 516 4280 556 4312
rect 588 4280 628 4312
rect 660 4280 700 4312
rect 732 4280 772 4312
rect 804 4280 844 4312
rect 876 4280 916 4312
rect 948 4280 1000 4312
rect 0 4240 1000 4280
rect 0 4208 52 4240
rect 84 4208 124 4240
rect 156 4208 196 4240
rect 228 4208 268 4240
rect 300 4208 340 4240
rect 372 4208 412 4240
rect 444 4208 484 4240
rect 516 4208 556 4240
rect 588 4208 628 4240
rect 660 4208 700 4240
rect 732 4208 772 4240
rect 804 4208 844 4240
rect 876 4208 916 4240
rect 948 4208 1000 4240
rect 0 4168 1000 4208
rect 0 4136 52 4168
rect 84 4136 124 4168
rect 156 4136 196 4168
rect 228 4136 268 4168
rect 300 4136 340 4168
rect 372 4136 412 4168
rect 444 4136 484 4168
rect 516 4136 556 4168
rect 588 4136 628 4168
rect 660 4136 700 4168
rect 732 4136 772 4168
rect 804 4136 844 4168
rect 876 4136 916 4168
rect 948 4136 1000 4168
rect 0 4096 1000 4136
rect 0 4064 52 4096
rect 84 4064 124 4096
rect 156 4064 196 4096
rect 228 4064 268 4096
rect 300 4064 340 4096
rect 372 4064 412 4096
rect 444 4064 484 4096
rect 516 4064 556 4096
rect 588 4064 628 4096
rect 660 4064 700 4096
rect 732 4064 772 4096
rect 804 4064 844 4096
rect 876 4064 916 4096
rect 948 4064 1000 4096
rect 0 4024 1000 4064
rect 0 3992 52 4024
rect 84 3992 124 4024
rect 156 3992 196 4024
rect 228 3992 268 4024
rect 300 3992 340 4024
rect 372 3992 412 4024
rect 444 3992 484 4024
rect 516 3992 556 4024
rect 588 3992 628 4024
rect 660 3992 700 4024
rect 732 3992 772 4024
rect 804 3992 844 4024
rect 876 3992 916 4024
rect 948 3992 1000 4024
rect 0 3952 1000 3992
rect 0 3920 52 3952
rect 84 3920 124 3952
rect 156 3920 196 3952
rect 228 3920 268 3952
rect 300 3920 340 3952
rect 372 3920 412 3952
rect 444 3920 484 3952
rect 516 3920 556 3952
rect 588 3920 628 3952
rect 660 3920 700 3952
rect 732 3920 772 3952
rect 804 3920 844 3952
rect 876 3920 916 3952
rect 948 3920 1000 3952
rect 0 3880 1000 3920
rect 0 3848 52 3880
rect 84 3848 124 3880
rect 156 3848 196 3880
rect 228 3848 268 3880
rect 300 3848 340 3880
rect 372 3848 412 3880
rect 444 3848 484 3880
rect 516 3848 556 3880
rect 588 3848 628 3880
rect 660 3848 700 3880
rect 732 3848 772 3880
rect 804 3848 844 3880
rect 876 3848 916 3880
rect 948 3848 1000 3880
rect 0 3808 1000 3848
rect 0 3776 52 3808
rect 84 3776 124 3808
rect 156 3776 196 3808
rect 228 3776 268 3808
rect 300 3776 340 3808
rect 372 3776 412 3808
rect 444 3776 484 3808
rect 516 3776 556 3808
rect 588 3776 628 3808
rect 660 3776 700 3808
rect 732 3776 772 3808
rect 804 3776 844 3808
rect 876 3776 916 3808
rect 948 3776 1000 3808
rect 0 3736 1000 3776
rect 0 3704 52 3736
rect 84 3704 124 3736
rect 156 3704 196 3736
rect 228 3704 268 3736
rect 300 3704 340 3736
rect 372 3704 412 3736
rect 444 3704 484 3736
rect 516 3704 556 3736
rect 588 3704 628 3736
rect 660 3704 700 3736
rect 732 3704 772 3736
rect 804 3704 844 3736
rect 876 3704 916 3736
rect 948 3704 1000 3736
rect 0 3664 1000 3704
rect 0 3632 52 3664
rect 84 3632 124 3664
rect 156 3632 196 3664
rect 228 3632 268 3664
rect 300 3632 340 3664
rect 372 3632 412 3664
rect 444 3632 484 3664
rect 516 3632 556 3664
rect 588 3632 628 3664
rect 660 3632 700 3664
rect 732 3632 772 3664
rect 804 3632 844 3664
rect 876 3632 916 3664
rect 948 3632 1000 3664
rect 0 3592 1000 3632
rect 0 3560 52 3592
rect 84 3560 124 3592
rect 156 3560 196 3592
rect 228 3560 268 3592
rect 300 3560 340 3592
rect 372 3560 412 3592
rect 444 3560 484 3592
rect 516 3560 556 3592
rect 588 3560 628 3592
rect 660 3560 700 3592
rect 732 3560 772 3592
rect 804 3560 844 3592
rect 876 3560 916 3592
rect 948 3560 1000 3592
rect 0 3520 1000 3560
rect 0 3488 52 3520
rect 84 3488 124 3520
rect 156 3488 196 3520
rect 228 3488 268 3520
rect 300 3488 340 3520
rect 372 3488 412 3520
rect 444 3488 484 3520
rect 516 3488 556 3520
rect 588 3488 628 3520
rect 660 3488 700 3520
rect 732 3488 772 3520
rect 804 3488 844 3520
rect 876 3488 916 3520
rect 948 3488 1000 3520
rect 0 3448 1000 3488
rect 0 3416 52 3448
rect 84 3416 124 3448
rect 156 3416 196 3448
rect 228 3416 268 3448
rect 300 3416 340 3448
rect 372 3416 412 3448
rect 444 3416 484 3448
rect 516 3416 556 3448
rect 588 3416 628 3448
rect 660 3416 700 3448
rect 732 3416 772 3448
rect 804 3416 844 3448
rect 876 3416 916 3448
rect 948 3416 1000 3448
rect 0 3376 1000 3416
rect 0 3344 52 3376
rect 84 3344 124 3376
rect 156 3344 196 3376
rect 228 3344 268 3376
rect 300 3344 340 3376
rect 372 3344 412 3376
rect 444 3344 484 3376
rect 516 3344 556 3376
rect 588 3344 628 3376
rect 660 3344 700 3376
rect 732 3344 772 3376
rect 804 3344 844 3376
rect 876 3344 916 3376
rect 948 3344 1000 3376
rect 0 3304 1000 3344
rect 0 3272 52 3304
rect 84 3272 124 3304
rect 156 3272 196 3304
rect 228 3272 268 3304
rect 300 3272 340 3304
rect 372 3272 412 3304
rect 444 3272 484 3304
rect 516 3272 556 3304
rect 588 3272 628 3304
rect 660 3272 700 3304
rect 732 3272 772 3304
rect 804 3272 844 3304
rect 876 3272 916 3304
rect 948 3272 1000 3304
rect 0 3232 1000 3272
rect 0 3200 52 3232
rect 84 3200 124 3232
rect 156 3200 196 3232
rect 228 3200 268 3232
rect 300 3200 340 3232
rect 372 3200 412 3232
rect 444 3200 484 3232
rect 516 3200 556 3232
rect 588 3200 628 3232
rect 660 3200 700 3232
rect 732 3200 772 3232
rect 804 3200 844 3232
rect 876 3200 916 3232
rect 948 3200 1000 3232
rect 0 3160 1000 3200
rect 0 3128 52 3160
rect 84 3128 124 3160
rect 156 3128 196 3160
rect 228 3128 268 3160
rect 300 3128 340 3160
rect 372 3128 412 3160
rect 444 3128 484 3160
rect 516 3128 556 3160
rect 588 3128 628 3160
rect 660 3128 700 3160
rect 732 3128 772 3160
rect 804 3128 844 3160
rect 876 3128 916 3160
rect 948 3128 1000 3160
rect 0 3088 1000 3128
rect 0 3056 52 3088
rect 84 3056 124 3088
rect 156 3056 196 3088
rect 228 3056 268 3088
rect 300 3056 340 3088
rect 372 3056 412 3088
rect 444 3056 484 3088
rect 516 3056 556 3088
rect 588 3056 628 3088
rect 660 3056 700 3088
rect 732 3056 772 3088
rect 804 3056 844 3088
rect 876 3056 916 3088
rect 948 3056 1000 3088
rect 0 3016 1000 3056
rect 0 2984 52 3016
rect 84 2984 124 3016
rect 156 2984 196 3016
rect 228 2984 268 3016
rect 300 2984 340 3016
rect 372 2984 412 3016
rect 444 2984 484 3016
rect 516 2984 556 3016
rect 588 2984 628 3016
rect 660 2984 700 3016
rect 732 2984 772 3016
rect 804 2984 844 3016
rect 876 2984 916 3016
rect 948 2984 1000 3016
rect 0 2944 1000 2984
rect 0 2912 52 2944
rect 84 2912 124 2944
rect 156 2912 196 2944
rect 228 2912 268 2944
rect 300 2912 340 2944
rect 372 2912 412 2944
rect 444 2912 484 2944
rect 516 2912 556 2944
rect 588 2912 628 2944
rect 660 2912 700 2944
rect 732 2912 772 2944
rect 804 2912 844 2944
rect 876 2912 916 2944
rect 948 2912 1000 2944
rect 0 2872 1000 2912
rect 0 2840 52 2872
rect 84 2840 124 2872
rect 156 2840 196 2872
rect 228 2840 268 2872
rect 300 2840 340 2872
rect 372 2840 412 2872
rect 444 2840 484 2872
rect 516 2840 556 2872
rect 588 2840 628 2872
rect 660 2840 700 2872
rect 732 2840 772 2872
rect 804 2840 844 2872
rect 876 2840 916 2872
rect 948 2840 1000 2872
rect 0 2800 1000 2840
rect 0 2768 52 2800
rect 84 2768 124 2800
rect 156 2768 196 2800
rect 228 2768 268 2800
rect 300 2768 340 2800
rect 372 2768 412 2800
rect 444 2768 484 2800
rect 516 2768 556 2800
rect 588 2768 628 2800
rect 660 2768 700 2800
rect 732 2768 772 2800
rect 804 2768 844 2800
rect 876 2768 916 2800
rect 948 2768 1000 2800
rect 0 2728 1000 2768
rect 0 2696 52 2728
rect 84 2696 124 2728
rect 156 2696 196 2728
rect 228 2696 268 2728
rect 300 2696 340 2728
rect 372 2696 412 2728
rect 444 2696 484 2728
rect 516 2696 556 2728
rect 588 2696 628 2728
rect 660 2696 700 2728
rect 732 2696 772 2728
rect 804 2696 844 2728
rect 876 2696 916 2728
rect 948 2696 1000 2728
rect 0 2656 1000 2696
rect 0 2624 52 2656
rect 84 2624 124 2656
rect 156 2624 196 2656
rect 228 2624 268 2656
rect 300 2624 340 2656
rect 372 2624 412 2656
rect 444 2624 484 2656
rect 516 2624 556 2656
rect 588 2624 628 2656
rect 660 2624 700 2656
rect 732 2624 772 2656
rect 804 2624 844 2656
rect 876 2624 916 2656
rect 948 2624 1000 2656
rect 0 2584 1000 2624
rect 0 2552 52 2584
rect 84 2552 124 2584
rect 156 2552 196 2584
rect 228 2552 268 2584
rect 300 2552 340 2584
rect 372 2552 412 2584
rect 444 2552 484 2584
rect 516 2552 556 2584
rect 588 2552 628 2584
rect 660 2552 700 2584
rect 732 2552 772 2584
rect 804 2552 844 2584
rect 876 2552 916 2584
rect 948 2552 1000 2584
rect 0 2512 1000 2552
rect 0 2480 52 2512
rect 84 2480 124 2512
rect 156 2480 196 2512
rect 228 2480 268 2512
rect 300 2480 340 2512
rect 372 2480 412 2512
rect 444 2480 484 2512
rect 516 2480 556 2512
rect 588 2480 628 2512
rect 660 2480 700 2512
rect 732 2480 772 2512
rect 804 2480 844 2512
rect 876 2480 916 2512
rect 948 2480 1000 2512
rect 0 2440 1000 2480
rect 0 2408 52 2440
rect 84 2408 124 2440
rect 156 2408 196 2440
rect 228 2408 268 2440
rect 300 2408 340 2440
rect 372 2408 412 2440
rect 444 2408 484 2440
rect 516 2408 556 2440
rect 588 2408 628 2440
rect 660 2408 700 2440
rect 732 2408 772 2440
rect 804 2408 844 2440
rect 876 2408 916 2440
rect 948 2408 1000 2440
rect 0 2368 1000 2408
rect 0 2336 52 2368
rect 84 2336 124 2368
rect 156 2336 196 2368
rect 228 2336 268 2368
rect 300 2336 340 2368
rect 372 2336 412 2368
rect 444 2336 484 2368
rect 516 2336 556 2368
rect 588 2336 628 2368
rect 660 2336 700 2368
rect 732 2336 772 2368
rect 804 2336 844 2368
rect 876 2336 916 2368
rect 948 2336 1000 2368
rect 0 2296 1000 2336
rect 0 2264 52 2296
rect 84 2264 124 2296
rect 156 2264 196 2296
rect 228 2264 268 2296
rect 300 2264 340 2296
rect 372 2264 412 2296
rect 444 2264 484 2296
rect 516 2264 556 2296
rect 588 2264 628 2296
rect 660 2264 700 2296
rect 732 2264 772 2296
rect 804 2264 844 2296
rect 876 2264 916 2296
rect 948 2264 1000 2296
rect 0 2224 1000 2264
rect 0 2192 52 2224
rect 84 2192 124 2224
rect 156 2192 196 2224
rect 228 2192 268 2224
rect 300 2192 340 2224
rect 372 2192 412 2224
rect 444 2192 484 2224
rect 516 2192 556 2224
rect 588 2192 628 2224
rect 660 2192 700 2224
rect 732 2192 772 2224
rect 804 2192 844 2224
rect 876 2192 916 2224
rect 948 2192 1000 2224
rect 0 2152 1000 2192
rect 0 2120 52 2152
rect 84 2120 124 2152
rect 156 2120 196 2152
rect 228 2120 268 2152
rect 300 2120 340 2152
rect 372 2120 412 2152
rect 444 2120 484 2152
rect 516 2120 556 2152
rect 588 2120 628 2152
rect 660 2120 700 2152
rect 732 2120 772 2152
rect 804 2120 844 2152
rect 876 2120 916 2152
rect 948 2120 1000 2152
rect 0 2080 1000 2120
rect 0 2048 52 2080
rect 84 2048 124 2080
rect 156 2048 196 2080
rect 228 2048 268 2080
rect 300 2048 340 2080
rect 372 2048 412 2080
rect 444 2048 484 2080
rect 516 2048 556 2080
rect 588 2048 628 2080
rect 660 2048 700 2080
rect 732 2048 772 2080
rect 804 2048 844 2080
rect 876 2048 916 2080
rect 948 2048 1000 2080
rect 0 2008 1000 2048
rect 0 1976 52 2008
rect 84 1976 124 2008
rect 156 1976 196 2008
rect 228 1976 268 2008
rect 300 1976 340 2008
rect 372 1976 412 2008
rect 444 1976 484 2008
rect 516 1976 556 2008
rect 588 1976 628 2008
rect 660 1976 700 2008
rect 732 1976 772 2008
rect 804 1976 844 2008
rect 876 1976 916 2008
rect 948 1976 1000 2008
rect 0 1936 1000 1976
rect 0 1904 52 1936
rect 84 1904 124 1936
rect 156 1904 196 1936
rect 228 1904 268 1936
rect 300 1904 340 1936
rect 372 1904 412 1936
rect 444 1904 484 1936
rect 516 1904 556 1936
rect 588 1904 628 1936
rect 660 1904 700 1936
rect 732 1904 772 1936
rect 804 1904 844 1936
rect 876 1904 916 1936
rect 948 1904 1000 1936
rect 0 1864 1000 1904
rect 0 1832 52 1864
rect 84 1832 124 1864
rect 156 1832 196 1864
rect 228 1832 268 1864
rect 300 1832 340 1864
rect 372 1832 412 1864
rect 444 1832 484 1864
rect 516 1832 556 1864
rect 588 1832 628 1864
rect 660 1832 700 1864
rect 732 1832 772 1864
rect 804 1832 844 1864
rect 876 1832 916 1864
rect 948 1832 1000 1864
rect 0 1792 1000 1832
rect 0 1760 52 1792
rect 84 1760 124 1792
rect 156 1760 196 1792
rect 228 1760 268 1792
rect 300 1760 340 1792
rect 372 1760 412 1792
rect 444 1760 484 1792
rect 516 1760 556 1792
rect 588 1760 628 1792
rect 660 1760 700 1792
rect 732 1760 772 1792
rect 804 1760 844 1792
rect 876 1760 916 1792
rect 948 1760 1000 1792
rect 0 1720 1000 1760
rect 0 1688 52 1720
rect 84 1688 124 1720
rect 156 1688 196 1720
rect 228 1688 268 1720
rect 300 1688 340 1720
rect 372 1688 412 1720
rect 444 1688 484 1720
rect 516 1688 556 1720
rect 588 1688 628 1720
rect 660 1688 700 1720
rect 732 1688 772 1720
rect 804 1688 844 1720
rect 876 1688 916 1720
rect 948 1688 1000 1720
rect 0 1648 1000 1688
rect 0 1616 52 1648
rect 84 1616 124 1648
rect 156 1616 196 1648
rect 228 1616 268 1648
rect 300 1616 340 1648
rect 372 1616 412 1648
rect 444 1616 484 1648
rect 516 1616 556 1648
rect 588 1616 628 1648
rect 660 1616 700 1648
rect 732 1616 772 1648
rect 804 1616 844 1648
rect 876 1616 916 1648
rect 948 1616 1000 1648
rect 0 1576 1000 1616
rect 0 1544 52 1576
rect 84 1544 124 1576
rect 156 1544 196 1576
rect 228 1544 268 1576
rect 300 1544 340 1576
rect 372 1544 412 1576
rect 444 1544 484 1576
rect 516 1544 556 1576
rect 588 1544 628 1576
rect 660 1544 700 1576
rect 732 1544 772 1576
rect 804 1544 844 1576
rect 876 1544 916 1576
rect 948 1544 1000 1576
rect 0 1504 1000 1544
rect 0 1472 52 1504
rect 84 1472 124 1504
rect 156 1472 196 1504
rect 228 1472 268 1504
rect 300 1472 340 1504
rect 372 1472 412 1504
rect 444 1472 484 1504
rect 516 1472 556 1504
rect 588 1472 628 1504
rect 660 1472 700 1504
rect 732 1472 772 1504
rect 804 1472 844 1504
rect 876 1472 916 1504
rect 948 1472 1000 1504
rect 0 1432 1000 1472
rect 0 1400 52 1432
rect 84 1400 124 1432
rect 156 1400 196 1432
rect 228 1400 268 1432
rect 300 1400 340 1432
rect 372 1400 412 1432
rect 444 1400 484 1432
rect 516 1400 556 1432
rect 588 1400 628 1432
rect 660 1400 700 1432
rect 732 1400 772 1432
rect 804 1400 844 1432
rect 876 1400 916 1432
rect 948 1400 1000 1432
rect 0 1360 1000 1400
rect 0 1328 52 1360
rect 84 1328 124 1360
rect 156 1328 196 1360
rect 228 1328 268 1360
rect 300 1328 340 1360
rect 372 1328 412 1360
rect 444 1328 484 1360
rect 516 1328 556 1360
rect 588 1328 628 1360
rect 660 1328 700 1360
rect 732 1328 772 1360
rect 804 1328 844 1360
rect 876 1328 916 1360
rect 948 1328 1000 1360
rect 0 1288 1000 1328
rect 0 1256 52 1288
rect 84 1256 124 1288
rect 156 1256 196 1288
rect 228 1256 268 1288
rect 300 1256 340 1288
rect 372 1256 412 1288
rect 444 1256 484 1288
rect 516 1256 556 1288
rect 588 1256 628 1288
rect 660 1256 700 1288
rect 732 1256 772 1288
rect 804 1256 844 1288
rect 876 1256 916 1288
rect 948 1256 1000 1288
rect 0 1200 1000 1256
<< metal3 >>
rect 0 32000 1000 35600
rect 0 28000 1000 31600
rect 0 25200 1000 26800
rect 0 18700 1000 23800
rect 0 13200 1000 18300
rect 0 6900 1000 12000
rect 0 1400 1000 6500
<< metal4 >>
rect 0 32440 1000 35600
rect 0 28000 1000 31160
rect 0 25200 1000 26800
rect 0 18700 1000 23800
rect 0 13200 1000 18300
rect 0 6900 1000 12000
rect 0 1400 1000 6500
<< metal5 >>
rect 0 32000 1000 35600
rect 0 28000 1000 31600
rect 0 25200 1000 26800
rect 0 18700 1000 23800
rect 0 13200 1000 18300
rect 0 6900 1000 12000
rect 0 1400 1000 6500
<< metal6 >>
rect 0 32000 1000 35600
rect 0 28000 1000 31600
rect 0 25200 1000 26800
rect 0 18700 1000 23800
rect 0 13200 1000 18300
rect 0 6900 1000 12000
rect 0 1400 1000 6500
<< metal7 >>
rect 0 25500 1000 26500
rect 0 19000 1000 23500
rect 0 13500 1000 18000
rect 0 7200 1000 11700
rect 0 1700 1000 6200
<< labels >>
rlabel metal3 s 0 32000 1000 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 1000 31600 4 vss
port 1 nsew
rlabel metal3 s 0 18700 1000 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 13200 1000 18300 4 iovdd
port 4 nsew
rlabel metal3 s 0 25200 1000 26800 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 1000 6500 4 iovss
port 3 nsew
rlabel metal3 s 0 6900 1000 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 1000 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 1000 35600 4 vss
port 1 nsew
rlabel metal4 s 0 18700 1000 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 13200 1000 18300 4 iovdd
port 4 nsew
rlabel metal4 s 0 25200 1000 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 1000 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 6900 1000 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 1000 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 1000 35600 4 vss
port 1 nsew
rlabel metal5 s 0 18700 1000 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 13200 1000 18300 4 iovdd
port 4 nsew
rlabel metal5 s 0 25200 1000 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 1000 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 6900 1000 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 1000 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 1000 35600 4 vss
port 1 nsew
rlabel metal6 s 0 18700 1000 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 13200 1000 18300 4 iovdd
port 4 nsew
rlabel metal6 s 0 25200 1000 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 1000 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 6900 1000 12000 4 iovss
port 3 nsew
rlabel metal7 s 0 13500 1000 18000 4 iovdd
port 4 nsew
rlabel metal7 s 0 19000 1000 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 1700 1000 6200 4 iovss
port 3 nsew
rlabel metal7 s 0 7200 1000 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 25500 1000 26500 4 iovss
port 3 nsew
flabel comment s 212 17744 212 17744 0 FreeSans 400 0 0 0 sub!
flabel comment s 219 22802 219 22802 0 FreeSans 400 0 0 0 sub!
flabel comment s 225 27708 225 27708 0 FreeSans 400 0 0 0 sub!
flabel comment s 534 31400 534 31400 0 FreeSans 400 0 0 0 sub!
flabel metal1 s 420 6226 622 6405 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 374 7940 588 8102 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 124 17524 268 17586 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 124 22628 268 22690 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 124 27517 268 27579 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 183 31384 273 31416 0 FreeSans 400 0 0 0 vss
port 1 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 1000 36000
string GDS_END 63852602
string GDS_FILE sg13g2_io.gds
string GDS_START 63578298
<< end >>
