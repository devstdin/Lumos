magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2124 18124 7008
<< nwell >>
rect -124 4692 16124 5008
rect -124 192 192 4692
rect 15808 192 16124 4692
rect -124 -124 16124 192
<< pwell >>
rect 334 4430 15666 4550
rect 334 454 454 4430
rect 880 4122 1028 4430
rect 1451 454 14549 4430
rect 15546 454 15666 4430
rect 334 334 15666 454
<< hvnmos >>
rect 1571 3454 1691 4334
rect 1927 3454 2047 4334
rect 2175 3454 2295 4334
rect 2531 3454 2651 4334
rect 2779 3454 2899 4334
rect 3135 3454 3255 4334
rect 3383 3454 3503 4334
rect 3739 3454 3859 4334
rect 3987 3454 4107 4334
rect 4343 3454 4463 4334
rect 4591 3454 4711 4334
rect 4947 3454 5067 4334
rect 5195 3454 5315 4334
rect 5551 3454 5671 4334
rect 5799 3454 5919 4334
rect 6155 3454 6275 4334
rect 6403 3454 6523 4334
rect 6759 3454 6879 4334
rect 7007 3454 7127 4334
rect 7363 3454 7483 4334
rect 7611 3454 7731 4334
rect 7967 3454 8087 4334
rect 8215 3454 8335 4334
rect 8571 3454 8691 4334
rect 8819 3454 8939 4334
rect 9175 3454 9295 4334
rect 9423 3454 9543 4334
rect 9779 3454 9899 4334
rect 10027 3454 10147 4334
rect 10383 3454 10503 4334
rect 10631 3454 10751 4334
rect 10987 3454 11107 4334
rect 11235 3454 11355 4334
rect 11591 3454 11711 4334
rect 11839 3454 11959 4334
rect 12195 3454 12315 4334
rect 12443 3454 12563 4334
rect 12799 3454 12919 4334
rect 13047 3454 13167 4334
rect 13403 3454 13523 4334
rect 13651 3454 13771 4334
rect 14007 3454 14127 4334
rect 14255 3454 14375 4334
rect 1571 2486 1691 3366
rect 1927 2486 2047 3366
rect 2175 2486 2295 3366
rect 2531 2486 2651 3366
rect 2779 2486 2899 3366
rect 3135 2486 3255 3366
rect 3383 2486 3503 3366
rect 3739 2486 3859 3366
rect 3987 2486 4107 3366
rect 4343 2486 4463 3366
rect 4591 2486 4711 3366
rect 4947 2486 5067 3366
rect 5195 2486 5315 3366
rect 5551 2486 5671 3366
rect 5799 2486 5919 3366
rect 6155 2486 6275 3366
rect 6403 2486 6523 3366
rect 6759 2486 6879 3366
rect 7007 2486 7127 3366
rect 7363 2486 7483 3366
rect 7611 2486 7731 3366
rect 7967 2486 8087 3366
rect 8215 2486 8335 3366
rect 8571 2486 8691 3366
rect 8819 2486 8939 3366
rect 9175 2486 9295 3366
rect 9423 2486 9543 3366
rect 9779 2486 9899 3366
rect 10027 2486 10147 3366
rect 10383 2486 10503 3366
rect 10631 2486 10751 3366
rect 10987 2486 11107 3366
rect 11235 2486 11355 3366
rect 11591 2486 11711 3366
rect 11839 2486 11959 3366
rect 12195 2486 12315 3366
rect 12443 2486 12563 3366
rect 12799 2486 12919 3366
rect 13047 2486 13167 3366
rect 13403 2486 13523 3366
rect 13651 2486 13771 3366
rect 14007 2486 14127 3366
rect 14255 2486 14375 3366
rect 1571 1518 1691 2398
rect 1927 1518 2047 2398
rect 2175 1518 2295 2398
rect 2531 1518 2651 2398
rect 2779 1518 2899 2398
rect 3135 1518 3255 2398
rect 3383 1518 3503 2398
rect 3739 1518 3859 2398
rect 3987 1518 4107 2398
rect 4343 1518 4463 2398
rect 4591 1518 4711 2398
rect 4947 1518 5067 2398
rect 5195 1518 5315 2398
rect 5551 1518 5671 2398
rect 5799 1518 5919 2398
rect 6155 1518 6275 2398
rect 6403 1518 6523 2398
rect 6759 1518 6879 2398
rect 7007 1518 7127 2398
rect 7363 1518 7483 2398
rect 7611 1518 7731 2398
rect 7967 1518 8087 2398
rect 8215 1518 8335 2398
rect 8571 1518 8691 2398
rect 8819 1518 8939 2398
rect 9175 1518 9295 2398
rect 9423 1518 9543 2398
rect 9779 1518 9899 2398
rect 10027 1518 10147 2398
rect 10383 1518 10503 2398
rect 10631 1518 10751 2398
rect 10987 1518 11107 2398
rect 11235 1518 11355 2398
rect 11591 1518 11711 2398
rect 11839 1518 11959 2398
rect 12195 1518 12315 2398
rect 12443 1518 12563 2398
rect 12799 1518 12919 2398
rect 13047 1518 13167 2398
rect 13403 1518 13523 2398
rect 13651 1518 13771 2398
rect 14007 1518 14127 2398
rect 14255 1518 14375 2398
rect 1571 550 1691 1430
rect 1927 550 2047 1430
rect 2175 550 2295 1430
rect 2531 550 2651 1430
rect 2779 550 2899 1430
rect 3135 550 3255 1430
rect 3383 550 3503 1430
rect 3739 550 3859 1430
rect 3987 550 4107 1430
rect 4343 550 4463 1430
rect 4591 550 4711 1430
rect 4947 550 5067 1430
rect 5195 550 5315 1430
rect 5551 550 5671 1430
rect 5799 550 5919 1430
rect 6155 550 6275 1430
rect 6403 550 6523 1430
rect 6759 550 6879 1430
rect 7007 550 7127 1430
rect 7363 550 7483 1430
rect 7611 550 7731 1430
rect 7967 550 8087 1430
rect 8215 550 8335 1430
rect 8571 550 8691 1430
rect 8819 550 8939 1430
rect 9175 550 9295 1430
rect 9423 550 9543 1430
rect 9779 550 9899 1430
rect 10027 550 10147 1430
rect 10383 550 10503 1430
rect 10631 550 10751 1430
rect 10987 550 11107 1430
rect 11235 550 11355 1430
rect 11591 550 11711 1430
rect 11839 550 11959 1430
rect 12195 550 12315 1430
rect 12443 550 12563 1430
rect 12799 550 12919 1430
rect 13047 550 13167 1430
rect 13403 550 13523 1430
rect 13651 550 13771 1430
rect 14007 550 14127 1430
rect 14255 550 14375 1430
<< hvndiff >>
rect 1477 4318 1571 4334
rect 1477 4286 1491 4318
rect 1523 4286 1571 4318
rect 1477 4250 1571 4286
rect 1477 4218 1491 4250
rect 1523 4218 1571 4250
rect 1477 4182 1571 4218
rect 1477 4150 1491 4182
rect 1523 4150 1571 4182
rect 1477 4114 1571 4150
rect 1477 4082 1491 4114
rect 1523 4082 1571 4114
rect 1477 4046 1571 4082
rect 1477 4014 1491 4046
rect 1523 4014 1571 4046
rect 1477 3978 1571 4014
rect 1477 3946 1491 3978
rect 1523 3946 1571 3978
rect 1477 3910 1571 3946
rect 1477 3878 1491 3910
rect 1523 3878 1571 3910
rect 1477 3842 1571 3878
rect 1477 3810 1491 3842
rect 1523 3810 1571 3842
rect 1477 3774 1571 3810
rect 1477 3742 1491 3774
rect 1523 3742 1571 3774
rect 1477 3706 1571 3742
rect 1477 3674 1491 3706
rect 1523 3674 1571 3706
rect 1477 3638 1571 3674
rect 1477 3606 1491 3638
rect 1523 3606 1571 3638
rect 1477 3570 1571 3606
rect 1477 3538 1491 3570
rect 1523 3538 1571 3570
rect 1477 3502 1571 3538
rect 1477 3470 1491 3502
rect 1523 3470 1571 3502
rect 1477 3454 1571 3470
rect 1691 4318 1927 4334
rect 1691 4286 1793 4318
rect 1825 4286 1927 4318
rect 1691 4250 1927 4286
rect 1691 4218 1793 4250
rect 1825 4218 1927 4250
rect 1691 4182 1927 4218
rect 1691 4150 1793 4182
rect 1825 4150 1927 4182
rect 1691 4114 1927 4150
rect 1691 4082 1793 4114
rect 1825 4082 1927 4114
rect 1691 4046 1927 4082
rect 1691 4014 1793 4046
rect 1825 4014 1927 4046
rect 1691 3978 1927 4014
rect 1691 3946 1793 3978
rect 1825 3946 1927 3978
rect 1691 3910 1927 3946
rect 1691 3878 1793 3910
rect 1825 3878 1927 3910
rect 1691 3842 1927 3878
rect 1691 3810 1793 3842
rect 1825 3810 1927 3842
rect 1691 3774 1927 3810
rect 1691 3742 1793 3774
rect 1825 3742 1927 3774
rect 1691 3706 1927 3742
rect 1691 3674 1793 3706
rect 1825 3674 1927 3706
rect 1691 3638 1927 3674
rect 1691 3606 1793 3638
rect 1825 3606 1927 3638
rect 1691 3570 1927 3606
rect 1691 3538 1793 3570
rect 1825 3538 1927 3570
rect 1691 3502 1927 3538
rect 1691 3470 1793 3502
rect 1825 3470 1927 3502
rect 1691 3454 1927 3470
rect 2047 4318 2175 4334
rect 2047 4286 2095 4318
rect 2127 4286 2175 4318
rect 2047 4250 2175 4286
rect 2047 4218 2095 4250
rect 2127 4218 2175 4250
rect 2047 4182 2175 4218
rect 2047 4150 2095 4182
rect 2127 4150 2175 4182
rect 2047 4114 2175 4150
rect 2047 4082 2095 4114
rect 2127 4082 2175 4114
rect 2047 4046 2175 4082
rect 2047 4014 2095 4046
rect 2127 4014 2175 4046
rect 2047 3978 2175 4014
rect 2047 3946 2095 3978
rect 2127 3946 2175 3978
rect 2047 3910 2175 3946
rect 2047 3878 2095 3910
rect 2127 3878 2175 3910
rect 2047 3842 2175 3878
rect 2047 3810 2095 3842
rect 2127 3810 2175 3842
rect 2047 3774 2175 3810
rect 2047 3742 2095 3774
rect 2127 3742 2175 3774
rect 2047 3706 2175 3742
rect 2047 3674 2095 3706
rect 2127 3674 2175 3706
rect 2047 3638 2175 3674
rect 2047 3606 2095 3638
rect 2127 3606 2175 3638
rect 2047 3570 2175 3606
rect 2047 3538 2095 3570
rect 2127 3538 2175 3570
rect 2047 3502 2175 3538
rect 2047 3470 2095 3502
rect 2127 3470 2175 3502
rect 2047 3454 2175 3470
rect 2295 4318 2531 4334
rect 2295 4286 2397 4318
rect 2429 4286 2531 4318
rect 2295 4250 2531 4286
rect 2295 4218 2397 4250
rect 2429 4218 2531 4250
rect 2295 4182 2531 4218
rect 2295 4150 2397 4182
rect 2429 4150 2531 4182
rect 2295 4114 2531 4150
rect 2295 4082 2397 4114
rect 2429 4082 2531 4114
rect 2295 4046 2531 4082
rect 2295 4014 2397 4046
rect 2429 4014 2531 4046
rect 2295 3978 2531 4014
rect 2295 3946 2397 3978
rect 2429 3946 2531 3978
rect 2295 3910 2531 3946
rect 2295 3878 2397 3910
rect 2429 3878 2531 3910
rect 2295 3842 2531 3878
rect 2295 3810 2397 3842
rect 2429 3810 2531 3842
rect 2295 3774 2531 3810
rect 2295 3742 2397 3774
rect 2429 3742 2531 3774
rect 2295 3706 2531 3742
rect 2295 3674 2397 3706
rect 2429 3674 2531 3706
rect 2295 3638 2531 3674
rect 2295 3606 2397 3638
rect 2429 3606 2531 3638
rect 2295 3570 2531 3606
rect 2295 3538 2397 3570
rect 2429 3538 2531 3570
rect 2295 3502 2531 3538
rect 2295 3470 2397 3502
rect 2429 3470 2531 3502
rect 2295 3454 2531 3470
rect 2651 4318 2779 4334
rect 2651 4286 2699 4318
rect 2731 4286 2779 4318
rect 2651 4250 2779 4286
rect 2651 4218 2699 4250
rect 2731 4218 2779 4250
rect 2651 4182 2779 4218
rect 2651 4150 2699 4182
rect 2731 4150 2779 4182
rect 2651 4114 2779 4150
rect 2651 4082 2699 4114
rect 2731 4082 2779 4114
rect 2651 4046 2779 4082
rect 2651 4014 2699 4046
rect 2731 4014 2779 4046
rect 2651 3978 2779 4014
rect 2651 3946 2699 3978
rect 2731 3946 2779 3978
rect 2651 3910 2779 3946
rect 2651 3878 2699 3910
rect 2731 3878 2779 3910
rect 2651 3842 2779 3878
rect 2651 3810 2699 3842
rect 2731 3810 2779 3842
rect 2651 3774 2779 3810
rect 2651 3742 2699 3774
rect 2731 3742 2779 3774
rect 2651 3706 2779 3742
rect 2651 3674 2699 3706
rect 2731 3674 2779 3706
rect 2651 3638 2779 3674
rect 2651 3606 2699 3638
rect 2731 3606 2779 3638
rect 2651 3570 2779 3606
rect 2651 3538 2699 3570
rect 2731 3538 2779 3570
rect 2651 3502 2779 3538
rect 2651 3470 2699 3502
rect 2731 3470 2779 3502
rect 2651 3454 2779 3470
rect 2899 4318 3135 4334
rect 2899 4286 3001 4318
rect 3033 4286 3135 4318
rect 2899 4250 3135 4286
rect 2899 4218 3001 4250
rect 3033 4218 3135 4250
rect 2899 4182 3135 4218
rect 2899 4150 3001 4182
rect 3033 4150 3135 4182
rect 2899 4114 3135 4150
rect 2899 4082 3001 4114
rect 3033 4082 3135 4114
rect 2899 4046 3135 4082
rect 2899 4014 3001 4046
rect 3033 4014 3135 4046
rect 2899 3978 3135 4014
rect 2899 3946 3001 3978
rect 3033 3946 3135 3978
rect 2899 3910 3135 3946
rect 2899 3878 3001 3910
rect 3033 3878 3135 3910
rect 2899 3842 3135 3878
rect 2899 3810 3001 3842
rect 3033 3810 3135 3842
rect 2899 3774 3135 3810
rect 2899 3742 3001 3774
rect 3033 3742 3135 3774
rect 2899 3706 3135 3742
rect 2899 3674 3001 3706
rect 3033 3674 3135 3706
rect 2899 3638 3135 3674
rect 2899 3606 3001 3638
rect 3033 3606 3135 3638
rect 2899 3570 3135 3606
rect 2899 3538 3001 3570
rect 3033 3538 3135 3570
rect 2899 3502 3135 3538
rect 2899 3470 3001 3502
rect 3033 3470 3135 3502
rect 2899 3454 3135 3470
rect 3255 4318 3383 4334
rect 3255 4286 3303 4318
rect 3335 4286 3383 4318
rect 3255 4250 3383 4286
rect 3255 4218 3303 4250
rect 3335 4218 3383 4250
rect 3255 4182 3383 4218
rect 3255 4150 3303 4182
rect 3335 4150 3383 4182
rect 3255 4114 3383 4150
rect 3255 4082 3303 4114
rect 3335 4082 3383 4114
rect 3255 4046 3383 4082
rect 3255 4014 3303 4046
rect 3335 4014 3383 4046
rect 3255 3978 3383 4014
rect 3255 3946 3303 3978
rect 3335 3946 3383 3978
rect 3255 3910 3383 3946
rect 3255 3878 3303 3910
rect 3335 3878 3383 3910
rect 3255 3842 3383 3878
rect 3255 3810 3303 3842
rect 3335 3810 3383 3842
rect 3255 3774 3383 3810
rect 3255 3742 3303 3774
rect 3335 3742 3383 3774
rect 3255 3706 3383 3742
rect 3255 3674 3303 3706
rect 3335 3674 3383 3706
rect 3255 3638 3383 3674
rect 3255 3606 3303 3638
rect 3335 3606 3383 3638
rect 3255 3570 3383 3606
rect 3255 3538 3303 3570
rect 3335 3538 3383 3570
rect 3255 3502 3383 3538
rect 3255 3470 3303 3502
rect 3335 3470 3383 3502
rect 3255 3454 3383 3470
rect 3503 4318 3739 4334
rect 3503 4286 3605 4318
rect 3637 4286 3739 4318
rect 3503 4250 3739 4286
rect 3503 4218 3605 4250
rect 3637 4218 3739 4250
rect 3503 4182 3739 4218
rect 3503 4150 3605 4182
rect 3637 4150 3739 4182
rect 3503 4114 3739 4150
rect 3503 4082 3605 4114
rect 3637 4082 3739 4114
rect 3503 4046 3739 4082
rect 3503 4014 3605 4046
rect 3637 4014 3739 4046
rect 3503 3978 3739 4014
rect 3503 3946 3605 3978
rect 3637 3946 3739 3978
rect 3503 3910 3739 3946
rect 3503 3878 3605 3910
rect 3637 3878 3739 3910
rect 3503 3842 3739 3878
rect 3503 3810 3605 3842
rect 3637 3810 3739 3842
rect 3503 3774 3739 3810
rect 3503 3742 3605 3774
rect 3637 3742 3739 3774
rect 3503 3706 3739 3742
rect 3503 3674 3605 3706
rect 3637 3674 3739 3706
rect 3503 3638 3739 3674
rect 3503 3606 3605 3638
rect 3637 3606 3739 3638
rect 3503 3570 3739 3606
rect 3503 3538 3605 3570
rect 3637 3538 3739 3570
rect 3503 3502 3739 3538
rect 3503 3470 3605 3502
rect 3637 3470 3739 3502
rect 3503 3454 3739 3470
rect 3859 4318 3987 4334
rect 3859 4286 3907 4318
rect 3939 4286 3987 4318
rect 3859 4250 3987 4286
rect 3859 4218 3907 4250
rect 3939 4218 3987 4250
rect 3859 4182 3987 4218
rect 3859 4150 3907 4182
rect 3939 4150 3987 4182
rect 3859 4114 3987 4150
rect 3859 4082 3907 4114
rect 3939 4082 3987 4114
rect 3859 4046 3987 4082
rect 3859 4014 3907 4046
rect 3939 4014 3987 4046
rect 3859 3978 3987 4014
rect 3859 3946 3907 3978
rect 3939 3946 3987 3978
rect 3859 3910 3987 3946
rect 3859 3878 3907 3910
rect 3939 3878 3987 3910
rect 3859 3842 3987 3878
rect 3859 3810 3907 3842
rect 3939 3810 3987 3842
rect 3859 3774 3987 3810
rect 3859 3742 3907 3774
rect 3939 3742 3987 3774
rect 3859 3706 3987 3742
rect 3859 3674 3907 3706
rect 3939 3674 3987 3706
rect 3859 3638 3987 3674
rect 3859 3606 3907 3638
rect 3939 3606 3987 3638
rect 3859 3570 3987 3606
rect 3859 3538 3907 3570
rect 3939 3538 3987 3570
rect 3859 3502 3987 3538
rect 3859 3470 3907 3502
rect 3939 3470 3987 3502
rect 3859 3454 3987 3470
rect 4107 4318 4343 4334
rect 4107 4286 4209 4318
rect 4241 4286 4343 4318
rect 4107 4250 4343 4286
rect 4107 4218 4209 4250
rect 4241 4218 4343 4250
rect 4107 4182 4343 4218
rect 4107 4150 4209 4182
rect 4241 4150 4343 4182
rect 4107 4114 4343 4150
rect 4107 4082 4209 4114
rect 4241 4082 4343 4114
rect 4107 4046 4343 4082
rect 4107 4014 4209 4046
rect 4241 4014 4343 4046
rect 4107 3978 4343 4014
rect 4107 3946 4209 3978
rect 4241 3946 4343 3978
rect 4107 3910 4343 3946
rect 4107 3878 4209 3910
rect 4241 3878 4343 3910
rect 4107 3842 4343 3878
rect 4107 3810 4209 3842
rect 4241 3810 4343 3842
rect 4107 3774 4343 3810
rect 4107 3742 4209 3774
rect 4241 3742 4343 3774
rect 4107 3706 4343 3742
rect 4107 3674 4209 3706
rect 4241 3674 4343 3706
rect 4107 3638 4343 3674
rect 4107 3606 4209 3638
rect 4241 3606 4343 3638
rect 4107 3570 4343 3606
rect 4107 3538 4209 3570
rect 4241 3538 4343 3570
rect 4107 3502 4343 3538
rect 4107 3470 4209 3502
rect 4241 3470 4343 3502
rect 4107 3454 4343 3470
rect 4463 4318 4591 4334
rect 4463 4286 4511 4318
rect 4543 4286 4591 4318
rect 4463 4250 4591 4286
rect 4463 4218 4511 4250
rect 4543 4218 4591 4250
rect 4463 4182 4591 4218
rect 4463 4150 4511 4182
rect 4543 4150 4591 4182
rect 4463 4114 4591 4150
rect 4463 4082 4511 4114
rect 4543 4082 4591 4114
rect 4463 4046 4591 4082
rect 4463 4014 4511 4046
rect 4543 4014 4591 4046
rect 4463 3978 4591 4014
rect 4463 3946 4511 3978
rect 4543 3946 4591 3978
rect 4463 3910 4591 3946
rect 4463 3878 4511 3910
rect 4543 3878 4591 3910
rect 4463 3842 4591 3878
rect 4463 3810 4511 3842
rect 4543 3810 4591 3842
rect 4463 3774 4591 3810
rect 4463 3742 4511 3774
rect 4543 3742 4591 3774
rect 4463 3706 4591 3742
rect 4463 3674 4511 3706
rect 4543 3674 4591 3706
rect 4463 3638 4591 3674
rect 4463 3606 4511 3638
rect 4543 3606 4591 3638
rect 4463 3570 4591 3606
rect 4463 3538 4511 3570
rect 4543 3538 4591 3570
rect 4463 3502 4591 3538
rect 4463 3470 4511 3502
rect 4543 3470 4591 3502
rect 4463 3454 4591 3470
rect 4711 4318 4947 4334
rect 4711 4286 4813 4318
rect 4845 4286 4947 4318
rect 4711 4250 4947 4286
rect 4711 4218 4813 4250
rect 4845 4218 4947 4250
rect 4711 4182 4947 4218
rect 4711 4150 4813 4182
rect 4845 4150 4947 4182
rect 4711 4114 4947 4150
rect 4711 4082 4813 4114
rect 4845 4082 4947 4114
rect 4711 4046 4947 4082
rect 4711 4014 4813 4046
rect 4845 4014 4947 4046
rect 4711 3978 4947 4014
rect 4711 3946 4813 3978
rect 4845 3946 4947 3978
rect 4711 3910 4947 3946
rect 4711 3878 4813 3910
rect 4845 3878 4947 3910
rect 4711 3842 4947 3878
rect 4711 3810 4813 3842
rect 4845 3810 4947 3842
rect 4711 3774 4947 3810
rect 4711 3742 4813 3774
rect 4845 3742 4947 3774
rect 4711 3706 4947 3742
rect 4711 3674 4813 3706
rect 4845 3674 4947 3706
rect 4711 3638 4947 3674
rect 4711 3606 4813 3638
rect 4845 3606 4947 3638
rect 4711 3570 4947 3606
rect 4711 3538 4813 3570
rect 4845 3538 4947 3570
rect 4711 3502 4947 3538
rect 4711 3470 4813 3502
rect 4845 3470 4947 3502
rect 4711 3454 4947 3470
rect 5067 4318 5195 4334
rect 5067 4286 5115 4318
rect 5147 4286 5195 4318
rect 5067 4250 5195 4286
rect 5067 4218 5115 4250
rect 5147 4218 5195 4250
rect 5067 4182 5195 4218
rect 5067 4150 5115 4182
rect 5147 4150 5195 4182
rect 5067 4114 5195 4150
rect 5067 4082 5115 4114
rect 5147 4082 5195 4114
rect 5067 4046 5195 4082
rect 5067 4014 5115 4046
rect 5147 4014 5195 4046
rect 5067 3978 5195 4014
rect 5067 3946 5115 3978
rect 5147 3946 5195 3978
rect 5067 3910 5195 3946
rect 5067 3878 5115 3910
rect 5147 3878 5195 3910
rect 5067 3842 5195 3878
rect 5067 3810 5115 3842
rect 5147 3810 5195 3842
rect 5067 3774 5195 3810
rect 5067 3742 5115 3774
rect 5147 3742 5195 3774
rect 5067 3706 5195 3742
rect 5067 3674 5115 3706
rect 5147 3674 5195 3706
rect 5067 3638 5195 3674
rect 5067 3606 5115 3638
rect 5147 3606 5195 3638
rect 5067 3570 5195 3606
rect 5067 3538 5115 3570
rect 5147 3538 5195 3570
rect 5067 3502 5195 3538
rect 5067 3470 5115 3502
rect 5147 3470 5195 3502
rect 5067 3454 5195 3470
rect 5315 4318 5551 4334
rect 5315 4286 5417 4318
rect 5449 4286 5551 4318
rect 5315 4250 5551 4286
rect 5315 4218 5417 4250
rect 5449 4218 5551 4250
rect 5315 4182 5551 4218
rect 5315 4150 5417 4182
rect 5449 4150 5551 4182
rect 5315 4114 5551 4150
rect 5315 4082 5417 4114
rect 5449 4082 5551 4114
rect 5315 4046 5551 4082
rect 5315 4014 5417 4046
rect 5449 4014 5551 4046
rect 5315 3978 5551 4014
rect 5315 3946 5417 3978
rect 5449 3946 5551 3978
rect 5315 3910 5551 3946
rect 5315 3878 5417 3910
rect 5449 3878 5551 3910
rect 5315 3842 5551 3878
rect 5315 3810 5417 3842
rect 5449 3810 5551 3842
rect 5315 3774 5551 3810
rect 5315 3742 5417 3774
rect 5449 3742 5551 3774
rect 5315 3706 5551 3742
rect 5315 3674 5417 3706
rect 5449 3674 5551 3706
rect 5315 3638 5551 3674
rect 5315 3606 5417 3638
rect 5449 3606 5551 3638
rect 5315 3570 5551 3606
rect 5315 3538 5417 3570
rect 5449 3538 5551 3570
rect 5315 3502 5551 3538
rect 5315 3470 5417 3502
rect 5449 3470 5551 3502
rect 5315 3454 5551 3470
rect 5671 4318 5799 4334
rect 5671 4286 5719 4318
rect 5751 4286 5799 4318
rect 5671 4250 5799 4286
rect 5671 4218 5719 4250
rect 5751 4218 5799 4250
rect 5671 4182 5799 4218
rect 5671 4150 5719 4182
rect 5751 4150 5799 4182
rect 5671 4114 5799 4150
rect 5671 4082 5719 4114
rect 5751 4082 5799 4114
rect 5671 4046 5799 4082
rect 5671 4014 5719 4046
rect 5751 4014 5799 4046
rect 5671 3978 5799 4014
rect 5671 3946 5719 3978
rect 5751 3946 5799 3978
rect 5671 3910 5799 3946
rect 5671 3878 5719 3910
rect 5751 3878 5799 3910
rect 5671 3842 5799 3878
rect 5671 3810 5719 3842
rect 5751 3810 5799 3842
rect 5671 3774 5799 3810
rect 5671 3742 5719 3774
rect 5751 3742 5799 3774
rect 5671 3706 5799 3742
rect 5671 3674 5719 3706
rect 5751 3674 5799 3706
rect 5671 3638 5799 3674
rect 5671 3606 5719 3638
rect 5751 3606 5799 3638
rect 5671 3570 5799 3606
rect 5671 3538 5719 3570
rect 5751 3538 5799 3570
rect 5671 3502 5799 3538
rect 5671 3470 5719 3502
rect 5751 3470 5799 3502
rect 5671 3454 5799 3470
rect 5919 4318 6155 4334
rect 5919 4286 6021 4318
rect 6053 4286 6155 4318
rect 5919 4250 6155 4286
rect 5919 4218 6021 4250
rect 6053 4218 6155 4250
rect 5919 4182 6155 4218
rect 5919 4150 6021 4182
rect 6053 4150 6155 4182
rect 5919 4114 6155 4150
rect 5919 4082 6021 4114
rect 6053 4082 6155 4114
rect 5919 4046 6155 4082
rect 5919 4014 6021 4046
rect 6053 4014 6155 4046
rect 5919 3978 6155 4014
rect 5919 3946 6021 3978
rect 6053 3946 6155 3978
rect 5919 3910 6155 3946
rect 5919 3878 6021 3910
rect 6053 3878 6155 3910
rect 5919 3842 6155 3878
rect 5919 3810 6021 3842
rect 6053 3810 6155 3842
rect 5919 3774 6155 3810
rect 5919 3742 6021 3774
rect 6053 3742 6155 3774
rect 5919 3706 6155 3742
rect 5919 3674 6021 3706
rect 6053 3674 6155 3706
rect 5919 3638 6155 3674
rect 5919 3606 6021 3638
rect 6053 3606 6155 3638
rect 5919 3570 6155 3606
rect 5919 3538 6021 3570
rect 6053 3538 6155 3570
rect 5919 3502 6155 3538
rect 5919 3470 6021 3502
rect 6053 3470 6155 3502
rect 5919 3454 6155 3470
rect 6275 4318 6403 4334
rect 6275 4286 6323 4318
rect 6355 4286 6403 4318
rect 6275 4250 6403 4286
rect 6275 4218 6323 4250
rect 6355 4218 6403 4250
rect 6275 4182 6403 4218
rect 6275 4150 6323 4182
rect 6355 4150 6403 4182
rect 6275 4114 6403 4150
rect 6275 4082 6323 4114
rect 6355 4082 6403 4114
rect 6275 4046 6403 4082
rect 6275 4014 6323 4046
rect 6355 4014 6403 4046
rect 6275 3978 6403 4014
rect 6275 3946 6323 3978
rect 6355 3946 6403 3978
rect 6275 3910 6403 3946
rect 6275 3878 6323 3910
rect 6355 3878 6403 3910
rect 6275 3842 6403 3878
rect 6275 3810 6323 3842
rect 6355 3810 6403 3842
rect 6275 3774 6403 3810
rect 6275 3742 6323 3774
rect 6355 3742 6403 3774
rect 6275 3706 6403 3742
rect 6275 3674 6323 3706
rect 6355 3674 6403 3706
rect 6275 3638 6403 3674
rect 6275 3606 6323 3638
rect 6355 3606 6403 3638
rect 6275 3570 6403 3606
rect 6275 3538 6323 3570
rect 6355 3538 6403 3570
rect 6275 3502 6403 3538
rect 6275 3470 6323 3502
rect 6355 3470 6403 3502
rect 6275 3454 6403 3470
rect 6523 4318 6759 4334
rect 6523 4286 6625 4318
rect 6657 4286 6759 4318
rect 6523 4250 6759 4286
rect 6523 4218 6625 4250
rect 6657 4218 6759 4250
rect 6523 4182 6759 4218
rect 6523 4150 6625 4182
rect 6657 4150 6759 4182
rect 6523 4114 6759 4150
rect 6523 4082 6625 4114
rect 6657 4082 6759 4114
rect 6523 4046 6759 4082
rect 6523 4014 6625 4046
rect 6657 4014 6759 4046
rect 6523 3978 6759 4014
rect 6523 3946 6625 3978
rect 6657 3946 6759 3978
rect 6523 3910 6759 3946
rect 6523 3878 6625 3910
rect 6657 3878 6759 3910
rect 6523 3842 6759 3878
rect 6523 3810 6625 3842
rect 6657 3810 6759 3842
rect 6523 3774 6759 3810
rect 6523 3742 6625 3774
rect 6657 3742 6759 3774
rect 6523 3706 6759 3742
rect 6523 3674 6625 3706
rect 6657 3674 6759 3706
rect 6523 3638 6759 3674
rect 6523 3606 6625 3638
rect 6657 3606 6759 3638
rect 6523 3570 6759 3606
rect 6523 3538 6625 3570
rect 6657 3538 6759 3570
rect 6523 3502 6759 3538
rect 6523 3470 6625 3502
rect 6657 3470 6759 3502
rect 6523 3454 6759 3470
rect 6879 4318 7007 4334
rect 6879 4286 6927 4318
rect 6959 4286 7007 4318
rect 6879 4250 7007 4286
rect 6879 4218 6927 4250
rect 6959 4218 7007 4250
rect 6879 4182 7007 4218
rect 6879 4150 6927 4182
rect 6959 4150 7007 4182
rect 6879 4114 7007 4150
rect 6879 4082 6927 4114
rect 6959 4082 7007 4114
rect 6879 4046 7007 4082
rect 6879 4014 6927 4046
rect 6959 4014 7007 4046
rect 6879 3978 7007 4014
rect 6879 3946 6927 3978
rect 6959 3946 7007 3978
rect 6879 3910 7007 3946
rect 6879 3878 6927 3910
rect 6959 3878 7007 3910
rect 6879 3842 7007 3878
rect 6879 3810 6927 3842
rect 6959 3810 7007 3842
rect 6879 3774 7007 3810
rect 6879 3742 6927 3774
rect 6959 3742 7007 3774
rect 6879 3706 7007 3742
rect 6879 3674 6927 3706
rect 6959 3674 7007 3706
rect 6879 3638 7007 3674
rect 6879 3606 6927 3638
rect 6959 3606 7007 3638
rect 6879 3570 7007 3606
rect 6879 3538 6927 3570
rect 6959 3538 7007 3570
rect 6879 3502 7007 3538
rect 6879 3470 6927 3502
rect 6959 3470 7007 3502
rect 6879 3454 7007 3470
rect 7127 4318 7363 4334
rect 7127 4286 7229 4318
rect 7261 4286 7363 4318
rect 7127 4250 7363 4286
rect 7127 4218 7229 4250
rect 7261 4218 7363 4250
rect 7127 4182 7363 4218
rect 7127 4150 7229 4182
rect 7261 4150 7363 4182
rect 7127 4114 7363 4150
rect 7127 4082 7229 4114
rect 7261 4082 7363 4114
rect 7127 4046 7363 4082
rect 7127 4014 7229 4046
rect 7261 4014 7363 4046
rect 7127 3978 7363 4014
rect 7127 3946 7229 3978
rect 7261 3946 7363 3978
rect 7127 3910 7363 3946
rect 7127 3878 7229 3910
rect 7261 3878 7363 3910
rect 7127 3842 7363 3878
rect 7127 3810 7229 3842
rect 7261 3810 7363 3842
rect 7127 3774 7363 3810
rect 7127 3742 7229 3774
rect 7261 3742 7363 3774
rect 7127 3706 7363 3742
rect 7127 3674 7229 3706
rect 7261 3674 7363 3706
rect 7127 3638 7363 3674
rect 7127 3606 7229 3638
rect 7261 3606 7363 3638
rect 7127 3570 7363 3606
rect 7127 3538 7229 3570
rect 7261 3538 7363 3570
rect 7127 3502 7363 3538
rect 7127 3470 7229 3502
rect 7261 3470 7363 3502
rect 7127 3454 7363 3470
rect 7483 4318 7611 4334
rect 7483 4286 7531 4318
rect 7563 4286 7611 4318
rect 7483 4250 7611 4286
rect 7483 4218 7531 4250
rect 7563 4218 7611 4250
rect 7483 4182 7611 4218
rect 7483 4150 7531 4182
rect 7563 4150 7611 4182
rect 7483 4114 7611 4150
rect 7483 4082 7531 4114
rect 7563 4082 7611 4114
rect 7483 4046 7611 4082
rect 7483 4014 7531 4046
rect 7563 4014 7611 4046
rect 7483 3978 7611 4014
rect 7483 3946 7531 3978
rect 7563 3946 7611 3978
rect 7483 3910 7611 3946
rect 7483 3878 7531 3910
rect 7563 3878 7611 3910
rect 7483 3842 7611 3878
rect 7483 3810 7531 3842
rect 7563 3810 7611 3842
rect 7483 3774 7611 3810
rect 7483 3742 7531 3774
rect 7563 3742 7611 3774
rect 7483 3706 7611 3742
rect 7483 3674 7531 3706
rect 7563 3674 7611 3706
rect 7483 3638 7611 3674
rect 7483 3606 7531 3638
rect 7563 3606 7611 3638
rect 7483 3570 7611 3606
rect 7483 3538 7531 3570
rect 7563 3538 7611 3570
rect 7483 3502 7611 3538
rect 7483 3470 7531 3502
rect 7563 3470 7611 3502
rect 7483 3454 7611 3470
rect 7731 4318 7967 4334
rect 7731 4286 7833 4318
rect 7865 4286 7967 4318
rect 7731 4250 7967 4286
rect 7731 4218 7833 4250
rect 7865 4218 7967 4250
rect 7731 4182 7967 4218
rect 7731 4150 7833 4182
rect 7865 4150 7967 4182
rect 7731 4114 7967 4150
rect 7731 4082 7833 4114
rect 7865 4082 7967 4114
rect 7731 4046 7967 4082
rect 7731 4014 7833 4046
rect 7865 4014 7967 4046
rect 7731 3978 7967 4014
rect 7731 3946 7833 3978
rect 7865 3946 7967 3978
rect 7731 3910 7967 3946
rect 7731 3878 7833 3910
rect 7865 3878 7967 3910
rect 7731 3842 7967 3878
rect 7731 3810 7833 3842
rect 7865 3810 7967 3842
rect 7731 3774 7967 3810
rect 7731 3742 7833 3774
rect 7865 3742 7967 3774
rect 7731 3706 7967 3742
rect 7731 3674 7833 3706
rect 7865 3674 7967 3706
rect 7731 3638 7967 3674
rect 7731 3606 7833 3638
rect 7865 3606 7967 3638
rect 7731 3570 7967 3606
rect 7731 3538 7833 3570
rect 7865 3538 7967 3570
rect 7731 3502 7967 3538
rect 7731 3470 7833 3502
rect 7865 3470 7967 3502
rect 7731 3454 7967 3470
rect 8087 4318 8215 4334
rect 8087 4286 8135 4318
rect 8167 4286 8215 4318
rect 8087 4250 8215 4286
rect 8087 4218 8135 4250
rect 8167 4218 8215 4250
rect 8087 4182 8215 4218
rect 8087 4150 8135 4182
rect 8167 4150 8215 4182
rect 8087 4114 8215 4150
rect 8087 4082 8135 4114
rect 8167 4082 8215 4114
rect 8087 4046 8215 4082
rect 8087 4014 8135 4046
rect 8167 4014 8215 4046
rect 8087 3978 8215 4014
rect 8087 3946 8135 3978
rect 8167 3946 8215 3978
rect 8087 3910 8215 3946
rect 8087 3878 8135 3910
rect 8167 3878 8215 3910
rect 8087 3842 8215 3878
rect 8087 3810 8135 3842
rect 8167 3810 8215 3842
rect 8087 3774 8215 3810
rect 8087 3742 8135 3774
rect 8167 3742 8215 3774
rect 8087 3706 8215 3742
rect 8087 3674 8135 3706
rect 8167 3674 8215 3706
rect 8087 3638 8215 3674
rect 8087 3606 8135 3638
rect 8167 3606 8215 3638
rect 8087 3570 8215 3606
rect 8087 3538 8135 3570
rect 8167 3538 8215 3570
rect 8087 3502 8215 3538
rect 8087 3470 8135 3502
rect 8167 3470 8215 3502
rect 8087 3454 8215 3470
rect 8335 4318 8571 4334
rect 8335 4286 8437 4318
rect 8469 4286 8571 4318
rect 8335 4250 8571 4286
rect 8335 4218 8437 4250
rect 8469 4218 8571 4250
rect 8335 4182 8571 4218
rect 8335 4150 8437 4182
rect 8469 4150 8571 4182
rect 8335 4114 8571 4150
rect 8335 4082 8437 4114
rect 8469 4082 8571 4114
rect 8335 4046 8571 4082
rect 8335 4014 8437 4046
rect 8469 4014 8571 4046
rect 8335 3978 8571 4014
rect 8335 3946 8437 3978
rect 8469 3946 8571 3978
rect 8335 3910 8571 3946
rect 8335 3878 8437 3910
rect 8469 3878 8571 3910
rect 8335 3842 8571 3878
rect 8335 3810 8437 3842
rect 8469 3810 8571 3842
rect 8335 3774 8571 3810
rect 8335 3742 8437 3774
rect 8469 3742 8571 3774
rect 8335 3706 8571 3742
rect 8335 3674 8437 3706
rect 8469 3674 8571 3706
rect 8335 3638 8571 3674
rect 8335 3606 8437 3638
rect 8469 3606 8571 3638
rect 8335 3570 8571 3606
rect 8335 3538 8437 3570
rect 8469 3538 8571 3570
rect 8335 3502 8571 3538
rect 8335 3470 8437 3502
rect 8469 3470 8571 3502
rect 8335 3454 8571 3470
rect 8691 4318 8819 4334
rect 8691 4286 8739 4318
rect 8771 4286 8819 4318
rect 8691 4250 8819 4286
rect 8691 4218 8739 4250
rect 8771 4218 8819 4250
rect 8691 4182 8819 4218
rect 8691 4150 8739 4182
rect 8771 4150 8819 4182
rect 8691 4114 8819 4150
rect 8691 4082 8739 4114
rect 8771 4082 8819 4114
rect 8691 4046 8819 4082
rect 8691 4014 8739 4046
rect 8771 4014 8819 4046
rect 8691 3978 8819 4014
rect 8691 3946 8739 3978
rect 8771 3946 8819 3978
rect 8691 3910 8819 3946
rect 8691 3878 8739 3910
rect 8771 3878 8819 3910
rect 8691 3842 8819 3878
rect 8691 3810 8739 3842
rect 8771 3810 8819 3842
rect 8691 3774 8819 3810
rect 8691 3742 8739 3774
rect 8771 3742 8819 3774
rect 8691 3706 8819 3742
rect 8691 3674 8739 3706
rect 8771 3674 8819 3706
rect 8691 3638 8819 3674
rect 8691 3606 8739 3638
rect 8771 3606 8819 3638
rect 8691 3570 8819 3606
rect 8691 3538 8739 3570
rect 8771 3538 8819 3570
rect 8691 3502 8819 3538
rect 8691 3470 8739 3502
rect 8771 3470 8819 3502
rect 8691 3454 8819 3470
rect 8939 4318 9175 4334
rect 8939 4286 9041 4318
rect 9073 4286 9175 4318
rect 8939 4250 9175 4286
rect 8939 4218 9041 4250
rect 9073 4218 9175 4250
rect 8939 4182 9175 4218
rect 8939 4150 9041 4182
rect 9073 4150 9175 4182
rect 8939 4114 9175 4150
rect 8939 4082 9041 4114
rect 9073 4082 9175 4114
rect 8939 4046 9175 4082
rect 8939 4014 9041 4046
rect 9073 4014 9175 4046
rect 8939 3978 9175 4014
rect 8939 3946 9041 3978
rect 9073 3946 9175 3978
rect 8939 3910 9175 3946
rect 8939 3878 9041 3910
rect 9073 3878 9175 3910
rect 8939 3842 9175 3878
rect 8939 3810 9041 3842
rect 9073 3810 9175 3842
rect 8939 3774 9175 3810
rect 8939 3742 9041 3774
rect 9073 3742 9175 3774
rect 8939 3706 9175 3742
rect 8939 3674 9041 3706
rect 9073 3674 9175 3706
rect 8939 3638 9175 3674
rect 8939 3606 9041 3638
rect 9073 3606 9175 3638
rect 8939 3570 9175 3606
rect 8939 3538 9041 3570
rect 9073 3538 9175 3570
rect 8939 3502 9175 3538
rect 8939 3470 9041 3502
rect 9073 3470 9175 3502
rect 8939 3454 9175 3470
rect 9295 4318 9423 4334
rect 9295 4286 9343 4318
rect 9375 4286 9423 4318
rect 9295 4250 9423 4286
rect 9295 4218 9343 4250
rect 9375 4218 9423 4250
rect 9295 4182 9423 4218
rect 9295 4150 9343 4182
rect 9375 4150 9423 4182
rect 9295 4114 9423 4150
rect 9295 4082 9343 4114
rect 9375 4082 9423 4114
rect 9295 4046 9423 4082
rect 9295 4014 9343 4046
rect 9375 4014 9423 4046
rect 9295 3978 9423 4014
rect 9295 3946 9343 3978
rect 9375 3946 9423 3978
rect 9295 3910 9423 3946
rect 9295 3878 9343 3910
rect 9375 3878 9423 3910
rect 9295 3842 9423 3878
rect 9295 3810 9343 3842
rect 9375 3810 9423 3842
rect 9295 3774 9423 3810
rect 9295 3742 9343 3774
rect 9375 3742 9423 3774
rect 9295 3706 9423 3742
rect 9295 3674 9343 3706
rect 9375 3674 9423 3706
rect 9295 3638 9423 3674
rect 9295 3606 9343 3638
rect 9375 3606 9423 3638
rect 9295 3570 9423 3606
rect 9295 3538 9343 3570
rect 9375 3538 9423 3570
rect 9295 3502 9423 3538
rect 9295 3470 9343 3502
rect 9375 3470 9423 3502
rect 9295 3454 9423 3470
rect 9543 4318 9779 4334
rect 9543 4286 9645 4318
rect 9677 4286 9779 4318
rect 9543 4250 9779 4286
rect 9543 4218 9645 4250
rect 9677 4218 9779 4250
rect 9543 4182 9779 4218
rect 9543 4150 9645 4182
rect 9677 4150 9779 4182
rect 9543 4114 9779 4150
rect 9543 4082 9645 4114
rect 9677 4082 9779 4114
rect 9543 4046 9779 4082
rect 9543 4014 9645 4046
rect 9677 4014 9779 4046
rect 9543 3978 9779 4014
rect 9543 3946 9645 3978
rect 9677 3946 9779 3978
rect 9543 3910 9779 3946
rect 9543 3878 9645 3910
rect 9677 3878 9779 3910
rect 9543 3842 9779 3878
rect 9543 3810 9645 3842
rect 9677 3810 9779 3842
rect 9543 3774 9779 3810
rect 9543 3742 9645 3774
rect 9677 3742 9779 3774
rect 9543 3706 9779 3742
rect 9543 3674 9645 3706
rect 9677 3674 9779 3706
rect 9543 3638 9779 3674
rect 9543 3606 9645 3638
rect 9677 3606 9779 3638
rect 9543 3570 9779 3606
rect 9543 3538 9645 3570
rect 9677 3538 9779 3570
rect 9543 3502 9779 3538
rect 9543 3470 9645 3502
rect 9677 3470 9779 3502
rect 9543 3454 9779 3470
rect 9899 4318 10027 4334
rect 9899 4286 9947 4318
rect 9979 4286 10027 4318
rect 9899 4250 10027 4286
rect 9899 4218 9947 4250
rect 9979 4218 10027 4250
rect 9899 4182 10027 4218
rect 9899 4150 9947 4182
rect 9979 4150 10027 4182
rect 9899 4114 10027 4150
rect 9899 4082 9947 4114
rect 9979 4082 10027 4114
rect 9899 4046 10027 4082
rect 9899 4014 9947 4046
rect 9979 4014 10027 4046
rect 9899 3978 10027 4014
rect 9899 3946 9947 3978
rect 9979 3946 10027 3978
rect 9899 3910 10027 3946
rect 9899 3878 9947 3910
rect 9979 3878 10027 3910
rect 9899 3842 10027 3878
rect 9899 3810 9947 3842
rect 9979 3810 10027 3842
rect 9899 3774 10027 3810
rect 9899 3742 9947 3774
rect 9979 3742 10027 3774
rect 9899 3706 10027 3742
rect 9899 3674 9947 3706
rect 9979 3674 10027 3706
rect 9899 3638 10027 3674
rect 9899 3606 9947 3638
rect 9979 3606 10027 3638
rect 9899 3570 10027 3606
rect 9899 3538 9947 3570
rect 9979 3538 10027 3570
rect 9899 3502 10027 3538
rect 9899 3470 9947 3502
rect 9979 3470 10027 3502
rect 9899 3454 10027 3470
rect 10147 4318 10383 4334
rect 10147 4286 10249 4318
rect 10281 4286 10383 4318
rect 10147 4250 10383 4286
rect 10147 4218 10249 4250
rect 10281 4218 10383 4250
rect 10147 4182 10383 4218
rect 10147 4150 10249 4182
rect 10281 4150 10383 4182
rect 10147 4114 10383 4150
rect 10147 4082 10249 4114
rect 10281 4082 10383 4114
rect 10147 4046 10383 4082
rect 10147 4014 10249 4046
rect 10281 4014 10383 4046
rect 10147 3978 10383 4014
rect 10147 3946 10249 3978
rect 10281 3946 10383 3978
rect 10147 3910 10383 3946
rect 10147 3878 10249 3910
rect 10281 3878 10383 3910
rect 10147 3842 10383 3878
rect 10147 3810 10249 3842
rect 10281 3810 10383 3842
rect 10147 3774 10383 3810
rect 10147 3742 10249 3774
rect 10281 3742 10383 3774
rect 10147 3706 10383 3742
rect 10147 3674 10249 3706
rect 10281 3674 10383 3706
rect 10147 3638 10383 3674
rect 10147 3606 10249 3638
rect 10281 3606 10383 3638
rect 10147 3570 10383 3606
rect 10147 3538 10249 3570
rect 10281 3538 10383 3570
rect 10147 3502 10383 3538
rect 10147 3470 10249 3502
rect 10281 3470 10383 3502
rect 10147 3454 10383 3470
rect 10503 4318 10631 4334
rect 10503 4286 10551 4318
rect 10583 4286 10631 4318
rect 10503 4250 10631 4286
rect 10503 4218 10551 4250
rect 10583 4218 10631 4250
rect 10503 4182 10631 4218
rect 10503 4150 10551 4182
rect 10583 4150 10631 4182
rect 10503 4114 10631 4150
rect 10503 4082 10551 4114
rect 10583 4082 10631 4114
rect 10503 4046 10631 4082
rect 10503 4014 10551 4046
rect 10583 4014 10631 4046
rect 10503 3978 10631 4014
rect 10503 3946 10551 3978
rect 10583 3946 10631 3978
rect 10503 3910 10631 3946
rect 10503 3878 10551 3910
rect 10583 3878 10631 3910
rect 10503 3842 10631 3878
rect 10503 3810 10551 3842
rect 10583 3810 10631 3842
rect 10503 3774 10631 3810
rect 10503 3742 10551 3774
rect 10583 3742 10631 3774
rect 10503 3706 10631 3742
rect 10503 3674 10551 3706
rect 10583 3674 10631 3706
rect 10503 3638 10631 3674
rect 10503 3606 10551 3638
rect 10583 3606 10631 3638
rect 10503 3570 10631 3606
rect 10503 3538 10551 3570
rect 10583 3538 10631 3570
rect 10503 3502 10631 3538
rect 10503 3470 10551 3502
rect 10583 3470 10631 3502
rect 10503 3454 10631 3470
rect 10751 4318 10987 4334
rect 10751 4286 10853 4318
rect 10885 4286 10987 4318
rect 10751 4250 10987 4286
rect 10751 4218 10853 4250
rect 10885 4218 10987 4250
rect 10751 4182 10987 4218
rect 10751 4150 10853 4182
rect 10885 4150 10987 4182
rect 10751 4114 10987 4150
rect 10751 4082 10853 4114
rect 10885 4082 10987 4114
rect 10751 4046 10987 4082
rect 10751 4014 10853 4046
rect 10885 4014 10987 4046
rect 10751 3978 10987 4014
rect 10751 3946 10853 3978
rect 10885 3946 10987 3978
rect 10751 3910 10987 3946
rect 10751 3878 10853 3910
rect 10885 3878 10987 3910
rect 10751 3842 10987 3878
rect 10751 3810 10853 3842
rect 10885 3810 10987 3842
rect 10751 3774 10987 3810
rect 10751 3742 10853 3774
rect 10885 3742 10987 3774
rect 10751 3706 10987 3742
rect 10751 3674 10853 3706
rect 10885 3674 10987 3706
rect 10751 3638 10987 3674
rect 10751 3606 10853 3638
rect 10885 3606 10987 3638
rect 10751 3570 10987 3606
rect 10751 3538 10853 3570
rect 10885 3538 10987 3570
rect 10751 3502 10987 3538
rect 10751 3470 10853 3502
rect 10885 3470 10987 3502
rect 10751 3454 10987 3470
rect 11107 4318 11235 4334
rect 11107 4286 11155 4318
rect 11187 4286 11235 4318
rect 11107 4250 11235 4286
rect 11107 4218 11155 4250
rect 11187 4218 11235 4250
rect 11107 4182 11235 4218
rect 11107 4150 11155 4182
rect 11187 4150 11235 4182
rect 11107 4114 11235 4150
rect 11107 4082 11155 4114
rect 11187 4082 11235 4114
rect 11107 4046 11235 4082
rect 11107 4014 11155 4046
rect 11187 4014 11235 4046
rect 11107 3978 11235 4014
rect 11107 3946 11155 3978
rect 11187 3946 11235 3978
rect 11107 3910 11235 3946
rect 11107 3878 11155 3910
rect 11187 3878 11235 3910
rect 11107 3842 11235 3878
rect 11107 3810 11155 3842
rect 11187 3810 11235 3842
rect 11107 3774 11235 3810
rect 11107 3742 11155 3774
rect 11187 3742 11235 3774
rect 11107 3706 11235 3742
rect 11107 3674 11155 3706
rect 11187 3674 11235 3706
rect 11107 3638 11235 3674
rect 11107 3606 11155 3638
rect 11187 3606 11235 3638
rect 11107 3570 11235 3606
rect 11107 3538 11155 3570
rect 11187 3538 11235 3570
rect 11107 3502 11235 3538
rect 11107 3470 11155 3502
rect 11187 3470 11235 3502
rect 11107 3454 11235 3470
rect 11355 4318 11591 4334
rect 11355 4286 11457 4318
rect 11489 4286 11591 4318
rect 11355 4250 11591 4286
rect 11355 4218 11457 4250
rect 11489 4218 11591 4250
rect 11355 4182 11591 4218
rect 11355 4150 11457 4182
rect 11489 4150 11591 4182
rect 11355 4114 11591 4150
rect 11355 4082 11457 4114
rect 11489 4082 11591 4114
rect 11355 4046 11591 4082
rect 11355 4014 11457 4046
rect 11489 4014 11591 4046
rect 11355 3978 11591 4014
rect 11355 3946 11457 3978
rect 11489 3946 11591 3978
rect 11355 3910 11591 3946
rect 11355 3878 11457 3910
rect 11489 3878 11591 3910
rect 11355 3842 11591 3878
rect 11355 3810 11457 3842
rect 11489 3810 11591 3842
rect 11355 3774 11591 3810
rect 11355 3742 11457 3774
rect 11489 3742 11591 3774
rect 11355 3706 11591 3742
rect 11355 3674 11457 3706
rect 11489 3674 11591 3706
rect 11355 3638 11591 3674
rect 11355 3606 11457 3638
rect 11489 3606 11591 3638
rect 11355 3570 11591 3606
rect 11355 3538 11457 3570
rect 11489 3538 11591 3570
rect 11355 3502 11591 3538
rect 11355 3470 11457 3502
rect 11489 3470 11591 3502
rect 11355 3454 11591 3470
rect 11711 4318 11839 4334
rect 11711 4286 11759 4318
rect 11791 4286 11839 4318
rect 11711 4250 11839 4286
rect 11711 4218 11759 4250
rect 11791 4218 11839 4250
rect 11711 4182 11839 4218
rect 11711 4150 11759 4182
rect 11791 4150 11839 4182
rect 11711 4114 11839 4150
rect 11711 4082 11759 4114
rect 11791 4082 11839 4114
rect 11711 4046 11839 4082
rect 11711 4014 11759 4046
rect 11791 4014 11839 4046
rect 11711 3978 11839 4014
rect 11711 3946 11759 3978
rect 11791 3946 11839 3978
rect 11711 3910 11839 3946
rect 11711 3878 11759 3910
rect 11791 3878 11839 3910
rect 11711 3842 11839 3878
rect 11711 3810 11759 3842
rect 11791 3810 11839 3842
rect 11711 3774 11839 3810
rect 11711 3742 11759 3774
rect 11791 3742 11839 3774
rect 11711 3706 11839 3742
rect 11711 3674 11759 3706
rect 11791 3674 11839 3706
rect 11711 3638 11839 3674
rect 11711 3606 11759 3638
rect 11791 3606 11839 3638
rect 11711 3570 11839 3606
rect 11711 3538 11759 3570
rect 11791 3538 11839 3570
rect 11711 3502 11839 3538
rect 11711 3470 11759 3502
rect 11791 3470 11839 3502
rect 11711 3454 11839 3470
rect 11959 4318 12195 4334
rect 11959 4286 12061 4318
rect 12093 4286 12195 4318
rect 11959 4250 12195 4286
rect 11959 4218 12061 4250
rect 12093 4218 12195 4250
rect 11959 4182 12195 4218
rect 11959 4150 12061 4182
rect 12093 4150 12195 4182
rect 11959 4114 12195 4150
rect 11959 4082 12061 4114
rect 12093 4082 12195 4114
rect 11959 4046 12195 4082
rect 11959 4014 12061 4046
rect 12093 4014 12195 4046
rect 11959 3978 12195 4014
rect 11959 3946 12061 3978
rect 12093 3946 12195 3978
rect 11959 3910 12195 3946
rect 11959 3878 12061 3910
rect 12093 3878 12195 3910
rect 11959 3842 12195 3878
rect 11959 3810 12061 3842
rect 12093 3810 12195 3842
rect 11959 3774 12195 3810
rect 11959 3742 12061 3774
rect 12093 3742 12195 3774
rect 11959 3706 12195 3742
rect 11959 3674 12061 3706
rect 12093 3674 12195 3706
rect 11959 3638 12195 3674
rect 11959 3606 12061 3638
rect 12093 3606 12195 3638
rect 11959 3570 12195 3606
rect 11959 3538 12061 3570
rect 12093 3538 12195 3570
rect 11959 3502 12195 3538
rect 11959 3470 12061 3502
rect 12093 3470 12195 3502
rect 11959 3454 12195 3470
rect 12315 4318 12443 4334
rect 12315 4286 12363 4318
rect 12395 4286 12443 4318
rect 12315 4250 12443 4286
rect 12315 4218 12363 4250
rect 12395 4218 12443 4250
rect 12315 4182 12443 4218
rect 12315 4150 12363 4182
rect 12395 4150 12443 4182
rect 12315 4114 12443 4150
rect 12315 4082 12363 4114
rect 12395 4082 12443 4114
rect 12315 4046 12443 4082
rect 12315 4014 12363 4046
rect 12395 4014 12443 4046
rect 12315 3978 12443 4014
rect 12315 3946 12363 3978
rect 12395 3946 12443 3978
rect 12315 3910 12443 3946
rect 12315 3878 12363 3910
rect 12395 3878 12443 3910
rect 12315 3842 12443 3878
rect 12315 3810 12363 3842
rect 12395 3810 12443 3842
rect 12315 3774 12443 3810
rect 12315 3742 12363 3774
rect 12395 3742 12443 3774
rect 12315 3706 12443 3742
rect 12315 3674 12363 3706
rect 12395 3674 12443 3706
rect 12315 3638 12443 3674
rect 12315 3606 12363 3638
rect 12395 3606 12443 3638
rect 12315 3570 12443 3606
rect 12315 3538 12363 3570
rect 12395 3538 12443 3570
rect 12315 3502 12443 3538
rect 12315 3470 12363 3502
rect 12395 3470 12443 3502
rect 12315 3454 12443 3470
rect 12563 4318 12799 4334
rect 12563 4286 12665 4318
rect 12697 4286 12799 4318
rect 12563 4250 12799 4286
rect 12563 4218 12665 4250
rect 12697 4218 12799 4250
rect 12563 4182 12799 4218
rect 12563 4150 12665 4182
rect 12697 4150 12799 4182
rect 12563 4114 12799 4150
rect 12563 4082 12665 4114
rect 12697 4082 12799 4114
rect 12563 4046 12799 4082
rect 12563 4014 12665 4046
rect 12697 4014 12799 4046
rect 12563 3978 12799 4014
rect 12563 3946 12665 3978
rect 12697 3946 12799 3978
rect 12563 3910 12799 3946
rect 12563 3878 12665 3910
rect 12697 3878 12799 3910
rect 12563 3842 12799 3878
rect 12563 3810 12665 3842
rect 12697 3810 12799 3842
rect 12563 3774 12799 3810
rect 12563 3742 12665 3774
rect 12697 3742 12799 3774
rect 12563 3706 12799 3742
rect 12563 3674 12665 3706
rect 12697 3674 12799 3706
rect 12563 3638 12799 3674
rect 12563 3606 12665 3638
rect 12697 3606 12799 3638
rect 12563 3570 12799 3606
rect 12563 3538 12665 3570
rect 12697 3538 12799 3570
rect 12563 3502 12799 3538
rect 12563 3470 12665 3502
rect 12697 3470 12799 3502
rect 12563 3454 12799 3470
rect 12919 4318 13047 4334
rect 12919 4286 12967 4318
rect 12999 4286 13047 4318
rect 12919 4250 13047 4286
rect 12919 4218 12967 4250
rect 12999 4218 13047 4250
rect 12919 4182 13047 4218
rect 12919 4150 12967 4182
rect 12999 4150 13047 4182
rect 12919 4114 13047 4150
rect 12919 4082 12967 4114
rect 12999 4082 13047 4114
rect 12919 4046 13047 4082
rect 12919 4014 12967 4046
rect 12999 4014 13047 4046
rect 12919 3978 13047 4014
rect 12919 3946 12967 3978
rect 12999 3946 13047 3978
rect 12919 3910 13047 3946
rect 12919 3878 12967 3910
rect 12999 3878 13047 3910
rect 12919 3842 13047 3878
rect 12919 3810 12967 3842
rect 12999 3810 13047 3842
rect 12919 3774 13047 3810
rect 12919 3742 12967 3774
rect 12999 3742 13047 3774
rect 12919 3706 13047 3742
rect 12919 3674 12967 3706
rect 12999 3674 13047 3706
rect 12919 3638 13047 3674
rect 12919 3606 12967 3638
rect 12999 3606 13047 3638
rect 12919 3570 13047 3606
rect 12919 3538 12967 3570
rect 12999 3538 13047 3570
rect 12919 3502 13047 3538
rect 12919 3470 12967 3502
rect 12999 3470 13047 3502
rect 12919 3454 13047 3470
rect 13167 4318 13403 4334
rect 13167 4286 13269 4318
rect 13301 4286 13403 4318
rect 13167 4250 13403 4286
rect 13167 4218 13269 4250
rect 13301 4218 13403 4250
rect 13167 4182 13403 4218
rect 13167 4150 13269 4182
rect 13301 4150 13403 4182
rect 13167 4114 13403 4150
rect 13167 4082 13269 4114
rect 13301 4082 13403 4114
rect 13167 4046 13403 4082
rect 13167 4014 13269 4046
rect 13301 4014 13403 4046
rect 13167 3978 13403 4014
rect 13167 3946 13269 3978
rect 13301 3946 13403 3978
rect 13167 3910 13403 3946
rect 13167 3878 13269 3910
rect 13301 3878 13403 3910
rect 13167 3842 13403 3878
rect 13167 3810 13269 3842
rect 13301 3810 13403 3842
rect 13167 3774 13403 3810
rect 13167 3742 13269 3774
rect 13301 3742 13403 3774
rect 13167 3706 13403 3742
rect 13167 3674 13269 3706
rect 13301 3674 13403 3706
rect 13167 3638 13403 3674
rect 13167 3606 13269 3638
rect 13301 3606 13403 3638
rect 13167 3570 13403 3606
rect 13167 3538 13269 3570
rect 13301 3538 13403 3570
rect 13167 3502 13403 3538
rect 13167 3470 13269 3502
rect 13301 3470 13403 3502
rect 13167 3454 13403 3470
rect 13523 4318 13651 4334
rect 13523 4286 13571 4318
rect 13603 4286 13651 4318
rect 13523 4250 13651 4286
rect 13523 4218 13571 4250
rect 13603 4218 13651 4250
rect 13523 4182 13651 4218
rect 13523 4150 13571 4182
rect 13603 4150 13651 4182
rect 13523 4114 13651 4150
rect 13523 4082 13571 4114
rect 13603 4082 13651 4114
rect 13523 4046 13651 4082
rect 13523 4014 13571 4046
rect 13603 4014 13651 4046
rect 13523 3978 13651 4014
rect 13523 3946 13571 3978
rect 13603 3946 13651 3978
rect 13523 3910 13651 3946
rect 13523 3878 13571 3910
rect 13603 3878 13651 3910
rect 13523 3842 13651 3878
rect 13523 3810 13571 3842
rect 13603 3810 13651 3842
rect 13523 3774 13651 3810
rect 13523 3742 13571 3774
rect 13603 3742 13651 3774
rect 13523 3706 13651 3742
rect 13523 3674 13571 3706
rect 13603 3674 13651 3706
rect 13523 3638 13651 3674
rect 13523 3606 13571 3638
rect 13603 3606 13651 3638
rect 13523 3570 13651 3606
rect 13523 3538 13571 3570
rect 13603 3538 13651 3570
rect 13523 3502 13651 3538
rect 13523 3470 13571 3502
rect 13603 3470 13651 3502
rect 13523 3454 13651 3470
rect 13771 4318 14007 4334
rect 13771 4286 13873 4318
rect 13905 4286 14007 4318
rect 13771 4250 14007 4286
rect 13771 4218 13873 4250
rect 13905 4218 14007 4250
rect 13771 4182 14007 4218
rect 13771 4150 13873 4182
rect 13905 4150 14007 4182
rect 13771 4114 14007 4150
rect 13771 4082 13873 4114
rect 13905 4082 14007 4114
rect 13771 4046 14007 4082
rect 13771 4014 13873 4046
rect 13905 4014 14007 4046
rect 13771 3978 14007 4014
rect 13771 3946 13873 3978
rect 13905 3946 14007 3978
rect 13771 3910 14007 3946
rect 13771 3878 13873 3910
rect 13905 3878 14007 3910
rect 13771 3842 14007 3878
rect 13771 3810 13873 3842
rect 13905 3810 14007 3842
rect 13771 3774 14007 3810
rect 13771 3742 13873 3774
rect 13905 3742 14007 3774
rect 13771 3706 14007 3742
rect 13771 3674 13873 3706
rect 13905 3674 14007 3706
rect 13771 3638 14007 3674
rect 13771 3606 13873 3638
rect 13905 3606 14007 3638
rect 13771 3570 14007 3606
rect 13771 3538 13873 3570
rect 13905 3538 14007 3570
rect 13771 3502 14007 3538
rect 13771 3470 13873 3502
rect 13905 3470 14007 3502
rect 13771 3454 14007 3470
rect 14127 4318 14255 4334
rect 14127 4286 14175 4318
rect 14207 4286 14255 4318
rect 14127 4250 14255 4286
rect 14127 4218 14175 4250
rect 14207 4218 14255 4250
rect 14127 4182 14255 4218
rect 14127 4150 14175 4182
rect 14207 4150 14255 4182
rect 14127 4114 14255 4150
rect 14127 4082 14175 4114
rect 14207 4082 14255 4114
rect 14127 4046 14255 4082
rect 14127 4014 14175 4046
rect 14207 4014 14255 4046
rect 14127 3978 14255 4014
rect 14127 3946 14175 3978
rect 14207 3946 14255 3978
rect 14127 3910 14255 3946
rect 14127 3878 14175 3910
rect 14207 3878 14255 3910
rect 14127 3842 14255 3878
rect 14127 3810 14175 3842
rect 14207 3810 14255 3842
rect 14127 3774 14255 3810
rect 14127 3742 14175 3774
rect 14207 3742 14255 3774
rect 14127 3706 14255 3742
rect 14127 3674 14175 3706
rect 14207 3674 14255 3706
rect 14127 3638 14255 3674
rect 14127 3606 14175 3638
rect 14207 3606 14255 3638
rect 14127 3570 14255 3606
rect 14127 3538 14175 3570
rect 14207 3538 14255 3570
rect 14127 3502 14255 3538
rect 14127 3470 14175 3502
rect 14207 3470 14255 3502
rect 14127 3454 14255 3470
rect 14375 4318 14523 4334
rect 14375 4286 14477 4318
rect 14509 4286 14523 4318
rect 14375 4250 14523 4286
rect 14375 4218 14477 4250
rect 14509 4218 14523 4250
rect 14375 4182 14523 4218
rect 14375 4150 14477 4182
rect 14509 4150 14523 4182
rect 14375 4114 14523 4150
rect 14375 4082 14477 4114
rect 14509 4082 14523 4114
rect 14375 4046 14523 4082
rect 14375 4014 14477 4046
rect 14509 4014 14523 4046
rect 14375 3978 14523 4014
rect 14375 3946 14477 3978
rect 14509 3946 14523 3978
rect 14375 3910 14523 3946
rect 14375 3878 14477 3910
rect 14509 3878 14523 3910
rect 14375 3842 14523 3878
rect 14375 3810 14477 3842
rect 14509 3810 14523 3842
rect 14375 3774 14523 3810
rect 14375 3742 14477 3774
rect 14509 3742 14523 3774
rect 14375 3706 14523 3742
rect 14375 3674 14477 3706
rect 14509 3674 14523 3706
rect 14375 3638 14523 3674
rect 14375 3606 14477 3638
rect 14509 3606 14523 3638
rect 14375 3570 14523 3606
rect 14375 3538 14477 3570
rect 14509 3538 14523 3570
rect 14375 3502 14523 3538
rect 14375 3470 14477 3502
rect 14509 3470 14523 3502
rect 14375 3454 14523 3470
rect 1477 3350 1571 3366
rect 1477 3318 1491 3350
rect 1523 3318 1571 3350
rect 1477 3282 1571 3318
rect 1477 3250 1491 3282
rect 1523 3250 1571 3282
rect 1477 3214 1571 3250
rect 1477 3182 1491 3214
rect 1523 3182 1571 3214
rect 1477 3146 1571 3182
rect 1477 3114 1491 3146
rect 1523 3114 1571 3146
rect 1477 3078 1571 3114
rect 1477 3046 1491 3078
rect 1523 3046 1571 3078
rect 1477 3010 1571 3046
rect 1477 2978 1491 3010
rect 1523 2978 1571 3010
rect 1477 2942 1571 2978
rect 1477 2910 1491 2942
rect 1523 2910 1571 2942
rect 1477 2874 1571 2910
rect 1477 2842 1491 2874
rect 1523 2842 1571 2874
rect 1477 2806 1571 2842
rect 1477 2774 1491 2806
rect 1523 2774 1571 2806
rect 1477 2738 1571 2774
rect 1477 2706 1491 2738
rect 1523 2706 1571 2738
rect 1477 2670 1571 2706
rect 1477 2638 1491 2670
rect 1523 2638 1571 2670
rect 1477 2602 1571 2638
rect 1477 2570 1491 2602
rect 1523 2570 1571 2602
rect 1477 2534 1571 2570
rect 1477 2502 1491 2534
rect 1523 2502 1571 2534
rect 1477 2486 1571 2502
rect 1691 3350 1927 3366
rect 1691 3318 1793 3350
rect 1825 3318 1927 3350
rect 1691 3282 1927 3318
rect 1691 3250 1793 3282
rect 1825 3250 1927 3282
rect 1691 3214 1927 3250
rect 1691 3182 1793 3214
rect 1825 3182 1927 3214
rect 1691 3146 1927 3182
rect 1691 3114 1793 3146
rect 1825 3114 1927 3146
rect 1691 3078 1927 3114
rect 1691 3046 1793 3078
rect 1825 3046 1927 3078
rect 1691 3010 1927 3046
rect 1691 2978 1793 3010
rect 1825 2978 1927 3010
rect 1691 2942 1927 2978
rect 1691 2910 1793 2942
rect 1825 2910 1927 2942
rect 1691 2874 1927 2910
rect 1691 2842 1793 2874
rect 1825 2842 1927 2874
rect 1691 2806 1927 2842
rect 1691 2774 1793 2806
rect 1825 2774 1927 2806
rect 1691 2738 1927 2774
rect 1691 2706 1793 2738
rect 1825 2706 1927 2738
rect 1691 2670 1927 2706
rect 1691 2638 1793 2670
rect 1825 2638 1927 2670
rect 1691 2602 1927 2638
rect 1691 2570 1793 2602
rect 1825 2570 1927 2602
rect 1691 2534 1927 2570
rect 1691 2502 1793 2534
rect 1825 2502 1927 2534
rect 1691 2486 1927 2502
rect 2047 3350 2175 3366
rect 2047 3318 2095 3350
rect 2127 3318 2175 3350
rect 2047 3282 2175 3318
rect 2047 3250 2095 3282
rect 2127 3250 2175 3282
rect 2047 3214 2175 3250
rect 2047 3182 2095 3214
rect 2127 3182 2175 3214
rect 2047 3146 2175 3182
rect 2047 3114 2095 3146
rect 2127 3114 2175 3146
rect 2047 3078 2175 3114
rect 2047 3046 2095 3078
rect 2127 3046 2175 3078
rect 2047 3010 2175 3046
rect 2047 2978 2095 3010
rect 2127 2978 2175 3010
rect 2047 2942 2175 2978
rect 2047 2910 2095 2942
rect 2127 2910 2175 2942
rect 2047 2874 2175 2910
rect 2047 2842 2095 2874
rect 2127 2842 2175 2874
rect 2047 2806 2175 2842
rect 2047 2774 2095 2806
rect 2127 2774 2175 2806
rect 2047 2738 2175 2774
rect 2047 2706 2095 2738
rect 2127 2706 2175 2738
rect 2047 2670 2175 2706
rect 2047 2638 2095 2670
rect 2127 2638 2175 2670
rect 2047 2602 2175 2638
rect 2047 2570 2095 2602
rect 2127 2570 2175 2602
rect 2047 2534 2175 2570
rect 2047 2502 2095 2534
rect 2127 2502 2175 2534
rect 2047 2486 2175 2502
rect 2295 3350 2531 3366
rect 2295 3318 2397 3350
rect 2429 3318 2531 3350
rect 2295 3282 2531 3318
rect 2295 3250 2397 3282
rect 2429 3250 2531 3282
rect 2295 3214 2531 3250
rect 2295 3182 2397 3214
rect 2429 3182 2531 3214
rect 2295 3146 2531 3182
rect 2295 3114 2397 3146
rect 2429 3114 2531 3146
rect 2295 3078 2531 3114
rect 2295 3046 2397 3078
rect 2429 3046 2531 3078
rect 2295 3010 2531 3046
rect 2295 2978 2397 3010
rect 2429 2978 2531 3010
rect 2295 2942 2531 2978
rect 2295 2910 2397 2942
rect 2429 2910 2531 2942
rect 2295 2874 2531 2910
rect 2295 2842 2397 2874
rect 2429 2842 2531 2874
rect 2295 2806 2531 2842
rect 2295 2774 2397 2806
rect 2429 2774 2531 2806
rect 2295 2738 2531 2774
rect 2295 2706 2397 2738
rect 2429 2706 2531 2738
rect 2295 2670 2531 2706
rect 2295 2638 2397 2670
rect 2429 2638 2531 2670
rect 2295 2602 2531 2638
rect 2295 2570 2397 2602
rect 2429 2570 2531 2602
rect 2295 2534 2531 2570
rect 2295 2502 2397 2534
rect 2429 2502 2531 2534
rect 2295 2486 2531 2502
rect 2651 3350 2779 3366
rect 2651 3318 2699 3350
rect 2731 3318 2779 3350
rect 2651 3282 2779 3318
rect 2651 3250 2699 3282
rect 2731 3250 2779 3282
rect 2651 3214 2779 3250
rect 2651 3182 2699 3214
rect 2731 3182 2779 3214
rect 2651 3146 2779 3182
rect 2651 3114 2699 3146
rect 2731 3114 2779 3146
rect 2651 3078 2779 3114
rect 2651 3046 2699 3078
rect 2731 3046 2779 3078
rect 2651 3010 2779 3046
rect 2651 2978 2699 3010
rect 2731 2978 2779 3010
rect 2651 2942 2779 2978
rect 2651 2910 2699 2942
rect 2731 2910 2779 2942
rect 2651 2874 2779 2910
rect 2651 2842 2699 2874
rect 2731 2842 2779 2874
rect 2651 2806 2779 2842
rect 2651 2774 2699 2806
rect 2731 2774 2779 2806
rect 2651 2738 2779 2774
rect 2651 2706 2699 2738
rect 2731 2706 2779 2738
rect 2651 2670 2779 2706
rect 2651 2638 2699 2670
rect 2731 2638 2779 2670
rect 2651 2602 2779 2638
rect 2651 2570 2699 2602
rect 2731 2570 2779 2602
rect 2651 2534 2779 2570
rect 2651 2502 2699 2534
rect 2731 2502 2779 2534
rect 2651 2486 2779 2502
rect 2899 3350 3135 3366
rect 2899 3318 3001 3350
rect 3033 3318 3135 3350
rect 2899 3282 3135 3318
rect 2899 3250 3001 3282
rect 3033 3250 3135 3282
rect 2899 3214 3135 3250
rect 2899 3182 3001 3214
rect 3033 3182 3135 3214
rect 2899 3146 3135 3182
rect 2899 3114 3001 3146
rect 3033 3114 3135 3146
rect 2899 3078 3135 3114
rect 2899 3046 3001 3078
rect 3033 3046 3135 3078
rect 2899 3010 3135 3046
rect 2899 2978 3001 3010
rect 3033 2978 3135 3010
rect 2899 2942 3135 2978
rect 2899 2910 3001 2942
rect 3033 2910 3135 2942
rect 2899 2874 3135 2910
rect 2899 2842 3001 2874
rect 3033 2842 3135 2874
rect 2899 2806 3135 2842
rect 2899 2774 3001 2806
rect 3033 2774 3135 2806
rect 2899 2738 3135 2774
rect 2899 2706 3001 2738
rect 3033 2706 3135 2738
rect 2899 2670 3135 2706
rect 2899 2638 3001 2670
rect 3033 2638 3135 2670
rect 2899 2602 3135 2638
rect 2899 2570 3001 2602
rect 3033 2570 3135 2602
rect 2899 2534 3135 2570
rect 2899 2502 3001 2534
rect 3033 2502 3135 2534
rect 2899 2486 3135 2502
rect 3255 3350 3383 3366
rect 3255 3318 3303 3350
rect 3335 3318 3383 3350
rect 3255 3282 3383 3318
rect 3255 3250 3303 3282
rect 3335 3250 3383 3282
rect 3255 3214 3383 3250
rect 3255 3182 3303 3214
rect 3335 3182 3383 3214
rect 3255 3146 3383 3182
rect 3255 3114 3303 3146
rect 3335 3114 3383 3146
rect 3255 3078 3383 3114
rect 3255 3046 3303 3078
rect 3335 3046 3383 3078
rect 3255 3010 3383 3046
rect 3255 2978 3303 3010
rect 3335 2978 3383 3010
rect 3255 2942 3383 2978
rect 3255 2910 3303 2942
rect 3335 2910 3383 2942
rect 3255 2874 3383 2910
rect 3255 2842 3303 2874
rect 3335 2842 3383 2874
rect 3255 2806 3383 2842
rect 3255 2774 3303 2806
rect 3335 2774 3383 2806
rect 3255 2738 3383 2774
rect 3255 2706 3303 2738
rect 3335 2706 3383 2738
rect 3255 2670 3383 2706
rect 3255 2638 3303 2670
rect 3335 2638 3383 2670
rect 3255 2602 3383 2638
rect 3255 2570 3303 2602
rect 3335 2570 3383 2602
rect 3255 2534 3383 2570
rect 3255 2502 3303 2534
rect 3335 2502 3383 2534
rect 3255 2486 3383 2502
rect 3503 3350 3739 3366
rect 3503 3318 3605 3350
rect 3637 3318 3739 3350
rect 3503 3282 3739 3318
rect 3503 3250 3605 3282
rect 3637 3250 3739 3282
rect 3503 3214 3739 3250
rect 3503 3182 3605 3214
rect 3637 3182 3739 3214
rect 3503 3146 3739 3182
rect 3503 3114 3605 3146
rect 3637 3114 3739 3146
rect 3503 3078 3739 3114
rect 3503 3046 3605 3078
rect 3637 3046 3739 3078
rect 3503 3010 3739 3046
rect 3503 2978 3605 3010
rect 3637 2978 3739 3010
rect 3503 2942 3739 2978
rect 3503 2910 3605 2942
rect 3637 2910 3739 2942
rect 3503 2874 3739 2910
rect 3503 2842 3605 2874
rect 3637 2842 3739 2874
rect 3503 2806 3739 2842
rect 3503 2774 3605 2806
rect 3637 2774 3739 2806
rect 3503 2738 3739 2774
rect 3503 2706 3605 2738
rect 3637 2706 3739 2738
rect 3503 2670 3739 2706
rect 3503 2638 3605 2670
rect 3637 2638 3739 2670
rect 3503 2602 3739 2638
rect 3503 2570 3605 2602
rect 3637 2570 3739 2602
rect 3503 2534 3739 2570
rect 3503 2502 3605 2534
rect 3637 2502 3739 2534
rect 3503 2486 3739 2502
rect 3859 3350 3987 3366
rect 3859 3318 3907 3350
rect 3939 3318 3987 3350
rect 3859 3282 3987 3318
rect 3859 3250 3907 3282
rect 3939 3250 3987 3282
rect 3859 3214 3987 3250
rect 3859 3182 3907 3214
rect 3939 3182 3987 3214
rect 3859 3146 3987 3182
rect 3859 3114 3907 3146
rect 3939 3114 3987 3146
rect 3859 3078 3987 3114
rect 3859 3046 3907 3078
rect 3939 3046 3987 3078
rect 3859 3010 3987 3046
rect 3859 2978 3907 3010
rect 3939 2978 3987 3010
rect 3859 2942 3987 2978
rect 3859 2910 3907 2942
rect 3939 2910 3987 2942
rect 3859 2874 3987 2910
rect 3859 2842 3907 2874
rect 3939 2842 3987 2874
rect 3859 2806 3987 2842
rect 3859 2774 3907 2806
rect 3939 2774 3987 2806
rect 3859 2738 3987 2774
rect 3859 2706 3907 2738
rect 3939 2706 3987 2738
rect 3859 2670 3987 2706
rect 3859 2638 3907 2670
rect 3939 2638 3987 2670
rect 3859 2602 3987 2638
rect 3859 2570 3907 2602
rect 3939 2570 3987 2602
rect 3859 2534 3987 2570
rect 3859 2502 3907 2534
rect 3939 2502 3987 2534
rect 3859 2486 3987 2502
rect 4107 3350 4343 3366
rect 4107 3318 4209 3350
rect 4241 3318 4343 3350
rect 4107 3282 4343 3318
rect 4107 3250 4209 3282
rect 4241 3250 4343 3282
rect 4107 3214 4343 3250
rect 4107 3182 4209 3214
rect 4241 3182 4343 3214
rect 4107 3146 4343 3182
rect 4107 3114 4209 3146
rect 4241 3114 4343 3146
rect 4107 3078 4343 3114
rect 4107 3046 4209 3078
rect 4241 3046 4343 3078
rect 4107 3010 4343 3046
rect 4107 2978 4209 3010
rect 4241 2978 4343 3010
rect 4107 2942 4343 2978
rect 4107 2910 4209 2942
rect 4241 2910 4343 2942
rect 4107 2874 4343 2910
rect 4107 2842 4209 2874
rect 4241 2842 4343 2874
rect 4107 2806 4343 2842
rect 4107 2774 4209 2806
rect 4241 2774 4343 2806
rect 4107 2738 4343 2774
rect 4107 2706 4209 2738
rect 4241 2706 4343 2738
rect 4107 2670 4343 2706
rect 4107 2638 4209 2670
rect 4241 2638 4343 2670
rect 4107 2602 4343 2638
rect 4107 2570 4209 2602
rect 4241 2570 4343 2602
rect 4107 2534 4343 2570
rect 4107 2502 4209 2534
rect 4241 2502 4343 2534
rect 4107 2486 4343 2502
rect 4463 3350 4591 3366
rect 4463 3318 4511 3350
rect 4543 3318 4591 3350
rect 4463 3282 4591 3318
rect 4463 3250 4511 3282
rect 4543 3250 4591 3282
rect 4463 3214 4591 3250
rect 4463 3182 4511 3214
rect 4543 3182 4591 3214
rect 4463 3146 4591 3182
rect 4463 3114 4511 3146
rect 4543 3114 4591 3146
rect 4463 3078 4591 3114
rect 4463 3046 4511 3078
rect 4543 3046 4591 3078
rect 4463 3010 4591 3046
rect 4463 2978 4511 3010
rect 4543 2978 4591 3010
rect 4463 2942 4591 2978
rect 4463 2910 4511 2942
rect 4543 2910 4591 2942
rect 4463 2874 4591 2910
rect 4463 2842 4511 2874
rect 4543 2842 4591 2874
rect 4463 2806 4591 2842
rect 4463 2774 4511 2806
rect 4543 2774 4591 2806
rect 4463 2738 4591 2774
rect 4463 2706 4511 2738
rect 4543 2706 4591 2738
rect 4463 2670 4591 2706
rect 4463 2638 4511 2670
rect 4543 2638 4591 2670
rect 4463 2602 4591 2638
rect 4463 2570 4511 2602
rect 4543 2570 4591 2602
rect 4463 2534 4591 2570
rect 4463 2502 4511 2534
rect 4543 2502 4591 2534
rect 4463 2486 4591 2502
rect 4711 3350 4947 3366
rect 4711 3318 4813 3350
rect 4845 3318 4947 3350
rect 4711 3282 4947 3318
rect 4711 3250 4813 3282
rect 4845 3250 4947 3282
rect 4711 3214 4947 3250
rect 4711 3182 4813 3214
rect 4845 3182 4947 3214
rect 4711 3146 4947 3182
rect 4711 3114 4813 3146
rect 4845 3114 4947 3146
rect 4711 3078 4947 3114
rect 4711 3046 4813 3078
rect 4845 3046 4947 3078
rect 4711 3010 4947 3046
rect 4711 2978 4813 3010
rect 4845 2978 4947 3010
rect 4711 2942 4947 2978
rect 4711 2910 4813 2942
rect 4845 2910 4947 2942
rect 4711 2874 4947 2910
rect 4711 2842 4813 2874
rect 4845 2842 4947 2874
rect 4711 2806 4947 2842
rect 4711 2774 4813 2806
rect 4845 2774 4947 2806
rect 4711 2738 4947 2774
rect 4711 2706 4813 2738
rect 4845 2706 4947 2738
rect 4711 2670 4947 2706
rect 4711 2638 4813 2670
rect 4845 2638 4947 2670
rect 4711 2602 4947 2638
rect 4711 2570 4813 2602
rect 4845 2570 4947 2602
rect 4711 2534 4947 2570
rect 4711 2502 4813 2534
rect 4845 2502 4947 2534
rect 4711 2486 4947 2502
rect 5067 3350 5195 3366
rect 5067 3318 5115 3350
rect 5147 3318 5195 3350
rect 5067 3282 5195 3318
rect 5067 3250 5115 3282
rect 5147 3250 5195 3282
rect 5067 3214 5195 3250
rect 5067 3182 5115 3214
rect 5147 3182 5195 3214
rect 5067 3146 5195 3182
rect 5067 3114 5115 3146
rect 5147 3114 5195 3146
rect 5067 3078 5195 3114
rect 5067 3046 5115 3078
rect 5147 3046 5195 3078
rect 5067 3010 5195 3046
rect 5067 2978 5115 3010
rect 5147 2978 5195 3010
rect 5067 2942 5195 2978
rect 5067 2910 5115 2942
rect 5147 2910 5195 2942
rect 5067 2874 5195 2910
rect 5067 2842 5115 2874
rect 5147 2842 5195 2874
rect 5067 2806 5195 2842
rect 5067 2774 5115 2806
rect 5147 2774 5195 2806
rect 5067 2738 5195 2774
rect 5067 2706 5115 2738
rect 5147 2706 5195 2738
rect 5067 2670 5195 2706
rect 5067 2638 5115 2670
rect 5147 2638 5195 2670
rect 5067 2602 5195 2638
rect 5067 2570 5115 2602
rect 5147 2570 5195 2602
rect 5067 2534 5195 2570
rect 5067 2502 5115 2534
rect 5147 2502 5195 2534
rect 5067 2486 5195 2502
rect 5315 3350 5551 3366
rect 5315 3318 5417 3350
rect 5449 3318 5551 3350
rect 5315 3282 5551 3318
rect 5315 3250 5417 3282
rect 5449 3250 5551 3282
rect 5315 3214 5551 3250
rect 5315 3182 5417 3214
rect 5449 3182 5551 3214
rect 5315 3146 5551 3182
rect 5315 3114 5417 3146
rect 5449 3114 5551 3146
rect 5315 3078 5551 3114
rect 5315 3046 5417 3078
rect 5449 3046 5551 3078
rect 5315 3010 5551 3046
rect 5315 2978 5417 3010
rect 5449 2978 5551 3010
rect 5315 2942 5551 2978
rect 5315 2910 5417 2942
rect 5449 2910 5551 2942
rect 5315 2874 5551 2910
rect 5315 2842 5417 2874
rect 5449 2842 5551 2874
rect 5315 2806 5551 2842
rect 5315 2774 5417 2806
rect 5449 2774 5551 2806
rect 5315 2738 5551 2774
rect 5315 2706 5417 2738
rect 5449 2706 5551 2738
rect 5315 2670 5551 2706
rect 5315 2638 5417 2670
rect 5449 2638 5551 2670
rect 5315 2602 5551 2638
rect 5315 2570 5417 2602
rect 5449 2570 5551 2602
rect 5315 2534 5551 2570
rect 5315 2502 5417 2534
rect 5449 2502 5551 2534
rect 5315 2486 5551 2502
rect 5671 3350 5799 3366
rect 5671 3318 5719 3350
rect 5751 3318 5799 3350
rect 5671 3282 5799 3318
rect 5671 3250 5719 3282
rect 5751 3250 5799 3282
rect 5671 3214 5799 3250
rect 5671 3182 5719 3214
rect 5751 3182 5799 3214
rect 5671 3146 5799 3182
rect 5671 3114 5719 3146
rect 5751 3114 5799 3146
rect 5671 3078 5799 3114
rect 5671 3046 5719 3078
rect 5751 3046 5799 3078
rect 5671 3010 5799 3046
rect 5671 2978 5719 3010
rect 5751 2978 5799 3010
rect 5671 2942 5799 2978
rect 5671 2910 5719 2942
rect 5751 2910 5799 2942
rect 5671 2874 5799 2910
rect 5671 2842 5719 2874
rect 5751 2842 5799 2874
rect 5671 2806 5799 2842
rect 5671 2774 5719 2806
rect 5751 2774 5799 2806
rect 5671 2738 5799 2774
rect 5671 2706 5719 2738
rect 5751 2706 5799 2738
rect 5671 2670 5799 2706
rect 5671 2638 5719 2670
rect 5751 2638 5799 2670
rect 5671 2602 5799 2638
rect 5671 2570 5719 2602
rect 5751 2570 5799 2602
rect 5671 2534 5799 2570
rect 5671 2502 5719 2534
rect 5751 2502 5799 2534
rect 5671 2486 5799 2502
rect 5919 3350 6155 3366
rect 5919 3318 6021 3350
rect 6053 3318 6155 3350
rect 5919 3282 6155 3318
rect 5919 3250 6021 3282
rect 6053 3250 6155 3282
rect 5919 3214 6155 3250
rect 5919 3182 6021 3214
rect 6053 3182 6155 3214
rect 5919 3146 6155 3182
rect 5919 3114 6021 3146
rect 6053 3114 6155 3146
rect 5919 3078 6155 3114
rect 5919 3046 6021 3078
rect 6053 3046 6155 3078
rect 5919 3010 6155 3046
rect 5919 2978 6021 3010
rect 6053 2978 6155 3010
rect 5919 2942 6155 2978
rect 5919 2910 6021 2942
rect 6053 2910 6155 2942
rect 5919 2874 6155 2910
rect 5919 2842 6021 2874
rect 6053 2842 6155 2874
rect 5919 2806 6155 2842
rect 5919 2774 6021 2806
rect 6053 2774 6155 2806
rect 5919 2738 6155 2774
rect 5919 2706 6021 2738
rect 6053 2706 6155 2738
rect 5919 2670 6155 2706
rect 5919 2638 6021 2670
rect 6053 2638 6155 2670
rect 5919 2602 6155 2638
rect 5919 2570 6021 2602
rect 6053 2570 6155 2602
rect 5919 2534 6155 2570
rect 5919 2502 6021 2534
rect 6053 2502 6155 2534
rect 5919 2486 6155 2502
rect 6275 3350 6403 3366
rect 6275 3318 6323 3350
rect 6355 3318 6403 3350
rect 6275 3282 6403 3318
rect 6275 3250 6323 3282
rect 6355 3250 6403 3282
rect 6275 3214 6403 3250
rect 6275 3182 6323 3214
rect 6355 3182 6403 3214
rect 6275 3146 6403 3182
rect 6275 3114 6323 3146
rect 6355 3114 6403 3146
rect 6275 3078 6403 3114
rect 6275 3046 6323 3078
rect 6355 3046 6403 3078
rect 6275 3010 6403 3046
rect 6275 2978 6323 3010
rect 6355 2978 6403 3010
rect 6275 2942 6403 2978
rect 6275 2910 6323 2942
rect 6355 2910 6403 2942
rect 6275 2874 6403 2910
rect 6275 2842 6323 2874
rect 6355 2842 6403 2874
rect 6275 2806 6403 2842
rect 6275 2774 6323 2806
rect 6355 2774 6403 2806
rect 6275 2738 6403 2774
rect 6275 2706 6323 2738
rect 6355 2706 6403 2738
rect 6275 2670 6403 2706
rect 6275 2638 6323 2670
rect 6355 2638 6403 2670
rect 6275 2602 6403 2638
rect 6275 2570 6323 2602
rect 6355 2570 6403 2602
rect 6275 2534 6403 2570
rect 6275 2502 6323 2534
rect 6355 2502 6403 2534
rect 6275 2486 6403 2502
rect 6523 3350 6759 3366
rect 6523 3318 6625 3350
rect 6657 3318 6759 3350
rect 6523 3282 6759 3318
rect 6523 3250 6625 3282
rect 6657 3250 6759 3282
rect 6523 3214 6759 3250
rect 6523 3182 6625 3214
rect 6657 3182 6759 3214
rect 6523 3146 6759 3182
rect 6523 3114 6625 3146
rect 6657 3114 6759 3146
rect 6523 3078 6759 3114
rect 6523 3046 6625 3078
rect 6657 3046 6759 3078
rect 6523 3010 6759 3046
rect 6523 2978 6625 3010
rect 6657 2978 6759 3010
rect 6523 2942 6759 2978
rect 6523 2910 6625 2942
rect 6657 2910 6759 2942
rect 6523 2874 6759 2910
rect 6523 2842 6625 2874
rect 6657 2842 6759 2874
rect 6523 2806 6759 2842
rect 6523 2774 6625 2806
rect 6657 2774 6759 2806
rect 6523 2738 6759 2774
rect 6523 2706 6625 2738
rect 6657 2706 6759 2738
rect 6523 2670 6759 2706
rect 6523 2638 6625 2670
rect 6657 2638 6759 2670
rect 6523 2602 6759 2638
rect 6523 2570 6625 2602
rect 6657 2570 6759 2602
rect 6523 2534 6759 2570
rect 6523 2502 6625 2534
rect 6657 2502 6759 2534
rect 6523 2486 6759 2502
rect 6879 3350 7007 3366
rect 6879 3318 6927 3350
rect 6959 3318 7007 3350
rect 6879 3282 7007 3318
rect 6879 3250 6927 3282
rect 6959 3250 7007 3282
rect 6879 3214 7007 3250
rect 6879 3182 6927 3214
rect 6959 3182 7007 3214
rect 6879 3146 7007 3182
rect 6879 3114 6927 3146
rect 6959 3114 7007 3146
rect 6879 3078 7007 3114
rect 6879 3046 6927 3078
rect 6959 3046 7007 3078
rect 6879 3010 7007 3046
rect 6879 2978 6927 3010
rect 6959 2978 7007 3010
rect 6879 2942 7007 2978
rect 6879 2910 6927 2942
rect 6959 2910 7007 2942
rect 6879 2874 7007 2910
rect 6879 2842 6927 2874
rect 6959 2842 7007 2874
rect 6879 2806 7007 2842
rect 6879 2774 6927 2806
rect 6959 2774 7007 2806
rect 6879 2738 7007 2774
rect 6879 2706 6927 2738
rect 6959 2706 7007 2738
rect 6879 2670 7007 2706
rect 6879 2638 6927 2670
rect 6959 2638 7007 2670
rect 6879 2602 7007 2638
rect 6879 2570 6927 2602
rect 6959 2570 7007 2602
rect 6879 2534 7007 2570
rect 6879 2502 6927 2534
rect 6959 2502 7007 2534
rect 6879 2486 7007 2502
rect 7127 3350 7363 3366
rect 7127 3318 7229 3350
rect 7261 3318 7363 3350
rect 7127 3282 7363 3318
rect 7127 3250 7229 3282
rect 7261 3250 7363 3282
rect 7127 3214 7363 3250
rect 7127 3182 7229 3214
rect 7261 3182 7363 3214
rect 7127 3146 7363 3182
rect 7127 3114 7229 3146
rect 7261 3114 7363 3146
rect 7127 3078 7363 3114
rect 7127 3046 7229 3078
rect 7261 3046 7363 3078
rect 7127 3010 7363 3046
rect 7127 2978 7229 3010
rect 7261 2978 7363 3010
rect 7127 2942 7363 2978
rect 7127 2910 7229 2942
rect 7261 2910 7363 2942
rect 7127 2874 7363 2910
rect 7127 2842 7229 2874
rect 7261 2842 7363 2874
rect 7127 2806 7363 2842
rect 7127 2774 7229 2806
rect 7261 2774 7363 2806
rect 7127 2738 7363 2774
rect 7127 2706 7229 2738
rect 7261 2706 7363 2738
rect 7127 2670 7363 2706
rect 7127 2638 7229 2670
rect 7261 2638 7363 2670
rect 7127 2602 7363 2638
rect 7127 2570 7229 2602
rect 7261 2570 7363 2602
rect 7127 2534 7363 2570
rect 7127 2502 7229 2534
rect 7261 2502 7363 2534
rect 7127 2486 7363 2502
rect 7483 3350 7611 3366
rect 7483 3318 7531 3350
rect 7563 3318 7611 3350
rect 7483 3282 7611 3318
rect 7483 3250 7531 3282
rect 7563 3250 7611 3282
rect 7483 3214 7611 3250
rect 7483 3182 7531 3214
rect 7563 3182 7611 3214
rect 7483 3146 7611 3182
rect 7483 3114 7531 3146
rect 7563 3114 7611 3146
rect 7483 3078 7611 3114
rect 7483 3046 7531 3078
rect 7563 3046 7611 3078
rect 7483 3010 7611 3046
rect 7483 2978 7531 3010
rect 7563 2978 7611 3010
rect 7483 2942 7611 2978
rect 7483 2910 7531 2942
rect 7563 2910 7611 2942
rect 7483 2874 7611 2910
rect 7483 2842 7531 2874
rect 7563 2842 7611 2874
rect 7483 2806 7611 2842
rect 7483 2774 7531 2806
rect 7563 2774 7611 2806
rect 7483 2738 7611 2774
rect 7483 2706 7531 2738
rect 7563 2706 7611 2738
rect 7483 2670 7611 2706
rect 7483 2638 7531 2670
rect 7563 2638 7611 2670
rect 7483 2602 7611 2638
rect 7483 2570 7531 2602
rect 7563 2570 7611 2602
rect 7483 2534 7611 2570
rect 7483 2502 7531 2534
rect 7563 2502 7611 2534
rect 7483 2486 7611 2502
rect 7731 3350 7967 3366
rect 7731 3318 7833 3350
rect 7865 3318 7967 3350
rect 7731 3282 7967 3318
rect 7731 3250 7833 3282
rect 7865 3250 7967 3282
rect 7731 3214 7967 3250
rect 7731 3182 7833 3214
rect 7865 3182 7967 3214
rect 7731 3146 7967 3182
rect 7731 3114 7833 3146
rect 7865 3114 7967 3146
rect 7731 3078 7967 3114
rect 7731 3046 7833 3078
rect 7865 3046 7967 3078
rect 7731 3010 7967 3046
rect 7731 2978 7833 3010
rect 7865 2978 7967 3010
rect 7731 2942 7967 2978
rect 7731 2910 7833 2942
rect 7865 2910 7967 2942
rect 7731 2874 7967 2910
rect 7731 2842 7833 2874
rect 7865 2842 7967 2874
rect 7731 2806 7967 2842
rect 7731 2774 7833 2806
rect 7865 2774 7967 2806
rect 7731 2738 7967 2774
rect 7731 2706 7833 2738
rect 7865 2706 7967 2738
rect 7731 2670 7967 2706
rect 7731 2638 7833 2670
rect 7865 2638 7967 2670
rect 7731 2602 7967 2638
rect 7731 2570 7833 2602
rect 7865 2570 7967 2602
rect 7731 2534 7967 2570
rect 7731 2502 7833 2534
rect 7865 2502 7967 2534
rect 7731 2486 7967 2502
rect 8087 3350 8215 3366
rect 8087 3318 8135 3350
rect 8167 3318 8215 3350
rect 8087 3282 8215 3318
rect 8087 3250 8135 3282
rect 8167 3250 8215 3282
rect 8087 3214 8215 3250
rect 8087 3182 8135 3214
rect 8167 3182 8215 3214
rect 8087 3146 8215 3182
rect 8087 3114 8135 3146
rect 8167 3114 8215 3146
rect 8087 3078 8215 3114
rect 8087 3046 8135 3078
rect 8167 3046 8215 3078
rect 8087 3010 8215 3046
rect 8087 2978 8135 3010
rect 8167 2978 8215 3010
rect 8087 2942 8215 2978
rect 8087 2910 8135 2942
rect 8167 2910 8215 2942
rect 8087 2874 8215 2910
rect 8087 2842 8135 2874
rect 8167 2842 8215 2874
rect 8087 2806 8215 2842
rect 8087 2774 8135 2806
rect 8167 2774 8215 2806
rect 8087 2738 8215 2774
rect 8087 2706 8135 2738
rect 8167 2706 8215 2738
rect 8087 2670 8215 2706
rect 8087 2638 8135 2670
rect 8167 2638 8215 2670
rect 8087 2602 8215 2638
rect 8087 2570 8135 2602
rect 8167 2570 8215 2602
rect 8087 2534 8215 2570
rect 8087 2502 8135 2534
rect 8167 2502 8215 2534
rect 8087 2486 8215 2502
rect 8335 3350 8571 3366
rect 8335 3318 8437 3350
rect 8469 3318 8571 3350
rect 8335 3282 8571 3318
rect 8335 3250 8437 3282
rect 8469 3250 8571 3282
rect 8335 3214 8571 3250
rect 8335 3182 8437 3214
rect 8469 3182 8571 3214
rect 8335 3146 8571 3182
rect 8335 3114 8437 3146
rect 8469 3114 8571 3146
rect 8335 3078 8571 3114
rect 8335 3046 8437 3078
rect 8469 3046 8571 3078
rect 8335 3010 8571 3046
rect 8335 2978 8437 3010
rect 8469 2978 8571 3010
rect 8335 2942 8571 2978
rect 8335 2910 8437 2942
rect 8469 2910 8571 2942
rect 8335 2874 8571 2910
rect 8335 2842 8437 2874
rect 8469 2842 8571 2874
rect 8335 2806 8571 2842
rect 8335 2774 8437 2806
rect 8469 2774 8571 2806
rect 8335 2738 8571 2774
rect 8335 2706 8437 2738
rect 8469 2706 8571 2738
rect 8335 2670 8571 2706
rect 8335 2638 8437 2670
rect 8469 2638 8571 2670
rect 8335 2602 8571 2638
rect 8335 2570 8437 2602
rect 8469 2570 8571 2602
rect 8335 2534 8571 2570
rect 8335 2502 8437 2534
rect 8469 2502 8571 2534
rect 8335 2486 8571 2502
rect 8691 3350 8819 3366
rect 8691 3318 8739 3350
rect 8771 3318 8819 3350
rect 8691 3282 8819 3318
rect 8691 3250 8739 3282
rect 8771 3250 8819 3282
rect 8691 3214 8819 3250
rect 8691 3182 8739 3214
rect 8771 3182 8819 3214
rect 8691 3146 8819 3182
rect 8691 3114 8739 3146
rect 8771 3114 8819 3146
rect 8691 3078 8819 3114
rect 8691 3046 8739 3078
rect 8771 3046 8819 3078
rect 8691 3010 8819 3046
rect 8691 2978 8739 3010
rect 8771 2978 8819 3010
rect 8691 2942 8819 2978
rect 8691 2910 8739 2942
rect 8771 2910 8819 2942
rect 8691 2874 8819 2910
rect 8691 2842 8739 2874
rect 8771 2842 8819 2874
rect 8691 2806 8819 2842
rect 8691 2774 8739 2806
rect 8771 2774 8819 2806
rect 8691 2738 8819 2774
rect 8691 2706 8739 2738
rect 8771 2706 8819 2738
rect 8691 2670 8819 2706
rect 8691 2638 8739 2670
rect 8771 2638 8819 2670
rect 8691 2602 8819 2638
rect 8691 2570 8739 2602
rect 8771 2570 8819 2602
rect 8691 2534 8819 2570
rect 8691 2502 8739 2534
rect 8771 2502 8819 2534
rect 8691 2486 8819 2502
rect 8939 3350 9175 3366
rect 8939 3318 9041 3350
rect 9073 3318 9175 3350
rect 8939 3282 9175 3318
rect 8939 3250 9041 3282
rect 9073 3250 9175 3282
rect 8939 3214 9175 3250
rect 8939 3182 9041 3214
rect 9073 3182 9175 3214
rect 8939 3146 9175 3182
rect 8939 3114 9041 3146
rect 9073 3114 9175 3146
rect 8939 3078 9175 3114
rect 8939 3046 9041 3078
rect 9073 3046 9175 3078
rect 8939 3010 9175 3046
rect 8939 2978 9041 3010
rect 9073 2978 9175 3010
rect 8939 2942 9175 2978
rect 8939 2910 9041 2942
rect 9073 2910 9175 2942
rect 8939 2874 9175 2910
rect 8939 2842 9041 2874
rect 9073 2842 9175 2874
rect 8939 2806 9175 2842
rect 8939 2774 9041 2806
rect 9073 2774 9175 2806
rect 8939 2738 9175 2774
rect 8939 2706 9041 2738
rect 9073 2706 9175 2738
rect 8939 2670 9175 2706
rect 8939 2638 9041 2670
rect 9073 2638 9175 2670
rect 8939 2602 9175 2638
rect 8939 2570 9041 2602
rect 9073 2570 9175 2602
rect 8939 2534 9175 2570
rect 8939 2502 9041 2534
rect 9073 2502 9175 2534
rect 8939 2486 9175 2502
rect 9295 3350 9423 3366
rect 9295 3318 9343 3350
rect 9375 3318 9423 3350
rect 9295 3282 9423 3318
rect 9295 3250 9343 3282
rect 9375 3250 9423 3282
rect 9295 3214 9423 3250
rect 9295 3182 9343 3214
rect 9375 3182 9423 3214
rect 9295 3146 9423 3182
rect 9295 3114 9343 3146
rect 9375 3114 9423 3146
rect 9295 3078 9423 3114
rect 9295 3046 9343 3078
rect 9375 3046 9423 3078
rect 9295 3010 9423 3046
rect 9295 2978 9343 3010
rect 9375 2978 9423 3010
rect 9295 2942 9423 2978
rect 9295 2910 9343 2942
rect 9375 2910 9423 2942
rect 9295 2874 9423 2910
rect 9295 2842 9343 2874
rect 9375 2842 9423 2874
rect 9295 2806 9423 2842
rect 9295 2774 9343 2806
rect 9375 2774 9423 2806
rect 9295 2738 9423 2774
rect 9295 2706 9343 2738
rect 9375 2706 9423 2738
rect 9295 2670 9423 2706
rect 9295 2638 9343 2670
rect 9375 2638 9423 2670
rect 9295 2602 9423 2638
rect 9295 2570 9343 2602
rect 9375 2570 9423 2602
rect 9295 2534 9423 2570
rect 9295 2502 9343 2534
rect 9375 2502 9423 2534
rect 9295 2486 9423 2502
rect 9543 3350 9779 3366
rect 9543 3318 9645 3350
rect 9677 3318 9779 3350
rect 9543 3282 9779 3318
rect 9543 3250 9645 3282
rect 9677 3250 9779 3282
rect 9543 3214 9779 3250
rect 9543 3182 9645 3214
rect 9677 3182 9779 3214
rect 9543 3146 9779 3182
rect 9543 3114 9645 3146
rect 9677 3114 9779 3146
rect 9543 3078 9779 3114
rect 9543 3046 9645 3078
rect 9677 3046 9779 3078
rect 9543 3010 9779 3046
rect 9543 2978 9645 3010
rect 9677 2978 9779 3010
rect 9543 2942 9779 2978
rect 9543 2910 9645 2942
rect 9677 2910 9779 2942
rect 9543 2874 9779 2910
rect 9543 2842 9645 2874
rect 9677 2842 9779 2874
rect 9543 2806 9779 2842
rect 9543 2774 9645 2806
rect 9677 2774 9779 2806
rect 9543 2738 9779 2774
rect 9543 2706 9645 2738
rect 9677 2706 9779 2738
rect 9543 2670 9779 2706
rect 9543 2638 9645 2670
rect 9677 2638 9779 2670
rect 9543 2602 9779 2638
rect 9543 2570 9645 2602
rect 9677 2570 9779 2602
rect 9543 2534 9779 2570
rect 9543 2502 9645 2534
rect 9677 2502 9779 2534
rect 9543 2486 9779 2502
rect 9899 3350 10027 3366
rect 9899 3318 9947 3350
rect 9979 3318 10027 3350
rect 9899 3282 10027 3318
rect 9899 3250 9947 3282
rect 9979 3250 10027 3282
rect 9899 3214 10027 3250
rect 9899 3182 9947 3214
rect 9979 3182 10027 3214
rect 9899 3146 10027 3182
rect 9899 3114 9947 3146
rect 9979 3114 10027 3146
rect 9899 3078 10027 3114
rect 9899 3046 9947 3078
rect 9979 3046 10027 3078
rect 9899 3010 10027 3046
rect 9899 2978 9947 3010
rect 9979 2978 10027 3010
rect 9899 2942 10027 2978
rect 9899 2910 9947 2942
rect 9979 2910 10027 2942
rect 9899 2874 10027 2910
rect 9899 2842 9947 2874
rect 9979 2842 10027 2874
rect 9899 2806 10027 2842
rect 9899 2774 9947 2806
rect 9979 2774 10027 2806
rect 9899 2738 10027 2774
rect 9899 2706 9947 2738
rect 9979 2706 10027 2738
rect 9899 2670 10027 2706
rect 9899 2638 9947 2670
rect 9979 2638 10027 2670
rect 9899 2602 10027 2638
rect 9899 2570 9947 2602
rect 9979 2570 10027 2602
rect 9899 2534 10027 2570
rect 9899 2502 9947 2534
rect 9979 2502 10027 2534
rect 9899 2486 10027 2502
rect 10147 3350 10383 3366
rect 10147 3318 10249 3350
rect 10281 3318 10383 3350
rect 10147 3282 10383 3318
rect 10147 3250 10249 3282
rect 10281 3250 10383 3282
rect 10147 3214 10383 3250
rect 10147 3182 10249 3214
rect 10281 3182 10383 3214
rect 10147 3146 10383 3182
rect 10147 3114 10249 3146
rect 10281 3114 10383 3146
rect 10147 3078 10383 3114
rect 10147 3046 10249 3078
rect 10281 3046 10383 3078
rect 10147 3010 10383 3046
rect 10147 2978 10249 3010
rect 10281 2978 10383 3010
rect 10147 2942 10383 2978
rect 10147 2910 10249 2942
rect 10281 2910 10383 2942
rect 10147 2874 10383 2910
rect 10147 2842 10249 2874
rect 10281 2842 10383 2874
rect 10147 2806 10383 2842
rect 10147 2774 10249 2806
rect 10281 2774 10383 2806
rect 10147 2738 10383 2774
rect 10147 2706 10249 2738
rect 10281 2706 10383 2738
rect 10147 2670 10383 2706
rect 10147 2638 10249 2670
rect 10281 2638 10383 2670
rect 10147 2602 10383 2638
rect 10147 2570 10249 2602
rect 10281 2570 10383 2602
rect 10147 2534 10383 2570
rect 10147 2502 10249 2534
rect 10281 2502 10383 2534
rect 10147 2486 10383 2502
rect 10503 3350 10631 3366
rect 10503 3318 10551 3350
rect 10583 3318 10631 3350
rect 10503 3282 10631 3318
rect 10503 3250 10551 3282
rect 10583 3250 10631 3282
rect 10503 3214 10631 3250
rect 10503 3182 10551 3214
rect 10583 3182 10631 3214
rect 10503 3146 10631 3182
rect 10503 3114 10551 3146
rect 10583 3114 10631 3146
rect 10503 3078 10631 3114
rect 10503 3046 10551 3078
rect 10583 3046 10631 3078
rect 10503 3010 10631 3046
rect 10503 2978 10551 3010
rect 10583 2978 10631 3010
rect 10503 2942 10631 2978
rect 10503 2910 10551 2942
rect 10583 2910 10631 2942
rect 10503 2874 10631 2910
rect 10503 2842 10551 2874
rect 10583 2842 10631 2874
rect 10503 2806 10631 2842
rect 10503 2774 10551 2806
rect 10583 2774 10631 2806
rect 10503 2738 10631 2774
rect 10503 2706 10551 2738
rect 10583 2706 10631 2738
rect 10503 2670 10631 2706
rect 10503 2638 10551 2670
rect 10583 2638 10631 2670
rect 10503 2602 10631 2638
rect 10503 2570 10551 2602
rect 10583 2570 10631 2602
rect 10503 2534 10631 2570
rect 10503 2502 10551 2534
rect 10583 2502 10631 2534
rect 10503 2486 10631 2502
rect 10751 3350 10987 3366
rect 10751 3318 10853 3350
rect 10885 3318 10987 3350
rect 10751 3282 10987 3318
rect 10751 3250 10853 3282
rect 10885 3250 10987 3282
rect 10751 3214 10987 3250
rect 10751 3182 10853 3214
rect 10885 3182 10987 3214
rect 10751 3146 10987 3182
rect 10751 3114 10853 3146
rect 10885 3114 10987 3146
rect 10751 3078 10987 3114
rect 10751 3046 10853 3078
rect 10885 3046 10987 3078
rect 10751 3010 10987 3046
rect 10751 2978 10853 3010
rect 10885 2978 10987 3010
rect 10751 2942 10987 2978
rect 10751 2910 10853 2942
rect 10885 2910 10987 2942
rect 10751 2874 10987 2910
rect 10751 2842 10853 2874
rect 10885 2842 10987 2874
rect 10751 2806 10987 2842
rect 10751 2774 10853 2806
rect 10885 2774 10987 2806
rect 10751 2738 10987 2774
rect 10751 2706 10853 2738
rect 10885 2706 10987 2738
rect 10751 2670 10987 2706
rect 10751 2638 10853 2670
rect 10885 2638 10987 2670
rect 10751 2602 10987 2638
rect 10751 2570 10853 2602
rect 10885 2570 10987 2602
rect 10751 2534 10987 2570
rect 10751 2502 10853 2534
rect 10885 2502 10987 2534
rect 10751 2486 10987 2502
rect 11107 3350 11235 3366
rect 11107 3318 11155 3350
rect 11187 3318 11235 3350
rect 11107 3282 11235 3318
rect 11107 3250 11155 3282
rect 11187 3250 11235 3282
rect 11107 3214 11235 3250
rect 11107 3182 11155 3214
rect 11187 3182 11235 3214
rect 11107 3146 11235 3182
rect 11107 3114 11155 3146
rect 11187 3114 11235 3146
rect 11107 3078 11235 3114
rect 11107 3046 11155 3078
rect 11187 3046 11235 3078
rect 11107 3010 11235 3046
rect 11107 2978 11155 3010
rect 11187 2978 11235 3010
rect 11107 2942 11235 2978
rect 11107 2910 11155 2942
rect 11187 2910 11235 2942
rect 11107 2874 11235 2910
rect 11107 2842 11155 2874
rect 11187 2842 11235 2874
rect 11107 2806 11235 2842
rect 11107 2774 11155 2806
rect 11187 2774 11235 2806
rect 11107 2738 11235 2774
rect 11107 2706 11155 2738
rect 11187 2706 11235 2738
rect 11107 2670 11235 2706
rect 11107 2638 11155 2670
rect 11187 2638 11235 2670
rect 11107 2602 11235 2638
rect 11107 2570 11155 2602
rect 11187 2570 11235 2602
rect 11107 2534 11235 2570
rect 11107 2502 11155 2534
rect 11187 2502 11235 2534
rect 11107 2486 11235 2502
rect 11355 3350 11591 3366
rect 11355 3318 11457 3350
rect 11489 3318 11591 3350
rect 11355 3282 11591 3318
rect 11355 3250 11457 3282
rect 11489 3250 11591 3282
rect 11355 3214 11591 3250
rect 11355 3182 11457 3214
rect 11489 3182 11591 3214
rect 11355 3146 11591 3182
rect 11355 3114 11457 3146
rect 11489 3114 11591 3146
rect 11355 3078 11591 3114
rect 11355 3046 11457 3078
rect 11489 3046 11591 3078
rect 11355 3010 11591 3046
rect 11355 2978 11457 3010
rect 11489 2978 11591 3010
rect 11355 2942 11591 2978
rect 11355 2910 11457 2942
rect 11489 2910 11591 2942
rect 11355 2874 11591 2910
rect 11355 2842 11457 2874
rect 11489 2842 11591 2874
rect 11355 2806 11591 2842
rect 11355 2774 11457 2806
rect 11489 2774 11591 2806
rect 11355 2738 11591 2774
rect 11355 2706 11457 2738
rect 11489 2706 11591 2738
rect 11355 2670 11591 2706
rect 11355 2638 11457 2670
rect 11489 2638 11591 2670
rect 11355 2602 11591 2638
rect 11355 2570 11457 2602
rect 11489 2570 11591 2602
rect 11355 2534 11591 2570
rect 11355 2502 11457 2534
rect 11489 2502 11591 2534
rect 11355 2486 11591 2502
rect 11711 3350 11839 3366
rect 11711 3318 11759 3350
rect 11791 3318 11839 3350
rect 11711 3282 11839 3318
rect 11711 3250 11759 3282
rect 11791 3250 11839 3282
rect 11711 3214 11839 3250
rect 11711 3182 11759 3214
rect 11791 3182 11839 3214
rect 11711 3146 11839 3182
rect 11711 3114 11759 3146
rect 11791 3114 11839 3146
rect 11711 3078 11839 3114
rect 11711 3046 11759 3078
rect 11791 3046 11839 3078
rect 11711 3010 11839 3046
rect 11711 2978 11759 3010
rect 11791 2978 11839 3010
rect 11711 2942 11839 2978
rect 11711 2910 11759 2942
rect 11791 2910 11839 2942
rect 11711 2874 11839 2910
rect 11711 2842 11759 2874
rect 11791 2842 11839 2874
rect 11711 2806 11839 2842
rect 11711 2774 11759 2806
rect 11791 2774 11839 2806
rect 11711 2738 11839 2774
rect 11711 2706 11759 2738
rect 11791 2706 11839 2738
rect 11711 2670 11839 2706
rect 11711 2638 11759 2670
rect 11791 2638 11839 2670
rect 11711 2602 11839 2638
rect 11711 2570 11759 2602
rect 11791 2570 11839 2602
rect 11711 2534 11839 2570
rect 11711 2502 11759 2534
rect 11791 2502 11839 2534
rect 11711 2486 11839 2502
rect 11959 3350 12195 3366
rect 11959 3318 12061 3350
rect 12093 3318 12195 3350
rect 11959 3282 12195 3318
rect 11959 3250 12061 3282
rect 12093 3250 12195 3282
rect 11959 3214 12195 3250
rect 11959 3182 12061 3214
rect 12093 3182 12195 3214
rect 11959 3146 12195 3182
rect 11959 3114 12061 3146
rect 12093 3114 12195 3146
rect 11959 3078 12195 3114
rect 11959 3046 12061 3078
rect 12093 3046 12195 3078
rect 11959 3010 12195 3046
rect 11959 2978 12061 3010
rect 12093 2978 12195 3010
rect 11959 2942 12195 2978
rect 11959 2910 12061 2942
rect 12093 2910 12195 2942
rect 11959 2874 12195 2910
rect 11959 2842 12061 2874
rect 12093 2842 12195 2874
rect 11959 2806 12195 2842
rect 11959 2774 12061 2806
rect 12093 2774 12195 2806
rect 11959 2738 12195 2774
rect 11959 2706 12061 2738
rect 12093 2706 12195 2738
rect 11959 2670 12195 2706
rect 11959 2638 12061 2670
rect 12093 2638 12195 2670
rect 11959 2602 12195 2638
rect 11959 2570 12061 2602
rect 12093 2570 12195 2602
rect 11959 2534 12195 2570
rect 11959 2502 12061 2534
rect 12093 2502 12195 2534
rect 11959 2486 12195 2502
rect 12315 3350 12443 3366
rect 12315 3318 12363 3350
rect 12395 3318 12443 3350
rect 12315 3282 12443 3318
rect 12315 3250 12363 3282
rect 12395 3250 12443 3282
rect 12315 3214 12443 3250
rect 12315 3182 12363 3214
rect 12395 3182 12443 3214
rect 12315 3146 12443 3182
rect 12315 3114 12363 3146
rect 12395 3114 12443 3146
rect 12315 3078 12443 3114
rect 12315 3046 12363 3078
rect 12395 3046 12443 3078
rect 12315 3010 12443 3046
rect 12315 2978 12363 3010
rect 12395 2978 12443 3010
rect 12315 2942 12443 2978
rect 12315 2910 12363 2942
rect 12395 2910 12443 2942
rect 12315 2874 12443 2910
rect 12315 2842 12363 2874
rect 12395 2842 12443 2874
rect 12315 2806 12443 2842
rect 12315 2774 12363 2806
rect 12395 2774 12443 2806
rect 12315 2738 12443 2774
rect 12315 2706 12363 2738
rect 12395 2706 12443 2738
rect 12315 2670 12443 2706
rect 12315 2638 12363 2670
rect 12395 2638 12443 2670
rect 12315 2602 12443 2638
rect 12315 2570 12363 2602
rect 12395 2570 12443 2602
rect 12315 2534 12443 2570
rect 12315 2502 12363 2534
rect 12395 2502 12443 2534
rect 12315 2486 12443 2502
rect 12563 3350 12799 3366
rect 12563 3318 12665 3350
rect 12697 3318 12799 3350
rect 12563 3282 12799 3318
rect 12563 3250 12665 3282
rect 12697 3250 12799 3282
rect 12563 3214 12799 3250
rect 12563 3182 12665 3214
rect 12697 3182 12799 3214
rect 12563 3146 12799 3182
rect 12563 3114 12665 3146
rect 12697 3114 12799 3146
rect 12563 3078 12799 3114
rect 12563 3046 12665 3078
rect 12697 3046 12799 3078
rect 12563 3010 12799 3046
rect 12563 2978 12665 3010
rect 12697 2978 12799 3010
rect 12563 2942 12799 2978
rect 12563 2910 12665 2942
rect 12697 2910 12799 2942
rect 12563 2874 12799 2910
rect 12563 2842 12665 2874
rect 12697 2842 12799 2874
rect 12563 2806 12799 2842
rect 12563 2774 12665 2806
rect 12697 2774 12799 2806
rect 12563 2738 12799 2774
rect 12563 2706 12665 2738
rect 12697 2706 12799 2738
rect 12563 2670 12799 2706
rect 12563 2638 12665 2670
rect 12697 2638 12799 2670
rect 12563 2602 12799 2638
rect 12563 2570 12665 2602
rect 12697 2570 12799 2602
rect 12563 2534 12799 2570
rect 12563 2502 12665 2534
rect 12697 2502 12799 2534
rect 12563 2486 12799 2502
rect 12919 3350 13047 3366
rect 12919 3318 12967 3350
rect 12999 3318 13047 3350
rect 12919 3282 13047 3318
rect 12919 3250 12967 3282
rect 12999 3250 13047 3282
rect 12919 3214 13047 3250
rect 12919 3182 12967 3214
rect 12999 3182 13047 3214
rect 12919 3146 13047 3182
rect 12919 3114 12967 3146
rect 12999 3114 13047 3146
rect 12919 3078 13047 3114
rect 12919 3046 12967 3078
rect 12999 3046 13047 3078
rect 12919 3010 13047 3046
rect 12919 2978 12967 3010
rect 12999 2978 13047 3010
rect 12919 2942 13047 2978
rect 12919 2910 12967 2942
rect 12999 2910 13047 2942
rect 12919 2874 13047 2910
rect 12919 2842 12967 2874
rect 12999 2842 13047 2874
rect 12919 2806 13047 2842
rect 12919 2774 12967 2806
rect 12999 2774 13047 2806
rect 12919 2738 13047 2774
rect 12919 2706 12967 2738
rect 12999 2706 13047 2738
rect 12919 2670 13047 2706
rect 12919 2638 12967 2670
rect 12999 2638 13047 2670
rect 12919 2602 13047 2638
rect 12919 2570 12967 2602
rect 12999 2570 13047 2602
rect 12919 2534 13047 2570
rect 12919 2502 12967 2534
rect 12999 2502 13047 2534
rect 12919 2486 13047 2502
rect 13167 3350 13403 3366
rect 13167 3318 13269 3350
rect 13301 3318 13403 3350
rect 13167 3282 13403 3318
rect 13167 3250 13269 3282
rect 13301 3250 13403 3282
rect 13167 3214 13403 3250
rect 13167 3182 13269 3214
rect 13301 3182 13403 3214
rect 13167 3146 13403 3182
rect 13167 3114 13269 3146
rect 13301 3114 13403 3146
rect 13167 3078 13403 3114
rect 13167 3046 13269 3078
rect 13301 3046 13403 3078
rect 13167 3010 13403 3046
rect 13167 2978 13269 3010
rect 13301 2978 13403 3010
rect 13167 2942 13403 2978
rect 13167 2910 13269 2942
rect 13301 2910 13403 2942
rect 13167 2874 13403 2910
rect 13167 2842 13269 2874
rect 13301 2842 13403 2874
rect 13167 2806 13403 2842
rect 13167 2774 13269 2806
rect 13301 2774 13403 2806
rect 13167 2738 13403 2774
rect 13167 2706 13269 2738
rect 13301 2706 13403 2738
rect 13167 2670 13403 2706
rect 13167 2638 13269 2670
rect 13301 2638 13403 2670
rect 13167 2602 13403 2638
rect 13167 2570 13269 2602
rect 13301 2570 13403 2602
rect 13167 2534 13403 2570
rect 13167 2502 13269 2534
rect 13301 2502 13403 2534
rect 13167 2486 13403 2502
rect 13523 3350 13651 3366
rect 13523 3318 13571 3350
rect 13603 3318 13651 3350
rect 13523 3282 13651 3318
rect 13523 3250 13571 3282
rect 13603 3250 13651 3282
rect 13523 3214 13651 3250
rect 13523 3182 13571 3214
rect 13603 3182 13651 3214
rect 13523 3146 13651 3182
rect 13523 3114 13571 3146
rect 13603 3114 13651 3146
rect 13523 3078 13651 3114
rect 13523 3046 13571 3078
rect 13603 3046 13651 3078
rect 13523 3010 13651 3046
rect 13523 2978 13571 3010
rect 13603 2978 13651 3010
rect 13523 2942 13651 2978
rect 13523 2910 13571 2942
rect 13603 2910 13651 2942
rect 13523 2874 13651 2910
rect 13523 2842 13571 2874
rect 13603 2842 13651 2874
rect 13523 2806 13651 2842
rect 13523 2774 13571 2806
rect 13603 2774 13651 2806
rect 13523 2738 13651 2774
rect 13523 2706 13571 2738
rect 13603 2706 13651 2738
rect 13523 2670 13651 2706
rect 13523 2638 13571 2670
rect 13603 2638 13651 2670
rect 13523 2602 13651 2638
rect 13523 2570 13571 2602
rect 13603 2570 13651 2602
rect 13523 2534 13651 2570
rect 13523 2502 13571 2534
rect 13603 2502 13651 2534
rect 13523 2486 13651 2502
rect 13771 3350 14007 3366
rect 13771 3318 13873 3350
rect 13905 3318 14007 3350
rect 13771 3282 14007 3318
rect 13771 3250 13873 3282
rect 13905 3250 14007 3282
rect 13771 3214 14007 3250
rect 13771 3182 13873 3214
rect 13905 3182 14007 3214
rect 13771 3146 14007 3182
rect 13771 3114 13873 3146
rect 13905 3114 14007 3146
rect 13771 3078 14007 3114
rect 13771 3046 13873 3078
rect 13905 3046 14007 3078
rect 13771 3010 14007 3046
rect 13771 2978 13873 3010
rect 13905 2978 14007 3010
rect 13771 2942 14007 2978
rect 13771 2910 13873 2942
rect 13905 2910 14007 2942
rect 13771 2874 14007 2910
rect 13771 2842 13873 2874
rect 13905 2842 14007 2874
rect 13771 2806 14007 2842
rect 13771 2774 13873 2806
rect 13905 2774 14007 2806
rect 13771 2738 14007 2774
rect 13771 2706 13873 2738
rect 13905 2706 14007 2738
rect 13771 2670 14007 2706
rect 13771 2638 13873 2670
rect 13905 2638 14007 2670
rect 13771 2602 14007 2638
rect 13771 2570 13873 2602
rect 13905 2570 14007 2602
rect 13771 2534 14007 2570
rect 13771 2502 13873 2534
rect 13905 2502 14007 2534
rect 13771 2486 14007 2502
rect 14127 3350 14255 3366
rect 14127 3318 14175 3350
rect 14207 3318 14255 3350
rect 14127 3282 14255 3318
rect 14127 3250 14175 3282
rect 14207 3250 14255 3282
rect 14127 3214 14255 3250
rect 14127 3182 14175 3214
rect 14207 3182 14255 3214
rect 14127 3146 14255 3182
rect 14127 3114 14175 3146
rect 14207 3114 14255 3146
rect 14127 3078 14255 3114
rect 14127 3046 14175 3078
rect 14207 3046 14255 3078
rect 14127 3010 14255 3046
rect 14127 2978 14175 3010
rect 14207 2978 14255 3010
rect 14127 2942 14255 2978
rect 14127 2910 14175 2942
rect 14207 2910 14255 2942
rect 14127 2874 14255 2910
rect 14127 2842 14175 2874
rect 14207 2842 14255 2874
rect 14127 2806 14255 2842
rect 14127 2774 14175 2806
rect 14207 2774 14255 2806
rect 14127 2738 14255 2774
rect 14127 2706 14175 2738
rect 14207 2706 14255 2738
rect 14127 2670 14255 2706
rect 14127 2638 14175 2670
rect 14207 2638 14255 2670
rect 14127 2602 14255 2638
rect 14127 2570 14175 2602
rect 14207 2570 14255 2602
rect 14127 2534 14255 2570
rect 14127 2502 14175 2534
rect 14207 2502 14255 2534
rect 14127 2486 14255 2502
rect 14375 3350 14523 3366
rect 14375 3318 14477 3350
rect 14509 3318 14523 3350
rect 14375 3282 14523 3318
rect 14375 3250 14477 3282
rect 14509 3250 14523 3282
rect 14375 3214 14523 3250
rect 14375 3182 14477 3214
rect 14509 3182 14523 3214
rect 14375 3146 14523 3182
rect 14375 3114 14477 3146
rect 14509 3114 14523 3146
rect 14375 3078 14523 3114
rect 14375 3046 14477 3078
rect 14509 3046 14523 3078
rect 14375 3010 14523 3046
rect 14375 2978 14477 3010
rect 14509 2978 14523 3010
rect 14375 2942 14523 2978
rect 14375 2910 14477 2942
rect 14509 2910 14523 2942
rect 14375 2874 14523 2910
rect 14375 2842 14477 2874
rect 14509 2842 14523 2874
rect 14375 2806 14523 2842
rect 14375 2774 14477 2806
rect 14509 2774 14523 2806
rect 14375 2738 14523 2774
rect 14375 2706 14477 2738
rect 14509 2706 14523 2738
rect 14375 2670 14523 2706
rect 14375 2638 14477 2670
rect 14509 2638 14523 2670
rect 14375 2602 14523 2638
rect 14375 2570 14477 2602
rect 14509 2570 14523 2602
rect 14375 2534 14523 2570
rect 14375 2502 14477 2534
rect 14509 2502 14523 2534
rect 14375 2486 14523 2502
rect 1477 2382 1571 2398
rect 1477 2350 1491 2382
rect 1523 2350 1571 2382
rect 1477 2314 1571 2350
rect 1477 2282 1491 2314
rect 1523 2282 1571 2314
rect 1477 2246 1571 2282
rect 1477 2214 1491 2246
rect 1523 2214 1571 2246
rect 1477 2178 1571 2214
rect 1477 2146 1491 2178
rect 1523 2146 1571 2178
rect 1477 2110 1571 2146
rect 1477 2078 1491 2110
rect 1523 2078 1571 2110
rect 1477 2042 1571 2078
rect 1477 2010 1491 2042
rect 1523 2010 1571 2042
rect 1477 1974 1571 2010
rect 1477 1942 1491 1974
rect 1523 1942 1571 1974
rect 1477 1906 1571 1942
rect 1477 1874 1491 1906
rect 1523 1874 1571 1906
rect 1477 1838 1571 1874
rect 1477 1806 1491 1838
rect 1523 1806 1571 1838
rect 1477 1770 1571 1806
rect 1477 1738 1491 1770
rect 1523 1738 1571 1770
rect 1477 1702 1571 1738
rect 1477 1670 1491 1702
rect 1523 1670 1571 1702
rect 1477 1634 1571 1670
rect 1477 1602 1491 1634
rect 1523 1602 1571 1634
rect 1477 1566 1571 1602
rect 1477 1534 1491 1566
rect 1523 1534 1571 1566
rect 1477 1518 1571 1534
rect 1691 2382 1927 2398
rect 1691 2350 1793 2382
rect 1825 2350 1927 2382
rect 1691 2314 1927 2350
rect 1691 2282 1793 2314
rect 1825 2282 1927 2314
rect 1691 2246 1927 2282
rect 1691 2214 1793 2246
rect 1825 2214 1927 2246
rect 1691 2178 1927 2214
rect 1691 2146 1793 2178
rect 1825 2146 1927 2178
rect 1691 2110 1927 2146
rect 1691 2078 1793 2110
rect 1825 2078 1927 2110
rect 1691 2042 1927 2078
rect 1691 2010 1793 2042
rect 1825 2010 1927 2042
rect 1691 1974 1927 2010
rect 1691 1942 1793 1974
rect 1825 1942 1927 1974
rect 1691 1906 1927 1942
rect 1691 1874 1793 1906
rect 1825 1874 1927 1906
rect 1691 1838 1927 1874
rect 1691 1806 1793 1838
rect 1825 1806 1927 1838
rect 1691 1770 1927 1806
rect 1691 1738 1793 1770
rect 1825 1738 1927 1770
rect 1691 1702 1927 1738
rect 1691 1670 1793 1702
rect 1825 1670 1927 1702
rect 1691 1634 1927 1670
rect 1691 1602 1793 1634
rect 1825 1602 1927 1634
rect 1691 1566 1927 1602
rect 1691 1534 1793 1566
rect 1825 1534 1927 1566
rect 1691 1518 1927 1534
rect 2047 2382 2175 2398
rect 2047 2350 2095 2382
rect 2127 2350 2175 2382
rect 2047 2314 2175 2350
rect 2047 2282 2095 2314
rect 2127 2282 2175 2314
rect 2047 2246 2175 2282
rect 2047 2214 2095 2246
rect 2127 2214 2175 2246
rect 2047 2178 2175 2214
rect 2047 2146 2095 2178
rect 2127 2146 2175 2178
rect 2047 2110 2175 2146
rect 2047 2078 2095 2110
rect 2127 2078 2175 2110
rect 2047 2042 2175 2078
rect 2047 2010 2095 2042
rect 2127 2010 2175 2042
rect 2047 1974 2175 2010
rect 2047 1942 2095 1974
rect 2127 1942 2175 1974
rect 2047 1906 2175 1942
rect 2047 1874 2095 1906
rect 2127 1874 2175 1906
rect 2047 1838 2175 1874
rect 2047 1806 2095 1838
rect 2127 1806 2175 1838
rect 2047 1770 2175 1806
rect 2047 1738 2095 1770
rect 2127 1738 2175 1770
rect 2047 1702 2175 1738
rect 2047 1670 2095 1702
rect 2127 1670 2175 1702
rect 2047 1634 2175 1670
rect 2047 1602 2095 1634
rect 2127 1602 2175 1634
rect 2047 1566 2175 1602
rect 2047 1534 2095 1566
rect 2127 1534 2175 1566
rect 2047 1518 2175 1534
rect 2295 2382 2531 2398
rect 2295 2350 2397 2382
rect 2429 2350 2531 2382
rect 2295 2314 2531 2350
rect 2295 2282 2397 2314
rect 2429 2282 2531 2314
rect 2295 2246 2531 2282
rect 2295 2214 2397 2246
rect 2429 2214 2531 2246
rect 2295 2178 2531 2214
rect 2295 2146 2397 2178
rect 2429 2146 2531 2178
rect 2295 2110 2531 2146
rect 2295 2078 2397 2110
rect 2429 2078 2531 2110
rect 2295 2042 2531 2078
rect 2295 2010 2397 2042
rect 2429 2010 2531 2042
rect 2295 1974 2531 2010
rect 2295 1942 2397 1974
rect 2429 1942 2531 1974
rect 2295 1906 2531 1942
rect 2295 1874 2397 1906
rect 2429 1874 2531 1906
rect 2295 1838 2531 1874
rect 2295 1806 2397 1838
rect 2429 1806 2531 1838
rect 2295 1770 2531 1806
rect 2295 1738 2397 1770
rect 2429 1738 2531 1770
rect 2295 1702 2531 1738
rect 2295 1670 2397 1702
rect 2429 1670 2531 1702
rect 2295 1634 2531 1670
rect 2295 1602 2397 1634
rect 2429 1602 2531 1634
rect 2295 1566 2531 1602
rect 2295 1534 2397 1566
rect 2429 1534 2531 1566
rect 2295 1518 2531 1534
rect 2651 2382 2779 2398
rect 2651 2350 2699 2382
rect 2731 2350 2779 2382
rect 2651 2314 2779 2350
rect 2651 2282 2699 2314
rect 2731 2282 2779 2314
rect 2651 2246 2779 2282
rect 2651 2214 2699 2246
rect 2731 2214 2779 2246
rect 2651 2178 2779 2214
rect 2651 2146 2699 2178
rect 2731 2146 2779 2178
rect 2651 2110 2779 2146
rect 2651 2078 2699 2110
rect 2731 2078 2779 2110
rect 2651 2042 2779 2078
rect 2651 2010 2699 2042
rect 2731 2010 2779 2042
rect 2651 1974 2779 2010
rect 2651 1942 2699 1974
rect 2731 1942 2779 1974
rect 2651 1906 2779 1942
rect 2651 1874 2699 1906
rect 2731 1874 2779 1906
rect 2651 1838 2779 1874
rect 2651 1806 2699 1838
rect 2731 1806 2779 1838
rect 2651 1770 2779 1806
rect 2651 1738 2699 1770
rect 2731 1738 2779 1770
rect 2651 1702 2779 1738
rect 2651 1670 2699 1702
rect 2731 1670 2779 1702
rect 2651 1634 2779 1670
rect 2651 1602 2699 1634
rect 2731 1602 2779 1634
rect 2651 1566 2779 1602
rect 2651 1534 2699 1566
rect 2731 1534 2779 1566
rect 2651 1518 2779 1534
rect 2899 2382 3135 2398
rect 2899 2350 3001 2382
rect 3033 2350 3135 2382
rect 2899 2314 3135 2350
rect 2899 2282 3001 2314
rect 3033 2282 3135 2314
rect 2899 2246 3135 2282
rect 2899 2214 3001 2246
rect 3033 2214 3135 2246
rect 2899 2178 3135 2214
rect 2899 2146 3001 2178
rect 3033 2146 3135 2178
rect 2899 2110 3135 2146
rect 2899 2078 3001 2110
rect 3033 2078 3135 2110
rect 2899 2042 3135 2078
rect 2899 2010 3001 2042
rect 3033 2010 3135 2042
rect 2899 1974 3135 2010
rect 2899 1942 3001 1974
rect 3033 1942 3135 1974
rect 2899 1906 3135 1942
rect 2899 1874 3001 1906
rect 3033 1874 3135 1906
rect 2899 1838 3135 1874
rect 2899 1806 3001 1838
rect 3033 1806 3135 1838
rect 2899 1770 3135 1806
rect 2899 1738 3001 1770
rect 3033 1738 3135 1770
rect 2899 1702 3135 1738
rect 2899 1670 3001 1702
rect 3033 1670 3135 1702
rect 2899 1634 3135 1670
rect 2899 1602 3001 1634
rect 3033 1602 3135 1634
rect 2899 1566 3135 1602
rect 2899 1534 3001 1566
rect 3033 1534 3135 1566
rect 2899 1518 3135 1534
rect 3255 2382 3383 2398
rect 3255 2350 3303 2382
rect 3335 2350 3383 2382
rect 3255 2314 3383 2350
rect 3255 2282 3303 2314
rect 3335 2282 3383 2314
rect 3255 2246 3383 2282
rect 3255 2214 3303 2246
rect 3335 2214 3383 2246
rect 3255 2178 3383 2214
rect 3255 2146 3303 2178
rect 3335 2146 3383 2178
rect 3255 2110 3383 2146
rect 3255 2078 3303 2110
rect 3335 2078 3383 2110
rect 3255 2042 3383 2078
rect 3255 2010 3303 2042
rect 3335 2010 3383 2042
rect 3255 1974 3383 2010
rect 3255 1942 3303 1974
rect 3335 1942 3383 1974
rect 3255 1906 3383 1942
rect 3255 1874 3303 1906
rect 3335 1874 3383 1906
rect 3255 1838 3383 1874
rect 3255 1806 3303 1838
rect 3335 1806 3383 1838
rect 3255 1770 3383 1806
rect 3255 1738 3303 1770
rect 3335 1738 3383 1770
rect 3255 1702 3383 1738
rect 3255 1670 3303 1702
rect 3335 1670 3383 1702
rect 3255 1634 3383 1670
rect 3255 1602 3303 1634
rect 3335 1602 3383 1634
rect 3255 1566 3383 1602
rect 3255 1534 3303 1566
rect 3335 1534 3383 1566
rect 3255 1518 3383 1534
rect 3503 2382 3739 2398
rect 3503 2350 3605 2382
rect 3637 2350 3739 2382
rect 3503 2314 3739 2350
rect 3503 2282 3605 2314
rect 3637 2282 3739 2314
rect 3503 2246 3739 2282
rect 3503 2214 3605 2246
rect 3637 2214 3739 2246
rect 3503 2178 3739 2214
rect 3503 2146 3605 2178
rect 3637 2146 3739 2178
rect 3503 2110 3739 2146
rect 3503 2078 3605 2110
rect 3637 2078 3739 2110
rect 3503 2042 3739 2078
rect 3503 2010 3605 2042
rect 3637 2010 3739 2042
rect 3503 1974 3739 2010
rect 3503 1942 3605 1974
rect 3637 1942 3739 1974
rect 3503 1906 3739 1942
rect 3503 1874 3605 1906
rect 3637 1874 3739 1906
rect 3503 1838 3739 1874
rect 3503 1806 3605 1838
rect 3637 1806 3739 1838
rect 3503 1770 3739 1806
rect 3503 1738 3605 1770
rect 3637 1738 3739 1770
rect 3503 1702 3739 1738
rect 3503 1670 3605 1702
rect 3637 1670 3739 1702
rect 3503 1634 3739 1670
rect 3503 1602 3605 1634
rect 3637 1602 3739 1634
rect 3503 1566 3739 1602
rect 3503 1534 3605 1566
rect 3637 1534 3739 1566
rect 3503 1518 3739 1534
rect 3859 2382 3987 2398
rect 3859 2350 3907 2382
rect 3939 2350 3987 2382
rect 3859 2314 3987 2350
rect 3859 2282 3907 2314
rect 3939 2282 3987 2314
rect 3859 2246 3987 2282
rect 3859 2214 3907 2246
rect 3939 2214 3987 2246
rect 3859 2178 3987 2214
rect 3859 2146 3907 2178
rect 3939 2146 3987 2178
rect 3859 2110 3987 2146
rect 3859 2078 3907 2110
rect 3939 2078 3987 2110
rect 3859 2042 3987 2078
rect 3859 2010 3907 2042
rect 3939 2010 3987 2042
rect 3859 1974 3987 2010
rect 3859 1942 3907 1974
rect 3939 1942 3987 1974
rect 3859 1906 3987 1942
rect 3859 1874 3907 1906
rect 3939 1874 3987 1906
rect 3859 1838 3987 1874
rect 3859 1806 3907 1838
rect 3939 1806 3987 1838
rect 3859 1770 3987 1806
rect 3859 1738 3907 1770
rect 3939 1738 3987 1770
rect 3859 1702 3987 1738
rect 3859 1670 3907 1702
rect 3939 1670 3987 1702
rect 3859 1634 3987 1670
rect 3859 1602 3907 1634
rect 3939 1602 3987 1634
rect 3859 1566 3987 1602
rect 3859 1534 3907 1566
rect 3939 1534 3987 1566
rect 3859 1518 3987 1534
rect 4107 2382 4343 2398
rect 4107 2350 4209 2382
rect 4241 2350 4343 2382
rect 4107 2314 4343 2350
rect 4107 2282 4209 2314
rect 4241 2282 4343 2314
rect 4107 2246 4343 2282
rect 4107 2214 4209 2246
rect 4241 2214 4343 2246
rect 4107 2178 4343 2214
rect 4107 2146 4209 2178
rect 4241 2146 4343 2178
rect 4107 2110 4343 2146
rect 4107 2078 4209 2110
rect 4241 2078 4343 2110
rect 4107 2042 4343 2078
rect 4107 2010 4209 2042
rect 4241 2010 4343 2042
rect 4107 1974 4343 2010
rect 4107 1942 4209 1974
rect 4241 1942 4343 1974
rect 4107 1906 4343 1942
rect 4107 1874 4209 1906
rect 4241 1874 4343 1906
rect 4107 1838 4343 1874
rect 4107 1806 4209 1838
rect 4241 1806 4343 1838
rect 4107 1770 4343 1806
rect 4107 1738 4209 1770
rect 4241 1738 4343 1770
rect 4107 1702 4343 1738
rect 4107 1670 4209 1702
rect 4241 1670 4343 1702
rect 4107 1634 4343 1670
rect 4107 1602 4209 1634
rect 4241 1602 4343 1634
rect 4107 1566 4343 1602
rect 4107 1534 4209 1566
rect 4241 1534 4343 1566
rect 4107 1518 4343 1534
rect 4463 2382 4591 2398
rect 4463 2350 4511 2382
rect 4543 2350 4591 2382
rect 4463 2314 4591 2350
rect 4463 2282 4511 2314
rect 4543 2282 4591 2314
rect 4463 2246 4591 2282
rect 4463 2214 4511 2246
rect 4543 2214 4591 2246
rect 4463 2178 4591 2214
rect 4463 2146 4511 2178
rect 4543 2146 4591 2178
rect 4463 2110 4591 2146
rect 4463 2078 4511 2110
rect 4543 2078 4591 2110
rect 4463 2042 4591 2078
rect 4463 2010 4511 2042
rect 4543 2010 4591 2042
rect 4463 1974 4591 2010
rect 4463 1942 4511 1974
rect 4543 1942 4591 1974
rect 4463 1906 4591 1942
rect 4463 1874 4511 1906
rect 4543 1874 4591 1906
rect 4463 1838 4591 1874
rect 4463 1806 4511 1838
rect 4543 1806 4591 1838
rect 4463 1770 4591 1806
rect 4463 1738 4511 1770
rect 4543 1738 4591 1770
rect 4463 1702 4591 1738
rect 4463 1670 4511 1702
rect 4543 1670 4591 1702
rect 4463 1634 4591 1670
rect 4463 1602 4511 1634
rect 4543 1602 4591 1634
rect 4463 1566 4591 1602
rect 4463 1534 4511 1566
rect 4543 1534 4591 1566
rect 4463 1518 4591 1534
rect 4711 2382 4947 2398
rect 4711 2350 4813 2382
rect 4845 2350 4947 2382
rect 4711 2314 4947 2350
rect 4711 2282 4813 2314
rect 4845 2282 4947 2314
rect 4711 2246 4947 2282
rect 4711 2214 4813 2246
rect 4845 2214 4947 2246
rect 4711 2178 4947 2214
rect 4711 2146 4813 2178
rect 4845 2146 4947 2178
rect 4711 2110 4947 2146
rect 4711 2078 4813 2110
rect 4845 2078 4947 2110
rect 4711 2042 4947 2078
rect 4711 2010 4813 2042
rect 4845 2010 4947 2042
rect 4711 1974 4947 2010
rect 4711 1942 4813 1974
rect 4845 1942 4947 1974
rect 4711 1906 4947 1942
rect 4711 1874 4813 1906
rect 4845 1874 4947 1906
rect 4711 1838 4947 1874
rect 4711 1806 4813 1838
rect 4845 1806 4947 1838
rect 4711 1770 4947 1806
rect 4711 1738 4813 1770
rect 4845 1738 4947 1770
rect 4711 1702 4947 1738
rect 4711 1670 4813 1702
rect 4845 1670 4947 1702
rect 4711 1634 4947 1670
rect 4711 1602 4813 1634
rect 4845 1602 4947 1634
rect 4711 1566 4947 1602
rect 4711 1534 4813 1566
rect 4845 1534 4947 1566
rect 4711 1518 4947 1534
rect 5067 2382 5195 2398
rect 5067 2350 5115 2382
rect 5147 2350 5195 2382
rect 5067 2314 5195 2350
rect 5067 2282 5115 2314
rect 5147 2282 5195 2314
rect 5067 2246 5195 2282
rect 5067 2214 5115 2246
rect 5147 2214 5195 2246
rect 5067 2178 5195 2214
rect 5067 2146 5115 2178
rect 5147 2146 5195 2178
rect 5067 2110 5195 2146
rect 5067 2078 5115 2110
rect 5147 2078 5195 2110
rect 5067 2042 5195 2078
rect 5067 2010 5115 2042
rect 5147 2010 5195 2042
rect 5067 1974 5195 2010
rect 5067 1942 5115 1974
rect 5147 1942 5195 1974
rect 5067 1906 5195 1942
rect 5067 1874 5115 1906
rect 5147 1874 5195 1906
rect 5067 1838 5195 1874
rect 5067 1806 5115 1838
rect 5147 1806 5195 1838
rect 5067 1770 5195 1806
rect 5067 1738 5115 1770
rect 5147 1738 5195 1770
rect 5067 1702 5195 1738
rect 5067 1670 5115 1702
rect 5147 1670 5195 1702
rect 5067 1634 5195 1670
rect 5067 1602 5115 1634
rect 5147 1602 5195 1634
rect 5067 1566 5195 1602
rect 5067 1534 5115 1566
rect 5147 1534 5195 1566
rect 5067 1518 5195 1534
rect 5315 2382 5551 2398
rect 5315 2350 5417 2382
rect 5449 2350 5551 2382
rect 5315 2314 5551 2350
rect 5315 2282 5417 2314
rect 5449 2282 5551 2314
rect 5315 2246 5551 2282
rect 5315 2214 5417 2246
rect 5449 2214 5551 2246
rect 5315 2178 5551 2214
rect 5315 2146 5417 2178
rect 5449 2146 5551 2178
rect 5315 2110 5551 2146
rect 5315 2078 5417 2110
rect 5449 2078 5551 2110
rect 5315 2042 5551 2078
rect 5315 2010 5417 2042
rect 5449 2010 5551 2042
rect 5315 1974 5551 2010
rect 5315 1942 5417 1974
rect 5449 1942 5551 1974
rect 5315 1906 5551 1942
rect 5315 1874 5417 1906
rect 5449 1874 5551 1906
rect 5315 1838 5551 1874
rect 5315 1806 5417 1838
rect 5449 1806 5551 1838
rect 5315 1770 5551 1806
rect 5315 1738 5417 1770
rect 5449 1738 5551 1770
rect 5315 1702 5551 1738
rect 5315 1670 5417 1702
rect 5449 1670 5551 1702
rect 5315 1634 5551 1670
rect 5315 1602 5417 1634
rect 5449 1602 5551 1634
rect 5315 1566 5551 1602
rect 5315 1534 5417 1566
rect 5449 1534 5551 1566
rect 5315 1518 5551 1534
rect 5671 2382 5799 2398
rect 5671 2350 5719 2382
rect 5751 2350 5799 2382
rect 5671 2314 5799 2350
rect 5671 2282 5719 2314
rect 5751 2282 5799 2314
rect 5671 2246 5799 2282
rect 5671 2214 5719 2246
rect 5751 2214 5799 2246
rect 5671 2178 5799 2214
rect 5671 2146 5719 2178
rect 5751 2146 5799 2178
rect 5671 2110 5799 2146
rect 5671 2078 5719 2110
rect 5751 2078 5799 2110
rect 5671 2042 5799 2078
rect 5671 2010 5719 2042
rect 5751 2010 5799 2042
rect 5671 1974 5799 2010
rect 5671 1942 5719 1974
rect 5751 1942 5799 1974
rect 5671 1906 5799 1942
rect 5671 1874 5719 1906
rect 5751 1874 5799 1906
rect 5671 1838 5799 1874
rect 5671 1806 5719 1838
rect 5751 1806 5799 1838
rect 5671 1770 5799 1806
rect 5671 1738 5719 1770
rect 5751 1738 5799 1770
rect 5671 1702 5799 1738
rect 5671 1670 5719 1702
rect 5751 1670 5799 1702
rect 5671 1634 5799 1670
rect 5671 1602 5719 1634
rect 5751 1602 5799 1634
rect 5671 1566 5799 1602
rect 5671 1534 5719 1566
rect 5751 1534 5799 1566
rect 5671 1518 5799 1534
rect 5919 2382 6155 2398
rect 5919 2350 6021 2382
rect 6053 2350 6155 2382
rect 5919 2314 6155 2350
rect 5919 2282 6021 2314
rect 6053 2282 6155 2314
rect 5919 2246 6155 2282
rect 5919 2214 6021 2246
rect 6053 2214 6155 2246
rect 5919 2178 6155 2214
rect 5919 2146 6021 2178
rect 6053 2146 6155 2178
rect 5919 2110 6155 2146
rect 5919 2078 6021 2110
rect 6053 2078 6155 2110
rect 5919 2042 6155 2078
rect 5919 2010 6021 2042
rect 6053 2010 6155 2042
rect 5919 1974 6155 2010
rect 5919 1942 6021 1974
rect 6053 1942 6155 1974
rect 5919 1906 6155 1942
rect 5919 1874 6021 1906
rect 6053 1874 6155 1906
rect 5919 1838 6155 1874
rect 5919 1806 6021 1838
rect 6053 1806 6155 1838
rect 5919 1770 6155 1806
rect 5919 1738 6021 1770
rect 6053 1738 6155 1770
rect 5919 1702 6155 1738
rect 5919 1670 6021 1702
rect 6053 1670 6155 1702
rect 5919 1634 6155 1670
rect 5919 1602 6021 1634
rect 6053 1602 6155 1634
rect 5919 1566 6155 1602
rect 5919 1534 6021 1566
rect 6053 1534 6155 1566
rect 5919 1518 6155 1534
rect 6275 2382 6403 2398
rect 6275 2350 6323 2382
rect 6355 2350 6403 2382
rect 6275 2314 6403 2350
rect 6275 2282 6323 2314
rect 6355 2282 6403 2314
rect 6275 2246 6403 2282
rect 6275 2214 6323 2246
rect 6355 2214 6403 2246
rect 6275 2178 6403 2214
rect 6275 2146 6323 2178
rect 6355 2146 6403 2178
rect 6275 2110 6403 2146
rect 6275 2078 6323 2110
rect 6355 2078 6403 2110
rect 6275 2042 6403 2078
rect 6275 2010 6323 2042
rect 6355 2010 6403 2042
rect 6275 1974 6403 2010
rect 6275 1942 6323 1974
rect 6355 1942 6403 1974
rect 6275 1906 6403 1942
rect 6275 1874 6323 1906
rect 6355 1874 6403 1906
rect 6275 1838 6403 1874
rect 6275 1806 6323 1838
rect 6355 1806 6403 1838
rect 6275 1770 6403 1806
rect 6275 1738 6323 1770
rect 6355 1738 6403 1770
rect 6275 1702 6403 1738
rect 6275 1670 6323 1702
rect 6355 1670 6403 1702
rect 6275 1634 6403 1670
rect 6275 1602 6323 1634
rect 6355 1602 6403 1634
rect 6275 1566 6403 1602
rect 6275 1534 6323 1566
rect 6355 1534 6403 1566
rect 6275 1518 6403 1534
rect 6523 2382 6759 2398
rect 6523 2350 6625 2382
rect 6657 2350 6759 2382
rect 6523 2314 6759 2350
rect 6523 2282 6625 2314
rect 6657 2282 6759 2314
rect 6523 2246 6759 2282
rect 6523 2214 6625 2246
rect 6657 2214 6759 2246
rect 6523 2178 6759 2214
rect 6523 2146 6625 2178
rect 6657 2146 6759 2178
rect 6523 2110 6759 2146
rect 6523 2078 6625 2110
rect 6657 2078 6759 2110
rect 6523 2042 6759 2078
rect 6523 2010 6625 2042
rect 6657 2010 6759 2042
rect 6523 1974 6759 2010
rect 6523 1942 6625 1974
rect 6657 1942 6759 1974
rect 6523 1906 6759 1942
rect 6523 1874 6625 1906
rect 6657 1874 6759 1906
rect 6523 1838 6759 1874
rect 6523 1806 6625 1838
rect 6657 1806 6759 1838
rect 6523 1770 6759 1806
rect 6523 1738 6625 1770
rect 6657 1738 6759 1770
rect 6523 1702 6759 1738
rect 6523 1670 6625 1702
rect 6657 1670 6759 1702
rect 6523 1634 6759 1670
rect 6523 1602 6625 1634
rect 6657 1602 6759 1634
rect 6523 1566 6759 1602
rect 6523 1534 6625 1566
rect 6657 1534 6759 1566
rect 6523 1518 6759 1534
rect 6879 2382 7007 2398
rect 6879 2350 6927 2382
rect 6959 2350 7007 2382
rect 6879 2314 7007 2350
rect 6879 2282 6927 2314
rect 6959 2282 7007 2314
rect 6879 2246 7007 2282
rect 6879 2214 6927 2246
rect 6959 2214 7007 2246
rect 6879 2178 7007 2214
rect 6879 2146 6927 2178
rect 6959 2146 7007 2178
rect 6879 2110 7007 2146
rect 6879 2078 6927 2110
rect 6959 2078 7007 2110
rect 6879 2042 7007 2078
rect 6879 2010 6927 2042
rect 6959 2010 7007 2042
rect 6879 1974 7007 2010
rect 6879 1942 6927 1974
rect 6959 1942 7007 1974
rect 6879 1906 7007 1942
rect 6879 1874 6927 1906
rect 6959 1874 7007 1906
rect 6879 1838 7007 1874
rect 6879 1806 6927 1838
rect 6959 1806 7007 1838
rect 6879 1770 7007 1806
rect 6879 1738 6927 1770
rect 6959 1738 7007 1770
rect 6879 1702 7007 1738
rect 6879 1670 6927 1702
rect 6959 1670 7007 1702
rect 6879 1634 7007 1670
rect 6879 1602 6927 1634
rect 6959 1602 7007 1634
rect 6879 1566 7007 1602
rect 6879 1534 6927 1566
rect 6959 1534 7007 1566
rect 6879 1518 7007 1534
rect 7127 2382 7363 2398
rect 7127 2350 7229 2382
rect 7261 2350 7363 2382
rect 7127 2314 7363 2350
rect 7127 2282 7229 2314
rect 7261 2282 7363 2314
rect 7127 2246 7363 2282
rect 7127 2214 7229 2246
rect 7261 2214 7363 2246
rect 7127 2178 7363 2214
rect 7127 2146 7229 2178
rect 7261 2146 7363 2178
rect 7127 2110 7363 2146
rect 7127 2078 7229 2110
rect 7261 2078 7363 2110
rect 7127 2042 7363 2078
rect 7127 2010 7229 2042
rect 7261 2010 7363 2042
rect 7127 1974 7363 2010
rect 7127 1942 7229 1974
rect 7261 1942 7363 1974
rect 7127 1906 7363 1942
rect 7127 1874 7229 1906
rect 7261 1874 7363 1906
rect 7127 1838 7363 1874
rect 7127 1806 7229 1838
rect 7261 1806 7363 1838
rect 7127 1770 7363 1806
rect 7127 1738 7229 1770
rect 7261 1738 7363 1770
rect 7127 1702 7363 1738
rect 7127 1670 7229 1702
rect 7261 1670 7363 1702
rect 7127 1634 7363 1670
rect 7127 1602 7229 1634
rect 7261 1602 7363 1634
rect 7127 1566 7363 1602
rect 7127 1534 7229 1566
rect 7261 1534 7363 1566
rect 7127 1518 7363 1534
rect 7483 2382 7611 2398
rect 7483 2350 7531 2382
rect 7563 2350 7611 2382
rect 7483 2314 7611 2350
rect 7483 2282 7531 2314
rect 7563 2282 7611 2314
rect 7483 2246 7611 2282
rect 7483 2214 7531 2246
rect 7563 2214 7611 2246
rect 7483 2178 7611 2214
rect 7483 2146 7531 2178
rect 7563 2146 7611 2178
rect 7483 2110 7611 2146
rect 7483 2078 7531 2110
rect 7563 2078 7611 2110
rect 7483 2042 7611 2078
rect 7483 2010 7531 2042
rect 7563 2010 7611 2042
rect 7483 1974 7611 2010
rect 7483 1942 7531 1974
rect 7563 1942 7611 1974
rect 7483 1906 7611 1942
rect 7483 1874 7531 1906
rect 7563 1874 7611 1906
rect 7483 1838 7611 1874
rect 7483 1806 7531 1838
rect 7563 1806 7611 1838
rect 7483 1770 7611 1806
rect 7483 1738 7531 1770
rect 7563 1738 7611 1770
rect 7483 1702 7611 1738
rect 7483 1670 7531 1702
rect 7563 1670 7611 1702
rect 7483 1634 7611 1670
rect 7483 1602 7531 1634
rect 7563 1602 7611 1634
rect 7483 1566 7611 1602
rect 7483 1534 7531 1566
rect 7563 1534 7611 1566
rect 7483 1518 7611 1534
rect 7731 2382 7967 2398
rect 7731 2350 7833 2382
rect 7865 2350 7967 2382
rect 7731 2314 7967 2350
rect 7731 2282 7833 2314
rect 7865 2282 7967 2314
rect 7731 2246 7967 2282
rect 7731 2214 7833 2246
rect 7865 2214 7967 2246
rect 7731 2178 7967 2214
rect 7731 2146 7833 2178
rect 7865 2146 7967 2178
rect 7731 2110 7967 2146
rect 7731 2078 7833 2110
rect 7865 2078 7967 2110
rect 7731 2042 7967 2078
rect 7731 2010 7833 2042
rect 7865 2010 7967 2042
rect 7731 1974 7967 2010
rect 7731 1942 7833 1974
rect 7865 1942 7967 1974
rect 7731 1906 7967 1942
rect 7731 1874 7833 1906
rect 7865 1874 7967 1906
rect 7731 1838 7967 1874
rect 7731 1806 7833 1838
rect 7865 1806 7967 1838
rect 7731 1770 7967 1806
rect 7731 1738 7833 1770
rect 7865 1738 7967 1770
rect 7731 1702 7967 1738
rect 7731 1670 7833 1702
rect 7865 1670 7967 1702
rect 7731 1634 7967 1670
rect 7731 1602 7833 1634
rect 7865 1602 7967 1634
rect 7731 1566 7967 1602
rect 7731 1534 7833 1566
rect 7865 1534 7967 1566
rect 7731 1518 7967 1534
rect 8087 2382 8215 2398
rect 8087 2350 8135 2382
rect 8167 2350 8215 2382
rect 8087 2314 8215 2350
rect 8087 2282 8135 2314
rect 8167 2282 8215 2314
rect 8087 2246 8215 2282
rect 8087 2214 8135 2246
rect 8167 2214 8215 2246
rect 8087 2178 8215 2214
rect 8087 2146 8135 2178
rect 8167 2146 8215 2178
rect 8087 2110 8215 2146
rect 8087 2078 8135 2110
rect 8167 2078 8215 2110
rect 8087 2042 8215 2078
rect 8087 2010 8135 2042
rect 8167 2010 8215 2042
rect 8087 1974 8215 2010
rect 8087 1942 8135 1974
rect 8167 1942 8215 1974
rect 8087 1906 8215 1942
rect 8087 1874 8135 1906
rect 8167 1874 8215 1906
rect 8087 1838 8215 1874
rect 8087 1806 8135 1838
rect 8167 1806 8215 1838
rect 8087 1770 8215 1806
rect 8087 1738 8135 1770
rect 8167 1738 8215 1770
rect 8087 1702 8215 1738
rect 8087 1670 8135 1702
rect 8167 1670 8215 1702
rect 8087 1634 8215 1670
rect 8087 1602 8135 1634
rect 8167 1602 8215 1634
rect 8087 1566 8215 1602
rect 8087 1534 8135 1566
rect 8167 1534 8215 1566
rect 8087 1518 8215 1534
rect 8335 2382 8571 2398
rect 8335 2350 8437 2382
rect 8469 2350 8571 2382
rect 8335 2314 8571 2350
rect 8335 2282 8437 2314
rect 8469 2282 8571 2314
rect 8335 2246 8571 2282
rect 8335 2214 8437 2246
rect 8469 2214 8571 2246
rect 8335 2178 8571 2214
rect 8335 2146 8437 2178
rect 8469 2146 8571 2178
rect 8335 2110 8571 2146
rect 8335 2078 8437 2110
rect 8469 2078 8571 2110
rect 8335 2042 8571 2078
rect 8335 2010 8437 2042
rect 8469 2010 8571 2042
rect 8335 1974 8571 2010
rect 8335 1942 8437 1974
rect 8469 1942 8571 1974
rect 8335 1906 8571 1942
rect 8335 1874 8437 1906
rect 8469 1874 8571 1906
rect 8335 1838 8571 1874
rect 8335 1806 8437 1838
rect 8469 1806 8571 1838
rect 8335 1770 8571 1806
rect 8335 1738 8437 1770
rect 8469 1738 8571 1770
rect 8335 1702 8571 1738
rect 8335 1670 8437 1702
rect 8469 1670 8571 1702
rect 8335 1634 8571 1670
rect 8335 1602 8437 1634
rect 8469 1602 8571 1634
rect 8335 1566 8571 1602
rect 8335 1534 8437 1566
rect 8469 1534 8571 1566
rect 8335 1518 8571 1534
rect 8691 2382 8819 2398
rect 8691 2350 8739 2382
rect 8771 2350 8819 2382
rect 8691 2314 8819 2350
rect 8691 2282 8739 2314
rect 8771 2282 8819 2314
rect 8691 2246 8819 2282
rect 8691 2214 8739 2246
rect 8771 2214 8819 2246
rect 8691 2178 8819 2214
rect 8691 2146 8739 2178
rect 8771 2146 8819 2178
rect 8691 2110 8819 2146
rect 8691 2078 8739 2110
rect 8771 2078 8819 2110
rect 8691 2042 8819 2078
rect 8691 2010 8739 2042
rect 8771 2010 8819 2042
rect 8691 1974 8819 2010
rect 8691 1942 8739 1974
rect 8771 1942 8819 1974
rect 8691 1906 8819 1942
rect 8691 1874 8739 1906
rect 8771 1874 8819 1906
rect 8691 1838 8819 1874
rect 8691 1806 8739 1838
rect 8771 1806 8819 1838
rect 8691 1770 8819 1806
rect 8691 1738 8739 1770
rect 8771 1738 8819 1770
rect 8691 1702 8819 1738
rect 8691 1670 8739 1702
rect 8771 1670 8819 1702
rect 8691 1634 8819 1670
rect 8691 1602 8739 1634
rect 8771 1602 8819 1634
rect 8691 1566 8819 1602
rect 8691 1534 8739 1566
rect 8771 1534 8819 1566
rect 8691 1518 8819 1534
rect 8939 2382 9175 2398
rect 8939 2350 9041 2382
rect 9073 2350 9175 2382
rect 8939 2314 9175 2350
rect 8939 2282 9041 2314
rect 9073 2282 9175 2314
rect 8939 2246 9175 2282
rect 8939 2214 9041 2246
rect 9073 2214 9175 2246
rect 8939 2178 9175 2214
rect 8939 2146 9041 2178
rect 9073 2146 9175 2178
rect 8939 2110 9175 2146
rect 8939 2078 9041 2110
rect 9073 2078 9175 2110
rect 8939 2042 9175 2078
rect 8939 2010 9041 2042
rect 9073 2010 9175 2042
rect 8939 1974 9175 2010
rect 8939 1942 9041 1974
rect 9073 1942 9175 1974
rect 8939 1906 9175 1942
rect 8939 1874 9041 1906
rect 9073 1874 9175 1906
rect 8939 1838 9175 1874
rect 8939 1806 9041 1838
rect 9073 1806 9175 1838
rect 8939 1770 9175 1806
rect 8939 1738 9041 1770
rect 9073 1738 9175 1770
rect 8939 1702 9175 1738
rect 8939 1670 9041 1702
rect 9073 1670 9175 1702
rect 8939 1634 9175 1670
rect 8939 1602 9041 1634
rect 9073 1602 9175 1634
rect 8939 1566 9175 1602
rect 8939 1534 9041 1566
rect 9073 1534 9175 1566
rect 8939 1518 9175 1534
rect 9295 2382 9423 2398
rect 9295 2350 9343 2382
rect 9375 2350 9423 2382
rect 9295 2314 9423 2350
rect 9295 2282 9343 2314
rect 9375 2282 9423 2314
rect 9295 2246 9423 2282
rect 9295 2214 9343 2246
rect 9375 2214 9423 2246
rect 9295 2178 9423 2214
rect 9295 2146 9343 2178
rect 9375 2146 9423 2178
rect 9295 2110 9423 2146
rect 9295 2078 9343 2110
rect 9375 2078 9423 2110
rect 9295 2042 9423 2078
rect 9295 2010 9343 2042
rect 9375 2010 9423 2042
rect 9295 1974 9423 2010
rect 9295 1942 9343 1974
rect 9375 1942 9423 1974
rect 9295 1906 9423 1942
rect 9295 1874 9343 1906
rect 9375 1874 9423 1906
rect 9295 1838 9423 1874
rect 9295 1806 9343 1838
rect 9375 1806 9423 1838
rect 9295 1770 9423 1806
rect 9295 1738 9343 1770
rect 9375 1738 9423 1770
rect 9295 1702 9423 1738
rect 9295 1670 9343 1702
rect 9375 1670 9423 1702
rect 9295 1634 9423 1670
rect 9295 1602 9343 1634
rect 9375 1602 9423 1634
rect 9295 1566 9423 1602
rect 9295 1534 9343 1566
rect 9375 1534 9423 1566
rect 9295 1518 9423 1534
rect 9543 2382 9779 2398
rect 9543 2350 9645 2382
rect 9677 2350 9779 2382
rect 9543 2314 9779 2350
rect 9543 2282 9645 2314
rect 9677 2282 9779 2314
rect 9543 2246 9779 2282
rect 9543 2214 9645 2246
rect 9677 2214 9779 2246
rect 9543 2178 9779 2214
rect 9543 2146 9645 2178
rect 9677 2146 9779 2178
rect 9543 2110 9779 2146
rect 9543 2078 9645 2110
rect 9677 2078 9779 2110
rect 9543 2042 9779 2078
rect 9543 2010 9645 2042
rect 9677 2010 9779 2042
rect 9543 1974 9779 2010
rect 9543 1942 9645 1974
rect 9677 1942 9779 1974
rect 9543 1906 9779 1942
rect 9543 1874 9645 1906
rect 9677 1874 9779 1906
rect 9543 1838 9779 1874
rect 9543 1806 9645 1838
rect 9677 1806 9779 1838
rect 9543 1770 9779 1806
rect 9543 1738 9645 1770
rect 9677 1738 9779 1770
rect 9543 1702 9779 1738
rect 9543 1670 9645 1702
rect 9677 1670 9779 1702
rect 9543 1634 9779 1670
rect 9543 1602 9645 1634
rect 9677 1602 9779 1634
rect 9543 1566 9779 1602
rect 9543 1534 9645 1566
rect 9677 1534 9779 1566
rect 9543 1518 9779 1534
rect 9899 2382 10027 2398
rect 9899 2350 9947 2382
rect 9979 2350 10027 2382
rect 9899 2314 10027 2350
rect 9899 2282 9947 2314
rect 9979 2282 10027 2314
rect 9899 2246 10027 2282
rect 9899 2214 9947 2246
rect 9979 2214 10027 2246
rect 9899 2178 10027 2214
rect 9899 2146 9947 2178
rect 9979 2146 10027 2178
rect 9899 2110 10027 2146
rect 9899 2078 9947 2110
rect 9979 2078 10027 2110
rect 9899 2042 10027 2078
rect 9899 2010 9947 2042
rect 9979 2010 10027 2042
rect 9899 1974 10027 2010
rect 9899 1942 9947 1974
rect 9979 1942 10027 1974
rect 9899 1906 10027 1942
rect 9899 1874 9947 1906
rect 9979 1874 10027 1906
rect 9899 1838 10027 1874
rect 9899 1806 9947 1838
rect 9979 1806 10027 1838
rect 9899 1770 10027 1806
rect 9899 1738 9947 1770
rect 9979 1738 10027 1770
rect 9899 1702 10027 1738
rect 9899 1670 9947 1702
rect 9979 1670 10027 1702
rect 9899 1634 10027 1670
rect 9899 1602 9947 1634
rect 9979 1602 10027 1634
rect 9899 1566 10027 1602
rect 9899 1534 9947 1566
rect 9979 1534 10027 1566
rect 9899 1518 10027 1534
rect 10147 2382 10383 2398
rect 10147 2350 10249 2382
rect 10281 2350 10383 2382
rect 10147 2314 10383 2350
rect 10147 2282 10249 2314
rect 10281 2282 10383 2314
rect 10147 2246 10383 2282
rect 10147 2214 10249 2246
rect 10281 2214 10383 2246
rect 10147 2178 10383 2214
rect 10147 2146 10249 2178
rect 10281 2146 10383 2178
rect 10147 2110 10383 2146
rect 10147 2078 10249 2110
rect 10281 2078 10383 2110
rect 10147 2042 10383 2078
rect 10147 2010 10249 2042
rect 10281 2010 10383 2042
rect 10147 1974 10383 2010
rect 10147 1942 10249 1974
rect 10281 1942 10383 1974
rect 10147 1906 10383 1942
rect 10147 1874 10249 1906
rect 10281 1874 10383 1906
rect 10147 1838 10383 1874
rect 10147 1806 10249 1838
rect 10281 1806 10383 1838
rect 10147 1770 10383 1806
rect 10147 1738 10249 1770
rect 10281 1738 10383 1770
rect 10147 1702 10383 1738
rect 10147 1670 10249 1702
rect 10281 1670 10383 1702
rect 10147 1634 10383 1670
rect 10147 1602 10249 1634
rect 10281 1602 10383 1634
rect 10147 1566 10383 1602
rect 10147 1534 10249 1566
rect 10281 1534 10383 1566
rect 10147 1518 10383 1534
rect 10503 2382 10631 2398
rect 10503 2350 10551 2382
rect 10583 2350 10631 2382
rect 10503 2314 10631 2350
rect 10503 2282 10551 2314
rect 10583 2282 10631 2314
rect 10503 2246 10631 2282
rect 10503 2214 10551 2246
rect 10583 2214 10631 2246
rect 10503 2178 10631 2214
rect 10503 2146 10551 2178
rect 10583 2146 10631 2178
rect 10503 2110 10631 2146
rect 10503 2078 10551 2110
rect 10583 2078 10631 2110
rect 10503 2042 10631 2078
rect 10503 2010 10551 2042
rect 10583 2010 10631 2042
rect 10503 1974 10631 2010
rect 10503 1942 10551 1974
rect 10583 1942 10631 1974
rect 10503 1906 10631 1942
rect 10503 1874 10551 1906
rect 10583 1874 10631 1906
rect 10503 1838 10631 1874
rect 10503 1806 10551 1838
rect 10583 1806 10631 1838
rect 10503 1770 10631 1806
rect 10503 1738 10551 1770
rect 10583 1738 10631 1770
rect 10503 1702 10631 1738
rect 10503 1670 10551 1702
rect 10583 1670 10631 1702
rect 10503 1634 10631 1670
rect 10503 1602 10551 1634
rect 10583 1602 10631 1634
rect 10503 1566 10631 1602
rect 10503 1534 10551 1566
rect 10583 1534 10631 1566
rect 10503 1518 10631 1534
rect 10751 2382 10987 2398
rect 10751 2350 10853 2382
rect 10885 2350 10987 2382
rect 10751 2314 10987 2350
rect 10751 2282 10853 2314
rect 10885 2282 10987 2314
rect 10751 2246 10987 2282
rect 10751 2214 10853 2246
rect 10885 2214 10987 2246
rect 10751 2178 10987 2214
rect 10751 2146 10853 2178
rect 10885 2146 10987 2178
rect 10751 2110 10987 2146
rect 10751 2078 10853 2110
rect 10885 2078 10987 2110
rect 10751 2042 10987 2078
rect 10751 2010 10853 2042
rect 10885 2010 10987 2042
rect 10751 1974 10987 2010
rect 10751 1942 10853 1974
rect 10885 1942 10987 1974
rect 10751 1906 10987 1942
rect 10751 1874 10853 1906
rect 10885 1874 10987 1906
rect 10751 1838 10987 1874
rect 10751 1806 10853 1838
rect 10885 1806 10987 1838
rect 10751 1770 10987 1806
rect 10751 1738 10853 1770
rect 10885 1738 10987 1770
rect 10751 1702 10987 1738
rect 10751 1670 10853 1702
rect 10885 1670 10987 1702
rect 10751 1634 10987 1670
rect 10751 1602 10853 1634
rect 10885 1602 10987 1634
rect 10751 1566 10987 1602
rect 10751 1534 10853 1566
rect 10885 1534 10987 1566
rect 10751 1518 10987 1534
rect 11107 2382 11235 2398
rect 11107 2350 11155 2382
rect 11187 2350 11235 2382
rect 11107 2314 11235 2350
rect 11107 2282 11155 2314
rect 11187 2282 11235 2314
rect 11107 2246 11235 2282
rect 11107 2214 11155 2246
rect 11187 2214 11235 2246
rect 11107 2178 11235 2214
rect 11107 2146 11155 2178
rect 11187 2146 11235 2178
rect 11107 2110 11235 2146
rect 11107 2078 11155 2110
rect 11187 2078 11235 2110
rect 11107 2042 11235 2078
rect 11107 2010 11155 2042
rect 11187 2010 11235 2042
rect 11107 1974 11235 2010
rect 11107 1942 11155 1974
rect 11187 1942 11235 1974
rect 11107 1906 11235 1942
rect 11107 1874 11155 1906
rect 11187 1874 11235 1906
rect 11107 1838 11235 1874
rect 11107 1806 11155 1838
rect 11187 1806 11235 1838
rect 11107 1770 11235 1806
rect 11107 1738 11155 1770
rect 11187 1738 11235 1770
rect 11107 1702 11235 1738
rect 11107 1670 11155 1702
rect 11187 1670 11235 1702
rect 11107 1634 11235 1670
rect 11107 1602 11155 1634
rect 11187 1602 11235 1634
rect 11107 1566 11235 1602
rect 11107 1534 11155 1566
rect 11187 1534 11235 1566
rect 11107 1518 11235 1534
rect 11355 2382 11591 2398
rect 11355 2350 11457 2382
rect 11489 2350 11591 2382
rect 11355 2314 11591 2350
rect 11355 2282 11457 2314
rect 11489 2282 11591 2314
rect 11355 2246 11591 2282
rect 11355 2214 11457 2246
rect 11489 2214 11591 2246
rect 11355 2178 11591 2214
rect 11355 2146 11457 2178
rect 11489 2146 11591 2178
rect 11355 2110 11591 2146
rect 11355 2078 11457 2110
rect 11489 2078 11591 2110
rect 11355 2042 11591 2078
rect 11355 2010 11457 2042
rect 11489 2010 11591 2042
rect 11355 1974 11591 2010
rect 11355 1942 11457 1974
rect 11489 1942 11591 1974
rect 11355 1906 11591 1942
rect 11355 1874 11457 1906
rect 11489 1874 11591 1906
rect 11355 1838 11591 1874
rect 11355 1806 11457 1838
rect 11489 1806 11591 1838
rect 11355 1770 11591 1806
rect 11355 1738 11457 1770
rect 11489 1738 11591 1770
rect 11355 1702 11591 1738
rect 11355 1670 11457 1702
rect 11489 1670 11591 1702
rect 11355 1634 11591 1670
rect 11355 1602 11457 1634
rect 11489 1602 11591 1634
rect 11355 1566 11591 1602
rect 11355 1534 11457 1566
rect 11489 1534 11591 1566
rect 11355 1518 11591 1534
rect 11711 2382 11839 2398
rect 11711 2350 11759 2382
rect 11791 2350 11839 2382
rect 11711 2314 11839 2350
rect 11711 2282 11759 2314
rect 11791 2282 11839 2314
rect 11711 2246 11839 2282
rect 11711 2214 11759 2246
rect 11791 2214 11839 2246
rect 11711 2178 11839 2214
rect 11711 2146 11759 2178
rect 11791 2146 11839 2178
rect 11711 2110 11839 2146
rect 11711 2078 11759 2110
rect 11791 2078 11839 2110
rect 11711 2042 11839 2078
rect 11711 2010 11759 2042
rect 11791 2010 11839 2042
rect 11711 1974 11839 2010
rect 11711 1942 11759 1974
rect 11791 1942 11839 1974
rect 11711 1906 11839 1942
rect 11711 1874 11759 1906
rect 11791 1874 11839 1906
rect 11711 1838 11839 1874
rect 11711 1806 11759 1838
rect 11791 1806 11839 1838
rect 11711 1770 11839 1806
rect 11711 1738 11759 1770
rect 11791 1738 11839 1770
rect 11711 1702 11839 1738
rect 11711 1670 11759 1702
rect 11791 1670 11839 1702
rect 11711 1634 11839 1670
rect 11711 1602 11759 1634
rect 11791 1602 11839 1634
rect 11711 1566 11839 1602
rect 11711 1534 11759 1566
rect 11791 1534 11839 1566
rect 11711 1518 11839 1534
rect 11959 2382 12195 2398
rect 11959 2350 12061 2382
rect 12093 2350 12195 2382
rect 11959 2314 12195 2350
rect 11959 2282 12061 2314
rect 12093 2282 12195 2314
rect 11959 2246 12195 2282
rect 11959 2214 12061 2246
rect 12093 2214 12195 2246
rect 11959 2178 12195 2214
rect 11959 2146 12061 2178
rect 12093 2146 12195 2178
rect 11959 2110 12195 2146
rect 11959 2078 12061 2110
rect 12093 2078 12195 2110
rect 11959 2042 12195 2078
rect 11959 2010 12061 2042
rect 12093 2010 12195 2042
rect 11959 1974 12195 2010
rect 11959 1942 12061 1974
rect 12093 1942 12195 1974
rect 11959 1906 12195 1942
rect 11959 1874 12061 1906
rect 12093 1874 12195 1906
rect 11959 1838 12195 1874
rect 11959 1806 12061 1838
rect 12093 1806 12195 1838
rect 11959 1770 12195 1806
rect 11959 1738 12061 1770
rect 12093 1738 12195 1770
rect 11959 1702 12195 1738
rect 11959 1670 12061 1702
rect 12093 1670 12195 1702
rect 11959 1634 12195 1670
rect 11959 1602 12061 1634
rect 12093 1602 12195 1634
rect 11959 1566 12195 1602
rect 11959 1534 12061 1566
rect 12093 1534 12195 1566
rect 11959 1518 12195 1534
rect 12315 2382 12443 2398
rect 12315 2350 12363 2382
rect 12395 2350 12443 2382
rect 12315 2314 12443 2350
rect 12315 2282 12363 2314
rect 12395 2282 12443 2314
rect 12315 2246 12443 2282
rect 12315 2214 12363 2246
rect 12395 2214 12443 2246
rect 12315 2178 12443 2214
rect 12315 2146 12363 2178
rect 12395 2146 12443 2178
rect 12315 2110 12443 2146
rect 12315 2078 12363 2110
rect 12395 2078 12443 2110
rect 12315 2042 12443 2078
rect 12315 2010 12363 2042
rect 12395 2010 12443 2042
rect 12315 1974 12443 2010
rect 12315 1942 12363 1974
rect 12395 1942 12443 1974
rect 12315 1906 12443 1942
rect 12315 1874 12363 1906
rect 12395 1874 12443 1906
rect 12315 1838 12443 1874
rect 12315 1806 12363 1838
rect 12395 1806 12443 1838
rect 12315 1770 12443 1806
rect 12315 1738 12363 1770
rect 12395 1738 12443 1770
rect 12315 1702 12443 1738
rect 12315 1670 12363 1702
rect 12395 1670 12443 1702
rect 12315 1634 12443 1670
rect 12315 1602 12363 1634
rect 12395 1602 12443 1634
rect 12315 1566 12443 1602
rect 12315 1534 12363 1566
rect 12395 1534 12443 1566
rect 12315 1518 12443 1534
rect 12563 2382 12799 2398
rect 12563 2350 12665 2382
rect 12697 2350 12799 2382
rect 12563 2314 12799 2350
rect 12563 2282 12665 2314
rect 12697 2282 12799 2314
rect 12563 2246 12799 2282
rect 12563 2214 12665 2246
rect 12697 2214 12799 2246
rect 12563 2178 12799 2214
rect 12563 2146 12665 2178
rect 12697 2146 12799 2178
rect 12563 2110 12799 2146
rect 12563 2078 12665 2110
rect 12697 2078 12799 2110
rect 12563 2042 12799 2078
rect 12563 2010 12665 2042
rect 12697 2010 12799 2042
rect 12563 1974 12799 2010
rect 12563 1942 12665 1974
rect 12697 1942 12799 1974
rect 12563 1906 12799 1942
rect 12563 1874 12665 1906
rect 12697 1874 12799 1906
rect 12563 1838 12799 1874
rect 12563 1806 12665 1838
rect 12697 1806 12799 1838
rect 12563 1770 12799 1806
rect 12563 1738 12665 1770
rect 12697 1738 12799 1770
rect 12563 1702 12799 1738
rect 12563 1670 12665 1702
rect 12697 1670 12799 1702
rect 12563 1634 12799 1670
rect 12563 1602 12665 1634
rect 12697 1602 12799 1634
rect 12563 1566 12799 1602
rect 12563 1534 12665 1566
rect 12697 1534 12799 1566
rect 12563 1518 12799 1534
rect 12919 2382 13047 2398
rect 12919 2350 12967 2382
rect 12999 2350 13047 2382
rect 12919 2314 13047 2350
rect 12919 2282 12967 2314
rect 12999 2282 13047 2314
rect 12919 2246 13047 2282
rect 12919 2214 12967 2246
rect 12999 2214 13047 2246
rect 12919 2178 13047 2214
rect 12919 2146 12967 2178
rect 12999 2146 13047 2178
rect 12919 2110 13047 2146
rect 12919 2078 12967 2110
rect 12999 2078 13047 2110
rect 12919 2042 13047 2078
rect 12919 2010 12967 2042
rect 12999 2010 13047 2042
rect 12919 1974 13047 2010
rect 12919 1942 12967 1974
rect 12999 1942 13047 1974
rect 12919 1906 13047 1942
rect 12919 1874 12967 1906
rect 12999 1874 13047 1906
rect 12919 1838 13047 1874
rect 12919 1806 12967 1838
rect 12999 1806 13047 1838
rect 12919 1770 13047 1806
rect 12919 1738 12967 1770
rect 12999 1738 13047 1770
rect 12919 1702 13047 1738
rect 12919 1670 12967 1702
rect 12999 1670 13047 1702
rect 12919 1634 13047 1670
rect 12919 1602 12967 1634
rect 12999 1602 13047 1634
rect 12919 1566 13047 1602
rect 12919 1534 12967 1566
rect 12999 1534 13047 1566
rect 12919 1518 13047 1534
rect 13167 2382 13403 2398
rect 13167 2350 13269 2382
rect 13301 2350 13403 2382
rect 13167 2314 13403 2350
rect 13167 2282 13269 2314
rect 13301 2282 13403 2314
rect 13167 2246 13403 2282
rect 13167 2214 13269 2246
rect 13301 2214 13403 2246
rect 13167 2178 13403 2214
rect 13167 2146 13269 2178
rect 13301 2146 13403 2178
rect 13167 2110 13403 2146
rect 13167 2078 13269 2110
rect 13301 2078 13403 2110
rect 13167 2042 13403 2078
rect 13167 2010 13269 2042
rect 13301 2010 13403 2042
rect 13167 1974 13403 2010
rect 13167 1942 13269 1974
rect 13301 1942 13403 1974
rect 13167 1906 13403 1942
rect 13167 1874 13269 1906
rect 13301 1874 13403 1906
rect 13167 1838 13403 1874
rect 13167 1806 13269 1838
rect 13301 1806 13403 1838
rect 13167 1770 13403 1806
rect 13167 1738 13269 1770
rect 13301 1738 13403 1770
rect 13167 1702 13403 1738
rect 13167 1670 13269 1702
rect 13301 1670 13403 1702
rect 13167 1634 13403 1670
rect 13167 1602 13269 1634
rect 13301 1602 13403 1634
rect 13167 1566 13403 1602
rect 13167 1534 13269 1566
rect 13301 1534 13403 1566
rect 13167 1518 13403 1534
rect 13523 2382 13651 2398
rect 13523 2350 13571 2382
rect 13603 2350 13651 2382
rect 13523 2314 13651 2350
rect 13523 2282 13571 2314
rect 13603 2282 13651 2314
rect 13523 2246 13651 2282
rect 13523 2214 13571 2246
rect 13603 2214 13651 2246
rect 13523 2178 13651 2214
rect 13523 2146 13571 2178
rect 13603 2146 13651 2178
rect 13523 2110 13651 2146
rect 13523 2078 13571 2110
rect 13603 2078 13651 2110
rect 13523 2042 13651 2078
rect 13523 2010 13571 2042
rect 13603 2010 13651 2042
rect 13523 1974 13651 2010
rect 13523 1942 13571 1974
rect 13603 1942 13651 1974
rect 13523 1906 13651 1942
rect 13523 1874 13571 1906
rect 13603 1874 13651 1906
rect 13523 1838 13651 1874
rect 13523 1806 13571 1838
rect 13603 1806 13651 1838
rect 13523 1770 13651 1806
rect 13523 1738 13571 1770
rect 13603 1738 13651 1770
rect 13523 1702 13651 1738
rect 13523 1670 13571 1702
rect 13603 1670 13651 1702
rect 13523 1634 13651 1670
rect 13523 1602 13571 1634
rect 13603 1602 13651 1634
rect 13523 1566 13651 1602
rect 13523 1534 13571 1566
rect 13603 1534 13651 1566
rect 13523 1518 13651 1534
rect 13771 2382 14007 2398
rect 13771 2350 13873 2382
rect 13905 2350 14007 2382
rect 13771 2314 14007 2350
rect 13771 2282 13873 2314
rect 13905 2282 14007 2314
rect 13771 2246 14007 2282
rect 13771 2214 13873 2246
rect 13905 2214 14007 2246
rect 13771 2178 14007 2214
rect 13771 2146 13873 2178
rect 13905 2146 14007 2178
rect 13771 2110 14007 2146
rect 13771 2078 13873 2110
rect 13905 2078 14007 2110
rect 13771 2042 14007 2078
rect 13771 2010 13873 2042
rect 13905 2010 14007 2042
rect 13771 1974 14007 2010
rect 13771 1942 13873 1974
rect 13905 1942 14007 1974
rect 13771 1906 14007 1942
rect 13771 1874 13873 1906
rect 13905 1874 14007 1906
rect 13771 1838 14007 1874
rect 13771 1806 13873 1838
rect 13905 1806 14007 1838
rect 13771 1770 14007 1806
rect 13771 1738 13873 1770
rect 13905 1738 14007 1770
rect 13771 1702 14007 1738
rect 13771 1670 13873 1702
rect 13905 1670 14007 1702
rect 13771 1634 14007 1670
rect 13771 1602 13873 1634
rect 13905 1602 14007 1634
rect 13771 1566 14007 1602
rect 13771 1534 13873 1566
rect 13905 1534 14007 1566
rect 13771 1518 14007 1534
rect 14127 2382 14255 2398
rect 14127 2350 14175 2382
rect 14207 2350 14255 2382
rect 14127 2314 14255 2350
rect 14127 2282 14175 2314
rect 14207 2282 14255 2314
rect 14127 2246 14255 2282
rect 14127 2214 14175 2246
rect 14207 2214 14255 2246
rect 14127 2178 14255 2214
rect 14127 2146 14175 2178
rect 14207 2146 14255 2178
rect 14127 2110 14255 2146
rect 14127 2078 14175 2110
rect 14207 2078 14255 2110
rect 14127 2042 14255 2078
rect 14127 2010 14175 2042
rect 14207 2010 14255 2042
rect 14127 1974 14255 2010
rect 14127 1942 14175 1974
rect 14207 1942 14255 1974
rect 14127 1906 14255 1942
rect 14127 1874 14175 1906
rect 14207 1874 14255 1906
rect 14127 1838 14255 1874
rect 14127 1806 14175 1838
rect 14207 1806 14255 1838
rect 14127 1770 14255 1806
rect 14127 1738 14175 1770
rect 14207 1738 14255 1770
rect 14127 1702 14255 1738
rect 14127 1670 14175 1702
rect 14207 1670 14255 1702
rect 14127 1634 14255 1670
rect 14127 1602 14175 1634
rect 14207 1602 14255 1634
rect 14127 1566 14255 1602
rect 14127 1534 14175 1566
rect 14207 1534 14255 1566
rect 14127 1518 14255 1534
rect 14375 2382 14523 2398
rect 14375 2350 14477 2382
rect 14509 2350 14523 2382
rect 14375 2314 14523 2350
rect 14375 2282 14477 2314
rect 14509 2282 14523 2314
rect 14375 2246 14523 2282
rect 14375 2214 14477 2246
rect 14509 2214 14523 2246
rect 14375 2178 14523 2214
rect 14375 2146 14477 2178
rect 14509 2146 14523 2178
rect 14375 2110 14523 2146
rect 14375 2078 14477 2110
rect 14509 2078 14523 2110
rect 14375 2042 14523 2078
rect 14375 2010 14477 2042
rect 14509 2010 14523 2042
rect 14375 1974 14523 2010
rect 14375 1942 14477 1974
rect 14509 1942 14523 1974
rect 14375 1906 14523 1942
rect 14375 1874 14477 1906
rect 14509 1874 14523 1906
rect 14375 1838 14523 1874
rect 14375 1806 14477 1838
rect 14509 1806 14523 1838
rect 14375 1770 14523 1806
rect 14375 1738 14477 1770
rect 14509 1738 14523 1770
rect 14375 1702 14523 1738
rect 14375 1670 14477 1702
rect 14509 1670 14523 1702
rect 14375 1634 14523 1670
rect 14375 1602 14477 1634
rect 14509 1602 14523 1634
rect 14375 1566 14523 1602
rect 14375 1534 14477 1566
rect 14509 1534 14523 1566
rect 14375 1518 14523 1534
rect 1477 1414 1571 1430
rect 1477 1382 1491 1414
rect 1523 1382 1571 1414
rect 1477 1346 1571 1382
rect 1477 1314 1491 1346
rect 1523 1314 1571 1346
rect 1477 1278 1571 1314
rect 1477 1246 1491 1278
rect 1523 1246 1571 1278
rect 1477 1210 1571 1246
rect 1477 1178 1491 1210
rect 1523 1178 1571 1210
rect 1477 1142 1571 1178
rect 1477 1110 1491 1142
rect 1523 1110 1571 1142
rect 1477 1074 1571 1110
rect 1477 1042 1491 1074
rect 1523 1042 1571 1074
rect 1477 1006 1571 1042
rect 1477 974 1491 1006
rect 1523 974 1571 1006
rect 1477 938 1571 974
rect 1477 906 1491 938
rect 1523 906 1571 938
rect 1477 870 1571 906
rect 1477 838 1491 870
rect 1523 838 1571 870
rect 1477 802 1571 838
rect 1477 770 1491 802
rect 1523 770 1571 802
rect 1477 734 1571 770
rect 1477 702 1491 734
rect 1523 702 1571 734
rect 1477 666 1571 702
rect 1477 634 1491 666
rect 1523 634 1571 666
rect 1477 598 1571 634
rect 1477 566 1491 598
rect 1523 566 1571 598
rect 1477 550 1571 566
rect 1691 1414 1927 1430
rect 1691 1382 1793 1414
rect 1825 1382 1927 1414
rect 1691 1346 1927 1382
rect 1691 1314 1793 1346
rect 1825 1314 1927 1346
rect 1691 1278 1927 1314
rect 1691 1246 1793 1278
rect 1825 1246 1927 1278
rect 1691 1210 1927 1246
rect 1691 1178 1793 1210
rect 1825 1178 1927 1210
rect 1691 1142 1927 1178
rect 1691 1110 1793 1142
rect 1825 1110 1927 1142
rect 1691 1074 1927 1110
rect 1691 1042 1793 1074
rect 1825 1042 1927 1074
rect 1691 1006 1927 1042
rect 1691 974 1793 1006
rect 1825 974 1927 1006
rect 1691 938 1927 974
rect 1691 906 1793 938
rect 1825 906 1927 938
rect 1691 870 1927 906
rect 1691 838 1793 870
rect 1825 838 1927 870
rect 1691 802 1927 838
rect 1691 770 1793 802
rect 1825 770 1927 802
rect 1691 734 1927 770
rect 1691 702 1793 734
rect 1825 702 1927 734
rect 1691 666 1927 702
rect 1691 634 1793 666
rect 1825 634 1927 666
rect 1691 598 1927 634
rect 1691 566 1793 598
rect 1825 566 1927 598
rect 1691 550 1927 566
rect 2047 1414 2175 1430
rect 2047 1382 2095 1414
rect 2127 1382 2175 1414
rect 2047 1346 2175 1382
rect 2047 1314 2095 1346
rect 2127 1314 2175 1346
rect 2047 1278 2175 1314
rect 2047 1246 2095 1278
rect 2127 1246 2175 1278
rect 2047 1210 2175 1246
rect 2047 1178 2095 1210
rect 2127 1178 2175 1210
rect 2047 1142 2175 1178
rect 2047 1110 2095 1142
rect 2127 1110 2175 1142
rect 2047 1074 2175 1110
rect 2047 1042 2095 1074
rect 2127 1042 2175 1074
rect 2047 1006 2175 1042
rect 2047 974 2095 1006
rect 2127 974 2175 1006
rect 2047 938 2175 974
rect 2047 906 2095 938
rect 2127 906 2175 938
rect 2047 870 2175 906
rect 2047 838 2095 870
rect 2127 838 2175 870
rect 2047 802 2175 838
rect 2047 770 2095 802
rect 2127 770 2175 802
rect 2047 734 2175 770
rect 2047 702 2095 734
rect 2127 702 2175 734
rect 2047 666 2175 702
rect 2047 634 2095 666
rect 2127 634 2175 666
rect 2047 598 2175 634
rect 2047 566 2095 598
rect 2127 566 2175 598
rect 2047 550 2175 566
rect 2295 1414 2531 1430
rect 2295 1382 2397 1414
rect 2429 1382 2531 1414
rect 2295 1346 2531 1382
rect 2295 1314 2397 1346
rect 2429 1314 2531 1346
rect 2295 1278 2531 1314
rect 2295 1246 2397 1278
rect 2429 1246 2531 1278
rect 2295 1210 2531 1246
rect 2295 1178 2397 1210
rect 2429 1178 2531 1210
rect 2295 1142 2531 1178
rect 2295 1110 2397 1142
rect 2429 1110 2531 1142
rect 2295 1074 2531 1110
rect 2295 1042 2397 1074
rect 2429 1042 2531 1074
rect 2295 1006 2531 1042
rect 2295 974 2397 1006
rect 2429 974 2531 1006
rect 2295 938 2531 974
rect 2295 906 2397 938
rect 2429 906 2531 938
rect 2295 870 2531 906
rect 2295 838 2397 870
rect 2429 838 2531 870
rect 2295 802 2531 838
rect 2295 770 2397 802
rect 2429 770 2531 802
rect 2295 734 2531 770
rect 2295 702 2397 734
rect 2429 702 2531 734
rect 2295 666 2531 702
rect 2295 634 2397 666
rect 2429 634 2531 666
rect 2295 598 2531 634
rect 2295 566 2397 598
rect 2429 566 2531 598
rect 2295 550 2531 566
rect 2651 1414 2779 1430
rect 2651 1382 2699 1414
rect 2731 1382 2779 1414
rect 2651 1346 2779 1382
rect 2651 1314 2699 1346
rect 2731 1314 2779 1346
rect 2651 1278 2779 1314
rect 2651 1246 2699 1278
rect 2731 1246 2779 1278
rect 2651 1210 2779 1246
rect 2651 1178 2699 1210
rect 2731 1178 2779 1210
rect 2651 1142 2779 1178
rect 2651 1110 2699 1142
rect 2731 1110 2779 1142
rect 2651 1074 2779 1110
rect 2651 1042 2699 1074
rect 2731 1042 2779 1074
rect 2651 1006 2779 1042
rect 2651 974 2699 1006
rect 2731 974 2779 1006
rect 2651 938 2779 974
rect 2651 906 2699 938
rect 2731 906 2779 938
rect 2651 870 2779 906
rect 2651 838 2699 870
rect 2731 838 2779 870
rect 2651 802 2779 838
rect 2651 770 2699 802
rect 2731 770 2779 802
rect 2651 734 2779 770
rect 2651 702 2699 734
rect 2731 702 2779 734
rect 2651 666 2779 702
rect 2651 634 2699 666
rect 2731 634 2779 666
rect 2651 598 2779 634
rect 2651 566 2699 598
rect 2731 566 2779 598
rect 2651 550 2779 566
rect 2899 1414 3135 1430
rect 2899 1382 3001 1414
rect 3033 1382 3135 1414
rect 2899 1346 3135 1382
rect 2899 1314 3001 1346
rect 3033 1314 3135 1346
rect 2899 1278 3135 1314
rect 2899 1246 3001 1278
rect 3033 1246 3135 1278
rect 2899 1210 3135 1246
rect 2899 1178 3001 1210
rect 3033 1178 3135 1210
rect 2899 1142 3135 1178
rect 2899 1110 3001 1142
rect 3033 1110 3135 1142
rect 2899 1074 3135 1110
rect 2899 1042 3001 1074
rect 3033 1042 3135 1074
rect 2899 1006 3135 1042
rect 2899 974 3001 1006
rect 3033 974 3135 1006
rect 2899 938 3135 974
rect 2899 906 3001 938
rect 3033 906 3135 938
rect 2899 870 3135 906
rect 2899 838 3001 870
rect 3033 838 3135 870
rect 2899 802 3135 838
rect 2899 770 3001 802
rect 3033 770 3135 802
rect 2899 734 3135 770
rect 2899 702 3001 734
rect 3033 702 3135 734
rect 2899 666 3135 702
rect 2899 634 3001 666
rect 3033 634 3135 666
rect 2899 598 3135 634
rect 2899 566 3001 598
rect 3033 566 3135 598
rect 2899 550 3135 566
rect 3255 1414 3383 1430
rect 3255 1382 3303 1414
rect 3335 1382 3383 1414
rect 3255 1346 3383 1382
rect 3255 1314 3303 1346
rect 3335 1314 3383 1346
rect 3255 1278 3383 1314
rect 3255 1246 3303 1278
rect 3335 1246 3383 1278
rect 3255 1210 3383 1246
rect 3255 1178 3303 1210
rect 3335 1178 3383 1210
rect 3255 1142 3383 1178
rect 3255 1110 3303 1142
rect 3335 1110 3383 1142
rect 3255 1074 3383 1110
rect 3255 1042 3303 1074
rect 3335 1042 3383 1074
rect 3255 1006 3383 1042
rect 3255 974 3303 1006
rect 3335 974 3383 1006
rect 3255 938 3383 974
rect 3255 906 3303 938
rect 3335 906 3383 938
rect 3255 870 3383 906
rect 3255 838 3303 870
rect 3335 838 3383 870
rect 3255 802 3383 838
rect 3255 770 3303 802
rect 3335 770 3383 802
rect 3255 734 3383 770
rect 3255 702 3303 734
rect 3335 702 3383 734
rect 3255 666 3383 702
rect 3255 634 3303 666
rect 3335 634 3383 666
rect 3255 598 3383 634
rect 3255 566 3303 598
rect 3335 566 3383 598
rect 3255 550 3383 566
rect 3503 1414 3739 1430
rect 3503 1382 3605 1414
rect 3637 1382 3739 1414
rect 3503 1346 3739 1382
rect 3503 1314 3605 1346
rect 3637 1314 3739 1346
rect 3503 1278 3739 1314
rect 3503 1246 3605 1278
rect 3637 1246 3739 1278
rect 3503 1210 3739 1246
rect 3503 1178 3605 1210
rect 3637 1178 3739 1210
rect 3503 1142 3739 1178
rect 3503 1110 3605 1142
rect 3637 1110 3739 1142
rect 3503 1074 3739 1110
rect 3503 1042 3605 1074
rect 3637 1042 3739 1074
rect 3503 1006 3739 1042
rect 3503 974 3605 1006
rect 3637 974 3739 1006
rect 3503 938 3739 974
rect 3503 906 3605 938
rect 3637 906 3739 938
rect 3503 870 3739 906
rect 3503 838 3605 870
rect 3637 838 3739 870
rect 3503 802 3739 838
rect 3503 770 3605 802
rect 3637 770 3739 802
rect 3503 734 3739 770
rect 3503 702 3605 734
rect 3637 702 3739 734
rect 3503 666 3739 702
rect 3503 634 3605 666
rect 3637 634 3739 666
rect 3503 598 3739 634
rect 3503 566 3605 598
rect 3637 566 3739 598
rect 3503 550 3739 566
rect 3859 1414 3987 1430
rect 3859 1382 3907 1414
rect 3939 1382 3987 1414
rect 3859 1346 3987 1382
rect 3859 1314 3907 1346
rect 3939 1314 3987 1346
rect 3859 1278 3987 1314
rect 3859 1246 3907 1278
rect 3939 1246 3987 1278
rect 3859 1210 3987 1246
rect 3859 1178 3907 1210
rect 3939 1178 3987 1210
rect 3859 1142 3987 1178
rect 3859 1110 3907 1142
rect 3939 1110 3987 1142
rect 3859 1074 3987 1110
rect 3859 1042 3907 1074
rect 3939 1042 3987 1074
rect 3859 1006 3987 1042
rect 3859 974 3907 1006
rect 3939 974 3987 1006
rect 3859 938 3987 974
rect 3859 906 3907 938
rect 3939 906 3987 938
rect 3859 870 3987 906
rect 3859 838 3907 870
rect 3939 838 3987 870
rect 3859 802 3987 838
rect 3859 770 3907 802
rect 3939 770 3987 802
rect 3859 734 3987 770
rect 3859 702 3907 734
rect 3939 702 3987 734
rect 3859 666 3987 702
rect 3859 634 3907 666
rect 3939 634 3987 666
rect 3859 598 3987 634
rect 3859 566 3907 598
rect 3939 566 3987 598
rect 3859 550 3987 566
rect 4107 1414 4343 1430
rect 4107 1382 4209 1414
rect 4241 1382 4343 1414
rect 4107 1346 4343 1382
rect 4107 1314 4209 1346
rect 4241 1314 4343 1346
rect 4107 1278 4343 1314
rect 4107 1246 4209 1278
rect 4241 1246 4343 1278
rect 4107 1210 4343 1246
rect 4107 1178 4209 1210
rect 4241 1178 4343 1210
rect 4107 1142 4343 1178
rect 4107 1110 4209 1142
rect 4241 1110 4343 1142
rect 4107 1074 4343 1110
rect 4107 1042 4209 1074
rect 4241 1042 4343 1074
rect 4107 1006 4343 1042
rect 4107 974 4209 1006
rect 4241 974 4343 1006
rect 4107 938 4343 974
rect 4107 906 4209 938
rect 4241 906 4343 938
rect 4107 870 4343 906
rect 4107 838 4209 870
rect 4241 838 4343 870
rect 4107 802 4343 838
rect 4107 770 4209 802
rect 4241 770 4343 802
rect 4107 734 4343 770
rect 4107 702 4209 734
rect 4241 702 4343 734
rect 4107 666 4343 702
rect 4107 634 4209 666
rect 4241 634 4343 666
rect 4107 598 4343 634
rect 4107 566 4209 598
rect 4241 566 4343 598
rect 4107 550 4343 566
rect 4463 1414 4591 1430
rect 4463 1382 4511 1414
rect 4543 1382 4591 1414
rect 4463 1346 4591 1382
rect 4463 1314 4511 1346
rect 4543 1314 4591 1346
rect 4463 1278 4591 1314
rect 4463 1246 4511 1278
rect 4543 1246 4591 1278
rect 4463 1210 4591 1246
rect 4463 1178 4511 1210
rect 4543 1178 4591 1210
rect 4463 1142 4591 1178
rect 4463 1110 4511 1142
rect 4543 1110 4591 1142
rect 4463 1074 4591 1110
rect 4463 1042 4511 1074
rect 4543 1042 4591 1074
rect 4463 1006 4591 1042
rect 4463 974 4511 1006
rect 4543 974 4591 1006
rect 4463 938 4591 974
rect 4463 906 4511 938
rect 4543 906 4591 938
rect 4463 870 4591 906
rect 4463 838 4511 870
rect 4543 838 4591 870
rect 4463 802 4591 838
rect 4463 770 4511 802
rect 4543 770 4591 802
rect 4463 734 4591 770
rect 4463 702 4511 734
rect 4543 702 4591 734
rect 4463 666 4591 702
rect 4463 634 4511 666
rect 4543 634 4591 666
rect 4463 598 4591 634
rect 4463 566 4511 598
rect 4543 566 4591 598
rect 4463 550 4591 566
rect 4711 1414 4947 1430
rect 4711 1382 4813 1414
rect 4845 1382 4947 1414
rect 4711 1346 4947 1382
rect 4711 1314 4813 1346
rect 4845 1314 4947 1346
rect 4711 1278 4947 1314
rect 4711 1246 4813 1278
rect 4845 1246 4947 1278
rect 4711 1210 4947 1246
rect 4711 1178 4813 1210
rect 4845 1178 4947 1210
rect 4711 1142 4947 1178
rect 4711 1110 4813 1142
rect 4845 1110 4947 1142
rect 4711 1074 4947 1110
rect 4711 1042 4813 1074
rect 4845 1042 4947 1074
rect 4711 1006 4947 1042
rect 4711 974 4813 1006
rect 4845 974 4947 1006
rect 4711 938 4947 974
rect 4711 906 4813 938
rect 4845 906 4947 938
rect 4711 870 4947 906
rect 4711 838 4813 870
rect 4845 838 4947 870
rect 4711 802 4947 838
rect 4711 770 4813 802
rect 4845 770 4947 802
rect 4711 734 4947 770
rect 4711 702 4813 734
rect 4845 702 4947 734
rect 4711 666 4947 702
rect 4711 634 4813 666
rect 4845 634 4947 666
rect 4711 598 4947 634
rect 4711 566 4813 598
rect 4845 566 4947 598
rect 4711 550 4947 566
rect 5067 1414 5195 1430
rect 5067 1382 5115 1414
rect 5147 1382 5195 1414
rect 5067 1346 5195 1382
rect 5067 1314 5115 1346
rect 5147 1314 5195 1346
rect 5067 1278 5195 1314
rect 5067 1246 5115 1278
rect 5147 1246 5195 1278
rect 5067 1210 5195 1246
rect 5067 1178 5115 1210
rect 5147 1178 5195 1210
rect 5067 1142 5195 1178
rect 5067 1110 5115 1142
rect 5147 1110 5195 1142
rect 5067 1074 5195 1110
rect 5067 1042 5115 1074
rect 5147 1042 5195 1074
rect 5067 1006 5195 1042
rect 5067 974 5115 1006
rect 5147 974 5195 1006
rect 5067 938 5195 974
rect 5067 906 5115 938
rect 5147 906 5195 938
rect 5067 870 5195 906
rect 5067 838 5115 870
rect 5147 838 5195 870
rect 5067 802 5195 838
rect 5067 770 5115 802
rect 5147 770 5195 802
rect 5067 734 5195 770
rect 5067 702 5115 734
rect 5147 702 5195 734
rect 5067 666 5195 702
rect 5067 634 5115 666
rect 5147 634 5195 666
rect 5067 598 5195 634
rect 5067 566 5115 598
rect 5147 566 5195 598
rect 5067 550 5195 566
rect 5315 1414 5551 1430
rect 5315 1382 5417 1414
rect 5449 1382 5551 1414
rect 5315 1346 5551 1382
rect 5315 1314 5417 1346
rect 5449 1314 5551 1346
rect 5315 1278 5551 1314
rect 5315 1246 5417 1278
rect 5449 1246 5551 1278
rect 5315 1210 5551 1246
rect 5315 1178 5417 1210
rect 5449 1178 5551 1210
rect 5315 1142 5551 1178
rect 5315 1110 5417 1142
rect 5449 1110 5551 1142
rect 5315 1074 5551 1110
rect 5315 1042 5417 1074
rect 5449 1042 5551 1074
rect 5315 1006 5551 1042
rect 5315 974 5417 1006
rect 5449 974 5551 1006
rect 5315 938 5551 974
rect 5315 906 5417 938
rect 5449 906 5551 938
rect 5315 870 5551 906
rect 5315 838 5417 870
rect 5449 838 5551 870
rect 5315 802 5551 838
rect 5315 770 5417 802
rect 5449 770 5551 802
rect 5315 734 5551 770
rect 5315 702 5417 734
rect 5449 702 5551 734
rect 5315 666 5551 702
rect 5315 634 5417 666
rect 5449 634 5551 666
rect 5315 598 5551 634
rect 5315 566 5417 598
rect 5449 566 5551 598
rect 5315 550 5551 566
rect 5671 1414 5799 1430
rect 5671 1382 5719 1414
rect 5751 1382 5799 1414
rect 5671 1346 5799 1382
rect 5671 1314 5719 1346
rect 5751 1314 5799 1346
rect 5671 1278 5799 1314
rect 5671 1246 5719 1278
rect 5751 1246 5799 1278
rect 5671 1210 5799 1246
rect 5671 1178 5719 1210
rect 5751 1178 5799 1210
rect 5671 1142 5799 1178
rect 5671 1110 5719 1142
rect 5751 1110 5799 1142
rect 5671 1074 5799 1110
rect 5671 1042 5719 1074
rect 5751 1042 5799 1074
rect 5671 1006 5799 1042
rect 5671 974 5719 1006
rect 5751 974 5799 1006
rect 5671 938 5799 974
rect 5671 906 5719 938
rect 5751 906 5799 938
rect 5671 870 5799 906
rect 5671 838 5719 870
rect 5751 838 5799 870
rect 5671 802 5799 838
rect 5671 770 5719 802
rect 5751 770 5799 802
rect 5671 734 5799 770
rect 5671 702 5719 734
rect 5751 702 5799 734
rect 5671 666 5799 702
rect 5671 634 5719 666
rect 5751 634 5799 666
rect 5671 598 5799 634
rect 5671 566 5719 598
rect 5751 566 5799 598
rect 5671 550 5799 566
rect 5919 1414 6155 1430
rect 5919 1382 6021 1414
rect 6053 1382 6155 1414
rect 5919 1346 6155 1382
rect 5919 1314 6021 1346
rect 6053 1314 6155 1346
rect 5919 1278 6155 1314
rect 5919 1246 6021 1278
rect 6053 1246 6155 1278
rect 5919 1210 6155 1246
rect 5919 1178 6021 1210
rect 6053 1178 6155 1210
rect 5919 1142 6155 1178
rect 5919 1110 6021 1142
rect 6053 1110 6155 1142
rect 5919 1074 6155 1110
rect 5919 1042 6021 1074
rect 6053 1042 6155 1074
rect 5919 1006 6155 1042
rect 5919 974 6021 1006
rect 6053 974 6155 1006
rect 5919 938 6155 974
rect 5919 906 6021 938
rect 6053 906 6155 938
rect 5919 870 6155 906
rect 5919 838 6021 870
rect 6053 838 6155 870
rect 5919 802 6155 838
rect 5919 770 6021 802
rect 6053 770 6155 802
rect 5919 734 6155 770
rect 5919 702 6021 734
rect 6053 702 6155 734
rect 5919 666 6155 702
rect 5919 634 6021 666
rect 6053 634 6155 666
rect 5919 598 6155 634
rect 5919 566 6021 598
rect 6053 566 6155 598
rect 5919 550 6155 566
rect 6275 1414 6403 1430
rect 6275 1382 6323 1414
rect 6355 1382 6403 1414
rect 6275 1346 6403 1382
rect 6275 1314 6323 1346
rect 6355 1314 6403 1346
rect 6275 1278 6403 1314
rect 6275 1246 6323 1278
rect 6355 1246 6403 1278
rect 6275 1210 6403 1246
rect 6275 1178 6323 1210
rect 6355 1178 6403 1210
rect 6275 1142 6403 1178
rect 6275 1110 6323 1142
rect 6355 1110 6403 1142
rect 6275 1074 6403 1110
rect 6275 1042 6323 1074
rect 6355 1042 6403 1074
rect 6275 1006 6403 1042
rect 6275 974 6323 1006
rect 6355 974 6403 1006
rect 6275 938 6403 974
rect 6275 906 6323 938
rect 6355 906 6403 938
rect 6275 870 6403 906
rect 6275 838 6323 870
rect 6355 838 6403 870
rect 6275 802 6403 838
rect 6275 770 6323 802
rect 6355 770 6403 802
rect 6275 734 6403 770
rect 6275 702 6323 734
rect 6355 702 6403 734
rect 6275 666 6403 702
rect 6275 634 6323 666
rect 6355 634 6403 666
rect 6275 598 6403 634
rect 6275 566 6323 598
rect 6355 566 6403 598
rect 6275 550 6403 566
rect 6523 1414 6759 1430
rect 6523 1382 6625 1414
rect 6657 1382 6759 1414
rect 6523 1346 6759 1382
rect 6523 1314 6625 1346
rect 6657 1314 6759 1346
rect 6523 1278 6759 1314
rect 6523 1246 6625 1278
rect 6657 1246 6759 1278
rect 6523 1210 6759 1246
rect 6523 1178 6625 1210
rect 6657 1178 6759 1210
rect 6523 1142 6759 1178
rect 6523 1110 6625 1142
rect 6657 1110 6759 1142
rect 6523 1074 6759 1110
rect 6523 1042 6625 1074
rect 6657 1042 6759 1074
rect 6523 1006 6759 1042
rect 6523 974 6625 1006
rect 6657 974 6759 1006
rect 6523 938 6759 974
rect 6523 906 6625 938
rect 6657 906 6759 938
rect 6523 870 6759 906
rect 6523 838 6625 870
rect 6657 838 6759 870
rect 6523 802 6759 838
rect 6523 770 6625 802
rect 6657 770 6759 802
rect 6523 734 6759 770
rect 6523 702 6625 734
rect 6657 702 6759 734
rect 6523 666 6759 702
rect 6523 634 6625 666
rect 6657 634 6759 666
rect 6523 598 6759 634
rect 6523 566 6625 598
rect 6657 566 6759 598
rect 6523 550 6759 566
rect 6879 1414 7007 1430
rect 6879 1382 6927 1414
rect 6959 1382 7007 1414
rect 6879 1346 7007 1382
rect 6879 1314 6927 1346
rect 6959 1314 7007 1346
rect 6879 1278 7007 1314
rect 6879 1246 6927 1278
rect 6959 1246 7007 1278
rect 6879 1210 7007 1246
rect 6879 1178 6927 1210
rect 6959 1178 7007 1210
rect 6879 1142 7007 1178
rect 6879 1110 6927 1142
rect 6959 1110 7007 1142
rect 6879 1074 7007 1110
rect 6879 1042 6927 1074
rect 6959 1042 7007 1074
rect 6879 1006 7007 1042
rect 6879 974 6927 1006
rect 6959 974 7007 1006
rect 6879 938 7007 974
rect 6879 906 6927 938
rect 6959 906 7007 938
rect 6879 870 7007 906
rect 6879 838 6927 870
rect 6959 838 7007 870
rect 6879 802 7007 838
rect 6879 770 6927 802
rect 6959 770 7007 802
rect 6879 734 7007 770
rect 6879 702 6927 734
rect 6959 702 7007 734
rect 6879 666 7007 702
rect 6879 634 6927 666
rect 6959 634 7007 666
rect 6879 598 7007 634
rect 6879 566 6927 598
rect 6959 566 7007 598
rect 6879 550 7007 566
rect 7127 1414 7363 1430
rect 7127 1382 7229 1414
rect 7261 1382 7363 1414
rect 7127 1346 7363 1382
rect 7127 1314 7229 1346
rect 7261 1314 7363 1346
rect 7127 1278 7363 1314
rect 7127 1246 7229 1278
rect 7261 1246 7363 1278
rect 7127 1210 7363 1246
rect 7127 1178 7229 1210
rect 7261 1178 7363 1210
rect 7127 1142 7363 1178
rect 7127 1110 7229 1142
rect 7261 1110 7363 1142
rect 7127 1074 7363 1110
rect 7127 1042 7229 1074
rect 7261 1042 7363 1074
rect 7127 1006 7363 1042
rect 7127 974 7229 1006
rect 7261 974 7363 1006
rect 7127 938 7363 974
rect 7127 906 7229 938
rect 7261 906 7363 938
rect 7127 870 7363 906
rect 7127 838 7229 870
rect 7261 838 7363 870
rect 7127 802 7363 838
rect 7127 770 7229 802
rect 7261 770 7363 802
rect 7127 734 7363 770
rect 7127 702 7229 734
rect 7261 702 7363 734
rect 7127 666 7363 702
rect 7127 634 7229 666
rect 7261 634 7363 666
rect 7127 598 7363 634
rect 7127 566 7229 598
rect 7261 566 7363 598
rect 7127 550 7363 566
rect 7483 1414 7611 1430
rect 7483 1382 7531 1414
rect 7563 1382 7611 1414
rect 7483 1346 7611 1382
rect 7483 1314 7531 1346
rect 7563 1314 7611 1346
rect 7483 1278 7611 1314
rect 7483 1246 7531 1278
rect 7563 1246 7611 1278
rect 7483 1210 7611 1246
rect 7483 1178 7531 1210
rect 7563 1178 7611 1210
rect 7483 1142 7611 1178
rect 7483 1110 7531 1142
rect 7563 1110 7611 1142
rect 7483 1074 7611 1110
rect 7483 1042 7531 1074
rect 7563 1042 7611 1074
rect 7483 1006 7611 1042
rect 7483 974 7531 1006
rect 7563 974 7611 1006
rect 7483 938 7611 974
rect 7483 906 7531 938
rect 7563 906 7611 938
rect 7483 870 7611 906
rect 7483 838 7531 870
rect 7563 838 7611 870
rect 7483 802 7611 838
rect 7483 770 7531 802
rect 7563 770 7611 802
rect 7483 734 7611 770
rect 7483 702 7531 734
rect 7563 702 7611 734
rect 7483 666 7611 702
rect 7483 634 7531 666
rect 7563 634 7611 666
rect 7483 598 7611 634
rect 7483 566 7531 598
rect 7563 566 7611 598
rect 7483 550 7611 566
rect 7731 1414 7967 1430
rect 7731 1382 7833 1414
rect 7865 1382 7967 1414
rect 7731 1346 7967 1382
rect 7731 1314 7833 1346
rect 7865 1314 7967 1346
rect 7731 1278 7967 1314
rect 7731 1246 7833 1278
rect 7865 1246 7967 1278
rect 7731 1210 7967 1246
rect 7731 1178 7833 1210
rect 7865 1178 7967 1210
rect 7731 1142 7967 1178
rect 7731 1110 7833 1142
rect 7865 1110 7967 1142
rect 7731 1074 7967 1110
rect 7731 1042 7833 1074
rect 7865 1042 7967 1074
rect 7731 1006 7967 1042
rect 7731 974 7833 1006
rect 7865 974 7967 1006
rect 7731 938 7967 974
rect 7731 906 7833 938
rect 7865 906 7967 938
rect 7731 870 7967 906
rect 7731 838 7833 870
rect 7865 838 7967 870
rect 7731 802 7967 838
rect 7731 770 7833 802
rect 7865 770 7967 802
rect 7731 734 7967 770
rect 7731 702 7833 734
rect 7865 702 7967 734
rect 7731 666 7967 702
rect 7731 634 7833 666
rect 7865 634 7967 666
rect 7731 598 7967 634
rect 7731 566 7833 598
rect 7865 566 7967 598
rect 7731 550 7967 566
rect 8087 1414 8215 1430
rect 8087 1382 8135 1414
rect 8167 1382 8215 1414
rect 8087 1346 8215 1382
rect 8087 1314 8135 1346
rect 8167 1314 8215 1346
rect 8087 1278 8215 1314
rect 8087 1246 8135 1278
rect 8167 1246 8215 1278
rect 8087 1210 8215 1246
rect 8087 1178 8135 1210
rect 8167 1178 8215 1210
rect 8087 1142 8215 1178
rect 8087 1110 8135 1142
rect 8167 1110 8215 1142
rect 8087 1074 8215 1110
rect 8087 1042 8135 1074
rect 8167 1042 8215 1074
rect 8087 1006 8215 1042
rect 8087 974 8135 1006
rect 8167 974 8215 1006
rect 8087 938 8215 974
rect 8087 906 8135 938
rect 8167 906 8215 938
rect 8087 870 8215 906
rect 8087 838 8135 870
rect 8167 838 8215 870
rect 8087 802 8215 838
rect 8087 770 8135 802
rect 8167 770 8215 802
rect 8087 734 8215 770
rect 8087 702 8135 734
rect 8167 702 8215 734
rect 8087 666 8215 702
rect 8087 634 8135 666
rect 8167 634 8215 666
rect 8087 598 8215 634
rect 8087 566 8135 598
rect 8167 566 8215 598
rect 8087 550 8215 566
rect 8335 1414 8571 1430
rect 8335 1382 8437 1414
rect 8469 1382 8571 1414
rect 8335 1346 8571 1382
rect 8335 1314 8437 1346
rect 8469 1314 8571 1346
rect 8335 1278 8571 1314
rect 8335 1246 8437 1278
rect 8469 1246 8571 1278
rect 8335 1210 8571 1246
rect 8335 1178 8437 1210
rect 8469 1178 8571 1210
rect 8335 1142 8571 1178
rect 8335 1110 8437 1142
rect 8469 1110 8571 1142
rect 8335 1074 8571 1110
rect 8335 1042 8437 1074
rect 8469 1042 8571 1074
rect 8335 1006 8571 1042
rect 8335 974 8437 1006
rect 8469 974 8571 1006
rect 8335 938 8571 974
rect 8335 906 8437 938
rect 8469 906 8571 938
rect 8335 870 8571 906
rect 8335 838 8437 870
rect 8469 838 8571 870
rect 8335 802 8571 838
rect 8335 770 8437 802
rect 8469 770 8571 802
rect 8335 734 8571 770
rect 8335 702 8437 734
rect 8469 702 8571 734
rect 8335 666 8571 702
rect 8335 634 8437 666
rect 8469 634 8571 666
rect 8335 598 8571 634
rect 8335 566 8437 598
rect 8469 566 8571 598
rect 8335 550 8571 566
rect 8691 1414 8819 1430
rect 8691 1382 8739 1414
rect 8771 1382 8819 1414
rect 8691 1346 8819 1382
rect 8691 1314 8739 1346
rect 8771 1314 8819 1346
rect 8691 1278 8819 1314
rect 8691 1246 8739 1278
rect 8771 1246 8819 1278
rect 8691 1210 8819 1246
rect 8691 1178 8739 1210
rect 8771 1178 8819 1210
rect 8691 1142 8819 1178
rect 8691 1110 8739 1142
rect 8771 1110 8819 1142
rect 8691 1074 8819 1110
rect 8691 1042 8739 1074
rect 8771 1042 8819 1074
rect 8691 1006 8819 1042
rect 8691 974 8739 1006
rect 8771 974 8819 1006
rect 8691 938 8819 974
rect 8691 906 8739 938
rect 8771 906 8819 938
rect 8691 870 8819 906
rect 8691 838 8739 870
rect 8771 838 8819 870
rect 8691 802 8819 838
rect 8691 770 8739 802
rect 8771 770 8819 802
rect 8691 734 8819 770
rect 8691 702 8739 734
rect 8771 702 8819 734
rect 8691 666 8819 702
rect 8691 634 8739 666
rect 8771 634 8819 666
rect 8691 598 8819 634
rect 8691 566 8739 598
rect 8771 566 8819 598
rect 8691 550 8819 566
rect 8939 1414 9175 1430
rect 8939 1382 9041 1414
rect 9073 1382 9175 1414
rect 8939 1346 9175 1382
rect 8939 1314 9041 1346
rect 9073 1314 9175 1346
rect 8939 1278 9175 1314
rect 8939 1246 9041 1278
rect 9073 1246 9175 1278
rect 8939 1210 9175 1246
rect 8939 1178 9041 1210
rect 9073 1178 9175 1210
rect 8939 1142 9175 1178
rect 8939 1110 9041 1142
rect 9073 1110 9175 1142
rect 8939 1074 9175 1110
rect 8939 1042 9041 1074
rect 9073 1042 9175 1074
rect 8939 1006 9175 1042
rect 8939 974 9041 1006
rect 9073 974 9175 1006
rect 8939 938 9175 974
rect 8939 906 9041 938
rect 9073 906 9175 938
rect 8939 870 9175 906
rect 8939 838 9041 870
rect 9073 838 9175 870
rect 8939 802 9175 838
rect 8939 770 9041 802
rect 9073 770 9175 802
rect 8939 734 9175 770
rect 8939 702 9041 734
rect 9073 702 9175 734
rect 8939 666 9175 702
rect 8939 634 9041 666
rect 9073 634 9175 666
rect 8939 598 9175 634
rect 8939 566 9041 598
rect 9073 566 9175 598
rect 8939 550 9175 566
rect 9295 1414 9423 1430
rect 9295 1382 9343 1414
rect 9375 1382 9423 1414
rect 9295 1346 9423 1382
rect 9295 1314 9343 1346
rect 9375 1314 9423 1346
rect 9295 1278 9423 1314
rect 9295 1246 9343 1278
rect 9375 1246 9423 1278
rect 9295 1210 9423 1246
rect 9295 1178 9343 1210
rect 9375 1178 9423 1210
rect 9295 1142 9423 1178
rect 9295 1110 9343 1142
rect 9375 1110 9423 1142
rect 9295 1074 9423 1110
rect 9295 1042 9343 1074
rect 9375 1042 9423 1074
rect 9295 1006 9423 1042
rect 9295 974 9343 1006
rect 9375 974 9423 1006
rect 9295 938 9423 974
rect 9295 906 9343 938
rect 9375 906 9423 938
rect 9295 870 9423 906
rect 9295 838 9343 870
rect 9375 838 9423 870
rect 9295 802 9423 838
rect 9295 770 9343 802
rect 9375 770 9423 802
rect 9295 734 9423 770
rect 9295 702 9343 734
rect 9375 702 9423 734
rect 9295 666 9423 702
rect 9295 634 9343 666
rect 9375 634 9423 666
rect 9295 598 9423 634
rect 9295 566 9343 598
rect 9375 566 9423 598
rect 9295 550 9423 566
rect 9543 1414 9779 1430
rect 9543 1382 9645 1414
rect 9677 1382 9779 1414
rect 9543 1346 9779 1382
rect 9543 1314 9645 1346
rect 9677 1314 9779 1346
rect 9543 1278 9779 1314
rect 9543 1246 9645 1278
rect 9677 1246 9779 1278
rect 9543 1210 9779 1246
rect 9543 1178 9645 1210
rect 9677 1178 9779 1210
rect 9543 1142 9779 1178
rect 9543 1110 9645 1142
rect 9677 1110 9779 1142
rect 9543 1074 9779 1110
rect 9543 1042 9645 1074
rect 9677 1042 9779 1074
rect 9543 1006 9779 1042
rect 9543 974 9645 1006
rect 9677 974 9779 1006
rect 9543 938 9779 974
rect 9543 906 9645 938
rect 9677 906 9779 938
rect 9543 870 9779 906
rect 9543 838 9645 870
rect 9677 838 9779 870
rect 9543 802 9779 838
rect 9543 770 9645 802
rect 9677 770 9779 802
rect 9543 734 9779 770
rect 9543 702 9645 734
rect 9677 702 9779 734
rect 9543 666 9779 702
rect 9543 634 9645 666
rect 9677 634 9779 666
rect 9543 598 9779 634
rect 9543 566 9645 598
rect 9677 566 9779 598
rect 9543 550 9779 566
rect 9899 1414 10027 1430
rect 9899 1382 9947 1414
rect 9979 1382 10027 1414
rect 9899 1346 10027 1382
rect 9899 1314 9947 1346
rect 9979 1314 10027 1346
rect 9899 1278 10027 1314
rect 9899 1246 9947 1278
rect 9979 1246 10027 1278
rect 9899 1210 10027 1246
rect 9899 1178 9947 1210
rect 9979 1178 10027 1210
rect 9899 1142 10027 1178
rect 9899 1110 9947 1142
rect 9979 1110 10027 1142
rect 9899 1074 10027 1110
rect 9899 1042 9947 1074
rect 9979 1042 10027 1074
rect 9899 1006 10027 1042
rect 9899 974 9947 1006
rect 9979 974 10027 1006
rect 9899 938 10027 974
rect 9899 906 9947 938
rect 9979 906 10027 938
rect 9899 870 10027 906
rect 9899 838 9947 870
rect 9979 838 10027 870
rect 9899 802 10027 838
rect 9899 770 9947 802
rect 9979 770 10027 802
rect 9899 734 10027 770
rect 9899 702 9947 734
rect 9979 702 10027 734
rect 9899 666 10027 702
rect 9899 634 9947 666
rect 9979 634 10027 666
rect 9899 598 10027 634
rect 9899 566 9947 598
rect 9979 566 10027 598
rect 9899 550 10027 566
rect 10147 1414 10383 1430
rect 10147 1382 10249 1414
rect 10281 1382 10383 1414
rect 10147 1346 10383 1382
rect 10147 1314 10249 1346
rect 10281 1314 10383 1346
rect 10147 1278 10383 1314
rect 10147 1246 10249 1278
rect 10281 1246 10383 1278
rect 10147 1210 10383 1246
rect 10147 1178 10249 1210
rect 10281 1178 10383 1210
rect 10147 1142 10383 1178
rect 10147 1110 10249 1142
rect 10281 1110 10383 1142
rect 10147 1074 10383 1110
rect 10147 1042 10249 1074
rect 10281 1042 10383 1074
rect 10147 1006 10383 1042
rect 10147 974 10249 1006
rect 10281 974 10383 1006
rect 10147 938 10383 974
rect 10147 906 10249 938
rect 10281 906 10383 938
rect 10147 870 10383 906
rect 10147 838 10249 870
rect 10281 838 10383 870
rect 10147 802 10383 838
rect 10147 770 10249 802
rect 10281 770 10383 802
rect 10147 734 10383 770
rect 10147 702 10249 734
rect 10281 702 10383 734
rect 10147 666 10383 702
rect 10147 634 10249 666
rect 10281 634 10383 666
rect 10147 598 10383 634
rect 10147 566 10249 598
rect 10281 566 10383 598
rect 10147 550 10383 566
rect 10503 1414 10631 1430
rect 10503 1382 10551 1414
rect 10583 1382 10631 1414
rect 10503 1346 10631 1382
rect 10503 1314 10551 1346
rect 10583 1314 10631 1346
rect 10503 1278 10631 1314
rect 10503 1246 10551 1278
rect 10583 1246 10631 1278
rect 10503 1210 10631 1246
rect 10503 1178 10551 1210
rect 10583 1178 10631 1210
rect 10503 1142 10631 1178
rect 10503 1110 10551 1142
rect 10583 1110 10631 1142
rect 10503 1074 10631 1110
rect 10503 1042 10551 1074
rect 10583 1042 10631 1074
rect 10503 1006 10631 1042
rect 10503 974 10551 1006
rect 10583 974 10631 1006
rect 10503 938 10631 974
rect 10503 906 10551 938
rect 10583 906 10631 938
rect 10503 870 10631 906
rect 10503 838 10551 870
rect 10583 838 10631 870
rect 10503 802 10631 838
rect 10503 770 10551 802
rect 10583 770 10631 802
rect 10503 734 10631 770
rect 10503 702 10551 734
rect 10583 702 10631 734
rect 10503 666 10631 702
rect 10503 634 10551 666
rect 10583 634 10631 666
rect 10503 598 10631 634
rect 10503 566 10551 598
rect 10583 566 10631 598
rect 10503 550 10631 566
rect 10751 1414 10987 1430
rect 10751 1382 10853 1414
rect 10885 1382 10987 1414
rect 10751 1346 10987 1382
rect 10751 1314 10853 1346
rect 10885 1314 10987 1346
rect 10751 1278 10987 1314
rect 10751 1246 10853 1278
rect 10885 1246 10987 1278
rect 10751 1210 10987 1246
rect 10751 1178 10853 1210
rect 10885 1178 10987 1210
rect 10751 1142 10987 1178
rect 10751 1110 10853 1142
rect 10885 1110 10987 1142
rect 10751 1074 10987 1110
rect 10751 1042 10853 1074
rect 10885 1042 10987 1074
rect 10751 1006 10987 1042
rect 10751 974 10853 1006
rect 10885 974 10987 1006
rect 10751 938 10987 974
rect 10751 906 10853 938
rect 10885 906 10987 938
rect 10751 870 10987 906
rect 10751 838 10853 870
rect 10885 838 10987 870
rect 10751 802 10987 838
rect 10751 770 10853 802
rect 10885 770 10987 802
rect 10751 734 10987 770
rect 10751 702 10853 734
rect 10885 702 10987 734
rect 10751 666 10987 702
rect 10751 634 10853 666
rect 10885 634 10987 666
rect 10751 598 10987 634
rect 10751 566 10853 598
rect 10885 566 10987 598
rect 10751 550 10987 566
rect 11107 1414 11235 1430
rect 11107 1382 11155 1414
rect 11187 1382 11235 1414
rect 11107 1346 11235 1382
rect 11107 1314 11155 1346
rect 11187 1314 11235 1346
rect 11107 1278 11235 1314
rect 11107 1246 11155 1278
rect 11187 1246 11235 1278
rect 11107 1210 11235 1246
rect 11107 1178 11155 1210
rect 11187 1178 11235 1210
rect 11107 1142 11235 1178
rect 11107 1110 11155 1142
rect 11187 1110 11235 1142
rect 11107 1074 11235 1110
rect 11107 1042 11155 1074
rect 11187 1042 11235 1074
rect 11107 1006 11235 1042
rect 11107 974 11155 1006
rect 11187 974 11235 1006
rect 11107 938 11235 974
rect 11107 906 11155 938
rect 11187 906 11235 938
rect 11107 870 11235 906
rect 11107 838 11155 870
rect 11187 838 11235 870
rect 11107 802 11235 838
rect 11107 770 11155 802
rect 11187 770 11235 802
rect 11107 734 11235 770
rect 11107 702 11155 734
rect 11187 702 11235 734
rect 11107 666 11235 702
rect 11107 634 11155 666
rect 11187 634 11235 666
rect 11107 598 11235 634
rect 11107 566 11155 598
rect 11187 566 11235 598
rect 11107 550 11235 566
rect 11355 1414 11591 1430
rect 11355 1382 11457 1414
rect 11489 1382 11591 1414
rect 11355 1346 11591 1382
rect 11355 1314 11457 1346
rect 11489 1314 11591 1346
rect 11355 1278 11591 1314
rect 11355 1246 11457 1278
rect 11489 1246 11591 1278
rect 11355 1210 11591 1246
rect 11355 1178 11457 1210
rect 11489 1178 11591 1210
rect 11355 1142 11591 1178
rect 11355 1110 11457 1142
rect 11489 1110 11591 1142
rect 11355 1074 11591 1110
rect 11355 1042 11457 1074
rect 11489 1042 11591 1074
rect 11355 1006 11591 1042
rect 11355 974 11457 1006
rect 11489 974 11591 1006
rect 11355 938 11591 974
rect 11355 906 11457 938
rect 11489 906 11591 938
rect 11355 870 11591 906
rect 11355 838 11457 870
rect 11489 838 11591 870
rect 11355 802 11591 838
rect 11355 770 11457 802
rect 11489 770 11591 802
rect 11355 734 11591 770
rect 11355 702 11457 734
rect 11489 702 11591 734
rect 11355 666 11591 702
rect 11355 634 11457 666
rect 11489 634 11591 666
rect 11355 598 11591 634
rect 11355 566 11457 598
rect 11489 566 11591 598
rect 11355 550 11591 566
rect 11711 1414 11839 1430
rect 11711 1382 11759 1414
rect 11791 1382 11839 1414
rect 11711 1346 11839 1382
rect 11711 1314 11759 1346
rect 11791 1314 11839 1346
rect 11711 1278 11839 1314
rect 11711 1246 11759 1278
rect 11791 1246 11839 1278
rect 11711 1210 11839 1246
rect 11711 1178 11759 1210
rect 11791 1178 11839 1210
rect 11711 1142 11839 1178
rect 11711 1110 11759 1142
rect 11791 1110 11839 1142
rect 11711 1074 11839 1110
rect 11711 1042 11759 1074
rect 11791 1042 11839 1074
rect 11711 1006 11839 1042
rect 11711 974 11759 1006
rect 11791 974 11839 1006
rect 11711 938 11839 974
rect 11711 906 11759 938
rect 11791 906 11839 938
rect 11711 870 11839 906
rect 11711 838 11759 870
rect 11791 838 11839 870
rect 11711 802 11839 838
rect 11711 770 11759 802
rect 11791 770 11839 802
rect 11711 734 11839 770
rect 11711 702 11759 734
rect 11791 702 11839 734
rect 11711 666 11839 702
rect 11711 634 11759 666
rect 11791 634 11839 666
rect 11711 598 11839 634
rect 11711 566 11759 598
rect 11791 566 11839 598
rect 11711 550 11839 566
rect 11959 1414 12195 1430
rect 11959 1382 12061 1414
rect 12093 1382 12195 1414
rect 11959 1346 12195 1382
rect 11959 1314 12061 1346
rect 12093 1314 12195 1346
rect 11959 1278 12195 1314
rect 11959 1246 12061 1278
rect 12093 1246 12195 1278
rect 11959 1210 12195 1246
rect 11959 1178 12061 1210
rect 12093 1178 12195 1210
rect 11959 1142 12195 1178
rect 11959 1110 12061 1142
rect 12093 1110 12195 1142
rect 11959 1074 12195 1110
rect 11959 1042 12061 1074
rect 12093 1042 12195 1074
rect 11959 1006 12195 1042
rect 11959 974 12061 1006
rect 12093 974 12195 1006
rect 11959 938 12195 974
rect 11959 906 12061 938
rect 12093 906 12195 938
rect 11959 870 12195 906
rect 11959 838 12061 870
rect 12093 838 12195 870
rect 11959 802 12195 838
rect 11959 770 12061 802
rect 12093 770 12195 802
rect 11959 734 12195 770
rect 11959 702 12061 734
rect 12093 702 12195 734
rect 11959 666 12195 702
rect 11959 634 12061 666
rect 12093 634 12195 666
rect 11959 598 12195 634
rect 11959 566 12061 598
rect 12093 566 12195 598
rect 11959 550 12195 566
rect 12315 1414 12443 1430
rect 12315 1382 12363 1414
rect 12395 1382 12443 1414
rect 12315 1346 12443 1382
rect 12315 1314 12363 1346
rect 12395 1314 12443 1346
rect 12315 1278 12443 1314
rect 12315 1246 12363 1278
rect 12395 1246 12443 1278
rect 12315 1210 12443 1246
rect 12315 1178 12363 1210
rect 12395 1178 12443 1210
rect 12315 1142 12443 1178
rect 12315 1110 12363 1142
rect 12395 1110 12443 1142
rect 12315 1074 12443 1110
rect 12315 1042 12363 1074
rect 12395 1042 12443 1074
rect 12315 1006 12443 1042
rect 12315 974 12363 1006
rect 12395 974 12443 1006
rect 12315 938 12443 974
rect 12315 906 12363 938
rect 12395 906 12443 938
rect 12315 870 12443 906
rect 12315 838 12363 870
rect 12395 838 12443 870
rect 12315 802 12443 838
rect 12315 770 12363 802
rect 12395 770 12443 802
rect 12315 734 12443 770
rect 12315 702 12363 734
rect 12395 702 12443 734
rect 12315 666 12443 702
rect 12315 634 12363 666
rect 12395 634 12443 666
rect 12315 598 12443 634
rect 12315 566 12363 598
rect 12395 566 12443 598
rect 12315 550 12443 566
rect 12563 1414 12799 1430
rect 12563 1382 12665 1414
rect 12697 1382 12799 1414
rect 12563 1346 12799 1382
rect 12563 1314 12665 1346
rect 12697 1314 12799 1346
rect 12563 1278 12799 1314
rect 12563 1246 12665 1278
rect 12697 1246 12799 1278
rect 12563 1210 12799 1246
rect 12563 1178 12665 1210
rect 12697 1178 12799 1210
rect 12563 1142 12799 1178
rect 12563 1110 12665 1142
rect 12697 1110 12799 1142
rect 12563 1074 12799 1110
rect 12563 1042 12665 1074
rect 12697 1042 12799 1074
rect 12563 1006 12799 1042
rect 12563 974 12665 1006
rect 12697 974 12799 1006
rect 12563 938 12799 974
rect 12563 906 12665 938
rect 12697 906 12799 938
rect 12563 870 12799 906
rect 12563 838 12665 870
rect 12697 838 12799 870
rect 12563 802 12799 838
rect 12563 770 12665 802
rect 12697 770 12799 802
rect 12563 734 12799 770
rect 12563 702 12665 734
rect 12697 702 12799 734
rect 12563 666 12799 702
rect 12563 634 12665 666
rect 12697 634 12799 666
rect 12563 598 12799 634
rect 12563 566 12665 598
rect 12697 566 12799 598
rect 12563 550 12799 566
rect 12919 1414 13047 1430
rect 12919 1382 12967 1414
rect 12999 1382 13047 1414
rect 12919 1346 13047 1382
rect 12919 1314 12967 1346
rect 12999 1314 13047 1346
rect 12919 1278 13047 1314
rect 12919 1246 12967 1278
rect 12999 1246 13047 1278
rect 12919 1210 13047 1246
rect 12919 1178 12967 1210
rect 12999 1178 13047 1210
rect 12919 1142 13047 1178
rect 12919 1110 12967 1142
rect 12999 1110 13047 1142
rect 12919 1074 13047 1110
rect 12919 1042 12967 1074
rect 12999 1042 13047 1074
rect 12919 1006 13047 1042
rect 12919 974 12967 1006
rect 12999 974 13047 1006
rect 12919 938 13047 974
rect 12919 906 12967 938
rect 12999 906 13047 938
rect 12919 870 13047 906
rect 12919 838 12967 870
rect 12999 838 13047 870
rect 12919 802 13047 838
rect 12919 770 12967 802
rect 12999 770 13047 802
rect 12919 734 13047 770
rect 12919 702 12967 734
rect 12999 702 13047 734
rect 12919 666 13047 702
rect 12919 634 12967 666
rect 12999 634 13047 666
rect 12919 598 13047 634
rect 12919 566 12967 598
rect 12999 566 13047 598
rect 12919 550 13047 566
rect 13167 1414 13403 1430
rect 13167 1382 13269 1414
rect 13301 1382 13403 1414
rect 13167 1346 13403 1382
rect 13167 1314 13269 1346
rect 13301 1314 13403 1346
rect 13167 1278 13403 1314
rect 13167 1246 13269 1278
rect 13301 1246 13403 1278
rect 13167 1210 13403 1246
rect 13167 1178 13269 1210
rect 13301 1178 13403 1210
rect 13167 1142 13403 1178
rect 13167 1110 13269 1142
rect 13301 1110 13403 1142
rect 13167 1074 13403 1110
rect 13167 1042 13269 1074
rect 13301 1042 13403 1074
rect 13167 1006 13403 1042
rect 13167 974 13269 1006
rect 13301 974 13403 1006
rect 13167 938 13403 974
rect 13167 906 13269 938
rect 13301 906 13403 938
rect 13167 870 13403 906
rect 13167 838 13269 870
rect 13301 838 13403 870
rect 13167 802 13403 838
rect 13167 770 13269 802
rect 13301 770 13403 802
rect 13167 734 13403 770
rect 13167 702 13269 734
rect 13301 702 13403 734
rect 13167 666 13403 702
rect 13167 634 13269 666
rect 13301 634 13403 666
rect 13167 598 13403 634
rect 13167 566 13269 598
rect 13301 566 13403 598
rect 13167 550 13403 566
rect 13523 1414 13651 1430
rect 13523 1382 13571 1414
rect 13603 1382 13651 1414
rect 13523 1346 13651 1382
rect 13523 1314 13571 1346
rect 13603 1314 13651 1346
rect 13523 1278 13651 1314
rect 13523 1246 13571 1278
rect 13603 1246 13651 1278
rect 13523 1210 13651 1246
rect 13523 1178 13571 1210
rect 13603 1178 13651 1210
rect 13523 1142 13651 1178
rect 13523 1110 13571 1142
rect 13603 1110 13651 1142
rect 13523 1074 13651 1110
rect 13523 1042 13571 1074
rect 13603 1042 13651 1074
rect 13523 1006 13651 1042
rect 13523 974 13571 1006
rect 13603 974 13651 1006
rect 13523 938 13651 974
rect 13523 906 13571 938
rect 13603 906 13651 938
rect 13523 870 13651 906
rect 13523 838 13571 870
rect 13603 838 13651 870
rect 13523 802 13651 838
rect 13523 770 13571 802
rect 13603 770 13651 802
rect 13523 734 13651 770
rect 13523 702 13571 734
rect 13603 702 13651 734
rect 13523 666 13651 702
rect 13523 634 13571 666
rect 13603 634 13651 666
rect 13523 598 13651 634
rect 13523 566 13571 598
rect 13603 566 13651 598
rect 13523 550 13651 566
rect 13771 1414 14007 1430
rect 13771 1382 13873 1414
rect 13905 1382 14007 1414
rect 13771 1346 14007 1382
rect 13771 1314 13873 1346
rect 13905 1314 14007 1346
rect 13771 1278 14007 1314
rect 13771 1246 13873 1278
rect 13905 1246 14007 1278
rect 13771 1210 14007 1246
rect 13771 1178 13873 1210
rect 13905 1178 14007 1210
rect 13771 1142 14007 1178
rect 13771 1110 13873 1142
rect 13905 1110 14007 1142
rect 13771 1074 14007 1110
rect 13771 1042 13873 1074
rect 13905 1042 14007 1074
rect 13771 1006 14007 1042
rect 13771 974 13873 1006
rect 13905 974 14007 1006
rect 13771 938 14007 974
rect 13771 906 13873 938
rect 13905 906 14007 938
rect 13771 870 14007 906
rect 13771 838 13873 870
rect 13905 838 14007 870
rect 13771 802 14007 838
rect 13771 770 13873 802
rect 13905 770 14007 802
rect 13771 734 14007 770
rect 13771 702 13873 734
rect 13905 702 14007 734
rect 13771 666 14007 702
rect 13771 634 13873 666
rect 13905 634 14007 666
rect 13771 598 14007 634
rect 13771 566 13873 598
rect 13905 566 14007 598
rect 13771 550 14007 566
rect 14127 1414 14255 1430
rect 14127 1382 14175 1414
rect 14207 1382 14255 1414
rect 14127 1346 14255 1382
rect 14127 1314 14175 1346
rect 14207 1314 14255 1346
rect 14127 1278 14255 1314
rect 14127 1246 14175 1278
rect 14207 1246 14255 1278
rect 14127 1210 14255 1246
rect 14127 1178 14175 1210
rect 14207 1178 14255 1210
rect 14127 1142 14255 1178
rect 14127 1110 14175 1142
rect 14207 1110 14255 1142
rect 14127 1074 14255 1110
rect 14127 1042 14175 1074
rect 14207 1042 14255 1074
rect 14127 1006 14255 1042
rect 14127 974 14175 1006
rect 14207 974 14255 1006
rect 14127 938 14255 974
rect 14127 906 14175 938
rect 14207 906 14255 938
rect 14127 870 14255 906
rect 14127 838 14175 870
rect 14207 838 14255 870
rect 14127 802 14255 838
rect 14127 770 14175 802
rect 14207 770 14255 802
rect 14127 734 14255 770
rect 14127 702 14175 734
rect 14207 702 14255 734
rect 14127 666 14255 702
rect 14127 634 14175 666
rect 14207 634 14255 666
rect 14127 598 14255 634
rect 14127 566 14175 598
rect 14207 566 14255 598
rect 14127 550 14255 566
rect 14375 1414 14523 1430
rect 14375 1382 14477 1414
rect 14509 1382 14523 1414
rect 14375 1346 14523 1382
rect 14375 1314 14477 1346
rect 14509 1314 14523 1346
rect 14375 1278 14523 1314
rect 14375 1246 14477 1278
rect 14509 1246 14523 1278
rect 14375 1210 14523 1246
rect 14375 1178 14477 1210
rect 14509 1178 14523 1210
rect 14375 1142 14523 1178
rect 14375 1110 14477 1142
rect 14509 1110 14523 1142
rect 14375 1074 14523 1110
rect 14375 1042 14477 1074
rect 14509 1042 14523 1074
rect 14375 1006 14523 1042
rect 14375 974 14477 1006
rect 14509 974 14523 1006
rect 14375 938 14523 974
rect 14375 906 14477 938
rect 14509 906 14523 938
rect 14375 870 14523 906
rect 14375 838 14477 870
rect 14509 838 14523 870
rect 14375 802 14523 838
rect 14375 770 14477 802
rect 14509 770 14523 802
rect 14375 734 14523 770
rect 14375 702 14477 734
rect 14509 702 14523 734
rect 14375 666 14523 702
rect 14375 634 14477 666
rect 14509 634 14523 666
rect 14375 598 14523 634
rect 14375 566 14477 598
rect 14509 566 14523 598
rect 14375 550 14523 566
<< hvndiffc >>
rect 1491 4286 1523 4318
rect 1491 4218 1523 4250
rect 1491 4150 1523 4182
rect 1491 4082 1523 4114
rect 1491 4014 1523 4046
rect 1491 3946 1523 3978
rect 1491 3878 1523 3910
rect 1491 3810 1523 3842
rect 1491 3742 1523 3774
rect 1491 3674 1523 3706
rect 1491 3606 1523 3638
rect 1491 3538 1523 3570
rect 1491 3470 1523 3502
rect 1793 4286 1825 4318
rect 1793 4218 1825 4250
rect 1793 4150 1825 4182
rect 1793 4082 1825 4114
rect 1793 4014 1825 4046
rect 1793 3946 1825 3978
rect 1793 3878 1825 3910
rect 1793 3810 1825 3842
rect 1793 3742 1825 3774
rect 1793 3674 1825 3706
rect 1793 3606 1825 3638
rect 1793 3538 1825 3570
rect 1793 3470 1825 3502
rect 2095 4286 2127 4318
rect 2095 4218 2127 4250
rect 2095 4150 2127 4182
rect 2095 4082 2127 4114
rect 2095 4014 2127 4046
rect 2095 3946 2127 3978
rect 2095 3878 2127 3910
rect 2095 3810 2127 3842
rect 2095 3742 2127 3774
rect 2095 3674 2127 3706
rect 2095 3606 2127 3638
rect 2095 3538 2127 3570
rect 2095 3470 2127 3502
rect 2397 4286 2429 4318
rect 2397 4218 2429 4250
rect 2397 4150 2429 4182
rect 2397 4082 2429 4114
rect 2397 4014 2429 4046
rect 2397 3946 2429 3978
rect 2397 3878 2429 3910
rect 2397 3810 2429 3842
rect 2397 3742 2429 3774
rect 2397 3674 2429 3706
rect 2397 3606 2429 3638
rect 2397 3538 2429 3570
rect 2397 3470 2429 3502
rect 2699 4286 2731 4318
rect 2699 4218 2731 4250
rect 2699 4150 2731 4182
rect 2699 4082 2731 4114
rect 2699 4014 2731 4046
rect 2699 3946 2731 3978
rect 2699 3878 2731 3910
rect 2699 3810 2731 3842
rect 2699 3742 2731 3774
rect 2699 3674 2731 3706
rect 2699 3606 2731 3638
rect 2699 3538 2731 3570
rect 2699 3470 2731 3502
rect 3001 4286 3033 4318
rect 3001 4218 3033 4250
rect 3001 4150 3033 4182
rect 3001 4082 3033 4114
rect 3001 4014 3033 4046
rect 3001 3946 3033 3978
rect 3001 3878 3033 3910
rect 3001 3810 3033 3842
rect 3001 3742 3033 3774
rect 3001 3674 3033 3706
rect 3001 3606 3033 3638
rect 3001 3538 3033 3570
rect 3001 3470 3033 3502
rect 3303 4286 3335 4318
rect 3303 4218 3335 4250
rect 3303 4150 3335 4182
rect 3303 4082 3335 4114
rect 3303 4014 3335 4046
rect 3303 3946 3335 3978
rect 3303 3878 3335 3910
rect 3303 3810 3335 3842
rect 3303 3742 3335 3774
rect 3303 3674 3335 3706
rect 3303 3606 3335 3638
rect 3303 3538 3335 3570
rect 3303 3470 3335 3502
rect 3605 4286 3637 4318
rect 3605 4218 3637 4250
rect 3605 4150 3637 4182
rect 3605 4082 3637 4114
rect 3605 4014 3637 4046
rect 3605 3946 3637 3978
rect 3605 3878 3637 3910
rect 3605 3810 3637 3842
rect 3605 3742 3637 3774
rect 3605 3674 3637 3706
rect 3605 3606 3637 3638
rect 3605 3538 3637 3570
rect 3605 3470 3637 3502
rect 3907 4286 3939 4318
rect 3907 4218 3939 4250
rect 3907 4150 3939 4182
rect 3907 4082 3939 4114
rect 3907 4014 3939 4046
rect 3907 3946 3939 3978
rect 3907 3878 3939 3910
rect 3907 3810 3939 3842
rect 3907 3742 3939 3774
rect 3907 3674 3939 3706
rect 3907 3606 3939 3638
rect 3907 3538 3939 3570
rect 3907 3470 3939 3502
rect 4209 4286 4241 4318
rect 4209 4218 4241 4250
rect 4209 4150 4241 4182
rect 4209 4082 4241 4114
rect 4209 4014 4241 4046
rect 4209 3946 4241 3978
rect 4209 3878 4241 3910
rect 4209 3810 4241 3842
rect 4209 3742 4241 3774
rect 4209 3674 4241 3706
rect 4209 3606 4241 3638
rect 4209 3538 4241 3570
rect 4209 3470 4241 3502
rect 4511 4286 4543 4318
rect 4511 4218 4543 4250
rect 4511 4150 4543 4182
rect 4511 4082 4543 4114
rect 4511 4014 4543 4046
rect 4511 3946 4543 3978
rect 4511 3878 4543 3910
rect 4511 3810 4543 3842
rect 4511 3742 4543 3774
rect 4511 3674 4543 3706
rect 4511 3606 4543 3638
rect 4511 3538 4543 3570
rect 4511 3470 4543 3502
rect 4813 4286 4845 4318
rect 4813 4218 4845 4250
rect 4813 4150 4845 4182
rect 4813 4082 4845 4114
rect 4813 4014 4845 4046
rect 4813 3946 4845 3978
rect 4813 3878 4845 3910
rect 4813 3810 4845 3842
rect 4813 3742 4845 3774
rect 4813 3674 4845 3706
rect 4813 3606 4845 3638
rect 4813 3538 4845 3570
rect 4813 3470 4845 3502
rect 5115 4286 5147 4318
rect 5115 4218 5147 4250
rect 5115 4150 5147 4182
rect 5115 4082 5147 4114
rect 5115 4014 5147 4046
rect 5115 3946 5147 3978
rect 5115 3878 5147 3910
rect 5115 3810 5147 3842
rect 5115 3742 5147 3774
rect 5115 3674 5147 3706
rect 5115 3606 5147 3638
rect 5115 3538 5147 3570
rect 5115 3470 5147 3502
rect 5417 4286 5449 4318
rect 5417 4218 5449 4250
rect 5417 4150 5449 4182
rect 5417 4082 5449 4114
rect 5417 4014 5449 4046
rect 5417 3946 5449 3978
rect 5417 3878 5449 3910
rect 5417 3810 5449 3842
rect 5417 3742 5449 3774
rect 5417 3674 5449 3706
rect 5417 3606 5449 3638
rect 5417 3538 5449 3570
rect 5417 3470 5449 3502
rect 5719 4286 5751 4318
rect 5719 4218 5751 4250
rect 5719 4150 5751 4182
rect 5719 4082 5751 4114
rect 5719 4014 5751 4046
rect 5719 3946 5751 3978
rect 5719 3878 5751 3910
rect 5719 3810 5751 3842
rect 5719 3742 5751 3774
rect 5719 3674 5751 3706
rect 5719 3606 5751 3638
rect 5719 3538 5751 3570
rect 5719 3470 5751 3502
rect 6021 4286 6053 4318
rect 6021 4218 6053 4250
rect 6021 4150 6053 4182
rect 6021 4082 6053 4114
rect 6021 4014 6053 4046
rect 6021 3946 6053 3978
rect 6021 3878 6053 3910
rect 6021 3810 6053 3842
rect 6021 3742 6053 3774
rect 6021 3674 6053 3706
rect 6021 3606 6053 3638
rect 6021 3538 6053 3570
rect 6021 3470 6053 3502
rect 6323 4286 6355 4318
rect 6323 4218 6355 4250
rect 6323 4150 6355 4182
rect 6323 4082 6355 4114
rect 6323 4014 6355 4046
rect 6323 3946 6355 3978
rect 6323 3878 6355 3910
rect 6323 3810 6355 3842
rect 6323 3742 6355 3774
rect 6323 3674 6355 3706
rect 6323 3606 6355 3638
rect 6323 3538 6355 3570
rect 6323 3470 6355 3502
rect 6625 4286 6657 4318
rect 6625 4218 6657 4250
rect 6625 4150 6657 4182
rect 6625 4082 6657 4114
rect 6625 4014 6657 4046
rect 6625 3946 6657 3978
rect 6625 3878 6657 3910
rect 6625 3810 6657 3842
rect 6625 3742 6657 3774
rect 6625 3674 6657 3706
rect 6625 3606 6657 3638
rect 6625 3538 6657 3570
rect 6625 3470 6657 3502
rect 6927 4286 6959 4318
rect 6927 4218 6959 4250
rect 6927 4150 6959 4182
rect 6927 4082 6959 4114
rect 6927 4014 6959 4046
rect 6927 3946 6959 3978
rect 6927 3878 6959 3910
rect 6927 3810 6959 3842
rect 6927 3742 6959 3774
rect 6927 3674 6959 3706
rect 6927 3606 6959 3638
rect 6927 3538 6959 3570
rect 6927 3470 6959 3502
rect 7229 4286 7261 4318
rect 7229 4218 7261 4250
rect 7229 4150 7261 4182
rect 7229 4082 7261 4114
rect 7229 4014 7261 4046
rect 7229 3946 7261 3978
rect 7229 3878 7261 3910
rect 7229 3810 7261 3842
rect 7229 3742 7261 3774
rect 7229 3674 7261 3706
rect 7229 3606 7261 3638
rect 7229 3538 7261 3570
rect 7229 3470 7261 3502
rect 7531 4286 7563 4318
rect 7531 4218 7563 4250
rect 7531 4150 7563 4182
rect 7531 4082 7563 4114
rect 7531 4014 7563 4046
rect 7531 3946 7563 3978
rect 7531 3878 7563 3910
rect 7531 3810 7563 3842
rect 7531 3742 7563 3774
rect 7531 3674 7563 3706
rect 7531 3606 7563 3638
rect 7531 3538 7563 3570
rect 7531 3470 7563 3502
rect 7833 4286 7865 4318
rect 7833 4218 7865 4250
rect 7833 4150 7865 4182
rect 7833 4082 7865 4114
rect 7833 4014 7865 4046
rect 7833 3946 7865 3978
rect 7833 3878 7865 3910
rect 7833 3810 7865 3842
rect 7833 3742 7865 3774
rect 7833 3674 7865 3706
rect 7833 3606 7865 3638
rect 7833 3538 7865 3570
rect 7833 3470 7865 3502
rect 8135 4286 8167 4318
rect 8135 4218 8167 4250
rect 8135 4150 8167 4182
rect 8135 4082 8167 4114
rect 8135 4014 8167 4046
rect 8135 3946 8167 3978
rect 8135 3878 8167 3910
rect 8135 3810 8167 3842
rect 8135 3742 8167 3774
rect 8135 3674 8167 3706
rect 8135 3606 8167 3638
rect 8135 3538 8167 3570
rect 8135 3470 8167 3502
rect 8437 4286 8469 4318
rect 8437 4218 8469 4250
rect 8437 4150 8469 4182
rect 8437 4082 8469 4114
rect 8437 4014 8469 4046
rect 8437 3946 8469 3978
rect 8437 3878 8469 3910
rect 8437 3810 8469 3842
rect 8437 3742 8469 3774
rect 8437 3674 8469 3706
rect 8437 3606 8469 3638
rect 8437 3538 8469 3570
rect 8437 3470 8469 3502
rect 8739 4286 8771 4318
rect 8739 4218 8771 4250
rect 8739 4150 8771 4182
rect 8739 4082 8771 4114
rect 8739 4014 8771 4046
rect 8739 3946 8771 3978
rect 8739 3878 8771 3910
rect 8739 3810 8771 3842
rect 8739 3742 8771 3774
rect 8739 3674 8771 3706
rect 8739 3606 8771 3638
rect 8739 3538 8771 3570
rect 8739 3470 8771 3502
rect 9041 4286 9073 4318
rect 9041 4218 9073 4250
rect 9041 4150 9073 4182
rect 9041 4082 9073 4114
rect 9041 4014 9073 4046
rect 9041 3946 9073 3978
rect 9041 3878 9073 3910
rect 9041 3810 9073 3842
rect 9041 3742 9073 3774
rect 9041 3674 9073 3706
rect 9041 3606 9073 3638
rect 9041 3538 9073 3570
rect 9041 3470 9073 3502
rect 9343 4286 9375 4318
rect 9343 4218 9375 4250
rect 9343 4150 9375 4182
rect 9343 4082 9375 4114
rect 9343 4014 9375 4046
rect 9343 3946 9375 3978
rect 9343 3878 9375 3910
rect 9343 3810 9375 3842
rect 9343 3742 9375 3774
rect 9343 3674 9375 3706
rect 9343 3606 9375 3638
rect 9343 3538 9375 3570
rect 9343 3470 9375 3502
rect 9645 4286 9677 4318
rect 9645 4218 9677 4250
rect 9645 4150 9677 4182
rect 9645 4082 9677 4114
rect 9645 4014 9677 4046
rect 9645 3946 9677 3978
rect 9645 3878 9677 3910
rect 9645 3810 9677 3842
rect 9645 3742 9677 3774
rect 9645 3674 9677 3706
rect 9645 3606 9677 3638
rect 9645 3538 9677 3570
rect 9645 3470 9677 3502
rect 9947 4286 9979 4318
rect 9947 4218 9979 4250
rect 9947 4150 9979 4182
rect 9947 4082 9979 4114
rect 9947 4014 9979 4046
rect 9947 3946 9979 3978
rect 9947 3878 9979 3910
rect 9947 3810 9979 3842
rect 9947 3742 9979 3774
rect 9947 3674 9979 3706
rect 9947 3606 9979 3638
rect 9947 3538 9979 3570
rect 9947 3470 9979 3502
rect 10249 4286 10281 4318
rect 10249 4218 10281 4250
rect 10249 4150 10281 4182
rect 10249 4082 10281 4114
rect 10249 4014 10281 4046
rect 10249 3946 10281 3978
rect 10249 3878 10281 3910
rect 10249 3810 10281 3842
rect 10249 3742 10281 3774
rect 10249 3674 10281 3706
rect 10249 3606 10281 3638
rect 10249 3538 10281 3570
rect 10249 3470 10281 3502
rect 10551 4286 10583 4318
rect 10551 4218 10583 4250
rect 10551 4150 10583 4182
rect 10551 4082 10583 4114
rect 10551 4014 10583 4046
rect 10551 3946 10583 3978
rect 10551 3878 10583 3910
rect 10551 3810 10583 3842
rect 10551 3742 10583 3774
rect 10551 3674 10583 3706
rect 10551 3606 10583 3638
rect 10551 3538 10583 3570
rect 10551 3470 10583 3502
rect 10853 4286 10885 4318
rect 10853 4218 10885 4250
rect 10853 4150 10885 4182
rect 10853 4082 10885 4114
rect 10853 4014 10885 4046
rect 10853 3946 10885 3978
rect 10853 3878 10885 3910
rect 10853 3810 10885 3842
rect 10853 3742 10885 3774
rect 10853 3674 10885 3706
rect 10853 3606 10885 3638
rect 10853 3538 10885 3570
rect 10853 3470 10885 3502
rect 11155 4286 11187 4318
rect 11155 4218 11187 4250
rect 11155 4150 11187 4182
rect 11155 4082 11187 4114
rect 11155 4014 11187 4046
rect 11155 3946 11187 3978
rect 11155 3878 11187 3910
rect 11155 3810 11187 3842
rect 11155 3742 11187 3774
rect 11155 3674 11187 3706
rect 11155 3606 11187 3638
rect 11155 3538 11187 3570
rect 11155 3470 11187 3502
rect 11457 4286 11489 4318
rect 11457 4218 11489 4250
rect 11457 4150 11489 4182
rect 11457 4082 11489 4114
rect 11457 4014 11489 4046
rect 11457 3946 11489 3978
rect 11457 3878 11489 3910
rect 11457 3810 11489 3842
rect 11457 3742 11489 3774
rect 11457 3674 11489 3706
rect 11457 3606 11489 3638
rect 11457 3538 11489 3570
rect 11457 3470 11489 3502
rect 11759 4286 11791 4318
rect 11759 4218 11791 4250
rect 11759 4150 11791 4182
rect 11759 4082 11791 4114
rect 11759 4014 11791 4046
rect 11759 3946 11791 3978
rect 11759 3878 11791 3910
rect 11759 3810 11791 3842
rect 11759 3742 11791 3774
rect 11759 3674 11791 3706
rect 11759 3606 11791 3638
rect 11759 3538 11791 3570
rect 11759 3470 11791 3502
rect 12061 4286 12093 4318
rect 12061 4218 12093 4250
rect 12061 4150 12093 4182
rect 12061 4082 12093 4114
rect 12061 4014 12093 4046
rect 12061 3946 12093 3978
rect 12061 3878 12093 3910
rect 12061 3810 12093 3842
rect 12061 3742 12093 3774
rect 12061 3674 12093 3706
rect 12061 3606 12093 3638
rect 12061 3538 12093 3570
rect 12061 3470 12093 3502
rect 12363 4286 12395 4318
rect 12363 4218 12395 4250
rect 12363 4150 12395 4182
rect 12363 4082 12395 4114
rect 12363 4014 12395 4046
rect 12363 3946 12395 3978
rect 12363 3878 12395 3910
rect 12363 3810 12395 3842
rect 12363 3742 12395 3774
rect 12363 3674 12395 3706
rect 12363 3606 12395 3638
rect 12363 3538 12395 3570
rect 12363 3470 12395 3502
rect 12665 4286 12697 4318
rect 12665 4218 12697 4250
rect 12665 4150 12697 4182
rect 12665 4082 12697 4114
rect 12665 4014 12697 4046
rect 12665 3946 12697 3978
rect 12665 3878 12697 3910
rect 12665 3810 12697 3842
rect 12665 3742 12697 3774
rect 12665 3674 12697 3706
rect 12665 3606 12697 3638
rect 12665 3538 12697 3570
rect 12665 3470 12697 3502
rect 12967 4286 12999 4318
rect 12967 4218 12999 4250
rect 12967 4150 12999 4182
rect 12967 4082 12999 4114
rect 12967 4014 12999 4046
rect 12967 3946 12999 3978
rect 12967 3878 12999 3910
rect 12967 3810 12999 3842
rect 12967 3742 12999 3774
rect 12967 3674 12999 3706
rect 12967 3606 12999 3638
rect 12967 3538 12999 3570
rect 12967 3470 12999 3502
rect 13269 4286 13301 4318
rect 13269 4218 13301 4250
rect 13269 4150 13301 4182
rect 13269 4082 13301 4114
rect 13269 4014 13301 4046
rect 13269 3946 13301 3978
rect 13269 3878 13301 3910
rect 13269 3810 13301 3842
rect 13269 3742 13301 3774
rect 13269 3674 13301 3706
rect 13269 3606 13301 3638
rect 13269 3538 13301 3570
rect 13269 3470 13301 3502
rect 13571 4286 13603 4318
rect 13571 4218 13603 4250
rect 13571 4150 13603 4182
rect 13571 4082 13603 4114
rect 13571 4014 13603 4046
rect 13571 3946 13603 3978
rect 13571 3878 13603 3910
rect 13571 3810 13603 3842
rect 13571 3742 13603 3774
rect 13571 3674 13603 3706
rect 13571 3606 13603 3638
rect 13571 3538 13603 3570
rect 13571 3470 13603 3502
rect 13873 4286 13905 4318
rect 13873 4218 13905 4250
rect 13873 4150 13905 4182
rect 13873 4082 13905 4114
rect 13873 4014 13905 4046
rect 13873 3946 13905 3978
rect 13873 3878 13905 3910
rect 13873 3810 13905 3842
rect 13873 3742 13905 3774
rect 13873 3674 13905 3706
rect 13873 3606 13905 3638
rect 13873 3538 13905 3570
rect 13873 3470 13905 3502
rect 14175 4286 14207 4318
rect 14175 4218 14207 4250
rect 14175 4150 14207 4182
rect 14175 4082 14207 4114
rect 14175 4014 14207 4046
rect 14175 3946 14207 3978
rect 14175 3878 14207 3910
rect 14175 3810 14207 3842
rect 14175 3742 14207 3774
rect 14175 3674 14207 3706
rect 14175 3606 14207 3638
rect 14175 3538 14207 3570
rect 14175 3470 14207 3502
rect 14477 4286 14509 4318
rect 14477 4218 14509 4250
rect 14477 4150 14509 4182
rect 14477 4082 14509 4114
rect 14477 4014 14509 4046
rect 14477 3946 14509 3978
rect 14477 3878 14509 3910
rect 14477 3810 14509 3842
rect 14477 3742 14509 3774
rect 14477 3674 14509 3706
rect 14477 3606 14509 3638
rect 14477 3538 14509 3570
rect 14477 3470 14509 3502
rect 1491 3318 1523 3350
rect 1491 3250 1523 3282
rect 1491 3182 1523 3214
rect 1491 3114 1523 3146
rect 1491 3046 1523 3078
rect 1491 2978 1523 3010
rect 1491 2910 1523 2942
rect 1491 2842 1523 2874
rect 1491 2774 1523 2806
rect 1491 2706 1523 2738
rect 1491 2638 1523 2670
rect 1491 2570 1523 2602
rect 1491 2502 1523 2534
rect 1793 3318 1825 3350
rect 1793 3250 1825 3282
rect 1793 3182 1825 3214
rect 1793 3114 1825 3146
rect 1793 3046 1825 3078
rect 1793 2978 1825 3010
rect 1793 2910 1825 2942
rect 1793 2842 1825 2874
rect 1793 2774 1825 2806
rect 1793 2706 1825 2738
rect 1793 2638 1825 2670
rect 1793 2570 1825 2602
rect 1793 2502 1825 2534
rect 2095 3318 2127 3350
rect 2095 3250 2127 3282
rect 2095 3182 2127 3214
rect 2095 3114 2127 3146
rect 2095 3046 2127 3078
rect 2095 2978 2127 3010
rect 2095 2910 2127 2942
rect 2095 2842 2127 2874
rect 2095 2774 2127 2806
rect 2095 2706 2127 2738
rect 2095 2638 2127 2670
rect 2095 2570 2127 2602
rect 2095 2502 2127 2534
rect 2397 3318 2429 3350
rect 2397 3250 2429 3282
rect 2397 3182 2429 3214
rect 2397 3114 2429 3146
rect 2397 3046 2429 3078
rect 2397 2978 2429 3010
rect 2397 2910 2429 2942
rect 2397 2842 2429 2874
rect 2397 2774 2429 2806
rect 2397 2706 2429 2738
rect 2397 2638 2429 2670
rect 2397 2570 2429 2602
rect 2397 2502 2429 2534
rect 2699 3318 2731 3350
rect 2699 3250 2731 3282
rect 2699 3182 2731 3214
rect 2699 3114 2731 3146
rect 2699 3046 2731 3078
rect 2699 2978 2731 3010
rect 2699 2910 2731 2942
rect 2699 2842 2731 2874
rect 2699 2774 2731 2806
rect 2699 2706 2731 2738
rect 2699 2638 2731 2670
rect 2699 2570 2731 2602
rect 2699 2502 2731 2534
rect 3001 3318 3033 3350
rect 3001 3250 3033 3282
rect 3001 3182 3033 3214
rect 3001 3114 3033 3146
rect 3001 3046 3033 3078
rect 3001 2978 3033 3010
rect 3001 2910 3033 2942
rect 3001 2842 3033 2874
rect 3001 2774 3033 2806
rect 3001 2706 3033 2738
rect 3001 2638 3033 2670
rect 3001 2570 3033 2602
rect 3001 2502 3033 2534
rect 3303 3318 3335 3350
rect 3303 3250 3335 3282
rect 3303 3182 3335 3214
rect 3303 3114 3335 3146
rect 3303 3046 3335 3078
rect 3303 2978 3335 3010
rect 3303 2910 3335 2942
rect 3303 2842 3335 2874
rect 3303 2774 3335 2806
rect 3303 2706 3335 2738
rect 3303 2638 3335 2670
rect 3303 2570 3335 2602
rect 3303 2502 3335 2534
rect 3605 3318 3637 3350
rect 3605 3250 3637 3282
rect 3605 3182 3637 3214
rect 3605 3114 3637 3146
rect 3605 3046 3637 3078
rect 3605 2978 3637 3010
rect 3605 2910 3637 2942
rect 3605 2842 3637 2874
rect 3605 2774 3637 2806
rect 3605 2706 3637 2738
rect 3605 2638 3637 2670
rect 3605 2570 3637 2602
rect 3605 2502 3637 2534
rect 3907 3318 3939 3350
rect 3907 3250 3939 3282
rect 3907 3182 3939 3214
rect 3907 3114 3939 3146
rect 3907 3046 3939 3078
rect 3907 2978 3939 3010
rect 3907 2910 3939 2942
rect 3907 2842 3939 2874
rect 3907 2774 3939 2806
rect 3907 2706 3939 2738
rect 3907 2638 3939 2670
rect 3907 2570 3939 2602
rect 3907 2502 3939 2534
rect 4209 3318 4241 3350
rect 4209 3250 4241 3282
rect 4209 3182 4241 3214
rect 4209 3114 4241 3146
rect 4209 3046 4241 3078
rect 4209 2978 4241 3010
rect 4209 2910 4241 2942
rect 4209 2842 4241 2874
rect 4209 2774 4241 2806
rect 4209 2706 4241 2738
rect 4209 2638 4241 2670
rect 4209 2570 4241 2602
rect 4209 2502 4241 2534
rect 4511 3318 4543 3350
rect 4511 3250 4543 3282
rect 4511 3182 4543 3214
rect 4511 3114 4543 3146
rect 4511 3046 4543 3078
rect 4511 2978 4543 3010
rect 4511 2910 4543 2942
rect 4511 2842 4543 2874
rect 4511 2774 4543 2806
rect 4511 2706 4543 2738
rect 4511 2638 4543 2670
rect 4511 2570 4543 2602
rect 4511 2502 4543 2534
rect 4813 3318 4845 3350
rect 4813 3250 4845 3282
rect 4813 3182 4845 3214
rect 4813 3114 4845 3146
rect 4813 3046 4845 3078
rect 4813 2978 4845 3010
rect 4813 2910 4845 2942
rect 4813 2842 4845 2874
rect 4813 2774 4845 2806
rect 4813 2706 4845 2738
rect 4813 2638 4845 2670
rect 4813 2570 4845 2602
rect 4813 2502 4845 2534
rect 5115 3318 5147 3350
rect 5115 3250 5147 3282
rect 5115 3182 5147 3214
rect 5115 3114 5147 3146
rect 5115 3046 5147 3078
rect 5115 2978 5147 3010
rect 5115 2910 5147 2942
rect 5115 2842 5147 2874
rect 5115 2774 5147 2806
rect 5115 2706 5147 2738
rect 5115 2638 5147 2670
rect 5115 2570 5147 2602
rect 5115 2502 5147 2534
rect 5417 3318 5449 3350
rect 5417 3250 5449 3282
rect 5417 3182 5449 3214
rect 5417 3114 5449 3146
rect 5417 3046 5449 3078
rect 5417 2978 5449 3010
rect 5417 2910 5449 2942
rect 5417 2842 5449 2874
rect 5417 2774 5449 2806
rect 5417 2706 5449 2738
rect 5417 2638 5449 2670
rect 5417 2570 5449 2602
rect 5417 2502 5449 2534
rect 5719 3318 5751 3350
rect 5719 3250 5751 3282
rect 5719 3182 5751 3214
rect 5719 3114 5751 3146
rect 5719 3046 5751 3078
rect 5719 2978 5751 3010
rect 5719 2910 5751 2942
rect 5719 2842 5751 2874
rect 5719 2774 5751 2806
rect 5719 2706 5751 2738
rect 5719 2638 5751 2670
rect 5719 2570 5751 2602
rect 5719 2502 5751 2534
rect 6021 3318 6053 3350
rect 6021 3250 6053 3282
rect 6021 3182 6053 3214
rect 6021 3114 6053 3146
rect 6021 3046 6053 3078
rect 6021 2978 6053 3010
rect 6021 2910 6053 2942
rect 6021 2842 6053 2874
rect 6021 2774 6053 2806
rect 6021 2706 6053 2738
rect 6021 2638 6053 2670
rect 6021 2570 6053 2602
rect 6021 2502 6053 2534
rect 6323 3318 6355 3350
rect 6323 3250 6355 3282
rect 6323 3182 6355 3214
rect 6323 3114 6355 3146
rect 6323 3046 6355 3078
rect 6323 2978 6355 3010
rect 6323 2910 6355 2942
rect 6323 2842 6355 2874
rect 6323 2774 6355 2806
rect 6323 2706 6355 2738
rect 6323 2638 6355 2670
rect 6323 2570 6355 2602
rect 6323 2502 6355 2534
rect 6625 3318 6657 3350
rect 6625 3250 6657 3282
rect 6625 3182 6657 3214
rect 6625 3114 6657 3146
rect 6625 3046 6657 3078
rect 6625 2978 6657 3010
rect 6625 2910 6657 2942
rect 6625 2842 6657 2874
rect 6625 2774 6657 2806
rect 6625 2706 6657 2738
rect 6625 2638 6657 2670
rect 6625 2570 6657 2602
rect 6625 2502 6657 2534
rect 6927 3318 6959 3350
rect 6927 3250 6959 3282
rect 6927 3182 6959 3214
rect 6927 3114 6959 3146
rect 6927 3046 6959 3078
rect 6927 2978 6959 3010
rect 6927 2910 6959 2942
rect 6927 2842 6959 2874
rect 6927 2774 6959 2806
rect 6927 2706 6959 2738
rect 6927 2638 6959 2670
rect 6927 2570 6959 2602
rect 6927 2502 6959 2534
rect 7229 3318 7261 3350
rect 7229 3250 7261 3282
rect 7229 3182 7261 3214
rect 7229 3114 7261 3146
rect 7229 3046 7261 3078
rect 7229 2978 7261 3010
rect 7229 2910 7261 2942
rect 7229 2842 7261 2874
rect 7229 2774 7261 2806
rect 7229 2706 7261 2738
rect 7229 2638 7261 2670
rect 7229 2570 7261 2602
rect 7229 2502 7261 2534
rect 7531 3318 7563 3350
rect 7531 3250 7563 3282
rect 7531 3182 7563 3214
rect 7531 3114 7563 3146
rect 7531 3046 7563 3078
rect 7531 2978 7563 3010
rect 7531 2910 7563 2942
rect 7531 2842 7563 2874
rect 7531 2774 7563 2806
rect 7531 2706 7563 2738
rect 7531 2638 7563 2670
rect 7531 2570 7563 2602
rect 7531 2502 7563 2534
rect 7833 3318 7865 3350
rect 7833 3250 7865 3282
rect 7833 3182 7865 3214
rect 7833 3114 7865 3146
rect 7833 3046 7865 3078
rect 7833 2978 7865 3010
rect 7833 2910 7865 2942
rect 7833 2842 7865 2874
rect 7833 2774 7865 2806
rect 7833 2706 7865 2738
rect 7833 2638 7865 2670
rect 7833 2570 7865 2602
rect 7833 2502 7865 2534
rect 8135 3318 8167 3350
rect 8135 3250 8167 3282
rect 8135 3182 8167 3214
rect 8135 3114 8167 3146
rect 8135 3046 8167 3078
rect 8135 2978 8167 3010
rect 8135 2910 8167 2942
rect 8135 2842 8167 2874
rect 8135 2774 8167 2806
rect 8135 2706 8167 2738
rect 8135 2638 8167 2670
rect 8135 2570 8167 2602
rect 8135 2502 8167 2534
rect 8437 3318 8469 3350
rect 8437 3250 8469 3282
rect 8437 3182 8469 3214
rect 8437 3114 8469 3146
rect 8437 3046 8469 3078
rect 8437 2978 8469 3010
rect 8437 2910 8469 2942
rect 8437 2842 8469 2874
rect 8437 2774 8469 2806
rect 8437 2706 8469 2738
rect 8437 2638 8469 2670
rect 8437 2570 8469 2602
rect 8437 2502 8469 2534
rect 8739 3318 8771 3350
rect 8739 3250 8771 3282
rect 8739 3182 8771 3214
rect 8739 3114 8771 3146
rect 8739 3046 8771 3078
rect 8739 2978 8771 3010
rect 8739 2910 8771 2942
rect 8739 2842 8771 2874
rect 8739 2774 8771 2806
rect 8739 2706 8771 2738
rect 8739 2638 8771 2670
rect 8739 2570 8771 2602
rect 8739 2502 8771 2534
rect 9041 3318 9073 3350
rect 9041 3250 9073 3282
rect 9041 3182 9073 3214
rect 9041 3114 9073 3146
rect 9041 3046 9073 3078
rect 9041 2978 9073 3010
rect 9041 2910 9073 2942
rect 9041 2842 9073 2874
rect 9041 2774 9073 2806
rect 9041 2706 9073 2738
rect 9041 2638 9073 2670
rect 9041 2570 9073 2602
rect 9041 2502 9073 2534
rect 9343 3318 9375 3350
rect 9343 3250 9375 3282
rect 9343 3182 9375 3214
rect 9343 3114 9375 3146
rect 9343 3046 9375 3078
rect 9343 2978 9375 3010
rect 9343 2910 9375 2942
rect 9343 2842 9375 2874
rect 9343 2774 9375 2806
rect 9343 2706 9375 2738
rect 9343 2638 9375 2670
rect 9343 2570 9375 2602
rect 9343 2502 9375 2534
rect 9645 3318 9677 3350
rect 9645 3250 9677 3282
rect 9645 3182 9677 3214
rect 9645 3114 9677 3146
rect 9645 3046 9677 3078
rect 9645 2978 9677 3010
rect 9645 2910 9677 2942
rect 9645 2842 9677 2874
rect 9645 2774 9677 2806
rect 9645 2706 9677 2738
rect 9645 2638 9677 2670
rect 9645 2570 9677 2602
rect 9645 2502 9677 2534
rect 9947 3318 9979 3350
rect 9947 3250 9979 3282
rect 9947 3182 9979 3214
rect 9947 3114 9979 3146
rect 9947 3046 9979 3078
rect 9947 2978 9979 3010
rect 9947 2910 9979 2942
rect 9947 2842 9979 2874
rect 9947 2774 9979 2806
rect 9947 2706 9979 2738
rect 9947 2638 9979 2670
rect 9947 2570 9979 2602
rect 9947 2502 9979 2534
rect 10249 3318 10281 3350
rect 10249 3250 10281 3282
rect 10249 3182 10281 3214
rect 10249 3114 10281 3146
rect 10249 3046 10281 3078
rect 10249 2978 10281 3010
rect 10249 2910 10281 2942
rect 10249 2842 10281 2874
rect 10249 2774 10281 2806
rect 10249 2706 10281 2738
rect 10249 2638 10281 2670
rect 10249 2570 10281 2602
rect 10249 2502 10281 2534
rect 10551 3318 10583 3350
rect 10551 3250 10583 3282
rect 10551 3182 10583 3214
rect 10551 3114 10583 3146
rect 10551 3046 10583 3078
rect 10551 2978 10583 3010
rect 10551 2910 10583 2942
rect 10551 2842 10583 2874
rect 10551 2774 10583 2806
rect 10551 2706 10583 2738
rect 10551 2638 10583 2670
rect 10551 2570 10583 2602
rect 10551 2502 10583 2534
rect 10853 3318 10885 3350
rect 10853 3250 10885 3282
rect 10853 3182 10885 3214
rect 10853 3114 10885 3146
rect 10853 3046 10885 3078
rect 10853 2978 10885 3010
rect 10853 2910 10885 2942
rect 10853 2842 10885 2874
rect 10853 2774 10885 2806
rect 10853 2706 10885 2738
rect 10853 2638 10885 2670
rect 10853 2570 10885 2602
rect 10853 2502 10885 2534
rect 11155 3318 11187 3350
rect 11155 3250 11187 3282
rect 11155 3182 11187 3214
rect 11155 3114 11187 3146
rect 11155 3046 11187 3078
rect 11155 2978 11187 3010
rect 11155 2910 11187 2942
rect 11155 2842 11187 2874
rect 11155 2774 11187 2806
rect 11155 2706 11187 2738
rect 11155 2638 11187 2670
rect 11155 2570 11187 2602
rect 11155 2502 11187 2534
rect 11457 3318 11489 3350
rect 11457 3250 11489 3282
rect 11457 3182 11489 3214
rect 11457 3114 11489 3146
rect 11457 3046 11489 3078
rect 11457 2978 11489 3010
rect 11457 2910 11489 2942
rect 11457 2842 11489 2874
rect 11457 2774 11489 2806
rect 11457 2706 11489 2738
rect 11457 2638 11489 2670
rect 11457 2570 11489 2602
rect 11457 2502 11489 2534
rect 11759 3318 11791 3350
rect 11759 3250 11791 3282
rect 11759 3182 11791 3214
rect 11759 3114 11791 3146
rect 11759 3046 11791 3078
rect 11759 2978 11791 3010
rect 11759 2910 11791 2942
rect 11759 2842 11791 2874
rect 11759 2774 11791 2806
rect 11759 2706 11791 2738
rect 11759 2638 11791 2670
rect 11759 2570 11791 2602
rect 11759 2502 11791 2534
rect 12061 3318 12093 3350
rect 12061 3250 12093 3282
rect 12061 3182 12093 3214
rect 12061 3114 12093 3146
rect 12061 3046 12093 3078
rect 12061 2978 12093 3010
rect 12061 2910 12093 2942
rect 12061 2842 12093 2874
rect 12061 2774 12093 2806
rect 12061 2706 12093 2738
rect 12061 2638 12093 2670
rect 12061 2570 12093 2602
rect 12061 2502 12093 2534
rect 12363 3318 12395 3350
rect 12363 3250 12395 3282
rect 12363 3182 12395 3214
rect 12363 3114 12395 3146
rect 12363 3046 12395 3078
rect 12363 2978 12395 3010
rect 12363 2910 12395 2942
rect 12363 2842 12395 2874
rect 12363 2774 12395 2806
rect 12363 2706 12395 2738
rect 12363 2638 12395 2670
rect 12363 2570 12395 2602
rect 12363 2502 12395 2534
rect 12665 3318 12697 3350
rect 12665 3250 12697 3282
rect 12665 3182 12697 3214
rect 12665 3114 12697 3146
rect 12665 3046 12697 3078
rect 12665 2978 12697 3010
rect 12665 2910 12697 2942
rect 12665 2842 12697 2874
rect 12665 2774 12697 2806
rect 12665 2706 12697 2738
rect 12665 2638 12697 2670
rect 12665 2570 12697 2602
rect 12665 2502 12697 2534
rect 12967 3318 12999 3350
rect 12967 3250 12999 3282
rect 12967 3182 12999 3214
rect 12967 3114 12999 3146
rect 12967 3046 12999 3078
rect 12967 2978 12999 3010
rect 12967 2910 12999 2942
rect 12967 2842 12999 2874
rect 12967 2774 12999 2806
rect 12967 2706 12999 2738
rect 12967 2638 12999 2670
rect 12967 2570 12999 2602
rect 12967 2502 12999 2534
rect 13269 3318 13301 3350
rect 13269 3250 13301 3282
rect 13269 3182 13301 3214
rect 13269 3114 13301 3146
rect 13269 3046 13301 3078
rect 13269 2978 13301 3010
rect 13269 2910 13301 2942
rect 13269 2842 13301 2874
rect 13269 2774 13301 2806
rect 13269 2706 13301 2738
rect 13269 2638 13301 2670
rect 13269 2570 13301 2602
rect 13269 2502 13301 2534
rect 13571 3318 13603 3350
rect 13571 3250 13603 3282
rect 13571 3182 13603 3214
rect 13571 3114 13603 3146
rect 13571 3046 13603 3078
rect 13571 2978 13603 3010
rect 13571 2910 13603 2942
rect 13571 2842 13603 2874
rect 13571 2774 13603 2806
rect 13571 2706 13603 2738
rect 13571 2638 13603 2670
rect 13571 2570 13603 2602
rect 13571 2502 13603 2534
rect 13873 3318 13905 3350
rect 13873 3250 13905 3282
rect 13873 3182 13905 3214
rect 13873 3114 13905 3146
rect 13873 3046 13905 3078
rect 13873 2978 13905 3010
rect 13873 2910 13905 2942
rect 13873 2842 13905 2874
rect 13873 2774 13905 2806
rect 13873 2706 13905 2738
rect 13873 2638 13905 2670
rect 13873 2570 13905 2602
rect 13873 2502 13905 2534
rect 14175 3318 14207 3350
rect 14175 3250 14207 3282
rect 14175 3182 14207 3214
rect 14175 3114 14207 3146
rect 14175 3046 14207 3078
rect 14175 2978 14207 3010
rect 14175 2910 14207 2942
rect 14175 2842 14207 2874
rect 14175 2774 14207 2806
rect 14175 2706 14207 2738
rect 14175 2638 14207 2670
rect 14175 2570 14207 2602
rect 14175 2502 14207 2534
rect 14477 3318 14509 3350
rect 14477 3250 14509 3282
rect 14477 3182 14509 3214
rect 14477 3114 14509 3146
rect 14477 3046 14509 3078
rect 14477 2978 14509 3010
rect 14477 2910 14509 2942
rect 14477 2842 14509 2874
rect 14477 2774 14509 2806
rect 14477 2706 14509 2738
rect 14477 2638 14509 2670
rect 14477 2570 14509 2602
rect 14477 2502 14509 2534
rect 1491 2350 1523 2382
rect 1491 2282 1523 2314
rect 1491 2214 1523 2246
rect 1491 2146 1523 2178
rect 1491 2078 1523 2110
rect 1491 2010 1523 2042
rect 1491 1942 1523 1974
rect 1491 1874 1523 1906
rect 1491 1806 1523 1838
rect 1491 1738 1523 1770
rect 1491 1670 1523 1702
rect 1491 1602 1523 1634
rect 1491 1534 1523 1566
rect 1793 2350 1825 2382
rect 1793 2282 1825 2314
rect 1793 2214 1825 2246
rect 1793 2146 1825 2178
rect 1793 2078 1825 2110
rect 1793 2010 1825 2042
rect 1793 1942 1825 1974
rect 1793 1874 1825 1906
rect 1793 1806 1825 1838
rect 1793 1738 1825 1770
rect 1793 1670 1825 1702
rect 1793 1602 1825 1634
rect 1793 1534 1825 1566
rect 2095 2350 2127 2382
rect 2095 2282 2127 2314
rect 2095 2214 2127 2246
rect 2095 2146 2127 2178
rect 2095 2078 2127 2110
rect 2095 2010 2127 2042
rect 2095 1942 2127 1974
rect 2095 1874 2127 1906
rect 2095 1806 2127 1838
rect 2095 1738 2127 1770
rect 2095 1670 2127 1702
rect 2095 1602 2127 1634
rect 2095 1534 2127 1566
rect 2397 2350 2429 2382
rect 2397 2282 2429 2314
rect 2397 2214 2429 2246
rect 2397 2146 2429 2178
rect 2397 2078 2429 2110
rect 2397 2010 2429 2042
rect 2397 1942 2429 1974
rect 2397 1874 2429 1906
rect 2397 1806 2429 1838
rect 2397 1738 2429 1770
rect 2397 1670 2429 1702
rect 2397 1602 2429 1634
rect 2397 1534 2429 1566
rect 2699 2350 2731 2382
rect 2699 2282 2731 2314
rect 2699 2214 2731 2246
rect 2699 2146 2731 2178
rect 2699 2078 2731 2110
rect 2699 2010 2731 2042
rect 2699 1942 2731 1974
rect 2699 1874 2731 1906
rect 2699 1806 2731 1838
rect 2699 1738 2731 1770
rect 2699 1670 2731 1702
rect 2699 1602 2731 1634
rect 2699 1534 2731 1566
rect 3001 2350 3033 2382
rect 3001 2282 3033 2314
rect 3001 2214 3033 2246
rect 3001 2146 3033 2178
rect 3001 2078 3033 2110
rect 3001 2010 3033 2042
rect 3001 1942 3033 1974
rect 3001 1874 3033 1906
rect 3001 1806 3033 1838
rect 3001 1738 3033 1770
rect 3001 1670 3033 1702
rect 3001 1602 3033 1634
rect 3001 1534 3033 1566
rect 3303 2350 3335 2382
rect 3303 2282 3335 2314
rect 3303 2214 3335 2246
rect 3303 2146 3335 2178
rect 3303 2078 3335 2110
rect 3303 2010 3335 2042
rect 3303 1942 3335 1974
rect 3303 1874 3335 1906
rect 3303 1806 3335 1838
rect 3303 1738 3335 1770
rect 3303 1670 3335 1702
rect 3303 1602 3335 1634
rect 3303 1534 3335 1566
rect 3605 2350 3637 2382
rect 3605 2282 3637 2314
rect 3605 2214 3637 2246
rect 3605 2146 3637 2178
rect 3605 2078 3637 2110
rect 3605 2010 3637 2042
rect 3605 1942 3637 1974
rect 3605 1874 3637 1906
rect 3605 1806 3637 1838
rect 3605 1738 3637 1770
rect 3605 1670 3637 1702
rect 3605 1602 3637 1634
rect 3605 1534 3637 1566
rect 3907 2350 3939 2382
rect 3907 2282 3939 2314
rect 3907 2214 3939 2246
rect 3907 2146 3939 2178
rect 3907 2078 3939 2110
rect 3907 2010 3939 2042
rect 3907 1942 3939 1974
rect 3907 1874 3939 1906
rect 3907 1806 3939 1838
rect 3907 1738 3939 1770
rect 3907 1670 3939 1702
rect 3907 1602 3939 1634
rect 3907 1534 3939 1566
rect 4209 2350 4241 2382
rect 4209 2282 4241 2314
rect 4209 2214 4241 2246
rect 4209 2146 4241 2178
rect 4209 2078 4241 2110
rect 4209 2010 4241 2042
rect 4209 1942 4241 1974
rect 4209 1874 4241 1906
rect 4209 1806 4241 1838
rect 4209 1738 4241 1770
rect 4209 1670 4241 1702
rect 4209 1602 4241 1634
rect 4209 1534 4241 1566
rect 4511 2350 4543 2382
rect 4511 2282 4543 2314
rect 4511 2214 4543 2246
rect 4511 2146 4543 2178
rect 4511 2078 4543 2110
rect 4511 2010 4543 2042
rect 4511 1942 4543 1974
rect 4511 1874 4543 1906
rect 4511 1806 4543 1838
rect 4511 1738 4543 1770
rect 4511 1670 4543 1702
rect 4511 1602 4543 1634
rect 4511 1534 4543 1566
rect 4813 2350 4845 2382
rect 4813 2282 4845 2314
rect 4813 2214 4845 2246
rect 4813 2146 4845 2178
rect 4813 2078 4845 2110
rect 4813 2010 4845 2042
rect 4813 1942 4845 1974
rect 4813 1874 4845 1906
rect 4813 1806 4845 1838
rect 4813 1738 4845 1770
rect 4813 1670 4845 1702
rect 4813 1602 4845 1634
rect 4813 1534 4845 1566
rect 5115 2350 5147 2382
rect 5115 2282 5147 2314
rect 5115 2214 5147 2246
rect 5115 2146 5147 2178
rect 5115 2078 5147 2110
rect 5115 2010 5147 2042
rect 5115 1942 5147 1974
rect 5115 1874 5147 1906
rect 5115 1806 5147 1838
rect 5115 1738 5147 1770
rect 5115 1670 5147 1702
rect 5115 1602 5147 1634
rect 5115 1534 5147 1566
rect 5417 2350 5449 2382
rect 5417 2282 5449 2314
rect 5417 2214 5449 2246
rect 5417 2146 5449 2178
rect 5417 2078 5449 2110
rect 5417 2010 5449 2042
rect 5417 1942 5449 1974
rect 5417 1874 5449 1906
rect 5417 1806 5449 1838
rect 5417 1738 5449 1770
rect 5417 1670 5449 1702
rect 5417 1602 5449 1634
rect 5417 1534 5449 1566
rect 5719 2350 5751 2382
rect 5719 2282 5751 2314
rect 5719 2214 5751 2246
rect 5719 2146 5751 2178
rect 5719 2078 5751 2110
rect 5719 2010 5751 2042
rect 5719 1942 5751 1974
rect 5719 1874 5751 1906
rect 5719 1806 5751 1838
rect 5719 1738 5751 1770
rect 5719 1670 5751 1702
rect 5719 1602 5751 1634
rect 5719 1534 5751 1566
rect 6021 2350 6053 2382
rect 6021 2282 6053 2314
rect 6021 2214 6053 2246
rect 6021 2146 6053 2178
rect 6021 2078 6053 2110
rect 6021 2010 6053 2042
rect 6021 1942 6053 1974
rect 6021 1874 6053 1906
rect 6021 1806 6053 1838
rect 6021 1738 6053 1770
rect 6021 1670 6053 1702
rect 6021 1602 6053 1634
rect 6021 1534 6053 1566
rect 6323 2350 6355 2382
rect 6323 2282 6355 2314
rect 6323 2214 6355 2246
rect 6323 2146 6355 2178
rect 6323 2078 6355 2110
rect 6323 2010 6355 2042
rect 6323 1942 6355 1974
rect 6323 1874 6355 1906
rect 6323 1806 6355 1838
rect 6323 1738 6355 1770
rect 6323 1670 6355 1702
rect 6323 1602 6355 1634
rect 6323 1534 6355 1566
rect 6625 2350 6657 2382
rect 6625 2282 6657 2314
rect 6625 2214 6657 2246
rect 6625 2146 6657 2178
rect 6625 2078 6657 2110
rect 6625 2010 6657 2042
rect 6625 1942 6657 1974
rect 6625 1874 6657 1906
rect 6625 1806 6657 1838
rect 6625 1738 6657 1770
rect 6625 1670 6657 1702
rect 6625 1602 6657 1634
rect 6625 1534 6657 1566
rect 6927 2350 6959 2382
rect 6927 2282 6959 2314
rect 6927 2214 6959 2246
rect 6927 2146 6959 2178
rect 6927 2078 6959 2110
rect 6927 2010 6959 2042
rect 6927 1942 6959 1974
rect 6927 1874 6959 1906
rect 6927 1806 6959 1838
rect 6927 1738 6959 1770
rect 6927 1670 6959 1702
rect 6927 1602 6959 1634
rect 6927 1534 6959 1566
rect 7229 2350 7261 2382
rect 7229 2282 7261 2314
rect 7229 2214 7261 2246
rect 7229 2146 7261 2178
rect 7229 2078 7261 2110
rect 7229 2010 7261 2042
rect 7229 1942 7261 1974
rect 7229 1874 7261 1906
rect 7229 1806 7261 1838
rect 7229 1738 7261 1770
rect 7229 1670 7261 1702
rect 7229 1602 7261 1634
rect 7229 1534 7261 1566
rect 7531 2350 7563 2382
rect 7531 2282 7563 2314
rect 7531 2214 7563 2246
rect 7531 2146 7563 2178
rect 7531 2078 7563 2110
rect 7531 2010 7563 2042
rect 7531 1942 7563 1974
rect 7531 1874 7563 1906
rect 7531 1806 7563 1838
rect 7531 1738 7563 1770
rect 7531 1670 7563 1702
rect 7531 1602 7563 1634
rect 7531 1534 7563 1566
rect 7833 2350 7865 2382
rect 7833 2282 7865 2314
rect 7833 2214 7865 2246
rect 7833 2146 7865 2178
rect 7833 2078 7865 2110
rect 7833 2010 7865 2042
rect 7833 1942 7865 1974
rect 7833 1874 7865 1906
rect 7833 1806 7865 1838
rect 7833 1738 7865 1770
rect 7833 1670 7865 1702
rect 7833 1602 7865 1634
rect 7833 1534 7865 1566
rect 8135 2350 8167 2382
rect 8135 2282 8167 2314
rect 8135 2214 8167 2246
rect 8135 2146 8167 2178
rect 8135 2078 8167 2110
rect 8135 2010 8167 2042
rect 8135 1942 8167 1974
rect 8135 1874 8167 1906
rect 8135 1806 8167 1838
rect 8135 1738 8167 1770
rect 8135 1670 8167 1702
rect 8135 1602 8167 1634
rect 8135 1534 8167 1566
rect 8437 2350 8469 2382
rect 8437 2282 8469 2314
rect 8437 2214 8469 2246
rect 8437 2146 8469 2178
rect 8437 2078 8469 2110
rect 8437 2010 8469 2042
rect 8437 1942 8469 1974
rect 8437 1874 8469 1906
rect 8437 1806 8469 1838
rect 8437 1738 8469 1770
rect 8437 1670 8469 1702
rect 8437 1602 8469 1634
rect 8437 1534 8469 1566
rect 8739 2350 8771 2382
rect 8739 2282 8771 2314
rect 8739 2214 8771 2246
rect 8739 2146 8771 2178
rect 8739 2078 8771 2110
rect 8739 2010 8771 2042
rect 8739 1942 8771 1974
rect 8739 1874 8771 1906
rect 8739 1806 8771 1838
rect 8739 1738 8771 1770
rect 8739 1670 8771 1702
rect 8739 1602 8771 1634
rect 8739 1534 8771 1566
rect 9041 2350 9073 2382
rect 9041 2282 9073 2314
rect 9041 2214 9073 2246
rect 9041 2146 9073 2178
rect 9041 2078 9073 2110
rect 9041 2010 9073 2042
rect 9041 1942 9073 1974
rect 9041 1874 9073 1906
rect 9041 1806 9073 1838
rect 9041 1738 9073 1770
rect 9041 1670 9073 1702
rect 9041 1602 9073 1634
rect 9041 1534 9073 1566
rect 9343 2350 9375 2382
rect 9343 2282 9375 2314
rect 9343 2214 9375 2246
rect 9343 2146 9375 2178
rect 9343 2078 9375 2110
rect 9343 2010 9375 2042
rect 9343 1942 9375 1974
rect 9343 1874 9375 1906
rect 9343 1806 9375 1838
rect 9343 1738 9375 1770
rect 9343 1670 9375 1702
rect 9343 1602 9375 1634
rect 9343 1534 9375 1566
rect 9645 2350 9677 2382
rect 9645 2282 9677 2314
rect 9645 2214 9677 2246
rect 9645 2146 9677 2178
rect 9645 2078 9677 2110
rect 9645 2010 9677 2042
rect 9645 1942 9677 1974
rect 9645 1874 9677 1906
rect 9645 1806 9677 1838
rect 9645 1738 9677 1770
rect 9645 1670 9677 1702
rect 9645 1602 9677 1634
rect 9645 1534 9677 1566
rect 9947 2350 9979 2382
rect 9947 2282 9979 2314
rect 9947 2214 9979 2246
rect 9947 2146 9979 2178
rect 9947 2078 9979 2110
rect 9947 2010 9979 2042
rect 9947 1942 9979 1974
rect 9947 1874 9979 1906
rect 9947 1806 9979 1838
rect 9947 1738 9979 1770
rect 9947 1670 9979 1702
rect 9947 1602 9979 1634
rect 9947 1534 9979 1566
rect 10249 2350 10281 2382
rect 10249 2282 10281 2314
rect 10249 2214 10281 2246
rect 10249 2146 10281 2178
rect 10249 2078 10281 2110
rect 10249 2010 10281 2042
rect 10249 1942 10281 1974
rect 10249 1874 10281 1906
rect 10249 1806 10281 1838
rect 10249 1738 10281 1770
rect 10249 1670 10281 1702
rect 10249 1602 10281 1634
rect 10249 1534 10281 1566
rect 10551 2350 10583 2382
rect 10551 2282 10583 2314
rect 10551 2214 10583 2246
rect 10551 2146 10583 2178
rect 10551 2078 10583 2110
rect 10551 2010 10583 2042
rect 10551 1942 10583 1974
rect 10551 1874 10583 1906
rect 10551 1806 10583 1838
rect 10551 1738 10583 1770
rect 10551 1670 10583 1702
rect 10551 1602 10583 1634
rect 10551 1534 10583 1566
rect 10853 2350 10885 2382
rect 10853 2282 10885 2314
rect 10853 2214 10885 2246
rect 10853 2146 10885 2178
rect 10853 2078 10885 2110
rect 10853 2010 10885 2042
rect 10853 1942 10885 1974
rect 10853 1874 10885 1906
rect 10853 1806 10885 1838
rect 10853 1738 10885 1770
rect 10853 1670 10885 1702
rect 10853 1602 10885 1634
rect 10853 1534 10885 1566
rect 11155 2350 11187 2382
rect 11155 2282 11187 2314
rect 11155 2214 11187 2246
rect 11155 2146 11187 2178
rect 11155 2078 11187 2110
rect 11155 2010 11187 2042
rect 11155 1942 11187 1974
rect 11155 1874 11187 1906
rect 11155 1806 11187 1838
rect 11155 1738 11187 1770
rect 11155 1670 11187 1702
rect 11155 1602 11187 1634
rect 11155 1534 11187 1566
rect 11457 2350 11489 2382
rect 11457 2282 11489 2314
rect 11457 2214 11489 2246
rect 11457 2146 11489 2178
rect 11457 2078 11489 2110
rect 11457 2010 11489 2042
rect 11457 1942 11489 1974
rect 11457 1874 11489 1906
rect 11457 1806 11489 1838
rect 11457 1738 11489 1770
rect 11457 1670 11489 1702
rect 11457 1602 11489 1634
rect 11457 1534 11489 1566
rect 11759 2350 11791 2382
rect 11759 2282 11791 2314
rect 11759 2214 11791 2246
rect 11759 2146 11791 2178
rect 11759 2078 11791 2110
rect 11759 2010 11791 2042
rect 11759 1942 11791 1974
rect 11759 1874 11791 1906
rect 11759 1806 11791 1838
rect 11759 1738 11791 1770
rect 11759 1670 11791 1702
rect 11759 1602 11791 1634
rect 11759 1534 11791 1566
rect 12061 2350 12093 2382
rect 12061 2282 12093 2314
rect 12061 2214 12093 2246
rect 12061 2146 12093 2178
rect 12061 2078 12093 2110
rect 12061 2010 12093 2042
rect 12061 1942 12093 1974
rect 12061 1874 12093 1906
rect 12061 1806 12093 1838
rect 12061 1738 12093 1770
rect 12061 1670 12093 1702
rect 12061 1602 12093 1634
rect 12061 1534 12093 1566
rect 12363 2350 12395 2382
rect 12363 2282 12395 2314
rect 12363 2214 12395 2246
rect 12363 2146 12395 2178
rect 12363 2078 12395 2110
rect 12363 2010 12395 2042
rect 12363 1942 12395 1974
rect 12363 1874 12395 1906
rect 12363 1806 12395 1838
rect 12363 1738 12395 1770
rect 12363 1670 12395 1702
rect 12363 1602 12395 1634
rect 12363 1534 12395 1566
rect 12665 2350 12697 2382
rect 12665 2282 12697 2314
rect 12665 2214 12697 2246
rect 12665 2146 12697 2178
rect 12665 2078 12697 2110
rect 12665 2010 12697 2042
rect 12665 1942 12697 1974
rect 12665 1874 12697 1906
rect 12665 1806 12697 1838
rect 12665 1738 12697 1770
rect 12665 1670 12697 1702
rect 12665 1602 12697 1634
rect 12665 1534 12697 1566
rect 12967 2350 12999 2382
rect 12967 2282 12999 2314
rect 12967 2214 12999 2246
rect 12967 2146 12999 2178
rect 12967 2078 12999 2110
rect 12967 2010 12999 2042
rect 12967 1942 12999 1974
rect 12967 1874 12999 1906
rect 12967 1806 12999 1838
rect 12967 1738 12999 1770
rect 12967 1670 12999 1702
rect 12967 1602 12999 1634
rect 12967 1534 12999 1566
rect 13269 2350 13301 2382
rect 13269 2282 13301 2314
rect 13269 2214 13301 2246
rect 13269 2146 13301 2178
rect 13269 2078 13301 2110
rect 13269 2010 13301 2042
rect 13269 1942 13301 1974
rect 13269 1874 13301 1906
rect 13269 1806 13301 1838
rect 13269 1738 13301 1770
rect 13269 1670 13301 1702
rect 13269 1602 13301 1634
rect 13269 1534 13301 1566
rect 13571 2350 13603 2382
rect 13571 2282 13603 2314
rect 13571 2214 13603 2246
rect 13571 2146 13603 2178
rect 13571 2078 13603 2110
rect 13571 2010 13603 2042
rect 13571 1942 13603 1974
rect 13571 1874 13603 1906
rect 13571 1806 13603 1838
rect 13571 1738 13603 1770
rect 13571 1670 13603 1702
rect 13571 1602 13603 1634
rect 13571 1534 13603 1566
rect 13873 2350 13905 2382
rect 13873 2282 13905 2314
rect 13873 2214 13905 2246
rect 13873 2146 13905 2178
rect 13873 2078 13905 2110
rect 13873 2010 13905 2042
rect 13873 1942 13905 1974
rect 13873 1874 13905 1906
rect 13873 1806 13905 1838
rect 13873 1738 13905 1770
rect 13873 1670 13905 1702
rect 13873 1602 13905 1634
rect 13873 1534 13905 1566
rect 14175 2350 14207 2382
rect 14175 2282 14207 2314
rect 14175 2214 14207 2246
rect 14175 2146 14207 2178
rect 14175 2078 14207 2110
rect 14175 2010 14207 2042
rect 14175 1942 14207 1974
rect 14175 1874 14207 1906
rect 14175 1806 14207 1838
rect 14175 1738 14207 1770
rect 14175 1670 14207 1702
rect 14175 1602 14207 1634
rect 14175 1534 14207 1566
rect 14477 2350 14509 2382
rect 14477 2282 14509 2314
rect 14477 2214 14509 2246
rect 14477 2146 14509 2178
rect 14477 2078 14509 2110
rect 14477 2010 14509 2042
rect 14477 1942 14509 1974
rect 14477 1874 14509 1906
rect 14477 1806 14509 1838
rect 14477 1738 14509 1770
rect 14477 1670 14509 1702
rect 14477 1602 14509 1634
rect 14477 1534 14509 1566
rect 1491 1382 1523 1414
rect 1491 1314 1523 1346
rect 1491 1246 1523 1278
rect 1491 1178 1523 1210
rect 1491 1110 1523 1142
rect 1491 1042 1523 1074
rect 1491 974 1523 1006
rect 1491 906 1523 938
rect 1491 838 1523 870
rect 1491 770 1523 802
rect 1491 702 1523 734
rect 1491 634 1523 666
rect 1491 566 1523 598
rect 1793 1382 1825 1414
rect 1793 1314 1825 1346
rect 1793 1246 1825 1278
rect 1793 1178 1825 1210
rect 1793 1110 1825 1142
rect 1793 1042 1825 1074
rect 1793 974 1825 1006
rect 1793 906 1825 938
rect 1793 838 1825 870
rect 1793 770 1825 802
rect 1793 702 1825 734
rect 1793 634 1825 666
rect 1793 566 1825 598
rect 2095 1382 2127 1414
rect 2095 1314 2127 1346
rect 2095 1246 2127 1278
rect 2095 1178 2127 1210
rect 2095 1110 2127 1142
rect 2095 1042 2127 1074
rect 2095 974 2127 1006
rect 2095 906 2127 938
rect 2095 838 2127 870
rect 2095 770 2127 802
rect 2095 702 2127 734
rect 2095 634 2127 666
rect 2095 566 2127 598
rect 2397 1382 2429 1414
rect 2397 1314 2429 1346
rect 2397 1246 2429 1278
rect 2397 1178 2429 1210
rect 2397 1110 2429 1142
rect 2397 1042 2429 1074
rect 2397 974 2429 1006
rect 2397 906 2429 938
rect 2397 838 2429 870
rect 2397 770 2429 802
rect 2397 702 2429 734
rect 2397 634 2429 666
rect 2397 566 2429 598
rect 2699 1382 2731 1414
rect 2699 1314 2731 1346
rect 2699 1246 2731 1278
rect 2699 1178 2731 1210
rect 2699 1110 2731 1142
rect 2699 1042 2731 1074
rect 2699 974 2731 1006
rect 2699 906 2731 938
rect 2699 838 2731 870
rect 2699 770 2731 802
rect 2699 702 2731 734
rect 2699 634 2731 666
rect 2699 566 2731 598
rect 3001 1382 3033 1414
rect 3001 1314 3033 1346
rect 3001 1246 3033 1278
rect 3001 1178 3033 1210
rect 3001 1110 3033 1142
rect 3001 1042 3033 1074
rect 3001 974 3033 1006
rect 3001 906 3033 938
rect 3001 838 3033 870
rect 3001 770 3033 802
rect 3001 702 3033 734
rect 3001 634 3033 666
rect 3001 566 3033 598
rect 3303 1382 3335 1414
rect 3303 1314 3335 1346
rect 3303 1246 3335 1278
rect 3303 1178 3335 1210
rect 3303 1110 3335 1142
rect 3303 1042 3335 1074
rect 3303 974 3335 1006
rect 3303 906 3335 938
rect 3303 838 3335 870
rect 3303 770 3335 802
rect 3303 702 3335 734
rect 3303 634 3335 666
rect 3303 566 3335 598
rect 3605 1382 3637 1414
rect 3605 1314 3637 1346
rect 3605 1246 3637 1278
rect 3605 1178 3637 1210
rect 3605 1110 3637 1142
rect 3605 1042 3637 1074
rect 3605 974 3637 1006
rect 3605 906 3637 938
rect 3605 838 3637 870
rect 3605 770 3637 802
rect 3605 702 3637 734
rect 3605 634 3637 666
rect 3605 566 3637 598
rect 3907 1382 3939 1414
rect 3907 1314 3939 1346
rect 3907 1246 3939 1278
rect 3907 1178 3939 1210
rect 3907 1110 3939 1142
rect 3907 1042 3939 1074
rect 3907 974 3939 1006
rect 3907 906 3939 938
rect 3907 838 3939 870
rect 3907 770 3939 802
rect 3907 702 3939 734
rect 3907 634 3939 666
rect 3907 566 3939 598
rect 4209 1382 4241 1414
rect 4209 1314 4241 1346
rect 4209 1246 4241 1278
rect 4209 1178 4241 1210
rect 4209 1110 4241 1142
rect 4209 1042 4241 1074
rect 4209 974 4241 1006
rect 4209 906 4241 938
rect 4209 838 4241 870
rect 4209 770 4241 802
rect 4209 702 4241 734
rect 4209 634 4241 666
rect 4209 566 4241 598
rect 4511 1382 4543 1414
rect 4511 1314 4543 1346
rect 4511 1246 4543 1278
rect 4511 1178 4543 1210
rect 4511 1110 4543 1142
rect 4511 1042 4543 1074
rect 4511 974 4543 1006
rect 4511 906 4543 938
rect 4511 838 4543 870
rect 4511 770 4543 802
rect 4511 702 4543 734
rect 4511 634 4543 666
rect 4511 566 4543 598
rect 4813 1382 4845 1414
rect 4813 1314 4845 1346
rect 4813 1246 4845 1278
rect 4813 1178 4845 1210
rect 4813 1110 4845 1142
rect 4813 1042 4845 1074
rect 4813 974 4845 1006
rect 4813 906 4845 938
rect 4813 838 4845 870
rect 4813 770 4845 802
rect 4813 702 4845 734
rect 4813 634 4845 666
rect 4813 566 4845 598
rect 5115 1382 5147 1414
rect 5115 1314 5147 1346
rect 5115 1246 5147 1278
rect 5115 1178 5147 1210
rect 5115 1110 5147 1142
rect 5115 1042 5147 1074
rect 5115 974 5147 1006
rect 5115 906 5147 938
rect 5115 838 5147 870
rect 5115 770 5147 802
rect 5115 702 5147 734
rect 5115 634 5147 666
rect 5115 566 5147 598
rect 5417 1382 5449 1414
rect 5417 1314 5449 1346
rect 5417 1246 5449 1278
rect 5417 1178 5449 1210
rect 5417 1110 5449 1142
rect 5417 1042 5449 1074
rect 5417 974 5449 1006
rect 5417 906 5449 938
rect 5417 838 5449 870
rect 5417 770 5449 802
rect 5417 702 5449 734
rect 5417 634 5449 666
rect 5417 566 5449 598
rect 5719 1382 5751 1414
rect 5719 1314 5751 1346
rect 5719 1246 5751 1278
rect 5719 1178 5751 1210
rect 5719 1110 5751 1142
rect 5719 1042 5751 1074
rect 5719 974 5751 1006
rect 5719 906 5751 938
rect 5719 838 5751 870
rect 5719 770 5751 802
rect 5719 702 5751 734
rect 5719 634 5751 666
rect 5719 566 5751 598
rect 6021 1382 6053 1414
rect 6021 1314 6053 1346
rect 6021 1246 6053 1278
rect 6021 1178 6053 1210
rect 6021 1110 6053 1142
rect 6021 1042 6053 1074
rect 6021 974 6053 1006
rect 6021 906 6053 938
rect 6021 838 6053 870
rect 6021 770 6053 802
rect 6021 702 6053 734
rect 6021 634 6053 666
rect 6021 566 6053 598
rect 6323 1382 6355 1414
rect 6323 1314 6355 1346
rect 6323 1246 6355 1278
rect 6323 1178 6355 1210
rect 6323 1110 6355 1142
rect 6323 1042 6355 1074
rect 6323 974 6355 1006
rect 6323 906 6355 938
rect 6323 838 6355 870
rect 6323 770 6355 802
rect 6323 702 6355 734
rect 6323 634 6355 666
rect 6323 566 6355 598
rect 6625 1382 6657 1414
rect 6625 1314 6657 1346
rect 6625 1246 6657 1278
rect 6625 1178 6657 1210
rect 6625 1110 6657 1142
rect 6625 1042 6657 1074
rect 6625 974 6657 1006
rect 6625 906 6657 938
rect 6625 838 6657 870
rect 6625 770 6657 802
rect 6625 702 6657 734
rect 6625 634 6657 666
rect 6625 566 6657 598
rect 6927 1382 6959 1414
rect 6927 1314 6959 1346
rect 6927 1246 6959 1278
rect 6927 1178 6959 1210
rect 6927 1110 6959 1142
rect 6927 1042 6959 1074
rect 6927 974 6959 1006
rect 6927 906 6959 938
rect 6927 838 6959 870
rect 6927 770 6959 802
rect 6927 702 6959 734
rect 6927 634 6959 666
rect 6927 566 6959 598
rect 7229 1382 7261 1414
rect 7229 1314 7261 1346
rect 7229 1246 7261 1278
rect 7229 1178 7261 1210
rect 7229 1110 7261 1142
rect 7229 1042 7261 1074
rect 7229 974 7261 1006
rect 7229 906 7261 938
rect 7229 838 7261 870
rect 7229 770 7261 802
rect 7229 702 7261 734
rect 7229 634 7261 666
rect 7229 566 7261 598
rect 7531 1382 7563 1414
rect 7531 1314 7563 1346
rect 7531 1246 7563 1278
rect 7531 1178 7563 1210
rect 7531 1110 7563 1142
rect 7531 1042 7563 1074
rect 7531 974 7563 1006
rect 7531 906 7563 938
rect 7531 838 7563 870
rect 7531 770 7563 802
rect 7531 702 7563 734
rect 7531 634 7563 666
rect 7531 566 7563 598
rect 7833 1382 7865 1414
rect 7833 1314 7865 1346
rect 7833 1246 7865 1278
rect 7833 1178 7865 1210
rect 7833 1110 7865 1142
rect 7833 1042 7865 1074
rect 7833 974 7865 1006
rect 7833 906 7865 938
rect 7833 838 7865 870
rect 7833 770 7865 802
rect 7833 702 7865 734
rect 7833 634 7865 666
rect 7833 566 7865 598
rect 8135 1382 8167 1414
rect 8135 1314 8167 1346
rect 8135 1246 8167 1278
rect 8135 1178 8167 1210
rect 8135 1110 8167 1142
rect 8135 1042 8167 1074
rect 8135 974 8167 1006
rect 8135 906 8167 938
rect 8135 838 8167 870
rect 8135 770 8167 802
rect 8135 702 8167 734
rect 8135 634 8167 666
rect 8135 566 8167 598
rect 8437 1382 8469 1414
rect 8437 1314 8469 1346
rect 8437 1246 8469 1278
rect 8437 1178 8469 1210
rect 8437 1110 8469 1142
rect 8437 1042 8469 1074
rect 8437 974 8469 1006
rect 8437 906 8469 938
rect 8437 838 8469 870
rect 8437 770 8469 802
rect 8437 702 8469 734
rect 8437 634 8469 666
rect 8437 566 8469 598
rect 8739 1382 8771 1414
rect 8739 1314 8771 1346
rect 8739 1246 8771 1278
rect 8739 1178 8771 1210
rect 8739 1110 8771 1142
rect 8739 1042 8771 1074
rect 8739 974 8771 1006
rect 8739 906 8771 938
rect 8739 838 8771 870
rect 8739 770 8771 802
rect 8739 702 8771 734
rect 8739 634 8771 666
rect 8739 566 8771 598
rect 9041 1382 9073 1414
rect 9041 1314 9073 1346
rect 9041 1246 9073 1278
rect 9041 1178 9073 1210
rect 9041 1110 9073 1142
rect 9041 1042 9073 1074
rect 9041 974 9073 1006
rect 9041 906 9073 938
rect 9041 838 9073 870
rect 9041 770 9073 802
rect 9041 702 9073 734
rect 9041 634 9073 666
rect 9041 566 9073 598
rect 9343 1382 9375 1414
rect 9343 1314 9375 1346
rect 9343 1246 9375 1278
rect 9343 1178 9375 1210
rect 9343 1110 9375 1142
rect 9343 1042 9375 1074
rect 9343 974 9375 1006
rect 9343 906 9375 938
rect 9343 838 9375 870
rect 9343 770 9375 802
rect 9343 702 9375 734
rect 9343 634 9375 666
rect 9343 566 9375 598
rect 9645 1382 9677 1414
rect 9645 1314 9677 1346
rect 9645 1246 9677 1278
rect 9645 1178 9677 1210
rect 9645 1110 9677 1142
rect 9645 1042 9677 1074
rect 9645 974 9677 1006
rect 9645 906 9677 938
rect 9645 838 9677 870
rect 9645 770 9677 802
rect 9645 702 9677 734
rect 9645 634 9677 666
rect 9645 566 9677 598
rect 9947 1382 9979 1414
rect 9947 1314 9979 1346
rect 9947 1246 9979 1278
rect 9947 1178 9979 1210
rect 9947 1110 9979 1142
rect 9947 1042 9979 1074
rect 9947 974 9979 1006
rect 9947 906 9979 938
rect 9947 838 9979 870
rect 9947 770 9979 802
rect 9947 702 9979 734
rect 9947 634 9979 666
rect 9947 566 9979 598
rect 10249 1382 10281 1414
rect 10249 1314 10281 1346
rect 10249 1246 10281 1278
rect 10249 1178 10281 1210
rect 10249 1110 10281 1142
rect 10249 1042 10281 1074
rect 10249 974 10281 1006
rect 10249 906 10281 938
rect 10249 838 10281 870
rect 10249 770 10281 802
rect 10249 702 10281 734
rect 10249 634 10281 666
rect 10249 566 10281 598
rect 10551 1382 10583 1414
rect 10551 1314 10583 1346
rect 10551 1246 10583 1278
rect 10551 1178 10583 1210
rect 10551 1110 10583 1142
rect 10551 1042 10583 1074
rect 10551 974 10583 1006
rect 10551 906 10583 938
rect 10551 838 10583 870
rect 10551 770 10583 802
rect 10551 702 10583 734
rect 10551 634 10583 666
rect 10551 566 10583 598
rect 10853 1382 10885 1414
rect 10853 1314 10885 1346
rect 10853 1246 10885 1278
rect 10853 1178 10885 1210
rect 10853 1110 10885 1142
rect 10853 1042 10885 1074
rect 10853 974 10885 1006
rect 10853 906 10885 938
rect 10853 838 10885 870
rect 10853 770 10885 802
rect 10853 702 10885 734
rect 10853 634 10885 666
rect 10853 566 10885 598
rect 11155 1382 11187 1414
rect 11155 1314 11187 1346
rect 11155 1246 11187 1278
rect 11155 1178 11187 1210
rect 11155 1110 11187 1142
rect 11155 1042 11187 1074
rect 11155 974 11187 1006
rect 11155 906 11187 938
rect 11155 838 11187 870
rect 11155 770 11187 802
rect 11155 702 11187 734
rect 11155 634 11187 666
rect 11155 566 11187 598
rect 11457 1382 11489 1414
rect 11457 1314 11489 1346
rect 11457 1246 11489 1278
rect 11457 1178 11489 1210
rect 11457 1110 11489 1142
rect 11457 1042 11489 1074
rect 11457 974 11489 1006
rect 11457 906 11489 938
rect 11457 838 11489 870
rect 11457 770 11489 802
rect 11457 702 11489 734
rect 11457 634 11489 666
rect 11457 566 11489 598
rect 11759 1382 11791 1414
rect 11759 1314 11791 1346
rect 11759 1246 11791 1278
rect 11759 1178 11791 1210
rect 11759 1110 11791 1142
rect 11759 1042 11791 1074
rect 11759 974 11791 1006
rect 11759 906 11791 938
rect 11759 838 11791 870
rect 11759 770 11791 802
rect 11759 702 11791 734
rect 11759 634 11791 666
rect 11759 566 11791 598
rect 12061 1382 12093 1414
rect 12061 1314 12093 1346
rect 12061 1246 12093 1278
rect 12061 1178 12093 1210
rect 12061 1110 12093 1142
rect 12061 1042 12093 1074
rect 12061 974 12093 1006
rect 12061 906 12093 938
rect 12061 838 12093 870
rect 12061 770 12093 802
rect 12061 702 12093 734
rect 12061 634 12093 666
rect 12061 566 12093 598
rect 12363 1382 12395 1414
rect 12363 1314 12395 1346
rect 12363 1246 12395 1278
rect 12363 1178 12395 1210
rect 12363 1110 12395 1142
rect 12363 1042 12395 1074
rect 12363 974 12395 1006
rect 12363 906 12395 938
rect 12363 838 12395 870
rect 12363 770 12395 802
rect 12363 702 12395 734
rect 12363 634 12395 666
rect 12363 566 12395 598
rect 12665 1382 12697 1414
rect 12665 1314 12697 1346
rect 12665 1246 12697 1278
rect 12665 1178 12697 1210
rect 12665 1110 12697 1142
rect 12665 1042 12697 1074
rect 12665 974 12697 1006
rect 12665 906 12697 938
rect 12665 838 12697 870
rect 12665 770 12697 802
rect 12665 702 12697 734
rect 12665 634 12697 666
rect 12665 566 12697 598
rect 12967 1382 12999 1414
rect 12967 1314 12999 1346
rect 12967 1246 12999 1278
rect 12967 1178 12999 1210
rect 12967 1110 12999 1142
rect 12967 1042 12999 1074
rect 12967 974 12999 1006
rect 12967 906 12999 938
rect 12967 838 12999 870
rect 12967 770 12999 802
rect 12967 702 12999 734
rect 12967 634 12999 666
rect 12967 566 12999 598
rect 13269 1382 13301 1414
rect 13269 1314 13301 1346
rect 13269 1246 13301 1278
rect 13269 1178 13301 1210
rect 13269 1110 13301 1142
rect 13269 1042 13301 1074
rect 13269 974 13301 1006
rect 13269 906 13301 938
rect 13269 838 13301 870
rect 13269 770 13301 802
rect 13269 702 13301 734
rect 13269 634 13301 666
rect 13269 566 13301 598
rect 13571 1382 13603 1414
rect 13571 1314 13603 1346
rect 13571 1246 13603 1278
rect 13571 1178 13603 1210
rect 13571 1110 13603 1142
rect 13571 1042 13603 1074
rect 13571 974 13603 1006
rect 13571 906 13603 938
rect 13571 838 13603 870
rect 13571 770 13603 802
rect 13571 702 13603 734
rect 13571 634 13603 666
rect 13571 566 13603 598
rect 13873 1382 13905 1414
rect 13873 1314 13905 1346
rect 13873 1246 13905 1278
rect 13873 1178 13905 1210
rect 13873 1110 13905 1142
rect 13873 1042 13905 1074
rect 13873 974 13905 1006
rect 13873 906 13905 938
rect 13873 838 13905 870
rect 13873 770 13905 802
rect 13873 702 13905 734
rect 13873 634 13905 666
rect 13873 566 13905 598
rect 14175 1382 14207 1414
rect 14175 1314 14207 1346
rect 14175 1246 14207 1278
rect 14175 1178 14207 1210
rect 14175 1110 14207 1142
rect 14175 1042 14207 1074
rect 14175 974 14207 1006
rect 14175 906 14207 938
rect 14175 838 14207 870
rect 14175 770 14207 802
rect 14175 702 14207 734
rect 14175 634 14207 666
rect 14175 566 14207 598
rect 14477 1382 14509 1414
rect 14477 1314 14509 1346
rect 14477 1246 14509 1278
rect 14477 1178 14509 1210
rect 14477 1110 14509 1142
rect 14477 1042 14509 1074
rect 14477 974 14509 1006
rect 14477 906 14509 938
rect 14477 838 14509 870
rect 14477 770 14509 802
rect 14477 702 14509 734
rect 14477 634 14509 666
rect 14477 566 14509 598
<< psubdiff >>
rect 360 4506 15640 4524
rect 360 4474 402 4506
rect 434 4474 470 4506
rect 502 4474 538 4506
rect 570 4474 606 4506
rect 638 4474 674 4506
rect 706 4474 742 4506
rect 774 4474 810 4506
rect 842 4474 878 4506
rect 910 4474 946 4506
rect 978 4474 1014 4506
rect 1046 4474 1082 4506
rect 1114 4474 1150 4506
rect 1182 4474 1218 4506
rect 1250 4474 1286 4506
rect 1318 4474 1354 4506
rect 1386 4474 1422 4506
rect 1454 4474 1490 4506
rect 1522 4474 1558 4506
rect 1590 4474 1626 4506
rect 1658 4474 1694 4506
rect 1726 4474 1762 4506
rect 1794 4474 1830 4506
rect 1862 4474 1898 4506
rect 1930 4474 1966 4506
rect 1998 4474 2034 4506
rect 2066 4474 2102 4506
rect 2134 4474 2170 4506
rect 2202 4474 2238 4506
rect 2270 4474 2306 4506
rect 2338 4474 2374 4506
rect 2406 4474 2442 4506
rect 2474 4474 2510 4506
rect 2542 4474 2578 4506
rect 2610 4474 2646 4506
rect 2678 4474 2714 4506
rect 2746 4474 2782 4506
rect 2814 4474 2850 4506
rect 2882 4474 2918 4506
rect 2950 4474 2986 4506
rect 3018 4474 3054 4506
rect 3086 4474 3122 4506
rect 3154 4474 3190 4506
rect 3222 4474 3258 4506
rect 3290 4474 3326 4506
rect 3358 4474 3394 4506
rect 3426 4474 3462 4506
rect 3494 4474 3530 4506
rect 3562 4474 3598 4506
rect 3630 4474 3666 4506
rect 3698 4474 3734 4506
rect 3766 4474 3802 4506
rect 3834 4474 3870 4506
rect 3902 4474 3938 4506
rect 3970 4474 4006 4506
rect 4038 4474 4074 4506
rect 4106 4474 4142 4506
rect 4174 4474 4210 4506
rect 4242 4474 4278 4506
rect 4310 4474 4346 4506
rect 4378 4474 4414 4506
rect 4446 4474 4482 4506
rect 4514 4474 4550 4506
rect 4582 4474 4618 4506
rect 4650 4474 4686 4506
rect 4718 4474 4754 4506
rect 4786 4474 4822 4506
rect 4854 4474 4890 4506
rect 4922 4474 4958 4506
rect 4990 4474 5026 4506
rect 5058 4474 5094 4506
rect 5126 4474 5162 4506
rect 5194 4474 5230 4506
rect 5262 4474 5298 4506
rect 5330 4474 5366 4506
rect 5398 4474 5434 4506
rect 5466 4474 5502 4506
rect 5534 4474 5570 4506
rect 5602 4474 5638 4506
rect 5670 4474 5706 4506
rect 5738 4474 5774 4506
rect 5806 4474 5842 4506
rect 5874 4474 5910 4506
rect 5942 4474 5978 4506
rect 6010 4474 6046 4506
rect 6078 4474 6114 4506
rect 6146 4474 6182 4506
rect 6214 4474 6250 4506
rect 6282 4474 6318 4506
rect 6350 4474 6386 4506
rect 6418 4474 6454 4506
rect 6486 4474 6522 4506
rect 6554 4474 6590 4506
rect 6622 4474 6658 4506
rect 6690 4474 6726 4506
rect 6758 4474 6794 4506
rect 6826 4474 6862 4506
rect 6894 4474 6930 4506
rect 6962 4474 6998 4506
rect 7030 4474 7066 4506
rect 7098 4474 7134 4506
rect 7166 4474 7202 4506
rect 7234 4474 7270 4506
rect 7302 4474 7338 4506
rect 7370 4474 7406 4506
rect 7438 4474 7474 4506
rect 7506 4474 7542 4506
rect 7574 4474 7610 4506
rect 7642 4474 7678 4506
rect 7710 4474 7746 4506
rect 7778 4474 7814 4506
rect 7846 4474 7882 4506
rect 7914 4474 7950 4506
rect 7982 4474 8018 4506
rect 8050 4474 8086 4506
rect 8118 4474 8154 4506
rect 8186 4474 8222 4506
rect 8254 4474 8290 4506
rect 8322 4474 8358 4506
rect 8390 4474 8426 4506
rect 8458 4474 8494 4506
rect 8526 4474 8562 4506
rect 8594 4474 8630 4506
rect 8662 4474 8698 4506
rect 8730 4474 8766 4506
rect 8798 4474 8834 4506
rect 8866 4474 8902 4506
rect 8934 4474 8970 4506
rect 9002 4474 9038 4506
rect 9070 4474 9106 4506
rect 9138 4474 9174 4506
rect 9206 4474 9242 4506
rect 9274 4474 9310 4506
rect 9342 4474 9378 4506
rect 9410 4474 9446 4506
rect 9478 4474 9514 4506
rect 9546 4474 9582 4506
rect 9614 4474 9650 4506
rect 9682 4474 9718 4506
rect 9750 4474 9786 4506
rect 9818 4474 9854 4506
rect 9886 4474 9922 4506
rect 9954 4474 9990 4506
rect 10022 4474 10058 4506
rect 10090 4474 10126 4506
rect 10158 4474 10194 4506
rect 10226 4474 10262 4506
rect 10294 4474 10330 4506
rect 10362 4474 10398 4506
rect 10430 4474 10466 4506
rect 10498 4474 10534 4506
rect 10566 4474 10602 4506
rect 10634 4474 10670 4506
rect 10702 4474 10738 4506
rect 10770 4474 10806 4506
rect 10838 4474 10874 4506
rect 10906 4474 10942 4506
rect 10974 4474 11010 4506
rect 11042 4474 11078 4506
rect 11110 4474 11146 4506
rect 11178 4474 11214 4506
rect 11246 4474 11282 4506
rect 11314 4474 11350 4506
rect 11382 4474 11418 4506
rect 11450 4474 11486 4506
rect 11518 4474 11554 4506
rect 11586 4474 11622 4506
rect 11654 4474 11690 4506
rect 11722 4474 11758 4506
rect 11790 4474 11826 4506
rect 11858 4474 11894 4506
rect 11926 4474 11962 4506
rect 11994 4474 12030 4506
rect 12062 4474 12098 4506
rect 12130 4474 12166 4506
rect 12198 4474 12234 4506
rect 12266 4474 12302 4506
rect 12334 4474 12370 4506
rect 12402 4474 12438 4506
rect 12470 4474 12506 4506
rect 12538 4474 12574 4506
rect 12606 4474 12642 4506
rect 12674 4474 12710 4506
rect 12742 4474 12778 4506
rect 12810 4474 12846 4506
rect 12878 4474 12914 4506
rect 12946 4474 12982 4506
rect 13014 4474 13050 4506
rect 13082 4474 13118 4506
rect 13150 4474 13186 4506
rect 13218 4474 13254 4506
rect 13286 4474 13322 4506
rect 13354 4474 13390 4506
rect 13422 4474 13458 4506
rect 13490 4474 13526 4506
rect 13558 4474 13594 4506
rect 13626 4474 13662 4506
rect 13694 4474 13730 4506
rect 13762 4474 13798 4506
rect 13830 4474 13866 4506
rect 13898 4474 13934 4506
rect 13966 4474 14002 4506
rect 14034 4474 14070 4506
rect 14102 4474 14138 4506
rect 14170 4474 14206 4506
rect 14238 4474 14274 4506
rect 14306 4474 14342 4506
rect 14374 4474 14410 4506
rect 14442 4474 14478 4506
rect 14510 4474 14546 4506
rect 14578 4474 14614 4506
rect 14646 4474 14682 4506
rect 14714 4474 14750 4506
rect 14782 4474 14818 4506
rect 14850 4474 14886 4506
rect 14918 4474 14954 4506
rect 14986 4474 15022 4506
rect 15054 4474 15090 4506
rect 15122 4474 15158 4506
rect 15190 4474 15226 4506
rect 15258 4474 15294 4506
rect 15326 4474 15362 4506
rect 15394 4474 15430 4506
rect 15462 4474 15498 4506
rect 15530 4474 15566 4506
rect 15598 4474 15640 4506
rect 360 4456 15640 4474
rect 360 4396 428 4456
rect 360 4364 378 4396
rect 410 4364 428 4396
rect 360 4328 428 4364
rect 15572 4396 15640 4456
rect 15572 4364 15590 4396
rect 15622 4364 15640 4396
rect 360 4296 378 4328
rect 410 4296 428 4328
rect 360 4260 428 4296
rect 360 4228 378 4260
rect 410 4228 428 4260
rect 360 4192 428 4228
rect 360 4160 378 4192
rect 410 4160 428 4192
rect 360 4124 428 4160
rect 360 4092 378 4124
rect 410 4092 428 4124
rect 360 4056 428 4092
rect 360 4024 378 4056
rect 410 4024 428 4056
rect 360 3988 428 4024
rect 360 3956 378 3988
rect 410 3956 428 3988
rect 360 3920 428 3956
rect 360 3888 378 3920
rect 410 3888 428 3920
rect 360 3852 428 3888
rect 360 3820 378 3852
rect 410 3820 428 3852
rect 360 3784 428 3820
rect 360 3752 378 3784
rect 410 3752 428 3784
rect 360 3716 428 3752
rect 360 3684 378 3716
rect 410 3684 428 3716
rect 360 3648 428 3684
rect 360 3616 378 3648
rect 410 3616 428 3648
rect 360 3580 428 3616
rect 360 3548 378 3580
rect 410 3548 428 3580
rect 360 3512 428 3548
rect 360 3480 378 3512
rect 410 3480 428 3512
rect 360 3444 428 3480
rect 15572 4328 15640 4364
rect 15572 4296 15590 4328
rect 15622 4296 15640 4328
rect 15572 4260 15640 4296
rect 15572 4228 15590 4260
rect 15622 4228 15640 4260
rect 15572 4192 15640 4228
rect 15572 4160 15590 4192
rect 15622 4160 15640 4192
rect 15572 4124 15640 4160
rect 15572 4092 15590 4124
rect 15622 4092 15640 4124
rect 15572 4056 15640 4092
rect 15572 4024 15590 4056
rect 15622 4024 15640 4056
rect 15572 3988 15640 4024
rect 15572 3956 15590 3988
rect 15622 3956 15640 3988
rect 15572 3920 15640 3956
rect 15572 3888 15590 3920
rect 15622 3888 15640 3920
rect 15572 3852 15640 3888
rect 15572 3820 15590 3852
rect 15622 3820 15640 3852
rect 15572 3784 15640 3820
rect 15572 3752 15590 3784
rect 15622 3752 15640 3784
rect 15572 3716 15640 3752
rect 15572 3684 15590 3716
rect 15622 3684 15640 3716
rect 15572 3648 15640 3684
rect 15572 3616 15590 3648
rect 15622 3616 15640 3648
rect 15572 3580 15640 3616
rect 15572 3548 15590 3580
rect 15622 3548 15640 3580
rect 15572 3512 15640 3548
rect 15572 3480 15590 3512
rect 15622 3480 15640 3512
rect 360 3412 378 3444
rect 410 3412 428 3444
rect 360 3376 428 3412
rect 360 3344 378 3376
rect 410 3344 428 3376
rect 15572 3444 15640 3480
rect 15572 3412 15590 3444
rect 15622 3412 15640 3444
rect 15572 3376 15640 3412
rect 360 3308 428 3344
rect 360 3276 378 3308
rect 410 3276 428 3308
rect 360 3240 428 3276
rect 360 3208 378 3240
rect 410 3208 428 3240
rect 360 3172 428 3208
rect 360 3140 378 3172
rect 410 3140 428 3172
rect 360 3104 428 3140
rect 360 3072 378 3104
rect 410 3072 428 3104
rect 360 3036 428 3072
rect 360 3004 378 3036
rect 410 3004 428 3036
rect 360 2968 428 3004
rect 360 2936 378 2968
rect 410 2936 428 2968
rect 360 2900 428 2936
rect 360 2868 378 2900
rect 410 2868 428 2900
rect 360 2832 428 2868
rect 360 2800 378 2832
rect 410 2800 428 2832
rect 360 2764 428 2800
rect 360 2732 378 2764
rect 410 2732 428 2764
rect 360 2696 428 2732
rect 360 2664 378 2696
rect 410 2664 428 2696
rect 360 2628 428 2664
rect 360 2596 378 2628
rect 410 2596 428 2628
rect 360 2560 428 2596
rect 360 2528 378 2560
rect 410 2528 428 2560
rect 360 2492 428 2528
rect 360 2460 378 2492
rect 410 2460 428 2492
rect 15572 3344 15590 3376
rect 15622 3344 15640 3376
rect 15572 3308 15640 3344
rect 15572 3276 15590 3308
rect 15622 3276 15640 3308
rect 15572 3240 15640 3276
rect 15572 3208 15590 3240
rect 15622 3208 15640 3240
rect 15572 3172 15640 3208
rect 15572 3140 15590 3172
rect 15622 3140 15640 3172
rect 15572 3104 15640 3140
rect 15572 3072 15590 3104
rect 15622 3072 15640 3104
rect 15572 3036 15640 3072
rect 15572 3004 15590 3036
rect 15622 3004 15640 3036
rect 15572 2968 15640 3004
rect 15572 2936 15590 2968
rect 15622 2936 15640 2968
rect 15572 2900 15640 2936
rect 15572 2868 15590 2900
rect 15622 2868 15640 2900
rect 15572 2832 15640 2868
rect 15572 2800 15590 2832
rect 15622 2800 15640 2832
rect 15572 2764 15640 2800
rect 15572 2732 15590 2764
rect 15622 2732 15640 2764
rect 15572 2696 15640 2732
rect 15572 2664 15590 2696
rect 15622 2664 15640 2696
rect 15572 2628 15640 2664
rect 15572 2596 15590 2628
rect 15622 2596 15640 2628
rect 15572 2560 15640 2596
rect 15572 2528 15590 2560
rect 15622 2528 15640 2560
rect 15572 2492 15640 2528
rect 360 2424 428 2460
rect 360 2392 378 2424
rect 410 2392 428 2424
rect 15572 2460 15590 2492
rect 15622 2460 15640 2492
rect 15572 2424 15640 2460
rect 360 2356 428 2392
rect 360 2324 378 2356
rect 410 2324 428 2356
rect 360 2288 428 2324
rect 360 2256 378 2288
rect 410 2256 428 2288
rect 360 2220 428 2256
rect 360 2188 378 2220
rect 410 2188 428 2220
rect 360 2152 428 2188
rect 360 2120 378 2152
rect 410 2120 428 2152
rect 360 2084 428 2120
rect 360 2052 378 2084
rect 410 2052 428 2084
rect 360 2016 428 2052
rect 360 1984 378 2016
rect 410 1984 428 2016
rect 360 1948 428 1984
rect 360 1916 378 1948
rect 410 1916 428 1948
rect 360 1880 428 1916
rect 360 1848 378 1880
rect 410 1848 428 1880
rect 360 1812 428 1848
rect 360 1780 378 1812
rect 410 1780 428 1812
rect 360 1744 428 1780
rect 360 1712 378 1744
rect 410 1712 428 1744
rect 360 1676 428 1712
rect 360 1644 378 1676
rect 410 1644 428 1676
rect 360 1608 428 1644
rect 360 1576 378 1608
rect 410 1576 428 1608
rect 360 1540 428 1576
rect 360 1508 378 1540
rect 410 1508 428 1540
rect 15572 2392 15590 2424
rect 15622 2392 15640 2424
rect 15572 2356 15640 2392
rect 15572 2324 15590 2356
rect 15622 2324 15640 2356
rect 15572 2288 15640 2324
rect 15572 2256 15590 2288
rect 15622 2256 15640 2288
rect 15572 2220 15640 2256
rect 15572 2188 15590 2220
rect 15622 2188 15640 2220
rect 15572 2152 15640 2188
rect 15572 2120 15590 2152
rect 15622 2120 15640 2152
rect 15572 2084 15640 2120
rect 15572 2052 15590 2084
rect 15622 2052 15640 2084
rect 15572 2016 15640 2052
rect 15572 1984 15590 2016
rect 15622 1984 15640 2016
rect 15572 1948 15640 1984
rect 15572 1916 15590 1948
rect 15622 1916 15640 1948
rect 15572 1880 15640 1916
rect 15572 1848 15590 1880
rect 15622 1848 15640 1880
rect 15572 1812 15640 1848
rect 15572 1780 15590 1812
rect 15622 1780 15640 1812
rect 15572 1744 15640 1780
rect 15572 1712 15590 1744
rect 15622 1712 15640 1744
rect 15572 1676 15640 1712
rect 15572 1644 15590 1676
rect 15622 1644 15640 1676
rect 15572 1608 15640 1644
rect 15572 1576 15590 1608
rect 15622 1576 15640 1608
rect 15572 1540 15640 1576
rect 360 1472 428 1508
rect 360 1440 378 1472
rect 410 1440 428 1472
rect 360 1404 428 1440
rect 15572 1508 15590 1540
rect 15622 1508 15640 1540
rect 15572 1472 15640 1508
rect 15572 1440 15590 1472
rect 15622 1440 15640 1472
rect 360 1372 378 1404
rect 410 1372 428 1404
rect 360 1336 428 1372
rect 360 1304 378 1336
rect 410 1304 428 1336
rect 360 1268 428 1304
rect 360 1236 378 1268
rect 410 1236 428 1268
rect 360 1200 428 1236
rect 360 1168 378 1200
rect 410 1168 428 1200
rect 360 1132 428 1168
rect 360 1100 378 1132
rect 410 1100 428 1132
rect 360 1064 428 1100
rect 360 1032 378 1064
rect 410 1032 428 1064
rect 360 996 428 1032
rect 360 964 378 996
rect 410 964 428 996
rect 360 928 428 964
rect 360 896 378 928
rect 410 896 428 928
rect 360 860 428 896
rect 360 828 378 860
rect 410 828 428 860
rect 360 792 428 828
rect 360 760 378 792
rect 410 760 428 792
rect 360 724 428 760
rect 360 692 378 724
rect 410 692 428 724
rect 360 656 428 692
rect 360 624 378 656
rect 410 624 428 656
rect 360 588 428 624
rect 360 556 378 588
rect 410 556 428 588
rect 360 520 428 556
rect 15572 1404 15640 1440
rect 15572 1372 15590 1404
rect 15622 1372 15640 1404
rect 15572 1336 15640 1372
rect 15572 1304 15590 1336
rect 15622 1304 15640 1336
rect 15572 1268 15640 1304
rect 15572 1236 15590 1268
rect 15622 1236 15640 1268
rect 15572 1200 15640 1236
rect 15572 1168 15590 1200
rect 15622 1168 15640 1200
rect 15572 1132 15640 1168
rect 15572 1100 15590 1132
rect 15622 1100 15640 1132
rect 15572 1064 15640 1100
rect 15572 1032 15590 1064
rect 15622 1032 15640 1064
rect 15572 996 15640 1032
rect 15572 964 15590 996
rect 15622 964 15640 996
rect 15572 928 15640 964
rect 15572 896 15590 928
rect 15622 896 15640 928
rect 15572 860 15640 896
rect 15572 828 15590 860
rect 15622 828 15640 860
rect 15572 792 15640 828
rect 15572 760 15590 792
rect 15622 760 15640 792
rect 15572 724 15640 760
rect 15572 692 15590 724
rect 15622 692 15640 724
rect 15572 656 15640 692
rect 15572 624 15590 656
rect 15622 624 15640 656
rect 15572 588 15640 624
rect 15572 556 15590 588
rect 15622 556 15640 588
rect 360 488 378 520
rect 410 488 428 520
rect 360 428 428 488
rect 15572 520 15640 556
rect 15572 488 15590 520
rect 15622 488 15640 520
rect 15572 428 15640 488
rect 360 410 15640 428
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 360 15640 378
<< nsubdiff >>
rect 0 4866 16000 4884
rect 0 4834 28 4866
rect 60 4834 96 4866
rect 128 4834 164 4866
rect 196 4834 232 4866
rect 264 4834 300 4866
rect 332 4834 368 4866
rect 400 4834 436 4866
rect 468 4834 504 4866
rect 536 4834 572 4866
rect 604 4834 640 4866
rect 672 4834 708 4866
rect 740 4834 776 4866
rect 808 4834 844 4866
rect 876 4834 912 4866
rect 944 4834 980 4866
rect 1012 4834 1048 4866
rect 1080 4834 1116 4866
rect 1148 4834 1184 4866
rect 1216 4834 1252 4866
rect 1284 4834 1320 4866
rect 1352 4834 1388 4866
rect 1420 4834 1456 4866
rect 1488 4834 1524 4866
rect 1556 4834 1592 4866
rect 1624 4834 1660 4866
rect 1692 4834 1728 4866
rect 1760 4834 1796 4866
rect 1828 4834 1864 4866
rect 1896 4834 1932 4866
rect 1964 4834 2000 4866
rect 2032 4834 2068 4866
rect 2100 4834 2136 4866
rect 2168 4834 2204 4866
rect 2236 4834 2272 4866
rect 2304 4834 2340 4866
rect 2372 4834 2408 4866
rect 2440 4834 2476 4866
rect 2508 4834 2544 4866
rect 2576 4834 2612 4866
rect 2644 4834 2680 4866
rect 2712 4834 2748 4866
rect 2780 4834 2816 4866
rect 2848 4834 2884 4866
rect 2916 4834 2952 4866
rect 2984 4834 3020 4866
rect 3052 4834 3088 4866
rect 3120 4834 3156 4866
rect 3188 4834 3224 4866
rect 3256 4834 3292 4866
rect 3324 4834 3360 4866
rect 3392 4834 3428 4866
rect 3460 4834 3496 4866
rect 3528 4834 3564 4866
rect 3596 4834 3632 4866
rect 3664 4834 3700 4866
rect 3732 4834 3768 4866
rect 3800 4834 3836 4866
rect 3868 4834 3904 4866
rect 3936 4834 3972 4866
rect 4004 4834 4040 4866
rect 4072 4834 4108 4866
rect 4140 4834 4176 4866
rect 4208 4834 4244 4866
rect 4276 4834 4312 4866
rect 4344 4834 4380 4866
rect 4412 4834 4448 4866
rect 4480 4834 4516 4866
rect 4548 4834 4584 4866
rect 4616 4834 4652 4866
rect 4684 4834 4720 4866
rect 4752 4834 4788 4866
rect 4820 4834 4856 4866
rect 4888 4834 4924 4866
rect 4956 4834 4992 4866
rect 5024 4834 5060 4866
rect 5092 4834 5128 4866
rect 5160 4834 5196 4866
rect 5228 4834 5264 4866
rect 5296 4834 5332 4866
rect 5364 4834 5400 4866
rect 5432 4834 5468 4866
rect 5500 4834 5536 4866
rect 5568 4834 5604 4866
rect 5636 4834 5672 4866
rect 5704 4834 5740 4866
rect 5772 4834 5808 4866
rect 5840 4834 5876 4866
rect 5908 4834 5944 4866
rect 5976 4834 6012 4866
rect 6044 4834 6080 4866
rect 6112 4834 6148 4866
rect 6180 4834 6216 4866
rect 6248 4834 6284 4866
rect 6316 4834 6352 4866
rect 6384 4834 6420 4866
rect 6452 4834 6488 4866
rect 6520 4834 6556 4866
rect 6588 4834 6624 4866
rect 6656 4834 6692 4866
rect 6724 4834 6760 4866
rect 6792 4834 6828 4866
rect 6860 4834 6896 4866
rect 6928 4834 6964 4866
rect 6996 4834 7032 4866
rect 7064 4834 7100 4866
rect 7132 4834 7168 4866
rect 7200 4834 7236 4866
rect 7268 4834 7304 4866
rect 7336 4834 7372 4866
rect 7404 4834 7440 4866
rect 7472 4834 7508 4866
rect 7540 4834 7576 4866
rect 7608 4834 7644 4866
rect 7676 4834 7712 4866
rect 7744 4834 7780 4866
rect 7812 4834 7848 4866
rect 7880 4834 7916 4866
rect 7948 4834 7984 4866
rect 8016 4834 8052 4866
rect 8084 4834 8120 4866
rect 8152 4834 8188 4866
rect 8220 4834 8256 4866
rect 8288 4834 8324 4866
rect 8356 4834 8392 4866
rect 8424 4834 8460 4866
rect 8492 4834 8528 4866
rect 8560 4834 8596 4866
rect 8628 4834 8664 4866
rect 8696 4834 8732 4866
rect 8764 4834 8800 4866
rect 8832 4834 8868 4866
rect 8900 4834 8936 4866
rect 8968 4834 9004 4866
rect 9036 4834 9072 4866
rect 9104 4834 9140 4866
rect 9172 4834 9208 4866
rect 9240 4834 9276 4866
rect 9308 4834 9344 4866
rect 9376 4834 9412 4866
rect 9444 4834 9480 4866
rect 9512 4834 9548 4866
rect 9580 4834 9616 4866
rect 9648 4834 9684 4866
rect 9716 4834 9752 4866
rect 9784 4834 9820 4866
rect 9852 4834 9888 4866
rect 9920 4834 9956 4866
rect 9988 4834 10024 4866
rect 10056 4834 10092 4866
rect 10124 4834 10160 4866
rect 10192 4834 10228 4866
rect 10260 4834 10296 4866
rect 10328 4834 10364 4866
rect 10396 4834 10432 4866
rect 10464 4834 10500 4866
rect 10532 4834 10568 4866
rect 10600 4834 10636 4866
rect 10668 4834 10704 4866
rect 10736 4834 10772 4866
rect 10804 4834 10840 4866
rect 10872 4834 10908 4866
rect 10940 4834 10976 4866
rect 11008 4834 11044 4866
rect 11076 4834 11112 4866
rect 11144 4834 11180 4866
rect 11212 4834 11248 4866
rect 11280 4834 11316 4866
rect 11348 4834 11384 4866
rect 11416 4834 11452 4866
rect 11484 4834 11520 4866
rect 11552 4834 11588 4866
rect 11620 4834 11656 4866
rect 11688 4834 11724 4866
rect 11756 4834 11792 4866
rect 11824 4834 11860 4866
rect 11892 4834 11928 4866
rect 11960 4834 11996 4866
rect 12028 4834 12064 4866
rect 12096 4834 12132 4866
rect 12164 4834 12200 4866
rect 12232 4834 12268 4866
rect 12300 4834 12336 4866
rect 12368 4834 12404 4866
rect 12436 4834 12472 4866
rect 12504 4834 12540 4866
rect 12572 4834 12608 4866
rect 12640 4834 12676 4866
rect 12708 4834 12744 4866
rect 12776 4834 12812 4866
rect 12844 4834 12880 4866
rect 12912 4834 12948 4866
rect 12980 4834 13016 4866
rect 13048 4834 13084 4866
rect 13116 4834 13152 4866
rect 13184 4834 13220 4866
rect 13252 4834 13288 4866
rect 13320 4834 13356 4866
rect 13388 4834 13424 4866
rect 13456 4834 13492 4866
rect 13524 4834 13560 4866
rect 13592 4834 13628 4866
rect 13660 4834 13696 4866
rect 13728 4834 13764 4866
rect 13796 4834 13832 4866
rect 13864 4834 13900 4866
rect 13932 4834 13968 4866
rect 14000 4834 14036 4866
rect 14068 4834 14104 4866
rect 14136 4834 14172 4866
rect 14204 4834 14240 4866
rect 14272 4834 14308 4866
rect 14340 4834 14376 4866
rect 14408 4834 14444 4866
rect 14476 4834 14512 4866
rect 14544 4834 14580 4866
rect 14612 4834 14648 4866
rect 14680 4834 14716 4866
rect 14748 4834 14784 4866
rect 14816 4834 14852 4866
rect 14884 4834 14920 4866
rect 14952 4834 14988 4866
rect 15020 4834 15056 4866
rect 15088 4834 15124 4866
rect 15156 4834 15192 4866
rect 15224 4834 15260 4866
rect 15292 4834 15328 4866
rect 15360 4834 15396 4866
rect 15428 4834 15464 4866
rect 15496 4834 15532 4866
rect 15564 4834 15600 4866
rect 15632 4834 15668 4866
rect 15700 4834 15736 4866
rect 15768 4834 15804 4866
rect 15836 4834 15872 4866
rect 15904 4834 15940 4866
rect 15972 4834 16000 4866
rect 0 4816 16000 4834
rect 0 4770 68 4816
rect 0 4738 18 4770
rect 50 4738 68 4770
rect 0 4702 68 4738
rect 0 4670 18 4702
rect 50 4670 68 4702
rect 0 4634 68 4670
rect 0 4602 18 4634
rect 50 4602 68 4634
rect 0 4566 68 4602
rect 0 4534 18 4566
rect 50 4534 68 4566
rect 0 4498 68 4534
rect 15932 4770 16000 4816
rect 15932 4738 15950 4770
rect 15982 4738 16000 4770
rect 15932 4702 16000 4738
rect 15932 4670 15950 4702
rect 15982 4670 16000 4702
rect 15932 4634 16000 4670
rect 15932 4602 15950 4634
rect 15982 4602 16000 4634
rect 15932 4566 16000 4602
rect 15932 4534 15950 4566
rect 15982 4534 16000 4566
rect 0 4466 18 4498
rect 50 4466 68 4498
rect 0 4430 68 4466
rect 0 4398 18 4430
rect 50 4398 68 4430
rect 0 4362 68 4398
rect 0 4330 18 4362
rect 50 4330 68 4362
rect 0 4294 68 4330
rect 0 4262 18 4294
rect 50 4262 68 4294
rect 0 4226 68 4262
rect 0 4194 18 4226
rect 50 4194 68 4226
rect 0 4158 68 4194
rect 0 4126 18 4158
rect 50 4126 68 4158
rect 0 4090 68 4126
rect 0 4058 18 4090
rect 50 4058 68 4090
rect 0 4022 68 4058
rect 0 3990 18 4022
rect 50 3990 68 4022
rect 0 3954 68 3990
rect 0 3922 18 3954
rect 50 3922 68 3954
rect 0 3886 68 3922
rect 0 3854 18 3886
rect 50 3854 68 3886
rect 0 3818 68 3854
rect 0 3786 18 3818
rect 50 3786 68 3818
rect 0 3750 68 3786
rect 0 3718 18 3750
rect 50 3718 68 3750
rect 0 3682 68 3718
rect 0 3650 18 3682
rect 50 3650 68 3682
rect 0 3614 68 3650
rect 0 3582 18 3614
rect 50 3582 68 3614
rect 0 3546 68 3582
rect 0 3514 18 3546
rect 50 3514 68 3546
rect 0 3478 68 3514
rect 0 3446 18 3478
rect 50 3446 68 3478
rect 0 3410 68 3446
rect 0 3378 18 3410
rect 50 3378 68 3410
rect 0 3342 68 3378
rect 0 3310 18 3342
rect 50 3310 68 3342
rect 0 3274 68 3310
rect 0 3242 18 3274
rect 50 3242 68 3274
rect 0 3206 68 3242
rect 0 3174 18 3206
rect 50 3174 68 3206
rect 0 3138 68 3174
rect 0 3106 18 3138
rect 50 3106 68 3138
rect 0 3070 68 3106
rect 0 3038 18 3070
rect 50 3038 68 3070
rect 0 3002 68 3038
rect 0 2970 18 3002
rect 50 2970 68 3002
rect 0 2934 68 2970
rect 0 2902 18 2934
rect 50 2902 68 2934
rect 0 2866 68 2902
rect 0 2834 18 2866
rect 50 2834 68 2866
rect 0 2798 68 2834
rect 0 2766 18 2798
rect 50 2766 68 2798
rect 0 2730 68 2766
rect 0 2698 18 2730
rect 50 2698 68 2730
rect 0 2662 68 2698
rect 0 2630 18 2662
rect 50 2630 68 2662
rect 0 2594 68 2630
rect 0 2562 18 2594
rect 50 2562 68 2594
rect 0 2526 68 2562
rect 0 2494 18 2526
rect 50 2494 68 2526
rect 0 2458 68 2494
rect 0 2426 18 2458
rect 50 2426 68 2458
rect 0 2390 68 2426
rect 0 2358 18 2390
rect 50 2358 68 2390
rect 0 2322 68 2358
rect 0 2290 18 2322
rect 50 2290 68 2322
rect 0 2254 68 2290
rect 0 2222 18 2254
rect 50 2222 68 2254
rect 0 2186 68 2222
rect 0 2154 18 2186
rect 50 2154 68 2186
rect 0 2118 68 2154
rect 0 2086 18 2118
rect 50 2086 68 2118
rect 0 2050 68 2086
rect 0 2018 18 2050
rect 50 2018 68 2050
rect 0 1982 68 2018
rect 0 1950 18 1982
rect 50 1950 68 1982
rect 0 1914 68 1950
rect 0 1882 18 1914
rect 50 1882 68 1914
rect 0 1846 68 1882
rect 0 1814 18 1846
rect 50 1814 68 1846
rect 0 1778 68 1814
rect 0 1746 18 1778
rect 50 1746 68 1778
rect 0 1710 68 1746
rect 0 1678 18 1710
rect 50 1678 68 1710
rect 0 1642 68 1678
rect 0 1610 18 1642
rect 50 1610 68 1642
rect 0 1574 68 1610
rect 0 1542 18 1574
rect 50 1542 68 1574
rect 0 1506 68 1542
rect 0 1474 18 1506
rect 50 1474 68 1506
rect 0 1438 68 1474
rect 0 1406 18 1438
rect 50 1406 68 1438
rect 0 1370 68 1406
rect 0 1338 18 1370
rect 50 1338 68 1370
rect 0 1302 68 1338
rect 0 1270 18 1302
rect 50 1270 68 1302
rect 0 1234 68 1270
rect 0 1202 18 1234
rect 50 1202 68 1234
rect 0 1166 68 1202
rect 0 1134 18 1166
rect 50 1134 68 1166
rect 0 1098 68 1134
rect 0 1066 18 1098
rect 50 1066 68 1098
rect 0 1030 68 1066
rect 0 998 18 1030
rect 50 998 68 1030
rect 0 962 68 998
rect 0 930 18 962
rect 50 930 68 962
rect 0 894 68 930
rect 0 862 18 894
rect 50 862 68 894
rect 0 826 68 862
rect 0 794 18 826
rect 50 794 68 826
rect 0 758 68 794
rect 0 726 18 758
rect 50 726 68 758
rect 0 690 68 726
rect 0 658 18 690
rect 50 658 68 690
rect 0 622 68 658
rect 0 590 18 622
rect 50 590 68 622
rect 0 554 68 590
rect 0 522 18 554
rect 50 522 68 554
rect 0 486 68 522
rect 0 454 18 486
rect 50 454 68 486
rect 0 418 68 454
rect 0 386 18 418
rect 50 386 68 418
rect 0 350 68 386
rect 15932 4498 16000 4534
rect 15932 4466 15950 4498
rect 15982 4466 16000 4498
rect 15932 4430 16000 4466
rect 15932 4398 15950 4430
rect 15982 4398 16000 4430
rect 15932 4362 16000 4398
rect 15932 4330 15950 4362
rect 15982 4330 16000 4362
rect 15932 4294 16000 4330
rect 15932 4262 15950 4294
rect 15982 4262 16000 4294
rect 15932 4226 16000 4262
rect 15932 4194 15950 4226
rect 15982 4194 16000 4226
rect 15932 4158 16000 4194
rect 15932 4126 15950 4158
rect 15982 4126 16000 4158
rect 15932 4090 16000 4126
rect 15932 4058 15950 4090
rect 15982 4058 16000 4090
rect 15932 4022 16000 4058
rect 15932 3990 15950 4022
rect 15982 3990 16000 4022
rect 15932 3954 16000 3990
rect 15932 3922 15950 3954
rect 15982 3922 16000 3954
rect 15932 3886 16000 3922
rect 15932 3854 15950 3886
rect 15982 3854 16000 3886
rect 15932 3818 16000 3854
rect 15932 3786 15950 3818
rect 15982 3786 16000 3818
rect 15932 3750 16000 3786
rect 15932 3718 15950 3750
rect 15982 3718 16000 3750
rect 15932 3682 16000 3718
rect 15932 3650 15950 3682
rect 15982 3650 16000 3682
rect 15932 3614 16000 3650
rect 15932 3582 15950 3614
rect 15982 3582 16000 3614
rect 15932 3546 16000 3582
rect 15932 3514 15950 3546
rect 15982 3514 16000 3546
rect 15932 3478 16000 3514
rect 15932 3446 15950 3478
rect 15982 3446 16000 3478
rect 15932 3410 16000 3446
rect 15932 3378 15950 3410
rect 15982 3378 16000 3410
rect 15932 3342 16000 3378
rect 15932 3310 15950 3342
rect 15982 3310 16000 3342
rect 15932 3274 16000 3310
rect 15932 3242 15950 3274
rect 15982 3242 16000 3274
rect 15932 3206 16000 3242
rect 15932 3174 15950 3206
rect 15982 3174 16000 3206
rect 15932 3138 16000 3174
rect 15932 3106 15950 3138
rect 15982 3106 16000 3138
rect 15932 3070 16000 3106
rect 15932 3038 15950 3070
rect 15982 3038 16000 3070
rect 15932 3002 16000 3038
rect 15932 2970 15950 3002
rect 15982 2970 16000 3002
rect 15932 2934 16000 2970
rect 15932 2902 15950 2934
rect 15982 2902 16000 2934
rect 15932 2866 16000 2902
rect 15932 2834 15950 2866
rect 15982 2834 16000 2866
rect 15932 2798 16000 2834
rect 15932 2766 15950 2798
rect 15982 2766 16000 2798
rect 15932 2730 16000 2766
rect 15932 2698 15950 2730
rect 15982 2698 16000 2730
rect 15932 2662 16000 2698
rect 15932 2630 15950 2662
rect 15982 2630 16000 2662
rect 15932 2594 16000 2630
rect 15932 2562 15950 2594
rect 15982 2562 16000 2594
rect 15932 2526 16000 2562
rect 15932 2494 15950 2526
rect 15982 2494 16000 2526
rect 15932 2458 16000 2494
rect 15932 2426 15950 2458
rect 15982 2426 16000 2458
rect 15932 2390 16000 2426
rect 15932 2358 15950 2390
rect 15982 2358 16000 2390
rect 15932 2322 16000 2358
rect 15932 2290 15950 2322
rect 15982 2290 16000 2322
rect 15932 2254 16000 2290
rect 15932 2222 15950 2254
rect 15982 2222 16000 2254
rect 15932 2186 16000 2222
rect 15932 2154 15950 2186
rect 15982 2154 16000 2186
rect 15932 2118 16000 2154
rect 15932 2086 15950 2118
rect 15982 2086 16000 2118
rect 15932 2050 16000 2086
rect 15932 2018 15950 2050
rect 15982 2018 16000 2050
rect 15932 1982 16000 2018
rect 15932 1950 15950 1982
rect 15982 1950 16000 1982
rect 15932 1914 16000 1950
rect 15932 1882 15950 1914
rect 15982 1882 16000 1914
rect 15932 1846 16000 1882
rect 15932 1814 15950 1846
rect 15982 1814 16000 1846
rect 15932 1778 16000 1814
rect 15932 1746 15950 1778
rect 15982 1746 16000 1778
rect 15932 1710 16000 1746
rect 15932 1678 15950 1710
rect 15982 1678 16000 1710
rect 15932 1642 16000 1678
rect 15932 1610 15950 1642
rect 15982 1610 16000 1642
rect 15932 1574 16000 1610
rect 15932 1542 15950 1574
rect 15982 1542 16000 1574
rect 15932 1506 16000 1542
rect 15932 1474 15950 1506
rect 15982 1474 16000 1506
rect 15932 1438 16000 1474
rect 15932 1406 15950 1438
rect 15982 1406 16000 1438
rect 15932 1370 16000 1406
rect 15932 1338 15950 1370
rect 15982 1338 16000 1370
rect 15932 1302 16000 1338
rect 15932 1270 15950 1302
rect 15982 1270 16000 1302
rect 15932 1234 16000 1270
rect 15932 1202 15950 1234
rect 15982 1202 16000 1234
rect 15932 1166 16000 1202
rect 15932 1134 15950 1166
rect 15982 1134 16000 1166
rect 15932 1098 16000 1134
rect 15932 1066 15950 1098
rect 15982 1066 16000 1098
rect 15932 1030 16000 1066
rect 15932 998 15950 1030
rect 15982 998 16000 1030
rect 15932 962 16000 998
rect 15932 930 15950 962
rect 15982 930 16000 962
rect 15932 894 16000 930
rect 15932 862 15950 894
rect 15982 862 16000 894
rect 15932 826 16000 862
rect 15932 794 15950 826
rect 15982 794 16000 826
rect 15932 758 16000 794
rect 15932 726 15950 758
rect 15982 726 16000 758
rect 15932 690 16000 726
rect 15932 658 15950 690
rect 15982 658 16000 690
rect 15932 622 16000 658
rect 15932 590 15950 622
rect 15982 590 16000 622
rect 15932 554 16000 590
rect 15932 522 15950 554
rect 15982 522 16000 554
rect 15932 486 16000 522
rect 15932 454 15950 486
rect 15982 454 16000 486
rect 15932 418 16000 454
rect 15932 386 15950 418
rect 15982 386 16000 418
rect 0 318 18 350
rect 50 318 68 350
rect 0 282 68 318
rect 0 250 18 282
rect 50 250 68 282
rect 0 214 68 250
rect 0 182 18 214
rect 50 182 68 214
rect 0 146 68 182
rect 0 114 18 146
rect 50 114 68 146
rect 0 68 68 114
rect 15932 350 16000 386
rect 15932 318 15950 350
rect 15982 318 16000 350
rect 15932 282 16000 318
rect 15932 250 15950 282
rect 15982 250 16000 282
rect 15932 214 16000 250
rect 15932 182 15950 214
rect 15982 182 16000 214
rect 15932 146 16000 182
rect 15932 114 15950 146
rect 15982 114 16000 146
rect 15932 68 16000 114
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< psubdiffcont >>
rect 402 4474 434 4506
rect 470 4474 502 4506
rect 538 4474 570 4506
rect 606 4474 638 4506
rect 674 4474 706 4506
rect 742 4474 774 4506
rect 810 4474 842 4506
rect 878 4474 910 4506
rect 946 4474 978 4506
rect 1014 4474 1046 4506
rect 1082 4474 1114 4506
rect 1150 4474 1182 4506
rect 1218 4474 1250 4506
rect 1286 4474 1318 4506
rect 1354 4474 1386 4506
rect 1422 4474 1454 4506
rect 1490 4474 1522 4506
rect 1558 4474 1590 4506
rect 1626 4474 1658 4506
rect 1694 4474 1726 4506
rect 1762 4474 1794 4506
rect 1830 4474 1862 4506
rect 1898 4474 1930 4506
rect 1966 4474 1998 4506
rect 2034 4474 2066 4506
rect 2102 4474 2134 4506
rect 2170 4474 2202 4506
rect 2238 4474 2270 4506
rect 2306 4474 2338 4506
rect 2374 4474 2406 4506
rect 2442 4474 2474 4506
rect 2510 4474 2542 4506
rect 2578 4474 2610 4506
rect 2646 4474 2678 4506
rect 2714 4474 2746 4506
rect 2782 4474 2814 4506
rect 2850 4474 2882 4506
rect 2918 4474 2950 4506
rect 2986 4474 3018 4506
rect 3054 4474 3086 4506
rect 3122 4474 3154 4506
rect 3190 4474 3222 4506
rect 3258 4474 3290 4506
rect 3326 4474 3358 4506
rect 3394 4474 3426 4506
rect 3462 4474 3494 4506
rect 3530 4474 3562 4506
rect 3598 4474 3630 4506
rect 3666 4474 3698 4506
rect 3734 4474 3766 4506
rect 3802 4474 3834 4506
rect 3870 4474 3902 4506
rect 3938 4474 3970 4506
rect 4006 4474 4038 4506
rect 4074 4474 4106 4506
rect 4142 4474 4174 4506
rect 4210 4474 4242 4506
rect 4278 4474 4310 4506
rect 4346 4474 4378 4506
rect 4414 4474 4446 4506
rect 4482 4474 4514 4506
rect 4550 4474 4582 4506
rect 4618 4474 4650 4506
rect 4686 4474 4718 4506
rect 4754 4474 4786 4506
rect 4822 4474 4854 4506
rect 4890 4474 4922 4506
rect 4958 4474 4990 4506
rect 5026 4474 5058 4506
rect 5094 4474 5126 4506
rect 5162 4474 5194 4506
rect 5230 4474 5262 4506
rect 5298 4474 5330 4506
rect 5366 4474 5398 4506
rect 5434 4474 5466 4506
rect 5502 4474 5534 4506
rect 5570 4474 5602 4506
rect 5638 4474 5670 4506
rect 5706 4474 5738 4506
rect 5774 4474 5806 4506
rect 5842 4474 5874 4506
rect 5910 4474 5942 4506
rect 5978 4474 6010 4506
rect 6046 4474 6078 4506
rect 6114 4474 6146 4506
rect 6182 4474 6214 4506
rect 6250 4474 6282 4506
rect 6318 4474 6350 4506
rect 6386 4474 6418 4506
rect 6454 4474 6486 4506
rect 6522 4474 6554 4506
rect 6590 4474 6622 4506
rect 6658 4474 6690 4506
rect 6726 4474 6758 4506
rect 6794 4474 6826 4506
rect 6862 4474 6894 4506
rect 6930 4474 6962 4506
rect 6998 4474 7030 4506
rect 7066 4474 7098 4506
rect 7134 4474 7166 4506
rect 7202 4474 7234 4506
rect 7270 4474 7302 4506
rect 7338 4474 7370 4506
rect 7406 4474 7438 4506
rect 7474 4474 7506 4506
rect 7542 4474 7574 4506
rect 7610 4474 7642 4506
rect 7678 4474 7710 4506
rect 7746 4474 7778 4506
rect 7814 4474 7846 4506
rect 7882 4474 7914 4506
rect 7950 4474 7982 4506
rect 8018 4474 8050 4506
rect 8086 4474 8118 4506
rect 8154 4474 8186 4506
rect 8222 4474 8254 4506
rect 8290 4474 8322 4506
rect 8358 4474 8390 4506
rect 8426 4474 8458 4506
rect 8494 4474 8526 4506
rect 8562 4474 8594 4506
rect 8630 4474 8662 4506
rect 8698 4474 8730 4506
rect 8766 4474 8798 4506
rect 8834 4474 8866 4506
rect 8902 4474 8934 4506
rect 8970 4474 9002 4506
rect 9038 4474 9070 4506
rect 9106 4474 9138 4506
rect 9174 4474 9206 4506
rect 9242 4474 9274 4506
rect 9310 4474 9342 4506
rect 9378 4474 9410 4506
rect 9446 4474 9478 4506
rect 9514 4474 9546 4506
rect 9582 4474 9614 4506
rect 9650 4474 9682 4506
rect 9718 4474 9750 4506
rect 9786 4474 9818 4506
rect 9854 4474 9886 4506
rect 9922 4474 9954 4506
rect 9990 4474 10022 4506
rect 10058 4474 10090 4506
rect 10126 4474 10158 4506
rect 10194 4474 10226 4506
rect 10262 4474 10294 4506
rect 10330 4474 10362 4506
rect 10398 4474 10430 4506
rect 10466 4474 10498 4506
rect 10534 4474 10566 4506
rect 10602 4474 10634 4506
rect 10670 4474 10702 4506
rect 10738 4474 10770 4506
rect 10806 4474 10838 4506
rect 10874 4474 10906 4506
rect 10942 4474 10974 4506
rect 11010 4474 11042 4506
rect 11078 4474 11110 4506
rect 11146 4474 11178 4506
rect 11214 4474 11246 4506
rect 11282 4474 11314 4506
rect 11350 4474 11382 4506
rect 11418 4474 11450 4506
rect 11486 4474 11518 4506
rect 11554 4474 11586 4506
rect 11622 4474 11654 4506
rect 11690 4474 11722 4506
rect 11758 4474 11790 4506
rect 11826 4474 11858 4506
rect 11894 4474 11926 4506
rect 11962 4474 11994 4506
rect 12030 4474 12062 4506
rect 12098 4474 12130 4506
rect 12166 4474 12198 4506
rect 12234 4474 12266 4506
rect 12302 4474 12334 4506
rect 12370 4474 12402 4506
rect 12438 4474 12470 4506
rect 12506 4474 12538 4506
rect 12574 4474 12606 4506
rect 12642 4474 12674 4506
rect 12710 4474 12742 4506
rect 12778 4474 12810 4506
rect 12846 4474 12878 4506
rect 12914 4474 12946 4506
rect 12982 4474 13014 4506
rect 13050 4474 13082 4506
rect 13118 4474 13150 4506
rect 13186 4474 13218 4506
rect 13254 4474 13286 4506
rect 13322 4474 13354 4506
rect 13390 4474 13422 4506
rect 13458 4474 13490 4506
rect 13526 4474 13558 4506
rect 13594 4474 13626 4506
rect 13662 4474 13694 4506
rect 13730 4474 13762 4506
rect 13798 4474 13830 4506
rect 13866 4474 13898 4506
rect 13934 4474 13966 4506
rect 14002 4474 14034 4506
rect 14070 4474 14102 4506
rect 14138 4474 14170 4506
rect 14206 4474 14238 4506
rect 14274 4474 14306 4506
rect 14342 4474 14374 4506
rect 14410 4474 14442 4506
rect 14478 4474 14510 4506
rect 14546 4474 14578 4506
rect 14614 4474 14646 4506
rect 14682 4474 14714 4506
rect 14750 4474 14782 4506
rect 14818 4474 14850 4506
rect 14886 4474 14918 4506
rect 14954 4474 14986 4506
rect 15022 4474 15054 4506
rect 15090 4474 15122 4506
rect 15158 4474 15190 4506
rect 15226 4474 15258 4506
rect 15294 4474 15326 4506
rect 15362 4474 15394 4506
rect 15430 4474 15462 4506
rect 15498 4474 15530 4506
rect 15566 4474 15598 4506
rect 378 4364 410 4396
rect 15590 4364 15622 4396
rect 378 4296 410 4328
rect 378 4228 410 4260
rect 378 4160 410 4192
rect 378 4092 410 4124
rect 378 4024 410 4056
rect 378 3956 410 3988
rect 378 3888 410 3920
rect 378 3820 410 3852
rect 378 3752 410 3784
rect 378 3684 410 3716
rect 378 3616 410 3648
rect 378 3548 410 3580
rect 378 3480 410 3512
rect 15590 4296 15622 4328
rect 15590 4228 15622 4260
rect 15590 4160 15622 4192
rect 15590 4092 15622 4124
rect 15590 4024 15622 4056
rect 15590 3956 15622 3988
rect 15590 3888 15622 3920
rect 15590 3820 15622 3852
rect 15590 3752 15622 3784
rect 15590 3684 15622 3716
rect 15590 3616 15622 3648
rect 15590 3548 15622 3580
rect 15590 3480 15622 3512
rect 378 3412 410 3444
rect 378 3344 410 3376
rect 15590 3412 15622 3444
rect 378 3276 410 3308
rect 378 3208 410 3240
rect 378 3140 410 3172
rect 378 3072 410 3104
rect 378 3004 410 3036
rect 378 2936 410 2968
rect 378 2868 410 2900
rect 378 2800 410 2832
rect 378 2732 410 2764
rect 378 2664 410 2696
rect 378 2596 410 2628
rect 378 2528 410 2560
rect 378 2460 410 2492
rect 15590 3344 15622 3376
rect 15590 3276 15622 3308
rect 15590 3208 15622 3240
rect 15590 3140 15622 3172
rect 15590 3072 15622 3104
rect 15590 3004 15622 3036
rect 15590 2936 15622 2968
rect 15590 2868 15622 2900
rect 15590 2800 15622 2832
rect 15590 2732 15622 2764
rect 15590 2664 15622 2696
rect 15590 2596 15622 2628
rect 15590 2528 15622 2560
rect 378 2392 410 2424
rect 15590 2460 15622 2492
rect 378 2324 410 2356
rect 378 2256 410 2288
rect 378 2188 410 2220
rect 378 2120 410 2152
rect 378 2052 410 2084
rect 378 1984 410 2016
rect 378 1916 410 1948
rect 378 1848 410 1880
rect 378 1780 410 1812
rect 378 1712 410 1744
rect 378 1644 410 1676
rect 378 1576 410 1608
rect 378 1508 410 1540
rect 15590 2392 15622 2424
rect 15590 2324 15622 2356
rect 15590 2256 15622 2288
rect 15590 2188 15622 2220
rect 15590 2120 15622 2152
rect 15590 2052 15622 2084
rect 15590 1984 15622 2016
rect 15590 1916 15622 1948
rect 15590 1848 15622 1880
rect 15590 1780 15622 1812
rect 15590 1712 15622 1744
rect 15590 1644 15622 1676
rect 15590 1576 15622 1608
rect 378 1440 410 1472
rect 15590 1508 15622 1540
rect 15590 1440 15622 1472
rect 378 1372 410 1404
rect 378 1304 410 1336
rect 378 1236 410 1268
rect 378 1168 410 1200
rect 378 1100 410 1132
rect 378 1032 410 1064
rect 378 964 410 996
rect 378 896 410 928
rect 378 828 410 860
rect 378 760 410 792
rect 378 692 410 724
rect 378 624 410 656
rect 378 556 410 588
rect 15590 1372 15622 1404
rect 15590 1304 15622 1336
rect 15590 1236 15622 1268
rect 15590 1168 15622 1200
rect 15590 1100 15622 1132
rect 15590 1032 15622 1064
rect 15590 964 15622 996
rect 15590 896 15622 928
rect 15590 828 15622 860
rect 15590 760 15622 792
rect 15590 692 15622 724
rect 15590 624 15622 656
rect 15590 556 15622 588
rect 378 488 410 520
rect 15590 488 15622 520
rect 402 378 434 410
rect 470 378 502 410
rect 538 378 570 410
rect 606 378 638 410
rect 674 378 706 410
rect 742 378 774 410
rect 810 378 842 410
rect 878 378 910 410
rect 946 378 978 410
rect 1014 378 1046 410
rect 1082 378 1114 410
rect 1150 378 1182 410
rect 1218 378 1250 410
rect 1286 378 1318 410
rect 1354 378 1386 410
rect 1422 378 1454 410
rect 1490 378 1522 410
rect 1558 378 1590 410
rect 1626 378 1658 410
rect 1694 378 1726 410
rect 1762 378 1794 410
rect 1830 378 1862 410
rect 1898 378 1930 410
rect 1966 378 1998 410
rect 2034 378 2066 410
rect 2102 378 2134 410
rect 2170 378 2202 410
rect 2238 378 2270 410
rect 2306 378 2338 410
rect 2374 378 2406 410
rect 2442 378 2474 410
rect 2510 378 2542 410
rect 2578 378 2610 410
rect 2646 378 2678 410
rect 2714 378 2746 410
rect 2782 378 2814 410
rect 2850 378 2882 410
rect 2918 378 2950 410
rect 2986 378 3018 410
rect 3054 378 3086 410
rect 3122 378 3154 410
rect 3190 378 3222 410
rect 3258 378 3290 410
rect 3326 378 3358 410
rect 3394 378 3426 410
rect 3462 378 3494 410
rect 3530 378 3562 410
rect 3598 378 3630 410
rect 3666 378 3698 410
rect 3734 378 3766 410
rect 3802 378 3834 410
rect 3870 378 3902 410
rect 3938 378 3970 410
rect 4006 378 4038 410
rect 4074 378 4106 410
rect 4142 378 4174 410
rect 4210 378 4242 410
rect 4278 378 4310 410
rect 4346 378 4378 410
rect 4414 378 4446 410
rect 4482 378 4514 410
rect 4550 378 4582 410
rect 4618 378 4650 410
rect 4686 378 4718 410
rect 4754 378 4786 410
rect 4822 378 4854 410
rect 4890 378 4922 410
rect 4958 378 4990 410
rect 5026 378 5058 410
rect 5094 378 5126 410
rect 5162 378 5194 410
rect 5230 378 5262 410
rect 5298 378 5330 410
rect 5366 378 5398 410
rect 5434 378 5466 410
rect 5502 378 5534 410
rect 5570 378 5602 410
rect 5638 378 5670 410
rect 5706 378 5738 410
rect 5774 378 5806 410
rect 5842 378 5874 410
rect 5910 378 5942 410
rect 5978 378 6010 410
rect 6046 378 6078 410
rect 6114 378 6146 410
rect 6182 378 6214 410
rect 6250 378 6282 410
rect 6318 378 6350 410
rect 6386 378 6418 410
rect 6454 378 6486 410
rect 6522 378 6554 410
rect 6590 378 6622 410
rect 6658 378 6690 410
rect 6726 378 6758 410
rect 6794 378 6826 410
rect 6862 378 6894 410
rect 6930 378 6962 410
rect 6998 378 7030 410
rect 7066 378 7098 410
rect 7134 378 7166 410
rect 7202 378 7234 410
rect 7270 378 7302 410
rect 7338 378 7370 410
rect 7406 378 7438 410
rect 7474 378 7506 410
rect 7542 378 7574 410
rect 7610 378 7642 410
rect 7678 378 7710 410
rect 7746 378 7778 410
rect 7814 378 7846 410
rect 7882 378 7914 410
rect 7950 378 7982 410
rect 8018 378 8050 410
rect 8086 378 8118 410
rect 8154 378 8186 410
rect 8222 378 8254 410
rect 8290 378 8322 410
rect 8358 378 8390 410
rect 8426 378 8458 410
rect 8494 378 8526 410
rect 8562 378 8594 410
rect 8630 378 8662 410
rect 8698 378 8730 410
rect 8766 378 8798 410
rect 8834 378 8866 410
rect 8902 378 8934 410
rect 8970 378 9002 410
rect 9038 378 9070 410
rect 9106 378 9138 410
rect 9174 378 9206 410
rect 9242 378 9274 410
rect 9310 378 9342 410
rect 9378 378 9410 410
rect 9446 378 9478 410
rect 9514 378 9546 410
rect 9582 378 9614 410
rect 9650 378 9682 410
rect 9718 378 9750 410
rect 9786 378 9818 410
rect 9854 378 9886 410
rect 9922 378 9954 410
rect 9990 378 10022 410
rect 10058 378 10090 410
rect 10126 378 10158 410
rect 10194 378 10226 410
rect 10262 378 10294 410
rect 10330 378 10362 410
rect 10398 378 10430 410
rect 10466 378 10498 410
rect 10534 378 10566 410
rect 10602 378 10634 410
rect 10670 378 10702 410
rect 10738 378 10770 410
rect 10806 378 10838 410
rect 10874 378 10906 410
rect 10942 378 10974 410
rect 11010 378 11042 410
rect 11078 378 11110 410
rect 11146 378 11178 410
rect 11214 378 11246 410
rect 11282 378 11314 410
rect 11350 378 11382 410
rect 11418 378 11450 410
rect 11486 378 11518 410
rect 11554 378 11586 410
rect 11622 378 11654 410
rect 11690 378 11722 410
rect 11758 378 11790 410
rect 11826 378 11858 410
rect 11894 378 11926 410
rect 11962 378 11994 410
rect 12030 378 12062 410
rect 12098 378 12130 410
rect 12166 378 12198 410
rect 12234 378 12266 410
rect 12302 378 12334 410
rect 12370 378 12402 410
rect 12438 378 12470 410
rect 12506 378 12538 410
rect 12574 378 12606 410
rect 12642 378 12674 410
rect 12710 378 12742 410
rect 12778 378 12810 410
rect 12846 378 12878 410
rect 12914 378 12946 410
rect 12982 378 13014 410
rect 13050 378 13082 410
rect 13118 378 13150 410
rect 13186 378 13218 410
rect 13254 378 13286 410
rect 13322 378 13354 410
rect 13390 378 13422 410
rect 13458 378 13490 410
rect 13526 378 13558 410
rect 13594 378 13626 410
rect 13662 378 13694 410
rect 13730 378 13762 410
rect 13798 378 13830 410
rect 13866 378 13898 410
rect 13934 378 13966 410
rect 14002 378 14034 410
rect 14070 378 14102 410
rect 14138 378 14170 410
rect 14206 378 14238 410
rect 14274 378 14306 410
rect 14342 378 14374 410
rect 14410 378 14442 410
rect 14478 378 14510 410
rect 14546 378 14578 410
rect 14614 378 14646 410
rect 14682 378 14714 410
rect 14750 378 14782 410
rect 14818 378 14850 410
rect 14886 378 14918 410
rect 14954 378 14986 410
rect 15022 378 15054 410
rect 15090 378 15122 410
rect 15158 378 15190 410
rect 15226 378 15258 410
rect 15294 378 15326 410
rect 15362 378 15394 410
rect 15430 378 15462 410
rect 15498 378 15530 410
rect 15566 378 15598 410
<< nsubdiffcont >>
rect 28 4834 60 4866
rect 96 4834 128 4866
rect 164 4834 196 4866
rect 232 4834 264 4866
rect 300 4834 332 4866
rect 368 4834 400 4866
rect 436 4834 468 4866
rect 504 4834 536 4866
rect 572 4834 604 4866
rect 640 4834 672 4866
rect 708 4834 740 4866
rect 776 4834 808 4866
rect 844 4834 876 4866
rect 912 4834 944 4866
rect 980 4834 1012 4866
rect 1048 4834 1080 4866
rect 1116 4834 1148 4866
rect 1184 4834 1216 4866
rect 1252 4834 1284 4866
rect 1320 4834 1352 4866
rect 1388 4834 1420 4866
rect 1456 4834 1488 4866
rect 1524 4834 1556 4866
rect 1592 4834 1624 4866
rect 1660 4834 1692 4866
rect 1728 4834 1760 4866
rect 1796 4834 1828 4866
rect 1864 4834 1896 4866
rect 1932 4834 1964 4866
rect 2000 4834 2032 4866
rect 2068 4834 2100 4866
rect 2136 4834 2168 4866
rect 2204 4834 2236 4866
rect 2272 4834 2304 4866
rect 2340 4834 2372 4866
rect 2408 4834 2440 4866
rect 2476 4834 2508 4866
rect 2544 4834 2576 4866
rect 2612 4834 2644 4866
rect 2680 4834 2712 4866
rect 2748 4834 2780 4866
rect 2816 4834 2848 4866
rect 2884 4834 2916 4866
rect 2952 4834 2984 4866
rect 3020 4834 3052 4866
rect 3088 4834 3120 4866
rect 3156 4834 3188 4866
rect 3224 4834 3256 4866
rect 3292 4834 3324 4866
rect 3360 4834 3392 4866
rect 3428 4834 3460 4866
rect 3496 4834 3528 4866
rect 3564 4834 3596 4866
rect 3632 4834 3664 4866
rect 3700 4834 3732 4866
rect 3768 4834 3800 4866
rect 3836 4834 3868 4866
rect 3904 4834 3936 4866
rect 3972 4834 4004 4866
rect 4040 4834 4072 4866
rect 4108 4834 4140 4866
rect 4176 4834 4208 4866
rect 4244 4834 4276 4866
rect 4312 4834 4344 4866
rect 4380 4834 4412 4866
rect 4448 4834 4480 4866
rect 4516 4834 4548 4866
rect 4584 4834 4616 4866
rect 4652 4834 4684 4866
rect 4720 4834 4752 4866
rect 4788 4834 4820 4866
rect 4856 4834 4888 4866
rect 4924 4834 4956 4866
rect 4992 4834 5024 4866
rect 5060 4834 5092 4866
rect 5128 4834 5160 4866
rect 5196 4834 5228 4866
rect 5264 4834 5296 4866
rect 5332 4834 5364 4866
rect 5400 4834 5432 4866
rect 5468 4834 5500 4866
rect 5536 4834 5568 4866
rect 5604 4834 5636 4866
rect 5672 4834 5704 4866
rect 5740 4834 5772 4866
rect 5808 4834 5840 4866
rect 5876 4834 5908 4866
rect 5944 4834 5976 4866
rect 6012 4834 6044 4866
rect 6080 4834 6112 4866
rect 6148 4834 6180 4866
rect 6216 4834 6248 4866
rect 6284 4834 6316 4866
rect 6352 4834 6384 4866
rect 6420 4834 6452 4866
rect 6488 4834 6520 4866
rect 6556 4834 6588 4866
rect 6624 4834 6656 4866
rect 6692 4834 6724 4866
rect 6760 4834 6792 4866
rect 6828 4834 6860 4866
rect 6896 4834 6928 4866
rect 6964 4834 6996 4866
rect 7032 4834 7064 4866
rect 7100 4834 7132 4866
rect 7168 4834 7200 4866
rect 7236 4834 7268 4866
rect 7304 4834 7336 4866
rect 7372 4834 7404 4866
rect 7440 4834 7472 4866
rect 7508 4834 7540 4866
rect 7576 4834 7608 4866
rect 7644 4834 7676 4866
rect 7712 4834 7744 4866
rect 7780 4834 7812 4866
rect 7848 4834 7880 4866
rect 7916 4834 7948 4866
rect 7984 4834 8016 4866
rect 8052 4834 8084 4866
rect 8120 4834 8152 4866
rect 8188 4834 8220 4866
rect 8256 4834 8288 4866
rect 8324 4834 8356 4866
rect 8392 4834 8424 4866
rect 8460 4834 8492 4866
rect 8528 4834 8560 4866
rect 8596 4834 8628 4866
rect 8664 4834 8696 4866
rect 8732 4834 8764 4866
rect 8800 4834 8832 4866
rect 8868 4834 8900 4866
rect 8936 4834 8968 4866
rect 9004 4834 9036 4866
rect 9072 4834 9104 4866
rect 9140 4834 9172 4866
rect 9208 4834 9240 4866
rect 9276 4834 9308 4866
rect 9344 4834 9376 4866
rect 9412 4834 9444 4866
rect 9480 4834 9512 4866
rect 9548 4834 9580 4866
rect 9616 4834 9648 4866
rect 9684 4834 9716 4866
rect 9752 4834 9784 4866
rect 9820 4834 9852 4866
rect 9888 4834 9920 4866
rect 9956 4834 9988 4866
rect 10024 4834 10056 4866
rect 10092 4834 10124 4866
rect 10160 4834 10192 4866
rect 10228 4834 10260 4866
rect 10296 4834 10328 4866
rect 10364 4834 10396 4866
rect 10432 4834 10464 4866
rect 10500 4834 10532 4866
rect 10568 4834 10600 4866
rect 10636 4834 10668 4866
rect 10704 4834 10736 4866
rect 10772 4834 10804 4866
rect 10840 4834 10872 4866
rect 10908 4834 10940 4866
rect 10976 4834 11008 4866
rect 11044 4834 11076 4866
rect 11112 4834 11144 4866
rect 11180 4834 11212 4866
rect 11248 4834 11280 4866
rect 11316 4834 11348 4866
rect 11384 4834 11416 4866
rect 11452 4834 11484 4866
rect 11520 4834 11552 4866
rect 11588 4834 11620 4866
rect 11656 4834 11688 4866
rect 11724 4834 11756 4866
rect 11792 4834 11824 4866
rect 11860 4834 11892 4866
rect 11928 4834 11960 4866
rect 11996 4834 12028 4866
rect 12064 4834 12096 4866
rect 12132 4834 12164 4866
rect 12200 4834 12232 4866
rect 12268 4834 12300 4866
rect 12336 4834 12368 4866
rect 12404 4834 12436 4866
rect 12472 4834 12504 4866
rect 12540 4834 12572 4866
rect 12608 4834 12640 4866
rect 12676 4834 12708 4866
rect 12744 4834 12776 4866
rect 12812 4834 12844 4866
rect 12880 4834 12912 4866
rect 12948 4834 12980 4866
rect 13016 4834 13048 4866
rect 13084 4834 13116 4866
rect 13152 4834 13184 4866
rect 13220 4834 13252 4866
rect 13288 4834 13320 4866
rect 13356 4834 13388 4866
rect 13424 4834 13456 4866
rect 13492 4834 13524 4866
rect 13560 4834 13592 4866
rect 13628 4834 13660 4866
rect 13696 4834 13728 4866
rect 13764 4834 13796 4866
rect 13832 4834 13864 4866
rect 13900 4834 13932 4866
rect 13968 4834 14000 4866
rect 14036 4834 14068 4866
rect 14104 4834 14136 4866
rect 14172 4834 14204 4866
rect 14240 4834 14272 4866
rect 14308 4834 14340 4866
rect 14376 4834 14408 4866
rect 14444 4834 14476 4866
rect 14512 4834 14544 4866
rect 14580 4834 14612 4866
rect 14648 4834 14680 4866
rect 14716 4834 14748 4866
rect 14784 4834 14816 4866
rect 14852 4834 14884 4866
rect 14920 4834 14952 4866
rect 14988 4834 15020 4866
rect 15056 4834 15088 4866
rect 15124 4834 15156 4866
rect 15192 4834 15224 4866
rect 15260 4834 15292 4866
rect 15328 4834 15360 4866
rect 15396 4834 15428 4866
rect 15464 4834 15496 4866
rect 15532 4834 15564 4866
rect 15600 4834 15632 4866
rect 15668 4834 15700 4866
rect 15736 4834 15768 4866
rect 15804 4834 15836 4866
rect 15872 4834 15904 4866
rect 15940 4834 15972 4866
rect 18 4738 50 4770
rect 18 4670 50 4702
rect 18 4602 50 4634
rect 18 4534 50 4566
rect 15950 4738 15982 4770
rect 15950 4670 15982 4702
rect 15950 4602 15982 4634
rect 15950 4534 15982 4566
rect 18 4466 50 4498
rect 18 4398 50 4430
rect 18 4330 50 4362
rect 18 4262 50 4294
rect 18 4194 50 4226
rect 18 4126 50 4158
rect 18 4058 50 4090
rect 18 3990 50 4022
rect 18 3922 50 3954
rect 18 3854 50 3886
rect 18 3786 50 3818
rect 18 3718 50 3750
rect 18 3650 50 3682
rect 18 3582 50 3614
rect 18 3514 50 3546
rect 18 3446 50 3478
rect 18 3378 50 3410
rect 18 3310 50 3342
rect 18 3242 50 3274
rect 18 3174 50 3206
rect 18 3106 50 3138
rect 18 3038 50 3070
rect 18 2970 50 3002
rect 18 2902 50 2934
rect 18 2834 50 2866
rect 18 2766 50 2798
rect 18 2698 50 2730
rect 18 2630 50 2662
rect 18 2562 50 2594
rect 18 2494 50 2526
rect 18 2426 50 2458
rect 18 2358 50 2390
rect 18 2290 50 2322
rect 18 2222 50 2254
rect 18 2154 50 2186
rect 18 2086 50 2118
rect 18 2018 50 2050
rect 18 1950 50 1982
rect 18 1882 50 1914
rect 18 1814 50 1846
rect 18 1746 50 1778
rect 18 1678 50 1710
rect 18 1610 50 1642
rect 18 1542 50 1574
rect 18 1474 50 1506
rect 18 1406 50 1438
rect 18 1338 50 1370
rect 18 1270 50 1302
rect 18 1202 50 1234
rect 18 1134 50 1166
rect 18 1066 50 1098
rect 18 998 50 1030
rect 18 930 50 962
rect 18 862 50 894
rect 18 794 50 826
rect 18 726 50 758
rect 18 658 50 690
rect 18 590 50 622
rect 18 522 50 554
rect 18 454 50 486
rect 18 386 50 418
rect 15950 4466 15982 4498
rect 15950 4398 15982 4430
rect 15950 4330 15982 4362
rect 15950 4262 15982 4294
rect 15950 4194 15982 4226
rect 15950 4126 15982 4158
rect 15950 4058 15982 4090
rect 15950 3990 15982 4022
rect 15950 3922 15982 3954
rect 15950 3854 15982 3886
rect 15950 3786 15982 3818
rect 15950 3718 15982 3750
rect 15950 3650 15982 3682
rect 15950 3582 15982 3614
rect 15950 3514 15982 3546
rect 15950 3446 15982 3478
rect 15950 3378 15982 3410
rect 15950 3310 15982 3342
rect 15950 3242 15982 3274
rect 15950 3174 15982 3206
rect 15950 3106 15982 3138
rect 15950 3038 15982 3070
rect 15950 2970 15982 3002
rect 15950 2902 15982 2934
rect 15950 2834 15982 2866
rect 15950 2766 15982 2798
rect 15950 2698 15982 2730
rect 15950 2630 15982 2662
rect 15950 2562 15982 2594
rect 15950 2494 15982 2526
rect 15950 2426 15982 2458
rect 15950 2358 15982 2390
rect 15950 2290 15982 2322
rect 15950 2222 15982 2254
rect 15950 2154 15982 2186
rect 15950 2086 15982 2118
rect 15950 2018 15982 2050
rect 15950 1950 15982 1982
rect 15950 1882 15982 1914
rect 15950 1814 15982 1846
rect 15950 1746 15982 1778
rect 15950 1678 15982 1710
rect 15950 1610 15982 1642
rect 15950 1542 15982 1574
rect 15950 1474 15982 1506
rect 15950 1406 15982 1438
rect 15950 1338 15982 1370
rect 15950 1270 15982 1302
rect 15950 1202 15982 1234
rect 15950 1134 15982 1166
rect 15950 1066 15982 1098
rect 15950 998 15982 1030
rect 15950 930 15982 962
rect 15950 862 15982 894
rect 15950 794 15982 826
rect 15950 726 15982 758
rect 15950 658 15982 690
rect 15950 590 15982 622
rect 15950 522 15982 554
rect 15950 454 15982 486
rect 15950 386 15982 418
rect 18 318 50 350
rect 18 250 50 282
rect 18 182 50 214
rect 18 114 50 146
rect 15950 318 15982 350
rect 15950 250 15982 282
rect 15950 182 15982 214
rect 15950 114 15982 146
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< poly >>
rect 1571 4394 1691 4408
rect 1571 4362 1615 4394
rect 1647 4362 1691 4394
rect 1571 4334 1691 4362
rect 1927 4394 2047 4408
rect 1927 4362 1971 4394
rect 2003 4362 2047 4394
rect 1927 4334 2047 4362
rect 2175 4394 2295 4408
rect 2175 4362 2219 4394
rect 2251 4362 2295 4394
rect 2175 4334 2295 4362
rect 2531 4394 2651 4408
rect 2531 4362 2575 4394
rect 2607 4362 2651 4394
rect 2531 4334 2651 4362
rect 2779 4394 2899 4408
rect 2779 4362 2823 4394
rect 2855 4362 2899 4394
rect 2779 4334 2899 4362
rect 3135 4394 3255 4408
rect 3135 4362 3179 4394
rect 3211 4362 3255 4394
rect 3135 4334 3255 4362
rect 3383 4394 3503 4408
rect 3383 4362 3427 4394
rect 3459 4362 3503 4394
rect 3383 4334 3503 4362
rect 3739 4394 3859 4408
rect 3739 4362 3783 4394
rect 3815 4362 3859 4394
rect 3739 4334 3859 4362
rect 3987 4394 4107 4408
rect 3987 4362 4031 4394
rect 4063 4362 4107 4394
rect 3987 4334 4107 4362
rect 4343 4394 4463 4408
rect 4343 4362 4387 4394
rect 4419 4362 4463 4394
rect 4343 4334 4463 4362
rect 4591 4394 4711 4408
rect 4591 4362 4635 4394
rect 4667 4362 4711 4394
rect 4591 4334 4711 4362
rect 4947 4394 5067 4408
rect 4947 4362 4991 4394
rect 5023 4362 5067 4394
rect 4947 4334 5067 4362
rect 5195 4394 5315 4408
rect 5195 4362 5239 4394
rect 5271 4362 5315 4394
rect 5195 4334 5315 4362
rect 5551 4394 5671 4408
rect 5551 4362 5595 4394
rect 5627 4362 5671 4394
rect 5551 4334 5671 4362
rect 5799 4394 5919 4408
rect 5799 4362 5843 4394
rect 5875 4362 5919 4394
rect 5799 4334 5919 4362
rect 6155 4394 6275 4408
rect 6155 4362 6199 4394
rect 6231 4362 6275 4394
rect 6155 4334 6275 4362
rect 6403 4394 6523 4408
rect 6403 4362 6447 4394
rect 6479 4362 6523 4394
rect 6403 4334 6523 4362
rect 6759 4394 6879 4408
rect 6759 4362 6803 4394
rect 6835 4362 6879 4394
rect 6759 4334 6879 4362
rect 7007 4394 7127 4408
rect 7007 4362 7051 4394
rect 7083 4362 7127 4394
rect 7007 4334 7127 4362
rect 7363 4394 7483 4408
rect 7363 4362 7407 4394
rect 7439 4362 7483 4394
rect 7363 4334 7483 4362
rect 7611 4394 7731 4408
rect 7611 4362 7655 4394
rect 7687 4362 7731 4394
rect 7611 4334 7731 4362
rect 7967 4394 8087 4408
rect 7967 4362 8011 4394
rect 8043 4362 8087 4394
rect 7967 4334 8087 4362
rect 8215 4394 8335 4408
rect 8215 4362 8259 4394
rect 8291 4362 8335 4394
rect 8215 4334 8335 4362
rect 8571 4394 8691 4408
rect 8571 4362 8615 4394
rect 8647 4362 8691 4394
rect 8571 4334 8691 4362
rect 8819 4394 8939 4408
rect 8819 4362 8863 4394
rect 8895 4362 8939 4394
rect 8819 4334 8939 4362
rect 9175 4394 9295 4408
rect 9175 4362 9219 4394
rect 9251 4362 9295 4394
rect 9175 4334 9295 4362
rect 9423 4394 9543 4408
rect 9423 4362 9467 4394
rect 9499 4362 9543 4394
rect 9423 4334 9543 4362
rect 9779 4394 9899 4408
rect 9779 4362 9823 4394
rect 9855 4362 9899 4394
rect 9779 4334 9899 4362
rect 10027 4394 10147 4408
rect 10027 4362 10071 4394
rect 10103 4362 10147 4394
rect 10027 4334 10147 4362
rect 10383 4394 10503 4408
rect 10383 4362 10427 4394
rect 10459 4362 10503 4394
rect 10383 4334 10503 4362
rect 10631 4394 10751 4408
rect 10631 4362 10675 4394
rect 10707 4362 10751 4394
rect 10631 4334 10751 4362
rect 10987 4394 11107 4408
rect 10987 4362 11031 4394
rect 11063 4362 11107 4394
rect 10987 4334 11107 4362
rect 11235 4394 11355 4408
rect 11235 4362 11279 4394
rect 11311 4362 11355 4394
rect 11235 4334 11355 4362
rect 11591 4394 11711 4408
rect 11591 4362 11635 4394
rect 11667 4362 11711 4394
rect 11591 4334 11711 4362
rect 11839 4394 11959 4408
rect 11839 4362 11883 4394
rect 11915 4362 11959 4394
rect 11839 4334 11959 4362
rect 12195 4394 12315 4408
rect 12195 4362 12239 4394
rect 12271 4362 12315 4394
rect 12195 4334 12315 4362
rect 12443 4394 12563 4408
rect 12443 4362 12487 4394
rect 12519 4362 12563 4394
rect 12443 4334 12563 4362
rect 12799 4394 12919 4408
rect 12799 4362 12843 4394
rect 12875 4362 12919 4394
rect 12799 4334 12919 4362
rect 13047 4394 13167 4408
rect 13047 4362 13091 4394
rect 13123 4362 13167 4394
rect 13047 4334 13167 4362
rect 13403 4394 13523 4408
rect 13403 4362 13447 4394
rect 13479 4362 13523 4394
rect 13403 4334 13523 4362
rect 13651 4394 13771 4408
rect 13651 4362 13695 4394
rect 13727 4362 13771 4394
rect 13651 4334 13771 4362
rect 14007 4394 14127 4408
rect 14007 4362 14051 4394
rect 14083 4362 14127 4394
rect 14007 4334 14127 4362
rect 14255 4394 14375 4408
rect 14255 4362 14299 4394
rect 14331 4362 14375 4394
rect 14255 4334 14375 4362
rect 1571 3426 1691 3454
rect 1571 3394 1615 3426
rect 1647 3394 1691 3426
rect 1571 3366 1691 3394
rect 1927 3426 2047 3454
rect 1927 3394 1971 3426
rect 2003 3394 2047 3426
rect 1927 3366 2047 3394
rect 2175 3426 2295 3454
rect 2175 3394 2219 3426
rect 2251 3394 2295 3426
rect 2175 3366 2295 3394
rect 2531 3426 2651 3454
rect 2531 3394 2575 3426
rect 2607 3394 2651 3426
rect 2531 3366 2651 3394
rect 2779 3426 2899 3454
rect 2779 3394 2823 3426
rect 2855 3394 2899 3426
rect 2779 3366 2899 3394
rect 3135 3426 3255 3454
rect 3135 3394 3179 3426
rect 3211 3394 3255 3426
rect 3135 3366 3255 3394
rect 3383 3426 3503 3454
rect 3383 3394 3427 3426
rect 3459 3394 3503 3426
rect 3383 3366 3503 3394
rect 3739 3426 3859 3454
rect 3739 3394 3783 3426
rect 3815 3394 3859 3426
rect 3739 3366 3859 3394
rect 3987 3426 4107 3454
rect 3987 3394 4031 3426
rect 4063 3394 4107 3426
rect 3987 3366 4107 3394
rect 4343 3426 4463 3454
rect 4343 3394 4387 3426
rect 4419 3394 4463 3426
rect 4343 3366 4463 3394
rect 4591 3426 4711 3454
rect 4591 3394 4635 3426
rect 4667 3394 4711 3426
rect 4591 3366 4711 3394
rect 4947 3426 5067 3454
rect 4947 3394 4991 3426
rect 5023 3394 5067 3426
rect 4947 3366 5067 3394
rect 5195 3426 5315 3454
rect 5195 3394 5239 3426
rect 5271 3394 5315 3426
rect 5195 3366 5315 3394
rect 5551 3426 5671 3454
rect 5551 3394 5595 3426
rect 5627 3394 5671 3426
rect 5551 3366 5671 3394
rect 5799 3426 5919 3454
rect 5799 3394 5843 3426
rect 5875 3394 5919 3426
rect 5799 3366 5919 3394
rect 6155 3426 6275 3454
rect 6155 3394 6199 3426
rect 6231 3394 6275 3426
rect 6155 3366 6275 3394
rect 6403 3426 6523 3454
rect 6403 3394 6447 3426
rect 6479 3394 6523 3426
rect 6403 3366 6523 3394
rect 6759 3426 6879 3454
rect 6759 3394 6803 3426
rect 6835 3394 6879 3426
rect 6759 3366 6879 3394
rect 7007 3426 7127 3454
rect 7007 3394 7051 3426
rect 7083 3394 7127 3426
rect 7007 3366 7127 3394
rect 7363 3426 7483 3454
rect 7363 3394 7407 3426
rect 7439 3394 7483 3426
rect 7363 3366 7483 3394
rect 7611 3426 7731 3454
rect 7611 3394 7655 3426
rect 7687 3394 7731 3426
rect 7611 3366 7731 3394
rect 7967 3426 8087 3454
rect 7967 3394 8011 3426
rect 8043 3394 8087 3426
rect 7967 3366 8087 3394
rect 8215 3426 8335 3454
rect 8215 3394 8259 3426
rect 8291 3394 8335 3426
rect 8215 3366 8335 3394
rect 8571 3426 8691 3454
rect 8571 3394 8615 3426
rect 8647 3394 8691 3426
rect 8571 3366 8691 3394
rect 8819 3426 8939 3454
rect 8819 3394 8863 3426
rect 8895 3394 8939 3426
rect 8819 3366 8939 3394
rect 9175 3426 9295 3454
rect 9175 3394 9219 3426
rect 9251 3394 9295 3426
rect 9175 3366 9295 3394
rect 9423 3426 9543 3454
rect 9423 3394 9467 3426
rect 9499 3394 9543 3426
rect 9423 3366 9543 3394
rect 9779 3426 9899 3454
rect 9779 3394 9823 3426
rect 9855 3394 9899 3426
rect 9779 3366 9899 3394
rect 10027 3426 10147 3454
rect 10027 3394 10071 3426
rect 10103 3394 10147 3426
rect 10027 3366 10147 3394
rect 10383 3426 10503 3454
rect 10383 3394 10427 3426
rect 10459 3394 10503 3426
rect 10383 3366 10503 3394
rect 10631 3426 10751 3454
rect 10631 3394 10675 3426
rect 10707 3394 10751 3426
rect 10631 3366 10751 3394
rect 10987 3426 11107 3454
rect 10987 3394 11031 3426
rect 11063 3394 11107 3426
rect 10987 3366 11107 3394
rect 11235 3426 11355 3454
rect 11235 3394 11279 3426
rect 11311 3394 11355 3426
rect 11235 3366 11355 3394
rect 11591 3426 11711 3454
rect 11591 3394 11635 3426
rect 11667 3394 11711 3426
rect 11591 3366 11711 3394
rect 11839 3426 11959 3454
rect 11839 3394 11883 3426
rect 11915 3394 11959 3426
rect 11839 3366 11959 3394
rect 12195 3426 12315 3454
rect 12195 3394 12239 3426
rect 12271 3394 12315 3426
rect 12195 3366 12315 3394
rect 12443 3426 12563 3454
rect 12443 3394 12487 3426
rect 12519 3394 12563 3426
rect 12443 3366 12563 3394
rect 12799 3426 12919 3454
rect 12799 3394 12843 3426
rect 12875 3394 12919 3426
rect 12799 3366 12919 3394
rect 13047 3426 13167 3454
rect 13047 3394 13091 3426
rect 13123 3394 13167 3426
rect 13047 3366 13167 3394
rect 13403 3426 13523 3454
rect 13403 3394 13447 3426
rect 13479 3394 13523 3426
rect 13403 3366 13523 3394
rect 13651 3426 13771 3454
rect 13651 3394 13695 3426
rect 13727 3394 13771 3426
rect 13651 3366 13771 3394
rect 14007 3426 14127 3454
rect 14007 3394 14051 3426
rect 14083 3394 14127 3426
rect 14007 3366 14127 3394
rect 14255 3426 14375 3454
rect 14255 3394 14299 3426
rect 14331 3394 14375 3426
rect 14255 3366 14375 3394
rect 1571 2458 1691 2486
rect 1571 2426 1615 2458
rect 1647 2426 1691 2458
rect 1571 2398 1691 2426
rect 1927 2458 2047 2486
rect 1927 2426 1971 2458
rect 2003 2426 2047 2458
rect 1927 2398 2047 2426
rect 2175 2458 2295 2486
rect 2175 2426 2219 2458
rect 2251 2426 2295 2458
rect 2175 2398 2295 2426
rect 2531 2458 2651 2486
rect 2531 2426 2575 2458
rect 2607 2426 2651 2458
rect 2531 2398 2651 2426
rect 2779 2458 2899 2486
rect 2779 2426 2823 2458
rect 2855 2426 2899 2458
rect 2779 2398 2899 2426
rect 3135 2458 3255 2486
rect 3135 2426 3179 2458
rect 3211 2426 3255 2458
rect 3135 2398 3255 2426
rect 3383 2458 3503 2486
rect 3383 2426 3427 2458
rect 3459 2426 3503 2458
rect 3383 2398 3503 2426
rect 3739 2458 3859 2486
rect 3739 2426 3783 2458
rect 3815 2426 3859 2458
rect 3739 2398 3859 2426
rect 3987 2458 4107 2486
rect 3987 2426 4031 2458
rect 4063 2426 4107 2458
rect 3987 2398 4107 2426
rect 4343 2458 4463 2486
rect 4343 2426 4387 2458
rect 4419 2426 4463 2458
rect 4343 2398 4463 2426
rect 4591 2458 4711 2486
rect 4591 2426 4635 2458
rect 4667 2426 4711 2458
rect 4591 2398 4711 2426
rect 4947 2458 5067 2486
rect 4947 2426 4991 2458
rect 5023 2426 5067 2458
rect 4947 2398 5067 2426
rect 5195 2458 5315 2486
rect 5195 2426 5239 2458
rect 5271 2426 5315 2458
rect 5195 2398 5315 2426
rect 5551 2458 5671 2486
rect 5551 2426 5595 2458
rect 5627 2426 5671 2458
rect 5551 2398 5671 2426
rect 5799 2458 5919 2486
rect 5799 2426 5843 2458
rect 5875 2426 5919 2458
rect 5799 2398 5919 2426
rect 6155 2458 6275 2486
rect 6155 2426 6199 2458
rect 6231 2426 6275 2458
rect 6155 2398 6275 2426
rect 6403 2458 6523 2486
rect 6403 2426 6447 2458
rect 6479 2426 6523 2458
rect 6403 2398 6523 2426
rect 6759 2458 6879 2486
rect 6759 2426 6803 2458
rect 6835 2426 6879 2458
rect 6759 2398 6879 2426
rect 7007 2458 7127 2486
rect 7007 2426 7051 2458
rect 7083 2426 7127 2458
rect 7007 2398 7127 2426
rect 7363 2458 7483 2486
rect 7363 2426 7407 2458
rect 7439 2426 7483 2458
rect 7363 2398 7483 2426
rect 7611 2458 7731 2486
rect 7611 2426 7655 2458
rect 7687 2426 7731 2458
rect 7611 2398 7731 2426
rect 7967 2458 8087 2486
rect 7967 2426 8011 2458
rect 8043 2426 8087 2458
rect 7967 2398 8087 2426
rect 8215 2458 8335 2486
rect 8215 2426 8259 2458
rect 8291 2426 8335 2458
rect 8215 2398 8335 2426
rect 8571 2458 8691 2486
rect 8571 2426 8615 2458
rect 8647 2426 8691 2458
rect 8571 2398 8691 2426
rect 8819 2458 8939 2486
rect 8819 2426 8863 2458
rect 8895 2426 8939 2458
rect 8819 2398 8939 2426
rect 9175 2458 9295 2486
rect 9175 2426 9219 2458
rect 9251 2426 9295 2458
rect 9175 2398 9295 2426
rect 9423 2458 9543 2486
rect 9423 2426 9467 2458
rect 9499 2426 9543 2458
rect 9423 2398 9543 2426
rect 9779 2458 9899 2486
rect 9779 2426 9823 2458
rect 9855 2426 9899 2458
rect 9779 2398 9899 2426
rect 10027 2458 10147 2486
rect 10027 2426 10071 2458
rect 10103 2426 10147 2458
rect 10027 2398 10147 2426
rect 10383 2458 10503 2486
rect 10383 2426 10427 2458
rect 10459 2426 10503 2458
rect 10383 2398 10503 2426
rect 10631 2458 10751 2486
rect 10631 2426 10675 2458
rect 10707 2426 10751 2458
rect 10631 2398 10751 2426
rect 10987 2458 11107 2486
rect 10987 2426 11031 2458
rect 11063 2426 11107 2458
rect 10987 2398 11107 2426
rect 11235 2458 11355 2486
rect 11235 2426 11279 2458
rect 11311 2426 11355 2458
rect 11235 2398 11355 2426
rect 11591 2458 11711 2486
rect 11591 2426 11635 2458
rect 11667 2426 11711 2458
rect 11591 2398 11711 2426
rect 11839 2458 11959 2486
rect 11839 2426 11883 2458
rect 11915 2426 11959 2458
rect 11839 2398 11959 2426
rect 12195 2458 12315 2486
rect 12195 2426 12239 2458
rect 12271 2426 12315 2458
rect 12195 2398 12315 2426
rect 12443 2458 12563 2486
rect 12443 2426 12487 2458
rect 12519 2426 12563 2458
rect 12443 2398 12563 2426
rect 12799 2458 12919 2486
rect 12799 2426 12843 2458
rect 12875 2426 12919 2458
rect 12799 2398 12919 2426
rect 13047 2458 13167 2486
rect 13047 2426 13091 2458
rect 13123 2426 13167 2458
rect 13047 2398 13167 2426
rect 13403 2458 13523 2486
rect 13403 2426 13447 2458
rect 13479 2426 13523 2458
rect 13403 2398 13523 2426
rect 13651 2458 13771 2486
rect 13651 2426 13695 2458
rect 13727 2426 13771 2458
rect 13651 2398 13771 2426
rect 14007 2458 14127 2486
rect 14007 2426 14051 2458
rect 14083 2426 14127 2458
rect 14007 2398 14127 2426
rect 14255 2458 14375 2486
rect 14255 2426 14299 2458
rect 14331 2426 14375 2458
rect 14255 2398 14375 2426
rect 1571 1490 1691 1518
rect 1571 1458 1615 1490
rect 1647 1458 1691 1490
rect 1571 1430 1691 1458
rect 1927 1490 2047 1518
rect 1927 1458 1971 1490
rect 2003 1458 2047 1490
rect 1927 1430 2047 1458
rect 2175 1490 2295 1518
rect 2175 1458 2219 1490
rect 2251 1458 2295 1490
rect 2175 1430 2295 1458
rect 2531 1490 2651 1518
rect 2531 1458 2575 1490
rect 2607 1458 2651 1490
rect 2531 1430 2651 1458
rect 2779 1490 2899 1518
rect 2779 1458 2823 1490
rect 2855 1458 2899 1490
rect 2779 1430 2899 1458
rect 3135 1490 3255 1518
rect 3135 1458 3179 1490
rect 3211 1458 3255 1490
rect 3135 1430 3255 1458
rect 3383 1490 3503 1518
rect 3383 1458 3427 1490
rect 3459 1458 3503 1490
rect 3383 1430 3503 1458
rect 3739 1490 3859 1518
rect 3739 1458 3783 1490
rect 3815 1458 3859 1490
rect 3739 1430 3859 1458
rect 3987 1490 4107 1518
rect 3987 1458 4031 1490
rect 4063 1458 4107 1490
rect 3987 1430 4107 1458
rect 4343 1490 4463 1518
rect 4343 1458 4387 1490
rect 4419 1458 4463 1490
rect 4343 1430 4463 1458
rect 4591 1490 4711 1518
rect 4591 1458 4635 1490
rect 4667 1458 4711 1490
rect 4591 1430 4711 1458
rect 4947 1490 5067 1518
rect 4947 1458 4991 1490
rect 5023 1458 5067 1490
rect 4947 1430 5067 1458
rect 5195 1490 5315 1518
rect 5195 1458 5239 1490
rect 5271 1458 5315 1490
rect 5195 1430 5315 1458
rect 5551 1490 5671 1518
rect 5551 1458 5595 1490
rect 5627 1458 5671 1490
rect 5551 1430 5671 1458
rect 5799 1490 5919 1518
rect 5799 1458 5843 1490
rect 5875 1458 5919 1490
rect 5799 1430 5919 1458
rect 6155 1490 6275 1518
rect 6155 1458 6199 1490
rect 6231 1458 6275 1490
rect 6155 1430 6275 1458
rect 6403 1490 6523 1518
rect 6403 1458 6447 1490
rect 6479 1458 6523 1490
rect 6403 1430 6523 1458
rect 6759 1490 6879 1518
rect 6759 1458 6803 1490
rect 6835 1458 6879 1490
rect 6759 1430 6879 1458
rect 7007 1490 7127 1518
rect 7007 1458 7051 1490
rect 7083 1458 7127 1490
rect 7007 1430 7127 1458
rect 7363 1490 7483 1518
rect 7363 1458 7407 1490
rect 7439 1458 7483 1490
rect 7363 1430 7483 1458
rect 7611 1490 7731 1518
rect 7611 1458 7655 1490
rect 7687 1458 7731 1490
rect 7611 1430 7731 1458
rect 7967 1490 8087 1518
rect 7967 1458 8011 1490
rect 8043 1458 8087 1490
rect 7967 1430 8087 1458
rect 8215 1490 8335 1518
rect 8215 1458 8259 1490
rect 8291 1458 8335 1490
rect 8215 1430 8335 1458
rect 8571 1490 8691 1518
rect 8571 1458 8615 1490
rect 8647 1458 8691 1490
rect 8571 1430 8691 1458
rect 8819 1490 8939 1518
rect 8819 1458 8863 1490
rect 8895 1458 8939 1490
rect 8819 1430 8939 1458
rect 9175 1490 9295 1518
rect 9175 1458 9219 1490
rect 9251 1458 9295 1490
rect 9175 1430 9295 1458
rect 9423 1490 9543 1518
rect 9423 1458 9467 1490
rect 9499 1458 9543 1490
rect 9423 1430 9543 1458
rect 9779 1490 9899 1518
rect 9779 1458 9823 1490
rect 9855 1458 9899 1490
rect 9779 1430 9899 1458
rect 10027 1490 10147 1518
rect 10027 1458 10071 1490
rect 10103 1458 10147 1490
rect 10027 1430 10147 1458
rect 10383 1490 10503 1518
rect 10383 1458 10427 1490
rect 10459 1458 10503 1490
rect 10383 1430 10503 1458
rect 10631 1490 10751 1518
rect 10631 1458 10675 1490
rect 10707 1458 10751 1490
rect 10631 1430 10751 1458
rect 10987 1490 11107 1518
rect 10987 1458 11031 1490
rect 11063 1458 11107 1490
rect 10987 1430 11107 1458
rect 11235 1490 11355 1518
rect 11235 1458 11279 1490
rect 11311 1458 11355 1490
rect 11235 1430 11355 1458
rect 11591 1490 11711 1518
rect 11591 1458 11635 1490
rect 11667 1458 11711 1490
rect 11591 1430 11711 1458
rect 11839 1490 11959 1518
rect 11839 1458 11883 1490
rect 11915 1458 11959 1490
rect 11839 1430 11959 1458
rect 12195 1490 12315 1518
rect 12195 1458 12239 1490
rect 12271 1458 12315 1490
rect 12195 1430 12315 1458
rect 12443 1490 12563 1518
rect 12443 1458 12487 1490
rect 12519 1458 12563 1490
rect 12443 1430 12563 1458
rect 12799 1490 12919 1518
rect 12799 1458 12843 1490
rect 12875 1458 12919 1490
rect 12799 1430 12919 1458
rect 13047 1490 13167 1518
rect 13047 1458 13091 1490
rect 13123 1458 13167 1490
rect 13047 1430 13167 1458
rect 13403 1490 13523 1518
rect 13403 1458 13447 1490
rect 13479 1458 13523 1490
rect 13403 1430 13523 1458
rect 13651 1490 13771 1518
rect 13651 1458 13695 1490
rect 13727 1458 13771 1490
rect 13651 1430 13771 1458
rect 14007 1490 14127 1518
rect 14007 1458 14051 1490
rect 14083 1458 14127 1490
rect 14007 1430 14127 1458
rect 14255 1490 14375 1518
rect 14255 1458 14299 1490
rect 14331 1458 14375 1490
rect 14255 1430 14375 1458
rect 1571 522 1691 550
rect 1571 490 1615 522
rect 1647 490 1691 522
rect 1571 476 1691 490
rect 1927 522 2047 550
rect 1927 490 1971 522
rect 2003 490 2047 522
rect 1927 476 2047 490
rect 2175 522 2295 550
rect 2175 490 2219 522
rect 2251 490 2295 522
rect 2175 476 2295 490
rect 2531 522 2651 550
rect 2531 490 2575 522
rect 2607 490 2651 522
rect 2531 476 2651 490
rect 2779 522 2899 550
rect 2779 490 2823 522
rect 2855 490 2899 522
rect 2779 476 2899 490
rect 3135 522 3255 550
rect 3135 490 3179 522
rect 3211 490 3255 522
rect 3135 476 3255 490
rect 3383 522 3503 550
rect 3383 490 3427 522
rect 3459 490 3503 522
rect 3383 476 3503 490
rect 3739 522 3859 550
rect 3739 490 3783 522
rect 3815 490 3859 522
rect 3739 476 3859 490
rect 3987 522 4107 550
rect 3987 490 4031 522
rect 4063 490 4107 522
rect 3987 476 4107 490
rect 4343 522 4463 550
rect 4343 490 4387 522
rect 4419 490 4463 522
rect 4343 476 4463 490
rect 4591 522 4711 550
rect 4591 490 4635 522
rect 4667 490 4711 522
rect 4591 476 4711 490
rect 4947 522 5067 550
rect 4947 490 4991 522
rect 5023 490 5067 522
rect 4947 476 5067 490
rect 5195 522 5315 550
rect 5195 490 5239 522
rect 5271 490 5315 522
rect 5195 476 5315 490
rect 5551 522 5671 550
rect 5551 490 5595 522
rect 5627 490 5671 522
rect 5551 476 5671 490
rect 5799 522 5919 550
rect 5799 490 5843 522
rect 5875 490 5919 522
rect 5799 476 5919 490
rect 6155 522 6275 550
rect 6155 490 6199 522
rect 6231 490 6275 522
rect 6155 476 6275 490
rect 6403 522 6523 550
rect 6403 490 6447 522
rect 6479 490 6523 522
rect 6403 476 6523 490
rect 6759 522 6879 550
rect 6759 490 6803 522
rect 6835 490 6879 522
rect 6759 476 6879 490
rect 7007 522 7127 550
rect 7007 490 7051 522
rect 7083 490 7127 522
rect 7007 476 7127 490
rect 7363 522 7483 550
rect 7363 490 7407 522
rect 7439 490 7483 522
rect 7363 476 7483 490
rect 7611 522 7731 550
rect 7611 490 7655 522
rect 7687 490 7731 522
rect 7611 476 7731 490
rect 7967 522 8087 550
rect 7967 490 8011 522
rect 8043 490 8087 522
rect 7967 476 8087 490
rect 8215 522 8335 550
rect 8215 490 8259 522
rect 8291 490 8335 522
rect 8215 476 8335 490
rect 8571 522 8691 550
rect 8571 490 8615 522
rect 8647 490 8691 522
rect 8571 476 8691 490
rect 8819 522 8939 550
rect 8819 490 8863 522
rect 8895 490 8939 522
rect 8819 476 8939 490
rect 9175 522 9295 550
rect 9175 490 9219 522
rect 9251 490 9295 522
rect 9175 476 9295 490
rect 9423 522 9543 550
rect 9423 490 9467 522
rect 9499 490 9543 522
rect 9423 476 9543 490
rect 9779 522 9899 550
rect 9779 490 9823 522
rect 9855 490 9899 522
rect 9779 476 9899 490
rect 10027 522 10147 550
rect 10027 490 10071 522
rect 10103 490 10147 522
rect 10027 476 10147 490
rect 10383 522 10503 550
rect 10383 490 10427 522
rect 10459 490 10503 522
rect 10383 476 10503 490
rect 10631 522 10751 550
rect 10631 490 10675 522
rect 10707 490 10751 522
rect 10631 476 10751 490
rect 10987 522 11107 550
rect 10987 490 11031 522
rect 11063 490 11107 522
rect 10987 476 11107 490
rect 11235 522 11355 550
rect 11235 490 11279 522
rect 11311 490 11355 522
rect 11235 476 11355 490
rect 11591 522 11711 550
rect 11591 490 11635 522
rect 11667 490 11711 522
rect 11591 476 11711 490
rect 11839 522 11959 550
rect 11839 490 11883 522
rect 11915 490 11959 522
rect 11839 476 11959 490
rect 12195 522 12315 550
rect 12195 490 12239 522
rect 12271 490 12315 522
rect 12195 476 12315 490
rect 12443 522 12563 550
rect 12443 490 12487 522
rect 12519 490 12563 522
rect 12443 476 12563 490
rect 12799 522 12919 550
rect 12799 490 12843 522
rect 12875 490 12919 522
rect 12799 476 12919 490
rect 13047 522 13167 550
rect 13047 490 13091 522
rect 13123 490 13167 522
rect 13047 476 13167 490
rect 13403 522 13523 550
rect 13403 490 13447 522
rect 13479 490 13523 522
rect 13403 476 13523 490
rect 13651 522 13771 550
rect 13651 490 13695 522
rect 13727 490 13771 522
rect 13651 476 13771 490
rect 14007 522 14127 550
rect 14007 490 14051 522
rect 14083 490 14127 522
rect 14007 476 14127 490
rect 14255 522 14375 550
rect 14255 490 14299 522
rect 14331 490 14375 522
rect 14255 476 14375 490
<< polycont >>
rect 1615 4362 1647 4394
rect 1971 4362 2003 4394
rect 2219 4362 2251 4394
rect 2575 4362 2607 4394
rect 2823 4362 2855 4394
rect 3179 4362 3211 4394
rect 3427 4362 3459 4394
rect 3783 4362 3815 4394
rect 4031 4362 4063 4394
rect 4387 4362 4419 4394
rect 4635 4362 4667 4394
rect 4991 4362 5023 4394
rect 5239 4362 5271 4394
rect 5595 4362 5627 4394
rect 5843 4362 5875 4394
rect 6199 4362 6231 4394
rect 6447 4362 6479 4394
rect 6803 4362 6835 4394
rect 7051 4362 7083 4394
rect 7407 4362 7439 4394
rect 7655 4362 7687 4394
rect 8011 4362 8043 4394
rect 8259 4362 8291 4394
rect 8615 4362 8647 4394
rect 8863 4362 8895 4394
rect 9219 4362 9251 4394
rect 9467 4362 9499 4394
rect 9823 4362 9855 4394
rect 10071 4362 10103 4394
rect 10427 4362 10459 4394
rect 10675 4362 10707 4394
rect 11031 4362 11063 4394
rect 11279 4362 11311 4394
rect 11635 4362 11667 4394
rect 11883 4362 11915 4394
rect 12239 4362 12271 4394
rect 12487 4362 12519 4394
rect 12843 4362 12875 4394
rect 13091 4362 13123 4394
rect 13447 4362 13479 4394
rect 13695 4362 13727 4394
rect 14051 4362 14083 4394
rect 14299 4362 14331 4394
rect 1615 3394 1647 3426
rect 1971 3394 2003 3426
rect 2219 3394 2251 3426
rect 2575 3394 2607 3426
rect 2823 3394 2855 3426
rect 3179 3394 3211 3426
rect 3427 3394 3459 3426
rect 3783 3394 3815 3426
rect 4031 3394 4063 3426
rect 4387 3394 4419 3426
rect 4635 3394 4667 3426
rect 4991 3394 5023 3426
rect 5239 3394 5271 3426
rect 5595 3394 5627 3426
rect 5843 3394 5875 3426
rect 6199 3394 6231 3426
rect 6447 3394 6479 3426
rect 6803 3394 6835 3426
rect 7051 3394 7083 3426
rect 7407 3394 7439 3426
rect 7655 3394 7687 3426
rect 8011 3394 8043 3426
rect 8259 3394 8291 3426
rect 8615 3394 8647 3426
rect 8863 3394 8895 3426
rect 9219 3394 9251 3426
rect 9467 3394 9499 3426
rect 9823 3394 9855 3426
rect 10071 3394 10103 3426
rect 10427 3394 10459 3426
rect 10675 3394 10707 3426
rect 11031 3394 11063 3426
rect 11279 3394 11311 3426
rect 11635 3394 11667 3426
rect 11883 3394 11915 3426
rect 12239 3394 12271 3426
rect 12487 3394 12519 3426
rect 12843 3394 12875 3426
rect 13091 3394 13123 3426
rect 13447 3394 13479 3426
rect 13695 3394 13727 3426
rect 14051 3394 14083 3426
rect 14299 3394 14331 3426
rect 1615 2426 1647 2458
rect 1971 2426 2003 2458
rect 2219 2426 2251 2458
rect 2575 2426 2607 2458
rect 2823 2426 2855 2458
rect 3179 2426 3211 2458
rect 3427 2426 3459 2458
rect 3783 2426 3815 2458
rect 4031 2426 4063 2458
rect 4387 2426 4419 2458
rect 4635 2426 4667 2458
rect 4991 2426 5023 2458
rect 5239 2426 5271 2458
rect 5595 2426 5627 2458
rect 5843 2426 5875 2458
rect 6199 2426 6231 2458
rect 6447 2426 6479 2458
rect 6803 2426 6835 2458
rect 7051 2426 7083 2458
rect 7407 2426 7439 2458
rect 7655 2426 7687 2458
rect 8011 2426 8043 2458
rect 8259 2426 8291 2458
rect 8615 2426 8647 2458
rect 8863 2426 8895 2458
rect 9219 2426 9251 2458
rect 9467 2426 9499 2458
rect 9823 2426 9855 2458
rect 10071 2426 10103 2458
rect 10427 2426 10459 2458
rect 10675 2426 10707 2458
rect 11031 2426 11063 2458
rect 11279 2426 11311 2458
rect 11635 2426 11667 2458
rect 11883 2426 11915 2458
rect 12239 2426 12271 2458
rect 12487 2426 12519 2458
rect 12843 2426 12875 2458
rect 13091 2426 13123 2458
rect 13447 2426 13479 2458
rect 13695 2426 13727 2458
rect 14051 2426 14083 2458
rect 14299 2426 14331 2458
rect 1615 1458 1647 1490
rect 1971 1458 2003 1490
rect 2219 1458 2251 1490
rect 2575 1458 2607 1490
rect 2823 1458 2855 1490
rect 3179 1458 3211 1490
rect 3427 1458 3459 1490
rect 3783 1458 3815 1490
rect 4031 1458 4063 1490
rect 4387 1458 4419 1490
rect 4635 1458 4667 1490
rect 4991 1458 5023 1490
rect 5239 1458 5271 1490
rect 5595 1458 5627 1490
rect 5843 1458 5875 1490
rect 6199 1458 6231 1490
rect 6447 1458 6479 1490
rect 6803 1458 6835 1490
rect 7051 1458 7083 1490
rect 7407 1458 7439 1490
rect 7655 1458 7687 1490
rect 8011 1458 8043 1490
rect 8259 1458 8291 1490
rect 8615 1458 8647 1490
rect 8863 1458 8895 1490
rect 9219 1458 9251 1490
rect 9467 1458 9499 1490
rect 9823 1458 9855 1490
rect 10071 1458 10103 1490
rect 10427 1458 10459 1490
rect 10675 1458 10707 1490
rect 11031 1458 11063 1490
rect 11279 1458 11311 1490
rect 11635 1458 11667 1490
rect 11883 1458 11915 1490
rect 12239 1458 12271 1490
rect 12487 1458 12519 1490
rect 12843 1458 12875 1490
rect 13091 1458 13123 1490
rect 13447 1458 13479 1490
rect 13695 1458 13727 1490
rect 14051 1458 14083 1490
rect 14299 1458 14331 1490
rect 1615 490 1647 522
rect 1971 490 2003 522
rect 2219 490 2251 522
rect 2575 490 2607 522
rect 2823 490 2855 522
rect 3179 490 3211 522
rect 3427 490 3459 522
rect 3783 490 3815 522
rect 4031 490 4063 522
rect 4387 490 4419 522
rect 4635 490 4667 522
rect 4991 490 5023 522
rect 5239 490 5271 522
rect 5595 490 5627 522
rect 5843 490 5875 522
rect 6199 490 6231 522
rect 6447 490 6479 522
rect 6803 490 6835 522
rect 7051 490 7083 522
rect 7407 490 7439 522
rect 7655 490 7687 522
rect 8011 490 8043 522
rect 8259 490 8291 522
rect 8615 490 8647 522
rect 8863 490 8895 522
rect 9219 490 9251 522
rect 9467 490 9499 522
rect 9823 490 9855 522
rect 10071 490 10103 522
rect 10427 490 10459 522
rect 10675 490 10707 522
rect 11031 490 11063 522
rect 11279 490 11311 522
rect 11635 490 11667 522
rect 11883 490 11915 522
rect 12239 490 12271 522
rect 12487 490 12519 522
rect 12843 490 12875 522
rect 13091 490 13123 522
rect 13447 490 13479 522
rect 13695 490 13727 522
rect 14051 490 14083 522
rect 14299 490 14331 522
<< ndiode >>
rect 906 4212 1002 4244
rect 906 4180 938 4212
rect 970 4180 1002 4212
rect 906 4148 1002 4180
<< ndiodecont >>
rect 938 4180 970 4212
<< metal1 >>
rect 0 4866 16000 4884
rect 0 4834 28 4866
rect 60 4834 96 4866
rect 128 4834 164 4866
rect 196 4834 232 4866
rect 264 4834 300 4866
rect 332 4834 368 4866
rect 400 4834 436 4866
rect 468 4834 504 4866
rect 536 4834 572 4866
rect 604 4834 640 4866
rect 672 4834 708 4866
rect 740 4834 776 4866
rect 808 4834 844 4866
rect 876 4834 912 4866
rect 944 4834 980 4866
rect 1012 4834 1048 4866
rect 1080 4834 1116 4866
rect 1148 4834 1184 4866
rect 1216 4834 1252 4866
rect 1284 4834 1320 4866
rect 1352 4834 1388 4866
rect 1420 4834 1456 4866
rect 1488 4834 1524 4866
rect 1556 4834 1592 4866
rect 1624 4834 1660 4866
rect 1692 4834 1728 4866
rect 1760 4834 1796 4866
rect 1828 4834 1864 4866
rect 1896 4834 1932 4866
rect 1964 4834 2000 4866
rect 2032 4834 2068 4866
rect 2100 4834 2136 4866
rect 2168 4834 2204 4866
rect 2236 4834 2272 4866
rect 2304 4834 2340 4866
rect 2372 4834 2408 4866
rect 2440 4834 2476 4866
rect 2508 4834 2544 4866
rect 2576 4834 2612 4866
rect 2644 4834 2680 4866
rect 2712 4834 2748 4866
rect 2780 4834 2816 4866
rect 2848 4834 2884 4866
rect 2916 4834 2952 4866
rect 2984 4834 3020 4866
rect 3052 4834 3088 4866
rect 3120 4834 3156 4866
rect 3188 4834 3224 4866
rect 3256 4834 3292 4866
rect 3324 4834 3360 4866
rect 3392 4834 3428 4866
rect 3460 4834 3496 4866
rect 3528 4834 3564 4866
rect 3596 4834 3632 4866
rect 3664 4834 3700 4866
rect 3732 4834 3768 4866
rect 3800 4834 3836 4866
rect 3868 4834 3904 4866
rect 3936 4834 3972 4866
rect 4004 4834 4040 4866
rect 4072 4834 4108 4866
rect 4140 4834 4176 4866
rect 4208 4834 4244 4866
rect 4276 4834 4312 4866
rect 4344 4834 4380 4866
rect 4412 4834 4448 4866
rect 4480 4834 4516 4866
rect 4548 4834 4584 4866
rect 4616 4834 4652 4866
rect 4684 4834 4720 4866
rect 4752 4834 4788 4866
rect 4820 4834 4856 4866
rect 4888 4834 4924 4866
rect 4956 4834 4992 4866
rect 5024 4834 5060 4866
rect 5092 4834 5128 4866
rect 5160 4834 5196 4866
rect 5228 4834 5264 4866
rect 5296 4834 5332 4866
rect 5364 4834 5400 4866
rect 5432 4834 5468 4866
rect 5500 4834 5536 4866
rect 5568 4834 5604 4866
rect 5636 4834 5672 4866
rect 5704 4834 5740 4866
rect 5772 4834 5808 4866
rect 5840 4834 5876 4866
rect 5908 4834 5944 4866
rect 5976 4834 6012 4866
rect 6044 4834 6080 4866
rect 6112 4834 6148 4866
rect 6180 4834 6216 4866
rect 6248 4834 6284 4866
rect 6316 4834 6352 4866
rect 6384 4834 6420 4866
rect 6452 4834 6488 4866
rect 6520 4834 6556 4866
rect 6588 4834 6624 4866
rect 6656 4834 6692 4866
rect 6724 4834 6760 4866
rect 6792 4834 6828 4866
rect 6860 4834 6896 4866
rect 6928 4834 6964 4866
rect 6996 4834 7032 4866
rect 7064 4834 7100 4866
rect 7132 4834 7168 4866
rect 7200 4834 7236 4866
rect 7268 4834 7304 4866
rect 7336 4834 7372 4866
rect 7404 4834 7440 4866
rect 7472 4834 7508 4866
rect 7540 4834 7576 4866
rect 7608 4834 7644 4866
rect 7676 4834 7712 4866
rect 7744 4834 7780 4866
rect 7812 4834 7848 4866
rect 7880 4834 7916 4866
rect 7948 4834 7984 4866
rect 8016 4834 8052 4866
rect 8084 4834 8120 4866
rect 8152 4834 8188 4866
rect 8220 4834 8256 4866
rect 8288 4834 8324 4866
rect 8356 4834 8392 4866
rect 8424 4834 8460 4866
rect 8492 4834 8528 4866
rect 8560 4834 8596 4866
rect 8628 4834 8664 4866
rect 8696 4834 8732 4866
rect 8764 4834 8800 4866
rect 8832 4834 8868 4866
rect 8900 4834 8936 4866
rect 8968 4834 9004 4866
rect 9036 4834 9072 4866
rect 9104 4834 9140 4866
rect 9172 4834 9208 4866
rect 9240 4834 9276 4866
rect 9308 4834 9344 4866
rect 9376 4834 9412 4866
rect 9444 4834 9480 4866
rect 9512 4834 9548 4866
rect 9580 4834 9616 4866
rect 9648 4834 9684 4866
rect 9716 4834 9752 4866
rect 9784 4834 9820 4866
rect 9852 4834 9888 4866
rect 9920 4834 9956 4866
rect 9988 4834 10024 4866
rect 10056 4834 10092 4866
rect 10124 4834 10160 4866
rect 10192 4834 10228 4866
rect 10260 4834 10296 4866
rect 10328 4834 10364 4866
rect 10396 4834 10432 4866
rect 10464 4834 10500 4866
rect 10532 4834 10568 4866
rect 10600 4834 10636 4866
rect 10668 4834 10704 4866
rect 10736 4834 10772 4866
rect 10804 4834 10840 4866
rect 10872 4834 10908 4866
rect 10940 4834 10976 4866
rect 11008 4834 11044 4866
rect 11076 4834 11112 4866
rect 11144 4834 11180 4866
rect 11212 4834 11248 4866
rect 11280 4834 11316 4866
rect 11348 4834 11384 4866
rect 11416 4834 11452 4866
rect 11484 4834 11520 4866
rect 11552 4834 11588 4866
rect 11620 4834 11656 4866
rect 11688 4834 11724 4866
rect 11756 4834 11792 4866
rect 11824 4834 11860 4866
rect 11892 4834 11928 4866
rect 11960 4834 11996 4866
rect 12028 4834 12064 4866
rect 12096 4834 12132 4866
rect 12164 4834 12200 4866
rect 12232 4834 12268 4866
rect 12300 4834 12336 4866
rect 12368 4834 12404 4866
rect 12436 4834 12472 4866
rect 12504 4834 12540 4866
rect 12572 4834 12608 4866
rect 12640 4834 12676 4866
rect 12708 4834 12744 4866
rect 12776 4834 12812 4866
rect 12844 4834 12880 4866
rect 12912 4834 12948 4866
rect 12980 4834 13016 4866
rect 13048 4834 13084 4866
rect 13116 4834 13152 4866
rect 13184 4834 13220 4866
rect 13252 4834 13288 4866
rect 13320 4834 13356 4866
rect 13388 4834 13424 4866
rect 13456 4834 13492 4866
rect 13524 4834 13560 4866
rect 13592 4834 13628 4866
rect 13660 4834 13696 4866
rect 13728 4834 13764 4866
rect 13796 4834 13832 4866
rect 13864 4834 13900 4866
rect 13932 4834 13968 4866
rect 14000 4834 14036 4866
rect 14068 4834 14104 4866
rect 14136 4834 14172 4866
rect 14204 4834 14240 4866
rect 14272 4834 14308 4866
rect 14340 4834 14376 4866
rect 14408 4834 14444 4866
rect 14476 4834 14512 4866
rect 14544 4834 14580 4866
rect 14612 4834 14648 4866
rect 14680 4834 14716 4866
rect 14748 4834 14784 4866
rect 14816 4834 14852 4866
rect 14884 4834 14920 4866
rect 14952 4834 14988 4866
rect 15020 4834 15056 4866
rect 15088 4834 15124 4866
rect 15156 4834 15192 4866
rect 15224 4834 15260 4866
rect 15292 4834 15328 4866
rect 15360 4834 15396 4866
rect 15428 4834 15464 4866
rect 15496 4834 15532 4866
rect 15564 4834 15600 4866
rect 15632 4834 15668 4866
rect 15700 4834 15736 4866
rect 15768 4834 15804 4866
rect 15836 4834 15872 4866
rect 15904 4834 15940 4866
rect 15972 4834 16000 4866
rect 0 4816 16000 4834
rect 0 4770 68 4816
rect 0 4738 18 4770
rect 50 4738 68 4770
rect 0 4702 68 4738
rect 0 4670 18 4702
rect 50 4670 68 4702
rect 0 4634 68 4670
rect 0 4602 18 4634
rect 50 4602 68 4634
rect 0 4566 68 4602
rect 0 4534 18 4566
rect 50 4534 68 4566
rect 0 4498 68 4534
rect 15932 4770 16000 4816
rect 15932 4738 15950 4770
rect 15982 4738 16000 4770
rect 15932 4702 16000 4738
rect 15932 4670 15950 4702
rect 15982 4670 16000 4702
rect 15932 4634 16000 4670
rect 15932 4602 15950 4634
rect 15982 4602 16000 4634
rect 15932 4566 16000 4602
rect 15932 4534 15950 4566
rect 15982 4534 16000 4566
rect 0 4466 18 4498
rect 50 4466 68 4498
rect 0 4430 68 4466
rect 0 4398 18 4430
rect 50 4398 68 4430
rect 0 4362 68 4398
rect 0 4330 18 4362
rect 50 4330 68 4362
rect 0 4294 68 4330
rect 0 4262 18 4294
rect 50 4262 68 4294
rect 0 4226 68 4262
rect 0 4194 18 4226
rect 50 4194 68 4226
rect 0 4158 68 4194
rect 0 4126 18 4158
rect 50 4126 68 4158
rect 0 4090 68 4126
rect 0 4058 18 4090
rect 50 4058 68 4090
rect 0 4022 68 4058
rect 0 3990 18 4022
rect 50 3990 68 4022
rect 0 3954 68 3990
rect 0 3922 18 3954
rect 50 3922 68 3954
rect 0 3886 68 3922
rect 0 3854 18 3886
rect 50 3854 68 3886
rect 0 3818 68 3854
rect 0 3786 18 3818
rect 50 3786 68 3818
rect 0 3750 68 3786
rect 0 3718 18 3750
rect 50 3718 68 3750
rect 0 3682 68 3718
rect 0 3650 18 3682
rect 50 3650 68 3682
rect 0 3614 68 3650
rect 0 3582 18 3614
rect 50 3582 68 3614
rect 0 3546 68 3582
rect 0 3514 18 3546
rect 50 3514 68 3546
rect 0 3478 68 3514
rect 0 3446 18 3478
rect 50 3446 68 3478
rect 0 3410 68 3446
rect 0 3378 18 3410
rect 50 3378 68 3410
rect 0 3342 68 3378
rect 0 3310 18 3342
rect 50 3310 68 3342
rect 0 3274 68 3310
rect 0 3242 18 3274
rect 50 3242 68 3274
rect 0 3206 68 3242
rect 0 3174 18 3206
rect 50 3174 68 3206
rect 0 3138 68 3174
rect 0 3106 18 3138
rect 50 3106 68 3138
rect 0 3070 68 3106
rect 0 3038 18 3070
rect 50 3038 68 3070
rect 0 3002 68 3038
rect 0 2970 18 3002
rect 50 2970 68 3002
rect 0 2934 68 2970
rect 0 2902 18 2934
rect 50 2902 68 2934
rect 0 2866 68 2902
rect 0 2834 18 2866
rect 50 2834 68 2866
rect 0 2798 68 2834
rect 0 2766 18 2798
rect 50 2766 68 2798
rect 0 2730 68 2766
rect 0 2698 18 2730
rect 50 2698 68 2730
rect 0 2662 68 2698
rect 0 2630 18 2662
rect 50 2630 68 2662
rect 0 2594 68 2630
rect 0 2562 18 2594
rect 50 2562 68 2594
rect 0 2526 68 2562
rect 0 2494 18 2526
rect 50 2494 68 2526
rect 0 2458 68 2494
rect 0 2426 18 2458
rect 50 2426 68 2458
rect 0 2390 68 2426
rect 0 2358 18 2390
rect 50 2358 68 2390
rect 0 2322 68 2358
rect 0 2290 18 2322
rect 50 2290 68 2322
rect 0 2254 68 2290
rect 0 2222 18 2254
rect 50 2222 68 2254
rect 0 2186 68 2222
rect 0 2154 18 2186
rect 50 2154 68 2186
rect 0 2118 68 2154
rect 0 2086 18 2118
rect 50 2086 68 2118
rect 0 2050 68 2086
rect 0 2018 18 2050
rect 50 2018 68 2050
rect 0 1982 68 2018
rect 0 1950 18 1982
rect 50 1950 68 1982
rect 0 1914 68 1950
rect 0 1882 18 1914
rect 50 1882 68 1914
rect 0 1846 68 1882
rect 0 1814 18 1846
rect 50 1814 68 1846
rect 0 1778 68 1814
rect 0 1746 18 1778
rect 50 1746 68 1778
rect 0 1710 68 1746
rect 0 1678 18 1710
rect 50 1678 68 1710
rect 0 1642 68 1678
rect 0 1610 18 1642
rect 50 1610 68 1642
rect 0 1574 68 1610
rect 0 1542 18 1574
rect 50 1542 68 1574
rect 0 1506 68 1542
rect 0 1474 18 1506
rect 50 1474 68 1506
rect 0 1438 68 1474
rect 0 1406 18 1438
rect 50 1406 68 1438
rect 0 1370 68 1406
rect 0 1338 18 1370
rect 50 1338 68 1370
rect 0 1302 68 1338
rect 0 1270 18 1302
rect 50 1270 68 1302
rect 0 1234 68 1270
rect 0 1202 18 1234
rect 50 1202 68 1234
rect 0 1166 68 1202
rect 0 1134 18 1166
rect 50 1134 68 1166
rect 0 1098 68 1134
rect 0 1066 18 1098
rect 50 1066 68 1098
rect 0 1030 68 1066
rect 0 998 18 1030
rect 50 998 68 1030
rect 0 962 68 998
rect 0 930 18 962
rect 50 930 68 962
rect 0 894 68 930
rect 0 862 18 894
rect 50 862 68 894
rect 0 826 68 862
rect 0 794 18 826
rect 50 794 68 826
rect 0 758 68 794
rect 0 726 18 758
rect 50 726 68 758
rect 0 690 68 726
rect 0 658 18 690
rect 50 658 68 690
rect 0 622 68 658
rect 0 590 18 622
rect 50 590 68 622
rect 0 554 68 590
rect 0 522 18 554
rect 50 522 68 554
rect 0 486 68 522
rect 0 454 18 486
rect 50 454 68 486
rect 0 418 68 454
rect 0 386 18 418
rect 50 386 68 418
rect 0 350 68 386
rect 360 4510 15640 4524
rect 360 4506 1487 4510
rect 1527 4506 2091 4510
rect 2131 4506 2695 4510
rect 2735 4506 3299 4510
rect 3339 4506 3903 4510
rect 3943 4506 4507 4510
rect 4547 4506 5111 4510
rect 5151 4506 5715 4510
rect 5755 4506 6319 4510
rect 6359 4506 6923 4510
rect 6963 4506 7527 4510
rect 7567 4506 8131 4510
rect 8171 4506 8735 4510
rect 8775 4506 9339 4510
rect 9379 4506 9943 4510
rect 9983 4506 10547 4510
rect 10587 4506 11151 4510
rect 11191 4506 11755 4510
rect 11795 4506 12359 4510
rect 12399 4506 12963 4510
rect 13003 4506 13567 4510
rect 13607 4506 14171 4510
rect 14211 4506 15640 4510
rect 360 4474 402 4506
rect 434 4474 470 4506
rect 502 4474 538 4506
rect 570 4474 606 4506
rect 638 4474 674 4506
rect 706 4474 742 4506
rect 774 4474 810 4506
rect 842 4474 878 4506
rect 910 4474 946 4506
rect 978 4474 1014 4506
rect 1046 4474 1082 4506
rect 1114 4474 1150 4506
rect 1182 4474 1218 4506
rect 1250 4474 1286 4506
rect 1318 4474 1354 4506
rect 1386 4474 1422 4506
rect 1454 4474 1487 4506
rect 1527 4474 1558 4506
rect 1590 4474 1626 4506
rect 1658 4474 1694 4506
rect 1726 4474 1762 4506
rect 1794 4474 1830 4506
rect 1862 4474 1898 4506
rect 1930 4474 1966 4506
rect 1998 4474 2034 4506
rect 2066 4474 2091 4506
rect 2134 4474 2170 4506
rect 2202 4474 2238 4506
rect 2270 4474 2306 4506
rect 2338 4474 2374 4506
rect 2406 4474 2442 4506
rect 2474 4474 2510 4506
rect 2542 4474 2578 4506
rect 2610 4474 2646 4506
rect 2678 4474 2695 4506
rect 2746 4474 2782 4506
rect 2814 4474 2850 4506
rect 2882 4474 2918 4506
rect 2950 4474 2986 4506
rect 3018 4474 3054 4506
rect 3086 4474 3122 4506
rect 3154 4474 3190 4506
rect 3222 4474 3258 4506
rect 3290 4474 3299 4506
rect 3358 4474 3394 4506
rect 3426 4474 3462 4506
rect 3494 4474 3530 4506
rect 3562 4474 3598 4506
rect 3630 4474 3666 4506
rect 3698 4474 3734 4506
rect 3766 4474 3802 4506
rect 3834 4474 3870 4506
rect 3902 4474 3903 4506
rect 3970 4474 4006 4506
rect 4038 4474 4074 4506
rect 4106 4474 4142 4506
rect 4174 4474 4210 4506
rect 4242 4474 4278 4506
rect 4310 4474 4346 4506
rect 4378 4474 4414 4506
rect 4446 4474 4482 4506
rect 4547 4474 4550 4506
rect 4582 4474 4618 4506
rect 4650 4474 4686 4506
rect 4718 4474 4754 4506
rect 4786 4474 4822 4506
rect 4854 4474 4890 4506
rect 4922 4474 4958 4506
rect 4990 4474 5026 4506
rect 5058 4474 5094 4506
rect 5151 4474 5162 4506
rect 5194 4474 5230 4506
rect 5262 4474 5298 4506
rect 5330 4474 5366 4506
rect 5398 4474 5434 4506
rect 5466 4474 5502 4506
rect 5534 4474 5570 4506
rect 5602 4474 5638 4506
rect 5670 4474 5706 4506
rect 5755 4474 5774 4506
rect 5806 4474 5842 4506
rect 5874 4474 5910 4506
rect 5942 4474 5978 4506
rect 6010 4474 6046 4506
rect 6078 4474 6114 4506
rect 6146 4474 6182 4506
rect 6214 4474 6250 4506
rect 6282 4474 6318 4506
rect 6359 4474 6386 4506
rect 6418 4474 6454 4506
rect 6486 4474 6522 4506
rect 6554 4474 6590 4506
rect 6622 4474 6658 4506
rect 6690 4474 6726 4506
rect 6758 4474 6794 4506
rect 6826 4474 6862 4506
rect 6894 4474 6923 4506
rect 6963 4474 6998 4506
rect 7030 4474 7066 4506
rect 7098 4474 7134 4506
rect 7166 4474 7202 4506
rect 7234 4474 7270 4506
rect 7302 4474 7338 4506
rect 7370 4474 7406 4506
rect 7438 4474 7474 4506
rect 7506 4474 7527 4506
rect 7574 4474 7610 4506
rect 7642 4474 7678 4506
rect 7710 4474 7746 4506
rect 7778 4474 7814 4506
rect 7846 4474 7882 4506
rect 7914 4474 7950 4506
rect 7982 4474 8018 4506
rect 8050 4474 8086 4506
rect 8118 4474 8131 4506
rect 8186 4474 8222 4506
rect 8254 4474 8290 4506
rect 8322 4474 8358 4506
rect 8390 4474 8426 4506
rect 8458 4474 8494 4506
rect 8526 4474 8562 4506
rect 8594 4474 8630 4506
rect 8662 4474 8698 4506
rect 8730 4474 8735 4506
rect 8798 4474 8834 4506
rect 8866 4474 8902 4506
rect 8934 4474 8970 4506
rect 9002 4474 9038 4506
rect 9070 4474 9106 4506
rect 9138 4474 9174 4506
rect 9206 4474 9242 4506
rect 9274 4474 9310 4506
rect 9410 4474 9446 4506
rect 9478 4474 9514 4506
rect 9546 4474 9582 4506
rect 9614 4474 9650 4506
rect 9682 4474 9718 4506
rect 9750 4474 9786 4506
rect 9818 4474 9854 4506
rect 9886 4474 9922 4506
rect 9983 4474 9990 4506
rect 10022 4474 10058 4506
rect 10090 4474 10126 4506
rect 10158 4474 10194 4506
rect 10226 4474 10262 4506
rect 10294 4474 10330 4506
rect 10362 4474 10398 4506
rect 10430 4474 10466 4506
rect 10498 4474 10534 4506
rect 10587 4474 10602 4506
rect 10634 4474 10670 4506
rect 10702 4474 10738 4506
rect 10770 4474 10806 4506
rect 10838 4474 10874 4506
rect 10906 4474 10942 4506
rect 10974 4474 11010 4506
rect 11042 4474 11078 4506
rect 11110 4474 11146 4506
rect 11191 4474 11214 4506
rect 11246 4474 11282 4506
rect 11314 4474 11350 4506
rect 11382 4474 11418 4506
rect 11450 4474 11486 4506
rect 11518 4474 11554 4506
rect 11586 4474 11622 4506
rect 11654 4474 11690 4506
rect 11722 4474 11755 4506
rect 11795 4474 11826 4506
rect 11858 4474 11894 4506
rect 11926 4474 11962 4506
rect 11994 4474 12030 4506
rect 12062 4474 12098 4506
rect 12130 4474 12166 4506
rect 12198 4474 12234 4506
rect 12266 4474 12302 4506
rect 12334 4474 12359 4506
rect 12402 4474 12438 4506
rect 12470 4474 12506 4506
rect 12538 4474 12574 4506
rect 12606 4474 12642 4506
rect 12674 4474 12710 4506
rect 12742 4474 12778 4506
rect 12810 4474 12846 4506
rect 12878 4474 12914 4506
rect 12946 4474 12963 4506
rect 13014 4474 13050 4506
rect 13082 4474 13118 4506
rect 13150 4474 13186 4506
rect 13218 4474 13254 4506
rect 13286 4474 13322 4506
rect 13354 4474 13390 4506
rect 13422 4474 13458 4506
rect 13490 4474 13526 4506
rect 13558 4474 13567 4506
rect 13626 4474 13662 4506
rect 13694 4474 13730 4506
rect 13762 4474 13798 4506
rect 13830 4474 13866 4506
rect 13898 4474 13934 4506
rect 13966 4474 14002 4506
rect 14034 4474 14070 4506
rect 14102 4474 14138 4506
rect 14170 4474 14171 4506
rect 14238 4474 14274 4506
rect 14306 4474 14342 4506
rect 14374 4474 14410 4506
rect 14442 4474 14478 4506
rect 14510 4474 14546 4506
rect 14578 4474 14614 4506
rect 14646 4474 14682 4506
rect 14714 4474 14750 4506
rect 14782 4474 14818 4506
rect 14850 4474 14886 4506
rect 14918 4474 14954 4506
rect 14986 4474 15022 4506
rect 15054 4474 15090 4506
rect 15122 4474 15158 4506
rect 15190 4474 15226 4506
rect 15258 4474 15294 4506
rect 15326 4474 15362 4506
rect 15394 4474 15430 4506
rect 15462 4474 15498 4506
rect 15530 4474 15566 4506
rect 15598 4474 15640 4506
rect 360 4470 1487 4474
rect 1527 4470 2091 4474
rect 2131 4470 2695 4474
rect 2735 4470 3299 4474
rect 3339 4470 3903 4474
rect 3943 4470 4507 4474
rect 4547 4470 5111 4474
rect 5151 4470 5715 4474
rect 5755 4470 6319 4474
rect 6359 4470 6923 4474
rect 6963 4470 7527 4474
rect 7567 4470 8131 4474
rect 8171 4470 8735 4474
rect 8775 4470 9339 4474
rect 9379 4470 9943 4474
rect 9983 4470 10547 4474
rect 10587 4470 11151 4474
rect 11191 4470 11755 4474
rect 11795 4470 12359 4474
rect 12399 4470 12963 4474
rect 13003 4470 13567 4474
rect 13607 4470 14171 4474
rect 14211 4470 15640 4474
rect 360 4456 15640 4470
rect 360 4396 428 4456
rect 360 4364 378 4396
rect 410 4364 428 4396
rect 360 4328 428 4364
rect 360 4296 378 4328
rect 410 4296 428 4328
rect 360 4260 428 4296
rect 360 4228 378 4260
rect 410 4228 428 4260
rect 360 4192 428 4228
rect 932 4394 14331 4410
rect 932 4378 1615 4394
rect 932 4368 974 4378
rect 932 4246 933 4368
rect 973 4246 974 4368
rect 1647 4378 1971 4394
rect 932 4212 974 4246
rect 1486 4324 1528 4334
rect 360 4160 378 4192
rect 410 4160 428 4192
rect 928 4180 980 4212
rect 360 4124 428 4160
rect 360 4092 378 4124
rect 410 4092 428 4124
rect 360 4056 428 4092
rect 360 4024 378 4056
rect 410 4024 428 4056
rect 360 3988 428 4024
rect 360 3956 378 3988
rect 410 3956 428 3988
rect 360 3920 428 3956
rect 360 3888 378 3920
rect 410 3888 428 3920
rect 360 3852 428 3888
rect 360 3820 378 3852
rect 410 3820 428 3852
rect 360 3784 428 3820
rect 360 3752 378 3784
rect 410 3752 428 3784
rect 360 3716 428 3752
rect 360 3684 378 3716
rect 410 3684 428 3716
rect 360 3648 428 3684
rect 360 3616 378 3648
rect 410 3616 428 3648
rect 360 3580 428 3616
rect 360 3548 378 3580
rect 410 3548 428 3580
rect 360 3512 428 3548
rect 360 3480 378 3512
rect 410 3480 428 3512
rect 360 3444 428 3480
rect 1486 3464 1487 4324
rect 1527 3464 1528 4324
rect 1486 3454 1528 3464
rect 360 3412 378 3444
rect 410 3412 428 3444
rect 360 3376 428 3412
rect 360 3344 378 3376
rect 410 3344 428 3376
rect 1615 3426 1647 4362
rect 2003 4378 2219 4394
rect 1747 4324 1871 4334
rect 1747 3464 1748 4324
rect 1870 3464 1871 4324
rect 1747 3454 1871 3464
rect 360 3308 428 3344
rect 360 3276 378 3308
rect 410 3276 428 3308
rect 360 3240 428 3276
rect 360 3208 378 3240
rect 410 3208 428 3240
rect 360 3172 428 3208
rect 360 3140 378 3172
rect 410 3140 428 3172
rect 360 3104 428 3140
rect 360 3072 378 3104
rect 410 3072 428 3104
rect 360 3036 428 3072
rect 360 3004 378 3036
rect 410 3004 428 3036
rect 360 2968 428 3004
rect 360 2936 378 2968
rect 410 2936 428 2968
rect 360 2900 428 2936
rect 360 2868 378 2900
rect 410 2868 428 2900
rect 360 2832 428 2868
rect 360 2800 378 2832
rect 410 2800 428 2832
rect 360 2764 428 2800
rect 360 2732 378 2764
rect 410 2732 428 2764
rect 360 2696 428 2732
rect 360 2664 378 2696
rect 410 2664 428 2696
rect 360 2628 428 2664
rect 360 2596 378 2628
rect 410 2596 428 2628
rect 360 2560 428 2596
rect 360 2528 378 2560
rect 410 2528 428 2560
rect 360 2492 428 2528
rect 360 2460 378 2492
rect 410 2460 428 2492
rect 1486 3356 1528 3366
rect 1486 2496 1487 3356
rect 1527 2496 1528 3356
rect 1486 2486 1528 2496
rect 360 2424 428 2460
rect 360 2392 378 2424
rect 410 2392 428 2424
rect 1615 2458 1647 3394
rect 1971 3426 2003 4362
rect 2251 4378 2575 4394
rect 2090 4324 2132 4334
rect 2090 3464 2091 4324
rect 2131 3464 2132 4324
rect 2090 3454 2132 3464
rect 1747 3356 1871 3366
rect 1747 2496 1748 3356
rect 1870 2496 1871 3356
rect 1747 2486 1871 2496
rect 360 2356 428 2392
rect 360 2324 378 2356
rect 410 2324 428 2356
rect 360 2288 428 2324
rect 360 2256 378 2288
rect 410 2256 428 2288
rect 360 2220 428 2256
rect 360 2188 378 2220
rect 410 2188 428 2220
rect 360 2152 428 2188
rect 360 2120 378 2152
rect 410 2120 428 2152
rect 360 2084 428 2120
rect 360 2052 378 2084
rect 410 2052 428 2084
rect 360 2016 428 2052
rect 360 1984 378 2016
rect 410 1984 428 2016
rect 360 1948 428 1984
rect 360 1916 378 1948
rect 410 1916 428 1948
rect 360 1880 428 1916
rect 360 1848 378 1880
rect 410 1848 428 1880
rect 360 1812 428 1848
rect 360 1780 378 1812
rect 410 1780 428 1812
rect 360 1744 428 1780
rect 360 1712 378 1744
rect 410 1712 428 1744
rect 360 1676 428 1712
rect 360 1644 378 1676
rect 410 1644 428 1676
rect 360 1608 428 1644
rect 360 1576 378 1608
rect 410 1576 428 1608
rect 360 1540 428 1576
rect 360 1508 378 1540
rect 410 1508 428 1540
rect 1486 2388 1528 2398
rect 1486 1528 1487 2388
rect 1527 1528 1528 2388
rect 1486 1518 1528 1528
rect 360 1472 428 1508
rect 360 1440 378 1472
rect 410 1440 428 1472
rect 360 1404 428 1440
rect 1615 1490 1647 2426
rect 1971 2458 2003 3394
rect 2219 3426 2251 4362
rect 2607 4378 2823 4394
rect 2351 4324 2475 4334
rect 2351 3464 2352 4324
rect 2474 3464 2475 4324
rect 2351 3454 2475 3464
rect 2090 3356 2132 3366
rect 2090 2496 2091 3356
rect 2131 2496 2132 3356
rect 2090 2486 2132 2496
rect 1747 2388 1871 2398
rect 1747 1528 1748 2388
rect 1870 1528 1871 2388
rect 1747 1518 1871 1528
rect 360 1372 378 1404
rect 410 1372 428 1404
rect 360 1336 428 1372
rect 360 1304 378 1336
rect 410 1304 428 1336
rect 360 1268 428 1304
rect 360 1236 378 1268
rect 410 1236 428 1268
rect 360 1200 428 1236
rect 360 1168 378 1200
rect 410 1168 428 1200
rect 360 1132 428 1168
rect 360 1100 378 1132
rect 410 1100 428 1132
rect 360 1064 428 1100
rect 360 1032 378 1064
rect 410 1032 428 1064
rect 360 996 428 1032
rect 360 964 378 996
rect 410 964 428 996
rect 360 928 428 964
rect 360 896 378 928
rect 410 896 428 928
rect 360 860 428 896
rect 360 828 378 860
rect 410 828 428 860
rect 360 792 428 828
rect 360 760 378 792
rect 410 760 428 792
rect 360 724 428 760
rect 360 692 378 724
rect 410 692 428 724
rect 360 656 428 692
rect 360 624 378 656
rect 410 624 428 656
rect 360 588 428 624
rect 360 556 378 588
rect 410 556 428 588
rect 360 520 428 556
rect 1486 1420 1528 1430
rect 1486 560 1487 1420
rect 1527 560 1528 1420
rect 1486 550 1528 560
rect 360 488 378 520
rect 410 488 428 520
rect 360 428 428 488
rect 1615 522 1647 1458
rect 1971 1490 2003 2426
rect 2219 2458 2251 3394
rect 2575 3426 2607 4362
rect 2855 4378 3179 4394
rect 2694 4324 2736 4334
rect 2694 3464 2695 4324
rect 2735 3464 2736 4324
rect 2694 3454 2736 3464
rect 2351 3356 2475 3366
rect 2351 2496 2352 3356
rect 2474 2496 2475 3356
rect 2351 2486 2475 2496
rect 2090 2388 2132 2398
rect 2090 1528 2091 2388
rect 2131 1528 2132 2388
rect 2090 1518 2132 1528
rect 1747 1420 1871 1430
rect 1747 560 1748 1420
rect 1870 560 1871 1420
rect 1747 550 1871 560
rect 1615 474 1647 490
rect 1971 522 2003 1458
rect 2219 1490 2251 2426
rect 2575 2458 2607 3394
rect 2823 3426 2855 4362
rect 3211 4378 3427 4394
rect 2955 4324 3079 4334
rect 2955 3464 2956 4324
rect 3078 3464 3079 4324
rect 2955 3454 3079 3464
rect 2694 3356 2736 3366
rect 2694 2496 2695 3356
rect 2735 2496 2736 3356
rect 2694 2486 2736 2496
rect 2351 2388 2475 2398
rect 2351 1528 2352 2388
rect 2474 1528 2475 2388
rect 2351 1518 2475 1528
rect 2090 1420 2132 1430
rect 2090 560 2091 1420
rect 2131 560 2132 1420
rect 2090 550 2132 560
rect 1971 474 2003 490
rect 2219 522 2251 1458
rect 2575 1490 2607 2426
rect 2823 2458 2855 3394
rect 3179 3426 3211 4362
rect 3459 4378 3783 4394
rect 3298 4324 3340 4334
rect 3298 3464 3299 4324
rect 3339 3464 3340 4324
rect 3298 3454 3340 3464
rect 2955 3356 3079 3366
rect 2955 2496 2956 3356
rect 3078 2496 3079 3356
rect 2955 2486 3079 2496
rect 2694 2388 2736 2398
rect 2694 1528 2695 2388
rect 2735 1528 2736 2388
rect 2694 1518 2736 1528
rect 2351 1420 2475 1430
rect 2351 560 2352 1420
rect 2474 560 2475 1420
rect 2351 550 2475 560
rect 2219 474 2251 490
rect 2575 522 2607 1458
rect 2823 1490 2855 2426
rect 3179 2458 3211 3394
rect 3427 3426 3459 4362
rect 3815 4378 4031 4394
rect 3559 4324 3683 4334
rect 3559 3464 3560 4324
rect 3682 3464 3683 4324
rect 3559 3454 3683 3464
rect 3298 3356 3340 3366
rect 3298 2496 3299 3356
rect 3339 2496 3340 3356
rect 3298 2486 3340 2496
rect 2955 2388 3079 2398
rect 2955 1528 2956 2388
rect 3078 1528 3079 2388
rect 2955 1518 3079 1528
rect 2694 1420 2736 1430
rect 2694 560 2695 1420
rect 2735 560 2736 1420
rect 2694 550 2736 560
rect 2575 474 2607 490
rect 2823 522 2855 1458
rect 3179 1490 3211 2426
rect 3427 2458 3459 3394
rect 3783 3426 3815 4362
rect 4063 4378 4387 4394
rect 3902 4324 3944 4334
rect 3902 3464 3903 4324
rect 3943 3464 3944 4324
rect 3902 3454 3944 3464
rect 3559 3356 3683 3366
rect 3559 2496 3560 3356
rect 3682 2496 3683 3356
rect 3559 2486 3683 2496
rect 3298 2388 3340 2398
rect 3298 1528 3299 2388
rect 3339 1528 3340 2388
rect 3298 1518 3340 1528
rect 2955 1420 3079 1430
rect 2955 560 2956 1420
rect 3078 560 3079 1420
rect 2955 550 3079 560
rect 2823 474 2855 490
rect 3179 522 3211 1458
rect 3427 1490 3459 2426
rect 3783 2458 3815 3394
rect 4031 3426 4063 4362
rect 4419 4378 4635 4394
rect 4163 4324 4287 4334
rect 4163 3464 4164 4324
rect 4286 3464 4287 4324
rect 4163 3454 4287 3464
rect 3902 3356 3944 3366
rect 3902 2496 3903 3356
rect 3943 2496 3944 3356
rect 3902 2486 3944 2496
rect 3559 2388 3683 2398
rect 3559 1528 3560 2388
rect 3682 1528 3683 2388
rect 3559 1518 3683 1528
rect 3298 1420 3340 1430
rect 3298 560 3299 1420
rect 3339 560 3340 1420
rect 3298 550 3340 560
rect 3179 474 3211 490
rect 3427 522 3459 1458
rect 3783 1490 3815 2426
rect 4031 2458 4063 3394
rect 4387 3426 4419 4362
rect 4667 4378 4991 4394
rect 4506 4324 4548 4334
rect 4506 3464 4507 4324
rect 4547 3464 4548 4324
rect 4506 3454 4548 3464
rect 4163 3356 4287 3366
rect 4163 2496 4164 3356
rect 4286 2496 4287 3356
rect 4163 2486 4287 2496
rect 3902 2388 3944 2398
rect 3902 1528 3903 2388
rect 3943 1528 3944 2388
rect 3902 1518 3944 1528
rect 3559 1420 3683 1430
rect 3559 560 3560 1420
rect 3682 560 3683 1420
rect 3559 550 3683 560
rect 3427 474 3459 490
rect 3783 522 3815 1458
rect 4031 1490 4063 2426
rect 4387 2458 4419 3394
rect 4635 3426 4667 4362
rect 5023 4378 5239 4394
rect 4767 4324 4891 4334
rect 4767 3464 4768 4324
rect 4890 3464 4891 4324
rect 4767 3454 4891 3464
rect 4506 3356 4548 3366
rect 4506 2496 4507 3356
rect 4547 2496 4548 3356
rect 4506 2486 4548 2496
rect 4163 2388 4287 2398
rect 4163 1528 4164 2388
rect 4286 1528 4287 2388
rect 4163 1518 4287 1528
rect 3902 1420 3944 1430
rect 3902 560 3903 1420
rect 3943 560 3944 1420
rect 3902 550 3944 560
rect 3783 474 3815 490
rect 4031 522 4063 1458
rect 4387 1490 4419 2426
rect 4635 2458 4667 3394
rect 4991 3426 5023 4362
rect 5271 4378 5595 4394
rect 5110 4324 5152 4334
rect 5110 3464 5111 4324
rect 5151 3464 5152 4324
rect 5110 3454 5152 3464
rect 4767 3356 4891 3366
rect 4767 2496 4768 3356
rect 4890 2496 4891 3356
rect 4767 2486 4891 2496
rect 4506 2388 4548 2398
rect 4506 1528 4507 2388
rect 4547 1528 4548 2388
rect 4506 1518 4548 1528
rect 4163 1420 4287 1430
rect 4163 560 4164 1420
rect 4286 560 4287 1420
rect 4163 550 4287 560
rect 4031 474 4063 490
rect 4387 522 4419 1458
rect 4635 1490 4667 2426
rect 4991 2458 5023 3394
rect 5239 3426 5271 4362
rect 5627 4378 5843 4394
rect 5371 4324 5495 4334
rect 5371 3464 5372 4324
rect 5494 3464 5495 4324
rect 5371 3454 5495 3464
rect 5110 3356 5152 3366
rect 5110 2496 5111 3356
rect 5151 2496 5152 3356
rect 5110 2486 5152 2496
rect 4767 2388 4891 2398
rect 4767 1528 4768 2388
rect 4890 1528 4891 2388
rect 4767 1518 4891 1528
rect 4506 1420 4548 1430
rect 4506 560 4507 1420
rect 4547 560 4548 1420
rect 4506 550 4548 560
rect 4387 474 4419 490
rect 4635 522 4667 1458
rect 4991 1490 5023 2426
rect 5239 2458 5271 3394
rect 5595 3426 5627 4362
rect 5875 4378 6199 4394
rect 5714 4324 5756 4334
rect 5714 3464 5715 4324
rect 5755 3464 5756 4324
rect 5714 3454 5756 3464
rect 5371 3356 5495 3366
rect 5371 2496 5372 3356
rect 5494 2496 5495 3356
rect 5371 2486 5495 2496
rect 5110 2388 5152 2398
rect 5110 1528 5111 2388
rect 5151 1528 5152 2388
rect 5110 1518 5152 1528
rect 4767 1420 4891 1430
rect 4767 560 4768 1420
rect 4890 560 4891 1420
rect 4767 550 4891 560
rect 4635 474 4667 490
rect 4991 522 5023 1458
rect 5239 1490 5271 2426
rect 5595 2458 5627 3394
rect 5843 3426 5875 4362
rect 6231 4378 6447 4394
rect 5975 4324 6099 4334
rect 5975 3464 5976 4324
rect 6098 3464 6099 4324
rect 5975 3454 6099 3464
rect 5714 3356 5756 3366
rect 5714 2496 5715 3356
rect 5755 2496 5756 3356
rect 5714 2486 5756 2496
rect 5371 2388 5495 2398
rect 5371 1528 5372 2388
rect 5494 1528 5495 2388
rect 5371 1518 5495 1528
rect 5110 1420 5152 1430
rect 5110 560 5111 1420
rect 5151 560 5152 1420
rect 5110 550 5152 560
rect 4991 474 5023 490
rect 5239 522 5271 1458
rect 5595 1490 5627 2426
rect 5843 2458 5875 3394
rect 6199 3426 6231 4362
rect 6479 4378 6803 4394
rect 6318 4324 6360 4334
rect 6318 3464 6319 4324
rect 6359 3464 6360 4324
rect 6318 3454 6360 3464
rect 5975 3356 6099 3366
rect 5975 2496 5976 3356
rect 6098 2496 6099 3356
rect 5975 2486 6099 2496
rect 5714 2388 5756 2398
rect 5714 1528 5715 2388
rect 5755 1528 5756 2388
rect 5714 1518 5756 1528
rect 5371 1420 5495 1430
rect 5371 560 5372 1420
rect 5494 560 5495 1420
rect 5371 550 5495 560
rect 5239 474 5271 490
rect 5595 522 5627 1458
rect 5843 1490 5875 2426
rect 6199 2458 6231 3394
rect 6447 3426 6479 4362
rect 6835 4378 7051 4394
rect 6579 4324 6703 4334
rect 6579 3464 6580 4324
rect 6702 3464 6703 4324
rect 6579 3454 6703 3464
rect 6318 3356 6360 3366
rect 6318 2496 6319 3356
rect 6359 2496 6360 3356
rect 6318 2486 6360 2496
rect 5975 2388 6099 2398
rect 5975 1528 5976 2388
rect 6098 1528 6099 2388
rect 5975 1518 6099 1528
rect 5714 1420 5756 1430
rect 5714 560 5715 1420
rect 5755 560 5756 1420
rect 5714 550 5756 560
rect 5595 474 5627 490
rect 5843 522 5875 1458
rect 6199 1490 6231 2426
rect 6447 2458 6479 3394
rect 6803 3426 6835 4362
rect 7083 4378 7407 4394
rect 6922 4324 6964 4334
rect 6922 3464 6923 4324
rect 6963 3464 6964 4324
rect 6922 3454 6964 3464
rect 6579 3356 6703 3366
rect 6579 2496 6580 3356
rect 6702 2496 6703 3356
rect 6579 2486 6703 2496
rect 6318 2388 6360 2398
rect 6318 1528 6319 2388
rect 6359 1528 6360 2388
rect 6318 1518 6360 1528
rect 5975 1420 6099 1430
rect 5975 560 5976 1420
rect 6098 560 6099 1420
rect 5975 550 6099 560
rect 5843 474 5875 490
rect 6199 522 6231 1458
rect 6447 1490 6479 2426
rect 6803 2458 6835 3394
rect 7051 3426 7083 4362
rect 7439 4378 7655 4394
rect 7183 4324 7307 4334
rect 7183 3464 7184 4324
rect 7306 3464 7307 4324
rect 7183 3454 7307 3464
rect 6922 3356 6964 3366
rect 6922 2496 6923 3356
rect 6963 2496 6964 3356
rect 6922 2486 6964 2496
rect 6579 2388 6703 2398
rect 6579 1528 6580 2388
rect 6702 1528 6703 2388
rect 6579 1518 6703 1528
rect 6318 1420 6360 1430
rect 6318 560 6319 1420
rect 6359 560 6360 1420
rect 6318 550 6360 560
rect 6199 474 6231 490
rect 6447 522 6479 1458
rect 6803 1490 6835 2426
rect 7051 2458 7083 3394
rect 7407 3426 7439 4362
rect 7687 4378 8011 4394
rect 7526 4324 7568 4334
rect 7526 3464 7527 4324
rect 7567 3464 7568 4324
rect 7526 3454 7568 3464
rect 7183 3356 7307 3366
rect 7183 2496 7184 3356
rect 7306 2496 7307 3356
rect 7183 2486 7307 2496
rect 6922 2388 6964 2398
rect 6922 1528 6923 2388
rect 6963 1528 6964 2388
rect 6922 1518 6964 1528
rect 6579 1420 6703 1430
rect 6579 560 6580 1420
rect 6702 560 6703 1420
rect 6579 550 6703 560
rect 6447 474 6479 490
rect 6803 522 6835 1458
rect 7051 1490 7083 2426
rect 7407 2458 7439 3394
rect 7655 3426 7687 4362
rect 8043 4378 8259 4394
rect 7787 4324 7911 4334
rect 7787 3464 7788 4324
rect 7910 3464 7911 4324
rect 7787 3454 7911 3464
rect 7526 3356 7568 3366
rect 7526 2496 7527 3356
rect 7567 2496 7568 3356
rect 7526 2486 7568 2496
rect 7183 2388 7307 2398
rect 7183 1528 7184 2388
rect 7306 1528 7307 2388
rect 7183 1518 7307 1528
rect 6922 1420 6964 1430
rect 6922 560 6923 1420
rect 6963 560 6964 1420
rect 6922 550 6964 560
rect 6803 474 6835 490
rect 7051 522 7083 1458
rect 7407 1490 7439 2426
rect 7655 2458 7687 3394
rect 8011 3426 8043 4362
rect 8291 4378 8615 4394
rect 8130 4324 8172 4334
rect 8130 3464 8131 4324
rect 8171 3464 8172 4324
rect 8130 3454 8172 3464
rect 7787 3356 7911 3366
rect 7787 2496 7788 3356
rect 7910 2496 7911 3356
rect 7787 2486 7911 2496
rect 7526 2388 7568 2398
rect 7526 1528 7527 2388
rect 7567 1528 7568 2388
rect 7526 1518 7568 1528
rect 7183 1420 7307 1430
rect 7183 560 7184 1420
rect 7306 560 7307 1420
rect 7183 550 7307 560
rect 7051 474 7083 490
rect 7407 522 7439 1458
rect 7655 1490 7687 2426
rect 8011 2458 8043 3394
rect 8259 3426 8291 4362
rect 8647 4378 8863 4394
rect 8391 4324 8515 4334
rect 8391 3464 8392 4324
rect 8514 3464 8515 4324
rect 8391 3454 8515 3464
rect 8130 3356 8172 3366
rect 8130 2496 8131 3356
rect 8171 2496 8172 3356
rect 8130 2486 8172 2496
rect 7787 2388 7911 2398
rect 7787 1528 7788 2388
rect 7910 1528 7911 2388
rect 7787 1518 7911 1528
rect 7526 1420 7568 1430
rect 7526 560 7527 1420
rect 7567 560 7568 1420
rect 7526 550 7568 560
rect 7407 474 7439 490
rect 7655 522 7687 1458
rect 8011 1490 8043 2426
rect 8259 2458 8291 3394
rect 8615 3426 8647 4362
rect 8895 4378 9219 4394
rect 8734 4324 8776 4334
rect 8734 3464 8735 4324
rect 8775 3464 8776 4324
rect 8734 3454 8776 3464
rect 8391 3356 8515 3366
rect 8391 2496 8392 3356
rect 8514 2496 8515 3356
rect 8391 2486 8515 2496
rect 8130 2388 8172 2398
rect 8130 1528 8131 2388
rect 8171 1528 8172 2388
rect 8130 1518 8172 1528
rect 7787 1420 7911 1430
rect 7787 560 7788 1420
rect 7910 560 7911 1420
rect 7787 550 7911 560
rect 7655 474 7687 490
rect 8011 522 8043 1458
rect 8259 1490 8291 2426
rect 8615 2458 8647 3394
rect 8863 3426 8895 4362
rect 9251 4378 9467 4394
rect 8995 4324 9119 4334
rect 8995 3464 8996 4324
rect 9118 3464 9119 4324
rect 8995 3454 9119 3464
rect 8734 3356 8776 3366
rect 8734 2496 8735 3356
rect 8775 2496 8776 3356
rect 8734 2486 8776 2496
rect 8391 2388 8515 2398
rect 8391 1528 8392 2388
rect 8514 1528 8515 2388
rect 8391 1518 8515 1528
rect 8130 1420 8172 1430
rect 8130 560 8131 1420
rect 8171 560 8172 1420
rect 8130 550 8172 560
rect 8011 474 8043 490
rect 8259 522 8291 1458
rect 8615 1490 8647 2426
rect 8863 2458 8895 3394
rect 9219 3426 9251 4362
rect 9499 4378 9823 4394
rect 9338 4324 9380 4334
rect 9338 3464 9339 4324
rect 9379 3464 9380 4324
rect 9338 3454 9380 3464
rect 8995 3356 9119 3366
rect 8995 2496 8996 3356
rect 9118 2496 9119 3356
rect 8995 2486 9119 2496
rect 8734 2388 8776 2398
rect 8734 1528 8735 2388
rect 8775 1528 8776 2388
rect 8734 1518 8776 1528
rect 8391 1420 8515 1430
rect 8391 560 8392 1420
rect 8514 560 8515 1420
rect 8391 550 8515 560
rect 8259 474 8291 490
rect 8615 522 8647 1458
rect 8863 1490 8895 2426
rect 9219 2458 9251 3394
rect 9467 3426 9499 4362
rect 9855 4378 10071 4394
rect 9599 4324 9723 4334
rect 9599 3464 9600 4324
rect 9722 3464 9723 4324
rect 9599 3454 9723 3464
rect 9338 3356 9380 3366
rect 9338 2496 9339 3356
rect 9379 2496 9380 3356
rect 9338 2486 9380 2496
rect 8995 2388 9119 2398
rect 8995 1528 8996 2388
rect 9118 1528 9119 2388
rect 8995 1518 9119 1528
rect 8734 1420 8776 1430
rect 8734 560 8735 1420
rect 8775 560 8776 1420
rect 8734 550 8776 560
rect 8615 474 8647 490
rect 8863 522 8895 1458
rect 9219 1490 9251 2426
rect 9467 2458 9499 3394
rect 9823 3426 9855 4362
rect 10103 4378 10427 4394
rect 9942 4324 9984 4334
rect 9942 3464 9943 4324
rect 9983 3464 9984 4324
rect 9942 3454 9984 3464
rect 9599 3356 9723 3366
rect 9599 2496 9600 3356
rect 9722 2496 9723 3356
rect 9599 2486 9723 2496
rect 9338 2388 9380 2398
rect 9338 1528 9339 2388
rect 9379 1528 9380 2388
rect 9338 1518 9380 1528
rect 8995 1420 9119 1430
rect 8995 560 8996 1420
rect 9118 560 9119 1420
rect 8995 550 9119 560
rect 8863 474 8895 490
rect 9219 522 9251 1458
rect 9467 1490 9499 2426
rect 9823 2458 9855 3394
rect 10071 3426 10103 4362
rect 10459 4378 10675 4394
rect 10203 4324 10327 4334
rect 10203 3464 10204 4324
rect 10326 3464 10327 4324
rect 10203 3454 10327 3464
rect 9942 3356 9984 3366
rect 9942 2496 9943 3356
rect 9983 2496 9984 3356
rect 9942 2486 9984 2496
rect 9599 2388 9723 2398
rect 9599 1528 9600 2388
rect 9722 1528 9723 2388
rect 9599 1518 9723 1528
rect 9338 1420 9380 1430
rect 9338 560 9339 1420
rect 9379 560 9380 1420
rect 9338 550 9380 560
rect 9219 474 9251 490
rect 9467 522 9499 1458
rect 9823 1490 9855 2426
rect 10071 2458 10103 3394
rect 10427 3426 10459 4362
rect 10707 4378 11031 4394
rect 10546 4324 10588 4334
rect 10546 3464 10547 4324
rect 10587 3464 10588 4324
rect 10546 3454 10588 3464
rect 10203 3356 10327 3366
rect 10203 2496 10204 3356
rect 10326 2496 10327 3356
rect 10203 2486 10327 2496
rect 9942 2388 9984 2398
rect 9942 1528 9943 2388
rect 9983 1528 9984 2388
rect 9942 1518 9984 1528
rect 9599 1420 9723 1430
rect 9599 560 9600 1420
rect 9722 560 9723 1420
rect 9599 550 9723 560
rect 9467 474 9499 490
rect 9823 522 9855 1458
rect 10071 1490 10103 2426
rect 10427 2458 10459 3394
rect 10675 3426 10707 4362
rect 11063 4378 11279 4394
rect 10807 4324 10931 4334
rect 10807 3464 10808 4324
rect 10930 3464 10931 4324
rect 10807 3454 10931 3464
rect 10546 3356 10588 3366
rect 10546 2496 10547 3356
rect 10587 2496 10588 3356
rect 10546 2486 10588 2496
rect 10203 2388 10327 2398
rect 10203 1528 10204 2388
rect 10326 1528 10327 2388
rect 10203 1518 10327 1528
rect 9942 1420 9984 1430
rect 9942 560 9943 1420
rect 9983 560 9984 1420
rect 9942 550 9984 560
rect 9823 474 9855 490
rect 10071 522 10103 1458
rect 10427 1490 10459 2426
rect 10675 2458 10707 3394
rect 11031 3426 11063 4362
rect 11311 4378 11635 4394
rect 11150 4324 11192 4334
rect 11150 3464 11151 4324
rect 11191 3464 11192 4324
rect 11150 3454 11192 3464
rect 10807 3356 10931 3366
rect 10807 2496 10808 3356
rect 10930 2496 10931 3356
rect 10807 2486 10931 2496
rect 10546 2388 10588 2398
rect 10546 1528 10547 2388
rect 10587 1528 10588 2388
rect 10546 1518 10588 1528
rect 10203 1420 10327 1430
rect 10203 560 10204 1420
rect 10326 560 10327 1420
rect 10203 550 10327 560
rect 10071 474 10103 490
rect 10427 522 10459 1458
rect 10675 1490 10707 2426
rect 11031 2458 11063 3394
rect 11279 3426 11311 4362
rect 11667 4378 11883 4394
rect 11411 4324 11535 4334
rect 11411 3464 11412 4324
rect 11534 3464 11535 4324
rect 11411 3454 11535 3464
rect 11150 3356 11192 3366
rect 11150 2496 11151 3356
rect 11191 2496 11192 3356
rect 11150 2486 11192 2496
rect 10807 2388 10931 2398
rect 10807 1528 10808 2388
rect 10930 1528 10931 2388
rect 10807 1518 10931 1528
rect 10546 1420 10588 1430
rect 10546 560 10547 1420
rect 10587 560 10588 1420
rect 10546 550 10588 560
rect 10427 474 10459 490
rect 10675 522 10707 1458
rect 11031 1490 11063 2426
rect 11279 2458 11311 3394
rect 11635 3426 11667 4362
rect 11915 4378 12239 4394
rect 11754 4324 11796 4334
rect 11754 3464 11755 4324
rect 11795 3464 11796 4324
rect 11754 3454 11796 3464
rect 11411 3356 11535 3366
rect 11411 2496 11412 3356
rect 11534 2496 11535 3356
rect 11411 2486 11535 2496
rect 11150 2388 11192 2398
rect 11150 1528 11151 2388
rect 11191 1528 11192 2388
rect 11150 1518 11192 1528
rect 10807 1420 10931 1430
rect 10807 560 10808 1420
rect 10930 560 10931 1420
rect 10807 550 10931 560
rect 10675 474 10707 490
rect 11031 522 11063 1458
rect 11279 1490 11311 2426
rect 11635 2458 11667 3394
rect 11883 3426 11915 4362
rect 12271 4378 12487 4394
rect 12015 4324 12139 4334
rect 12015 3464 12016 4324
rect 12138 3464 12139 4324
rect 12015 3454 12139 3464
rect 11754 3356 11796 3366
rect 11754 2496 11755 3356
rect 11795 2496 11796 3356
rect 11754 2486 11796 2496
rect 11411 2388 11535 2398
rect 11411 1528 11412 2388
rect 11534 1528 11535 2388
rect 11411 1518 11535 1528
rect 11150 1420 11192 1430
rect 11150 560 11151 1420
rect 11191 560 11192 1420
rect 11150 550 11192 560
rect 11031 474 11063 490
rect 11279 522 11311 1458
rect 11635 1490 11667 2426
rect 11883 2458 11915 3394
rect 12239 3426 12271 4362
rect 12519 4378 12843 4394
rect 12358 4324 12400 4334
rect 12358 3464 12359 4324
rect 12399 3464 12400 4324
rect 12358 3454 12400 3464
rect 12015 3356 12139 3366
rect 12015 2496 12016 3356
rect 12138 2496 12139 3356
rect 12015 2486 12139 2496
rect 11754 2388 11796 2398
rect 11754 1528 11755 2388
rect 11795 1528 11796 2388
rect 11754 1518 11796 1528
rect 11411 1420 11535 1430
rect 11411 560 11412 1420
rect 11534 560 11535 1420
rect 11411 550 11535 560
rect 11279 474 11311 490
rect 11635 522 11667 1458
rect 11883 1490 11915 2426
rect 12239 2458 12271 3394
rect 12487 3426 12519 4362
rect 12875 4378 13091 4394
rect 12619 4324 12743 4334
rect 12619 3464 12620 4324
rect 12742 3464 12743 4324
rect 12619 3454 12743 3464
rect 12358 3356 12400 3366
rect 12358 2496 12359 3356
rect 12399 2496 12400 3356
rect 12358 2486 12400 2496
rect 12015 2388 12139 2398
rect 12015 1528 12016 2388
rect 12138 1528 12139 2388
rect 12015 1518 12139 1528
rect 11754 1420 11796 1430
rect 11754 560 11755 1420
rect 11795 560 11796 1420
rect 11754 550 11796 560
rect 11635 474 11667 490
rect 11883 522 11915 1458
rect 12239 1490 12271 2426
rect 12487 2458 12519 3394
rect 12843 3426 12875 4362
rect 13123 4378 13447 4394
rect 12962 4324 13004 4334
rect 12962 3464 12963 4324
rect 13003 3464 13004 4324
rect 12962 3454 13004 3464
rect 12619 3356 12743 3366
rect 12619 2496 12620 3356
rect 12742 2496 12743 3356
rect 12619 2486 12743 2496
rect 12358 2388 12400 2398
rect 12358 1528 12359 2388
rect 12399 1528 12400 2388
rect 12358 1518 12400 1528
rect 12015 1420 12139 1430
rect 12015 560 12016 1420
rect 12138 560 12139 1420
rect 12015 550 12139 560
rect 11883 474 11915 490
rect 12239 522 12271 1458
rect 12487 1490 12519 2426
rect 12843 2458 12875 3394
rect 13091 3426 13123 4362
rect 13479 4378 13695 4394
rect 13223 4324 13347 4334
rect 13223 3464 13224 4324
rect 13346 3464 13347 4324
rect 13223 3454 13347 3464
rect 12962 3356 13004 3366
rect 12962 2496 12963 3356
rect 13003 2496 13004 3356
rect 12962 2486 13004 2496
rect 12619 2388 12743 2398
rect 12619 1528 12620 2388
rect 12742 1528 12743 2388
rect 12619 1518 12743 1528
rect 12358 1420 12400 1430
rect 12358 560 12359 1420
rect 12399 560 12400 1420
rect 12358 550 12400 560
rect 12239 474 12271 490
rect 12487 522 12519 1458
rect 12843 1490 12875 2426
rect 13091 2458 13123 3394
rect 13447 3426 13479 4362
rect 13727 4378 14051 4394
rect 13566 4324 13608 4334
rect 13566 3464 13567 4324
rect 13607 3464 13608 4324
rect 13566 3454 13608 3464
rect 13223 3356 13347 3366
rect 13223 2496 13224 3356
rect 13346 2496 13347 3356
rect 13223 2486 13347 2496
rect 12962 2388 13004 2398
rect 12962 1528 12963 2388
rect 13003 1528 13004 2388
rect 12962 1518 13004 1528
rect 12619 1420 12743 1430
rect 12619 560 12620 1420
rect 12742 560 12743 1420
rect 12619 550 12743 560
rect 12487 474 12519 490
rect 12843 522 12875 1458
rect 13091 1490 13123 2426
rect 13447 2458 13479 3394
rect 13695 3426 13727 4362
rect 14083 4378 14299 4394
rect 13827 4324 13951 4334
rect 13827 3464 13828 4324
rect 13950 3464 13951 4324
rect 13827 3454 13951 3464
rect 13566 3356 13608 3366
rect 13566 2496 13567 3356
rect 13607 2496 13608 3356
rect 13566 2486 13608 2496
rect 13223 2388 13347 2398
rect 13223 1528 13224 2388
rect 13346 1528 13347 2388
rect 13223 1518 13347 1528
rect 12962 1420 13004 1430
rect 12962 560 12963 1420
rect 13003 560 13004 1420
rect 12962 550 13004 560
rect 12843 474 12875 490
rect 13091 522 13123 1458
rect 13447 1490 13479 2426
rect 13695 2458 13727 3394
rect 14051 3426 14083 4362
rect 14170 4324 14212 4334
rect 14170 3464 14171 4324
rect 14211 3464 14212 4324
rect 14170 3454 14212 3464
rect 13827 3356 13951 3366
rect 13827 2496 13828 3356
rect 13950 2496 13951 3356
rect 13827 2486 13951 2496
rect 13566 2388 13608 2398
rect 13566 1528 13567 2388
rect 13607 1528 13608 2388
rect 13566 1518 13608 1528
rect 13223 1420 13347 1430
rect 13223 560 13224 1420
rect 13346 560 13347 1420
rect 13223 550 13347 560
rect 13091 474 13123 490
rect 13447 522 13479 1458
rect 13695 1490 13727 2426
rect 14051 2458 14083 3394
rect 14299 3426 14331 4362
rect 15572 4396 15640 4456
rect 15572 4364 15590 4396
rect 15622 4364 15640 4396
rect 14431 4324 14555 4334
rect 14431 3464 14432 4324
rect 14554 3464 14555 4324
rect 14431 3454 14555 3464
rect 15572 4328 15640 4364
rect 15572 4296 15590 4328
rect 15622 4296 15640 4328
rect 15572 4260 15640 4296
rect 15572 4228 15590 4260
rect 15622 4228 15640 4260
rect 15572 4192 15640 4228
rect 15572 4160 15590 4192
rect 15622 4160 15640 4192
rect 15572 4124 15640 4160
rect 15572 4092 15590 4124
rect 15622 4092 15640 4124
rect 15572 4056 15640 4092
rect 15572 4024 15590 4056
rect 15622 4024 15640 4056
rect 15572 3988 15640 4024
rect 15572 3956 15590 3988
rect 15622 3956 15640 3988
rect 15572 3920 15640 3956
rect 15572 3888 15590 3920
rect 15622 3888 15640 3920
rect 15572 3852 15640 3888
rect 15572 3820 15590 3852
rect 15622 3820 15640 3852
rect 15572 3784 15640 3820
rect 15572 3752 15590 3784
rect 15622 3752 15640 3784
rect 15572 3716 15640 3752
rect 15572 3684 15590 3716
rect 15622 3684 15640 3716
rect 15572 3648 15640 3684
rect 15572 3616 15590 3648
rect 15622 3616 15640 3648
rect 15572 3580 15640 3616
rect 15572 3548 15590 3580
rect 15622 3548 15640 3580
rect 15572 3512 15640 3548
rect 15572 3480 15590 3512
rect 15622 3480 15640 3512
rect 14170 3356 14212 3366
rect 14170 2496 14171 3356
rect 14211 2496 14212 3356
rect 14170 2486 14212 2496
rect 13827 2388 13951 2398
rect 13827 1528 13828 2388
rect 13950 1528 13951 2388
rect 13827 1518 13951 1528
rect 13566 1420 13608 1430
rect 13566 560 13567 1420
rect 13607 560 13608 1420
rect 13566 550 13608 560
rect 13447 474 13479 490
rect 13695 522 13727 1458
rect 14051 1490 14083 2426
rect 14299 2458 14331 3394
rect 15572 3444 15640 3480
rect 15572 3412 15590 3444
rect 15622 3412 15640 3444
rect 15572 3376 15640 3412
rect 14431 3356 14555 3366
rect 14431 2496 14432 3356
rect 14554 2496 14555 3356
rect 14431 2486 14555 2496
rect 15572 3344 15590 3376
rect 15622 3344 15640 3376
rect 15572 3308 15640 3344
rect 15572 3276 15590 3308
rect 15622 3276 15640 3308
rect 15572 3240 15640 3276
rect 15572 3208 15590 3240
rect 15622 3208 15640 3240
rect 15572 3172 15640 3208
rect 15572 3140 15590 3172
rect 15622 3140 15640 3172
rect 15572 3104 15640 3140
rect 15572 3072 15590 3104
rect 15622 3072 15640 3104
rect 15572 3036 15640 3072
rect 15572 3004 15590 3036
rect 15622 3004 15640 3036
rect 15572 2968 15640 3004
rect 15572 2936 15590 2968
rect 15622 2936 15640 2968
rect 15572 2900 15640 2936
rect 15572 2868 15590 2900
rect 15622 2868 15640 2900
rect 15572 2832 15640 2868
rect 15572 2800 15590 2832
rect 15622 2800 15640 2832
rect 15572 2764 15640 2800
rect 15572 2732 15590 2764
rect 15622 2732 15640 2764
rect 15572 2696 15640 2732
rect 15572 2664 15590 2696
rect 15622 2664 15640 2696
rect 15572 2628 15640 2664
rect 15572 2596 15590 2628
rect 15622 2596 15640 2628
rect 15572 2560 15640 2596
rect 15572 2528 15590 2560
rect 15622 2528 15640 2560
rect 15572 2492 15640 2528
rect 14170 2388 14212 2398
rect 14170 1528 14171 2388
rect 14211 1528 14212 2388
rect 14170 1518 14212 1528
rect 13827 1420 13951 1430
rect 13827 560 13828 1420
rect 13950 560 13951 1420
rect 13827 550 13951 560
rect 13695 474 13727 490
rect 14051 522 14083 1458
rect 14299 1490 14331 2426
rect 15572 2460 15590 2492
rect 15622 2460 15640 2492
rect 15572 2424 15640 2460
rect 14431 2388 14555 2398
rect 14431 1528 14432 2388
rect 14554 1528 14555 2388
rect 14431 1518 14555 1528
rect 15572 2392 15590 2424
rect 15622 2392 15640 2424
rect 15572 2356 15640 2392
rect 15572 2324 15590 2356
rect 15622 2324 15640 2356
rect 15572 2288 15640 2324
rect 15572 2256 15590 2288
rect 15622 2256 15640 2288
rect 15572 2220 15640 2256
rect 15572 2188 15590 2220
rect 15622 2188 15640 2220
rect 15572 2152 15640 2188
rect 15572 2120 15590 2152
rect 15622 2120 15640 2152
rect 15572 2084 15640 2120
rect 15572 2052 15590 2084
rect 15622 2052 15640 2084
rect 15572 2016 15640 2052
rect 15572 1984 15590 2016
rect 15622 1984 15640 2016
rect 15572 1948 15640 1984
rect 15572 1916 15590 1948
rect 15622 1916 15640 1948
rect 15572 1880 15640 1916
rect 15572 1848 15590 1880
rect 15622 1848 15640 1880
rect 15572 1812 15640 1848
rect 15572 1780 15590 1812
rect 15622 1780 15640 1812
rect 15572 1744 15640 1780
rect 15572 1712 15590 1744
rect 15622 1712 15640 1744
rect 15572 1676 15640 1712
rect 15572 1644 15590 1676
rect 15622 1644 15640 1676
rect 15572 1608 15640 1644
rect 15572 1576 15590 1608
rect 15622 1576 15640 1608
rect 15572 1540 15640 1576
rect 14170 1420 14212 1430
rect 14170 560 14171 1420
rect 14211 560 14212 1420
rect 14170 550 14212 560
rect 14051 474 14083 490
rect 14299 522 14331 1458
rect 15572 1508 15590 1540
rect 15622 1508 15640 1540
rect 15572 1472 15640 1508
rect 15572 1440 15590 1472
rect 15622 1440 15640 1472
rect 14431 1420 14555 1430
rect 14431 560 14432 1420
rect 14554 560 14555 1420
rect 14431 550 14555 560
rect 15572 1404 15640 1440
rect 15572 1372 15590 1404
rect 15622 1372 15640 1404
rect 15572 1336 15640 1372
rect 15572 1304 15590 1336
rect 15622 1304 15640 1336
rect 15572 1268 15640 1304
rect 15572 1236 15590 1268
rect 15622 1236 15640 1268
rect 15572 1200 15640 1236
rect 15572 1168 15590 1200
rect 15622 1168 15640 1200
rect 15572 1132 15640 1168
rect 15572 1100 15590 1132
rect 15622 1100 15640 1132
rect 15572 1064 15640 1100
rect 15572 1032 15590 1064
rect 15622 1032 15640 1064
rect 15572 996 15640 1032
rect 15572 964 15590 996
rect 15622 964 15640 996
rect 15572 928 15640 964
rect 15572 896 15590 928
rect 15622 896 15640 928
rect 15572 860 15640 896
rect 15572 828 15590 860
rect 15622 828 15640 860
rect 15572 792 15640 828
rect 15572 760 15590 792
rect 15622 760 15640 792
rect 15572 724 15640 760
rect 15572 692 15590 724
rect 15622 692 15640 724
rect 15572 656 15640 692
rect 15572 624 15590 656
rect 15622 624 15640 656
rect 15572 588 15640 624
rect 15572 556 15590 588
rect 15622 556 15640 588
rect 14299 474 14331 490
rect 15572 520 15640 556
rect 15572 488 15590 520
rect 15622 488 15640 520
rect 15572 428 15640 488
rect 360 414 15640 428
rect 360 410 1487 414
rect 1527 410 2091 414
rect 2131 410 2695 414
rect 2735 410 3299 414
rect 3339 410 3903 414
rect 3943 410 4507 414
rect 4547 410 5111 414
rect 5151 410 5715 414
rect 5755 410 6319 414
rect 6359 410 6923 414
rect 6963 410 7527 414
rect 7567 410 8131 414
rect 8171 410 8735 414
rect 8775 410 9339 414
rect 9379 410 9943 414
rect 9983 410 10547 414
rect 10587 410 11151 414
rect 11191 410 11755 414
rect 11795 410 12359 414
rect 12399 410 12963 414
rect 13003 410 13567 414
rect 13607 410 14171 414
rect 14211 410 15640 414
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1487 410
rect 1527 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2091 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2695 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3299 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3903 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4547 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5151 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5755 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6359 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6923 410
rect 6963 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7527 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8131 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8735 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9983 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10587 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11191 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11755 410
rect 11795 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12359 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12963 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13567 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14171 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 374 1487 378
rect 1527 374 2091 378
rect 2131 374 2695 378
rect 2735 374 3299 378
rect 3339 374 3903 378
rect 3943 374 4507 378
rect 4547 374 5111 378
rect 5151 374 5715 378
rect 5755 374 6319 378
rect 6359 374 6923 378
rect 6963 374 7527 378
rect 7567 374 8131 378
rect 8171 374 8735 378
rect 8775 374 9339 378
rect 9379 374 9943 378
rect 9983 374 10547 378
rect 10587 374 11151 378
rect 11191 374 11755 378
rect 11795 374 12359 378
rect 12399 374 12963 378
rect 13003 374 13567 378
rect 13607 374 14171 378
rect 14211 374 15640 378
rect 360 360 15640 374
rect 15932 4498 16000 4534
rect 15932 4466 15950 4498
rect 15982 4466 16000 4498
rect 15932 4430 16000 4466
rect 15932 4398 15950 4430
rect 15982 4398 16000 4430
rect 15932 4362 16000 4398
rect 15932 4330 15950 4362
rect 15982 4330 16000 4362
rect 15932 4294 16000 4330
rect 15932 4262 15950 4294
rect 15982 4262 16000 4294
rect 15932 4226 16000 4262
rect 15932 4194 15950 4226
rect 15982 4194 16000 4226
rect 15932 4158 16000 4194
rect 15932 4126 15950 4158
rect 15982 4126 16000 4158
rect 15932 4090 16000 4126
rect 15932 4058 15950 4090
rect 15982 4058 16000 4090
rect 15932 4022 16000 4058
rect 15932 3990 15950 4022
rect 15982 3990 16000 4022
rect 15932 3954 16000 3990
rect 15932 3922 15950 3954
rect 15982 3922 16000 3954
rect 15932 3886 16000 3922
rect 15932 3854 15950 3886
rect 15982 3854 16000 3886
rect 15932 3818 16000 3854
rect 15932 3786 15950 3818
rect 15982 3786 16000 3818
rect 15932 3750 16000 3786
rect 15932 3718 15950 3750
rect 15982 3718 16000 3750
rect 15932 3682 16000 3718
rect 15932 3650 15950 3682
rect 15982 3650 16000 3682
rect 15932 3614 16000 3650
rect 15932 3582 15950 3614
rect 15982 3582 16000 3614
rect 15932 3546 16000 3582
rect 15932 3514 15950 3546
rect 15982 3514 16000 3546
rect 15932 3478 16000 3514
rect 15932 3446 15950 3478
rect 15982 3446 16000 3478
rect 15932 3410 16000 3446
rect 15932 3378 15950 3410
rect 15982 3378 16000 3410
rect 15932 3342 16000 3378
rect 15932 3310 15950 3342
rect 15982 3310 16000 3342
rect 15932 3274 16000 3310
rect 15932 3242 15950 3274
rect 15982 3242 16000 3274
rect 15932 3206 16000 3242
rect 15932 3174 15950 3206
rect 15982 3174 16000 3206
rect 15932 3138 16000 3174
rect 15932 3106 15950 3138
rect 15982 3106 16000 3138
rect 15932 3070 16000 3106
rect 15932 3038 15950 3070
rect 15982 3038 16000 3070
rect 15932 3002 16000 3038
rect 15932 2970 15950 3002
rect 15982 2970 16000 3002
rect 15932 2934 16000 2970
rect 15932 2902 15950 2934
rect 15982 2902 16000 2934
rect 15932 2866 16000 2902
rect 15932 2834 15950 2866
rect 15982 2834 16000 2866
rect 15932 2798 16000 2834
rect 15932 2766 15950 2798
rect 15982 2766 16000 2798
rect 15932 2730 16000 2766
rect 15932 2698 15950 2730
rect 15982 2698 16000 2730
rect 15932 2662 16000 2698
rect 15932 2630 15950 2662
rect 15982 2630 16000 2662
rect 15932 2594 16000 2630
rect 15932 2562 15950 2594
rect 15982 2562 16000 2594
rect 15932 2526 16000 2562
rect 15932 2494 15950 2526
rect 15982 2494 16000 2526
rect 15932 2458 16000 2494
rect 15932 2426 15950 2458
rect 15982 2426 16000 2458
rect 15932 2390 16000 2426
rect 15932 2358 15950 2390
rect 15982 2358 16000 2390
rect 15932 2322 16000 2358
rect 15932 2290 15950 2322
rect 15982 2290 16000 2322
rect 15932 2254 16000 2290
rect 15932 2222 15950 2254
rect 15982 2222 16000 2254
rect 15932 2186 16000 2222
rect 15932 2154 15950 2186
rect 15982 2154 16000 2186
rect 15932 2118 16000 2154
rect 15932 2086 15950 2118
rect 15982 2086 16000 2118
rect 15932 2050 16000 2086
rect 15932 2018 15950 2050
rect 15982 2018 16000 2050
rect 15932 1982 16000 2018
rect 15932 1950 15950 1982
rect 15982 1950 16000 1982
rect 15932 1914 16000 1950
rect 15932 1882 15950 1914
rect 15982 1882 16000 1914
rect 15932 1846 16000 1882
rect 15932 1814 15950 1846
rect 15982 1814 16000 1846
rect 15932 1778 16000 1814
rect 15932 1746 15950 1778
rect 15982 1746 16000 1778
rect 15932 1710 16000 1746
rect 15932 1678 15950 1710
rect 15982 1678 16000 1710
rect 15932 1642 16000 1678
rect 15932 1610 15950 1642
rect 15982 1610 16000 1642
rect 15932 1574 16000 1610
rect 15932 1542 15950 1574
rect 15982 1542 16000 1574
rect 15932 1506 16000 1542
rect 15932 1474 15950 1506
rect 15982 1474 16000 1506
rect 15932 1438 16000 1474
rect 15932 1406 15950 1438
rect 15982 1406 16000 1438
rect 15932 1370 16000 1406
rect 15932 1338 15950 1370
rect 15982 1338 16000 1370
rect 15932 1302 16000 1338
rect 15932 1270 15950 1302
rect 15982 1270 16000 1302
rect 15932 1234 16000 1270
rect 15932 1202 15950 1234
rect 15982 1202 16000 1234
rect 15932 1166 16000 1202
rect 15932 1134 15950 1166
rect 15982 1134 16000 1166
rect 15932 1098 16000 1134
rect 15932 1066 15950 1098
rect 15982 1066 16000 1098
rect 15932 1030 16000 1066
rect 15932 998 15950 1030
rect 15982 998 16000 1030
rect 15932 962 16000 998
rect 15932 930 15950 962
rect 15982 930 16000 962
rect 15932 894 16000 930
rect 15932 862 15950 894
rect 15982 862 16000 894
rect 15932 826 16000 862
rect 15932 794 15950 826
rect 15982 794 16000 826
rect 15932 758 16000 794
rect 15932 726 15950 758
rect 15982 726 16000 758
rect 15932 690 16000 726
rect 15932 658 15950 690
rect 15982 658 16000 690
rect 15932 622 16000 658
rect 15932 590 15950 622
rect 15982 590 16000 622
rect 15932 554 16000 590
rect 15932 522 15950 554
rect 15982 522 16000 554
rect 15932 486 16000 522
rect 15932 454 15950 486
rect 15982 454 16000 486
rect 15932 418 16000 454
rect 15932 386 15950 418
rect 15982 386 16000 418
rect 0 318 18 350
rect 50 318 68 350
rect 0 282 68 318
rect 0 250 18 282
rect 50 250 68 282
rect 0 214 68 250
rect 0 182 18 214
rect 50 182 68 214
rect 0 146 68 182
rect 0 114 18 146
rect 50 114 68 146
rect 0 68 68 114
rect 15932 350 16000 386
rect 15932 318 15950 350
rect 15982 318 16000 350
rect 15932 282 16000 318
rect 15932 250 15950 282
rect 15982 250 16000 282
rect 15932 214 16000 250
rect 15932 182 15950 214
rect 15982 182 16000 214
rect 15932 146 16000 182
rect 15932 114 15950 146
rect 15982 114 16000 146
rect 15932 68 16000 114
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 1487 4506 1527 4510
rect 2091 4506 2131 4510
rect 2695 4506 2735 4510
rect 3299 4506 3339 4510
rect 3903 4506 3943 4510
rect 4507 4506 4547 4510
rect 5111 4506 5151 4510
rect 5715 4506 5755 4510
rect 6319 4506 6359 4510
rect 6923 4506 6963 4510
rect 7527 4506 7567 4510
rect 8131 4506 8171 4510
rect 8735 4506 8775 4510
rect 9339 4506 9379 4510
rect 9943 4506 9983 4510
rect 10547 4506 10587 4510
rect 11151 4506 11191 4510
rect 11755 4506 11795 4510
rect 12359 4506 12399 4510
rect 12963 4506 13003 4510
rect 13567 4506 13607 4510
rect 14171 4506 14211 4510
rect 1487 4474 1490 4506
rect 1490 4474 1522 4506
rect 1522 4474 1527 4506
rect 2091 4474 2102 4506
rect 2102 4474 2131 4506
rect 2695 4474 2714 4506
rect 2714 4474 2735 4506
rect 3299 4474 3326 4506
rect 3326 4474 3339 4506
rect 3903 4474 3938 4506
rect 3938 4474 3943 4506
rect 4507 4474 4514 4506
rect 4514 4474 4547 4506
rect 5111 4474 5126 4506
rect 5126 4474 5151 4506
rect 5715 4474 5738 4506
rect 5738 4474 5755 4506
rect 6319 4474 6350 4506
rect 6350 4474 6359 4506
rect 6923 4474 6930 4506
rect 6930 4474 6962 4506
rect 6962 4474 6963 4506
rect 7527 4474 7542 4506
rect 7542 4474 7567 4506
rect 8131 4474 8154 4506
rect 8154 4474 8171 4506
rect 8735 4474 8766 4506
rect 8766 4474 8775 4506
rect 9339 4474 9342 4506
rect 9342 4474 9378 4506
rect 9378 4474 9379 4506
rect 9943 4474 9954 4506
rect 9954 4474 9983 4506
rect 10547 4474 10566 4506
rect 10566 4474 10587 4506
rect 11151 4474 11178 4506
rect 11178 4474 11191 4506
rect 11755 4474 11758 4506
rect 11758 4474 11790 4506
rect 11790 4474 11795 4506
rect 12359 4474 12370 4506
rect 12370 4474 12399 4506
rect 12963 4474 12982 4506
rect 12982 4474 13003 4506
rect 13567 4474 13594 4506
rect 13594 4474 13607 4506
rect 14171 4474 14206 4506
rect 14206 4474 14211 4506
rect 1487 4470 1527 4474
rect 2091 4470 2131 4474
rect 2695 4470 2735 4474
rect 3299 4470 3339 4474
rect 3903 4470 3943 4474
rect 4507 4470 4547 4474
rect 5111 4470 5151 4474
rect 5715 4470 5755 4474
rect 6319 4470 6359 4474
rect 6923 4470 6963 4474
rect 7527 4470 7567 4474
rect 8131 4470 8171 4474
rect 8735 4470 8775 4474
rect 9339 4470 9379 4474
rect 9943 4470 9983 4474
rect 10547 4470 10587 4474
rect 11151 4470 11191 4474
rect 11755 4470 11795 4474
rect 12359 4470 12399 4474
rect 12963 4470 13003 4474
rect 13567 4470 13607 4474
rect 14171 4470 14211 4474
rect 933 4246 973 4368
rect 1487 4318 1527 4324
rect 1487 4286 1491 4318
rect 1491 4286 1523 4318
rect 1523 4286 1527 4318
rect 1487 4250 1527 4286
rect 1487 4218 1491 4250
rect 1491 4218 1523 4250
rect 1523 4218 1527 4250
rect 1487 4182 1527 4218
rect 1487 4150 1491 4182
rect 1491 4150 1523 4182
rect 1523 4150 1527 4182
rect 1487 4114 1527 4150
rect 1487 4082 1491 4114
rect 1491 4082 1523 4114
rect 1523 4082 1527 4114
rect 1487 4046 1527 4082
rect 1487 4014 1491 4046
rect 1491 4014 1523 4046
rect 1523 4014 1527 4046
rect 1487 3978 1527 4014
rect 1487 3946 1491 3978
rect 1491 3946 1523 3978
rect 1523 3946 1527 3978
rect 1487 3910 1527 3946
rect 1487 3878 1491 3910
rect 1491 3878 1523 3910
rect 1523 3878 1527 3910
rect 1487 3842 1527 3878
rect 1487 3810 1491 3842
rect 1491 3810 1523 3842
rect 1523 3810 1527 3842
rect 1487 3774 1527 3810
rect 1487 3742 1491 3774
rect 1491 3742 1523 3774
rect 1523 3742 1527 3774
rect 1487 3706 1527 3742
rect 1487 3674 1491 3706
rect 1491 3674 1523 3706
rect 1523 3674 1527 3706
rect 1487 3638 1527 3674
rect 1487 3606 1491 3638
rect 1491 3606 1523 3638
rect 1523 3606 1527 3638
rect 1487 3570 1527 3606
rect 1487 3538 1491 3570
rect 1491 3538 1523 3570
rect 1523 3538 1527 3570
rect 1487 3502 1527 3538
rect 1487 3470 1491 3502
rect 1491 3470 1523 3502
rect 1523 3470 1527 3502
rect 1487 3464 1527 3470
rect 1748 4318 1870 4324
rect 1748 4286 1793 4318
rect 1793 4286 1825 4318
rect 1825 4286 1870 4318
rect 1748 4250 1870 4286
rect 1748 4218 1793 4250
rect 1793 4218 1825 4250
rect 1825 4218 1870 4250
rect 1748 4182 1870 4218
rect 1748 4150 1793 4182
rect 1793 4150 1825 4182
rect 1825 4150 1870 4182
rect 1748 4114 1870 4150
rect 1748 4082 1793 4114
rect 1793 4082 1825 4114
rect 1825 4082 1870 4114
rect 1748 4046 1870 4082
rect 1748 4014 1793 4046
rect 1793 4014 1825 4046
rect 1825 4014 1870 4046
rect 1748 3978 1870 4014
rect 1748 3946 1793 3978
rect 1793 3946 1825 3978
rect 1825 3946 1870 3978
rect 1748 3910 1870 3946
rect 1748 3878 1793 3910
rect 1793 3878 1825 3910
rect 1825 3878 1870 3910
rect 1748 3842 1870 3878
rect 1748 3810 1793 3842
rect 1793 3810 1825 3842
rect 1825 3810 1870 3842
rect 1748 3774 1870 3810
rect 1748 3742 1793 3774
rect 1793 3742 1825 3774
rect 1825 3742 1870 3774
rect 1748 3706 1870 3742
rect 1748 3674 1793 3706
rect 1793 3674 1825 3706
rect 1825 3674 1870 3706
rect 1748 3638 1870 3674
rect 1748 3606 1793 3638
rect 1793 3606 1825 3638
rect 1825 3606 1870 3638
rect 1748 3570 1870 3606
rect 1748 3538 1793 3570
rect 1793 3538 1825 3570
rect 1825 3538 1870 3570
rect 1748 3502 1870 3538
rect 1748 3470 1793 3502
rect 1793 3470 1825 3502
rect 1825 3470 1870 3502
rect 1748 3464 1870 3470
rect 1487 3350 1527 3356
rect 1487 3318 1491 3350
rect 1491 3318 1523 3350
rect 1523 3318 1527 3350
rect 1487 3282 1527 3318
rect 1487 3250 1491 3282
rect 1491 3250 1523 3282
rect 1523 3250 1527 3282
rect 1487 3214 1527 3250
rect 1487 3182 1491 3214
rect 1491 3182 1523 3214
rect 1523 3182 1527 3214
rect 1487 3146 1527 3182
rect 1487 3114 1491 3146
rect 1491 3114 1523 3146
rect 1523 3114 1527 3146
rect 1487 3078 1527 3114
rect 1487 3046 1491 3078
rect 1491 3046 1523 3078
rect 1523 3046 1527 3078
rect 1487 3010 1527 3046
rect 1487 2978 1491 3010
rect 1491 2978 1523 3010
rect 1523 2978 1527 3010
rect 1487 2942 1527 2978
rect 1487 2910 1491 2942
rect 1491 2910 1523 2942
rect 1523 2910 1527 2942
rect 1487 2874 1527 2910
rect 1487 2842 1491 2874
rect 1491 2842 1523 2874
rect 1523 2842 1527 2874
rect 1487 2806 1527 2842
rect 1487 2774 1491 2806
rect 1491 2774 1523 2806
rect 1523 2774 1527 2806
rect 1487 2738 1527 2774
rect 1487 2706 1491 2738
rect 1491 2706 1523 2738
rect 1523 2706 1527 2738
rect 1487 2670 1527 2706
rect 1487 2638 1491 2670
rect 1491 2638 1523 2670
rect 1523 2638 1527 2670
rect 1487 2602 1527 2638
rect 1487 2570 1491 2602
rect 1491 2570 1523 2602
rect 1523 2570 1527 2602
rect 1487 2534 1527 2570
rect 1487 2502 1491 2534
rect 1491 2502 1523 2534
rect 1523 2502 1527 2534
rect 1487 2496 1527 2502
rect 2091 4318 2131 4324
rect 2091 4286 2095 4318
rect 2095 4286 2127 4318
rect 2127 4286 2131 4318
rect 2091 4250 2131 4286
rect 2091 4218 2095 4250
rect 2095 4218 2127 4250
rect 2127 4218 2131 4250
rect 2091 4182 2131 4218
rect 2091 4150 2095 4182
rect 2095 4150 2127 4182
rect 2127 4150 2131 4182
rect 2091 4114 2131 4150
rect 2091 4082 2095 4114
rect 2095 4082 2127 4114
rect 2127 4082 2131 4114
rect 2091 4046 2131 4082
rect 2091 4014 2095 4046
rect 2095 4014 2127 4046
rect 2127 4014 2131 4046
rect 2091 3978 2131 4014
rect 2091 3946 2095 3978
rect 2095 3946 2127 3978
rect 2127 3946 2131 3978
rect 2091 3910 2131 3946
rect 2091 3878 2095 3910
rect 2095 3878 2127 3910
rect 2127 3878 2131 3910
rect 2091 3842 2131 3878
rect 2091 3810 2095 3842
rect 2095 3810 2127 3842
rect 2127 3810 2131 3842
rect 2091 3774 2131 3810
rect 2091 3742 2095 3774
rect 2095 3742 2127 3774
rect 2127 3742 2131 3774
rect 2091 3706 2131 3742
rect 2091 3674 2095 3706
rect 2095 3674 2127 3706
rect 2127 3674 2131 3706
rect 2091 3638 2131 3674
rect 2091 3606 2095 3638
rect 2095 3606 2127 3638
rect 2127 3606 2131 3638
rect 2091 3570 2131 3606
rect 2091 3538 2095 3570
rect 2095 3538 2127 3570
rect 2127 3538 2131 3570
rect 2091 3502 2131 3538
rect 2091 3470 2095 3502
rect 2095 3470 2127 3502
rect 2127 3470 2131 3502
rect 2091 3464 2131 3470
rect 1748 3350 1870 3356
rect 1748 3318 1793 3350
rect 1793 3318 1825 3350
rect 1825 3318 1870 3350
rect 1748 3282 1870 3318
rect 1748 3250 1793 3282
rect 1793 3250 1825 3282
rect 1825 3250 1870 3282
rect 1748 3214 1870 3250
rect 1748 3182 1793 3214
rect 1793 3182 1825 3214
rect 1825 3182 1870 3214
rect 1748 3146 1870 3182
rect 1748 3114 1793 3146
rect 1793 3114 1825 3146
rect 1825 3114 1870 3146
rect 1748 3078 1870 3114
rect 1748 3046 1793 3078
rect 1793 3046 1825 3078
rect 1825 3046 1870 3078
rect 1748 3010 1870 3046
rect 1748 2978 1793 3010
rect 1793 2978 1825 3010
rect 1825 2978 1870 3010
rect 1748 2942 1870 2978
rect 1748 2910 1793 2942
rect 1793 2910 1825 2942
rect 1825 2910 1870 2942
rect 1748 2874 1870 2910
rect 1748 2842 1793 2874
rect 1793 2842 1825 2874
rect 1825 2842 1870 2874
rect 1748 2806 1870 2842
rect 1748 2774 1793 2806
rect 1793 2774 1825 2806
rect 1825 2774 1870 2806
rect 1748 2738 1870 2774
rect 1748 2706 1793 2738
rect 1793 2706 1825 2738
rect 1825 2706 1870 2738
rect 1748 2670 1870 2706
rect 1748 2638 1793 2670
rect 1793 2638 1825 2670
rect 1825 2638 1870 2670
rect 1748 2602 1870 2638
rect 1748 2570 1793 2602
rect 1793 2570 1825 2602
rect 1825 2570 1870 2602
rect 1748 2534 1870 2570
rect 1748 2502 1793 2534
rect 1793 2502 1825 2534
rect 1825 2502 1870 2534
rect 1748 2496 1870 2502
rect 1487 2382 1527 2388
rect 1487 2350 1491 2382
rect 1491 2350 1523 2382
rect 1523 2350 1527 2382
rect 1487 2314 1527 2350
rect 1487 2282 1491 2314
rect 1491 2282 1523 2314
rect 1523 2282 1527 2314
rect 1487 2246 1527 2282
rect 1487 2214 1491 2246
rect 1491 2214 1523 2246
rect 1523 2214 1527 2246
rect 1487 2178 1527 2214
rect 1487 2146 1491 2178
rect 1491 2146 1523 2178
rect 1523 2146 1527 2178
rect 1487 2110 1527 2146
rect 1487 2078 1491 2110
rect 1491 2078 1523 2110
rect 1523 2078 1527 2110
rect 1487 2042 1527 2078
rect 1487 2010 1491 2042
rect 1491 2010 1523 2042
rect 1523 2010 1527 2042
rect 1487 1974 1527 2010
rect 1487 1942 1491 1974
rect 1491 1942 1523 1974
rect 1523 1942 1527 1974
rect 1487 1906 1527 1942
rect 1487 1874 1491 1906
rect 1491 1874 1523 1906
rect 1523 1874 1527 1906
rect 1487 1838 1527 1874
rect 1487 1806 1491 1838
rect 1491 1806 1523 1838
rect 1523 1806 1527 1838
rect 1487 1770 1527 1806
rect 1487 1738 1491 1770
rect 1491 1738 1523 1770
rect 1523 1738 1527 1770
rect 1487 1702 1527 1738
rect 1487 1670 1491 1702
rect 1491 1670 1523 1702
rect 1523 1670 1527 1702
rect 1487 1634 1527 1670
rect 1487 1602 1491 1634
rect 1491 1602 1523 1634
rect 1523 1602 1527 1634
rect 1487 1566 1527 1602
rect 1487 1534 1491 1566
rect 1491 1534 1523 1566
rect 1523 1534 1527 1566
rect 1487 1528 1527 1534
rect 2352 4318 2474 4324
rect 2352 4286 2397 4318
rect 2397 4286 2429 4318
rect 2429 4286 2474 4318
rect 2352 4250 2474 4286
rect 2352 4218 2397 4250
rect 2397 4218 2429 4250
rect 2429 4218 2474 4250
rect 2352 4182 2474 4218
rect 2352 4150 2397 4182
rect 2397 4150 2429 4182
rect 2429 4150 2474 4182
rect 2352 4114 2474 4150
rect 2352 4082 2397 4114
rect 2397 4082 2429 4114
rect 2429 4082 2474 4114
rect 2352 4046 2474 4082
rect 2352 4014 2397 4046
rect 2397 4014 2429 4046
rect 2429 4014 2474 4046
rect 2352 3978 2474 4014
rect 2352 3946 2397 3978
rect 2397 3946 2429 3978
rect 2429 3946 2474 3978
rect 2352 3910 2474 3946
rect 2352 3878 2397 3910
rect 2397 3878 2429 3910
rect 2429 3878 2474 3910
rect 2352 3842 2474 3878
rect 2352 3810 2397 3842
rect 2397 3810 2429 3842
rect 2429 3810 2474 3842
rect 2352 3774 2474 3810
rect 2352 3742 2397 3774
rect 2397 3742 2429 3774
rect 2429 3742 2474 3774
rect 2352 3706 2474 3742
rect 2352 3674 2397 3706
rect 2397 3674 2429 3706
rect 2429 3674 2474 3706
rect 2352 3638 2474 3674
rect 2352 3606 2397 3638
rect 2397 3606 2429 3638
rect 2429 3606 2474 3638
rect 2352 3570 2474 3606
rect 2352 3538 2397 3570
rect 2397 3538 2429 3570
rect 2429 3538 2474 3570
rect 2352 3502 2474 3538
rect 2352 3470 2397 3502
rect 2397 3470 2429 3502
rect 2429 3470 2474 3502
rect 2352 3464 2474 3470
rect 2091 3350 2131 3356
rect 2091 3318 2095 3350
rect 2095 3318 2127 3350
rect 2127 3318 2131 3350
rect 2091 3282 2131 3318
rect 2091 3250 2095 3282
rect 2095 3250 2127 3282
rect 2127 3250 2131 3282
rect 2091 3214 2131 3250
rect 2091 3182 2095 3214
rect 2095 3182 2127 3214
rect 2127 3182 2131 3214
rect 2091 3146 2131 3182
rect 2091 3114 2095 3146
rect 2095 3114 2127 3146
rect 2127 3114 2131 3146
rect 2091 3078 2131 3114
rect 2091 3046 2095 3078
rect 2095 3046 2127 3078
rect 2127 3046 2131 3078
rect 2091 3010 2131 3046
rect 2091 2978 2095 3010
rect 2095 2978 2127 3010
rect 2127 2978 2131 3010
rect 2091 2942 2131 2978
rect 2091 2910 2095 2942
rect 2095 2910 2127 2942
rect 2127 2910 2131 2942
rect 2091 2874 2131 2910
rect 2091 2842 2095 2874
rect 2095 2842 2127 2874
rect 2127 2842 2131 2874
rect 2091 2806 2131 2842
rect 2091 2774 2095 2806
rect 2095 2774 2127 2806
rect 2127 2774 2131 2806
rect 2091 2738 2131 2774
rect 2091 2706 2095 2738
rect 2095 2706 2127 2738
rect 2127 2706 2131 2738
rect 2091 2670 2131 2706
rect 2091 2638 2095 2670
rect 2095 2638 2127 2670
rect 2127 2638 2131 2670
rect 2091 2602 2131 2638
rect 2091 2570 2095 2602
rect 2095 2570 2127 2602
rect 2127 2570 2131 2602
rect 2091 2534 2131 2570
rect 2091 2502 2095 2534
rect 2095 2502 2127 2534
rect 2127 2502 2131 2534
rect 2091 2496 2131 2502
rect 1748 2382 1870 2388
rect 1748 2350 1793 2382
rect 1793 2350 1825 2382
rect 1825 2350 1870 2382
rect 1748 2314 1870 2350
rect 1748 2282 1793 2314
rect 1793 2282 1825 2314
rect 1825 2282 1870 2314
rect 1748 2246 1870 2282
rect 1748 2214 1793 2246
rect 1793 2214 1825 2246
rect 1825 2214 1870 2246
rect 1748 2178 1870 2214
rect 1748 2146 1793 2178
rect 1793 2146 1825 2178
rect 1825 2146 1870 2178
rect 1748 2110 1870 2146
rect 1748 2078 1793 2110
rect 1793 2078 1825 2110
rect 1825 2078 1870 2110
rect 1748 2042 1870 2078
rect 1748 2010 1793 2042
rect 1793 2010 1825 2042
rect 1825 2010 1870 2042
rect 1748 1974 1870 2010
rect 1748 1942 1793 1974
rect 1793 1942 1825 1974
rect 1825 1942 1870 1974
rect 1748 1906 1870 1942
rect 1748 1874 1793 1906
rect 1793 1874 1825 1906
rect 1825 1874 1870 1906
rect 1748 1838 1870 1874
rect 1748 1806 1793 1838
rect 1793 1806 1825 1838
rect 1825 1806 1870 1838
rect 1748 1770 1870 1806
rect 1748 1738 1793 1770
rect 1793 1738 1825 1770
rect 1825 1738 1870 1770
rect 1748 1702 1870 1738
rect 1748 1670 1793 1702
rect 1793 1670 1825 1702
rect 1825 1670 1870 1702
rect 1748 1634 1870 1670
rect 1748 1602 1793 1634
rect 1793 1602 1825 1634
rect 1825 1602 1870 1634
rect 1748 1566 1870 1602
rect 1748 1534 1793 1566
rect 1793 1534 1825 1566
rect 1825 1534 1870 1566
rect 1748 1528 1870 1534
rect 1487 1414 1527 1420
rect 1487 1382 1491 1414
rect 1491 1382 1523 1414
rect 1523 1382 1527 1414
rect 1487 1346 1527 1382
rect 1487 1314 1491 1346
rect 1491 1314 1523 1346
rect 1523 1314 1527 1346
rect 1487 1278 1527 1314
rect 1487 1246 1491 1278
rect 1491 1246 1523 1278
rect 1523 1246 1527 1278
rect 1487 1210 1527 1246
rect 1487 1178 1491 1210
rect 1491 1178 1523 1210
rect 1523 1178 1527 1210
rect 1487 1142 1527 1178
rect 1487 1110 1491 1142
rect 1491 1110 1523 1142
rect 1523 1110 1527 1142
rect 1487 1074 1527 1110
rect 1487 1042 1491 1074
rect 1491 1042 1523 1074
rect 1523 1042 1527 1074
rect 1487 1006 1527 1042
rect 1487 974 1491 1006
rect 1491 974 1523 1006
rect 1523 974 1527 1006
rect 1487 938 1527 974
rect 1487 906 1491 938
rect 1491 906 1523 938
rect 1523 906 1527 938
rect 1487 870 1527 906
rect 1487 838 1491 870
rect 1491 838 1523 870
rect 1523 838 1527 870
rect 1487 802 1527 838
rect 1487 770 1491 802
rect 1491 770 1523 802
rect 1523 770 1527 802
rect 1487 734 1527 770
rect 1487 702 1491 734
rect 1491 702 1523 734
rect 1523 702 1527 734
rect 1487 666 1527 702
rect 1487 634 1491 666
rect 1491 634 1523 666
rect 1523 634 1527 666
rect 1487 598 1527 634
rect 1487 566 1491 598
rect 1491 566 1523 598
rect 1523 566 1527 598
rect 1487 560 1527 566
rect 2695 4318 2735 4324
rect 2695 4286 2699 4318
rect 2699 4286 2731 4318
rect 2731 4286 2735 4318
rect 2695 4250 2735 4286
rect 2695 4218 2699 4250
rect 2699 4218 2731 4250
rect 2731 4218 2735 4250
rect 2695 4182 2735 4218
rect 2695 4150 2699 4182
rect 2699 4150 2731 4182
rect 2731 4150 2735 4182
rect 2695 4114 2735 4150
rect 2695 4082 2699 4114
rect 2699 4082 2731 4114
rect 2731 4082 2735 4114
rect 2695 4046 2735 4082
rect 2695 4014 2699 4046
rect 2699 4014 2731 4046
rect 2731 4014 2735 4046
rect 2695 3978 2735 4014
rect 2695 3946 2699 3978
rect 2699 3946 2731 3978
rect 2731 3946 2735 3978
rect 2695 3910 2735 3946
rect 2695 3878 2699 3910
rect 2699 3878 2731 3910
rect 2731 3878 2735 3910
rect 2695 3842 2735 3878
rect 2695 3810 2699 3842
rect 2699 3810 2731 3842
rect 2731 3810 2735 3842
rect 2695 3774 2735 3810
rect 2695 3742 2699 3774
rect 2699 3742 2731 3774
rect 2731 3742 2735 3774
rect 2695 3706 2735 3742
rect 2695 3674 2699 3706
rect 2699 3674 2731 3706
rect 2731 3674 2735 3706
rect 2695 3638 2735 3674
rect 2695 3606 2699 3638
rect 2699 3606 2731 3638
rect 2731 3606 2735 3638
rect 2695 3570 2735 3606
rect 2695 3538 2699 3570
rect 2699 3538 2731 3570
rect 2731 3538 2735 3570
rect 2695 3502 2735 3538
rect 2695 3470 2699 3502
rect 2699 3470 2731 3502
rect 2731 3470 2735 3502
rect 2695 3464 2735 3470
rect 2352 3350 2474 3356
rect 2352 3318 2397 3350
rect 2397 3318 2429 3350
rect 2429 3318 2474 3350
rect 2352 3282 2474 3318
rect 2352 3250 2397 3282
rect 2397 3250 2429 3282
rect 2429 3250 2474 3282
rect 2352 3214 2474 3250
rect 2352 3182 2397 3214
rect 2397 3182 2429 3214
rect 2429 3182 2474 3214
rect 2352 3146 2474 3182
rect 2352 3114 2397 3146
rect 2397 3114 2429 3146
rect 2429 3114 2474 3146
rect 2352 3078 2474 3114
rect 2352 3046 2397 3078
rect 2397 3046 2429 3078
rect 2429 3046 2474 3078
rect 2352 3010 2474 3046
rect 2352 2978 2397 3010
rect 2397 2978 2429 3010
rect 2429 2978 2474 3010
rect 2352 2942 2474 2978
rect 2352 2910 2397 2942
rect 2397 2910 2429 2942
rect 2429 2910 2474 2942
rect 2352 2874 2474 2910
rect 2352 2842 2397 2874
rect 2397 2842 2429 2874
rect 2429 2842 2474 2874
rect 2352 2806 2474 2842
rect 2352 2774 2397 2806
rect 2397 2774 2429 2806
rect 2429 2774 2474 2806
rect 2352 2738 2474 2774
rect 2352 2706 2397 2738
rect 2397 2706 2429 2738
rect 2429 2706 2474 2738
rect 2352 2670 2474 2706
rect 2352 2638 2397 2670
rect 2397 2638 2429 2670
rect 2429 2638 2474 2670
rect 2352 2602 2474 2638
rect 2352 2570 2397 2602
rect 2397 2570 2429 2602
rect 2429 2570 2474 2602
rect 2352 2534 2474 2570
rect 2352 2502 2397 2534
rect 2397 2502 2429 2534
rect 2429 2502 2474 2534
rect 2352 2496 2474 2502
rect 2091 2382 2131 2388
rect 2091 2350 2095 2382
rect 2095 2350 2127 2382
rect 2127 2350 2131 2382
rect 2091 2314 2131 2350
rect 2091 2282 2095 2314
rect 2095 2282 2127 2314
rect 2127 2282 2131 2314
rect 2091 2246 2131 2282
rect 2091 2214 2095 2246
rect 2095 2214 2127 2246
rect 2127 2214 2131 2246
rect 2091 2178 2131 2214
rect 2091 2146 2095 2178
rect 2095 2146 2127 2178
rect 2127 2146 2131 2178
rect 2091 2110 2131 2146
rect 2091 2078 2095 2110
rect 2095 2078 2127 2110
rect 2127 2078 2131 2110
rect 2091 2042 2131 2078
rect 2091 2010 2095 2042
rect 2095 2010 2127 2042
rect 2127 2010 2131 2042
rect 2091 1974 2131 2010
rect 2091 1942 2095 1974
rect 2095 1942 2127 1974
rect 2127 1942 2131 1974
rect 2091 1906 2131 1942
rect 2091 1874 2095 1906
rect 2095 1874 2127 1906
rect 2127 1874 2131 1906
rect 2091 1838 2131 1874
rect 2091 1806 2095 1838
rect 2095 1806 2127 1838
rect 2127 1806 2131 1838
rect 2091 1770 2131 1806
rect 2091 1738 2095 1770
rect 2095 1738 2127 1770
rect 2127 1738 2131 1770
rect 2091 1702 2131 1738
rect 2091 1670 2095 1702
rect 2095 1670 2127 1702
rect 2127 1670 2131 1702
rect 2091 1634 2131 1670
rect 2091 1602 2095 1634
rect 2095 1602 2127 1634
rect 2127 1602 2131 1634
rect 2091 1566 2131 1602
rect 2091 1534 2095 1566
rect 2095 1534 2127 1566
rect 2127 1534 2131 1566
rect 2091 1528 2131 1534
rect 1748 1414 1870 1420
rect 1748 1382 1793 1414
rect 1793 1382 1825 1414
rect 1825 1382 1870 1414
rect 1748 1346 1870 1382
rect 1748 1314 1793 1346
rect 1793 1314 1825 1346
rect 1825 1314 1870 1346
rect 1748 1278 1870 1314
rect 1748 1246 1793 1278
rect 1793 1246 1825 1278
rect 1825 1246 1870 1278
rect 1748 1210 1870 1246
rect 1748 1178 1793 1210
rect 1793 1178 1825 1210
rect 1825 1178 1870 1210
rect 1748 1142 1870 1178
rect 1748 1110 1793 1142
rect 1793 1110 1825 1142
rect 1825 1110 1870 1142
rect 1748 1074 1870 1110
rect 1748 1042 1793 1074
rect 1793 1042 1825 1074
rect 1825 1042 1870 1074
rect 1748 1006 1870 1042
rect 1748 974 1793 1006
rect 1793 974 1825 1006
rect 1825 974 1870 1006
rect 1748 938 1870 974
rect 1748 906 1793 938
rect 1793 906 1825 938
rect 1825 906 1870 938
rect 1748 870 1870 906
rect 1748 838 1793 870
rect 1793 838 1825 870
rect 1825 838 1870 870
rect 1748 802 1870 838
rect 1748 770 1793 802
rect 1793 770 1825 802
rect 1825 770 1870 802
rect 1748 734 1870 770
rect 1748 702 1793 734
rect 1793 702 1825 734
rect 1825 702 1870 734
rect 1748 666 1870 702
rect 1748 634 1793 666
rect 1793 634 1825 666
rect 1825 634 1870 666
rect 1748 598 1870 634
rect 1748 566 1793 598
rect 1793 566 1825 598
rect 1825 566 1870 598
rect 1748 560 1870 566
rect 2956 4318 3078 4324
rect 2956 4286 3001 4318
rect 3001 4286 3033 4318
rect 3033 4286 3078 4318
rect 2956 4250 3078 4286
rect 2956 4218 3001 4250
rect 3001 4218 3033 4250
rect 3033 4218 3078 4250
rect 2956 4182 3078 4218
rect 2956 4150 3001 4182
rect 3001 4150 3033 4182
rect 3033 4150 3078 4182
rect 2956 4114 3078 4150
rect 2956 4082 3001 4114
rect 3001 4082 3033 4114
rect 3033 4082 3078 4114
rect 2956 4046 3078 4082
rect 2956 4014 3001 4046
rect 3001 4014 3033 4046
rect 3033 4014 3078 4046
rect 2956 3978 3078 4014
rect 2956 3946 3001 3978
rect 3001 3946 3033 3978
rect 3033 3946 3078 3978
rect 2956 3910 3078 3946
rect 2956 3878 3001 3910
rect 3001 3878 3033 3910
rect 3033 3878 3078 3910
rect 2956 3842 3078 3878
rect 2956 3810 3001 3842
rect 3001 3810 3033 3842
rect 3033 3810 3078 3842
rect 2956 3774 3078 3810
rect 2956 3742 3001 3774
rect 3001 3742 3033 3774
rect 3033 3742 3078 3774
rect 2956 3706 3078 3742
rect 2956 3674 3001 3706
rect 3001 3674 3033 3706
rect 3033 3674 3078 3706
rect 2956 3638 3078 3674
rect 2956 3606 3001 3638
rect 3001 3606 3033 3638
rect 3033 3606 3078 3638
rect 2956 3570 3078 3606
rect 2956 3538 3001 3570
rect 3001 3538 3033 3570
rect 3033 3538 3078 3570
rect 2956 3502 3078 3538
rect 2956 3470 3001 3502
rect 3001 3470 3033 3502
rect 3033 3470 3078 3502
rect 2956 3464 3078 3470
rect 2695 3350 2735 3356
rect 2695 3318 2699 3350
rect 2699 3318 2731 3350
rect 2731 3318 2735 3350
rect 2695 3282 2735 3318
rect 2695 3250 2699 3282
rect 2699 3250 2731 3282
rect 2731 3250 2735 3282
rect 2695 3214 2735 3250
rect 2695 3182 2699 3214
rect 2699 3182 2731 3214
rect 2731 3182 2735 3214
rect 2695 3146 2735 3182
rect 2695 3114 2699 3146
rect 2699 3114 2731 3146
rect 2731 3114 2735 3146
rect 2695 3078 2735 3114
rect 2695 3046 2699 3078
rect 2699 3046 2731 3078
rect 2731 3046 2735 3078
rect 2695 3010 2735 3046
rect 2695 2978 2699 3010
rect 2699 2978 2731 3010
rect 2731 2978 2735 3010
rect 2695 2942 2735 2978
rect 2695 2910 2699 2942
rect 2699 2910 2731 2942
rect 2731 2910 2735 2942
rect 2695 2874 2735 2910
rect 2695 2842 2699 2874
rect 2699 2842 2731 2874
rect 2731 2842 2735 2874
rect 2695 2806 2735 2842
rect 2695 2774 2699 2806
rect 2699 2774 2731 2806
rect 2731 2774 2735 2806
rect 2695 2738 2735 2774
rect 2695 2706 2699 2738
rect 2699 2706 2731 2738
rect 2731 2706 2735 2738
rect 2695 2670 2735 2706
rect 2695 2638 2699 2670
rect 2699 2638 2731 2670
rect 2731 2638 2735 2670
rect 2695 2602 2735 2638
rect 2695 2570 2699 2602
rect 2699 2570 2731 2602
rect 2731 2570 2735 2602
rect 2695 2534 2735 2570
rect 2695 2502 2699 2534
rect 2699 2502 2731 2534
rect 2731 2502 2735 2534
rect 2695 2496 2735 2502
rect 2352 2382 2474 2388
rect 2352 2350 2397 2382
rect 2397 2350 2429 2382
rect 2429 2350 2474 2382
rect 2352 2314 2474 2350
rect 2352 2282 2397 2314
rect 2397 2282 2429 2314
rect 2429 2282 2474 2314
rect 2352 2246 2474 2282
rect 2352 2214 2397 2246
rect 2397 2214 2429 2246
rect 2429 2214 2474 2246
rect 2352 2178 2474 2214
rect 2352 2146 2397 2178
rect 2397 2146 2429 2178
rect 2429 2146 2474 2178
rect 2352 2110 2474 2146
rect 2352 2078 2397 2110
rect 2397 2078 2429 2110
rect 2429 2078 2474 2110
rect 2352 2042 2474 2078
rect 2352 2010 2397 2042
rect 2397 2010 2429 2042
rect 2429 2010 2474 2042
rect 2352 1974 2474 2010
rect 2352 1942 2397 1974
rect 2397 1942 2429 1974
rect 2429 1942 2474 1974
rect 2352 1906 2474 1942
rect 2352 1874 2397 1906
rect 2397 1874 2429 1906
rect 2429 1874 2474 1906
rect 2352 1838 2474 1874
rect 2352 1806 2397 1838
rect 2397 1806 2429 1838
rect 2429 1806 2474 1838
rect 2352 1770 2474 1806
rect 2352 1738 2397 1770
rect 2397 1738 2429 1770
rect 2429 1738 2474 1770
rect 2352 1702 2474 1738
rect 2352 1670 2397 1702
rect 2397 1670 2429 1702
rect 2429 1670 2474 1702
rect 2352 1634 2474 1670
rect 2352 1602 2397 1634
rect 2397 1602 2429 1634
rect 2429 1602 2474 1634
rect 2352 1566 2474 1602
rect 2352 1534 2397 1566
rect 2397 1534 2429 1566
rect 2429 1534 2474 1566
rect 2352 1528 2474 1534
rect 2091 1414 2131 1420
rect 2091 1382 2095 1414
rect 2095 1382 2127 1414
rect 2127 1382 2131 1414
rect 2091 1346 2131 1382
rect 2091 1314 2095 1346
rect 2095 1314 2127 1346
rect 2127 1314 2131 1346
rect 2091 1278 2131 1314
rect 2091 1246 2095 1278
rect 2095 1246 2127 1278
rect 2127 1246 2131 1278
rect 2091 1210 2131 1246
rect 2091 1178 2095 1210
rect 2095 1178 2127 1210
rect 2127 1178 2131 1210
rect 2091 1142 2131 1178
rect 2091 1110 2095 1142
rect 2095 1110 2127 1142
rect 2127 1110 2131 1142
rect 2091 1074 2131 1110
rect 2091 1042 2095 1074
rect 2095 1042 2127 1074
rect 2127 1042 2131 1074
rect 2091 1006 2131 1042
rect 2091 974 2095 1006
rect 2095 974 2127 1006
rect 2127 974 2131 1006
rect 2091 938 2131 974
rect 2091 906 2095 938
rect 2095 906 2127 938
rect 2127 906 2131 938
rect 2091 870 2131 906
rect 2091 838 2095 870
rect 2095 838 2127 870
rect 2127 838 2131 870
rect 2091 802 2131 838
rect 2091 770 2095 802
rect 2095 770 2127 802
rect 2127 770 2131 802
rect 2091 734 2131 770
rect 2091 702 2095 734
rect 2095 702 2127 734
rect 2127 702 2131 734
rect 2091 666 2131 702
rect 2091 634 2095 666
rect 2095 634 2127 666
rect 2127 634 2131 666
rect 2091 598 2131 634
rect 2091 566 2095 598
rect 2095 566 2127 598
rect 2127 566 2131 598
rect 2091 560 2131 566
rect 3299 4318 3339 4324
rect 3299 4286 3303 4318
rect 3303 4286 3335 4318
rect 3335 4286 3339 4318
rect 3299 4250 3339 4286
rect 3299 4218 3303 4250
rect 3303 4218 3335 4250
rect 3335 4218 3339 4250
rect 3299 4182 3339 4218
rect 3299 4150 3303 4182
rect 3303 4150 3335 4182
rect 3335 4150 3339 4182
rect 3299 4114 3339 4150
rect 3299 4082 3303 4114
rect 3303 4082 3335 4114
rect 3335 4082 3339 4114
rect 3299 4046 3339 4082
rect 3299 4014 3303 4046
rect 3303 4014 3335 4046
rect 3335 4014 3339 4046
rect 3299 3978 3339 4014
rect 3299 3946 3303 3978
rect 3303 3946 3335 3978
rect 3335 3946 3339 3978
rect 3299 3910 3339 3946
rect 3299 3878 3303 3910
rect 3303 3878 3335 3910
rect 3335 3878 3339 3910
rect 3299 3842 3339 3878
rect 3299 3810 3303 3842
rect 3303 3810 3335 3842
rect 3335 3810 3339 3842
rect 3299 3774 3339 3810
rect 3299 3742 3303 3774
rect 3303 3742 3335 3774
rect 3335 3742 3339 3774
rect 3299 3706 3339 3742
rect 3299 3674 3303 3706
rect 3303 3674 3335 3706
rect 3335 3674 3339 3706
rect 3299 3638 3339 3674
rect 3299 3606 3303 3638
rect 3303 3606 3335 3638
rect 3335 3606 3339 3638
rect 3299 3570 3339 3606
rect 3299 3538 3303 3570
rect 3303 3538 3335 3570
rect 3335 3538 3339 3570
rect 3299 3502 3339 3538
rect 3299 3470 3303 3502
rect 3303 3470 3335 3502
rect 3335 3470 3339 3502
rect 3299 3464 3339 3470
rect 2956 3350 3078 3356
rect 2956 3318 3001 3350
rect 3001 3318 3033 3350
rect 3033 3318 3078 3350
rect 2956 3282 3078 3318
rect 2956 3250 3001 3282
rect 3001 3250 3033 3282
rect 3033 3250 3078 3282
rect 2956 3214 3078 3250
rect 2956 3182 3001 3214
rect 3001 3182 3033 3214
rect 3033 3182 3078 3214
rect 2956 3146 3078 3182
rect 2956 3114 3001 3146
rect 3001 3114 3033 3146
rect 3033 3114 3078 3146
rect 2956 3078 3078 3114
rect 2956 3046 3001 3078
rect 3001 3046 3033 3078
rect 3033 3046 3078 3078
rect 2956 3010 3078 3046
rect 2956 2978 3001 3010
rect 3001 2978 3033 3010
rect 3033 2978 3078 3010
rect 2956 2942 3078 2978
rect 2956 2910 3001 2942
rect 3001 2910 3033 2942
rect 3033 2910 3078 2942
rect 2956 2874 3078 2910
rect 2956 2842 3001 2874
rect 3001 2842 3033 2874
rect 3033 2842 3078 2874
rect 2956 2806 3078 2842
rect 2956 2774 3001 2806
rect 3001 2774 3033 2806
rect 3033 2774 3078 2806
rect 2956 2738 3078 2774
rect 2956 2706 3001 2738
rect 3001 2706 3033 2738
rect 3033 2706 3078 2738
rect 2956 2670 3078 2706
rect 2956 2638 3001 2670
rect 3001 2638 3033 2670
rect 3033 2638 3078 2670
rect 2956 2602 3078 2638
rect 2956 2570 3001 2602
rect 3001 2570 3033 2602
rect 3033 2570 3078 2602
rect 2956 2534 3078 2570
rect 2956 2502 3001 2534
rect 3001 2502 3033 2534
rect 3033 2502 3078 2534
rect 2956 2496 3078 2502
rect 2695 2382 2735 2388
rect 2695 2350 2699 2382
rect 2699 2350 2731 2382
rect 2731 2350 2735 2382
rect 2695 2314 2735 2350
rect 2695 2282 2699 2314
rect 2699 2282 2731 2314
rect 2731 2282 2735 2314
rect 2695 2246 2735 2282
rect 2695 2214 2699 2246
rect 2699 2214 2731 2246
rect 2731 2214 2735 2246
rect 2695 2178 2735 2214
rect 2695 2146 2699 2178
rect 2699 2146 2731 2178
rect 2731 2146 2735 2178
rect 2695 2110 2735 2146
rect 2695 2078 2699 2110
rect 2699 2078 2731 2110
rect 2731 2078 2735 2110
rect 2695 2042 2735 2078
rect 2695 2010 2699 2042
rect 2699 2010 2731 2042
rect 2731 2010 2735 2042
rect 2695 1974 2735 2010
rect 2695 1942 2699 1974
rect 2699 1942 2731 1974
rect 2731 1942 2735 1974
rect 2695 1906 2735 1942
rect 2695 1874 2699 1906
rect 2699 1874 2731 1906
rect 2731 1874 2735 1906
rect 2695 1838 2735 1874
rect 2695 1806 2699 1838
rect 2699 1806 2731 1838
rect 2731 1806 2735 1838
rect 2695 1770 2735 1806
rect 2695 1738 2699 1770
rect 2699 1738 2731 1770
rect 2731 1738 2735 1770
rect 2695 1702 2735 1738
rect 2695 1670 2699 1702
rect 2699 1670 2731 1702
rect 2731 1670 2735 1702
rect 2695 1634 2735 1670
rect 2695 1602 2699 1634
rect 2699 1602 2731 1634
rect 2731 1602 2735 1634
rect 2695 1566 2735 1602
rect 2695 1534 2699 1566
rect 2699 1534 2731 1566
rect 2731 1534 2735 1566
rect 2695 1528 2735 1534
rect 2352 1414 2474 1420
rect 2352 1382 2397 1414
rect 2397 1382 2429 1414
rect 2429 1382 2474 1414
rect 2352 1346 2474 1382
rect 2352 1314 2397 1346
rect 2397 1314 2429 1346
rect 2429 1314 2474 1346
rect 2352 1278 2474 1314
rect 2352 1246 2397 1278
rect 2397 1246 2429 1278
rect 2429 1246 2474 1278
rect 2352 1210 2474 1246
rect 2352 1178 2397 1210
rect 2397 1178 2429 1210
rect 2429 1178 2474 1210
rect 2352 1142 2474 1178
rect 2352 1110 2397 1142
rect 2397 1110 2429 1142
rect 2429 1110 2474 1142
rect 2352 1074 2474 1110
rect 2352 1042 2397 1074
rect 2397 1042 2429 1074
rect 2429 1042 2474 1074
rect 2352 1006 2474 1042
rect 2352 974 2397 1006
rect 2397 974 2429 1006
rect 2429 974 2474 1006
rect 2352 938 2474 974
rect 2352 906 2397 938
rect 2397 906 2429 938
rect 2429 906 2474 938
rect 2352 870 2474 906
rect 2352 838 2397 870
rect 2397 838 2429 870
rect 2429 838 2474 870
rect 2352 802 2474 838
rect 2352 770 2397 802
rect 2397 770 2429 802
rect 2429 770 2474 802
rect 2352 734 2474 770
rect 2352 702 2397 734
rect 2397 702 2429 734
rect 2429 702 2474 734
rect 2352 666 2474 702
rect 2352 634 2397 666
rect 2397 634 2429 666
rect 2429 634 2474 666
rect 2352 598 2474 634
rect 2352 566 2397 598
rect 2397 566 2429 598
rect 2429 566 2474 598
rect 2352 560 2474 566
rect 3560 4318 3682 4324
rect 3560 4286 3605 4318
rect 3605 4286 3637 4318
rect 3637 4286 3682 4318
rect 3560 4250 3682 4286
rect 3560 4218 3605 4250
rect 3605 4218 3637 4250
rect 3637 4218 3682 4250
rect 3560 4182 3682 4218
rect 3560 4150 3605 4182
rect 3605 4150 3637 4182
rect 3637 4150 3682 4182
rect 3560 4114 3682 4150
rect 3560 4082 3605 4114
rect 3605 4082 3637 4114
rect 3637 4082 3682 4114
rect 3560 4046 3682 4082
rect 3560 4014 3605 4046
rect 3605 4014 3637 4046
rect 3637 4014 3682 4046
rect 3560 3978 3682 4014
rect 3560 3946 3605 3978
rect 3605 3946 3637 3978
rect 3637 3946 3682 3978
rect 3560 3910 3682 3946
rect 3560 3878 3605 3910
rect 3605 3878 3637 3910
rect 3637 3878 3682 3910
rect 3560 3842 3682 3878
rect 3560 3810 3605 3842
rect 3605 3810 3637 3842
rect 3637 3810 3682 3842
rect 3560 3774 3682 3810
rect 3560 3742 3605 3774
rect 3605 3742 3637 3774
rect 3637 3742 3682 3774
rect 3560 3706 3682 3742
rect 3560 3674 3605 3706
rect 3605 3674 3637 3706
rect 3637 3674 3682 3706
rect 3560 3638 3682 3674
rect 3560 3606 3605 3638
rect 3605 3606 3637 3638
rect 3637 3606 3682 3638
rect 3560 3570 3682 3606
rect 3560 3538 3605 3570
rect 3605 3538 3637 3570
rect 3637 3538 3682 3570
rect 3560 3502 3682 3538
rect 3560 3470 3605 3502
rect 3605 3470 3637 3502
rect 3637 3470 3682 3502
rect 3560 3464 3682 3470
rect 3299 3350 3339 3356
rect 3299 3318 3303 3350
rect 3303 3318 3335 3350
rect 3335 3318 3339 3350
rect 3299 3282 3339 3318
rect 3299 3250 3303 3282
rect 3303 3250 3335 3282
rect 3335 3250 3339 3282
rect 3299 3214 3339 3250
rect 3299 3182 3303 3214
rect 3303 3182 3335 3214
rect 3335 3182 3339 3214
rect 3299 3146 3339 3182
rect 3299 3114 3303 3146
rect 3303 3114 3335 3146
rect 3335 3114 3339 3146
rect 3299 3078 3339 3114
rect 3299 3046 3303 3078
rect 3303 3046 3335 3078
rect 3335 3046 3339 3078
rect 3299 3010 3339 3046
rect 3299 2978 3303 3010
rect 3303 2978 3335 3010
rect 3335 2978 3339 3010
rect 3299 2942 3339 2978
rect 3299 2910 3303 2942
rect 3303 2910 3335 2942
rect 3335 2910 3339 2942
rect 3299 2874 3339 2910
rect 3299 2842 3303 2874
rect 3303 2842 3335 2874
rect 3335 2842 3339 2874
rect 3299 2806 3339 2842
rect 3299 2774 3303 2806
rect 3303 2774 3335 2806
rect 3335 2774 3339 2806
rect 3299 2738 3339 2774
rect 3299 2706 3303 2738
rect 3303 2706 3335 2738
rect 3335 2706 3339 2738
rect 3299 2670 3339 2706
rect 3299 2638 3303 2670
rect 3303 2638 3335 2670
rect 3335 2638 3339 2670
rect 3299 2602 3339 2638
rect 3299 2570 3303 2602
rect 3303 2570 3335 2602
rect 3335 2570 3339 2602
rect 3299 2534 3339 2570
rect 3299 2502 3303 2534
rect 3303 2502 3335 2534
rect 3335 2502 3339 2534
rect 3299 2496 3339 2502
rect 2956 2382 3078 2388
rect 2956 2350 3001 2382
rect 3001 2350 3033 2382
rect 3033 2350 3078 2382
rect 2956 2314 3078 2350
rect 2956 2282 3001 2314
rect 3001 2282 3033 2314
rect 3033 2282 3078 2314
rect 2956 2246 3078 2282
rect 2956 2214 3001 2246
rect 3001 2214 3033 2246
rect 3033 2214 3078 2246
rect 2956 2178 3078 2214
rect 2956 2146 3001 2178
rect 3001 2146 3033 2178
rect 3033 2146 3078 2178
rect 2956 2110 3078 2146
rect 2956 2078 3001 2110
rect 3001 2078 3033 2110
rect 3033 2078 3078 2110
rect 2956 2042 3078 2078
rect 2956 2010 3001 2042
rect 3001 2010 3033 2042
rect 3033 2010 3078 2042
rect 2956 1974 3078 2010
rect 2956 1942 3001 1974
rect 3001 1942 3033 1974
rect 3033 1942 3078 1974
rect 2956 1906 3078 1942
rect 2956 1874 3001 1906
rect 3001 1874 3033 1906
rect 3033 1874 3078 1906
rect 2956 1838 3078 1874
rect 2956 1806 3001 1838
rect 3001 1806 3033 1838
rect 3033 1806 3078 1838
rect 2956 1770 3078 1806
rect 2956 1738 3001 1770
rect 3001 1738 3033 1770
rect 3033 1738 3078 1770
rect 2956 1702 3078 1738
rect 2956 1670 3001 1702
rect 3001 1670 3033 1702
rect 3033 1670 3078 1702
rect 2956 1634 3078 1670
rect 2956 1602 3001 1634
rect 3001 1602 3033 1634
rect 3033 1602 3078 1634
rect 2956 1566 3078 1602
rect 2956 1534 3001 1566
rect 3001 1534 3033 1566
rect 3033 1534 3078 1566
rect 2956 1528 3078 1534
rect 2695 1414 2735 1420
rect 2695 1382 2699 1414
rect 2699 1382 2731 1414
rect 2731 1382 2735 1414
rect 2695 1346 2735 1382
rect 2695 1314 2699 1346
rect 2699 1314 2731 1346
rect 2731 1314 2735 1346
rect 2695 1278 2735 1314
rect 2695 1246 2699 1278
rect 2699 1246 2731 1278
rect 2731 1246 2735 1278
rect 2695 1210 2735 1246
rect 2695 1178 2699 1210
rect 2699 1178 2731 1210
rect 2731 1178 2735 1210
rect 2695 1142 2735 1178
rect 2695 1110 2699 1142
rect 2699 1110 2731 1142
rect 2731 1110 2735 1142
rect 2695 1074 2735 1110
rect 2695 1042 2699 1074
rect 2699 1042 2731 1074
rect 2731 1042 2735 1074
rect 2695 1006 2735 1042
rect 2695 974 2699 1006
rect 2699 974 2731 1006
rect 2731 974 2735 1006
rect 2695 938 2735 974
rect 2695 906 2699 938
rect 2699 906 2731 938
rect 2731 906 2735 938
rect 2695 870 2735 906
rect 2695 838 2699 870
rect 2699 838 2731 870
rect 2731 838 2735 870
rect 2695 802 2735 838
rect 2695 770 2699 802
rect 2699 770 2731 802
rect 2731 770 2735 802
rect 2695 734 2735 770
rect 2695 702 2699 734
rect 2699 702 2731 734
rect 2731 702 2735 734
rect 2695 666 2735 702
rect 2695 634 2699 666
rect 2699 634 2731 666
rect 2731 634 2735 666
rect 2695 598 2735 634
rect 2695 566 2699 598
rect 2699 566 2731 598
rect 2731 566 2735 598
rect 2695 560 2735 566
rect 3903 4318 3943 4324
rect 3903 4286 3907 4318
rect 3907 4286 3939 4318
rect 3939 4286 3943 4318
rect 3903 4250 3943 4286
rect 3903 4218 3907 4250
rect 3907 4218 3939 4250
rect 3939 4218 3943 4250
rect 3903 4182 3943 4218
rect 3903 4150 3907 4182
rect 3907 4150 3939 4182
rect 3939 4150 3943 4182
rect 3903 4114 3943 4150
rect 3903 4082 3907 4114
rect 3907 4082 3939 4114
rect 3939 4082 3943 4114
rect 3903 4046 3943 4082
rect 3903 4014 3907 4046
rect 3907 4014 3939 4046
rect 3939 4014 3943 4046
rect 3903 3978 3943 4014
rect 3903 3946 3907 3978
rect 3907 3946 3939 3978
rect 3939 3946 3943 3978
rect 3903 3910 3943 3946
rect 3903 3878 3907 3910
rect 3907 3878 3939 3910
rect 3939 3878 3943 3910
rect 3903 3842 3943 3878
rect 3903 3810 3907 3842
rect 3907 3810 3939 3842
rect 3939 3810 3943 3842
rect 3903 3774 3943 3810
rect 3903 3742 3907 3774
rect 3907 3742 3939 3774
rect 3939 3742 3943 3774
rect 3903 3706 3943 3742
rect 3903 3674 3907 3706
rect 3907 3674 3939 3706
rect 3939 3674 3943 3706
rect 3903 3638 3943 3674
rect 3903 3606 3907 3638
rect 3907 3606 3939 3638
rect 3939 3606 3943 3638
rect 3903 3570 3943 3606
rect 3903 3538 3907 3570
rect 3907 3538 3939 3570
rect 3939 3538 3943 3570
rect 3903 3502 3943 3538
rect 3903 3470 3907 3502
rect 3907 3470 3939 3502
rect 3939 3470 3943 3502
rect 3903 3464 3943 3470
rect 3560 3350 3682 3356
rect 3560 3318 3605 3350
rect 3605 3318 3637 3350
rect 3637 3318 3682 3350
rect 3560 3282 3682 3318
rect 3560 3250 3605 3282
rect 3605 3250 3637 3282
rect 3637 3250 3682 3282
rect 3560 3214 3682 3250
rect 3560 3182 3605 3214
rect 3605 3182 3637 3214
rect 3637 3182 3682 3214
rect 3560 3146 3682 3182
rect 3560 3114 3605 3146
rect 3605 3114 3637 3146
rect 3637 3114 3682 3146
rect 3560 3078 3682 3114
rect 3560 3046 3605 3078
rect 3605 3046 3637 3078
rect 3637 3046 3682 3078
rect 3560 3010 3682 3046
rect 3560 2978 3605 3010
rect 3605 2978 3637 3010
rect 3637 2978 3682 3010
rect 3560 2942 3682 2978
rect 3560 2910 3605 2942
rect 3605 2910 3637 2942
rect 3637 2910 3682 2942
rect 3560 2874 3682 2910
rect 3560 2842 3605 2874
rect 3605 2842 3637 2874
rect 3637 2842 3682 2874
rect 3560 2806 3682 2842
rect 3560 2774 3605 2806
rect 3605 2774 3637 2806
rect 3637 2774 3682 2806
rect 3560 2738 3682 2774
rect 3560 2706 3605 2738
rect 3605 2706 3637 2738
rect 3637 2706 3682 2738
rect 3560 2670 3682 2706
rect 3560 2638 3605 2670
rect 3605 2638 3637 2670
rect 3637 2638 3682 2670
rect 3560 2602 3682 2638
rect 3560 2570 3605 2602
rect 3605 2570 3637 2602
rect 3637 2570 3682 2602
rect 3560 2534 3682 2570
rect 3560 2502 3605 2534
rect 3605 2502 3637 2534
rect 3637 2502 3682 2534
rect 3560 2496 3682 2502
rect 3299 2382 3339 2388
rect 3299 2350 3303 2382
rect 3303 2350 3335 2382
rect 3335 2350 3339 2382
rect 3299 2314 3339 2350
rect 3299 2282 3303 2314
rect 3303 2282 3335 2314
rect 3335 2282 3339 2314
rect 3299 2246 3339 2282
rect 3299 2214 3303 2246
rect 3303 2214 3335 2246
rect 3335 2214 3339 2246
rect 3299 2178 3339 2214
rect 3299 2146 3303 2178
rect 3303 2146 3335 2178
rect 3335 2146 3339 2178
rect 3299 2110 3339 2146
rect 3299 2078 3303 2110
rect 3303 2078 3335 2110
rect 3335 2078 3339 2110
rect 3299 2042 3339 2078
rect 3299 2010 3303 2042
rect 3303 2010 3335 2042
rect 3335 2010 3339 2042
rect 3299 1974 3339 2010
rect 3299 1942 3303 1974
rect 3303 1942 3335 1974
rect 3335 1942 3339 1974
rect 3299 1906 3339 1942
rect 3299 1874 3303 1906
rect 3303 1874 3335 1906
rect 3335 1874 3339 1906
rect 3299 1838 3339 1874
rect 3299 1806 3303 1838
rect 3303 1806 3335 1838
rect 3335 1806 3339 1838
rect 3299 1770 3339 1806
rect 3299 1738 3303 1770
rect 3303 1738 3335 1770
rect 3335 1738 3339 1770
rect 3299 1702 3339 1738
rect 3299 1670 3303 1702
rect 3303 1670 3335 1702
rect 3335 1670 3339 1702
rect 3299 1634 3339 1670
rect 3299 1602 3303 1634
rect 3303 1602 3335 1634
rect 3335 1602 3339 1634
rect 3299 1566 3339 1602
rect 3299 1534 3303 1566
rect 3303 1534 3335 1566
rect 3335 1534 3339 1566
rect 3299 1528 3339 1534
rect 2956 1414 3078 1420
rect 2956 1382 3001 1414
rect 3001 1382 3033 1414
rect 3033 1382 3078 1414
rect 2956 1346 3078 1382
rect 2956 1314 3001 1346
rect 3001 1314 3033 1346
rect 3033 1314 3078 1346
rect 2956 1278 3078 1314
rect 2956 1246 3001 1278
rect 3001 1246 3033 1278
rect 3033 1246 3078 1278
rect 2956 1210 3078 1246
rect 2956 1178 3001 1210
rect 3001 1178 3033 1210
rect 3033 1178 3078 1210
rect 2956 1142 3078 1178
rect 2956 1110 3001 1142
rect 3001 1110 3033 1142
rect 3033 1110 3078 1142
rect 2956 1074 3078 1110
rect 2956 1042 3001 1074
rect 3001 1042 3033 1074
rect 3033 1042 3078 1074
rect 2956 1006 3078 1042
rect 2956 974 3001 1006
rect 3001 974 3033 1006
rect 3033 974 3078 1006
rect 2956 938 3078 974
rect 2956 906 3001 938
rect 3001 906 3033 938
rect 3033 906 3078 938
rect 2956 870 3078 906
rect 2956 838 3001 870
rect 3001 838 3033 870
rect 3033 838 3078 870
rect 2956 802 3078 838
rect 2956 770 3001 802
rect 3001 770 3033 802
rect 3033 770 3078 802
rect 2956 734 3078 770
rect 2956 702 3001 734
rect 3001 702 3033 734
rect 3033 702 3078 734
rect 2956 666 3078 702
rect 2956 634 3001 666
rect 3001 634 3033 666
rect 3033 634 3078 666
rect 2956 598 3078 634
rect 2956 566 3001 598
rect 3001 566 3033 598
rect 3033 566 3078 598
rect 2956 560 3078 566
rect 4164 4318 4286 4324
rect 4164 4286 4209 4318
rect 4209 4286 4241 4318
rect 4241 4286 4286 4318
rect 4164 4250 4286 4286
rect 4164 4218 4209 4250
rect 4209 4218 4241 4250
rect 4241 4218 4286 4250
rect 4164 4182 4286 4218
rect 4164 4150 4209 4182
rect 4209 4150 4241 4182
rect 4241 4150 4286 4182
rect 4164 4114 4286 4150
rect 4164 4082 4209 4114
rect 4209 4082 4241 4114
rect 4241 4082 4286 4114
rect 4164 4046 4286 4082
rect 4164 4014 4209 4046
rect 4209 4014 4241 4046
rect 4241 4014 4286 4046
rect 4164 3978 4286 4014
rect 4164 3946 4209 3978
rect 4209 3946 4241 3978
rect 4241 3946 4286 3978
rect 4164 3910 4286 3946
rect 4164 3878 4209 3910
rect 4209 3878 4241 3910
rect 4241 3878 4286 3910
rect 4164 3842 4286 3878
rect 4164 3810 4209 3842
rect 4209 3810 4241 3842
rect 4241 3810 4286 3842
rect 4164 3774 4286 3810
rect 4164 3742 4209 3774
rect 4209 3742 4241 3774
rect 4241 3742 4286 3774
rect 4164 3706 4286 3742
rect 4164 3674 4209 3706
rect 4209 3674 4241 3706
rect 4241 3674 4286 3706
rect 4164 3638 4286 3674
rect 4164 3606 4209 3638
rect 4209 3606 4241 3638
rect 4241 3606 4286 3638
rect 4164 3570 4286 3606
rect 4164 3538 4209 3570
rect 4209 3538 4241 3570
rect 4241 3538 4286 3570
rect 4164 3502 4286 3538
rect 4164 3470 4209 3502
rect 4209 3470 4241 3502
rect 4241 3470 4286 3502
rect 4164 3464 4286 3470
rect 3903 3350 3943 3356
rect 3903 3318 3907 3350
rect 3907 3318 3939 3350
rect 3939 3318 3943 3350
rect 3903 3282 3943 3318
rect 3903 3250 3907 3282
rect 3907 3250 3939 3282
rect 3939 3250 3943 3282
rect 3903 3214 3943 3250
rect 3903 3182 3907 3214
rect 3907 3182 3939 3214
rect 3939 3182 3943 3214
rect 3903 3146 3943 3182
rect 3903 3114 3907 3146
rect 3907 3114 3939 3146
rect 3939 3114 3943 3146
rect 3903 3078 3943 3114
rect 3903 3046 3907 3078
rect 3907 3046 3939 3078
rect 3939 3046 3943 3078
rect 3903 3010 3943 3046
rect 3903 2978 3907 3010
rect 3907 2978 3939 3010
rect 3939 2978 3943 3010
rect 3903 2942 3943 2978
rect 3903 2910 3907 2942
rect 3907 2910 3939 2942
rect 3939 2910 3943 2942
rect 3903 2874 3943 2910
rect 3903 2842 3907 2874
rect 3907 2842 3939 2874
rect 3939 2842 3943 2874
rect 3903 2806 3943 2842
rect 3903 2774 3907 2806
rect 3907 2774 3939 2806
rect 3939 2774 3943 2806
rect 3903 2738 3943 2774
rect 3903 2706 3907 2738
rect 3907 2706 3939 2738
rect 3939 2706 3943 2738
rect 3903 2670 3943 2706
rect 3903 2638 3907 2670
rect 3907 2638 3939 2670
rect 3939 2638 3943 2670
rect 3903 2602 3943 2638
rect 3903 2570 3907 2602
rect 3907 2570 3939 2602
rect 3939 2570 3943 2602
rect 3903 2534 3943 2570
rect 3903 2502 3907 2534
rect 3907 2502 3939 2534
rect 3939 2502 3943 2534
rect 3903 2496 3943 2502
rect 3560 2382 3682 2388
rect 3560 2350 3605 2382
rect 3605 2350 3637 2382
rect 3637 2350 3682 2382
rect 3560 2314 3682 2350
rect 3560 2282 3605 2314
rect 3605 2282 3637 2314
rect 3637 2282 3682 2314
rect 3560 2246 3682 2282
rect 3560 2214 3605 2246
rect 3605 2214 3637 2246
rect 3637 2214 3682 2246
rect 3560 2178 3682 2214
rect 3560 2146 3605 2178
rect 3605 2146 3637 2178
rect 3637 2146 3682 2178
rect 3560 2110 3682 2146
rect 3560 2078 3605 2110
rect 3605 2078 3637 2110
rect 3637 2078 3682 2110
rect 3560 2042 3682 2078
rect 3560 2010 3605 2042
rect 3605 2010 3637 2042
rect 3637 2010 3682 2042
rect 3560 1974 3682 2010
rect 3560 1942 3605 1974
rect 3605 1942 3637 1974
rect 3637 1942 3682 1974
rect 3560 1906 3682 1942
rect 3560 1874 3605 1906
rect 3605 1874 3637 1906
rect 3637 1874 3682 1906
rect 3560 1838 3682 1874
rect 3560 1806 3605 1838
rect 3605 1806 3637 1838
rect 3637 1806 3682 1838
rect 3560 1770 3682 1806
rect 3560 1738 3605 1770
rect 3605 1738 3637 1770
rect 3637 1738 3682 1770
rect 3560 1702 3682 1738
rect 3560 1670 3605 1702
rect 3605 1670 3637 1702
rect 3637 1670 3682 1702
rect 3560 1634 3682 1670
rect 3560 1602 3605 1634
rect 3605 1602 3637 1634
rect 3637 1602 3682 1634
rect 3560 1566 3682 1602
rect 3560 1534 3605 1566
rect 3605 1534 3637 1566
rect 3637 1534 3682 1566
rect 3560 1528 3682 1534
rect 3299 1414 3339 1420
rect 3299 1382 3303 1414
rect 3303 1382 3335 1414
rect 3335 1382 3339 1414
rect 3299 1346 3339 1382
rect 3299 1314 3303 1346
rect 3303 1314 3335 1346
rect 3335 1314 3339 1346
rect 3299 1278 3339 1314
rect 3299 1246 3303 1278
rect 3303 1246 3335 1278
rect 3335 1246 3339 1278
rect 3299 1210 3339 1246
rect 3299 1178 3303 1210
rect 3303 1178 3335 1210
rect 3335 1178 3339 1210
rect 3299 1142 3339 1178
rect 3299 1110 3303 1142
rect 3303 1110 3335 1142
rect 3335 1110 3339 1142
rect 3299 1074 3339 1110
rect 3299 1042 3303 1074
rect 3303 1042 3335 1074
rect 3335 1042 3339 1074
rect 3299 1006 3339 1042
rect 3299 974 3303 1006
rect 3303 974 3335 1006
rect 3335 974 3339 1006
rect 3299 938 3339 974
rect 3299 906 3303 938
rect 3303 906 3335 938
rect 3335 906 3339 938
rect 3299 870 3339 906
rect 3299 838 3303 870
rect 3303 838 3335 870
rect 3335 838 3339 870
rect 3299 802 3339 838
rect 3299 770 3303 802
rect 3303 770 3335 802
rect 3335 770 3339 802
rect 3299 734 3339 770
rect 3299 702 3303 734
rect 3303 702 3335 734
rect 3335 702 3339 734
rect 3299 666 3339 702
rect 3299 634 3303 666
rect 3303 634 3335 666
rect 3335 634 3339 666
rect 3299 598 3339 634
rect 3299 566 3303 598
rect 3303 566 3335 598
rect 3335 566 3339 598
rect 3299 560 3339 566
rect 4507 4318 4547 4324
rect 4507 4286 4511 4318
rect 4511 4286 4543 4318
rect 4543 4286 4547 4318
rect 4507 4250 4547 4286
rect 4507 4218 4511 4250
rect 4511 4218 4543 4250
rect 4543 4218 4547 4250
rect 4507 4182 4547 4218
rect 4507 4150 4511 4182
rect 4511 4150 4543 4182
rect 4543 4150 4547 4182
rect 4507 4114 4547 4150
rect 4507 4082 4511 4114
rect 4511 4082 4543 4114
rect 4543 4082 4547 4114
rect 4507 4046 4547 4082
rect 4507 4014 4511 4046
rect 4511 4014 4543 4046
rect 4543 4014 4547 4046
rect 4507 3978 4547 4014
rect 4507 3946 4511 3978
rect 4511 3946 4543 3978
rect 4543 3946 4547 3978
rect 4507 3910 4547 3946
rect 4507 3878 4511 3910
rect 4511 3878 4543 3910
rect 4543 3878 4547 3910
rect 4507 3842 4547 3878
rect 4507 3810 4511 3842
rect 4511 3810 4543 3842
rect 4543 3810 4547 3842
rect 4507 3774 4547 3810
rect 4507 3742 4511 3774
rect 4511 3742 4543 3774
rect 4543 3742 4547 3774
rect 4507 3706 4547 3742
rect 4507 3674 4511 3706
rect 4511 3674 4543 3706
rect 4543 3674 4547 3706
rect 4507 3638 4547 3674
rect 4507 3606 4511 3638
rect 4511 3606 4543 3638
rect 4543 3606 4547 3638
rect 4507 3570 4547 3606
rect 4507 3538 4511 3570
rect 4511 3538 4543 3570
rect 4543 3538 4547 3570
rect 4507 3502 4547 3538
rect 4507 3470 4511 3502
rect 4511 3470 4543 3502
rect 4543 3470 4547 3502
rect 4507 3464 4547 3470
rect 4164 3350 4286 3356
rect 4164 3318 4209 3350
rect 4209 3318 4241 3350
rect 4241 3318 4286 3350
rect 4164 3282 4286 3318
rect 4164 3250 4209 3282
rect 4209 3250 4241 3282
rect 4241 3250 4286 3282
rect 4164 3214 4286 3250
rect 4164 3182 4209 3214
rect 4209 3182 4241 3214
rect 4241 3182 4286 3214
rect 4164 3146 4286 3182
rect 4164 3114 4209 3146
rect 4209 3114 4241 3146
rect 4241 3114 4286 3146
rect 4164 3078 4286 3114
rect 4164 3046 4209 3078
rect 4209 3046 4241 3078
rect 4241 3046 4286 3078
rect 4164 3010 4286 3046
rect 4164 2978 4209 3010
rect 4209 2978 4241 3010
rect 4241 2978 4286 3010
rect 4164 2942 4286 2978
rect 4164 2910 4209 2942
rect 4209 2910 4241 2942
rect 4241 2910 4286 2942
rect 4164 2874 4286 2910
rect 4164 2842 4209 2874
rect 4209 2842 4241 2874
rect 4241 2842 4286 2874
rect 4164 2806 4286 2842
rect 4164 2774 4209 2806
rect 4209 2774 4241 2806
rect 4241 2774 4286 2806
rect 4164 2738 4286 2774
rect 4164 2706 4209 2738
rect 4209 2706 4241 2738
rect 4241 2706 4286 2738
rect 4164 2670 4286 2706
rect 4164 2638 4209 2670
rect 4209 2638 4241 2670
rect 4241 2638 4286 2670
rect 4164 2602 4286 2638
rect 4164 2570 4209 2602
rect 4209 2570 4241 2602
rect 4241 2570 4286 2602
rect 4164 2534 4286 2570
rect 4164 2502 4209 2534
rect 4209 2502 4241 2534
rect 4241 2502 4286 2534
rect 4164 2496 4286 2502
rect 3903 2382 3943 2388
rect 3903 2350 3907 2382
rect 3907 2350 3939 2382
rect 3939 2350 3943 2382
rect 3903 2314 3943 2350
rect 3903 2282 3907 2314
rect 3907 2282 3939 2314
rect 3939 2282 3943 2314
rect 3903 2246 3943 2282
rect 3903 2214 3907 2246
rect 3907 2214 3939 2246
rect 3939 2214 3943 2246
rect 3903 2178 3943 2214
rect 3903 2146 3907 2178
rect 3907 2146 3939 2178
rect 3939 2146 3943 2178
rect 3903 2110 3943 2146
rect 3903 2078 3907 2110
rect 3907 2078 3939 2110
rect 3939 2078 3943 2110
rect 3903 2042 3943 2078
rect 3903 2010 3907 2042
rect 3907 2010 3939 2042
rect 3939 2010 3943 2042
rect 3903 1974 3943 2010
rect 3903 1942 3907 1974
rect 3907 1942 3939 1974
rect 3939 1942 3943 1974
rect 3903 1906 3943 1942
rect 3903 1874 3907 1906
rect 3907 1874 3939 1906
rect 3939 1874 3943 1906
rect 3903 1838 3943 1874
rect 3903 1806 3907 1838
rect 3907 1806 3939 1838
rect 3939 1806 3943 1838
rect 3903 1770 3943 1806
rect 3903 1738 3907 1770
rect 3907 1738 3939 1770
rect 3939 1738 3943 1770
rect 3903 1702 3943 1738
rect 3903 1670 3907 1702
rect 3907 1670 3939 1702
rect 3939 1670 3943 1702
rect 3903 1634 3943 1670
rect 3903 1602 3907 1634
rect 3907 1602 3939 1634
rect 3939 1602 3943 1634
rect 3903 1566 3943 1602
rect 3903 1534 3907 1566
rect 3907 1534 3939 1566
rect 3939 1534 3943 1566
rect 3903 1528 3943 1534
rect 3560 1414 3682 1420
rect 3560 1382 3605 1414
rect 3605 1382 3637 1414
rect 3637 1382 3682 1414
rect 3560 1346 3682 1382
rect 3560 1314 3605 1346
rect 3605 1314 3637 1346
rect 3637 1314 3682 1346
rect 3560 1278 3682 1314
rect 3560 1246 3605 1278
rect 3605 1246 3637 1278
rect 3637 1246 3682 1278
rect 3560 1210 3682 1246
rect 3560 1178 3605 1210
rect 3605 1178 3637 1210
rect 3637 1178 3682 1210
rect 3560 1142 3682 1178
rect 3560 1110 3605 1142
rect 3605 1110 3637 1142
rect 3637 1110 3682 1142
rect 3560 1074 3682 1110
rect 3560 1042 3605 1074
rect 3605 1042 3637 1074
rect 3637 1042 3682 1074
rect 3560 1006 3682 1042
rect 3560 974 3605 1006
rect 3605 974 3637 1006
rect 3637 974 3682 1006
rect 3560 938 3682 974
rect 3560 906 3605 938
rect 3605 906 3637 938
rect 3637 906 3682 938
rect 3560 870 3682 906
rect 3560 838 3605 870
rect 3605 838 3637 870
rect 3637 838 3682 870
rect 3560 802 3682 838
rect 3560 770 3605 802
rect 3605 770 3637 802
rect 3637 770 3682 802
rect 3560 734 3682 770
rect 3560 702 3605 734
rect 3605 702 3637 734
rect 3637 702 3682 734
rect 3560 666 3682 702
rect 3560 634 3605 666
rect 3605 634 3637 666
rect 3637 634 3682 666
rect 3560 598 3682 634
rect 3560 566 3605 598
rect 3605 566 3637 598
rect 3637 566 3682 598
rect 3560 560 3682 566
rect 4768 4318 4890 4324
rect 4768 4286 4813 4318
rect 4813 4286 4845 4318
rect 4845 4286 4890 4318
rect 4768 4250 4890 4286
rect 4768 4218 4813 4250
rect 4813 4218 4845 4250
rect 4845 4218 4890 4250
rect 4768 4182 4890 4218
rect 4768 4150 4813 4182
rect 4813 4150 4845 4182
rect 4845 4150 4890 4182
rect 4768 4114 4890 4150
rect 4768 4082 4813 4114
rect 4813 4082 4845 4114
rect 4845 4082 4890 4114
rect 4768 4046 4890 4082
rect 4768 4014 4813 4046
rect 4813 4014 4845 4046
rect 4845 4014 4890 4046
rect 4768 3978 4890 4014
rect 4768 3946 4813 3978
rect 4813 3946 4845 3978
rect 4845 3946 4890 3978
rect 4768 3910 4890 3946
rect 4768 3878 4813 3910
rect 4813 3878 4845 3910
rect 4845 3878 4890 3910
rect 4768 3842 4890 3878
rect 4768 3810 4813 3842
rect 4813 3810 4845 3842
rect 4845 3810 4890 3842
rect 4768 3774 4890 3810
rect 4768 3742 4813 3774
rect 4813 3742 4845 3774
rect 4845 3742 4890 3774
rect 4768 3706 4890 3742
rect 4768 3674 4813 3706
rect 4813 3674 4845 3706
rect 4845 3674 4890 3706
rect 4768 3638 4890 3674
rect 4768 3606 4813 3638
rect 4813 3606 4845 3638
rect 4845 3606 4890 3638
rect 4768 3570 4890 3606
rect 4768 3538 4813 3570
rect 4813 3538 4845 3570
rect 4845 3538 4890 3570
rect 4768 3502 4890 3538
rect 4768 3470 4813 3502
rect 4813 3470 4845 3502
rect 4845 3470 4890 3502
rect 4768 3464 4890 3470
rect 4507 3350 4547 3356
rect 4507 3318 4511 3350
rect 4511 3318 4543 3350
rect 4543 3318 4547 3350
rect 4507 3282 4547 3318
rect 4507 3250 4511 3282
rect 4511 3250 4543 3282
rect 4543 3250 4547 3282
rect 4507 3214 4547 3250
rect 4507 3182 4511 3214
rect 4511 3182 4543 3214
rect 4543 3182 4547 3214
rect 4507 3146 4547 3182
rect 4507 3114 4511 3146
rect 4511 3114 4543 3146
rect 4543 3114 4547 3146
rect 4507 3078 4547 3114
rect 4507 3046 4511 3078
rect 4511 3046 4543 3078
rect 4543 3046 4547 3078
rect 4507 3010 4547 3046
rect 4507 2978 4511 3010
rect 4511 2978 4543 3010
rect 4543 2978 4547 3010
rect 4507 2942 4547 2978
rect 4507 2910 4511 2942
rect 4511 2910 4543 2942
rect 4543 2910 4547 2942
rect 4507 2874 4547 2910
rect 4507 2842 4511 2874
rect 4511 2842 4543 2874
rect 4543 2842 4547 2874
rect 4507 2806 4547 2842
rect 4507 2774 4511 2806
rect 4511 2774 4543 2806
rect 4543 2774 4547 2806
rect 4507 2738 4547 2774
rect 4507 2706 4511 2738
rect 4511 2706 4543 2738
rect 4543 2706 4547 2738
rect 4507 2670 4547 2706
rect 4507 2638 4511 2670
rect 4511 2638 4543 2670
rect 4543 2638 4547 2670
rect 4507 2602 4547 2638
rect 4507 2570 4511 2602
rect 4511 2570 4543 2602
rect 4543 2570 4547 2602
rect 4507 2534 4547 2570
rect 4507 2502 4511 2534
rect 4511 2502 4543 2534
rect 4543 2502 4547 2534
rect 4507 2496 4547 2502
rect 4164 2382 4286 2388
rect 4164 2350 4209 2382
rect 4209 2350 4241 2382
rect 4241 2350 4286 2382
rect 4164 2314 4286 2350
rect 4164 2282 4209 2314
rect 4209 2282 4241 2314
rect 4241 2282 4286 2314
rect 4164 2246 4286 2282
rect 4164 2214 4209 2246
rect 4209 2214 4241 2246
rect 4241 2214 4286 2246
rect 4164 2178 4286 2214
rect 4164 2146 4209 2178
rect 4209 2146 4241 2178
rect 4241 2146 4286 2178
rect 4164 2110 4286 2146
rect 4164 2078 4209 2110
rect 4209 2078 4241 2110
rect 4241 2078 4286 2110
rect 4164 2042 4286 2078
rect 4164 2010 4209 2042
rect 4209 2010 4241 2042
rect 4241 2010 4286 2042
rect 4164 1974 4286 2010
rect 4164 1942 4209 1974
rect 4209 1942 4241 1974
rect 4241 1942 4286 1974
rect 4164 1906 4286 1942
rect 4164 1874 4209 1906
rect 4209 1874 4241 1906
rect 4241 1874 4286 1906
rect 4164 1838 4286 1874
rect 4164 1806 4209 1838
rect 4209 1806 4241 1838
rect 4241 1806 4286 1838
rect 4164 1770 4286 1806
rect 4164 1738 4209 1770
rect 4209 1738 4241 1770
rect 4241 1738 4286 1770
rect 4164 1702 4286 1738
rect 4164 1670 4209 1702
rect 4209 1670 4241 1702
rect 4241 1670 4286 1702
rect 4164 1634 4286 1670
rect 4164 1602 4209 1634
rect 4209 1602 4241 1634
rect 4241 1602 4286 1634
rect 4164 1566 4286 1602
rect 4164 1534 4209 1566
rect 4209 1534 4241 1566
rect 4241 1534 4286 1566
rect 4164 1528 4286 1534
rect 3903 1414 3943 1420
rect 3903 1382 3907 1414
rect 3907 1382 3939 1414
rect 3939 1382 3943 1414
rect 3903 1346 3943 1382
rect 3903 1314 3907 1346
rect 3907 1314 3939 1346
rect 3939 1314 3943 1346
rect 3903 1278 3943 1314
rect 3903 1246 3907 1278
rect 3907 1246 3939 1278
rect 3939 1246 3943 1278
rect 3903 1210 3943 1246
rect 3903 1178 3907 1210
rect 3907 1178 3939 1210
rect 3939 1178 3943 1210
rect 3903 1142 3943 1178
rect 3903 1110 3907 1142
rect 3907 1110 3939 1142
rect 3939 1110 3943 1142
rect 3903 1074 3943 1110
rect 3903 1042 3907 1074
rect 3907 1042 3939 1074
rect 3939 1042 3943 1074
rect 3903 1006 3943 1042
rect 3903 974 3907 1006
rect 3907 974 3939 1006
rect 3939 974 3943 1006
rect 3903 938 3943 974
rect 3903 906 3907 938
rect 3907 906 3939 938
rect 3939 906 3943 938
rect 3903 870 3943 906
rect 3903 838 3907 870
rect 3907 838 3939 870
rect 3939 838 3943 870
rect 3903 802 3943 838
rect 3903 770 3907 802
rect 3907 770 3939 802
rect 3939 770 3943 802
rect 3903 734 3943 770
rect 3903 702 3907 734
rect 3907 702 3939 734
rect 3939 702 3943 734
rect 3903 666 3943 702
rect 3903 634 3907 666
rect 3907 634 3939 666
rect 3939 634 3943 666
rect 3903 598 3943 634
rect 3903 566 3907 598
rect 3907 566 3939 598
rect 3939 566 3943 598
rect 3903 560 3943 566
rect 5111 4318 5151 4324
rect 5111 4286 5115 4318
rect 5115 4286 5147 4318
rect 5147 4286 5151 4318
rect 5111 4250 5151 4286
rect 5111 4218 5115 4250
rect 5115 4218 5147 4250
rect 5147 4218 5151 4250
rect 5111 4182 5151 4218
rect 5111 4150 5115 4182
rect 5115 4150 5147 4182
rect 5147 4150 5151 4182
rect 5111 4114 5151 4150
rect 5111 4082 5115 4114
rect 5115 4082 5147 4114
rect 5147 4082 5151 4114
rect 5111 4046 5151 4082
rect 5111 4014 5115 4046
rect 5115 4014 5147 4046
rect 5147 4014 5151 4046
rect 5111 3978 5151 4014
rect 5111 3946 5115 3978
rect 5115 3946 5147 3978
rect 5147 3946 5151 3978
rect 5111 3910 5151 3946
rect 5111 3878 5115 3910
rect 5115 3878 5147 3910
rect 5147 3878 5151 3910
rect 5111 3842 5151 3878
rect 5111 3810 5115 3842
rect 5115 3810 5147 3842
rect 5147 3810 5151 3842
rect 5111 3774 5151 3810
rect 5111 3742 5115 3774
rect 5115 3742 5147 3774
rect 5147 3742 5151 3774
rect 5111 3706 5151 3742
rect 5111 3674 5115 3706
rect 5115 3674 5147 3706
rect 5147 3674 5151 3706
rect 5111 3638 5151 3674
rect 5111 3606 5115 3638
rect 5115 3606 5147 3638
rect 5147 3606 5151 3638
rect 5111 3570 5151 3606
rect 5111 3538 5115 3570
rect 5115 3538 5147 3570
rect 5147 3538 5151 3570
rect 5111 3502 5151 3538
rect 5111 3470 5115 3502
rect 5115 3470 5147 3502
rect 5147 3470 5151 3502
rect 5111 3464 5151 3470
rect 4768 3350 4890 3356
rect 4768 3318 4813 3350
rect 4813 3318 4845 3350
rect 4845 3318 4890 3350
rect 4768 3282 4890 3318
rect 4768 3250 4813 3282
rect 4813 3250 4845 3282
rect 4845 3250 4890 3282
rect 4768 3214 4890 3250
rect 4768 3182 4813 3214
rect 4813 3182 4845 3214
rect 4845 3182 4890 3214
rect 4768 3146 4890 3182
rect 4768 3114 4813 3146
rect 4813 3114 4845 3146
rect 4845 3114 4890 3146
rect 4768 3078 4890 3114
rect 4768 3046 4813 3078
rect 4813 3046 4845 3078
rect 4845 3046 4890 3078
rect 4768 3010 4890 3046
rect 4768 2978 4813 3010
rect 4813 2978 4845 3010
rect 4845 2978 4890 3010
rect 4768 2942 4890 2978
rect 4768 2910 4813 2942
rect 4813 2910 4845 2942
rect 4845 2910 4890 2942
rect 4768 2874 4890 2910
rect 4768 2842 4813 2874
rect 4813 2842 4845 2874
rect 4845 2842 4890 2874
rect 4768 2806 4890 2842
rect 4768 2774 4813 2806
rect 4813 2774 4845 2806
rect 4845 2774 4890 2806
rect 4768 2738 4890 2774
rect 4768 2706 4813 2738
rect 4813 2706 4845 2738
rect 4845 2706 4890 2738
rect 4768 2670 4890 2706
rect 4768 2638 4813 2670
rect 4813 2638 4845 2670
rect 4845 2638 4890 2670
rect 4768 2602 4890 2638
rect 4768 2570 4813 2602
rect 4813 2570 4845 2602
rect 4845 2570 4890 2602
rect 4768 2534 4890 2570
rect 4768 2502 4813 2534
rect 4813 2502 4845 2534
rect 4845 2502 4890 2534
rect 4768 2496 4890 2502
rect 4507 2382 4547 2388
rect 4507 2350 4511 2382
rect 4511 2350 4543 2382
rect 4543 2350 4547 2382
rect 4507 2314 4547 2350
rect 4507 2282 4511 2314
rect 4511 2282 4543 2314
rect 4543 2282 4547 2314
rect 4507 2246 4547 2282
rect 4507 2214 4511 2246
rect 4511 2214 4543 2246
rect 4543 2214 4547 2246
rect 4507 2178 4547 2214
rect 4507 2146 4511 2178
rect 4511 2146 4543 2178
rect 4543 2146 4547 2178
rect 4507 2110 4547 2146
rect 4507 2078 4511 2110
rect 4511 2078 4543 2110
rect 4543 2078 4547 2110
rect 4507 2042 4547 2078
rect 4507 2010 4511 2042
rect 4511 2010 4543 2042
rect 4543 2010 4547 2042
rect 4507 1974 4547 2010
rect 4507 1942 4511 1974
rect 4511 1942 4543 1974
rect 4543 1942 4547 1974
rect 4507 1906 4547 1942
rect 4507 1874 4511 1906
rect 4511 1874 4543 1906
rect 4543 1874 4547 1906
rect 4507 1838 4547 1874
rect 4507 1806 4511 1838
rect 4511 1806 4543 1838
rect 4543 1806 4547 1838
rect 4507 1770 4547 1806
rect 4507 1738 4511 1770
rect 4511 1738 4543 1770
rect 4543 1738 4547 1770
rect 4507 1702 4547 1738
rect 4507 1670 4511 1702
rect 4511 1670 4543 1702
rect 4543 1670 4547 1702
rect 4507 1634 4547 1670
rect 4507 1602 4511 1634
rect 4511 1602 4543 1634
rect 4543 1602 4547 1634
rect 4507 1566 4547 1602
rect 4507 1534 4511 1566
rect 4511 1534 4543 1566
rect 4543 1534 4547 1566
rect 4507 1528 4547 1534
rect 4164 1414 4286 1420
rect 4164 1382 4209 1414
rect 4209 1382 4241 1414
rect 4241 1382 4286 1414
rect 4164 1346 4286 1382
rect 4164 1314 4209 1346
rect 4209 1314 4241 1346
rect 4241 1314 4286 1346
rect 4164 1278 4286 1314
rect 4164 1246 4209 1278
rect 4209 1246 4241 1278
rect 4241 1246 4286 1278
rect 4164 1210 4286 1246
rect 4164 1178 4209 1210
rect 4209 1178 4241 1210
rect 4241 1178 4286 1210
rect 4164 1142 4286 1178
rect 4164 1110 4209 1142
rect 4209 1110 4241 1142
rect 4241 1110 4286 1142
rect 4164 1074 4286 1110
rect 4164 1042 4209 1074
rect 4209 1042 4241 1074
rect 4241 1042 4286 1074
rect 4164 1006 4286 1042
rect 4164 974 4209 1006
rect 4209 974 4241 1006
rect 4241 974 4286 1006
rect 4164 938 4286 974
rect 4164 906 4209 938
rect 4209 906 4241 938
rect 4241 906 4286 938
rect 4164 870 4286 906
rect 4164 838 4209 870
rect 4209 838 4241 870
rect 4241 838 4286 870
rect 4164 802 4286 838
rect 4164 770 4209 802
rect 4209 770 4241 802
rect 4241 770 4286 802
rect 4164 734 4286 770
rect 4164 702 4209 734
rect 4209 702 4241 734
rect 4241 702 4286 734
rect 4164 666 4286 702
rect 4164 634 4209 666
rect 4209 634 4241 666
rect 4241 634 4286 666
rect 4164 598 4286 634
rect 4164 566 4209 598
rect 4209 566 4241 598
rect 4241 566 4286 598
rect 4164 560 4286 566
rect 5372 4318 5494 4324
rect 5372 4286 5417 4318
rect 5417 4286 5449 4318
rect 5449 4286 5494 4318
rect 5372 4250 5494 4286
rect 5372 4218 5417 4250
rect 5417 4218 5449 4250
rect 5449 4218 5494 4250
rect 5372 4182 5494 4218
rect 5372 4150 5417 4182
rect 5417 4150 5449 4182
rect 5449 4150 5494 4182
rect 5372 4114 5494 4150
rect 5372 4082 5417 4114
rect 5417 4082 5449 4114
rect 5449 4082 5494 4114
rect 5372 4046 5494 4082
rect 5372 4014 5417 4046
rect 5417 4014 5449 4046
rect 5449 4014 5494 4046
rect 5372 3978 5494 4014
rect 5372 3946 5417 3978
rect 5417 3946 5449 3978
rect 5449 3946 5494 3978
rect 5372 3910 5494 3946
rect 5372 3878 5417 3910
rect 5417 3878 5449 3910
rect 5449 3878 5494 3910
rect 5372 3842 5494 3878
rect 5372 3810 5417 3842
rect 5417 3810 5449 3842
rect 5449 3810 5494 3842
rect 5372 3774 5494 3810
rect 5372 3742 5417 3774
rect 5417 3742 5449 3774
rect 5449 3742 5494 3774
rect 5372 3706 5494 3742
rect 5372 3674 5417 3706
rect 5417 3674 5449 3706
rect 5449 3674 5494 3706
rect 5372 3638 5494 3674
rect 5372 3606 5417 3638
rect 5417 3606 5449 3638
rect 5449 3606 5494 3638
rect 5372 3570 5494 3606
rect 5372 3538 5417 3570
rect 5417 3538 5449 3570
rect 5449 3538 5494 3570
rect 5372 3502 5494 3538
rect 5372 3470 5417 3502
rect 5417 3470 5449 3502
rect 5449 3470 5494 3502
rect 5372 3464 5494 3470
rect 5111 3350 5151 3356
rect 5111 3318 5115 3350
rect 5115 3318 5147 3350
rect 5147 3318 5151 3350
rect 5111 3282 5151 3318
rect 5111 3250 5115 3282
rect 5115 3250 5147 3282
rect 5147 3250 5151 3282
rect 5111 3214 5151 3250
rect 5111 3182 5115 3214
rect 5115 3182 5147 3214
rect 5147 3182 5151 3214
rect 5111 3146 5151 3182
rect 5111 3114 5115 3146
rect 5115 3114 5147 3146
rect 5147 3114 5151 3146
rect 5111 3078 5151 3114
rect 5111 3046 5115 3078
rect 5115 3046 5147 3078
rect 5147 3046 5151 3078
rect 5111 3010 5151 3046
rect 5111 2978 5115 3010
rect 5115 2978 5147 3010
rect 5147 2978 5151 3010
rect 5111 2942 5151 2978
rect 5111 2910 5115 2942
rect 5115 2910 5147 2942
rect 5147 2910 5151 2942
rect 5111 2874 5151 2910
rect 5111 2842 5115 2874
rect 5115 2842 5147 2874
rect 5147 2842 5151 2874
rect 5111 2806 5151 2842
rect 5111 2774 5115 2806
rect 5115 2774 5147 2806
rect 5147 2774 5151 2806
rect 5111 2738 5151 2774
rect 5111 2706 5115 2738
rect 5115 2706 5147 2738
rect 5147 2706 5151 2738
rect 5111 2670 5151 2706
rect 5111 2638 5115 2670
rect 5115 2638 5147 2670
rect 5147 2638 5151 2670
rect 5111 2602 5151 2638
rect 5111 2570 5115 2602
rect 5115 2570 5147 2602
rect 5147 2570 5151 2602
rect 5111 2534 5151 2570
rect 5111 2502 5115 2534
rect 5115 2502 5147 2534
rect 5147 2502 5151 2534
rect 5111 2496 5151 2502
rect 4768 2382 4890 2388
rect 4768 2350 4813 2382
rect 4813 2350 4845 2382
rect 4845 2350 4890 2382
rect 4768 2314 4890 2350
rect 4768 2282 4813 2314
rect 4813 2282 4845 2314
rect 4845 2282 4890 2314
rect 4768 2246 4890 2282
rect 4768 2214 4813 2246
rect 4813 2214 4845 2246
rect 4845 2214 4890 2246
rect 4768 2178 4890 2214
rect 4768 2146 4813 2178
rect 4813 2146 4845 2178
rect 4845 2146 4890 2178
rect 4768 2110 4890 2146
rect 4768 2078 4813 2110
rect 4813 2078 4845 2110
rect 4845 2078 4890 2110
rect 4768 2042 4890 2078
rect 4768 2010 4813 2042
rect 4813 2010 4845 2042
rect 4845 2010 4890 2042
rect 4768 1974 4890 2010
rect 4768 1942 4813 1974
rect 4813 1942 4845 1974
rect 4845 1942 4890 1974
rect 4768 1906 4890 1942
rect 4768 1874 4813 1906
rect 4813 1874 4845 1906
rect 4845 1874 4890 1906
rect 4768 1838 4890 1874
rect 4768 1806 4813 1838
rect 4813 1806 4845 1838
rect 4845 1806 4890 1838
rect 4768 1770 4890 1806
rect 4768 1738 4813 1770
rect 4813 1738 4845 1770
rect 4845 1738 4890 1770
rect 4768 1702 4890 1738
rect 4768 1670 4813 1702
rect 4813 1670 4845 1702
rect 4845 1670 4890 1702
rect 4768 1634 4890 1670
rect 4768 1602 4813 1634
rect 4813 1602 4845 1634
rect 4845 1602 4890 1634
rect 4768 1566 4890 1602
rect 4768 1534 4813 1566
rect 4813 1534 4845 1566
rect 4845 1534 4890 1566
rect 4768 1528 4890 1534
rect 4507 1414 4547 1420
rect 4507 1382 4511 1414
rect 4511 1382 4543 1414
rect 4543 1382 4547 1414
rect 4507 1346 4547 1382
rect 4507 1314 4511 1346
rect 4511 1314 4543 1346
rect 4543 1314 4547 1346
rect 4507 1278 4547 1314
rect 4507 1246 4511 1278
rect 4511 1246 4543 1278
rect 4543 1246 4547 1278
rect 4507 1210 4547 1246
rect 4507 1178 4511 1210
rect 4511 1178 4543 1210
rect 4543 1178 4547 1210
rect 4507 1142 4547 1178
rect 4507 1110 4511 1142
rect 4511 1110 4543 1142
rect 4543 1110 4547 1142
rect 4507 1074 4547 1110
rect 4507 1042 4511 1074
rect 4511 1042 4543 1074
rect 4543 1042 4547 1074
rect 4507 1006 4547 1042
rect 4507 974 4511 1006
rect 4511 974 4543 1006
rect 4543 974 4547 1006
rect 4507 938 4547 974
rect 4507 906 4511 938
rect 4511 906 4543 938
rect 4543 906 4547 938
rect 4507 870 4547 906
rect 4507 838 4511 870
rect 4511 838 4543 870
rect 4543 838 4547 870
rect 4507 802 4547 838
rect 4507 770 4511 802
rect 4511 770 4543 802
rect 4543 770 4547 802
rect 4507 734 4547 770
rect 4507 702 4511 734
rect 4511 702 4543 734
rect 4543 702 4547 734
rect 4507 666 4547 702
rect 4507 634 4511 666
rect 4511 634 4543 666
rect 4543 634 4547 666
rect 4507 598 4547 634
rect 4507 566 4511 598
rect 4511 566 4543 598
rect 4543 566 4547 598
rect 4507 560 4547 566
rect 5715 4318 5755 4324
rect 5715 4286 5719 4318
rect 5719 4286 5751 4318
rect 5751 4286 5755 4318
rect 5715 4250 5755 4286
rect 5715 4218 5719 4250
rect 5719 4218 5751 4250
rect 5751 4218 5755 4250
rect 5715 4182 5755 4218
rect 5715 4150 5719 4182
rect 5719 4150 5751 4182
rect 5751 4150 5755 4182
rect 5715 4114 5755 4150
rect 5715 4082 5719 4114
rect 5719 4082 5751 4114
rect 5751 4082 5755 4114
rect 5715 4046 5755 4082
rect 5715 4014 5719 4046
rect 5719 4014 5751 4046
rect 5751 4014 5755 4046
rect 5715 3978 5755 4014
rect 5715 3946 5719 3978
rect 5719 3946 5751 3978
rect 5751 3946 5755 3978
rect 5715 3910 5755 3946
rect 5715 3878 5719 3910
rect 5719 3878 5751 3910
rect 5751 3878 5755 3910
rect 5715 3842 5755 3878
rect 5715 3810 5719 3842
rect 5719 3810 5751 3842
rect 5751 3810 5755 3842
rect 5715 3774 5755 3810
rect 5715 3742 5719 3774
rect 5719 3742 5751 3774
rect 5751 3742 5755 3774
rect 5715 3706 5755 3742
rect 5715 3674 5719 3706
rect 5719 3674 5751 3706
rect 5751 3674 5755 3706
rect 5715 3638 5755 3674
rect 5715 3606 5719 3638
rect 5719 3606 5751 3638
rect 5751 3606 5755 3638
rect 5715 3570 5755 3606
rect 5715 3538 5719 3570
rect 5719 3538 5751 3570
rect 5751 3538 5755 3570
rect 5715 3502 5755 3538
rect 5715 3470 5719 3502
rect 5719 3470 5751 3502
rect 5751 3470 5755 3502
rect 5715 3464 5755 3470
rect 5372 3350 5494 3356
rect 5372 3318 5417 3350
rect 5417 3318 5449 3350
rect 5449 3318 5494 3350
rect 5372 3282 5494 3318
rect 5372 3250 5417 3282
rect 5417 3250 5449 3282
rect 5449 3250 5494 3282
rect 5372 3214 5494 3250
rect 5372 3182 5417 3214
rect 5417 3182 5449 3214
rect 5449 3182 5494 3214
rect 5372 3146 5494 3182
rect 5372 3114 5417 3146
rect 5417 3114 5449 3146
rect 5449 3114 5494 3146
rect 5372 3078 5494 3114
rect 5372 3046 5417 3078
rect 5417 3046 5449 3078
rect 5449 3046 5494 3078
rect 5372 3010 5494 3046
rect 5372 2978 5417 3010
rect 5417 2978 5449 3010
rect 5449 2978 5494 3010
rect 5372 2942 5494 2978
rect 5372 2910 5417 2942
rect 5417 2910 5449 2942
rect 5449 2910 5494 2942
rect 5372 2874 5494 2910
rect 5372 2842 5417 2874
rect 5417 2842 5449 2874
rect 5449 2842 5494 2874
rect 5372 2806 5494 2842
rect 5372 2774 5417 2806
rect 5417 2774 5449 2806
rect 5449 2774 5494 2806
rect 5372 2738 5494 2774
rect 5372 2706 5417 2738
rect 5417 2706 5449 2738
rect 5449 2706 5494 2738
rect 5372 2670 5494 2706
rect 5372 2638 5417 2670
rect 5417 2638 5449 2670
rect 5449 2638 5494 2670
rect 5372 2602 5494 2638
rect 5372 2570 5417 2602
rect 5417 2570 5449 2602
rect 5449 2570 5494 2602
rect 5372 2534 5494 2570
rect 5372 2502 5417 2534
rect 5417 2502 5449 2534
rect 5449 2502 5494 2534
rect 5372 2496 5494 2502
rect 5111 2382 5151 2388
rect 5111 2350 5115 2382
rect 5115 2350 5147 2382
rect 5147 2350 5151 2382
rect 5111 2314 5151 2350
rect 5111 2282 5115 2314
rect 5115 2282 5147 2314
rect 5147 2282 5151 2314
rect 5111 2246 5151 2282
rect 5111 2214 5115 2246
rect 5115 2214 5147 2246
rect 5147 2214 5151 2246
rect 5111 2178 5151 2214
rect 5111 2146 5115 2178
rect 5115 2146 5147 2178
rect 5147 2146 5151 2178
rect 5111 2110 5151 2146
rect 5111 2078 5115 2110
rect 5115 2078 5147 2110
rect 5147 2078 5151 2110
rect 5111 2042 5151 2078
rect 5111 2010 5115 2042
rect 5115 2010 5147 2042
rect 5147 2010 5151 2042
rect 5111 1974 5151 2010
rect 5111 1942 5115 1974
rect 5115 1942 5147 1974
rect 5147 1942 5151 1974
rect 5111 1906 5151 1942
rect 5111 1874 5115 1906
rect 5115 1874 5147 1906
rect 5147 1874 5151 1906
rect 5111 1838 5151 1874
rect 5111 1806 5115 1838
rect 5115 1806 5147 1838
rect 5147 1806 5151 1838
rect 5111 1770 5151 1806
rect 5111 1738 5115 1770
rect 5115 1738 5147 1770
rect 5147 1738 5151 1770
rect 5111 1702 5151 1738
rect 5111 1670 5115 1702
rect 5115 1670 5147 1702
rect 5147 1670 5151 1702
rect 5111 1634 5151 1670
rect 5111 1602 5115 1634
rect 5115 1602 5147 1634
rect 5147 1602 5151 1634
rect 5111 1566 5151 1602
rect 5111 1534 5115 1566
rect 5115 1534 5147 1566
rect 5147 1534 5151 1566
rect 5111 1528 5151 1534
rect 4768 1414 4890 1420
rect 4768 1382 4813 1414
rect 4813 1382 4845 1414
rect 4845 1382 4890 1414
rect 4768 1346 4890 1382
rect 4768 1314 4813 1346
rect 4813 1314 4845 1346
rect 4845 1314 4890 1346
rect 4768 1278 4890 1314
rect 4768 1246 4813 1278
rect 4813 1246 4845 1278
rect 4845 1246 4890 1278
rect 4768 1210 4890 1246
rect 4768 1178 4813 1210
rect 4813 1178 4845 1210
rect 4845 1178 4890 1210
rect 4768 1142 4890 1178
rect 4768 1110 4813 1142
rect 4813 1110 4845 1142
rect 4845 1110 4890 1142
rect 4768 1074 4890 1110
rect 4768 1042 4813 1074
rect 4813 1042 4845 1074
rect 4845 1042 4890 1074
rect 4768 1006 4890 1042
rect 4768 974 4813 1006
rect 4813 974 4845 1006
rect 4845 974 4890 1006
rect 4768 938 4890 974
rect 4768 906 4813 938
rect 4813 906 4845 938
rect 4845 906 4890 938
rect 4768 870 4890 906
rect 4768 838 4813 870
rect 4813 838 4845 870
rect 4845 838 4890 870
rect 4768 802 4890 838
rect 4768 770 4813 802
rect 4813 770 4845 802
rect 4845 770 4890 802
rect 4768 734 4890 770
rect 4768 702 4813 734
rect 4813 702 4845 734
rect 4845 702 4890 734
rect 4768 666 4890 702
rect 4768 634 4813 666
rect 4813 634 4845 666
rect 4845 634 4890 666
rect 4768 598 4890 634
rect 4768 566 4813 598
rect 4813 566 4845 598
rect 4845 566 4890 598
rect 4768 560 4890 566
rect 5976 4318 6098 4324
rect 5976 4286 6021 4318
rect 6021 4286 6053 4318
rect 6053 4286 6098 4318
rect 5976 4250 6098 4286
rect 5976 4218 6021 4250
rect 6021 4218 6053 4250
rect 6053 4218 6098 4250
rect 5976 4182 6098 4218
rect 5976 4150 6021 4182
rect 6021 4150 6053 4182
rect 6053 4150 6098 4182
rect 5976 4114 6098 4150
rect 5976 4082 6021 4114
rect 6021 4082 6053 4114
rect 6053 4082 6098 4114
rect 5976 4046 6098 4082
rect 5976 4014 6021 4046
rect 6021 4014 6053 4046
rect 6053 4014 6098 4046
rect 5976 3978 6098 4014
rect 5976 3946 6021 3978
rect 6021 3946 6053 3978
rect 6053 3946 6098 3978
rect 5976 3910 6098 3946
rect 5976 3878 6021 3910
rect 6021 3878 6053 3910
rect 6053 3878 6098 3910
rect 5976 3842 6098 3878
rect 5976 3810 6021 3842
rect 6021 3810 6053 3842
rect 6053 3810 6098 3842
rect 5976 3774 6098 3810
rect 5976 3742 6021 3774
rect 6021 3742 6053 3774
rect 6053 3742 6098 3774
rect 5976 3706 6098 3742
rect 5976 3674 6021 3706
rect 6021 3674 6053 3706
rect 6053 3674 6098 3706
rect 5976 3638 6098 3674
rect 5976 3606 6021 3638
rect 6021 3606 6053 3638
rect 6053 3606 6098 3638
rect 5976 3570 6098 3606
rect 5976 3538 6021 3570
rect 6021 3538 6053 3570
rect 6053 3538 6098 3570
rect 5976 3502 6098 3538
rect 5976 3470 6021 3502
rect 6021 3470 6053 3502
rect 6053 3470 6098 3502
rect 5976 3464 6098 3470
rect 5715 3350 5755 3356
rect 5715 3318 5719 3350
rect 5719 3318 5751 3350
rect 5751 3318 5755 3350
rect 5715 3282 5755 3318
rect 5715 3250 5719 3282
rect 5719 3250 5751 3282
rect 5751 3250 5755 3282
rect 5715 3214 5755 3250
rect 5715 3182 5719 3214
rect 5719 3182 5751 3214
rect 5751 3182 5755 3214
rect 5715 3146 5755 3182
rect 5715 3114 5719 3146
rect 5719 3114 5751 3146
rect 5751 3114 5755 3146
rect 5715 3078 5755 3114
rect 5715 3046 5719 3078
rect 5719 3046 5751 3078
rect 5751 3046 5755 3078
rect 5715 3010 5755 3046
rect 5715 2978 5719 3010
rect 5719 2978 5751 3010
rect 5751 2978 5755 3010
rect 5715 2942 5755 2978
rect 5715 2910 5719 2942
rect 5719 2910 5751 2942
rect 5751 2910 5755 2942
rect 5715 2874 5755 2910
rect 5715 2842 5719 2874
rect 5719 2842 5751 2874
rect 5751 2842 5755 2874
rect 5715 2806 5755 2842
rect 5715 2774 5719 2806
rect 5719 2774 5751 2806
rect 5751 2774 5755 2806
rect 5715 2738 5755 2774
rect 5715 2706 5719 2738
rect 5719 2706 5751 2738
rect 5751 2706 5755 2738
rect 5715 2670 5755 2706
rect 5715 2638 5719 2670
rect 5719 2638 5751 2670
rect 5751 2638 5755 2670
rect 5715 2602 5755 2638
rect 5715 2570 5719 2602
rect 5719 2570 5751 2602
rect 5751 2570 5755 2602
rect 5715 2534 5755 2570
rect 5715 2502 5719 2534
rect 5719 2502 5751 2534
rect 5751 2502 5755 2534
rect 5715 2496 5755 2502
rect 5372 2382 5494 2388
rect 5372 2350 5417 2382
rect 5417 2350 5449 2382
rect 5449 2350 5494 2382
rect 5372 2314 5494 2350
rect 5372 2282 5417 2314
rect 5417 2282 5449 2314
rect 5449 2282 5494 2314
rect 5372 2246 5494 2282
rect 5372 2214 5417 2246
rect 5417 2214 5449 2246
rect 5449 2214 5494 2246
rect 5372 2178 5494 2214
rect 5372 2146 5417 2178
rect 5417 2146 5449 2178
rect 5449 2146 5494 2178
rect 5372 2110 5494 2146
rect 5372 2078 5417 2110
rect 5417 2078 5449 2110
rect 5449 2078 5494 2110
rect 5372 2042 5494 2078
rect 5372 2010 5417 2042
rect 5417 2010 5449 2042
rect 5449 2010 5494 2042
rect 5372 1974 5494 2010
rect 5372 1942 5417 1974
rect 5417 1942 5449 1974
rect 5449 1942 5494 1974
rect 5372 1906 5494 1942
rect 5372 1874 5417 1906
rect 5417 1874 5449 1906
rect 5449 1874 5494 1906
rect 5372 1838 5494 1874
rect 5372 1806 5417 1838
rect 5417 1806 5449 1838
rect 5449 1806 5494 1838
rect 5372 1770 5494 1806
rect 5372 1738 5417 1770
rect 5417 1738 5449 1770
rect 5449 1738 5494 1770
rect 5372 1702 5494 1738
rect 5372 1670 5417 1702
rect 5417 1670 5449 1702
rect 5449 1670 5494 1702
rect 5372 1634 5494 1670
rect 5372 1602 5417 1634
rect 5417 1602 5449 1634
rect 5449 1602 5494 1634
rect 5372 1566 5494 1602
rect 5372 1534 5417 1566
rect 5417 1534 5449 1566
rect 5449 1534 5494 1566
rect 5372 1528 5494 1534
rect 5111 1414 5151 1420
rect 5111 1382 5115 1414
rect 5115 1382 5147 1414
rect 5147 1382 5151 1414
rect 5111 1346 5151 1382
rect 5111 1314 5115 1346
rect 5115 1314 5147 1346
rect 5147 1314 5151 1346
rect 5111 1278 5151 1314
rect 5111 1246 5115 1278
rect 5115 1246 5147 1278
rect 5147 1246 5151 1278
rect 5111 1210 5151 1246
rect 5111 1178 5115 1210
rect 5115 1178 5147 1210
rect 5147 1178 5151 1210
rect 5111 1142 5151 1178
rect 5111 1110 5115 1142
rect 5115 1110 5147 1142
rect 5147 1110 5151 1142
rect 5111 1074 5151 1110
rect 5111 1042 5115 1074
rect 5115 1042 5147 1074
rect 5147 1042 5151 1074
rect 5111 1006 5151 1042
rect 5111 974 5115 1006
rect 5115 974 5147 1006
rect 5147 974 5151 1006
rect 5111 938 5151 974
rect 5111 906 5115 938
rect 5115 906 5147 938
rect 5147 906 5151 938
rect 5111 870 5151 906
rect 5111 838 5115 870
rect 5115 838 5147 870
rect 5147 838 5151 870
rect 5111 802 5151 838
rect 5111 770 5115 802
rect 5115 770 5147 802
rect 5147 770 5151 802
rect 5111 734 5151 770
rect 5111 702 5115 734
rect 5115 702 5147 734
rect 5147 702 5151 734
rect 5111 666 5151 702
rect 5111 634 5115 666
rect 5115 634 5147 666
rect 5147 634 5151 666
rect 5111 598 5151 634
rect 5111 566 5115 598
rect 5115 566 5147 598
rect 5147 566 5151 598
rect 5111 560 5151 566
rect 6319 4318 6359 4324
rect 6319 4286 6323 4318
rect 6323 4286 6355 4318
rect 6355 4286 6359 4318
rect 6319 4250 6359 4286
rect 6319 4218 6323 4250
rect 6323 4218 6355 4250
rect 6355 4218 6359 4250
rect 6319 4182 6359 4218
rect 6319 4150 6323 4182
rect 6323 4150 6355 4182
rect 6355 4150 6359 4182
rect 6319 4114 6359 4150
rect 6319 4082 6323 4114
rect 6323 4082 6355 4114
rect 6355 4082 6359 4114
rect 6319 4046 6359 4082
rect 6319 4014 6323 4046
rect 6323 4014 6355 4046
rect 6355 4014 6359 4046
rect 6319 3978 6359 4014
rect 6319 3946 6323 3978
rect 6323 3946 6355 3978
rect 6355 3946 6359 3978
rect 6319 3910 6359 3946
rect 6319 3878 6323 3910
rect 6323 3878 6355 3910
rect 6355 3878 6359 3910
rect 6319 3842 6359 3878
rect 6319 3810 6323 3842
rect 6323 3810 6355 3842
rect 6355 3810 6359 3842
rect 6319 3774 6359 3810
rect 6319 3742 6323 3774
rect 6323 3742 6355 3774
rect 6355 3742 6359 3774
rect 6319 3706 6359 3742
rect 6319 3674 6323 3706
rect 6323 3674 6355 3706
rect 6355 3674 6359 3706
rect 6319 3638 6359 3674
rect 6319 3606 6323 3638
rect 6323 3606 6355 3638
rect 6355 3606 6359 3638
rect 6319 3570 6359 3606
rect 6319 3538 6323 3570
rect 6323 3538 6355 3570
rect 6355 3538 6359 3570
rect 6319 3502 6359 3538
rect 6319 3470 6323 3502
rect 6323 3470 6355 3502
rect 6355 3470 6359 3502
rect 6319 3464 6359 3470
rect 5976 3350 6098 3356
rect 5976 3318 6021 3350
rect 6021 3318 6053 3350
rect 6053 3318 6098 3350
rect 5976 3282 6098 3318
rect 5976 3250 6021 3282
rect 6021 3250 6053 3282
rect 6053 3250 6098 3282
rect 5976 3214 6098 3250
rect 5976 3182 6021 3214
rect 6021 3182 6053 3214
rect 6053 3182 6098 3214
rect 5976 3146 6098 3182
rect 5976 3114 6021 3146
rect 6021 3114 6053 3146
rect 6053 3114 6098 3146
rect 5976 3078 6098 3114
rect 5976 3046 6021 3078
rect 6021 3046 6053 3078
rect 6053 3046 6098 3078
rect 5976 3010 6098 3046
rect 5976 2978 6021 3010
rect 6021 2978 6053 3010
rect 6053 2978 6098 3010
rect 5976 2942 6098 2978
rect 5976 2910 6021 2942
rect 6021 2910 6053 2942
rect 6053 2910 6098 2942
rect 5976 2874 6098 2910
rect 5976 2842 6021 2874
rect 6021 2842 6053 2874
rect 6053 2842 6098 2874
rect 5976 2806 6098 2842
rect 5976 2774 6021 2806
rect 6021 2774 6053 2806
rect 6053 2774 6098 2806
rect 5976 2738 6098 2774
rect 5976 2706 6021 2738
rect 6021 2706 6053 2738
rect 6053 2706 6098 2738
rect 5976 2670 6098 2706
rect 5976 2638 6021 2670
rect 6021 2638 6053 2670
rect 6053 2638 6098 2670
rect 5976 2602 6098 2638
rect 5976 2570 6021 2602
rect 6021 2570 6053 2602
rect 6053 2570 6098 2602
rect 5976 2534 6098 2570
rect 5976 2502 6021 2534
rect 6021 2502 6053 2534
rect 6053 2502 6098 2534
rect 5976 2496 6098 2502
rect 5715 2382 5755 2388
rect 5715 2350 5719 2382
rect 5719 2350 5751 2382
rect 5751 2350 5755 2382
rect 5715 2314 5755 2350
rect 5715 2282 5719 2314
rect 5719 2282 5751 2314
rect 5751 2282 5755 2314
rect 5715 2246 5755 2282
rect 5715 2214 5719 2246
rect 5719 2214 5751 2246
rect 5751 2214 5755 2246
rect 5715 2178 5755 2214
rect 5715 2146 5719 2178
rect 5719 2146 5751 2178
rect 5751 2146 5755 2178
rect 5715 2110 5755 2146
rect 5715 2078 5719 2110
rect 5719 2078 5751 2110
rect 5751 2078 5755 2110
rect 5715 2042 5755 2078
rect 5715 2010 5719 2042
rect 5719 2010 5751 2042
rect 5751 2010 5755 2042
rect 5715 1974 5755 2010
rect 5715 1942 5719 1974
rect 5719 1942 5751 1974
rect 5751 1942 5755 1974
rect 5715 1906 5755 1942
rect 5715 1874 5719 1906
rect 5719 1874 5751 1906
rect 5751 1874 5755 1906
rect 5715 1838 5755 1874
rect 5715 1806 5719 1838
rect 5719 1806 5751 1838
rect 5751 1806 5755 1838
rect 5715 1770 5755 1806
rect 5715 1738 5719 1770
rect 5719 1738 5751 1770
rect 5751 1738 5755 1770
rect 5715 1702 5755 1738
rect 5715 1670 5719 1702
rect 5719 1670 5751 1702
rect 5751 1670 5755 1702
rect 5715 1634 5755 1670
rect 5715 1602 5719 1634
rect 5719 1602 5751 1634
rect 5751 1602 5755 1634
rect 5715 1566 5755 1602
rect 5715 1534 5719 1566
rect 5719 1534 5751 1566
rect 5751 1534 5755 1566
rect 5715 1528 5755 1534
rect 5372 1414 5494 1420
rect 5372 1382 5417 1414
rect 5417 1382 5449 1414
rect 5449 1382 5494 1414
rect 5372 1346 5494 1382
rect 5372 1314 5417 1346
rect 5417 1314 5449 1346
rect 5449 1314 5494 1346
rect 5372 1278 5494 1314
rect 5372 1246 5417 1278
rect 5417 1246 5449 1278
rect 5449 1246 5494 1278
rect 5372 1210 5494 1246
rect 5372 1178 5417 1210
rect 5417 1178 5449 1210
rect 5449 1178 5494 1210
rect 5372 1142 5494 1178
rect 5372 1110 5417 1142
rect 5417 1110 5449 1142
rect 5449 1110 5494 1142
rect 5372 1074 5494 1110
rect 5372 1042 5417 1074
rect 5417 1042 5449 1074
rect 5449 1042 5494 1074
rect 5372 1006 5494 1042
rect 5372 974 5417 1006
rect 5417 974 5449 1006
rect 5449 974 5494 1006
rect 5372 938 5494 974
rect 5372 906 5417 938
rect 5417 906 5449 938
rect 5449 906 5494 938
rect 5372 870 5494 906
rect 5372 838 5417 870
rect 5417 838 5449 870
rect 5449 838 5494 870
rect 5372 802 5494 838
rect 5372 770 5417 802
rect 5417 770 5449 802
rect 5449 770 5494 802
rect 5372 734 5494 770
rect 5372 702 5417 734
rect 5417 702 5449 734
rect 5449 702 5494 734
rect 5372 666 5494 702
rect 5372 634 5417 666
rect 5417 634 5449 666
rect 5449 634 5494 666
rect 5372 598 5494 634
rect 5372 566 5417 598
rect 5417 566 5449 598
rect 5449 566 5494 598
rect 5372 560 5494 566
rect 6580 4318 6702 4324
rect 6580 4286 6625 4318
rect 6625 4286 6657 4318
rect 6657 4286 6702 4318
rect 6580 4250 6702 4286
rect 6580 4218 6625 4250
rect 6625 4218 6657 4250
rect 6657 4218 6702 4250
rect 6580 4182 6702 4218
rect 6580 4150 6625 4182
rect 6625 4150 6657 4182
rect 6657 4150 6702 4182
rect 6580 4114 6702 4150
rect 6580 4082 6625 4114
rect 6625 4082 6657 4114
rect 6657 4082 6702 4114
rect 6580 4046 6702 4082
rect 6580 4014 6625 4046
rect 6625 4014 6657 4046
rect 6657 4014 6702 4046
rect 6580 3978 6702 4014
rect 6580 3946 6625 3978
rect 6625 3946 6657 3978
rect 6657 3946 6702 3978
rect 6580 3910 6702 3946
rect 6580 3878 6625 3910
rect 6625 3878 6657 3910
rect 6657 3878 6702 3910
rect 6580 3842 6702 3878
rect 6580 3810 6625 3842
rect 6625 3810 6657 3842
rect 6657 3810 6702 3842
rect 6580 3774 6702 3810
rect 6580 3742 6625 3774
rect 6625 3742 6657 3774
rect 6657 3742 6702 3774
rect 6580 3706 6702 3742
rect 6580 3674 6625 3706
rect 6625 3674 6657 3706
rect 6657 3674 6702 3706
rect 6580 3638 6702 3674
rect 6580 3606 6625 3638
rect 6625 3606 6657 3638
rect 6657 3606 6702 3638
rect 6580 3570 6702 3606
rect 6580 3538 6625 3570
rect 6625 3538 6657 3570
rect 6657 3538 6702 3570
rect 6580 3502 6702 3538
rect 6580 3470 6625 3502
rect 6625 3470 6657 3502
rect 6657 3470 6702 3502
rect 6580 3464 6702 3470
rect 6319 3350 6359 3356
rect 6319 3318 6323 3350
rect 6323 3318 6355 3350
rect 6355 3318 6359 3350
rect 6319 3282 6359 3318
rect 6319 3250 6323 3282
rect 6323 3250 6355 3282
rect 6355 3250 6359 3282
rect 6319 3214 6359 3250
rect 6319 3182 6323 3214
rect 6323 3182 6355 3214
rect 6355 3182 6359 3214
rect 6319 3146 6359 3182
rect 6319 3114 6323 3146
rect 6323 3114 6355 3146
rect 6355 3114 6359 3146
rect 6319 3078 6359 3114
rect 6319 3046 6323 3078
rect 6323 3046 6355 3078
rect 6355 3046 6359 3078
rect 6319 3010 6359 3046
rect 6319 2978 6323 3010
rect 6323 2978 6355 3010
rect 6355 2978 6359 3010
rect 6319 2942 6359 2978
rect 6319 2910 6323 2942
rect 6323 2910 6355 2942
rect 6355 2910 6359 2942
rect 6319 2874 6359 2910
rect 6319 2842 6323 2874
rect 6323 2842 6355 2874
rect 6355 2842 6359 2874
rect 6319 2806 6359 2842
rect 6319 2774 6323 2806
rect 6323 2774 6355 2806
rect 6355 2774 6359 2806
rect 6319 2738 6359 2774
rect 6319 2706 6323 2738
rect 6323 2706 6355 2738
rect 6355 2706 6359 2738
rect 6319 2670 6359 2706
rect 6319 2638 6323 2670
rect 6323 2638 6355 2670
rect 6355 2638 6359 2670
rect 6319 2602 6359 2638
rect 6319 2570 6323 2602
rect 6323 2570 6355 2602
rect 6355 2570 6359 2602
rect 6319 2534 6359 2570
rect 6319 2502 6323 2534
rect 6323 2502 6355 2534
rect 6355 2502 6359 2534
rect 6319 2496 6359 2502
rect 5976 2382 6098 2388
rect 5976 2350 6021 2382
rect 6021 2350 6053 2382
rect 6053 2350 6098 2382
rect 5976 2314 6098 2350
rect 5976 2282 6021 2314
rect 6021 2282 6053 2314
rect 6053 2282 6098 2314
rect 5976 2246 6098 2282
rect 5976 2214 6021 2246
rect 6021 2214 6053 2246
rect 6053 2214 6098 2246
rect 5976 2178 6098 2214
rect 5976 2146 6021 2178
rect 6021 2146 6053 2178
rect 6053 2146 6098 2178
rect 5976 2110 6098 2146
rect 5976 2078 6021 2110
rect 6021 2078 6053 2110
rect 6053 2078 6098 2110
rect 5976 2042 6098 2078
rect 5976 2010 6021 2042
rect 6021 2010 6053 2042
rect 6053 2010 6098 2042
rect 5976 1974 6098 2010
rect 5976 1942 6021 1974
rect 6021 1942 6053 1974
rect 6053 1942 6098 1974
rect 5976 1906 6098 1942
rect 5976 1874 6021 1906
rect 6021 1874 6053 1906
rect 6053 1874 6098 1906
rect 5976 1838 6098 1874
rect 5976 1806 6021 1838
rect 6021 1806 6053 1838
rect 6053 1806 6098 1838
rect 5976 1770 6098 1806
rect 5976 1738 6021 1770
rect 6021 1738 6053 1770
rect 6053 1738 6098 1770
rect 5976 1702 6098 1738
rect 5976 1670 6021 1702
rect 6021 1670 6053 1702
rect 6053 1670 6098 1702
rect 5976 1634 6098 1670
rect 5976 1602 6021 1634
rect 6021 1602 6053 1634
rect 6053 1602 6098 1634
rect 5976 1566 6098 1602
rect 5976 1534 6021 1566
rect 6021 1534 6053 1566
rect 6053 1534 6098 1566
rect 5976 1528 6098 1534
rect 5715 1414 5755 1420
rect 5715 1382 5719 1414
rect 5719 1382 5751 1414
rect 5751 1382 5755 1414
rect 5715 1346 5755 1382
rect 5715 1314 5719 1346
rect 5719 1314 5751 1346
rect 5751 1314 5755 1346
rect 5715 1278 5755 1314
rect 5715 1246 5719 1278
rect 5719 1246 5751 1278
rect 5751 1246 5755 1278
rect 5715 1210 5755 1246
rect 5715 1178 5719 1210
rect 5719 1178 5751 1210
rect 5751 1178 5755 1210
rect 5715 1142 5755 1178
rect 5715 1110 5719 1142
rect 5719 1110 5751 1142
rect 5751 1110 5755 1142
rect 5715 1074 5755 1110
rect 5715 1042 5719 1074
rect 5719 1042 5751 1074
rect 5751 1042 5755 1074
rect 5715 1006 5755 1042
rect 5715 974 5719 1006
rect 5719 974 5751 1006
rect 5751 974 5755 1006
rect 5715 938 5755 974
rect 5715 906 5719 938
rect 5719 906 5751 938
rect 5751 906 5755 938
rect 5715 870 5755 906
rect 5715 838 5719 870
rect 5719 838 5751 870
rect 5751 838 5755 870
rect 5715 802 5755 838
rect 5715 770 5719 802
rect 5719 770 5751 802
rect 5751 770 5755 802
rect 5715 734 5755 770
rect 5715 702 5719 734
rect 5719 702 5751 734
rect 5751 702 5755 734
rect 5715 666 5755 702
rect 5715 634 5719 666
rect 5719 634 5751 666
rect 5751 634 5755 666
rect 5715 598 5755 634
rect 5715 566 5719 598
rect 5719 566 5751 598
rect 5751 566 5755 598
rect 5715 560 5755 566
rect 6923 4318 6963 4324
rect 6923 4286 6927 4318
rect 6927 4286 6959 4318
rect 6959 4286 6963 4318
rect 6923 4250 6963 4286
rect 6923 4218 6927 4250
rect 6927 4218 6959 4250
rect 6959 4218 6963 4250
rect 6923 4182 6963 4218
rect 6923 4150 6927 4182
rect 6927 4150 6959 4182
rect 6959 4150 6963 4182
rect 6923 4114 6963 4150
rect 6923 4082 6927 4114
rect 6927 4082 6959 4114
rect 6959 4082 6963 4114
rect 6923 4046 6963 4082
rect 6923 4014 6927 4046
rect 6927 4014 6959 4046
rect 6959 4014 6963 4046
rect 6923 3978 6963 4014
rect 6923 3946 6927 3978
rect 6927 3946 6959 3978
rect 6959 3946 6963 3978
rect 6923 3910 6963 3946
rect 6923 3878 6927 3910
rect 6927 3878 6959 3910
rect 6959 3878 6963 3910
rect 6923 3842 6963 3878
rect 6923 3810 6927 3842
rect 6927 3810 6959 3842
rect 6959 3810 6963 3842
rect 6923 3774 6963 3810
rect 6923 3742 6927 3774
rect 6927 3742 6959 3774
rect 6959 3742 6963 3774
rect 6923 3706 6963 3742
rect 6923 3674 6927 3706
rect 6927 3674 6959 3706
rect 6959 3674 6963 3706
rect 6923 3638 6963 3674
rect 6923 3606 6927 3638
rect 6927 3606 6959 3638
rect 6959 3606 6963 3638
rect 6923 3570 6963 3606
rect 6923 3538 6927 3570
rect 6927 3538 6959 3570
rect 6959 3538 6963 3570
rect 6923 3502 6963 3538
rect 6923 3470 6927 3502
rect 6927 3470 6959 3502
rect 6959 3470 6963 3502
rect 6923 3464 6963 3470
rect 6580 3350 6702 3356
rect 6580 3318 6625 3350
rect 6625 3318 6657 3350
rect 6657 3318 6702 3350
rect 6580 3282 6702 3318
rect 6580 3250 6625 3282
rect 6625 3250 6657 3282
rect 6657 3250 6702 3282
rect 6580 3214 6702 3250
rect 6580 3182 6625 3214
rect 6625 3182 6657 3214
rect 6657 3182 6702 3214
rect 6580 3146 6702 3182
rect 6580 3114 6625 3146
rect 6625 3114 6657 3146
rect 6657 3114 6702 3146
rect 6580 3078 6702 3114
rect 6580 3046 6625 3078
rect 6625 3046 6657 3078
rect 6657 3046 6702 3078
rect 6580 3010 6702 3046
rect 6580 2978 6625 3010
rect 6625 2978 6657 3010
rect 6657 2978 6702 3010
rect 6580 2942 6702 2978
rect 6580 2910 6625 2942
rect 6625 2910 6657 2942
rect 6657 2910 6702 2942
rect 6580 2874 6702 2910
rect 6580 2842 6625 2874
rect 6625 2842 6657 2874
rect 6657 2842 6702 2874
rect 6580 2806 6702 2842
rect 6580 2774 6625 2806
rect 6625 2774 6657 2806
rect 6657 2774 6702 2806
rect 6580 2738 6702 2774
rect 6580 2706 6625 2738
rect 6625 2706 6657 2738
rect 6657 2706 6702 2738
rect 6580 2670 6702 2706
rect 6580 2638 6625 2670
rect 6625 2638 6657 2670
rect 6657 2638 6702 2670
rect 6580 2602 6702 2638
rect 6580 2570 6625 2602
rect 6625 2570 6657 2602
rect 6657 2570 6702 2602
rect 6580 2534 6702 2570
rect 6580 2502 6625 2534
rect 6625 2502 6657 2534
rect 6657 2502 6702 2534
rect 6580 2496 6702 2502
rect 6319 2382 6359 2388
rect 6319 2350 6323 2382
rect 6323 2350 6355 2382
rect 6355 2350 6359 2382
rect 6319 2314 6359 2350
rect 6319 2282 6323 2314
rect 6323 2282 6355 2314
rect 6355 2282 6359 2314
rect 6319 2246 6359 2282
rect 6319 2214 6323 2246
rect 6323 2214 6355 2246
rect 6355 2214 6359 2246
rect 6319 2178 6359 2214
rect 6319 2146 6323 2178
rect 6323 2146 6355 2178
rect 6355 2146 6359 2178
rect 6319 2110 6359 2146
rect 6319 2078 6323 2110
rect 6323 2078 6355 2110
rect 6355 2078 6359 2110
rect 6319 2042 6359 2078
rect 6319 2010 6323 2042
rect 6323 2010 6355 2042
rect 6355 2010 6359 2042
rect 6319 1974 6359 2010
rect 6319 1942 6323 1974
rect 6323 1942 6355 1974
rect 6355 1942 6359 1974
rect 6319 1906 6359 1942
rect 6319 1874 6323 1906
rect 6323 1874 6355 1906
rect 6355 1874 6359 1906
rect 6319 1838 6359 1874
rect 6319 1806 6323 1838
rect 6323 1806 6355 1838
rect 6355 1806 6359 1838
rect 6319 1770 6359 1806
rect 6319 1738 6323 1770
rect 6323 1738 6355 1770
rect 6355 1738 6359 1770
rect 6319 1702 6359 1738
rect 6319 1670 6323 1702
rect 6323 1670 6355 1702
rect 6355 1670 6359 1702
rect 6319 1634 6359 1670
rect 6319 1602 6323 1634
rect 6323 1602 6355 1634
rect 6355 1602 6359 1634
rect 6319 1566 6359 1602
rect 6319 1534 6323 1566
rect 6323 1534 6355 1566
rect 6355 1534 6359 1566
rect 6319 1528 6359 1534
rect 5976 1414 6098 1420
rect 5976 1382 6021 1414
rect 6021 1382 6053 1414
rect 6053 1382 6098 1414
rect 5976 1346 6098 1382
rect 5976 1314 6021 1346
rect 6021 1314 6053 1346
rect 6053 1314 6098 1346
rect 5976 1278 6098 1314
rect 5976 1246 6021 1278
rect 6021 1246 6053 1278
rect 6053 1246 6098 1278
rect 5976 1210 6098 1246
rect 5976 1178 6021 1210
rect 6021 1178 6053 1210
rect 6053 1178 6098 1210
rect 5976 1142 6098 1178
rect 5976 1110 6021 1142
rect 6021 1110 6053 1142
rect 6053 1110 6098 1142
rect 5976 1074 6098 1110
rect 5976 1042 6021 1074
rect 6021 1042 6053 1074
rect 6053 1042 6098 1074
rect 5976 1006 6098 1042
rect 5976 974 6021 1006
rect 6021 974 6053 1006
rect 6053 974 6098 1006
rect 5976 938 6098 974
rect 5976 906 6021 938
rect 6021 906 6053 938
rect 6053 906 6098 938
rect 5976 870 6098 906
rect 5976 838 6021 870
rect 6021 838 6053 870
rect 6053 838 6098 870
rect 5976 802 6098 838
rect 5976 770 6021 802
rect 6021 770 6053 802
rect 6053 770 6098 802
rect 5976 734 6098 770
rect 5976 702 6021 734
rect 6021 702 6053 734
rect 6053 702 6098 734
rect 5976 666 6098 702
rect 5976 634 6021 666
rect 6021 634 6053 666
rect 6053 634 6098 666
rect 5976 598 6098 634
rect 5976 566 6021 598
rect 6021 566 6053 598
rect 6053 566 6098 598
rect 5976 560 6098 566
rect 7184 4318 7306 4324
rect 7184 4286 7229 4318
rect 7229 4286 7261 4318
rect 7261 4286 7306 4318
rect 7184 4250 7306 4286
rect 7184 4218 7229 4250
rect 7229 4218 7261 4250
rect 7261 4218 7306 4250
rect 7184 4182 7306 4218
rect 7184 4150 7229 4182
rect 7229 4150 7261 4182
rect 7261 4150 7306 4182
rect 7184 4114 7306 4150
rect 7184 4082 7229 4114
rect 7229 4082 7261 4114
rect 7261 4082 7306 4114
rect 7184 4046 7306 4082
rect 7184 4014 7229 4046
rect 7229 4014 7261 4046
rect 7261 4014 7306 4046
rect 7184 3978 7306 4014
rect 7184 3946 7229 3978
rect 7229 3946 7261 3978
rect 7261 3946 7306 3978
rect 7184 3910 7306 3946
rect 7184 3878 7229 3910
rect 7229 3878 7261 3910
rect 7261 3878 7306 3910
rect 7184 3842 7306 3878
rect 7184 3810 7229 3842
rect 7229 3810 7261 3842
rect 7261 3810 7306 3842
rect 7184 3774 7306 3810
rect 7184 3742 7229 3774
rect 7229 3742 7261 3774
rect 7261 3742 7306 3774
rect 7184 3706 7306 3742
rect 7184 3674 7229 3706
rect 7229 3674 7261 3706
rect 7261 3674 7306 3706
rect 7184 3638 7306 3674
rect 7184 3606 7229 3638
rect 7229 3606 7261 3638
rect 7261 3606 7306 3638
rect 7184 3570 7306 3606
rect 7184 3538 7229 3570
rect 7229 3538 7261 3570
rect 7261 3538 7306 3570
rect 7184 3502 7306 3538
rect 7184 3470 7229 3502
rect 7229 3470 7261 3502
rect 7261 3470 7306 3502
rect 7184 3464 7306 3470
rect 6923 3350 6963 3356
rect 6923 3318 6927 3350
rect 6927 3318 6959 3350
rect 6959 3318 6963 3350
rect 6923 3282 6963 3318
rect 6923 3250 6927 3282
rect 6927 3250 6959 3282
rect 6959 3250 6963 3282
rect 6923 3214 6963 3250
rect 6923 3182 6927 3214
rect 6927 3182 6959 3214
rect 6959 3182 6963 3214
rect 6923 3146 6963 3182
rect 6923 3114 6927 3146
rect 6927 3114 6959 3146
rect 6959 3114 6963 3146
rect 6923 3078 6963 3114
rect 6923 3046 6927 3078
rect 6927 3046 6959 3078
rect 6959 3046 6963 3078
rect 6923 3010 6963 3046
rect 6923 2978 6927 3010
rect 6927 2978 6959 3010
rect 6959 2978 6963 3010
rect 6923 2942 6963 2978
rect 6923 2910 6927 2942
rect 6927 2910 6959 2942
rect 6959 2910 6963 2942
rect 6923 2874 6963 2910
rect 6923 2842 6927 2874
rect 6927 2842 6959 2874
rect 6959 2842 6963 2874
rect 6923 2806 6963 2842
rect 6923 2774 6927 2806
rect 6927 2774 6959 2806
rect 6959 2774 6963 2806
rect 6923 2738 6963 2774
rect 6923 2706 6927 2738
rect 6927 2706 6959 2738
rect 6959 2706 6963 2738
rect 6923 2670 6963 2706
rect 6923 2638 6927 2670
rect 6927 2638 6959 2670
rect 6959 2638 6963 2670
rect 6923 2602 6963 2638
rect 6923 2570 6927 2602
rect 6927 2570 6959 2602
rect 6959 2570 6963 2602
rect 6923 2534 6963 2570
rect 6923 2502 6927 2534
rect 6927 2502 6959 2534
rect 6959 2502 6963 2534
rect 6923 2496 6963 2502
rect 6580 2382 6702 2388
rect 6580 2350 6625 2382
rect 6625 2350 6657 2382
rect 6657 2350 6702 2382
rect 6580 2314 6702 2350
rect 6580 2282 6625 2314
rect 6625 2282 6657 2314
rect 6657 2282 6702 2314
rect 6580 2246 6702 2282
rect 6580 2214 6625 2246
rect 6625 2214 6657 2246
rect 6657 2214 6702 2246
rect 6580 2178 6702 2214
rect 6580 2146 6625 2178
rect 6625 2146 6657 2178
rect 6657 2146 6702 2178
rect 6580 2110 6702 2146
rect 6580 2078 6625 2110
rect 6625 2078 6657 2110
rect 6657 2078 6702 2110
rect 6580 2042 6702 2078
rect 6580 2010 6625 2042
rect 6625 2010 6657 2042
rect 6657 2010 6702 2042
rect 6580 1974 6702 2010
rect 6580 1942 6625 1974
rect 6625 1942 6657 1974
rect 6657 1942 6702 1974
rect 6580 1906 6702 1942
rect 6580 1874 6625 1906
rect 6625 1874 6657 1906
rect 6657 1874 6702 1906
rect 6580 1838 6702 1874
rect 6580 1806 6625 1838
rect 6625 1806 6657 1838
rect 6657 1806 6702 1838
rect 6580 1770 6702 1806
rect 6580 1738 6625 1770
rect 6625 1738 6657 1770
rect 6657 1738 6702 1770
rect 6580 1702 6702 1738
rect 6580 1670 6625 1702
rect 6625 1670 6657 1702
rect 6657 1670 6702 1702
rect 6580 1634 6702 1670
rect 6580 1602 6625 1634
rect 6625 1602 6657 1634
rect 6657 1602 6702 1634
rect 6580 1566 6702 1602
rect 6580 1534 6625 1566
rect 6625 1534 6657 1566
rect 6657 1534 6702 1566
rect 6580 1528 6702 1534
rect 6319 1414 6359 1420
rect 6319 1382 6323 1414
rect 6323 1382 6355 1414
rect 6355 1382 6359 1414
rect 6319 1346 6359 1382
rect 6319 1314 6323 1346
rect 6323 1314 6355 1346
rect 6355 1314 6359 1346
rect 6319 1278 6359 1314
rect 6319 1246 6323 1278
rect 6323 1246 6355 1278
rect 6355 1246 6359 1278
rect 6319 1210 6359 1246
rect 6319 1178 6323 1210
rect 6323 1178 6355 1210
rect 6355 1178 6359 1210
rect 6319 1142 6359 1178
rect 6319 1110 6323 1142
rect 6323 1110 6355 1142
rect 6355 1110 6359 1142
rect 6319 1074 6359 1110
rect 6319 1042 6323 1074
rect 6323 1042 6355 1074
rect 6355 1042 6359 1074
rect 6319 1006 6359 1042
rect 6319 974 6323 1006
rect 6323 974 6355 1006
rect 6355 974 6359 1006
rect 6319 938 6359 974
rect 6319 906 6323 938
rect 6323 906 6355 938
rect 6355 906 6359 938
rect 6319 870 6359 906
rect 6319 838 6323 870
rect 6323 838 6355 870
rect 6355 838 6359 870
rect 6319 802 6359 838
rect 6319 770 6323 802
rect 6323 770 6355 802
rect 6355 770 6359 802
rect 6319 734 6359 770
rect 6319 702 6323 734
rect 6323 702 6355 734
rect 6355 702 6359 734
rect 6319 666 6359 702
rect 6319 634 6323 666
rect 6323 634 6355 666
rect 6355 634 6359 666
rect 6319 598 6359 634
rect 6319 566 6323 598
rect 6323 566 6355 598
rect 6355 566 6359 598
rect 6319 560 6359 566
rect 7527 4318 7567 4324
rect 7527 4286 7531 4318
rect 7531 4286 7563 4318
rect 7563 4286 7567 4318
rect 7527 4250 7567 4286
rect 7527 4218 7531 4250
rect 7531 4218 7563 4250
rect 7563 4218 7567 4250
rect 7527 4182 7567 4218
rect 7527 4150 7531 4182
rect 7531 4150 7563 4182
rect 7563 4150 7567 4182
rect 7527 4114 7567 4150
rect 7527 4082 7531 4114
rect 7531 4082 7563 4114
rect 7563 4082 7567 4114
rect 7527 4046 7567 4082
rect 7527 4014 7531 4046
rect 7531 4014 7563 4046
rect 7563 4014 7567 4046
rect 7527 3978 7567 4014
rect 7527 3946 7531 3978
rect 7531 3946 7563 3978
rect 7563 3946 7567 3978
rect 7527 3910 7567 3946
rect 7527 3878 7531 3910
rect 7531 3878 7563 3910
rect 7563 3878 7567 3910
rect 7527 3842 7567 3878
rect 7527 3810 7531 3842
rect 7531 3810 7563 3842
rect 7563 3810 7567 3842
rect 7527 3774 7567 3810
rect 7527 3742 7531 3774
rect 7531 3742 7563 3774
rect 7563 3742 7567 3774
rect 7527 3706 7567 3742
rect 7527 3674 7531 3706
rect 7531 3674 7563 3706
rect 7563 3674 7567 3706
rect 7527 3638 7567 3674
rect 7527 3606 7531 3638
rect 7531 3606 7563 3638
rect 7563 3606 7567 3638
rect 7527 3570 7567 3606
rect 7527 3538 7531 3570
rect 7531 3538 7563 3570
rect 7563 3538 7567 3570
rect 7527 3502 7567 3538
rect 7527 3470 7531 3502
rect 7531 3470 7563 3502
rect 7563 3470 7567 3502
rect 7527 3464 7567 3470
rect 7184 3350 7306 3356
rect 7184 3318 7229 3350
rect 7229 3318 7261 3350
rect 7261 3318 7306 3350
rect 7184 3282 7306 3318
rect 7184 3250 7229 3282
rect 7229 3250 7261 3282
rect 7261 3250 7306 3282
rect 7184 3214 7306 3250
rect 7184 3182 7229 3214
rect 7229 3182 7261 3214
rect 7261 3182 7306 3214
rect 7184 3146 7306 3182
rect 7184 3114 7229 3146
rect 7229 3114 7261 3146
rect 7261 3114 7306 3146
rect 7184 3078 7306 3114
rect 7184 3046 7229 3078
rect 7229 3046 7261 3078
rect 7261 3046 7306 3078
rect 7184 3010 7306 3046
rect 7184 2978 7229 3010
rect 7229 2978 7261 3010
rect 7261 2978 7306 3010
rect 7184 2942 7306 2978
rect 7184 2910 7229 2942
rect 7229 2910 7261 2942
rect 7261 2910 7306 2942
rect 7184 2874 7306 2910
rect 7184 2842 7229 2874
rect 7229 2842 7261 2874
rect 7261 2842 7306 2874
rect 7184 2806 7306 2842
rect 7184 2774 7229 2806
rect 7229 2774 7261 2806
rect 7261 2774 7306 2806
rect 7184 2738 7306 2774
rect 7184 2706 7229 2738
rect 7229 2706 7261 2738
rect 7261 2706 7306 2738
rect 7184 2670 7306 2706
rect 7184 2638 7229 2670
rect 7229 2638 7261 2670
rect 7261 2638 7306 2670
rect 7184 2602 7306 2638
rect 7184 2570 7229 2602
rect 7229 2570 7261 2602
rect 7261 2570 7306 2602
rect 7184 2534 7306 2570
rect 7184 2502 7229 2534
rect 7229 2502 7261 2534
rect 7261 2502 7306 2534
rect 7184 2496 7306 2502
rect 6923 2382 6963 2388
rect 6923 2350 6927 2382
rect 6927 2350 6959 2382
rect 6959 2350 6963 2382
rect 6923 2314 6963 2350
rect 6923 2282 6927 2314
rect 6927 2282 6959 2314
rect 6959 2282 6963 2314
rect 6923 2246 6963 2282
rect 6923 2214 6927 2246
rect 6927 2214 6959 2246
rect 6959 2214 6963 2246
rect 6923 2178 6963 2214
rect 6923 2146 6927 2178
rect 6927 2146 6959 2178
rect 6959 2146 6963 2178
rect 6923 2110 6963 2146
rect 6923 2078 6927 2110
rect 6927 2078 6959 2110
rect 6959 2078 6963 2110
rect 6923 2042 6963 2078
rect 6923 2010 6927 2042
rect 6927 2010 6959 2042
rect 6959 2010 6963 2042
rect 6923 1974 6963 2010
rect 6923 1942 6927 1974
rect 6927 1942 6959 1974
rect 6959 1942 6963 1974
rect 6923 1906 6963 1942
rect 6923 1874 6927 1906
rect 6927 1874 6959 1906
rect 6959 1874 6963 1906
rect 6923 1838 6963 1874
rect 6923 1806 6927 1838
rect 6927 1806 6959 1838
rect 6959 1806 6963 1838
rect 6923 1770 6963 1806
rect 6923 1738 6927 1770
rect 6927 1738 6959 1770
rect 6959 1738 6963 1770
rect 6923 1702 6963 1738
rect 6923 1670 6927 1702
rect 6927 1670 6959 1702
rect 6959 1670 6963 1702
rect 6923 1634 6963 1670
rect 6923 1602 6927 1634
rect 6927 1602 6959 1634
rect 6959 1602 6963 1634
rect 6923 1566 6963 1602
rect 6923 1534 6927 1566
rect 6927 1534 6959 1566
rect 6959 1534 6963 1566
rect 6923 1528 6963 1534
rect 6580 1414 6702 1420
rect 6580 1382 6625 1414
rect 6625 1382 6657 1414
rect 6657 1382 6702 1414
rect 6580 1346 6702 1382
rect 6580 1314 6625 1346
rect 6625 1314 6657 1346
rect 6657 1314 6702 1346
rect 6580 1278 6702 1314
rect 6580 1246 6625 1278
rect 6625 1246 6657 1278
rect 6657 1246 6702 1278
rect 6580 1210 6702 1246
rect 6580 1178 6625 1210
rect 6625 1178 6657 1210
rect 6657 1178 6702 1210
rect 6580 1142 6702 1178
rect 6580 1110 6625 1142
rect 6625 1110 6657 1142
rect 6657 1110 6702 1142
rect 6580 1074 6702 1110
rect 6580 1042 6625 1074
rect 6625 1042 6657 1074
rect 6657 1042 6702 1074
rect 6580 1006 6702 1042
rect 6580 974 6625 1006
rect 6625 974 6657 1006
rect 6657 974 6702 1006
rect 6580 938 6702 974
rect 6580 906 6625 938
rect 6625 906 6657 938
rect 6657 906 6702 938
rect 6580 870 6702 906
rect 6580 838 6625 870
rect 6625 838 6657 870
rect 6657 838 6702 870
rect 6580 802 6702 838
rect 6580 770 6625 802
rect 6625 770 6657 802
rect 6657 770 6702 802
rect 6580 734 6702 770
rect 6580 702 6625 734
rect 6625 702 6657 734
rect 6657 702 6702 734
rect 6580 666 6702 702
rect 6580 634 6625 666
rect 6625 634 6657 666
rect 6657 634 6702 666
rect 6580 598 6702 634
rect 6580 566 6625 598
rect 6625 566 6657 598
rect 6657 566 6702 598
rect 6580 560 6702 566
rect 7788 4318 7910 4324
rect 7788 4286 7833 4318
rect 7833 4286 7865 4318
rect 7865 4286 7910 4318
rect 7788 4250 7910 4286
rect 7788 4218 7833 4250
rect 7833 4218 7865 4250
rect 7865 4218 7910 4250
rect 7788 4182 7910 4218
rect 7788 4150 7833 4182
rect 7833 4150 7865 4182
rect 7865 4150 7910 4182
rect 7788 4114 7910 4150
rect 7788 4082 7833 4114
rect 7833 4082 7865 4114
rect 7865 4082 7910 4114
rect 7788 4046 7910 4082
rect 7788 4014 7833 4046
rect 7833 4014 7865 4046
rect 7865 4014 7910 4046
rect 7788 3978 7910 4014
rect 7788 3946 7833 3978
rect 7833 3946 7865 3978
rect 7865 3946 7910 3978
rect 7788 3910 7910 3946
rect 7788 3878 7833 3910
rect 7833 3878 7865 3910
rect 7865 3878 7910 3910
rect 7788 3842 7910 3878
rect 7788 3810 7833 3842
rect 7833 3810 7865 3842
rect 7865 3810 7910 3842
rect 7788 3774 7910 3810
rect 7788 3742 7833 3774
rect 7833 3742 7865 3774
rect 7865 3742 7910 3774
rect 7788 3706 7910 3742
rect 7788 3674 7833 3706
rect 7833 3674 7865 3706
rect 7865 3674 7910 3706
rect 7788 3638 7910 3674
rect 7788 3606 7833 3638
rect 7833 3606 7865 3638
rect 7865 3606 7910 3638
rect 7788 3570 7910 3606
rect 7788 3538 7833 3570
rect 7833 3538 7865 3570
rect 7865 3538 7910 3570
rect 7788 3502 7910 3538
rect 7788 3470 7833 3502
rect 7833 3470 7865 3502
rect 7865 3470 7910 3502
rect 7788 3464 7910 3470
rect 7527 3350 7567 3356
rect 7527 3318 7531 3350
rect 7531 3318 7563 3350
rect 7563 3318 7567 3350
rect 7527 3282 7567 3318
rect 7527 3250 7531 3282
rect 7531 3250 7563 3282
rect 7563 3250 7567 3282
rect 7527 3214 7567 3250
rect 7527 3182 7531 3214
rect 7531 3182 7563 3214
rect 7563 3182 7567 3214
rect 7527 3146 7567 3182
rect 7527 3114 7531 3146
rect 7531 3114 7563 3146
rect 7563 3114 7567 3146
rect 7527 3078 7567 3114
rect 7527 3046 7531 3078
rect 7531 3046 7563 3078
rect 7563 3046 7567 3078
rect 7527 3010 7567 3046
rect 7527 2978 7531 3010
rect 7531 2978 7563 3010
rect 7563 2978 7567 3010
rect 7527 2942 7567 2978
rect 7527 2910 7531 2942
rect 7531 2910 7563 2942
rect 7563 2910 7567 2942
rect 7527 2874 7567 2910
rect 7527 2842 7531 2874
rect 7531 2842 7563 2874
rect 7563 2842 7567 2874
rect 7527 2806 7567 2842
rect 7527 2774 7531 2806
rect 7531 2774 7563 2806
rect 7563 2774 7567 2806
rect 7527 2738 7567 2774
rect 7527 2706 7531 2738
rect 7531 2706 7563 2738
rect 7563 2706 7567 2738
rect 7527 2670 7567 2706
rect 7527 2638 7531 2670
rect 7531 2638 7563 2670
rect 7563 2638 7567 2670
rect 7527 2602 7567 2638
rect 7527 2570 7531 2602
rect 7531 2570 7563 2602
rect 7563 2570 7567 2602
rect 7527 2534 7567 2570
rect 7527 2502 7531 2534
rect 7531 2502 7563 2534
rect 7563 2502 7567 2534
rect 7527 2496 7567 2502
rect 7184 2382 7306 2388
rect 7184 2350 7229 2382
rect 7229 2350 7261 2382
rect 7261 2350 7306 2382
rect 7184 2314 7306 2350
rect 7184 2282 7229 2314
rect 7229 2282 7261 2314
rect 7261 2282 7306 2314
rect 7184 2246 7306 2282
rect 7184 2214 7229 2246
rect 7229 2214 7261 2246
rect 7261 2214 7306 2246
rect 7184 2178 7306 2214
rect 7184 2146 7229 2178
rect 7229 2146 7261 2178
rect 7261 2146 7306 2178
rect 7184 2110 7306 2146
rect 7184 2078 7229 2110
rect 7229 2078 7261 2110
rect 7261 2078 7306 2110
rect 7184 2042 7306 2078
rect 7184 2010 7229 2042
rect 7229 2010 7261 2042
rect 7261 2010 7306 2042
rect 7184 1974 7306 2010
rect 7184 1942 7229 1974
rect 7229 1942 7261 1974
rect 7261 1942 7306 1974
rect 7184 1906 7306 1942
rect 7184 1874 7229 1906
rect 7229 1874 7261 1906
rect 7261 1874 7306 1906
rect 7184 1838 7306 1874
rect 7184 1806 7229 1838
rect 7229 1806 7261 1838
rect 7261 1806 7306 1838
rect 7184 1770 7306 1806
rect 7184 1738 7229 1770
rect 7229 1738 7261 1770
rect 7261 1738 7306 1770
rect 7184 1702 7306 1738
rect 7184 1670 7229 1702
rect 7229 1670 7261 1702
rect 7261 1670 7306 1702
rect 7184 1634 7306 1670
rect 7184 1602 7229 1634
rect 7229 1602 7261 1634
rect 7261 1602 7306 1634
rect 7184 1566 7306 1602
rect 7184 1534 7229 1566
rect 7229 1534 7261 1566
rect 7261 1534 7306 1566
rect 7184 1528 7306 1534
rect 6923 1414 6963 1420
rect 6923 1382 6927 1414
rect 6927 1382 6959 1414
rect 6959 1382 6963 1414
rect 6923 1346 6963 1382
rect 6923 1314 6927 1346
rect 6927 1314 6959 1346
rect 6959 1314 6963 1346
rect 6923 1278 6963 1314
rect 6923 1246 6927 1278
rect 6927 1246 6959 1278
rect 6959 1246 6963 1278
rect 6923 1210 6963 1246
rect 6923 1178 6927 1210
rect 6927 1178 6959 1210
rect 6959 1178 6963 1210
rect 6923 1142 6963 1178
rect 6923 1110 6927 1142
rect 6927 1110 6959 1142
rect 6959 1110 6963 1142
rect 6923 1074 6963 1110
rect 6923 1042 6927 1074
rect 6927 1042 6959 1074
rect 6959 1042 6963 1074
rect 6923 1006 6963 1042
rect 6923 974 6927 1006
rect 6927 974 6959 1006
rect 6959 974 6963 1006
rect 6923 938 6963 974
rect 6923 906 6927 938
rect 6927 906 6959 938
rect 6959 906 6963 938
rect 6923 870 6963 906
rect 6923 838 6927 870
rect 6927 838 6959 870
rect 6959 838 6963 870
rect 6923 802 6963 838
rect 6923 770 6927 802
rect 6927 770 6959 802
rect 6959 770 6963 802
rect 6923 734 6963 770
rect 6923 702 6927 734
rect 6927 702 6959 734
rect 6959 702 6963 734
rect 6923 666 6963 702
rect 6923 634 6927 666
rect 6927 634 6959 666
rect 6959 634 6963 666
rect 6923 598 6963 634
rect 6923 566 6927 598
rect 6927 566 6959 598
rect 6959 566 6963 598
rect 6923 560 6963 566
rect 8131 4318 8171 4324
rect 8131 4286 8135 4318
rect 8135 4286 8167 4318
rect 8167 4286 8171 4318
rect 8131 4250 8171 4286
rect 8131 4218 8135 4250
rect 8135 4218 8167 4250
rect 8167 4218 8171 4250
rect 8131 4182 8171 4218
rect 8131 4150 8135 4182
rect 8135 4150 8167 4182
rect 8167 4150 8171 4182
rect 8131 4114 8171 4150
rect 8131 4082 8135 4114
rect 8135 4082 8167 4114
rect 8167 4082 8171 4114
rect 8131 4046 8171 4082
rect 8131 4014 8135 4046
rect 8135 4014 8167 4046
rect 8167 4014 8171 4046
rect 8131 3978 8171 4014
rect 8131 3946 8135 3978
rect 8135 3946 8167 3978
rect 8167 3946 8171 3978
rect 8131 3910 8171 3946
rect 8131 3878 8135 3910
rect 8135 3878 8167 3910
rect 8167 3878 8171 3910
rect 8131 3842 8171 3878
rect 8131 3810 8135 3842
rect 8135 3810 8167 3842
rect 8167 3810 8171 3842
rect 8131 3774 8171 3810
rect 8131 3742 8135 3774
rect 8135 3742 8167 3774
rect 8167 3742 8171 3774
rect 8131 3706 8171 3742
rect 8131 3674 8135 3706
rect 8135 3674 8167 3706
rect 8167 3674 8171 3706
rect 8131 3638 8171 3674
rect 8131 3606 8135 3638
rect 8135 3606 8167 3638
rect 8167 3606 8171 3638
rect 8131 3570 8171 3606
rect 8131 3538 8135 3570
rect 8135 3538 8167 3570
rect 8167 3538 8171 3570
rect 8131 3502 8171 3538
rect 8131 3470 8135 3502
rect 8135 3470 8167 3502
rect 8167 3470 8171 3502
rect 8131 3464 8171 3470
rect 7788 3350 7910 3356
rect 7788 3318 7833 3350
rect 7833 3318 7865 3350
rect 7865 3318 7910 3350
rect 7788 3282 7910 3318
rect 7788 3250 7833 3282
rect 7833 3250 7865 3282
rect 7865 3250 7910 3282
rect 7788 3214 7910 3250
rect 7788 3182 7833 3214
rect 7833 3182 7865 3214
rect 7865 3182 7910 3214
rect 7788 3146 7910 3182
rect 7788 3114 7833 3146
rect 7833 3114 7865 3146
rect 7865 3114 7910 3146
rect 7788 3078 7910 3114
rect 7788 3046 7833 3078
rect 7833 3046 7865 3078
rect 7865 3046 7910 3078
rect 7788 3010 7910 3046
rect 7788 2978 7833 3010
rect 7833 2978 7865 3010
rect 7865 2978 7910 3010
rect 7788 2942 7910 2978
rect 7788 2910 7833 2942
rect 7833 2910 7865 2942
rect 7865 2910 7910 2942
rect 7788 2874 7910 2910
rect 7788 2842 7833 2874
rect 7833 2842 7865 2874
rect 7865 2842 7910 2874
rect 7788 2806 7910 2842
rect 7788 2774 7833 2806
rect 7833 2774 7865 2806
rect 7865 2774 7910 2806
rect 7788 2738 7910 2774
rect 7788 2706 7833 2738
rect 7833 2706 7865 2738
rect 7865 2706 7910 2738
rect 7788 2670 7910 2706
rect 7788 2638 7833 2670
rect 7833 2638 7865 2670
rect 7865 2638 7910 2670
rect 7788 2602 7910 2638
rect 7788 2570 7833 2602
rect 7833 2570 7865 2602
rect 7865 2570 7910 2602
rect 7788 2534 7910 2570
rect 7788 2502 7833 2534
rect 7833 2502 7865 2534
rect 7865 2502 7910 2534
rect 7788 2496 7910 2502
rect 7527 2382 7567 2388
rect 7527 2350 7531 2382
rect 7531 2350 7563 2382
rect 7563 2350 7567 2382
rect 7527 2314 7567 2350
rect 7527 2282 7531 2314
rect 7531 2282 7563 2314
rect 7563 2282 7567 2314
rect 7527 2246 7567 2282
rect 7527 2214 7531 2246
rect 7531 2214 7563 2246
rect 7563 2214 7567 2246
rect 7527 2178 7567 2214
rect 7527 2146 7531 2178
rect 7531 2146 7563 2178
rect 7563 2146 7567 2178
rect 7527 2110 7567 2146
rect 7527 2078 7531 2110
rect 7531 2078 7563 2110
rect 7563 2078 7567 2110
rect 7527 2042 7567 2078
rect 7527 2010 7531 2042
rect 7531 2010 7563 2042
rect 7563 2010 7567 2042
rect 7527 1974 7567 2010
rect 7527 1942 7531 1974
rect 7531 1942 7563 1974
rect 7563 1942 7567 1974
rect 7527 1906 7567 1942
rect 7527 1874 7531 1906
rect 7531 1874 7563 1906
rect 7563 1874 7567 1906
rect 7527 1838 7567 1874
rect 7527 1806 7531 1838
rect 7531 1806 7563 1838
rect 7563 1806 7567 1838
rect 7527 1770 7567 1806
rect 7527 1738 7531 1770
rect 7531 1738 7563 1770
rect 7563 1738 7567 1770
rect 7527 1702 7567 1738
rect 7527 1670 7531 1702
rect 7531 1670 7563 1702
rect 7563 1670 7567 1702
rect 7527 1634 7567 1670
rect 7527 1602 7531 1634
rect 7531 1602 7563 1634
rect 7563 1602 7567 1634
rect 7527 1566 7567 1602
rect 7527 1534 7531 1566
rect 7531 1534 7563 1566
rect 7563 1534 7567 1566
rect 7527 1528 7567 1534
rect 7184 1414 7306 1420
rect 7184 1382 7229 1414
rect 7229 1382 7261 1414
rect 7261 1382 7306 1414
rect 7184 1346 7306 1382
rect 7184 1314 7229 1346
rect 7229 1314 7261 1346
rect 7261 1314 7306 1346
rect 7184 1278 7306 1314
rect 7184 1246 7229 1278
rect 7229 1246 7261 1278
rect 7261 1246 7306 1278
rect 7184 1210 7306 1246
rect 7184 1178 7229 1210
rect 7229 1178 7261 1210
rect 7261 1178 7306 1210
rect 7184 1142 7306 1178
rect 7184 1110 7229 1142
rect 7229 1110 7261 1142
rect 7261 1110 7306 1142
rect 7184 1074 7306 1110
rect 7184 1042 7229 1074
rect 7229 1042 7261 1074
rect 7261 1042 7306 1074
rect 7184 1006 7306 1042
rect 7184 974 7229 1006
rect 7229 974 7261 1006
rect 7261 974 7306 1006
rect 7184 938 7306 974
rect 7184 906 7229 938
rect 7229 906 7261 938
rect 7261 906 7306 938
rect 7184 870 7306 906
rect 7184 838 7229 870
rect 7229 838 7261 870
rect 7261 838 7306 870
rect 7184 802 7306 838
rect 7184 770 7229 802
rect 7229 770 7261 802
rect 7261 770 7306 802
rect 7184 734 7306 770
rect 7184 702 7229 734
rect 7229 702 7261 734
rect 7261 702 7306 734
rect 7184 666 7306 702
rect 7184 634 7229 666
rect 7229 634 7261 666
rect 7261 634 7306 666
rect 7184 598 7306 634
rect 7184 566 7229 598
rect 7229 566 7261 598
rect 7261 566 7306 598
rect 7184 560 7306 566
rect 8392 4318 8514 4324
rect 8392 4286 8437 4318
rect 8437 4286 8469 4318
rect 8469 4286 8514 4318
rect 8392 4250 8514 4286
rect 8392 4218 8437 4250
rect 8437 4218 8469 4250
rect 8469 4218 8514 4250
rect 8392 4182 8514 4218
rect 8392 4150 8437 4182
rect 8437 4150 8469 4182
rect 8469 4150 8514 4182
rect 8392 4114 8514 4150
rect 8392 4082 8437 4114
rect 8437 4082 8469 4114
rect 8469 4082 8514 4114
rect 8392 4046 8514 4082
rect 8392 4014 8437 4046
rect 8437 4014 8469 4046
rect 8469 4014 8514 4046
rect 8392 3978 8514 4014
rect 8392 3946 8437 3978
rect 8437 3946 8469 3978
rect 8469 3946 8514 3978
rect 8392 3910 8514 3946
rect 8392 3878 8437 3910
rect 8437 3878 8469 3910
rect 8469 3878 8514 3910
rect 8392 3842 8514 3878
rect 8392 3810 8437 3842
rect 8437 3810 8469 3842
rect 8469 3810 8514 3842
rect 8392 3774 8514 3810
rect 8392 3742 8437 3774
rect 8437 3742 8469 3774
rect 8469 3742 8514 3774
rect 8392 3706 8514 3742
rect 8392 3674 8437 3706
rect 8437 3674 8469 3706
rect 8469 3674 8514 3706
rect 8392 3638 8514 3674
rect 8392 3606 8437 3638
rect 8437 3606 8469 3638
rect 8469 3606 8514 3638
rect 8392 3570 8514 3606
rect 8392 3538 8437 3570
rect 8437 3538 8469 3570
rect 8469 3538 8514 3570
rect 8392 3502 8514 3538
rect 8392 3470 8437 3502
rect 8437 3470 8469 3502
rect 8469 3470 8514 3502
rect 8392 3464 8514 3470
rect 8131 3350 8171 3356
rect 8131 3318 8135 3350
rect 8135 3318 8167 3350
rect 8167 3318 8171 3350
rect 8131 3282 8171 3318
rect 8131 3250 8135 3282
rect 8135 3250 8167 3282
rect 8167 3250 8171 3282
rect 8131 3214 8171 3250
rect 8131 3182 8135 3214
rect 8135 3182 8167 3214
rect 8167 3182 8171 3214
rect 8131 3146 8171 3182
rect 8131 3114 8135 3146
rect 8135 3114 8167 3146
rect 8167 3114 8171 3146
rect 8131 3078 8171 3114
rect 8131 3046 8135 3078
rect 8135 3046 8167 3078
rect 8167 3046 8171 3078
rect 8131 3010 8171 3046
rect 8131 2978 8135 3010
rect 8135 2978 8167 3010
rect 8167 2978 8171 3010
rect 8131 2942 8171 2978
rect 8131 2910 8135 2942
rect 8135 2910 8167 2942
rect 8167 2910 8171 2942
rect 8131 2874 8171 2910
rect 8131 2842 8135 2874
rect 8135 2842 8167 2874
rect 8167 2842 8171 2874
rect 8131 2806 8171 2842
rect 8131 2774 8135 2806
rect 8135 2774 8167 2806
rect 8167 2774 8171 2806
rect 8131 2738 8171 2774
rect 8131 2706 8135 2738
rect 8135 2706 8167 2738
rect 8167 2706 8171 2738
rect 8131 2670 8171 2706
rect 8131 2638 8135 2670
rect 8135 2638 8167 2670
rect 8167 2638 8171 2670
rect 8131 2602 8171 2638
rect 8131 2570 8135 2602
rect 8135 2570 8167 2602
rect 8167 2570 8171 2602
rect 8131 2534 8171 2570
rect 8131 2502 8135 2534
rect 8135 2502 8167 2534
rect 8167 2502 8171 2534
rect 8131 2496 8171 2502
rect 7788 2382 7910 2388
rect 7788 2350 7833 2382
rect 7833 2350 7865 2382
rect 7865 2350 7910 2382
rect 7788 2314 7910 2350
rect 7788 2282 7833 2314
rect 7833 2282 7865 2314
rect 7865 2282 7910 2314
rect 7788 2246 7910 2282
rect 7788 2214 7833 2246
rect 7833 2214 7865 2246
rect 7865 2214 7910 2246
rect 7788 2178 7910 2214
rect 7788 2146 7833 2178
rect 7833 2146 7865 2178
rect 7865 2146 7910 2178
rect 7788 2110 7910 2146
rect 7788 2078 7833 2110
rect 7833 2078 7865 2110
rect 7865 2078 7910 2110
rect 7788 2042 7910 2078
rect 7788 2010 7833 2042
rect 7833 2010 7865 2042
rect 7865 2010 7910 2042
rect 7788 1974 7910 2010
rect 7788 1942 7833 1974
rect 7833 1942 7865 1974
rect 7865 1942 7910 1974
rect 7788 1906 7910 1942
rect 7788 1874 7833 1906
rect 7833 1874 7865 1906
rect 7865 1874 7910 1906
rect 7788 1838 7910 1874
rect 7788 1806 7833 1838
rect 7833 1806 7865 1838
rect 7865 1806 7910 1838
rect 7788 1770 7910 1806
rect 7788 1738 7833 1770
rect 7833 1738 7865 1770
rect 7865 1738 7910 1770
rect 7788 1702 7910 1738
rect 7788 1670 7833 1702
rect 7833 1670 7865 1702
rect 7865 1670 7910 1702
rect 7788 1634 7910 1670
rect 7788 1602 7833 1634
rect 7833 1602 7865 1634
rect 7865 1602 7910 1634
rect 7788 1566 7910 1602
rect 7788 1534 7833 1566
rect 7833 1534 7865 1566
rect 7865 1534 7910 1566
rect 7788 1528 7910 1534
rect 7527 1414 7567 1420
rect 7527 1382 7531 1414
rect 7531 1382 7563 1414
rect 7563 1382 7567 1414
rect 7527 1346 7567 1382
rect 7527 1314 7531 1346
rect 7531 1314 7563 1346
rect 7563 1314 7567 1346
rect 7527 1278 7567 1314
rect 7527 1246 7531 1278
rect 7531 1246 7563 1278
rect 7563 1246 7567 1278
rect 7527 1210 7567 1246
rect 7527 1178 7531 1210
rect 7531 1178 7563 1210
rect 7563 1178 7567 1210
rect 7527 1142 7567 1178
rect 7527 1110 7531 1142
rect 7531 1110 7563 1142
rect 7563 1110 7567 1142
rect 7527 1074 7567 1110
rect 7527 1042 7531 1074
rect 7531 1042 7563 1074
rect 7563 1042 7567 1074
rect 7527 1006 7567 1042
rect 7527 974 7531 1006
rect 7531 974 7563 1006
rect 7563 974 7567 1006
rect 7527 938 7567 974
rect 7527 906 7531 938
rect 7531 906 7563 938
rect 7563 906 7567 938
rect 7527 870 7567 906
rect 7527 838 7531 870
rect 7531 838 7563 870
rect 7563 838 7567 870
rect 7527 802 7567 838
rect 7527 770 7531 802
rect 7531 770 7563 802
rect 7563 770 7567 802
rect 7527 734 7567 770
rect 7527 702 7531 734
rect 7531 702 7563 734
rect 7563 702 7567 734
rect 7527 666 7567 702
rect 7527 634 7531 666
rect 7531 634 7563 666
rect 7563 634 7567 666
rect 7527 598 7567 634
rect 7527 566 7531 598
rect 7531 566 7563 598
rect 7563 566 7567 598
rect 7527 560 7567 566
rect 8735 4318 8775 4324
rect 8735 4286 8739 4318
rect 8739 4286 8771 4318
rect 8771 4286 8775 4318
rect 8735 4250 8775 4286
rect 8735 4218 8739 4250
rect 8739 4218 8771 4250
rect 8771 4218 8775 4250
rect 8735 4182 8775 4218
rect 8735 4150 8739 4182
rect 8739 4150 8771 4182
rect 8771 4150 8775 4182
rect 8735 4114 8775 4150
rect 8735 4082 8739 4114
rect 8739 4082 8771 4114
rect 8771 4082 8775 4114
rect 8735 4046 8775 4082
rect 8735 4014 8739 4046
rect 8739 4014 8771 4046
rect 8771 4014 8775 4046
rect 8735 3978 8775 4014
rect 8735 3946 8739 3978
rect 8739 3946 8771 3978
rect 8771 3946 8775 3978
rect 8735 3910 8775 3946
rect 8735 3878 8739 3910
rect 8739 3878 8771 3910
rect 8771 3878 8775 3910
rect 8735 3842 8775 3878
rect 8735 3810 8739 3842
rect 8739 3810 8771 3842
rect 8771 3810 8775 3842
rect 8735 3774 8775 3810
rect 8735 3742 8739 3774
rect 8739 3742 8771 3774
rect 8771 3742 8775 3774
rect 8735 3706 8775 3742
rect 8735 3674 8739 3706
rect 8739 3674 8771 3706
rect 8771 3674 8775 3706
rect 8735 3638 8775 3674
rect 8735 3606 8739 3638
rect 8739 3606 8771 3638
rect 8771 3606 8775 3638
rect 8735 3570 8775 3606
rect 8735 3538 8739 3570
rect 8739 3538 8771 3570
rect 8771 3538 8775 3570
rect 8735 3502 8775 3538
rect 8735 3470 8739 3502
rect 8739 3470 8771 3502
rect 8771 3470 8775 3502
rect 8735 3464 8775 3470
rect 8392 3350 8514 3356
rect 8392 3318 8437 3350
rect 8437 3318 8469 3350
rect 8469 3318 8514 3350
rect 8392 3282 8514 3318
rect 8392 3250 8437 3282
rect 8437 3250 8469 3282
rect 8469 3250 8514 3282
rect 8392 3214 8514 3250
rect 8392 3182 8437 3214
rect 8437 3182 8469 3214
rect 8469 3182 8514 3214
rect 8392 3146 8514 3182
rect 8392 3114 8437 3146
rect 8437 3114 8469 3146
rect 8469 3114 8514 3146
rect 8392 3078 8514 3114
rect 8392 3046 8437 3078
rect 8437 3046 8469 3078
rect 8469 3046 8514 3078
rect 8392 3010 8514 3046
rect 8392 2978 8437 3010
rect 8437 2978 8469 3010
rect 8469 2978 8514 3010
rect 8392 2942 8514 2978
rect 8392 2910 8437 2942
rect 8437 2910 8469 2942
rect 8469 2910 8514 2942
rect 8392 2874 8514 2910
rect 8392 2842 8437 2874
rect 8437 2842 8469 2874
rect 8469 2842 8514 2874
rect 8392 2806 8514 2842
rect 8392 2774 8437 2806
rect 8437 2774 8469 2806
rect 8469 2774 8514 2806
rect 8392 2738 8514 2774
rect 8392 2706 8437 2738
rect 8437 2706 8469 2738
rect 8469 2706 8514 2738
rect 8392 2670 8514 2706
rect 8392 2638 8437 2670
rect 8437 2638 8469 2670
rect 8469 2638 8514 2670
rect 8392 2602 8514 2638
rect 8392 2570 8437 2602
rect 8437 2570 8469 2602
rect 8469 2570 8514 2602
rect 8392 2534 8514 2570
rect 8392 2502 8437 2534
rect 8437 2502 8469 2534
rect 8469 2502 8514 2534
rect 8392 2496 8514 2502
rect 8131 2382 8171 2388
rect 8131 2350 8135 2382
rect 8135 2350 8167 2382
rect 8167 2350 8171 2382
rect 8131 2314 8171 2350
rect 8131 2282 8135 2314
rect 8135 2282 8167 2314
rect 8167 2282 8171 2314
rect 8131 2246 8171 2282
rect 8131 2214 8135 2246
rect 8135 2214 8167 2246
rect 8167 2214 8171 2246
rect 8131 2178 8171 2214
rect 8131 2146 8135 2178
rect 8135 2146 8167 2178
rect 8167 2146 8171 2178
rect 8131 2110 8171 2146
rect 8131 2078 8135 2110
rect 8135 2078 8167 2110
rect 8167 2078 8171 2110
rect 8131 2042 8171 2078
rect 8131 2010 8135 2042
rect 8135 2010 8167 2042
rect 8167 2010 8171 2042
rect 8131 1974 8171 2010
rect 8131 1942 8135 1974
rect 8135 1942 8167 1974
rect 8167 1942 8171 1974
rect 8131 1906 8171 1942
rect 8131 1874 8135 1906
rect 8135 1874 8167 1906
rect 8167 1874 8171 1906
rect 8131 1838 8171 1874
rect 8131 1806 8135 1838
rect 8135 1806 8167 1838
rect 8167 1806 8171 1838
rect 8131 1770 8171 1806
rect 8131 1738 8135 1770
rect 8135 1738 8167 1770
rect 8167 1738 8171 1770
rect 8131 1702 8171 1738
rect 8131 1670 8135 1702
rect 8135 1670 8167 1702
rect 8167 1670 8171 1702
rect 8131 1634 8171 1670
rect 8131 1602 8135 1634
rect 8135 1602 8167 1634
rect 8167 1602 8171 1634
rect 8131 1566 8171 1602
rect 8131 1534 8135 1566
rect 8135 1534 8167 1566
rect 8167 1534 8171 1566
rect 8131 1528 8171 1534
rect 7788 1414 7910 1420
rect 7788 1382 7833 1414
rect 7833 1382 7865 1414
rect 7865 1382 7910 1414
rect 7788 1346 7910 1382
rect 7788 1314 7833 1346
rect 7833 1314 7865 1346
rect 7865 1314 7910 1346
rect 7788 1278 7910 1314
rect 7788 1246 7833 1278
rect 7833 1246 7865 1278
rect 7865 1246 7910 1278
rect 7788 1210 7910 1246
rect 7788 1178 7833 1210
rect 7833 1178 7865 1210
rect 7865 1178 7910 1210
rect 7788 1142 7910 1178
rect 7788 1110 7833 1142
rect 7833 1110 7865 1142
rect 7865 1110 7910 1142
rect 7788 1074 7910 1110
rect 7788 1042 7833 1074
rect 7833 1042 7865 1074
rect 7865 1042 7910 1074
rect 7788 1006 7910 1042
rect 7788 974 7833 1006
rect 7833 974 7865 1006
rect 7865 974 7910 1006
rect 7788 938 7910 974
rect 7788 906 7833 938
rect 7833 906 7865 938
rect 7865 906 7910 938
rect 7788 870 7910 906
rect 7788 838 7833 870
rect 7833 838 7865 870
rect 7865 838 7910 870
rect 7788 802 7910 838
rect 7788 770 7833 802
rect 7833 770 7865 802
rect 7865 770 7910 802
rect 7788 734 7910 770
rect 7788 702 7833 734
rect 7833 702 7865 734
rect 7865 702 7910 734
rect 7788 666 7910 702
rect 7788 634 7833 666
rect 7833 634 7865 666
rect 7865 634 7910 666
rect 7788 598 7910 634
rect 7788 566 7833 598
rect 7833 566 7865 598
rect 7865 566 7910 598
rect 7788 560 7910 566
rect 8996 4318 9118 4324
rect 8996 4286 9041 4318
rect 9041 4286 9073 4318
rect 9073 4286 9118 4318
rect 8996 4250 9118 4286
rect 8996 4218 9041 4250
rect 9041 4218 9073 4250
rect 9073 4218 9118 4250
rect 8996 4182 9118 4218
rect 8996 4150 9041 4182
rect 9041 4150 9073 4182
rect 9073 4150 9118 4182
rect 8996 4114 9118 4150
rect 8996 4082 9041 4114
rect 9041 4082 9073 4114
rect 9073 4082 9118 4114
rect 8996 4046 9118 4082
rect 8996 4014 9041 4046
rect 9041 4014 9073 4046
rect 9073 4014 9118 4046
rect 8996 3978 9118 4014
rect 8996 3946 9041 3978
rect 9041 3946 9073 3978
rect 9073 3946 9118 3978
rect 8996 3910 9118 3946
rect 8996 3878 9041 3910
rect 9041 3878 9073 3910
rect 9073 3878 9118 3910
rect 8996 3842 9118 3878
rect 8996 3810 9041 3842
rect 9041 3810 9073 3842
rect 9073 3810 9118 3842
rect 8996 3774 9118 3810
rect 8996 3742 9041 3774
rect 9041 3742 9073 3774
rect 9073 3742 9118 3774
rect 8996 3706 9118 3742
rect 8996 3674 9041 3706
rect 9041 3674 9073 3706
rect 9073 3674 9118 3706
rect 8996 3638 9118 3674
rect 8996 3606 9041 3638
rect 9041 3606 9073 3638
rect 9073 3606 9118 3638
rect 8996 3570 9118 3606
rect 8996 3538 9041 3570
rect 9041 3538 9073 3570
rect 9073 3538 9118 3570
rect 8996 3502 9118 3538
rect 8996 3470 9041 3502
rect 9041 3470 9073 3502
rect 9073 3470 9118 3502
rect 8996 3464 9118 3470
rect 8735 3350 8775 3356
rect 8735 3318 8739 3350
rect 8739 3318 8771 3350
rect 8771 3318 8775 3350
rect 8735 3282 8775 3318
rect 8735 3250 8739 3282
rect 8739 3250 8771 3282
rect 8771 3250 8775 3282
rect 8735 3214 8775 3250
rect 8735 3182 8739 3214
rect 8739 3182 8771 3214
rect 8771 3182 8775 3214
rect 8735 3146 8775 3182
rect 8735 3114 8739 3146
rect 8739 3114 8771 3146
rect 8771 3114 8775 3146
rect 8735 3078 8775 3114
rect 8735 3046 8739 3078
rect 8739 3046 8771 3078
rect 8771 3046 8775 3078
rect 8735 3010 8775 3046
rect 8735 2978 8739 3010
rect 8739 2978 8771 3010
rect 8771 2978 8775 3010
rect 8735 2942 8775 2978
rect 8735 2910 8739 2942
rect 8739 2910 8771 2942
rect 8771 2910 8775 2942
rect 8735 2874 8775 2910
rect 8735 2842 8739 2874
rect 8739 2842 8771 2874
rect 8771 2842 8775 2874
rect 8735 2806 8775 2842
rect 8735 2774 8739 2806
rect 8739 2774 8771 2806
rect 8771 2774 8775 2806
rect 8735 2738 8775 2774
rect 8735 2706 8739 2738
rect 8739 2706 8771 2738
rect 8771 2706 8775 2738
rect 8735 2670 8775 2706
rect 8735 2638 8739 2670
rect 8739 2638 8771 2670
rect 8771 2638 8775 2670
rect 8735 2602 8775 2638
rect 8735 2570 8739 2602
rect 8739 2570 8771 2602
rect 8771 2570 8775 2602
rect 8735 2534 8775 2570
rect 8735 2502 8739 2534
rect 8739 2502 8771 2534
rect 8771 2502 8775 2534
rect 8735 2496 8775 2502
rect 8392 2382 8514 2388
rect 8392 2350 8437 2382
rect 8437 2350 8469 2382
rect 8469 2350 8514 2382
rect 8392 2314 8514 2350
rect 8392 2282 8437 2314
rect 8437 2282 8469 2314
rect 8469 2282 8514 2314
rect 8392 2246 8514 2282
rect 8392 2214 8437 2246
rect 8437 2214 8469 2246
rect 8469 2214 8514 2246
rect 8392 2178 8514 2214
rect 8392 2146 8437 2178
rect 8437 2146 8469 2178
rect 8469 2146 8514 2178
rect 8392 2110 8514 2146
rect 8392 2078 8437 2110
rect 8437 2078 8469 2110
rect 8469 2078 8514 2110
rect 8392 2042 8514 2078
rect 8392 2010 8437 2042
rect 8437 2010 8469 2042
rect 8469 2010 8514 2042
rect 8392 1974 8514 2010
rect 8392 1942 8437 1974
rect 8437 1942 8469 1974
rect 8469 1942 8514 1974
rect 8392 1906 8514 1942
rect 8392 1874 8437 1906
rect 8437 1874 8469 1906
rect 8469 1874 8514 1906
rect 8392 1838 8514 1874
rect 8392 1806 8437 1838
rect 8437 1806 8469 1838
rect 8469 1806 8514 1838
rect 8392 1770 8514 1806
rect 8392 1738 8437 1770
rect 8437 1738 8469 1770
rect 8469 1738 8514 1770
rect 8392 1702 8514 1738
rect 8392 1670 8437 1702
rect 8437 1670 8469 1702
rect 8469 1670 8514 1702
rect 8392 1634 8514 1670
rect 8392 1602 8437 1634
rect 8437 1602 8469 1634
rect 8469 1602 8514 1634
rect 8392 1566 8514 1602
rect 8392 1534 8437 1566
rect 8437 1534 8469 1566
rect 8469 1534 8514 1566
rect 8392 1528 8514 1534
rect 8131 1414 8171 1420
rect 8131 1382 8135 1414
rect 8135 1382 8167 1414
rect 8167 1382 8171 1414
rect 8131 1346 8171 1382
rect 8131 1314 8135 1346
rect 8135 1314 8167 1346
rect 8167 1314 8171 1346
rect 8131 1278 8171 1314
rect 8131 1246 8135 1278
rect 8135 1246 8167 1278
rect 8167 1246 8171 1278
rect 8131 1210 8171 1246
rect 8131 1178 8135 1210
rect 8135 1178 8167 1210
rect 8167 1178 8171 1210
rect 8131 1142 8171 1178
rect 8131 1110 8135 1142
rect 8135 1110 8167 1142
rect 8167 1110 8171 1142
rect 8131 1074 8171 1110
rect 8131 1042 8135 1074
rect 8135 1042 8167 1074
rect 8167 1042 8171 1074
rect 8131 1006 8171 1042
rect 8131 974 8135 1006
rect 8135 974 8167 1006
rect 8167 974 8171 1006
rect 8131 938 8171 974
rect 8131 906 8135 938
rect 8135 906 8167 938
rect 8167 906 8171 938
rect 8131 870 8171 906
rect 8131 838 8135 870
rect 8135 838 8167 870
rect 8167 838 8171 870
rect 8131 802 8171 838
rect 8131 770 8135 802
rect 8135 770 8167 802
rect 8167 770 8171 802
rect 8131 734 8171 770
rect 8131 702 8135 734
rect 8135 702 8167 734
rect 8167 702 8171 734
rect 8131 666 8171 702
rect 8131 634 8135 666
rect 8135 634 8167 666
rect 8167 634 8171 666
rect 8131 598 8171 634
rect 8131 566 8135 598
rect 8135 566 8167 598
rect 8167 566 8171 598
rect 8131 560 8171 566
rect 9339 4318 9379 4324
rect 9339 4286 9343 4318
rect 9343 4286 9375 4318
rect 9375 4286 9379 4318
rect 9339 4250 9379 4286
rect 9339 4218 9343 4250
rect 9343 4218 9375 4250
rect 9375 4218 9379 4250
rect 9339 4182 9379 4218
rect 9339 4150 9343 4182
rect 9343 4150 9375 4182
rect 9375 4150 9379 4182
rect 9339 4114 9379 4150
rect 9339 4082 9343 4114
rect 9343 4082 9375 4114
rect 9375 4082 9379 4114
rect 9339 4046 9379 4082
rect 9339 4014 9343 4046
rect 9343 4014 9375 4046
rect 9375 4014 9379 4046
rect 9339 3978 9379 4014
rect 9339 3946 9343 3978
rect 9343 3946 9375 3978
rect 9375 3946 9379 3978
rect 9339 3910 9379 3946
rect 9339 3878 9343 3910
rect 9343 3878 9375 3910
rect 9375 3878 9379 3910
rect 9339 3842 9379 3878
rect 9339 3810 9343 3842
rect 9343 3810 9375 3842
rect 9375 3810 9379 3842
rect 9339 3774 9379 3810
rect 9339 3742 9343 3774
rect 9343 3742 9375 3774
rect 9375 3742 9379 3774
rect 9339 3706 9379 3742
rect 9339 3674 9343 3706
rect 9343 3674 9375 3706
rect 9375 3674 9379 3706
rect 9339 3638 9379 3674
rect 9339 3606 9343 3638
rect 9343 3606 9375 3638
rect 9375 3606 9379 3638
rect 9339 3570 9379 3606
rect 9339 3538 9343 3570
rect 9343 3538 9375 3570
rect 9375 3538 9379 3570
rect 9339 3502 9379 3538
rect 9339 3470 9343 3502
rect 9343 3470 9375 3502
rect 9375 3470 9379 3502
rect 9339 3464 9379 3470
rect 8996 3350 9118 3356
rect 8996 3318 9041 3350
rect 9041 3318 9073 3350
rect 9073 3318 9118 3350
rect 8996 3282 9118 3318
rect 8996 3250 9041 3282
rect 9041 3250 9073 3282
rect 9073 3250 9118 3282
rect 8996 3214 9118 3250
rect 8996 3182 9041 3214
rect 9041 3182 9073 3214
rect 9073 3182 9118 3214
rect 8996 3146 9118 3182
rect 8996 3114 9041 3146
rect 9041 3114 9073 3146
rect 9073 3114 9118 3146
rect 8996 3078 9118 3114
rect 8996 3046 9041 3078
rect 9041 3046 9073 3078
rect 9073 3046 9118 3078
rect 8996 3010 9118 3046
rect 8996 2978 9041 3010
rect 9041 2978 9073 3010
rect 9073 2978 9118 3010
rect 8996 2942 9118 2978
rect 8996 2910 9041 2942
rect 9041 2910 9073 2942
rect 9073 2910 9118 2942
rect 8996 2874 9118 2910
rect 8996 2842 9041 2874
rect 9041 2842 9073 2874
rect 9073 2842 9118 2874
rect 8996 2806 9118 2842
rect 8996 2774 9041 2806
rect 9041 2774 9073 2806
rect 9073 2774 9118 2806
rect 8996 2738 9118 2774
rect 8996 2706 9041 2738
rect 9041 2706 9073 2738
rect 9073 2706 9118 2738
rect 8996 2670 9118 2706
rect 8996 2638 9041 2670
rect 9041 2638 9073 2670
rect 9073 2638 9118 2670
rect 8996 2602 9118 2638
rect 8996 2570 9041 2602
rect 9041 2570 9073 2602
rect 9073 2570 9118 2602
rect 8996 2534 9118 2570
rect 8996 2502 9041 2534
rect 9041 2502 9073 2534
rect 9073 2502 9118 2534
rect 8996 2496 9118 2502
rect 8735 2382 8775 2388
rect 8735 2350 8739 2382
rect 8739 2350 8771 2382
rect 8771 2350 8775 2382
rect 8735 2314 8775 2350
rect 8735 2282 8739 2314
rect 8739 2282 8771 2314
rect 8771 2282 8775 2314
rect 8735 2246 8775 2282
rect 8735 2214 8739 2246
rect 8739 2214 8771 2246
rect 8771 2214 8775 2246
rect 8735 2178 8775 2214
rect 8735 2146 8739 2178
rect 8739 2146 8771 2178
rect 8771 2146 8775 2178
rect 8735 2110 8775 2146
rect 8735 2078 8739 2110
rect 8739 2078 8771 2110
rect 8771 2078 8775 2110
rect 8735 2042 8775 2078
rect 8735 2010 8739 2042
rect 8739 2010 8771 2042
rect 8771 2010 8775 2042
rect 8735 1974 8775 2010
rect 8735 1942 8739 1974
rect 8739 1942 8771 1974
rect 8771 1942 8775 1974
rect 8735 1906 8775 1942
rect 8735 1874 8739 1906
rect 8739 1874 8771 1906
rect 8771 1874 8775 1906
rect 8735 1838 8775 1874
rect 8735 1806 8739 1838
rect 8739 1806 8771 1838
rect 8771 1806 8775 1838
rect 8735 1770 8775 1806
rect 8735 1738 8739 1770
rect 8739 1738 8771 1770
rect 8771 1738 8775 1770
rect 8735 1702 8775 1738
rect 8735 1670 8739 1702
rect 8739 1670 8771 1702
rect 8771 1670 8775 1702
rect 8735 1634 8775 1670
rect 8735 1602 8739 1634
rect 8739 1602 8771 1634
rect 8771 1602 8775 1634
rect 8735 1566 8775 1602
rect 8735 1534 8739 1566
rect 8739 1534 8771 1566
rect 8771 1534 8775 1566
rect 8735 1528 8775 1534
rect 8392 1414 8514 1420
rect 8392 1382 8437 1414
rect 8437 1382 8469 1414
rect 8469 1382 8514 1414
rect 8392 1346 8514 1382
rect 8392 1314 8437 1346
rect 8437 1314 8469 1346
rect 8469 1314 8514 1346
rect 8392 1278 8514 1314
rect 8392 1246 8437 1278
rect 8437 1246 8469 1278
rect 8469 1246 8514 1278
rect 8392 1210 8514 1246
rect 8392 1178 8437 1210
rect 8437 1178 8469 1210
rect 8469 1178 8514 1210
rect 8392 1142 8514 1178
rect 8392 1110 8437 1142
rect 8437 1110 8469 1142
rect 8469 1110 8514 1142
rect 8392 1074 8514 1110
rect 8392 1042 8437 1074
rect 8437 1042 8469 1074
rect 8469 1042 8514 1074
rect 8392 1006 8514 1042
rect 8392 974 8437 1006
rect 8437 974 8469 1006
rect 8469 974 8514 1006
rect 8392 938 8514 974
rect 8392 906 8437 938
rect 8437 906 8469 938
rect 8469 906 8514 938
rect 8392 870 8514 906
rect 8392 838 8437 870
rect 8437 838 8469 870
rect 8469 838 8514 870
rect 8392 802 8514 838
rect 8392 770 8437 802
rect 8437 770 8469 802
rect 8469 770 8514 802
rect 8392 734 8514 770
rect 8392 702 8437 734
rect 8437 702 8469 734
rect 8469 702 8514 734
rect 8392 666 8514 702
rect 8392 634 8437 666
rect 8437 634 8469 666
rect 8469 634 8514 666
rect 8392 598 8514 634
rect 8392 566 8437 598
rect 8437 566 8469 598
rect 8469 566 8514 598
rect 8392 560 8514 566
rect 9600 4318 9722 4324
rect 9600 4286 9645 4318
rect 9645 4286 9677 4318
rect 9677 4286 9722 4318
rect 9600 4250 9722 4286
rect 9600 4218 9645 4250
rect 9645 4218 9677 4250
rect 9677 4218 9722 4250
rect 9600 4182 9722 4218
rect 9600 4150 9645 4182
rect 9645 4150 9677 4182
rect 9677 4150 9722 4182
rect 9600 4114 9722 4150
rect 9600 4082 9645 4114
rect 9645 4082 9677 4114
rect 9677 4082 9722 4114
rect 9600 4046 9722 4082
rect 9600 4014 9645 4046
rect 9645 4014 9677 4046
rect 9677 4014 9722 4046
rect 9600 3978 9722 4014
rect 9600 3946 9645 3978
rect 9645 3946 9677 3978
rect 9677 3946 9722 3978
rect 9600 3910 9722 3946
rect 9600 3878 9645 3910
rect 9645 3878 9677 3910
rect 9677 3878 9722 3910
rect 9600 3842 9722 3878
rect 9600 3810 9645 3842
rect 9645 3810 9677 3842
rect 9677 3810 9722 3842
rect 9600 3774 9722 3810
rect 9600 3742 9645 3774
rect 9645 3742 9677 3774
rect 9677 3742 9722 3774
rect 9600 3706 9722 3742
rect 9600 3674 9645 3706
rect 9645 3674 9677 3706
rect 9677 3674 9722 3706
rect 9600 3638 9722 3674
rect 9600 3606 9645 3638
rect 9645 3606 9677 3638
rect 9677 3606 9722 3638
rect 9600 3570 9722 3606
rect 9600 3538 9645 3570
rect 9645 3538 9677 3570
rect 9677 3538 9722 3570
rect 9600 3502 9722 3538
rect 9600 3470 9645 3502
rect 9645 3470 9677 3502
rect 9677 3470 9722 3502
rect 9600 3464 9722 3470
rect 9339 3350 9379 3356
rect 9339 3318 9343 3350
rect 9343 3318 9375 3350
rect 9375 3318 9379 3350
rect 9339 3282 9379 3318
rect 9339 3250 9343 3282
rect 9343 3250 9375 3282
rect 9375 3250 9379 3282
rect 9339 3214 9379 3250
rect 9339 3182 9343 3214
rect 9343 3182 9375 3214
rect 9375 3182 9379 3214
rect 9339 3146 9379 3182
rect 9339 3114 9343 3146
rect 9343 3114 9375 3146
rect 9375 3114 9379 3146
rect 9339 3078 9379 3114
rect 9339 3046 9343 3078
rect 9343 3046 9375 3078
rect 9375 3046 9379 3078
rect 9339 3010 9379 3046
rect 9339 2978 9343 3010
rect 9343 2978 9375 3010
rect 9375 2978 9379 3010
rect 9339 2942 9379 2978
rect 9339 2910 9343 2942
rect 9343 2910 9375 2942
rect 9375 2910 9379 2942
rect 9339 2874 9379 2910
rect 9339 2842 9343 2874
rect 9343 2842 9375 2874
rect 9375 2842 9379 2874
rect 9339 2806 9379 2842
rect 9339 2774 9343 2806
rect 9343 2774 9375 2806
rect 9375 2774 9379 2806
rect 9339 2738 9379 2774
rect 9339 2706 9343 2738
rect 9343 2706 9375 2738
rect 9375 2706 9379 2738
rect 9339 2670 9379 2706
rect 9339 2638 9343 2670
rect 9343 2638 9375 2670
rect 9375 2638 9379 2670
rect 9339 2602 9379 2638
rect 9339 2570 9343 2602
rect 9343 2570 9375 2602
rect 9375 2570 9379 2602
rect 9339 2534 9379 2570
rect 9339 2502 9343 2534
rect 9343 2502 9375 2534
rect 9375 2502 9379 2534
rect 9339 2496 9379 2502
rect 8996 2382 9118 2388
rect 8996 2350 9041 2382
rect 9041 2350 9073 2382
rect 9073 2350 9118 2382
rect 8996 2314 9118 2350
rect 8996 2282 9041 2314
rect 9041 2282 9073 2314
rect 9073 2282 9118 2314
rect 8996 2246 9118 2282
rect 8996 2214 9041 2246
rect 9041 2214 9073 2246
rect 9073 2214 9118 2246
rect 8996 2178 9118 2214
rect 8996 2146 9041 2178
rect 9041 2146 9073 2178
rect 9073 2146 9118 2178
rect 8996 2110 9118 2146
rect 8996 2078 9041 2110
rect 9041 2078 9073 2110
rect 9073 2078 9118 2110
rect 8996 2042 9118 2078
rect 8996 2010 9041 2042
rect 9041 2010 9073 2042
rect 9073 2010 9118 2042
rect 8996 1974 9118 2010
rect 8996 1942 9041 1974
rect 9041 1942 9073 1974
rect 9073 1942 9118 1974
rect 8996 1906 9118 1942
rect 8996 1874 9041 1906
rect 9041 1874 9073 1906
rect 9073 1874 9118 1906
rect 8996 1838 9118 1874
rect 8996 1806 9041 1838
rect 9041 1806 9073 1838
rect 9073 1806 9118 1838
rect 8996 1770 9118 1806
rect 8996 1738 9041 1770
rect 9041 1738 9073 1770
rect 9073 1738 9118 1770
rect 8996 1702 9118 1738
rect 8996 1670 9041 1702
rect 9041 1670 9073 1702
rect 9073 1670 9118 1702
rect 8996 1634 9118 1670
rect 8996 1602 9041 1634
rect 9041 1602 9073 1634
rect 9073 1602 9118 1634
rect 8996 1566 9118 1602
rect 8996 1534 9041 1566
rect 9041 1534 9073 1566
rect 9073 1534 9118 1566
rect 8996 1528 9118 1534
rect 8735 1414 8775 1420
rect 8735 1382 8739 1414
rect 8739 1382 8771 1414
rect 8771 1382 8775 1414
rect 8735 1346 8775 1382
rect 8735 1314 8739 1346
rect 8739 1314 8771 1346
rect 8771 1314 8775 1346
rect 8735 1278 8775 1314
rect 8735 1246 8739 1278
rect 8739 1246 8771 1278
rect 8771 1246 8775 1278
rect 8735 1210 8775 1246
rect 8735 1178 8739 1210
rect 8739 1178 8771 1210
rect 8771 1178 8775 1210
rect 8735 1142 8775 1178
rect 8735 1110 8739 1142
rect 8739 1110 8771 1142
rect 8771 1110 8775 1142
rect 8735 1074 8775 1110
rect 8735 1042 8739 1074
rect 8739 1042 8771 1074
rect 8771 1042 8775 1074
rect 8735 1006 8775 1042
rect 8735 974 8739 1006
rect 8739 974 8771 1006
rect 8771 974 8775 1006
rect 8735 938 8775 974
rect 8735 906 8739 938
rect 8739 906 8771 938
rect 8771 906 8775 938
rect 8735 870 8775 906
rect 8735 838 8739 870
rect 8739 838 8771 870
rect 8771 838 8775 870
rect 8735 802 8775 838
rect 8735 770 8739 802
rect 8739 770 8771 802
rect 8771 770 8775 802
rect 8735 734 8775 770
rect 8735 702 8739 734
rect 8739 702 8771 734
rect 8771 702 8775 734
rect 8735 666 8775 702
rect 8735 634 8739 666
rect 8739 634 8771 666
rect 8771 634 8775 666
rect 8735 598 8775 634
rect 8735 566 8739 598
rect 8739 566 8771 598
rect 8771 566 8775 598
rect 8735 560 8775 566
rect 9943 4318 9983 4324
rect 9943 4286 9947 4318
rect 9947 4286 9979 4318
rect 9979 4286 9983 4318
rect 9943 4250 9983 4286
rect 9943 4218 9947 4250
rect 9947 4218 9979 4250
rect 9979 4218 9983 4250
rect 9943 4182 9983 4218
rect 9943 4150 9947 4182
rect 9947 4150 9979 4182
rect 9979 4150 9983 4182
rect 9943 4114 9983 4150
rect 9943 4082 9947 4114
rect 9947 4082 9979 4114
rect 9979 4082 9983 4114
rect 9943 4046 9983 4082
rect 9943 4014 9947 4046
rect 9947 4014 9979 4046
rect 9979 4014 9983 4046
rect 9943 3978 9983 4014
rect 9943 3946 9947 3978
rect 9947 3946 9979 3978
rect 9979 3946 9983 3978
rect 9943 3910 9983 3946
rect 9943 3878 9947 3910
rect 9947 3878 9979 3910
rect 9979 3878 9983 3910
rect 9943 3842 9983 3878
rect 9943 3810 9947 3842
rect 9947 3810 9979 3842
rect 9979 3810 9983 3842
rect 9943 3774 9983 3810
rect 9943 3742 9947 3774
rect 9947 3742 9979 3774
rect 9979 3742 9983 3774
rect 9943 3706 9983 3742
rect 9943 3674 9947 3706
rect 9947 3674 9979 3706
rect 9979 3674 9983 3706
rect 9943 3638 9983 3674
rect 9943 3606 9947 3638
rect 9947 3606 9979 3638
rect 9979 3606 9983 3638
rect 9943 3570 9983 3606
rect 9943 3538 9947 3570
rect 9947 3538 9979 3570
rect 9979 3538 9983 3570
rect 9943 3502 9983 3538
rect 9943 3470 9947 3502
rect 9947 3470 9979 3502
rect 9979 3470 9983 3502
rect 9943 3464 9983 3470
rect 9600 3350 9722 3356
rect 9600 3318 9645 3350
rect 9645 3318 9677 3350
rect 9677 3318 9722 3350
rect 9600 3282 9722 3318
rect 9600 3250 9645 3282
rect 9645 3250 9677 3282
rect 9677 3250 9722 3282
rect 9600 3214 9722 3250
rect 9600 3182 9645 3214
rect 9645 3182 9677 3214
rect 9677 3182 9722 3214
rect 9600 3146 9722 3182
rect 9600 3114 9645 3146
rect 9645 3114 9677 3146
rect 9677 3114 9722 3146
rect 9600 3078 9722 3114
rect 9600 3046 9645 3078
rect 9645 3046 9677 3078
rect 9677 3046 9722 3078
rect 9600 3010 9722 3046
rect 9600 2978 9645 3010
rect 9645 2978 9677 3010
rect 9677 2978 9722 3010
rect 9600 2942 9722 2978
rect 9600 2910 9645 2942
rect 9645 2910 9677 2942
rect 9677 2910 9722 2942
rect 9600 2874 9722 2910
rect 9600 2842 9645 2874
rect 9645 2842 9677 2874
rect 9677 2842 9722 2874
rect 9600 2806 9722 2842
rect 9600 2774 9645 2806
rect 9645 2774 9677 2806
rect 9677 2774 9722 2806
rect 9600 2738 9722 2774
rect 9600 2706 9645 2738
rect 9645 2706 9677 2738
rect 9677 2706 9722 2738
rect 9600 2670 9722 2706
rect 9600 2638 9645 2670
rect 9645 2638 9677 2670
rect 9677 2638 9722 2670
rect 9600 2602 9722 2638
rect 9600 2570 9645 2602
rect 9645 2570 9677 2602
rect 9677 2570 9722 2602
rect 9600 2534 9722 2570
rect 9600 2502 9645 2534
rect 9645 2502 9677 2534
rect 9677 2502 9722 2534
rect 9600 2496 9722 2502
rect 9339 2382 9379 2388
rect 9339 2350 9343 2382
rect 9343 2350 9375 2382
rect 9375 2350 9379 2382
rect 9339 2314 9379 2350
rect 9339 2282 9343 2314
rect 9343 2282 9375 2314
rect 9375 2282 9379 2314
rect 9339 2246 9379 2282
rect 9339 2214 9343 2246
rect 9343 2214 9375 2246
rect 9375 2214 9379 2246
rect 9339 2178 9379 2214
rect 9339 2146 9343 2178
rect 9343 2146 9375 2178
rect 9375 2146 9379 2178
rect 9339 2110 9379 2146
rect 9339 2078 9343 2110
rect 9343 2078 9375 2110
rect 9375 2078 9379 2110
rect 9339 2042 9379 2078
rect 9339 2010 9343 2042
rect 9343 2010 9375 2042
rect 9375 2010 9379 2042
rect 9339 1974 9379 2010
rect 9339 1942 9343 1974
rect 9343 1942 9375 1974
rect 9375 1942 9379 1974
rect 9339 1906 9379 1942
rect 9339 1874 9343 1906
rect 9343 1874 9375 1906
rect 9375 1874 9379 1906
rect 9339 1838 9379 1874
rect 9339 1806 9343 1838
rect 9343 1806 9375 1838
rect 9375 1806 9379 1838
rect 9339 1770 9379 1806
rect 9339 1738 9343 1770
rect 9343 1738 9375 1770
rect 9375 1738 9379 1770
rect 9339 1702 9379 1738
rect 9339 1670 9343 1702
rect 9343 1670 9375 1702
rect 9375 1670 9379 1702
rect 9339 1634 9379 1670
rect 9339 1602 9343 1634
rect 9343 1602 9375 1634
rect 9375 1602 9379 1634
rect 9339 1566 9379 1602
rect 9339 1534 9343 1566
rect 9343 1534 9375 1566
rect 9375 1534 9379 1566
rect 9339 1528 9379 1534
rect 8996 1414 9118 1420
rect 8996 1382 9041 1414
rect 9041 1382 9073 1414
rect 9073 1382 9118 1414
rect 8996 1346 9118 1382
rect 8996 1314 9041 1346
rect 9041 1314 9073 1346
rect 9073 1314 9118 1346
rect 8996 1278 9118 1314
rect 8996 1246 9041 1278
rect 9041 1246 9073 1278
rect 9073 1246 9118 1278
rect 8996 1210 9118 1246
rect 8996 1178 9041 1210
rect 9041 1178 9073 1210
rect 9073 1178 9118 1210
rect 8996 1142 9118 1178
rect 8996 1110 9041 1142
rect 9041 1110 9073 1142
rect 9073 1110 9118 1142
rect 8996 1074 9118 1110
rect 8996 1042 9041 1074
rect 9041 1042 9073 1074
rect 9073 1042 9118 1074
rect 8996 1006 9118 1042
rect 8996 974 9041 1006
rect 9041 974 9073 1006
rect 9073 974 9118 1006
rect 8996 938 9118 974
rect 8996 906 9041 938
rect 9041 906 9073 938
rect 9073 906 9118 938
rect 8996 870 9118 906
rect 8996 838 9041 870
rect 9041 838 9073 870
rect 9073 838 9118 870
rect 8996 802 9118 838
rect 8996 770 9041 802
rect 9041 770 9073 802
rect 9073 770 9118 802
rect 8996 734 9118 770
rect 8996 702 9041 734
rect 9041 702 9073 734
rect 9073 702 9118 734
rect 8996 666 9118 702
rect 8996 634 9041 666
rect 9041 634 9073 666
rect 9073 634 9118 666
rect 8996 598 9118 634
rect 8996 566 9041 598
rect 9041 566 9073 598
rect 9073 566 9118 598
rect 8996 560 9118 566
rect 10204 4318 10326 4324
rect 10204 4286 10249 4318
rect 10249 4286 10281 4318
rect 10281 4286 10326 4318
rect 10204 4250 10326 4286
rect 10204 4218 10249 4250
rect 10249 4218 10281 4250
rect 10281 4218 10326 4250
rect 10204 4182 10326 4218
rect 10204 4150 10249 4182
rect 10249 4150 10281 4182
rect 10281 4150 10326 4182
rect 10204 4114 10326 4150
rect 10204 4082 10249 4114
rect 10249 4082 10281 4114
rect 10281 4082 10326 4114
rect 10204 4046 10326 4082
rect 10204 4014 10249 4046
rect 10249 4014 10281 4046
rect 10281 4014 10326 4046
rect 10204 3978 10326 4014
rect 10204 3946 10249 3978
rect 10249 3946 10281 3978
rect 10281 3946 10326 3978
rect 10204 3910 10326 3946
rect 10204 3878 10249 3910
rect 10249 3878 10281 3910
rect 10281 3878 10326 3910
rect 10204 3842 10326 3878
rect 10204 3810 10249 3842
rect 10249 3810 10281 3842
rect 10281 3810 10326 3842
rect 10204 3774 10326 3810
rect 10204 3742 10249 3774
rect 10249 3742 10281 3774
rect 10281 3742 10326 3774
rect 10204 3706 10326 3742
rect 10204 3674 10249 3706
rect 10249 3674 10281 3706
rect 10281 3674 10326 3706
rect 10204 3638 10326 3674
rect 10204 3606 10249 3638
rect 10249 3606 10281 3638
rect 10281 3606 10326 3638
rect 10204 3570 10326 3606
rect 10204 3538 10249 3570
rect 10249 3538 10281 3570
rect 10281 3538 10326 3570
rect 10204 3502 10326 3538
rect 10204 3470 10249 3502
rect 10249 3470 10281 3502
rect 10281 3470 10326 3502
rect 10204 3464 10326 3470
rect 9943 3350 9983 3356
rect 9943 3318 9947 3350
rect 9947 3318 9979 3350
rect 9979 3318 9983 3350
rect 9943 3282 9983 3318
rect 9943 3250 9947 3282
rect 9947 3250 9979 3282
rect 9979 3250 9983 3282
rect 9943 3214 9983 3250
rect 9943 3182 9947 3214
rect 9947 3182 9979 3214
rect 9979 3182 9983 3214
rect 9943 3146 9983 3182
rect 9943 3114 9947 3146
rect 9947 3114 9979 3146
rect 9979 3114 9983 3146
rect 9943 3078 9983 3114
rect 9943 3046 9947 3078
rect 9947 3046 9979 3078
rect 9979 3046 9983 3078
rect 9943 3010 9983 3046
rect 9943 2978 9947 3010
rect 9947 2978 9979 3010
rect 9979 2978 9983 3010
rect 9943 2942 9983 2978
rect 9943 2910 9947 2942
rect 9947 2910 9979 2942
rect 9979 2910 9983 2942
rect 9943 2874 9983 2910
rect 9943 2842 9947 2874
rect 9947 2842 9979 2874
rect 9979 2842 9983 2874
rect 9943 2806 9983 2842
rect 9943 2774 9947 2806
rect 9947 2774 9979 2806
rect 9979 2774 9983 2806
rect 9943 2738 9983 2774
rect 9943 2706 9947 2738
rect 9947 2706 9979 2738
rect 9979 2706 9983 2738
rect 9943 2670 9983 2706
rect 9943 2638 9947 2670
rect 9947 2638 9979 2670
rect 9979 2638 9983 2670
rect 9943 2602 9983 2638
rect 9943 2570 9947 2602
rect 9947 2570 9979 2602
rect 9979 2570 9983 2602
rect 9943 2534 9983 2570
rect 9943 2502 9947 2534
rect 9947 2502 9979 2534
rect 9979 2502 9983 2534
rect 9943 2496 9983 2502
rect 9600 2382 9722 2388
rect 9600 2350 9645 2382
rect 9645 2350 9677 2382
rect 9677 2350 9722 2382
rect 9600 2314 9722 2350
rect 9600 2282 9645 2314
rect 9645 2282 9677 2314
rect 9677 2282 9722 2314
rect 9600 2246 9722 2282
rect 9600 2214 9645 2246
rect 9645 2214 9677 2246
rect 9677 2214 9722 2246
rect 9600 2178 9722 2214
rect 9600 2146 9645 2178
rect 9645 2146 9677 2178
rect 9677 2146 9722 2178
rect 9600 2110 9722 2146
rect 9600 2078 9645 2110
rect 9645 2078 9677 2110
rect 9677 2078 9722 2110
rect 9600 2042 9722 2078
rect 9600 2010 9645 2042
rect 9645 2010 9677 2042
rect 9677 2010 9722 2042
rect 9600 1974 9722 2010
rect 9600 1942 9645 1974
rect 9645 1942 9677 1974
rect 9677 1942 9722 1974
rect 9600 1906 9722 1942
rect 9600 1874 9645 1906
rect 9645 1874 9677 1906
rect 9677 1874 9722 1906
rect 9600 1838 9722 1874
rect 9600 1806 9645 1838
rect 9645 1806 9677 1838
rect 9677 1806 9722 1838
rect 9600 1770 9722 1806
rect 9600 1738 9645 1770
rect 9645 1738 9677 1770
rect 9677 1738 9722 1770
rect 9600 1702 9722 1738
rect 9600 1670 9645 1702
rect 9645 1670 9677 1702
rect 9677 1670 9722 1702
rect 9600 1634 9722 1670
rect 9600 1602 9645 1634
rect 9645 1602 9677 1634
rect 9677 1602 9722 1634
rect 9600 1566 9722 1602
rect 9600 1534 9645 1566
rect 9645 1534 9677 1566
rect 9677 1534 9722 1566
rect 9600 1528 9722 1534
rect 9339 1414 9379 1420
rect 9339 1382 9343 1414
rect 9343 1382 9375 1414
rect 9375 1382 9379 1414
rect 9339 1346 9379 1382
rect 9339 1314 9343 1346
rect 9343 1314 9375 1346
rect 9375 1314 9379 1346
rect 9339 1278 9379 1314
rect 9339 1246 9343 1278
rect 9343 1246 9375 1278
rect 9375 1246 9379 1278
rect 9339 1210 9379 1246
rect 9339 1178 9343 1210
rect 9343 1178 9375 1210
rect 9375 1178 9379 1210
rect 9339 1142 9379 1178
rect 9339 1110 9343 1142
rect 9343 1110 9375 1142
rect 9375 1110 9379 1142
rect 9339 1074 9379 1110
rect 9339 1042 9343 1074
rect 9343 1042 9375 1074
rect 9375 1042 9379 1074
rect 9339 1006 9379 1042
rect 9339 974 9343 1006
rect 9343 974 9375 1006
rect 9375 974 9379 1006
rect 9339 938 9379 974
rect 9339 906 9343 938
rect 9343 906 9375 938
rect 9375 906 9379 938
rect 9339 870 9379 906
rect 9339 838 9343 870
rect 9343 838 9375 870
rect 9375 838 9379 870
rect 9339 802 9379 838
rect 9339 770 9343 802
rect 9343 770 9375 802
rect 9375 770 9379 802
rect 9339 734 9379 770
rect 9339 702 9343 734
rect 9343 702 9375 734
rect 9375 702 9379 734
rect 9339 666 9379 702
rect 9339 634 9343 666
rect 9343 634 9375 666
rect 9375 634 9379 666
rect 9339 598 9379 634
rect 9339 566 9343 598
rect 9343 566 9375 598
rect 9375 566 9379 598
rect 9339 560 9379 566
rect 10547 4318 10587 4324
rect 10547 4286 10551 4318
rect 10551 4286 10583 4318
rect 10583 4286 10587 4318
rect 10547 4250 10587 4286
rect 10547 4218 10551 4250
rect 10551 4218 10583 4250
rect 10583 4218 10587 4250
rect 10547 4182 10587 4218
rect 10547 4150 10551 4182
rect 10551 4150 10583 4182
rect 10583 4150 10587 4182
rect 10547 4114 10587 4150
rect 10547 4082 10551 4114
rect 10551 4082 10583 4114
rect 10583 4082 10587 4114
rect 10547 4046 10587 4082
rect 10547 4014 10551 4046
rect 10551 4014 10583 4046
rect 10583 4014 10587 4046
rect 10547 3978 10587 4014
rect 10547 3946 10551 3978
rect 10551 3946 10583 3978
rect 10583 3946 10587 3978
rect 10547 3910 10587 3946
rect 10547 3878 10551 3910
rect 10551 3878 10583 3910
rect 10583 3878 10587 3910
rect 10547 3842 10587 3878
rect 10547 3810 10551 3842
rect 10551 3810 10583 3842
rect 10583 3810 10587 3842
rect 10547 3774 10587 3810
rect 10547 3742 10551 3774
rect 10551 3742 10583 3774
rect 10583 3742 10587 3774
rect 10547 3706 10587 3742
rect 10547 3674 10551 3706
rect 10551 3674 10583 3706
rect 10583 3674 10587 3706
rect 10547 3638 10587 3674
rect 10547 3606 10551 3638
rect 10551 3606 10583 3638
rect 10583 3606 10587 3638
rect 10547 3570 10587 3606
rect 10547 3538 10551 3570
rect 10551 3538 10583 3570
rect 10583 3538 10587 3570
rect 10547 3502 10587 3538
rect 10547 3470 10551 3502
rect 10551 3470 10583 3502
rect 10583 3470 10587 3502
rect 10547 3464 10587 3470
rect 10204 3350 10326 3356
rect 10204 3318 10249 3350
rect 10249 3318 10281 3350
rect 10281 3318 10326 3350
rect 10204 3282 10326 3318
rect 10204 3250 10249 3282
rect 10249 3250 10281 3282
rect 10281 3250 10326 3282
rect 10204 3214 10326 3250
rect 10204 3182 10249 3214
rect 10249 3182 10281 3214
rect 10281 3182 10326 3214
rect 10204 3146 10326 3182
rect 10204 3114 10249 3146
rect 10249 3114 10281 3146
rect 10281 3114 10326 3146
rect 10204 3078 10326 3114
rect 10204 3046 10249 3078
rect 10249 3046 10281 3078
rect 10281 3046 10326 3078
rect 10204 3010 10326 3046
rect 10204 2978 10249 3010
rect 10249 2978 10281 3010
rect 10281 2978 10326 3010
rect 10204 2942 10326 2978
rect 10204 2910 10249 2942
rect 10249 2910 10281 2942
rect 10281 2910 10326 2942
rect 10204 2874 10326 2910
rect 10204 2842 10249 2874
rect 10249 2842 10281 2874
rect 10281 2842 10326 2874
rect 10204 2806 10326 2842
rect 10204 2774 10249 2806
rect 10249 2774 10281 2806
rect 10281 2774 10326 2806
rect 10204 2738 10326 2774
rect 10204 2706 10249 2738
rect 10249 2706 10281 2738
rect 10281 2706 10326 2738
rect 10204 2670 10326 2706
rect 10204 2638 10249 2670
rect 10249 2638 10281 2670
rect 10281 2638 10326 2670
rect 10204 2602 10326 2638
rect 10204 2570 10249 2602
rect 10249 2570 10281 2602
rect 10281 2570 10326 2602
rect 10204 2534 10326 2570
rect 10204 2502 10249 2534
rect 10249 2502 10281 2534
rect 10281 2502 10326 2534
rect 10204 2496 10326 2502
rect 9943 2382 9983 2388
rect 9943 2350 9947 2382
rect 9947 2350 9979 2382
rect 9979 2350 9983 2382
rect 9943 2314 9983 2350
rect 9943 2282 9947 2314
rect 9947 2282 9979 2314
rect 9979 2282 9983 2314
rect 9943 2246 9983 2282
rect 9943 2214 9947 2246
rect 9947 2214 9979 2246
rect 9979 2214 9983 2246
rect 9943 2178 9983 2214
rect 9943 2146 9947 2178
rect 9947 2146 9979 2178
rect 9979 2146 9983 2178
rect 9943 2110 9983 2146
rect 9943 2078 9947 2110
rect 9947 2078 9979 2110
rect 9979 2078 9983 2110
rect 9943 2042 9983 2078
rect 9943 2010 9947 2042
rect 9947 2010 9979 2042
rect 9979 2010 9983 2042
rect 9943 1974 9983 2010
rect 9943 1942 9947 1974
rect 9947 1942 9979 1974
rect 9979 1942 9983 1974
rect 9943 1906 9983 1942
rect 9943 1874 9947 1906
rect 9947 1874 9979 1906
rect 9979 1874 9983 1906
rect 9943 1838 9983 1874
rect 9943 1806 9947 1838
rect 9947 1806 9979 1838
rect 9979 1806 9983 1838
rect 9943 1770 9983 1806
rect 9943 1738 9947 1770
rect 9947 1738 9979 1770
rect 9979 1738 9983 1770
rect 9943 1702 9983 1738
rect 9943 1670 9947 1702
rect 9947 1670 9979 1702
rect 9979 1670 9983 1702
rect 9943 1634 9983 1670
rect 9943 1602 9947 1634
rect 9947 1602 9979 1634
rect 9979 1602 9983 1634
rect 9943 1566 9983 1602
rect 9943 1534 9947 1566
rect 9947 1534 9979 1566
rect 9979 1534 9983 1566
rect 9943 1528 9983 1534
rect 9600 1414 9722 1420
rect 9600 1382 9645 1414
rect 9645 1382 9677 1414
rect 9677 1382 9722 1414
rect 9600 1346 9722 1382
rect 9600 1314 9645 1346
rect 9645 1314 9677 1346
rect 9677 1314 9722 1346
rect 9600 1278 9722 1314
rect 9600 1246 9645 1278
rect 9645 1246 9677 1278
rect 9677 1246 9722 1278
rect 9600 1210 9722 1246
rect 9600 1178 9645 1210
rect 9645 1178 9677 1210
rect 9677 1178 9722 1210
rect 9600 1142 9722 1178
rect 9600 1110 9645 1142
rect 9645 1110 9677 1142
rect 9677 1110 9722 1142
rect 9600 1074 9722 1110
rect 9600 1042 9645 1074
rect 9645 1042 9677 1074
rect 9677 1042 9722 1074
rect 9600 1006 9722 1042
rect 9600 974 9645 1006
rect 9645 974 9677 1006
rect 9677 974 9722 1006
rect 9600 938 9722 974
rect 9600 906 9645 938
rect 9645 906 9677 938
rect 9677 906 9722 938
rect 9600 870 9722 906
rect 9600 838 9645 870
rect 9645 838 9677 870
rect 9677 838 9722 870
rect 9600 802 9722 838
rect 9600 770 9645 802
rect 9645 770 9677 802
rect 9677 770 9722 802
rect 9600 734 9722 770
rect 9600 702 9645 734
rect 9645 702 9677 734
rect 9677 702 9722 734
rect 9600 666 9722 702
rect 9600 634 9645 666
rect 9645 634 9677 666
rect 9677 634 9722 666
rect 9600 598 9722 634
rect 9600 566 9645 598
rect 9645 566 9677 598
rect 9677 566 9722 598
rect 9600 560 9722 566
rect 10808 4318 10930 4324
rect 10808 4286 10853 4318
rect 10853 4286 10885 4318
rect 10885 4286 10930 4318
rect 10808 4250 10930 4286
rect 10808 4218 10853 4250
rect 10853 4218 10885 4250
rect 10885 4218 10930 4250
rect 10808 4182 10930 4218
rect 10808 4150 10853 4182
rect 10853 4150 10885 4182
rect 10885 4150 10930 4182
rect 10808 4114 10930 4150
rect 10808 4082 10853 4114
rect 10853 4082 10885 4114
rect 10885 4082 10930 4114
rect 10808 4046 10930 4082
rect 10808 4014 10853 4046
rect 10853 4014 10885 4046
rect 10885 4014 10930 4046
rect 10808 3978 10930 4014
rect 10808 3946 10853 3978
rect 10853 3946 10885 3978
rect 10885 3946 10930 3978
rect 10808 3910 10930 3946
rect 10808 3878 10853 3910
rect 10853 3878 10885 3910
rect 10885 3878 10930 3910
rect 10808 3842 10930 3878
rect 10808 3810 10853 3842
rect 10853 3810 10885 3842
rect 10885 3810 10930 3842
rect 10808 3774 10930 3810
rect 10808 3742 10853 3774
rect 10853 3742 10885 3774
rect 10885 3742 10930 3774
rect 10808 3706 10930 3742
rect 10808 3674 10853 3706
rect 10853 3674 10885 3706
rect 10885 3674 10930 3706
rect 10808 3638 10930 3674
rect 10808 3606 10853 3638
rect 10853 3606 10885 3638
rect 10885 3606 10930 3638
rect 10808 3570 10930 3606
rect 10808 3538 10853 3570
rect 10853 3538 10885 3570
rect 10885 3538 10930 3570
rect 10808 3502 10930 3538
rect 10808 3470 10853 3502
rect 10853 3470 10885 3502
rect 10885 3470 10930 3502
rect 10808 3464 10930 3470
rect 10547 3350 10587 3356
rect 10547 3318 10551 3350
rect 10551 3318 10583 3350
rect 10583 3318 10587 3350
rect 10547 3282 10587 3318
rect 10547 3250 10551 3282
rect 10551 3250 10583 3282
rect 10583 3250 10587 3282
rect 10547 3214 10587 3250
rect 10547 3182 10551 3214
rect 10551 3182 10583 3214
rect 10583 3182 10587 3214
rect 10547 3146 10587 3182
rect 10547 3114 10551 3146
rect 10551 3114 10583 3146
rect 10583 3114 10587 3146
rect 10547 3078 10587 3114
rect 10547 3046 10551 3078
rect 10551 3046 10583 3078
rect 10583 3046 10587 3078
rect 10547 3010 10587 3046
rect 10547 2978 10551 3010
rect 10551 2978 10583 3010
rect 10583 2978 10587 3010
rect 10547 2942 10587 2978
rect 10547 2910 10551 2942
rect 10551 2910 10583 2942
rect 10583 2910 10587 2942
rect 10547 2874 10587 2910
rect 10547 2842 10551 2874
rect 10551 2842 10583 2874
rect 10583 2842 10587 2874
rect 10547 2806 10587 2842
rect 10547 2774 10551 2806
rect 10551 2774 10583 2806
rect 10583 2774 10587 2806
rect 10547 2738 10587 2774
rect 10547 2706 10551 2738
rect 10551 2706 10583 2738
rect 10583 2706 10587 2738
rect 10547 2670 10587 2706
rect 10547 2638 10551 2670
rect 10551 2638 10583 2670
rect 10583 2638 10587 2670
rect 10547 2602 10587 2638
rect 10547 2570 10551 2602
rect 10551 2570 10583 2602
rect 10583 2570 10587 2602
rect 10547 2534 10587 2570
rect 10547 2502 10551 2534
rect 10551 2502 10583 2534
rect 10583 2502 10587 2534
rect 10547 2496 10587 2502
rect 10204 2382 10326 2388
rect 10204 2350 10249 2382
rect 10249 2350 10281 2382
rect 10281 2350 10326 2382
rect 10204 2314 10326 2350
rect 10204 2282 10249 2314
rect 10249 2282 10281 2314
rect 10281 2282 10326 2314
rect 10204 2246 10326 2282
rect 10204 2214 10249 2246
rect 10249 2214 10281 2246
rect 10281 2214 10326 2246
rect 10204 2178 10326 2214
rect 10204 2146 10249 2178
rect 10249 2146 10281 2178
rect 10281 2146 10326 2178
rect 10204 2110 10326 2146
rect 10204 2078 10249 2110
rect 10249 2078 10281 2110
rect 10281 2078 10326 2110
rect 10204 2042 10326 2078
rect 10204 2010 10249 2042
rect 10249 2010 10281 2042
rect 10281 2010 10326 2042
rect 10204 1974 10326 2010
rect 10204 1942 10249 1974
rect 10249 1942 10281 1974
rect 10281 1942 10326 1974
rect 10204 1906 10326 1942
rect 10204 1874 10249 1906
rect 10249 1874 10281 1906
rect 10281 1874 10326 1906
rect 10204 1838 10326 1874
rect 10204 1806 10249 1838
rect 10249 1806 10281 1838
rect 10281 1806 10326 1838
rect 10204 1770 10326 1806
rect 10204 1738 10249 1770
rect 10249 1738 10281 1770
rect 10281 1738 10326 1770
rect 10204 1702 10326 1738
rect 10204 1670 10249 1702
rect 10249 1670 10281 1702
rect 10281 1670 10326 1702
rect 10204 1634 10326 1670
rect 10204 1602 10249 1634
rect 10249 1602 10281 1634
rect 10281 1602 10326 1634
rect 10204 1566 10326 1602
rect 10204 1534 10249 1566
rect 10249 1534 10281 1566
rect 10281 1534 10326 1566
rect 10204 1528 10326 1534
rect 9943 1414 9983 1420
rect 9943 1382 9947 1414
rect 9947 1382 9979 1414
rect 9979 1382 9983 1414
rect 9943 1346 9983 1382
rect 9943 1314 9947 1346
rect 9947 1314 9979 1346
rect 9979 1314 9983 1346
rect 9943 1278 9983 1314
rect 9943 1246 9947 1278
rect 9947 1246 9979 1278
rect 9979 1246 9983 1278
rect 9943 1210 9983 1246
rect 9943 1178 9947 1210
rect 9947 1178 9979 1210
rect 9979 1178 9983 1210
rect 9943 1142 9983 1178
rect 9943 1110 9947 1142
rect 9947 1110 9979 1142
rect 9979 1110 9983 1142
rect 9943 1074 9983 1110
rect 9943 1042 9947 1074
rect 9947 1042 9979 1074
rect 9979 1042 9983 1074
rect 9943 1006 9983 1042
rect 9943 974 9947 1006
rect 9947 974 9979 1006
rect 9979 974 9983 1006
rect 9943 938 9983 974
rect 9943 906 9947 938
rect 9947 906 9979 938
rect 9979 906 9983 938
rect 9943 870 9983 906
rect 9943 838 9947 870
rect 9947 838 9979 870
rect 9979 838 9983 870
rect 9943 802 9983 838
rect 9943 770 9947 802
rect 9947 770 9979 802
rect 9979 770 9983 802
rect 9943 734 9983 770
rect 9943 702 9947 734
rect 9947 702 9979 734
rect 9979 702 9983 734
rect 9943 666 9983 702
rect 9943 634 9947 666
rect 9947 634 9979 666
rect 9979 634 9983 666
rect 9943 598 9983 634
rect 9943 566 9947 598
rect 9947 566 9979 598
rect 9979 566 9983 598
rect 9943 560 9983 566
rect 11151 4318 11191 4324
rect 11151 4286 11155 4318
rect 11155 4286 11187 4318
rect 11187 4286 11191 4318
rect 11151 4250 11191 4286
rect 11151 4218 11155 4250
rect 11155 4218 11187 4250
rect 11187 4218 11191 4250
rect 11151 4182 11191 4218
rect 11151 4150 11155 4182
rect 11155 4150 11187 4182
rect 11187 4150 11191 4182
rect 11151 4114 11191 4150
rect 11151 4082 11155 4114
rect 11155 4082 11187 4114
rect 11187 4082 11191 4114
rect 11151 4046 11191 4082
rect 11151 4014 11155 4046
rect 11155 4014 11187 4046
rect 11187 4014 11191 4046
rect 11151 3978 11191 4014
rect 11151 3946 11155 3978
rect 11155 3946 11187 3978
rect 11187 3946 11191 3978
rect 11151 3910 11191 3946
rect 11151 3878 11155 3910
rect 11155 3878 11187 3910
rect 11187 3878 11191 3910
rect 11151 3842 11191 3878
rect 11151 3810 11155 3842
rect 11155 3810 11187 3842
rect 11187 3810 11191 3842
rect 11151 3774 11191 3810
rect 11151 3742 11155 3774
rect 11155 3742 11187 3774
rect 11187 3742 11191 3774
rect 11151 3706 11191 3742
rect 11151 3674 11155 3706
rect 11155 3674 11187 3706
rect 11187 3674 11191 3706
rect 11151 3638 11191 3674
rect 11151 3606 11155 3638
rect 11155 3606 11187 3638
rect 11187 3606 11191 3638
rect 11151 3570 11191 3606
rect 11151 3538 11155 3570
rect 11155 3538 11187 3570
rect 11187 3538 11191 3570
rect 11151 3502 11191 3538
rect 11151 3470 11155 3502
rect 11155 3470 11187 3502
rect 11187 3470 11191 3502
rect 11151 3464 11191 3470
rect 10808 3350 10930 3356
rect 10808 3318 10853 3350
rect 10853 3318 10885 3350
rect 10885 3318 10930 3350
rect 10808 3282 10930 3318
rect 10808 3250 10853 3282
rect 10853 3250 10885 3282
rect 10885 3250 10930 3282
rect 10808 3214 10930 3250
rect 10808 3182 10853 3214
rect 10853 3182 10885 3214
rect 10885 3182 10930 3214
rect 10808 3146 10930 3182
rect 10808 3114 10853 3146
rect 10853 3114 10885 3146
rect 10885 3114 10930 3146
rect 10808 3078 10930 3114
rect 10808 3046 10853 3078
rect 10853 3046 10885 3078
rect 10885 3046 10930 3078
rect 10808 3010 10930 3046
rect 10808 2978 10853 3010
rect 10853 2978 10885 3010
rect 10885 2978 10930 3010
rect 10808 2942 10930 2978
rect 10808 2910 10853 2942
rect 10853 2910 10885 2942
rect 10885 2910 10930 2942
rect 10808 2874 10930 2910
rect 10808 2842 10853 2874
rect 10853 2842 10885 2874
rect 10885 2842 10930 2874
rect 10808 2806 10930 2842
rect 10808 2774 10853 2806
rect 10853 2774 10885 2806
rect 10885 2774 10930 2806
rect 10808 2738 10930 2774
rect 10808 2706 10853 2738
rect 10853 2706 10885 2738
rect 10885 2706 10930 2738
rect 10808 2670 10930 2706
rect 10808 2638 10853 2670
rect 10853 2638 10885 2670
rect 10885 2638 10930 2670
rect 10808 2602 10930 2638
rect 10808 2570 10853 2602
rect 10853 2570 10885 2602
rect 10885 2570 10930 2602
rect 10808 2534 10930 2570
rect 10808 2502 10853 2534
rect 10853 2502 10885 2534
rect 10885 2502 10930 2534
rect 10808 2496 10930 2502
rect 10547 2382 10587 2388
rect 10547 2350 10551 2382
rect 10551 2350 10583 2382
rect 10583 2350 10587 2382
rect 10547 2314 10587 2350
rect 10547 2282 10551 2314
rect 10551 2282 10583 2314
rect 10583 2282 10587 2314
rect 10547 2246 10587 2282
rect 10547 2214 10551 2246
rect 10551 2214 10583 2246
rect 10583 2214 10587 2246
rect 10547 2178 10587 2214
rect 10547 2146 10551 2178
rect 10551 2146 10583 2178
rect 10583 2146 10587 2178
rect 10547 2110 10587 2146
rect 10547 2078 10551 2110
rect 10551 2078 10583 2110
rect 10583 2078 10587 2110
rect 10547 2042 10587 2078
rect 10547 2010 10551 2042
rect 10551 2010 10583 2042
rect 10583 2010 10587 2042
rect 10547 1974 10587 2010
rect 10547 1942 10551 1974
rect 10551 1942 10583 1974
rect 10583 1942 10587 1974
rect 10547 1906 10587 1942
rect 10547 1874 10551 1906
rect 10551 1874 10583 1906
rect 10583 1874 10587 1906
rect 10547 1838 10587 1874
rect 10547 1806 10551 1838
rect 10551 1806 10583 1838
rect 10583 1806 10587 1838
rect 10547 1770 10587 1806
rect 10547 1738 10551 1770
rect 10551 1738 10583 1770
rect 10583 1738 10587 1770
rect 10547 1702 10587 1738
rect 10547 1670 10551 1702
rect 10551 1670 10583 1702
rect 10583 1670 10587 1702
rect 10547 1634 10587 1670
rect 10547 1602 10551 1634
rect 10551 1602 10583 1634
rect 10583 1602 10587 1634
rect 10547 1566 10587 1602
rect 10547 1534 10551 1566
rect 10551 1534 10583 1566
rect 10583 1534 10587 1566
rect 10547 1528 10587 1534
rect 10204 1414 10326 1420
rect 10204 1382 10249 1414
rect 10249 1382 10281 1414
rect 10281 1382 10326 1414
rect 10204 1346 10326 1382
rect 10204 1314 10249 1346
rect 10249 1314 10281 1346
rect 10281 1314 10326 1346
rect 10204 1278 10326 1314
rect 10204 1246 10249 1278
rect 10249 1246 10281 1278
rect 10281 1246 10326 1278
rect 10204 1210 10326 1246
rect 10204 1178 10249 1210
rect 10249 1178 10281 1210
rect 10281 1178 10326 1210
rect 10204 1142 10326 1178
rect 10204 1110 10249 1142
rect 10249 1110 10281 1142
rect 10281 1110 10326 1142
rect 10204 1074 10326 1110
rect 10204 1042 10249 1074
rect 10249 1042 10281 1074
rect 10281 1042 10326 1074
rect 10204 1006 10326 1042
rect 10204 974 10249 1006
rect 10249 974 10281 1006
rect 10281 974 10326 1006
rect 10204 938 10326 974
rect 10204 906 10249 938
rect 10249 906 10281 938
rect 10281 906 10326 938
rect 10204 870 10326 906
rect 10204 838 10249 870
rect 10249 838 10281 870
rect 10281 838 10326 870
rect 10204 802 10326 838
rect 10204 770 10249 802
rect 10249 770 10281 802
rect 10281 770 10326 802
rect 10204 734 10326 770
rect 10204 702 10249 734
rect 10249 702 10281 734
rect 10281 702 10326 734
rect 10204 666 10326 702
rect 10204 634 10249 666
rect 10249 634 10281 666
rect 10281 634 10326 666
rect 10204 598 10326 634
rect 10204 566 10249 598
rect 10249 566 10281 598
rect 10281 566 10326 598
rect 10204 560 10326 566
rect 11412 4318 11534 4324
rect 11412 4286 11457 4318
rect 11457 4286 11489 4318
rect 11489 4286 11534 4318
rect 11412 4250 11534 4286
rect 11412 4218 11457 4250
rect 11457 4218 11489 4250
rect 11489 4218 11534 4250
rect 11412 4182 11534 4218
rect 11412 4150 11457 4182
rect 11457 4150 11489 4182
rect 11489 4150 11534 4182
rect 11412 4114 11534 4150
rect 11412 4082 11457 4114
rect 11457 4082 11489 4114
rect 11489 4082 11534 4114
rect 11412 4046 11534 4082
rect 11412 4014 11457 4046
rect 11457 4014 11489 4046
rect 11489 4014 11534 4046
rect 11412 3978 11534 4014
rect 11412 3946 11457 3978
rect 11457 3946 11489 3978
rect 11489 3946 11534 3978
rect 11412 3910 11534 3946
rect 11412 3878 11457 3910
rect 11457 3878 11489 3910
rect 11489 3878 11534 3910
rect 11412 3842 11534 3878
rect 11412 3810 11457 3842
rect 11457 3810 11489 3842
rect 11489 3810 11534 3842
rect 11412 3774 11534 3810
rect 11412 3742 11457 3774
rect 11457 3742 11489 3774
rect 11489 3742 11534 3774
rect 11412 3706 11534 3742
rect 11412 3674 11457 3706
rect 11457 3674 11489 3706
rect 11489 3674 11534 3706
rect 11412 3638 11534 3674
rect 11412 3606 11457 3638
rect 11457 3606 11489 3638
rect 11489 3606 11534 3638
rect 11412 3570 11534 3606
rect 11412 3538 11457 3570
rect 11457 3538 11489 3570
rect 11489 3538 11534 3570
rect 11412 3502 11534 3538
rect 11412 3470 11457 3502
rect 11457 3470 11489 3502
rect 11489 3470 11534 3502
rect 11412 3464 11534 3470
rect 11151 3350 11191 3356
rect 11151 3318 11155 3350
rect 11155 3318 11187 3350
rect 11187 3318 11191 3350
rect 11151 3282 11191 3318
rect 11151 3250 11155 3282
rect 11155 3250 11187 3282
rect 11187 3250 11191 3282
rect 11151 3214 11191 3250
rect 11151 3182 11155 3214
rect 11155 3182 11187 3214
rect 11187 3182 11191 3214
rect 11151 3146 11191 3182
rect 11151 3114 11155 3146
rect 11155 3114 11187 3146
rect 11187 3114 11191 3146
rect 11151 3078 11191 3114
rect 11151 3046 11155 3078
rect 11155 3046 11187 3078
rect 11187 3046 11191 3078
rect 11151 3010 11191 3046
rect 11151 2978 11155 3010
rect 11155 2978 11187 3010
rect 11187 2978 11191 3010
rect 11151 2942 11191 2978
rect 11151 2910 11155 2942
rect 11155 2910 11187 2942
rect 11187 2910 11191 2942
rect 11151 2874 11191 2910
rect 11151 2842 11155 2874
rect 11155 2842 11187 2874
rect 11187 2842 11191 2874
rect 11151 2806 11191 2842
rect 11151 2774 11155 2806
rect 11155 2774 11187 2806
rect 11187 2774 11191 2806
rect 11151 2738 11191 2774
rect 11151 2706 11155 2738
rect 11155 2706 11187 2738
rect 11187 2706 11191 2738
rect 11151 2670 11191 2706
rect 11151 2638 11155 2670
rect 11155 2638 11187 2670
rect 11187 2638 11191 2670
rect 11151 2602 11191 2638
rect 11151 2570 11155 2602
rect 11155 2570 11187 2602
rect 11187 2570 11191 2602
rect 11151 2534 11191 2570
rect 11151 2502 11155 2534
rect 11155 2502 11187 2534
rect 11187 2502 11191 2534
rect 11151 2496 11191 2502
rect 10808 2382 10930 2388
rect 10808 2350 10853 2382
rect 10853 2350 10885 2382
rect 10885 2350 10930 2382
rect 10808 2314 10930 2350
rect 10808 2282 10853 2314
rect 10853 2282 10885 2314
rect 10885 2282 10930 2314
rect 10808 2246 10930 2282
rect 10808 2214 10853 2246
rect 10853 2214 10885 2246
rect 10885 2214 10930 2246
rect 10808 2178 10930 2214
rect 10808 2146 10853 2178
rect 10853 2146 10885 2178
rect 10885 2146 10930 2178
rect 10808 2110 10930 2146
rect 10808 2078 10853 2110
rect 10853 2078 10885 2110
rect 10885 2078 10930 2110
rect 10808 2042 10930 2078
rect 10808 2010 10853 2042
rect 10853 2010 10885 2042
rect 10885 2010 10930 2042
rect 10808 1974 10930 2010
rect 10808 1942 10853 1974
rect 10853 1942 10885 1974
rect 10885 1942 10930 1974
rect 10808 1906 10930 1942
rect 10808 1874 10853 1906
rect 10853 1874 10885 1906
rect 10885 1874 10930 1906
rect 10808 1838 10930 1874
rect 10808 1806 10853 1838
rect 10853 1806 10885 1838
rect 10885 1806 10930 1838
rect 10808 1770 10930 1806
rect 10808 1738 10853 1770
rect 10853 1738 10885 1770
rect 10885 1738 10930 1770
rect 10808 1702 10930 1738
rect 10808 1670 10853 1702
rect 10853 1670 10885 1702
rect 10885 1670 10930 1702
rect 10808 1634 10930 1670
rect 10808 1602 10853 1634
rect 10853 1602 10885 1634
rect 10885 1602 10930 1634
rect 10808 1566 10930 1602
rect 10808 1534 10853 1566
rect 10853 1534 10885 1566
rect 10885 1534 10930 1566
rect 10808 1528 10930 1534
rect 10547 1414 10587 1420
rect 10547 1382 10551 1414
rect 10551 1382 10583 1414
rect 10583 1382 10587 1414
rect 10547 1346 10587 1382
rect 10547 1314 10551 1346
rect 10551 1314 10583 1346
rect 10583 1314 10587 1346
rect 10547 1278 10587 1314
rect 10547 1246 10551 1278
rect 10551 1246 10583 1278
rect 10583 1246 10587 1278
rect 10547 1210 10587 1246
rect 10547 1178 10551 1210
rect 10551 1178 10583 1210
rect 10583 1178 10587 1210
rect 10547 1142 10587 1178
rect 10547 1110 10551 1142
rect 10551 1110 10583 1142
rect 10583 1110 10587 1142
rect 10547 1074 10587 1110
rect 10547 1042 10551 1074
rect 10551 1042 10583 1074
rect 10583 1042 10587 1074
rect 10547 1006 10587 1042
rect 10547 974 10551 1006
rect 10551 974 10583 1006
rect 10583 974 10587 1006
rect 10547 938 10587 974
rect 10547 906 10551 938
rect 10551 906 10583 938
rect 10583 906 10587 938
rect 10547 870 10587 906
rect 10547 838 10551 870
rect 10551 838 10583 870
rect 10583 838 10587 870
rect 10547 802 10587 838
rect 10547 770 10551 802
rect 10551 770 10583 802
rect 10583 770 10587 802
rect 10547 734 10587 770
rect 10547 702 10551 734
rect 10551 702 10583 734
rect 10583 702 10587 734
rect 10547 666 10587 702
rect 10547 634 10551 666
rect 10551 634 10583 666
rect 10583 634 10587 666
rect 10547 598 10587 634
rect 10547 566 10551 598
rect 10551 566 10583 598
rect 10583 566 10587 598
rect 10547 560 10587 566
rect 11755 4318 11795 4324
rect 11755 4286 11759 4318
rect 11759 4286 11791 4318
rect 11791 4286 11795 4318
rect 11755 4250 11795 4286
rect 11755 4218 11759 4250
rect 11759 4218 11791 4250
rect 11791 4218 11795 4250
rect 11755 4182 11795 4218
rect 11755 4150 11759 4182
rect 11759 4150 11791 4182
rect 11791 4150 11795 4182
rect 11755 4114 11795 4150
rect 11755 4082 11759 4114
rect 11759 4082 11791 4114
rect 11791 4082 11795 4114
rect 11755 4046 11795 4082
rect 11755 4014 11759 4046
rect 11759 4014 11791 4046
rect 11791 4014 11795 4046
rect 11755 3978 11795 4014
rect 11755 3946 11759 3978
rect 11759 3946 11791 3978
rect 11791 3946 11795 3978
rect 11755 3910 11795 3946
rect 11755 3878 11759 3910
rect 11759 3878 11791 3910
rect 11791 3878 11795 3910
rect 11755 3842 11795 3878
rect 11755 3810 11759 3842
rect 11759 3810 11791 3842
rect 11791 3810 11795 3842
rect 11755 3774 11795 3810
rect 11755 3742 11759 3774
rect 11759 3742 11791 3774
rect 11791 3742 11795 3774
rect 11755 3706 11795 3742
rect 11755 3674 11759 3706
rect 11759 3674 11791 3706
rect 11791 3674 11795 3706
rect 11755 3638 11795 3674
rect 11755 3606 11759 3638
rect 11759 3606 11791 3638
rect 11791 3606 11795 3638
rect 11755 3570 11795 3606
rect 11755 3538 11759 3570
rect 11759 3538 11791 3570
rect 11791 3538 11795 3570
rect 11755 3502 11795 3538
rect 11755 3470 11759 3502
rect 11759 3470 11791 3502
rect 11791 3470 11795 3502
rect 11755 3464 11795 3470
rect 11412 3350 11534 3356
rect 11412 3318 11457 3350
rect 11457 3318 11489 3350
rect 11489 3318 11534 3350
rect 11412 3282 11534 3318
rect 11412 3250 11457 3282
rect 11457 3250 11489 3282
rect 11489 3250 11534 3282
rect 11412 3214 11534 3250
rect 11412 3182 11457 3214
rect 11457 3182 11489 3214
rect 11489 3182 11534 3214
rect 11412 3146 11534 3182
rect 11412 3114 11457 3146
rect 11457 3114 11489 3146
rect 11489 3114 11534 3146
rect 11412 3078 11534 3114
rect 11412 3046 11457 3078
rect 11457 3046 11489 3078
rect 11489 3046 11534 3078
rect 11412 3010 11534 3046
rect 11412 2978 11457 3010
rect 11457 2978 11489 3010
rect 11489 2978 11534 3010
rect 11412 2942 11534 2978
rect 11412 2910 11457 2942
rect 11457 2910 11489 2942
rect 11489 2910 11534 2942
rect 11412 2874 11534 2910
rect 11412 2842 11457 2874
rect 11457 2842 11489 2874
rect 11489 2842 11534 2874
rect 11412 2806 11534 2842
rect 11412 2774 11457 2806
rect 11457 2774 11489 2806
rect 11489 2774 11534 2806
rect 11412 2738 11534 2774
rect 11412 2706 11457 2738
rect 11457 2706 11489 2738
rect 11489 2706 11534 2738
rect 11412 2670 11534 2706
rect 11412 2638 11457 2670
rect 11457 2638 11489 2670
rect 11489 2638 11534 2670
rect 11412 2602 11534 2638
rect 11412 2570 11457 2602
rect 11457 2570 11489 2602
rect 11489 2570 11534 2602
rect 11412 2534 11534 2570
rect 11412 2502 11457 2534
rect 11457 2502 11489 2534
rect 11489 2502 11534 2534
rect 11412 2496 11534 2502
rect 11151 2382 11191 2388
rect 11151 2350 11155 2382
rect 11155 2350 11187 2382
rect 11187 2350 11191 2382
rect 11151 2314 11191 2350
rect 11151 2282 11155 2314
rect 11155 2282 11187 2314
rect 11187 2282 11191 2314
rect 11151 2246 11191 2282
rect 11151 2214 11155 2246
rect 11155 2214 11187 2246
rect 11187 2214 11191 2246
rect 11151 2178 11191 2214
rect 11151 2146 11155 2178
rect 11155 2146 11187 2178
rect 11187 2146 11191 2178
rect 11151 2110 11191 2146
rect 11151 2078 11155 2110
rect 11155 2078 11187 2110
rect 11187 2078 11191 2110
rect 11151 2042 11191 2078
rect 11151 2010 11155 2042
rect 11155 2010 11187 2042
rect 11187 2010 11191 2042
rect 11151 1974 11191 2010
rect 11151 1942 11155 1974
rect 11155 1942 11187 1974
rect 11187 1942 11191 1974
rect 11151 1906 11191 1942
rect 11151 1874 11155 1906
rect 11155 1874 11187 1906
rect 11187 1874 11191 1906
rect 11151 1838 11191 1874
rect 11151 1806 11155 1838
rect 11155 1806 11187 1838
rect 11187 1806 11191 1838
rect 11151 1770 11191 1806
rect 11151 1738 11155 1770
rect 11155 1738 11187 1770
rect 11187 1738 11191 1770
rect 11151 1702 11191 1738
rect 11151 1670 11155 1702
rect 11155 1670 11187 1702
rect 11187 1670 11191 1702
rect 11151 1634 11191 1670
rect 11151 1602 11155 1634
rect 11155 1602 11187 1634
rect 11187 1602 11191 1634
rect 11151 1566 11191 1602
rect 11151 1534 11155 1566
rect 11155 1534 11187 1566
rect 11187 1534 11191 1566
rect 11151 1528 11191 1534
rect 10808 1414 10930 1420
rect 10808 1382 10853 1414
rect 10853 1382 10885 1414
rect 10885 1382 10930 1414
rect 10808 1346 10930 1382
rect 10808 1314 10853 1346
rect 10853 1314 10885 1346
rect 10885 1314 10930 1346
rect 10808 1278 10930 1314
rect 10808 1246 10853 1278
rect 10853 1246 10885 1278
rect 10885 1246 10930 1278
rect 10808 1210 10930 1246
rect 10808 1178 10853 1210
rect 10853 1178 10885 1210
rect 10885 1178 10930 1210
rect 10808 1142 10930 1178
rect 10808 1110 10853 1142
rect 10853 1110 10885 1142
rect 10885 1110 10930 1142
rect 10808 1074 10930 1110
rect 10808 1042 10853 1074
rect 10853 1042 10885 1074
rect 10885 1042 10930 1074
rect 10808 1006 10930 1042
rect 10808 974 10853 1006
rect 10853 974 10885 1006
rect 10885 974 10930 1006
rect 10808 938 10930 974
rect 10808 906 10853 938
rect 10853 906 10885 938
rect 10885 906 10930 938
rect 10808 870 10930 906
rect 10808 838 10853 870
rect 10853 838 10885 870
rect 10885 838 10930 870
rect 10808 802 10930 838
rect 10808 770 10853 802
rect 10853 770 10885 802
rect 10885 770 10930 802
rect 10808 734 10930 770
rect 10808 702 10853 734
rect 10853 702 10885 734
rect 10885 702 10930 734
rect 10808 666 10930 702
rect 10808 634 10853 666
rect 10853 634 10885 666
rect 10885 634 10930 666
rect 10808 598 10930 634
rect 10808 566 10853 598
rect 10853 566 10885 598
rect 10885 566 10930 598
rect 10808 560 10930 566
rect 12016 4318 12138 4324
rect 12016 4286 12061 4318
rect 12061 4286 12093 4318
rect 12093 4286 12138 4318
rect 12016 4250 12138 4286
rect 12016 4218 12061 4250
rect 12061 4218 12093 4250
rect 12093 4218 12138 4250
rect 12016 4182 12138 4218
rect 12016 4150 12061 4182
rect 12061 4150 12093 4182
rect 12093 4150 12138 4182
rect 12016 4114 12138 4150
rect 12016 4082 12061 4114
rect 12061 4082 12093 4114
rect 12093 4082 12138 4114
rect 12016 4046 12138 4082
rect 12016 4014 12061 4046
rect 12061 4014 12093 4046
rect 12093 4014 12138 4046
rect 12016 3978 12138 4014
rect 12016 3946 12061 3978
rect 12061 3946 12093 3978
rect 12093 3946 12138 3978
rect 12016 3910 12138 3946
rect 12016 3878 12061 3910
rect 12061 3878 12093 3910
rect 12093 3878 12138 3910
rect 12016 3842 12138 3878
rect 12016 3810 12061 3842
rect 12061 3810 12093 3842
rect 12093 3810 12138 3842
rect 12016 3774 12138 3810
rect 12016 3742 12061 3774
rect 12061 3742 12093 3774
rect 12093 3742 12138 3774
rect 12016 3706 12138 3742
rect 12016 3674 12061 3706
rect 12061 3674 12093 3706
rect 12093 3674 12138 3706
rect 12016 3638 12138 3674
rect 12016 3606 12061 3638
rect 12061 3606 12093 3638
rect 12093 3606 12138 3638
rect 12016 3570 12138 3606
rect 12016 3538 12061 3570
rect 12061 3538 12093 3570
rect 12093 3538 12138 3570
rect 12016 3502 12138 3538
rect 12016 3470 12061 3502
rect 12061 3470 12093 3502
rect 12093 3470 12138 3502
rect 12016 3464 12138 3470
rect 11755 3350 11795 3356
rect 11755 3318 11759 3350
rect 11759 3318 11791 3350
rect 11791 3318 11795 3350
rect 11755 3282 11795 3318
rect 11755 3250 11759 3282
rect 11759 3250 11791 3282
rect 11791 3250 11795 3282
rect 11755 3214 11795 3250
rect 11755 3182 11759 3214
rect 11759 3182 11791 3214
rect 11791 3182 11795 3214
rect 11755 3146 11795 3182
rect 11755 3114 11759 3146
rect 11759 3114 11791 3146
rect 11791 3114 11795 3146
rect 11755 3078 11795 3114
rect 11755 3046 11759 3078
rect 11759 3046 11791 3078
rect 11791 3046 11795 3078
rect 11755 3010 11795 3046
rect 11755 2978 11759 3010
rect 11759 2978 11791 3010
rect 11791 2978 11795 3010
rect 11755 2942 11795 2978
rect 11755 2910 11759 2942
rect 11759 2910 11791 2942
rect 11791 2910 11795 2942
rect 11755 2874 11795 2910
rect 11755 2842 11759 2874
rect 11759 2842 11791 2874
rect 11791 2842 11795 2874
rect 11755 2806 11795 2842
rect 11755 2774 11759 2806
rect 11759 2774 11791 2806
rect 11791 2774 11795 2806
rect 11755 2738 11795 2774
rect 11755 2706 11759 2738
rect 11759 2706 11791 2738
rect 11791 2706 11795 2738
rect 11755 2670 11795 2706
rect 11755 2638 11759 2670
rect 11759 2638 11791 2670
rect 11791 2638 11795 2670
rect 11755 2602 11795 2638
rect 11755 2570 11759 2602
rect 11759 2570 11791 2602
rect 11791 2570 11795 2602
rect 11755 2534 11795 2570
rect 11755 2502 11759 2534
rect 11759 2502 11791 2534
rect 11791 2502 11795 2534
rect 11755 2496 11795 2502
rect 11412 2382 11534 2388
rect 11412 2350 11457 2382
rect 11457 2350 11489 2382
rect 11489 2350 11534 2382
rect 11412 2314 11534 2350
rect 11412 2282 11457 2314
rect 11457 2282 11489 2314
rect 11489 2282 11534 2314
rect 11412 2246 11534 2282
rect 11412 2214 11457 2246
rect 11457 2214 11489 2246
rect 11489 2214 11534 2246
rect 11412 2178 11534 2214
rect 11412 2146 11457 2178
rect 11457 2146 11489 2178
rect 11489 2146 11534 2178
rect 11412 2110 11534 2146
rect 11412 2078 11457 2110
rect 11457 2078 11489 2110
rect 11489 2078 11534 2110
rect 11412 2042 11534 2078
rect 11412 2010 11457 2042
rect 11457 2010 11489 2042
rect 11489 2010 11534 2042
rect 11412 1974 11534 2010
rect 11412 1942 11457 1974
rect 11457 1942 11489 1974
rect 11489 1942 11534 1974
rect 11412 1906 11534 1942
rect 11412 1874 11457 1906
rect 11457 1874 11489 1906
rect 11489 1874 11534 1906
rect 11412 1838 11534 1874
rect 11412 1806 11457 1838
rect 11457 1806 11489 1838
rect 11489 1806 11534 1838
rect 11412 1770 11534 1806
rect 11412 1738 11457 1770
rect 11457 1738 11489 1770
rect 11489 1738 11534 1770
rect 11412 1702 11534 1738
rect 11412 1670 11457 1702
rect 11457 1670 11489 1702
rect 11489 1670 11534 1702
rect 11412 1634 11534 1670
rect 11412 1602 11457 1634
rect 11457 1602 11489 1634
rect 11489 1602 11534 1634
rect 11412 1566 11534 1602
rect 11412 1534 11457 1566
rect 11457 1534 11489 1566
rect 11489 1534 11534 1566
rect 11412 1528 11534 1534
rect 11151 1414 11191 1420
rect 11151 1382 11155 1414
rect 11155 1382 11187 1414
rect 11187 1382 11191 1414
rect 11151 1346 11191 1382
rect 11151 1314 11155 1346
rect 11155 1314 11187 1346
rect 11187 1314 11191 1346
rect 11151 1278 11191 1314
rect 11151 1246 11155 1278
rect 11155 1246 11187 1278
rect 11187 1246 11191 1278
rect 11151 1210 11191 1246
rect 11151 1178 11155 1210
rect 11155 1178 11187 1210
rect 11187 1178 11191 1210
rect 11151 1142 11191 1178
rect 11151 1110 11155 1142
rect 11155 1110 11187 1142
rect 11187 1110 11191 1142
rect 11151 1074 11191 1110
rect 11151 1042 11155 1074
rect 11155 1042 11187 1074
rect 11187 1042 11191 1074
rect 11151 1006 11191 1042
rect 11151 974 11155 1006
rect 11155 974 11187 1006
rect 11187 974 11191 1006
rect 11151 938 11191 974
rect 11151 906 11155 938
rect 11155 906 11187 938
rect 11187 906 11191 938
rect 11151 870 11191 906
rect 11151 838 11155 870
rect 11155 838 11187 870
rect 11187 838 11191 870
rect 11151 802 11191 838
rect 11151 770 11155 802
rect 11155 770 11187 802
rect 11187 770 11191 802
rect 11151 734 11191 770
rect 11151 702 11155 734
rect 11155 702 11187 734
rect 11187 702 11191 734
rect 11151 666 11191 702
rect 11151 634 11155 666
rect 11155 634 11187 666
rect 11187 634 11191 666
rect 11151 598 11191 634
rect 11151 566 11155 598
rect 11155 566 11187 598
rect 11187 566 11191 598
rect 11151 560 11191 566
rect 12359 4318 12399 4324
rect 12359 4286 12363 4318
rect 12363 4286 12395 4318
rect 12395 4286 12399 4318
rect 12359 4250 12399 4286
rect 12359 4218 12363 4250
rect 12363 4218 12395 4250
rect 12395 4218 12399 4250
rect 12359 4182 12399 4218
rect 12359 4150 12363 4182
rect 12363 4150 12395 4182
rect 12395 4150 12399 4182
rect 12359 4114 12399 4150
rect 12359 4082 12363 4114
rect 12363 4082 12395 4114
rect 12395 4082 12399 4114
rect 12359 4046 12399 4082
rect 12359 4014 12363 4046
rect 12363 4014 12395 4046
rect 12395 4014 12399 4046
rect 12359 3978 12399 4014
rect 12359 3946 12363 3978
rect 12363 3946 12395 3978
rect 12395 3946 12399 3978
rect 12359 3910 12399 3946
rect 12359 3878 12363 3910
rect 12363 3878 12395 3910
rect 12395 3878 12399 3910
rect 12359 3842 12399 3878
rect 12359 3810 12363 3842
rect 12363 3810 12395 3842
rect 12395 3810 12399 3842
rect 12359 3774 12399 3810
rect 12359 3742 12363 3774
rect 12363 3742 12395 3774
rect 12395 3742 12399 3774
rect 12359 3706 12399 3742
rect 12359 3674 12363 3706
rect 12363 3674 12395 3706
rect 12395 3674 12399 3706
rect 12359 3638 12399 3674
rect 12359 3606 12363 3638
rect 12363 3606 12395 3638
rect 12395 3606 12399 3638
rect 12359 3570 12399 3606
rect 12359 3538 12363 3570
rect 12363 3538 12395 3570
rect 12395 3538 12399 3570
rect 12359 3502 12399 3538
rect 12359 3470 12363 3502
rect 12363 3470 12395 3502
rect 12395 3470 12399 3502
rect 12359 3464 12399 3470
rect 12016 3350 12138 3356
rect 12016 3318 12061 3350
rect 12061 3318 12093 3350
rect 12093 3318 12138 3350
rect 12016 3282 12138 3318
rect 12016 3250 12061 3282
rect 12061 3250 12093 3282
rect 12093 3250 12138 3282
rect 12016 3214 12138 3250
rect 12016 3182 12061 3214
rect 12061 3182 12093 3214
rect 12093 3182 12138 3214
rect 12016 3146 12138 3182
rect 12016 3114 12061 3146
rect 12061 3114 12093 3146
rect 12093 3114 12138 3146
rect 12016 3078 12138 3114
rect 12016 3046 12061 3078
rect 12061 3046 12093 3078
rect 12093 3046 12138 3078
rect 12016 3010 12138 3046
rect 12016 2978 12061 3010
rect 12061 2978 12093 3010
rect 12093 2978 12138 3010
rect 12016 2942 12138 2978
rect 12016 2910 12061 2942
rect 12061 2910 12093 2942
rect 12093 2910 12138 2942
rect 12016 2874 12138 2910
rect 12016 2842 12061 2874
rect 12061 2842 12093 2874
rect 12093 2842 12138 2874
rect 12016 2806 12138 2842
rect 12016 2774 12061 2806
rect 12061 2774 12093 2806
rect 12093 2774 12138 2806
rect 12016 2738 12138 2774
rect 12016 2706 12061 2738
rect 12061 2706 12093 2738
rect 12093 2706 12138 2738
rect 12016 2670 12138 2706
rect 12016 2638 12061 2670
rect 12061 2638 12093 2670
rect 12093 2638 12138 2670
rect 12016 2602 12138 2638
rect 12016 2570 12061 2602
rect 12061 2570 12093 2602
rect 12093 2570 12138 2602
rect 12016 2534 12138 2570
rect 12016 2502 12061 2534
rect 12061 2502 12093 2534
rect 12093 2502 12138 2534
rect 12016 2496 12138 2502
rect 11755 2382 11795 2388
rect 11755 2350 11759 2382
rect 11759 2350 11791 2382
rect 11791 2350 11795 2382
rect 11755 2314 11795 2350
rect 11755 2282 11759 2314
rect 11759 2282 11791 2314
rect 11791 2282 11795 2314
rect 11755 2246 11795 2282
rect 11755 2214 11759 2246
rect 11759 2214 11791 2246
rect 11791 2214 11795 2246
rect 11755 2178 11795 2214
rect 11755 2146 11759 2178
rect 11759 2146 11791 2178
rect 11791 2146 11795 2178
rect 11755 2110 11795 2146
rect 11755 2078 11759 2110
rect 11759 2078 11791 2110
rect 11791 2078 11795 2110
rect 11755 2042 11795 2078
rect 11755 2010 11759 2042
rect 11759 2010 11791 2042
rect 11791 2010 11795 2042
rect 11755 1974 11795 2010
rect 11755 1942 11759 1974
rect 11759 1942 11791 1974
rect 11791 1942 11795 1974
rect 11755 1906 11795 1942
rect 11755 1874 11759 1906
rect 11759 1874 11791 1906
rect 11791 1874 11795 1906
rect 11755 1838 11795 1874
rect 11755 1806 11759 1838
rect 11759 1806 11791 1838
rect 11791 1806 11795 1838
rect 11755 1770 11795 1806
rect 11755 1738 11759 1770
rect 11759 1738 11791 1770
rect 11791 1738 11795 1770
rect 11755 1702 11795 1738
rect 11755 1670 11759 1702
rect 11759 1670 11791 1702
rect 11791 1670 11795 1702
rect 11755 1634 11795 1670
rect 11755 1602 11759 1634
rect 11759 1602 11791 1634
rect 11791 1602 11795 1634
rect 11755 1566 11795 1602
rect 11755 1534 11759 1566
rect 11759 1534 11791 1566
rect 11791 1534 11795 1566
rect 11755 1528 11795 1534
rect 11412 1414 11534 1420
rect 11412 1382 11457 1414
rect 11457 1382 11489 1414
rect 11489 1382 11534 1414
rect 11412 1346 11534 1382
rect 11412 1314 11457 1346
rect 11457 1314 11489 1346
rect 11489 1314 11534 1346
rect 11412 1278 11534 1314
rect 11412 1246 11457 1278
rect 11457 1246 11489 1278
rect 11489 1246 11534 1278
rect 11412 1210 11534 1246
rect 11412 1178 11457 1210
rect 11457 1178 11489 1210
rect 11489 1178 11534 1210
rect 11412 1142 11534 1178
rect 11412 1110 11457 1142
rect 11457 1110 11489 1142
rect 11489 1110 11534 1142
rect 11412 1074 11534 1110
rect 11412 1042 11457 1074
rect 11457 1042 11489 1074
rect 11489 1042 11534 1074
rect 11412 1006 11534 1042
rect 11412 974 11457 1006
rect 11457 974 11489 1006
rect 11489 974 11534 1006
rect 11412 938 11534 974
rect 11412 906 11457 938
rect 11457 906 11489 938
rect 11489 906 11534 938
rect 11412 870 11534 906
rect 11412 838 11457 870
rect 11457 838 11489 870
rect 11489 838 11534 870
rect 11412 802 11534 838
rect 11412 770 11457 802
rect 11457 770 11489 802
rect 11489 770 11534 802
rect 11412 734 11534 770
rect 11412 702 11457 734
rect 11457 702 11489 734
rect 11489 702 11534 734
rect 11412 666 11534 702
rect 11412 634 11457 666
rect 11457 634 11489 666
rect 11489 634 11534 666
rect 11412 598 11534 634
rect 11412 566 11457 598
rect 11457 566 11489 598
rect 11489 566 11534 598
rect 11412 560 11534 566
rect 12620 4318 12742 4324
rect 12620 4286 12665 4318
rect 12665 4286 12697 4318
rect 12697 4286 12742 4318
rect 12620 4250 12742 4286
rect 12620 4218 12665 4250
rect 12665 4218 12697 4250
rect 12697 4218 12742 4250
rect 12620 4182 12742 4218
rect 12620 4150 12665 4182
rect 12665 4150 12697 4182
rect 12697 4150 12742 4182
rect 12620 4114 12742 4150
rect 12620 4082 12665 4114
rect 12665 4082 12697 4114
rect 12697 4082 12742 4114
rect 12620 4046 12742 4082
rect 12620 4014 12665 4046
rect 12665 4014 12697 4046
rect 12697 4014 12742 4046
rect 12620 3978 12742 4014
rect 12620 3946 12665 3978
rect 12665 3946 12697 3978
rect 12697 3946 12742 3978
rect 12620 3910 12742 3946
rect 12620 3878 12665 3910
rect 12665 3878 12697 3910
rect 12697 3878 12742 3910
rect 12620 3842 12742 3878
rect 12620 3810 12665 3842
rect 12665 3810 12697 3842
rect 12697 3810 12742 3842
rect 12620 3774 12742 3810
rect 12620 3742 12665 3774
rect 12665 3742 12697 3774
rect 12697 3742 12742 3774
rect 12620 3706 12742 3742
rect 12620 3674 12665 3706
rect 12665 3674 12697 3706
rect 12697 3674 12742 3706
rect 12620 3638 12742 3674
rect 12620 3606 12665 3638
rect 12665 3606 12697 3638
rect 12697 3606 12742 3638
rect 12620 3570 12742 3606
rect 12620 3538 12665 3570
rect 12665 3538 12697 3570
rect 12697 3538 12742 3570
rect 12620 3502 12742 3538
rect 12620 3470 12665 3502
rect 12665 3470 12697 3502
rect 12697 3470 12742 3502
rect 12620 3464 12742 3470
rect 12359 3350 12399 3356
rect 12359 3318 12363 3350
rect 12363 3318 12395 3350
rect 12395 3318 12399 3350
rect 12359 3282 12399 3318
rect 12359 3250 12363 3282
rect 12363 3250 12395 3282
rect 12395 3250 12399 3282
rect 12359 3214 12399 3250
rect 12359 3182 12363 3214
rect 12363 3182 12395 3214
rect 12395 3182 12399 3214
rect 12359 3146 12399 3182
rect 12359 3114 12363 3146
rect 12363 3114 12395 3146
rect 12395 3114 12399 3146
rect 12359 3078 12399 3114
rect 12359 3046 12363 3078
rect 12363 3046 12395 3078
rect 12395 3046 12399 3078
rect 12359 3010 12399 3046
rect 12359 2978 12363 3010
rect 12363 2978 12395 3010
rect 12395 2978 12399 3010
rect 12359 2942 12399 2978
rect 12359 2910 12363 2942
rect 12363 2910 12395 2942
rect 12395 2910 12399 2942
rect 12359 2874 12399 2910
rect 12359 2842 12363 2874
rect 12363 2842 12395 2874
rect 12395 2842 12399 2874
rect 12359 2806 12399 2842
rect 12359 2774 12363 2806
rect 12363 2774 12395 2806
rect 12395 2774 12399 2806
rect 12359 2738 12399 2774
rect 12359 2706 12363 2738
rect 12363 2706 12395 2738
rect 12395 2706 12399 2738
rect 12359 2670 12399 2706
rect 12359 2638 12363 2670
rect 12363 2638 12395 2670
rect 12395 2638 12399 2670
rect 12359 2602 12399 2638
rect 12359 2570 12363 2602
rect 12363 2570 12395 2602
rect 12395 2570 12399 2602
rect 12359 2534 12399 2570
rect 12359 2502 12363 2534
rect 12363 2502 12395 2534
rect 12395 2502 12399 2534
rect 12359 2496 12399 2502
rect 12016 2382 12138 2388
rect 12016 2350 12061 2382
rect 12061 2350 12093 2382
rect 12093 2350 12138 2382
rect 12016 2314 12138 2350
rect 12016 2282 12061 2314
rect 12061 2282 12093 2314
rect 12093 2282 12138 2314
rect 12016 2246 12138 2282
rect 12016 2214 12061 2246
rect 12061 2214 12093 2246
rect 12093 2214 12138 2246
rect 12016 2178 12138 2214
rect 12016 2146 12061 2178
rect 12061 2146 12093 2178
rect 12093 2146 12138 2178
rect 12016 2110 12138 2146
rect 12016 2078 12061 2110
rect 12061 2078 12093 2110
rect 12093 2078 12138 2110
rect 12016 2042 12138 2078
rect 12016 2010 12061 2042
rect 12061 2010 12093 2042
rect 12093 2010 12138 2042
rect 12016 1974 12138 2010
rect 12016 1942 12061 1974
rect 12061 1942 12093 1974
rect 12093 1942 12138 1974
rect 12016 1906 12138 1942
rect 12016 1874 12061 1906
rect 12061 1874 12093 1906
rect 12093 1874 12138 1906
rect 12016 1838 12138 1874
rect 12016 1806 12061 1838
rect 12061 1806 12093 1838
rect 12093 1806 12138 1838
rect 12016 1770 12138 1806
rect 12016 1738 12061 1770
rect 12061 1738 12093 1770
rect 12093 1738 12138 1770
rect 12016 1702 12138 1738
rect 12016 1670 12061 1702
rect 12061 1670 12093 1702
rect 12093 1670 12138 1702
rect 12016 1634 12138 1670
rect 12016 1602 12061 1634
rect 12061 1602 12093 1634
rect 12093 1602 12138 1634
rect 12016 1566 12138 1602
rect 12016 1534 12061 1566
rect 12061 1534 12093 1566
rect 12093 1534 12138 1566
rect 12016 1528 12138 1534
rect 11755 1414 11795 1420
rect 11755 1382 11759 1414
rect 11759 1382 11791 1414
rect 11791 1382 11795 1414
rect 11755 1346 11795 1382
rect 11755 1314 11759 1346
rect 11759 1314 11791 1346
rect 11791 1314 11795 1346
rect 11755 1278 11795 1314
rect 11755 1246 11759 1278
rect 11759 1246 11791 1278
rect 11791 1246 11795 1278
rect 11755 1210 11795 1246
rect 11755 1178 11759 1210
rect 11759 1178 11791 1210
rect 11791 1178 11795 1210
rect 11755 1142 11795 1178
rect 11755 1110 11759 1142
rect 11759 1110 11791 1142
rect 11791 1110 11795 1142
rect 11755 1074 11795 1110
rect 11755 1042 11759 1074
rect 11759 1042 11791 1074
rect 11791 1042 11795 1074
rect 11755 1006 11795 1042
rect 11755 974 11759 1006
rect 11759 974 11791 1006
rect 11791 974 11795 1006
rect 11755 938 11795 974
rect 11755 906 11759 938
rect 11759 906 11791 938
rect 11791 906 11795 938
rect 11755 870 11795 906
rect 11755 838 11759 870
rect 11759 838 11791 870
rect 11791 838 11795 870
rect 11755 802 11795 838
rect 11755 770 11759 802
rect 11759 770 11791 802
rect 11791 770 11795 802
rect 11755 734 11795 770
rect 11755 702 11759 734
rect 11759 702 11791 734
rect 11791 702 11795 734
rect 11755 666 11795 702
rect 11755 634 11759 666
rect 11759 634 11791 666
rect 11791 634 11795 666
rect 11755 598 11795 634
rect 11755 566 11759 598
rect 11759 566 11791 598
rect 11791 566 11795 598
rect 11755 560 11795 566
rect 12963 4318 13003 4324
rect 12963 4286 12967 4318
rect 12967 4286 12999 4318
rect 12999 4286 13003 4318
rect 12963 4250 13003 4286
rect 12963 4218 12967 4250
rect 12967 4218 12999 4250
rect 12999 4218 13003 4250
rect 12963 4182 13003 4218
rect 12963 4150 12967 4182
rect 12967 4150 12999 4182
rect 12999 4150 13003 4182
rect 12963 4114 13003 4150
rect 12963 4082 12967 4114
rect 12967 4082 12999 4114
rect 12999 4082 13003 4114
rect 12963 4046 13003 4082
rect 12963 4014 12967 4046
rect 12967 4014 12999 4046
rect 12999 4014 13003 4046
rect 12963 3978 13003 4014
rect 12963 3946 12967 3978
rect 12967 3946 12999 3978
rect 12999 3946 13003 3978
rect 12963 3910 13003 3946
rect 12963 3878 12967 3910
rect 12967 3878 12999 3910
rect 12999 3878 13003 3910
rect 12963 3842 13003 3878
rect 12963 3810 12967 3842
rect 12967 3810 12999 3842
rect 12999 3810 13003 3842
rect 12963 3774 13003 3810
rect 12963 3742 12967 3774
rect 12967 3742 12999 3774
rect 12999 3742 13003 3774
rect 12963 3706 13003 3742
rect 12963 3674 12967 3706
rect 12967 3674 12999 3706
rect 12999 3674 13003 3706
rect 12963 3638 13003 3674
rect 12963 3606 12967 3638
rect 12967 3606 12999 3638
rect 12999 3606 13003 3638
rect 12963 3570 13003 3606
rect 12963 3538 12967 3570
rect 12967 3538 12999 3570
rect 12999 3538 13003 3570
rect 12963 3502 13003 3538
rect 12963 3470 12967 3502
rect 12967 3470 12999 3502
rect 12999 3470 13003 3502
rect 12963 3464 13003 3470
rect 12620 3350 12742 3356
rect 12620 3318 12665 3350
rect 12665 3318 12697 3350
rect 12697 3318 12742 3350
rect 12620 3282 12742 3318
rect 12620 3250 12665 3282
rect 12665 3250 12697 3282
rect 12697 3250 12742 3282
rect 12620 3214 12742 3250
rect 12620 3182 12665 3214
rect 12665 3182 12697 3214
rect 12697 3182 12742 3214
rect 12620 3146 12742 3182
rect 12620 3114 12665 3146
rect 12665 3114 12697 3146
rect 12697 3114 12742 3146
rect 12620 3078 12742 3114
rect 12620 3046 12665 3078
rect 12665 3046 12697 3078
rect 12697 3046 12742 3078
rect 12620 3010 12742 3046
rect 12620 2978 12665 3010
rect 12665 2978 12697 3010
rect 12697 2978 12742 3010
rect 12620 2942 12742 2978
rect 12620 2910 12665 2942
rect 12665 2910 12697 2942
rect 12697 2910 12742 2942
rect 12620 2874 12742 2910
rect 12620 2842 12665 2874
rect 12665 2842 12697 2874
rect 12697 2842 12742 2874
rect 12620 2806 12742 2842
rect 12620 2774 12665 2806
rect 12665 2774 12697 2806
rect 12697 2774 12742 2806
rect 12620 2738 12742 2774
rect 12620 2706 12665 2738
rect 12665 2706 12697 2738
rect 12697 2706 12742 2738
rect 12620 2670 12742 2706
rect 12620 2638 12665 2670
rect 12665 2638 12697 2670
rect 12697 2638 12742 2670
rect 12620 2602 12742 2638
rect 12620 2570 12665 2602
rect 12665 2570 12697 2602
rect 12697 2570 12742 2602
rect 12620 2534 12742 2570
rect 12620 2502 12665 2534
rect 12665 2502 12697 2534
rect 12697 2502 12742 2534
rect 12620 2496 12742 2502
rect 12359 2382 12399 2388
rect 12359 2350 12363 2382
rect 12363 2350 12395 2382
rect 12395 2350 12399 2382
rect 12359 2314 12399 2350
rect 12359 2282 12363 2314
rect 12363 2282 12395 2314
rect 12395 2282 12399 2314
rect 12359 2246 12399 2282
rect 12359 2214 12363 2246
rect 12363 2214 12395 2246
rect 12395 2214 12399 2246
rect 12359 2178 12399 2214
rect 12359 2146 12363 2178
rect 12363 2146 12395 2178
rect 12395 2146 12399 2178
rect 12359 2110 12399 2146
rect 12359 2078 12363 2110
rect 12363 2078 12395 2110
rect 12395 2078 12399 2110
rect 12359 2042 12399 2078
rect 12359 2010 12363 2042
rect 12363 2010 12395 2042
rect 12395 2010 12399 2042
rect 12359 1974 12399 2010
rect 12359 1942 12363 1974
rect 12363 1942 12395 1974
rect 12395 1942 12399 1974
rect 12359 1906 12399 1942
rect 12359 1874 12363 1906
rect 12363 1874 12395 1906
rect 12395 1874 12399 1906
rect 12359 1838 12399 1874
rect 12359 1806 12363 1838
rect 12363 1806 12395 1838
rect 12395 1806 12399 1838
rect 12359 1770 12399 1806
rect 12359 1738 12363 1770
rect 12363 1738 12395 1770
rect 12395 1738 12399 1770
rect 12359 1702 12399 1738
rect 12359 1670 12363 1702
rect 12363 1670 12395 1702
rect 12395 1670 12399 1702
rect 12359 1634 12399 1670
rect 12359 1602 12363 1634
rect 12363 1602 12395 1634
rect 12395 1602 12399 1634
rect 12359 1566 12399 1602
rect 12359 1534 12363 1566
rect 12363 1534 12395 1566
rect 12395 1534 12399 1566
rect 12359 1528 12399 1534
rect 12016 1414 12138 1420
rect 12016 1382 12061 1414
rect 12061 1382 12093 1414
rect 12093 1382 12138 1414
rect 12016 1346 12138 1382
rect 12016 1314 12061 1346
rect 12061 1314 12093 1346
rect 12093 1314 12138 1346
rect 12016 1278 12138 1314
rect 12016 1246 12061 1278
rect 12061 1246 12093 1278
rect 12093 1246 12138 1278
rect 12016 1210 12138 1246
rect 12016 1178 12061 1210
rect 12061 1178 12093 1210
rect 12093 1178 12138 1210
rect 12016 1142 12138 1178
rect 12016 1110 12061 1142
rect 12061 1110 12093 1142
rect 12093 1110 12138 1142
rect 12016 1074 12138 1110
rect 12016 1042 12061 1074
rect 12061 1042 12093 1074
rect 12093 1042 12138 1074
rect 12016 1006 12138 1042
rect 12016 974 12061 1006
rect 12061 974 12093 1006
rect 12093 974 12138 1006
rect 12016 938 12138 974
rect 12016 906 12061 938
rect 12061 906 12093 938
rect 12093 906 12138 938
rect 12016 870 12138 906
rect 12016 838 12061 870
rect 12061 838 12093 870
rect 12093 838 12138 870
rect 12016 802 12138 838
rect 12016 770 12061 802
rect 12061 770 12093 802
rect 12093 770 12138 802
rect 12016 734 12138 770
rect 12016 702 12061 734
rect 12061 702 12093 734
rect 12093 702 12138 734
rect 12016 666 12138 702
rect 12016 634 12061 666
rect 12061 634 12093 666
rect 12093 634 12138 666
rect 12016 598 12138 634
rect 12016 566 12061 598
rect 12061 566 12093 598
rect 12093 566 12138 598
rect 12016 560 12138 566
rect 13224 4318 13346 4324
rect 13224 4286 13269 4318
rect 13269 4286 13301 4318
rect 13301 4286 13346 4318
rect 13224 4250 13346 4286
rect 13224 4218 13269 4250
rect 13269 4218 13301 4250
rect 13301 4218 13346 4250
rect 13224 4182 13346 4218
rect 13224 4150 13269 4182
rect 13269 4150 13301 4182
rect 13301 4150 13346 4182
rect 13224 4114 13346 4150
rect 13224 4082 13269 4114
rect 13269 4082 13301 4114
rect 13301 4082 13346 4114
rect 13224 4046 13346 4082
rect 13224 4014 13269 4046
rect 13269 4014 13301 4046
rect 13301 4014 13346 4046
rect 13224 3978 13346 4014
rect 13224 3946 13269 3978
rect 13269 3946 13301 3978
rect 13301 3946 13346 3978
rect 13224 3910 13346 3946
rect 13224 3878 13269 3910
rect 13269 3878 13301 3910
rect 13301 3878 13346 3910
rect 13224 3842 13346 3878
rect 13224 3810 13269 3842
rect 13269 3810 13301 3842
rect 13301 3810 13346 3842
rect 13224 3774 13346 3810
rect 13224 3742 13269 3774
rect 13269 3742 13301 3774
rect 13301 3742 13346 3774
rect 13224 3706 13346 3742
rect 13224 3674 13269 3706
rect 13269 3674 13301 3706
rect 13301 3674 13346 3706
rect 13224 3638 13346 3674
rect 13224 3606 13269 3638
rect 13269 3606 13301 3638
rect 13301 3606 13346 3638
rect 13224 3570 13346 3606
rect 13224 3538 13269 3570
rect 13269 3538 13301 3570
rect 13301 3538 13346 3570
rect 13224 3502 13346 3538
rect 13224 3470 13269 3502
rect 13269 3470 13301 3502
rect 13301 3470 13346 3502
rect 13224 3464 13346 3470
rect 12963 3350 13003 3356
rect 12963 3318 12967 3350
rect 12967 3318 12999 3350
rect 12999 3318 13003 3350
rect 12963 3282 13003 3318
rect 12963 3250 12967 3282
rect 12967 3250 12999 3282
rect 12999 3250 13003 3282
rect 12963 3214 13003 3250
rect 12963 3182 12967 3214
rect 12967 3182 12999 3214
rect 12999 3182 13003 3214
rect 12963 3146 13003 3182
rect 12963 3114 12967 3146
rect 12967 3114 12999 3146
rect 12999 3114 13003 3146
rect 12963 3078 13003 3114
rect 12963 3046 12967 3078
rect 12967 3046 12999 3078
rect 12999 3046 13003 3078
rect 12963 3010 13003 3046
rect 12963 2978 12967 3010
rect 12967 2978 12999 3010
rect 12999 2978 13003 3010
rect 12963 2942 13003 2978
rect 12963 2910 12967 2942
rect 12967 2910 12999 2942
rect 12999 2910 13003 2942
rect 12963 2874 13003 2910
rect 12963 2842 12967 2874
rect 12967 2842 12999 2874
rect 12999 2842 13003 2874
rect 12963 2806 13003 2842
rect 12963 2774 12967 2806
rect 12967 2774 12999 2806
rect 12999 2774 13003 2806
rect 12963 2738 13003 2774
rect 12963 2706 12967 2738
rect 12967 2706 12999 2738
rect 12999 2706 13003 2738
rect 12963 2670 13003 2706
rect 12963 2638 12967 2670
rect 12967 2638 12999 2670
rect 12999 2638 13003 2670
rect 12963 2602 13003 2638
rect 12963 2570 12967 2602
rect 12967 2570 12999 2602
rect 12999 2570 13003 2602
rect 12963 2534 13003 2570
rect 12963 2502 12967 2534
rect 12967 2502 12999 2534
rect 12999 2502 13003 2534
rect 12963 2496 13003 2502
rect 12620 2382 12742 2388
rect 12620 2350 12665 2382
rect 12665 2350 12697 2382
rect 12697 2350 12742 2382
rect 12620 2314 12742 2350
rect 12620 2282 12665 2314
rect 12665 2282 12697 2314
rect 12697 2282 12742 2314
rect 12620 2246 12742 2282
rect 12620 2214 12665 2246
rect 12665 2214 12697 2246
rect 12697 2214 12742 2246
rect 12620 2178 12742 2214
rect 12620 2146 12665 2178
rect 12665 2146 12697 2178
rect 12697 2146 12742 2178
rect 12620 2110 12742 2146
rect 12620 2078 12665 2110
rect 12665 2078 12697 2110
rect 12697 2078 12742 2110
rect 12620 2042 12742 2078
rect 12620 2010 12665 2042
rect 12665 2010 12697 2042
rect 12697 2010 12742 2042
rect 12620 1974 12742 2010
rect 12620 1942 12665 1974
rect 12665 1942 12697 1974
rect 12697 1942 12742 1974
rect 12620 1906 12742 1942
rect 12620 1874 12665 1906
rect 12665 1874 12697 1906
rect 12697 1874 12742 1906
rect 12620 1838 12742 1874
rect 12620 1806 12665 1838
rect 12665 1806 12697 1838
rect 12697 1806 12742 1838
rect 12620 1770 12742 1806
rect 12620 1738 12665 1770
rect 12665 1738 12697 1770
rect 12697 1738 12742 1770
rect 12620 1702 12742 1738
rect 12620 1670 12665 1702
rect 12665 1670 12697 1702
rect 12697 1670 12742 1702
rect 12620 1634 12742 1670
rect 12620 1602 12665 1634
rect 12665 1602 12697 1634
rect 12697 1602 12742 1634
rect 12620 1566 12742 1602
rect 12620 1534 12665 1566
rect 12665 1534 12697 1566
rect 12697 1534 12742 1566
rect 12620 1528 12742 1534
rect 12359 1414 12399 1420
rect 12359 1382 12363 1414
rect 12363 1382 12395 1414
rect 12395 1382 12399 1414
rect 12359 1346 12399 1382
rect 12359 1314 12363 1346
rect 12363 1314 12395 1346
rect 12395 1314 12399 1346
rect 12359 1278 12399 1314
rect 12359 1246 12363 1278
rect 12363 1246 12395 1278
rect 12395 1246 12399 1278
rect 12359 1210 12399 1246
rect 12359 1178 12363 1210
rect 12363 1178 12395 1210
rect 12395 1178 12399 1210
rect 12359 1142 12399 1178
rect 12359 1110 12363 1142
rect 12363 1110 12395 1142
rect 12395 1110 12399 1142
rect 12359 1074 12399 1110
rect 12359 1042 12363 1074
rect 12363 1042 12395 1074
rect 12395 1042 12399 1074
rect 12359 1006 12399 1042
rect 12359 974 12363 1006
rect 12363 974 12395 1006
rect 12395 974 12399 1006
rect 12359 938 12399 974
rect 12359 906 12363 938
rect 12363 906 12395 938
rect 12395 906 12399 938
rect 12359 870 12399 906
rect 12359 838 12363 870
rect 12363 838 12395 870
rect 12395 838 12399 870
rect 12359 802 12399 838
rect 12359 770 12363 802
rect 12363 770 12395 802
rect 12395 770 12399 802
rect 12359 734 12399 770
rect 12359 702 12363 734
rect 12363 702 12395 734
rect 12395 702 12399 734
rect 12359 666 12399 702
rect 12359 634 12363 666
rect 12363 634 12395 666
rect 12395 634 12399 666
rect 12359 598 12399 634
rect 12359 566 12363 598
rect 12363 566 12395 598
rect 12395 566 12399 598
rect 12359 560 12399 566
rect 13567 4318 13607 4324
rect 13567 4286 13571 4318
rect 13571 4286 13603 4318
rect 13603 4286 13607 4318
rect 13567 4250 13607 4286
rect 13567 4218 13571 4250
rect 13571 4218 13603 4250
rect 13603 4218 13607 4250
rect 13567 4182 13607 4218
rect 13567 4150 13571 4182
rect 13571 4150 13603 4182
rect 13603 4150 13607 4182
rect 13567 4114 13607 4150
rect 13567 4082 13571 4114
rect 13571 4082 13603 4114
rect 13603 4082 13607 4114
rect 13567 4046 13607 4082
rect 13567 4014 13571 4046
rect 13571 4014 13603 4046
rect 13603 4014 13607 4046
rect 13567 3978 13607 4014
rect 13567 3946 13571 3978
rect 13571 3946 13603 3978
rect 13603 3946 13607 3978
rect 13567 3910 13607 3946
rect 13567 3878 13571 3910
rect 13571 3878 13603 3910
rect 13603 3878 13607 3910
rect 13567 3842 13607 3878
rect 13567 3810 13571 3842
rect 13571 3810 13603 3842
rect 13603 3810 13607 3842
rect 13567 3774 13607 3810
rect 13567 3742 13571 3774
rect 13571 3742 13603 3774
rect 13603 3742 13607 3774
rect 13567 3706 13607 3742
rect 13567 3674 13571 3706
rect 13571 3674 13603 3706
rect 13603 3674 13607 3706
rect 13567 3638 13607 3674
rect 13567 3606 13571 3638
rect 13571 3606 13603 3638
rect 13603 3606 13607 3638
rect 13567 3570 13607 3606
rect 13567 3538 13571 3570
rect 13571 3538 13603 3570
rect 13603 3538 13607 3570
rect 13567 3502 13607 3538
rect 13567 3470 13571 3502
rect 13571 3470 13603 3502
rect 13603 3470 13607 3502
rect 13567 3464 13607 3470
rect 13224 3350 13346 3356
rect 13224 3318 13269 3350
rect 13269 3318 13301 3350
rect 13301 3318 13346 3350
rect 13224 3282 13346 3318
rect 13224 3250 13269 3282
rect 13269 3250 13301 3282
rect 13301 3250 13346 3282
rect 13224 3214 13346 3250
rect 13224 3182 13269 3214
rect 13269 3182 13301 3214
rect 13301 3182 13346 3214
rect 13224 3146 13346 3182
rect 13224 3114 13269 3146
rect 13269 3114 13301 3146
rect 13301 3114 13346 3146
rect 13224 3078 13346 3114
rect 13224 3046 13269 3078
rect 13269 3046 13301 3078
rect 13301 3046 13346 3078
rect 13224 3010 13346 3046
rect 13224 2978 13269 3010
rect 13269 2978 13301 3010
rect 13301 2978 13346 3010
rect 13224 2942 13346 2978
rect 13224 2910 13269 2942
rect 13269 2910 13301 2942
rect 13301 2910 13346 2942
rect 13224 2874 13346 2910
rect 13224 2842 13269 2874
rect 13269 2842 13301 2874
rect 13301 2842 13346 2874
rect 13224 2806 13346 2842
rect 13224 2774 13269 2806
rect 13269 2774 13301 2806
rect 13301 2774 13346 2806
rect 13224 2738 13346 2774
rect 13224 2706 13269 2738
rect 13269 2706 13301 2738
rect 13301 2706 13346 2738
rect 13224 2670 13346 2706
rect 13224 2638 13269 2670
rect 13269 2638 13301 2670
rect 13301 2638 13346 2670
rect 13224 2602 13346 2638
rect 13224 2570 13269 2602
rect 13269 2570 13301 2602
rect 13301 2570 13346 2602
rect 13224 2534 13346 2570
rect 13224 2502 13269 2534
rect 13269 2502 13301 2534
rect 13301 2502 13346 2534
rect 13224 2496 13346 2502
rect 12963 2382 13003 2388
rect 12963 2350 12967 2382
rect 12967 2350 12999 2382
rect 12999 2350 13003 2382
rect 12963 2314 13003 2350
rect 12963 2282 12967 2314
rect 12967 2282 12999 2314
rect 12999 2282 13003 2314
rect 12963 2246 13003 2282
rect 12963 2214 12967 2246
rect 12967 2214 12999 2246
rect 12999 2214 13003 2246
rect 12963 2178 13003 2214
rect 12963 2146 12967 2178
rect 12967 2146 12999 2178
rect 12999 2146 13003 2178
rect 12963 2110 13003 2146
rect 12963 2078 12967 2110
rect 12967 2078 12999 2110
rect 12999 2078 13003 2110
rect 12963 2042 13003 2078
rect 12963 2010 12967 2042
rect 12967 2010 12999 2042
rect 12999 2010 13003 2042
rect 12963 1974 13003 2010
rect 12963 1942 12967 1974
rect 12967 1942 12999 1974
rect 12999 1942 13003 1974
rect 12963 1906 13003 1942
rect 12963 1874 12967 1906
rect 12967 1874 12999 1906
rect 12999 1874 13003 1906
rect 12963 1838 13003 1874
rect 12963 1806 12967 1838
rect 12967 1806 12999 1838
rect 12999 1806 13003 1838
rect 12963 1770 13003 1806
rect 12963 1738 12967 1770
rect 12967 1738 12999 1770
rect 12999 1738 13003 1770
rect 12963 1702 13003 1738
rect 12963 1670 12967 1702
rect 12967 1670 12999 1702
rect 12999 1670 13003 1702
rect 12963 1634 13003 1670
rect 12963 1602 12967 1634
rect 12967 1602 12999 1634
rect 12999 1602 13003 1634
rect 12963 1566 13003 1602
rect 12963 1534 12967 1566
rect 12967 1534 12999 1566
rect 12999 1534 13003 1566
rect 12963 1528 13003 1534
rect 12620 1414 12742 1420
rect 12620 1382 12665 1414
rect 12665 1382 12697 1414
rect 12697 1382 12742 1414
rect 12620 1346 12742 1382
rect 12620 1314 12665 1346
rect 12665 1314 12697 1346
rect 12697 1314 12742 1346
rect 12620 1278 12742 1314
rect 12620 1246 12665 1278
rect 12665 1246 12697 1278
rect 12697 1246 12742 1278
rect 12620 1210 12742 1246
rect 12620 1178 12665 1210
rect 12665 1178 12697 1210
rect 12697 1178 12742 1210
rect 12620 1142 12742 1178
rect 12620 1110 12665 1142
rect 12665 1110 12697 1142
rect 12697 1110 12742 1142
rect 12620 1074 12742 1110
rect 12620 1042 12665 1074
rect 12665 1042 12697 1074
rect 12697 1042 12742 1074
rect 12620 1006 12742 1042
rect 12620 974 12665 1006
rect 12665 974 12697 1006
rect 12697 974 12742 1006
rect 12620 938 12742 974
rect 12620 906 12665 938
rect 12665 906 12697 938
rect 12697 906 12742 938
rect 12620 870 12742 906
rect 12620 838 12665 870
rect 12665 838 12697 870
rect 12697 838 12742 870
rect 12620 802 12742 838
rect 12620 770 12665 802
rect 12665 770 12697 802
rect 12697 770 12742 802
rect 12620 734 12742 770
rect 12620 702 12665 734
rect 12665 702 12697 734
rect 12697 702 12742 734
rect 12620 666 12742 702
rect 12620 634 12665 666
rect 12665 634 12697 666
rect 12697 634 12742 666
rect 12620 598 12742 634
rect 12620 566 12665 598
rect 12665 566 12697 598
rect 12697 566 12742 598
rect 12620 560 12742 566
rect 13828 4318 13950 4324
rect 13828 4286 13873 4318
rect 13873 4286 13905 4318
rect 13905 4286 13950 4318
rect 13828 4250 13950 4286
rect 13828 4218 13873 4250
rect 13873 4218 13905 4250
rect 13905 4218 13950 4250
rect 13828 4182 13950 4218
rect 13828 4150 13873 4182
rect 13873 4150 13905 4182
rect 13905 4150 13950 4182
rect 13828 4114 13950 4150
rect 13828 4082 13873 4114
rect 13873 4082 13905 4114
rect 13905 4082 13950 4114
rect 13828 4046 13950 4082
rect 13828 4014 13873 4046
rect 13873 4014 13905 4046
rect 13905 4014 13950 4046
rect 13828 3978 13950 4014
rect 13828 3946 13873 3978
rect 13873 3946 13905 3978
rect 13905 3946 13950 3978
rect 13828 3910 13950 3946
rect 13828 3878 13873 3910
rect 13873 3878 13905 3910
rect 13905 3878 13950 3910
rect 13828 3842 13950 3878
rect 13828 3810 13873 3842
rect 13873 3810 13905 3842
rect 13905 3810 13950 3842
rect 13828 3774 13950 3810
rect 13828 3742 13873 3774
rect 13873 3742 13905 3774
rect 13905 3742 13950 3774
rect 13828 3706 13950 3742
rect 13828 3674 13873 3706
rect 13873 3674 13905 3706
rect 13905 3674 13950 3706
rect 13828 3638 13950 3674
rect 13828 3606 13873 3638
rect 13873 3606 13905 3638
rect 13905 3606 13950 3638
rect 13828 3570 13950 3606
rect 13828 3538 13873 3570
rect 13873 3538 13905 3570
rect 13905 3538 13950 3570
rect 13828 3502 13950 3538
rect 13828 3470 13873 3502
rect 13873 3470 13905 3502
rect 13905 3470 13950 3502
rect 13828 3464 13950 3470
rect 13567 3350 13607 3356
rect 13567 3318 13571 3350
rect 13571 3318 13603 3350
rect 13603 3318 13607 3350
rect 13567 3282 13607 3318
rect 13567 3250 13571 3282
rect 13571 3250 13603 3282
rect 13603 3250 13607 3282
rect 13567 3214 13607 3250
rect 13567 3182 13571 3214
rect 13571 3182 13603 3214
rect 13603 3182 13607 3214
rect 13567 3146 13607 3182
rect 13567 3114 13571 3146
rect 13571 3114 13603 3146
rect 13603 3114 13607 3146
rect 13567 3078 13607 3114
rect 13567 3046 13571 3078
rect 13571 3046 13603 3078
rect 13603 3046 13607 3078
rect 13567 3010 13607 3046
rect 13567 2978 13571 3010
rect 13571 2978 13603 3010
rect 13603 2978 13607 3010
rect 13567 2942 13607 2978
rect 13567 2910 13571 2942
rect 13571 2910 13603 2942
rect 13603 2910 13607 2942
rect 13567 2874 13607 2910
rect 13567 2842 13571 2874
rect 13571 2842 13603 2874
rect 13603 2842 13607 2874
rect 13567 2806 13607 2842
rect 13567 2774 13571 2806
rect 13571 2774 13603 2806
rect 13603 2774 13607 2806
rect 13567 2738 13607 2774
rect 13567 2706 13571 2738
rect 13571 2706 13603 2738
rect 13603 2706 13607 2738
rect 13567 2670 13607 2706
rect 13567 2638 13571 2670
rect 13571 2638 13603 2670
rect 13603 2638 13607 2670
rect 13567 2602 13607 2638
rect 13567 2570 13571 2602
rect 13571 2570 13603 2602
rect 13603 2570 13607 2602
rect 13567 2534 13607 2570
rect 13567 2502 13571 2534
rect 13571 2502 13603 2534
rect 13603 2502 13607 2534
rect 13567 2496 13607 2502
rect 13224 2382 13346 2388
rect 13224 2350 13269 2382
rect 13269 2350 13301 2382
rect 13301 2350 13346 2382
rect 13224 2314 13346 2350
rect 13224 2282 13269 2314
rect 13269 2282 13301 2314
rect 13301 2282 13346 2314
rect 13224 2246 13346 2282
rect 13224 2214 13269 2246
rect 13269 2214 13301 2246
rect 13301 2214 13346 2246
rect 13224 2178 13346 2214
rect 13224 2146 13269 2178
rect 13269 2146 13301 2178
rect 13301 2146 13346 2178
rect 13224 2110 13346 2146
rect 13224 2078 13269 2110
rect 13269 2078 13301 2110
rect 13301 2078 13346 2110
rect 13224 2042 13346 2078
rect 13224 2010 13269 2042
rect 13269 2010 13301 2042
rect 13301 2010 13346 2042
rect 13224 1974 13346 2010
rect 13224 1942 13269 1974
rect 13269 1942 13301 1974
rect 13301 1942 13346 1974
rect 13224 1906 13346 1942
rect 13224 1874 13269 1906
rect 13269 1874 13301 1906
rect 13301 1874 13346 1906
rect 13224 1838 13346 1874
rect 13224 1806 13269 1838
rect 13269 1806 13301 1838
rect 13301 1806 13346 1838
rect 13224 1770 13346 1806
rect 13224 1738 13269 1770
rect 13269 1738 13301 1770
rect 13301 1738 13346 1770
rect 13224 1702 13346 1738
rect 13224 1670 13269 1702
rect 13269 1670 13301 1702
rect 13301 1670 13346 1702
rect 13224 1634 13346 1670
rect 13224 1602 13269 1634
rect 13269 1602 13301 1634
rect 13301 1602 13346 1634
rect 13224 1566 13346 1602
rect 13224 1534 13269 1566
rect 13269 1534 13301 1566
rect 13301 1534 13346 1566
rect 13224 1528 13346 1534
rect 12963 1414 13003 1420
rect 12963 1382 12967 1414
rect 12967 1382 12999 1414
rect 12999 1382 13003 1414
rect 12963 1346 13003 1382
rect 12963 1314 12967 1346
rect 12967 1314 12999 1346
rect 12999 1314 13003 1346
rect 12963 1278 13003 1314
rect 12963 1246 12967 1278
rect 12967 1246 12999 1278
rect 12999 1246 13003 1278
rect 12963 1210 13003 1246
rect 12963 1178 12967 1210
rect 12967 1178 12999 1210
rect 12999 1178 13003 1210
rect 12963 1142 13003 1178
rect 12963 1110 12967 1142
rect 12967 1110 12999 1142
rect 12999 1110 13003 1142
rect 12963 1074 13003 1110
rect 12963 1042 12967 1074
rect 12967 1042 12999 1074
rect 12999 1042 13003 1074
rect 12963 1006 13003 1042
rect 12963 974 12967 1006
rect 12967 974 12999 1006
rect 12999 974 13003 1006
rect 12963 938 13003 974
rect 12963 906 12967 938
rect 12967 906 12999 938
rect 12999 906 13003 938
rect 12963 870 13003 906
rect 12963 838 12967 870
rect 12967 838 12999 870
rect 12999 838 13003 870
rect 12963 802 13003 838
rect 12963 770 12967 802
rect 12967 770 12999 802
rect 12999 770 13003 802
rect 12963 734 13003 770
rect 12963 702 12967 734
rect 12967 702 12999 734
rect 12999 702 13003 734
rect 12963 666 13003 702
rect 12963 634 12967 666
rect 12967 634 12999 666
rect 12999 634 13003 666
rect 12963 598 13003 634
rect 12963 566 12967 598
rect 12967 566 12999 598
rect 12999 566 13003 598
rect 12963 560 13003 566
rect 14171 4318 14211 4324
rect 14171 4286 14175 4318
rect 14175 4286 14207 4318
rect 14207 4286 14211 4318
rect 14171 4250 14211 4286
rect 14171 4218 14175 4250
rect 14175 4218 14207 4250
rect 14207 4218 14211 4250
rect 14171 4182 14211 4218
rect 14171 4150 14175 4182
rect 14175 4150 14207 4182
rect 14207 4150 14211 4182
rect 14171 4114 14211 4150
rect 14171 4082 14175 4114
rect 14175 4082 14207 4114
rect 14207 4082 14211 4114
rect 14171 4046 14211 4082
rect 14171 4014 14175 4046
rect 14175 4014 14207 4046
rect 14207 4014 14211 4046
rect 14171 3978 14211 4014
rect 14171 3946 14175 3978
rect 14175 3946 14207 3978
rect 14207 3946 14211 3978
rect 14171 3910 14211 3946
rect 14171 3878 14175 3910
rect 14175 3878 14207 3910
rect 14207 3878 14211 3910
rect 14171 3842 14211 3878
rect 14171 3810 14175 3842
rect 14175 3810 14207 3842
rect 14207 3810 14211 3842
rect 14171 3774 14211 3810
rect 14171 3742 14175 3774
rect 14175 3742 14207 3774
rect 14207 3742 14211 3774
rect 14171 3706 14211 3742
rect 14171 3674 14175 3706
rect 14175 3674 14207 3706
rect 14207 3674 14211 3706
rect 14171 3638 14211 3674
rect 14171 3606 14175 3638
rect 14175 3606 14207 3638
rect 14207 3606 14211 3638
rect 14171 3570 14211 3606
rect 14171 3538 14175 3570
rect 14175 3538 14207 3570
rect 14207 3538 14211 3570
rect 14171 3502 14211 3538
rect 14171 3470 14175 3502
rect 14175 3470 14207 3502
rect 14207 3470 14211 3502
rect 14171 3464 14211 3470
rect 13828 3350 13950 3356
rect 13828 3318 13873 3350
rect 13873 3318 13905 3350
rect 13905 3318 13950 3350
rect 13828 3282 13950 3318
rect 13828 3250 13873 3282
rect 13873 3250 13905 3282
rect 13905 3250 13950 3282
rect 13828 3214 13950 3250
rect 13828 3182 13873 3214
rect 13873 3182 13905 3214
rect 13905 3182 13950 3214
rect 13828 3146 13950 3182
rect 13828 3114 13873 3146
rect 13873 3114 13905 3146
rect 13905 3114 13950 3146
rect 13828 3078 13950 3114
rect 13828 3046 13873 3078
rect 13873 3046 13905 3078
rect 13905 3046 13950 3078
rect 13828 3010 13950 3046
rect 13828 2978 13873 3010
rect 13873 2978 13905 3010
rect 13905 2978 13950 3010
rect 13828 2942 13950 2978
rect 13828 2910 13873 2942
rect 13873 2910 13905 2942
rect 13905 2910 13950 2942
rect 13828 2874 13950 2910
rect 13828 2842 13873 2874
rect 13873 2842 13905 2874
rect 13905 2842 13950 2874
rect 13828 2806 13950 2842
rect 13828 2774 13873 2806
rect 13873 2774 13905 2806
rect 13905 2774 13950 2806
rect 13828 2738 13950 2774
rect 13828 2706 13873 2738
rect 13873 2706 13905 2738
rect 13905 2706 13950 2738
rect 13828 2670 13950 2706
rect 13828 2638 13873 2670
rect 13873 2638 13905 2670
rect 13905 2638 13950 2670
rect 13828 2602 13950 2638
rect 13828 2570 13873 2602
rect 13873 2570 13905 2602
rect 13905 2570 13950 2602
rect 13828 2534 13950 2570
rect 13828 2502 13873 2534
rect 13873 2502 13905 2534
rect 13905 2502 13950 2534
rect 13828 2496 13950 2502
rect 13567 2382 13607 2388
rect 13567 2350 13571 2382
rect 13571 2350 13603 2382
rect 13603 2350 13607 2382
rect 13567 2314 13607 2350
rect 13567 2282 13571 2314
rect 13571 2282 13603 2314
rect 13603 2282 13607 2314
rect 13567 2246 13607 2282
rect 13567 2214 13571 2246
rect 13571 2214 13603 2246
rect 13603 2214 13607 2246
rect 13567 2178 13607 2214
rect 13567 2146 13571 2178
rect 13571 2146 13603 2178
rect 13603 2146 13607 2178
rect 13567 2110 13607 2146
rect 13567 2078 13571 2110
rect 13571 2078 13603 2110
rect 13603 2078 13607 2110
rect 13567 2042 13607 2078
rect 13567 2010 13571 2042
rect 13571 2010 13603 2042
rect 13603 2010 13607 2042
rect 13567 1974 13607 2010
rect 13567 1942 13571 1974
rect 13571 1942 13603 1974
rect 13603 1942 13607 1974
rect 13567 1906 13607 1942
rect 13567 1874 13571 1906
rect 13571 1874 13603 1906
rect 13603 1874 13607 1906
rect 13567 1838 13607 1874
rect 13567 1806 13571 1838
rect 13571 1806 13603 1838
rect 13603 1806 13607 1838
rect 13567 1770 13607 1806
rect 13567 1738 13571 1770
rect 13571 1738 13603 1770
rect 13603 1738 13607 1770
rect 13567 1702 13607 1738
rect 13567 1670 13571 1702
rect 13571 1670 13603 1702
rect 13603 1670 13607 1702
rect 13567 1634 13607 1670
rect 13567 1602 13571 1634
rect 13571 1602 13603 1634
rect 13603 1602 13607 1634
rect 13567 1566 13607 1602
rect 13567 1534 13571 1566
rect 13571 1534 13603 1566
rect 13603 1534 13607 1566
rect 13567 1528 13607 1534
rect 13224 1414 13346 1420
rect 13224 1382 13269 1414
rect 13269 1382 13301 1414
rect 13301 1382 13346 1414
rect 13224 1346 13346 1382
rect 13224 1314 13269 1346
rect 13269 1314 13301 1346
rect 13301 1314 13346 1346
rect 13224 1278 13346 1314
rect 13224 1246 13269 1278
rect 13269 1246 13301 1278
rect 13301 1246 13346 1278
rect 13224 1210 13346 1246
rect 13224 1178 13269 1210
rect 13269 1178 13301 1210
rect 13301 1178 13346 1210
rect 13224 1142 13346 1178
rect 13224 1110 13269 1142
rect 13269 1110 13301 1142
rect 13301 1110 13346 1142
rect 13224 1074 13346 1110
rect 13224 1042 13269 1074
rect 13269 1042 13301 1074
rect 13301 1042 13346 1074
rect 13224 1006 13346 1042
rect 13224 974 13269 1006
rect 13269 974 13301 1006
rect 13301 974 13346 1006
rect 13224 938 13346 974
rect 13224 906 13269 938
rect 13269 906 13301 938
rect 13301 906 13346 938
rect 13224 870 13346 906
rect 13224 838 13269 870
rect 13269 838 13301 870
rect 13301 838 13346 870
rect 13224 802 13346 838
rect 13224 770 13269 802
rect 13269 770 13301 802
rect 13301 770 13346 802
rect 13224 734 13346 770
rect 13224 702 13269 734
rect 13269 702 13301 734
rect 13301 702 13346 734
rect 13224 666 13346 702
rect 13224 634 13269 666
rect 13269 634 13301 666
rect 13301 634 13346 666
rect 13224 598 13346 634
rect 13224 566 13269 598
rect 13269 566 13301 598
rect 13301 566 13346 598
rect 13224 560 13346 566
rect 14432 4318 14554 4324
rect 14432 4286 14477 4318
rect 14477 4286 14509 4318
rect 14509 4286 14554 4318
rect 14432 4250 14554 4286
rect 14432 4218 14477 4250
rect 14477 4218 14509 4250
rect 14509 4218 14554 4250
rect 14432 4182 14554 4218
rect 14432 4150 14477 4182
rect 14477 4150 14509 4182
rect 14509 4150 14554 4182
rect 14432 4114 14554 4150
rect 14432 4082 14477 4114
rect 14477 4082 14509 4114
rect 14509 4082 14554 4114
rect 14432 4046 14554 4082
rect 14432 4014 14477 4046
rect 14477 4014 14509 4046
rect 14509 4014 14554 4046
rect 14432 3978 14554 4014
rect 14432 3946 14477 3978
rect 14477 3946 14509 3978
rect 14509 3946 14554 3978
rect 14432 3910 14554 3946
rect 14432 3878 14477 3910
rect 14477 3878 14509 3910
rect 14509 3878 14554 3910
rect 14432 3842 14554 3878
rect 14432 3810 14477 3842
rect 14477 3810 14509 3842
rect 14509 3810 14554 3842
rect 14432 3774 14554 3810
rect 14432 3742 14477 3774
rect 14477 3742 14509 3774
rect 14509 3742 14554 3774
rect 14432 3706 14554 3742
rect 14432 3674 14477 3706
rect 14477 3674 14509 3706
rect 14509 3674 14554 3706
rect 14432 3638 14554 3674
rect 14432 3606 14477 3638
rect 14477 3606 14509 3638
rect 14509 3606 14554 3638
rect 14432 3570 14554 3606
rect 14432 3538 14477 3570
rect 14477 3538 14509 3570
rect 14509 3538 14554 3570
rect 14432 3502 14554 3538
rect 14432 3470 14477 3502
rect 14477 3470 14509 3502
rect 14509 3470 14554 3502
rect 14432 3464 14554 3470
rect 14171 3350 14211 3356
rect 14171 3318 14175 3350
rect 14175 3318 14207 3350
rect 14207 3318 14211 3350
rect 14171 3282 14211 3318
rect 14171 3250 14175 3282
rect 14175 3250 14207 3282
rect 14207 3250 14211 3282
rect 14171 3214 14211 3250
rect 14171 3182 14175 3214
rect 14175 3182 14207 3214
rect 14207 3182 14211 3214
rect 14171 3146 14211 3182
rect 14171 3114 14175 3146
rect 14175 3114 14207 3146
rect 14207 3114 14211 3146
rect 14171 3078 14211 3114
rect 14171 3046 14175 3078
rect 14175 3046 14207 3078
rect 14207 3046 14211 3078
rect 14171 3010 14211 3046
rect 14171 2978 14175 3010
rect 14175 2978 14207 3010
rect 14207 2978 14211 3010
rect 14171 2942 14211 2978
rect 14171 2910 14175 2942
rect 14175 2910 14207 2942
rect 14207 2910 14211 2942
rect 14171 2874 14211 2910
rect 14171 2842 14175 2874
rect 14175 2842 14207 2874
rect 14207 2842 14211 2874
rect 14171 2806 14211 2842
rect 14171 2774 14175 2806
rect 14175 2774 14207 2806
rect 14207 2774 14211 2806
rect 14171 2738 14211 2774
rect 14171 2706 14175 2738
rect 14175 2706 14207 2738
rect 14207 2706 14211 2738
rect 14171 2670 14211 2706
rect 14171 2638 14175 2670
rect 14175 2638 14207 2670
rect 14207 2638 14211 2670
rect 14171 2602 14211 2638
rect 14171 2570 14175 2602
rect 14175 2570 14207 2602
rect 14207 2570 14211 2602
rect 14171 2534 14211 2570
rect 14171 2502 14175 2534
rect 14175 2502 14207 2534
rect 14207 2502 14211 2534
rect 14171 2496 14211 2502
rect 13828 2382 13950 2388
rect 13828 2350 13873 2382
rect 13873 2350 13905 2382
rect 13905 2350 13950 2382
rect 13828 2314 13950 2350
rect 13828 2282 13873 2314
rect 13873 2282 13905 2314
rect 13905 2282 13950 2314
rect 13828 2246 13950 2282
rect 13828 2214 13873 2246
rect 13873 2214 13905 2246
rect 13905 2214 13950 2246
rect 13828 2178 13950 2214
rect 13828 2146 13873 2178
rect 13873 2146 13905 2178
rect 13905 2146 13950 2178
rect 13828 2110 13950 2146
rect 13828 2078 13873 2110
rect 13873 2078 13905 2110
rect 13905 2078 13950 2110
rect 13828 2042 13950 2078
rect 13828 2010 13873 2042
rect 13873 2010 13905 2042
rect 13905 2010 13950 2042
rect 13828 1974 13950 2010
rect 13828 1942 13873 1974
rect 13873 1942 13905 1974
rect 13905 1942 13950 1974
rect 13828 1906 13950 1942
rect 13828 1874 13873 1906
rect 13873 1874 13905 1906
rect 13905 1874 13950 1906
rect 13828 1838 13950 1874
rect 13828 1806 13873 1838
rect 13873 1806 13905 1838
rect 13905 1806 13950 1838
rect 13828 1770 13950 1806
rect 13828 1738 13873 1770
rect 13873 1738 13905 1770
rect 13905 1738 13950 1770
rect 13828 1702 13950 1738
rect 13828 1670 13873 1702
rect 13873 1670 13905 1702
rect 13905 1670 13950 1702
rect 13828 1634 13950 1670
rect 13828 1602 13873 1634
rect 13873 1602 13905 1634
rect 13905 1602 13950 1634
rect 13828 1566 13950 1602
rect 13828 1534 13873 1566
rect 13873 1534 13905 1566
rect 13905 1534 13950 1566
rect 13828 1528 13950 1534
rect 13567 1414 13607 1420
rect 13567 1382 13571 1414
rect 13571 1382 13603 1414
rect 13603 1382 13607 1414
rect 13567 1346 13607 1382
rect 13567 1314 13571 1346
rect 13571 1314 13603 1346
rect 13603 1314 13607 1346
rect 13567 1278 13607 1314
rect 13567 1246 13571 1278
rect 13571 1246 13603 1278
rect 13603 1246 13607 1278
rect 13567 1210 13607 1246
rect 13567 1178 13571 1210
rect 13571 1178 13603 1210
rect 13603 1178 13607 1210
rect 13567 1142 13607 1178
rect 13567 1110 13571 1142
rect 13571 1110 13603 1142
rect 13603 1110 13607 1142
rect 13567 1074 13607 1110
rect 13567 1042 13571 1074
rect 13571 1042 13603 1074
rect 13603 1042 13607 1074
rect 13567 1006 13607 1042
rect 13567 974 13571 1006
rect 13571 974 13603 1006
rect 13603 974 13607 1006
rect 13567 938 13607 974
rect 13567 906 13571 938
rect 13571 906 13603 938
rect 13603 906 13607 938
rect 13567 870 13607 906
rect 13567 838 13571 870
rect 13571 838 13603 870
rect 13603 838 13607 870
rect 13567 802 13607 838
rect 13567 770 13571 802
rect 13571 770 13603 802
rect 13603 770 13607 802
rect 13567 734 13607 770
rect 13567 702 13571 734
rect 13571 702 13603 734
rect 13603 702 13607 734
rect 13567 666 13607 702
rect 13567 634 13571 666
rect 13571 634 13603 666
rect 13603 634 13607 666
rect 13567 598 13607 634
rect 13567 566 13571 598
rect 13571 566 13603 598
rect 13603 566 13607 598
rect 13567 560 13607 566
rect 14432 3350 14554 3356
rect 14432 3318 14477 3350
rect 14477 3318 14509 3350
rect 14509 3318 14554 3350
rect 14432 3282 14554 3318
rect 14432 3250 14477 3282
rect 14477 3250 14509 3282
rect 14509 3250 14554 3282
rect 14432 3214 14554 3250
rect 14432 3182 14477 3214
rect 14477 3182 14509 3214
rect 14509 3182 14554 3214
rect 14432 3146 14554 3182
rect 14432 3114 14477 3146
rect 14477 3114 14509 3146
rect 14509 3114 14554 3146
rect 14432 3078 14554 3114
rect 14432 3046 14477 3078
rect 14477 3046 14509 3078
rect 14509 3046 14554 3078
rect 14432 3010 14554 3046
rect 14432 2978 14477 3010
rect 14477 2978 14509 3010
rect 14509 2978 14554 3010
rect 14432 2942 14554 2978
rect 14432 2910 14477 2942
rect 14477 2910 14509 2942
rect 14509 2910 14554 2942
rect 14432 2874 14554 2910
rect 14432 2842 14477 2874
rect 14477 2842 14509 2874
rect 14509 2842 14554 2874
rect 14432 2806 14554 2842
rect 14432 2774 14477 2806
rect 14477 2774 14509 2806
rect 14509 2774 14554 2806
rect 14432 2738 14554 2774
rect 14432 2706 14477 2738
rect 14477 2706 14509 2738
rect 14509 2706 14554 2738
rect 14432 2670 14554 2706
rect 14432 2638 14477 2670
rect 14477 2638 14509 2670
rect 14509 2638 14554 2670
rect 14432 2602 14554 2638
rect 14432 2570 14477 2602
rect 14477 2570 14509 2602
rect 14509 2570 14554 2602
rect 14432 2534 14554 2570
rect 14432 2502 14477 2534
rect 14477 2502 14509 2534
rect 14509 2502 14554 2534
rect 14432 2496 14554 2502
rect 14171 2382 14211 2388
rect 14171 2350 14175 2382
rect 14175 2350 14207 2382
rect 14207 2350 14211 2382
rect 14171 2314 14211 2350
rect 14171 2282 14175 2314
rect 14175 2282 14207 2314
rect 14207 2282 14211 2314
rect 14171 2246 14211 2282
rect 14171 2214 14175 2246
rect 14175 2214 14207 2246
rect 14207 2214 14211 2246
rect 14171 2178 14211 2214
rect 14171 2146 14175 2178
rect 14175 2146 14207 2178
rect 14207 2146 14211 2178
rect 14171 2110 14211 2146
rect 14171 2078 14175 2110
rect 14175 2078 14207 2110
rect 14207 2078 14211 2110
rect 14171 2042 14211 2078
rect 14171 2010 14175 2042
rect 14175 2010 14207 2042
rect 14207 2010 14211 2042
rect 14171 1974 14211 2010
rect 14171 1942 14175 1974
rect 14175 1942 14207 1974
rect 14207 1942 14211 1974
rect 14171 1906 14211 1942
rect 14171 1874 14175 1906
rect 14175 1874 14207 1906
rect 14207 1874 14211 1906
rect 14171 1838 14211 1874
rect 14171 1806 14175 1838
rect 14175 1806 14207 1838
rect 14207 1806 14211 1838
rect 14171 1770 14211 1806
rect 14171 1738 14175 1770
rect 14175 1738 14207 1770
rect 14207 1738 14211 1770
rect 14171 1702 14211 1738
rect 14171 1670 14175 1702
rect 14175 1670 14207 1702
rect 14207 1670 14211 1702
rect 14171 1634 14211 1670
rect 14171 1602 14175 1634
rect 14175 1602 14207 1634
rect 14207 1602 14211 1634
rect 14171 1566 14211 1602
rect 14171 1534 14175 1566
rect 14175 1534 14207 1566
rect 14207 1534 14211 1566
rect 14171 1528 14211 1534
rect 13828 1414 13950 1420
rect 13828 1382 13873 1414
rect 13873 1382 13905 1414
rect 13905 1382 13950 1414
rect 13828 1346 13950 1382
rect 13828 1314 13873 1346
rect 13873 1314 13905 1346
rect 13905 1314 13950 1346
rect 13828 1278 13950 1314
rect 13828 1246 13873 1278
rect 13873 1246 13905 1278
rect 13905 1246 13950 1278
rect 13828 1210 13950 1246
rect 13828 1178 13873 1210
rect 13873 1178 13905 1210
rect 13905 1178 13950 1210
rect 13828 1142 13950 1178
rect 13828 1110 13873 1142
rect 13873 1110 13905 1142
rect 13905 1110 13950 1142
rect 13828 1074 13950 1110
rect 13828 1042 13873 1074
rect 13873 1042 13905 1074
rect 13905 1042 13950 1074
rect 13828 1006 13950 1042
rect 13828 974 13873 1006
rect 13873 974 13905 1006
rect 13905 974 13950 1006
rect 13828 938 13950 974
rect 13828 906 13873 938
rect 13873 906 13905 938
rect 13905 906 13950 938
rect 13828 870 13950 906
rect 13828 838 13873 870
rect 13873 838 13905 870
rect 13905 838 13950 870
rect 13828 802 13950 838
rect 13828 770 13873 802
rect 13873 770 13905 802
rect 13905 770 13950 802
rect 13828 734 13950 770
rect 13828 702 13873 734
rect 13873 702 13905 734
rect 13905 702 13950 734
rect 13828 666 13950 702
rect 13828 634 13873 666
rect 13873 634 13905 666
rect 13905 634 13950 666
rect 13828 598 13950 634
rect 13828 566 13873 598
rect 13873 566 13905 598
rect 13905 566 13950 598
rect 13828 560 13950 566
rect 14432 2382 14554 2388
rect 14432 2350 14477 2382
rect 14477 2350 14509 2382
rect 14509 2350 14554 2382
rect 14432 2314 14554 2350
rect 14432 2282 14477 2314
rect 14477 2282 14509 2314
rect 14509 2282 14554 2314
rect 14432 2246 14554 2282
rect 14432 2214 14477 2246
rect 14477 2214 14509 2246
rect 14509 2214 14554 2246
rect 14432 2178 14554 2214
rect 14432 2146 14477 2178
rect 14477 2146 14509 2178
rect 14509 2146 14554 2178
rect 14432 2110 14554 2146
rect 14432 2078 14477 2110
rect 14477 2078 14509 2110
rect 14509 2078 14554 2110
rect 14432 2042 14554 2078
rect 14432 2010 14477 2042
rect 14477 2010 14509 2042
rect 14509 2010 14554 2042
rect 14432 1974 14554 2010
rect 14432 1942 14477 1974
rect 14477 1942 14509 1974
rect 14509 1942 14554 1974
rect 14432 1906 14554 1942
rect 14432 1874 14477 1906
rect 14477 1874 14509 1906
rect 14509 1874 14554 1906
rect 14432 1838 14554 1874
rect 14432 1806 14477 1838
rect 14477 1806 14509 1838
rect 14509 1806 14554 1838
rect 14432 1770 14554 1806
rect 14432 1738 14477 1770
rect 14477 1738 14509 1770
rect 14509 1738 14554 1770
rect 14432 1702 14554 1738
rect 14432 1670 14477 1702
rect 14477 1670 14509 1702
rect 14509 1670 14554 1702
rect 14432 1634 14554 1670
rect 14432 1602 14477 1634
rect 14477 1602 14509 1634
rect 14509 1602 14554 1634
rect 14432 1566 14554 1602
rect 14432 1534 14477 1566
rect 14477 1534 14509 1566
rect 14509 1534 14554 1566
rect 14432 1528 14554 1534
rect 14171 1414 14211 1420
rect 14171 1382 14175 1414
rect 14175 1382 14207 1414
rect 14207 1382 14211 1414
rect 14171 1346 14211 1382
rect 14171 1314 14175 1346
rect 14175 1314 14207 1346
rect 14207 1314 14211 1346
rect 14171 1278 14211 1314
rect 14171 1246 14175 1278
rect 14175 1246 14207 1278
rect 14207 1246 14211 1278
rect 14171 1210 14211 1246
rect 14171 1178 14175 1210
rect 14175 1178 14207 1210
rect 14207 1178 14211 1210
rect 14171 1142 14211 1178
rect 14171 1110 14175 1142
rect 14175 1110 14207 1142
rect 14207 1110 14211 1142
rect 14171 1074 14211 1110
rect 14171 1042 14175 1074
rect 14175 1042 14207 1074
rect 14207 1042 14211 1074
rect 14171 1006 14211 1042
rect 14171 974 14175 1006
rect 14175 974 14207 1006
rect 14207 974 14211 1006
rect 14171 938 14211 974
rect 14171 906 14175 938
rect 14175 906 14207 938
rect 14207 906 14211 938
rect 14171 870 14211 906
rect 14171 838 14175 870
rect 14175 838 14207 870
rect 14207 838 14211 870
rect 14171 802 14211 838
rect 14171 770 14175 802
rect 14175 770 14207 802
rect 14207 770 14211 802
rect 14171 734 14211 770
rect 14171 702 14175 734
rect 14175 702 14207 734
rect 14207 702 14211 734
rect 14171 666 14211 702
rect 14171 634 14175 666
rect 14175 634 14207 666
rect 14207 634 14211 666
rect 14171 598 14211 634
rect 14171 566 14175 598
rect 14175 566 14207 598
rect 14207 566 14211 598
rect 14171 560 14211 566
rect 14432 1414 14554 1420
rect 14432 1382 14477 1414
rect 14477 1382 14509 1414
rect 14509 1382 14554 1414
rect 14432 1346 14554 1382
rect 14432 1314 14477 1346
rect 14477 1314 14509 1346
rect 14509 1314 14554 1346
rect 14432 1278 14554 1314
rect 14432 1246 14477 1278
rect 14477 1246 14509 1278
rect 14509 1246 14554 1278
rect 14432 1210 14554 1246
rect 14432 1178 14477 1210
rect 14477 1178 14509 1210
rect 14509 1178 14554 1210
rect 14432 1142 14554 1178
rect 14432 1110 14477 1142
rect 14477 1110 14509 1142
rect 14509 1110 14554 1142
rect 14432 1074 14554 1110
rect 14432 1042 14477 1074
rect 14477 1042 14509 1074
rect 14509 1042 14554 1074
rect 14432 1006 14554 1042
rect 14432 974 14477 1006
rect 14477 974 14509 1006
rect 14509 974 14554 1006
rect 14432 938 14554 974
rect 14432 906 14477 938
rect 14477 906 14509 938
rect 14509 906 14554 938
rect 14432 870 14554 906
rect 14432 838 14477 870
rect 14477 838 14509 870
rect 14509 838 14554 870
rect 14432 802 14554 838
rect 14432 770 14477 802
rect 14477 770 14509 802
rect 14509 770 14554 802
rect 14432 734 14554 770
rect 14432 702 14477 734
rect 14477 702 14509 734
rect 14509 702 14554 734
rect 14432 666 14554 702
rect 14432 634 14477 666
rect 14477 634 14509 666
rect 14509 634 14554 666
rect 14432 598 14554 634
rect 14432 566 14477 598
rect 14477 566 14509 598
rect 14509 566 14554 598
rect 14432 560 14554 566
rect 1487 410 1527 414
rect 2091 410 2131 414
rect 2695 410 2735 414
rect 3299 410 3339 414
rect 3903 410 3943 414
rect 4507 410 4547 414
rect 5111 410 5151 414
rect 5715 410 5755 414
rect 6319 410 6359 414
rect 6923 410 6963 414
rect 7527 410 7567 414
rect 8131 410 8171 414
rect 8735 410 8775 414
rect 9339 410 9379 414
rect 9943 410 9983 414
rect 10547 410 10587 414
rect 11151 410 11191 414
rect 11755 410 11795 414
rect 12359 410 12399 414
rect 12963 410 13003 414
rect 13567 410 13607 414
rect 14171 410 14211 414
rect 1487 378 1490 410
rect 1490 378 1522 410
rect 1522 378 1527 410
rect 2091 378 2102 410
rect 2102 378 2131 410
rect 2695 378 2714 410
rect 2714 378 2735 410
rect 3299 378 3326 410
rect 3326 378 3339 410
rect 3903 378 3938 410
rect 3938 378 3943 410
rect 4507 378 4514 410
rect 4514 378 4547 410
rect 5111 378 5126 410
rect 5126 378 5151 410
rect 5715 378 5738 410
rect 5738 378 5755 410
rect 6319 378 6350 410
rect 6350 378 6359 410
rect 6923 378 6930 410
rect 6930 378 6962 410
rect 6962 378 6963 410
rect 7527 378 7542 410
rect 7542 378 7567 410
rect 8131 378 8154 410
rect 8154 378 8171 410
rect 8735 378 8766 410
rect 8766 378 8775 410
rect 9339 378 9342 410
rect 9342 378 9378 410
rect 9378 378 9379 410
rect 9943 378 9954 410
rect 9954 378 9983 410
rect 10547 378 10566 410
rect 10566 378 10587 410
rect 11151 378 11178 410
rect 11178 378 11191 410
rect 11755 378 11758 410
rect 11758 378 11790 410
rect 11790 378 11795 410
rect 12359 378 12370 410
rect 12370 378 12399 410
rect 12963 378 12982 410
rect 12982 378 13003 410
rect 13567 378 13594 410
rect 13594 378 13607 410
rect 14171 378 14206 410
rect 14206 378 14211 410
rect 1487 374 1527 378
rect 2091 374 2131 378
rect 2695 374 2735 378
rect 3299 374 3339 378
rect 3903 374 3943 378
rect 4507 374 4547 378
rect 5111 374 5151 378
rect 5715 374 5755 378
rect 6319 374 6359 378
rect 6923 374 6963 378
rect 7527 374 7567 378
rect 8131 374 8171 378
rect 8735 374 8775 378
rect 9339 374 9379 378
rect 9943 374 9983 378
rect 10547 374 10587 378
rect 11151 374 11191 378
rect 11755 374 11795 378
rect 12359 374 12399 378
rect 12963 374 13003 378
rect 13567 374 13607 378
rect 14171 374 14211 378
<< metal2 >>
rect 933 4368 973 4884
rect 933 4237 973 4246
rect 1487 4840 1527 4884
rect 1748 4324 1870 4884
rect 1748 3356 1870 3464
rect 1748 2388 1870 2496
rect 1748 1420 1870 1528
rect 1748 551 1870 560
rect 2091 4840 2131 4884
rect 1487 0 1527 44
rect 2352 4324 2474 4884
rect 2352 3356 2474 3464
rect 2352 2388 2474 2496
rect 2352 1420 2474 1528
rect 2352 551 2474 560
rect 2695 4840 2735 4884
rect 2091 0 2131 44
rect 2956 4324 3078 4884
rect 2956 3356 3078 3464
rect 2956 2388 3078 2496
rect 2956 1420 3078 1528
rect 2956 551 3078 560
rect 3299 4840 3339 4884
rect 2695 0 2735 44
rect 3560 4324 3682 4884
rect 3560 3356 3682 3464
rect 3560 2388 3682 2496
rect 3560 1420 3682 1528
rect 3560 551 3682 560
rect 3903 4840 3943 4884
rect 3299 0 3339 44
rect 4164 4324 4286 4884
rect 4164 3356 4286 3464
rect 4164 2388 4286 2496
rect 4164 1420 4286 1528
rect 4164 551 4286 560
rect 4507 4840 4547 4884
rect 3903 0 3943 44
rect 4768 4324 4890 4884
rect 4768 3356 4890 3464
rect 4768 2388 4890 2496
rect 4768 1420 4890 1528
rect 4768 551 4890 560
rect 5111 4840 5151 4884
rect 4507 0 4547 44
rect 5372 4324 5494 4884
rect 5372 3356 5494 3464
rect 5372 2388 5494 2496
rect 5372 1420 5494 1528
rect 5372 551 5494 560
rect 5715 4840 5755 4884
rect 5111 0 5151 44
rect 5976 4324 6098 4884
rect 5976 3356 6098 3464
rect 5976 2388 6098 2496
rect 5976 1420 6098 1528
rect 5976 551 6098 560
rect 6319 4840 6359 4884
rect 5715 0 5755 44
rect 6580 4324 6702 4884
rect 6580 3356 6702 3464
rect 6580 2388 6702 2496
rect 6580 1420 6702 1528
rect 6580 551 6702 560
rect 6923 4840 6963 4884
rect 6319 0 6359 44
rect 7184 4324 7306 4884
rect 7184 3356 7306 3464
rect 7184 2388 7306 2496
rect 7184 1420 7306 1528
rect 7184 551 7306 560
rect 7527 4840 7567 4884
rect 6923 0 6963 44
rect 7788 4324 7910 4884
rect 7788 3356 7910 3464
rect 7788 2388 7910 2496
rect 7788 1420 7910 1528
rect 7788 551 7910 560
rect 8131 4840 8171 4884
rect 7527 0 7567 44
rect 8392 4324 8514 4884
rect 8392 3356 8514 3464
rect 8392 2388 8514 2496
rect 8392 1420 8514 1528
rect 8392 551 8514 560
rect 8735 4840 8775 4884
rect 8131 0 8171 44
rect 8996 4324 9118 4884
rect 8996 3356 9118 3464
rect 8996 2388 9118 2496
rect 8996 1420 9118 1528
rect 8996 551 9118 560
rect 9339 4840 9379 4884
rect 8735 0 8775 44
rect 9600 4324 9722 4884
rect 9600 3356 9722 3464
rect 9600 2388 9722 2496
rect 9600 1420 9722 1528
rect 9600 551 9722 560
rect 9943 4840 9983 4884
rect 9339 0 9379 44
rect 10204 4324 10326 4884
rect 10204 3356 10326 3464
rect 10204 2388 10326 2496
rect 10204 1420 10326 1528
rect 10204 551 10326 560
rect 10547 4840 10587 4884
rect 9943 0 9983 44
rect 10808 4324 10930 4884
rect 10808 3356 10930 3464
rect 10808 2388 10930 2496
rect 10808 1420 10930 1528
rect 10808 551 10930 560
rect 11151 4840 11191 4884
rect 10547 0 10587 44
rect 11412 4324 11534 4884
rect 11412 3356 11534 3464
rect 11412 2388 11534 2496
rect 11412 1420 11534 1528
rect 11412 551 11534 560
rect 11755 4840 11795 4884
rect 11151 0 11191 44
rect 12016 4324 12138 4884
rect 12016 3356 12138 3464
rect 12016 2388 12138 2496
rect 12016 1420 12138 1528
rect 12016 551 12138 560
rect 12359 4840 12399 4884
rect 11755 0 11795 44
rect 12620 4324 12742 4884
rect 12620 3356 12742 3464
rect 12620 2388 12742 2496
rect 12620 1420 12742 1528
rect 12620 551 12742 560
rect 12963 4840 13003 4884
rect 12359 0 12399 44
rect 13224 4324 13346 4884
rect 13224 3356 13346 3464
rect 13224 2388 13346 2496
rect 13224 1420 13346 1528
rect 13224 551 13346 560
rect 13567 4840 13607 4884
rect 12963 0 13003 44
rect 13828 4324 13950 4884
rect 13828 3356 13950 3464
rect 13828 2388 13950 2496
rect 13828 1420 13950 1528
rect 13828 551 13950 560
rect 14171 4840 14211 4884
rect 13567 0 13607 44
rect 14432 4324 14554 4884
rect 14432 3356 14554 3464
rect 14432 2388 14554 2496
rect 14432 1420 14554 1528
rect 14432 551 14554 560
rect 14171 0 14211 44
<< via2 >>
rect 1487 4510 1527 4840
rect 1487 4470 1527 4510
rect 1487 4324 1527 4470
rect 1487 3464 1527 4324
rect 1487 3356 1527 3464
rect 1487 2496 1527 3356
rect 1487 2388 1527 2496
rect 1487 1528 1527 2388
rect 1487 1420 1527 1528
rect 1487 560 1527 1420
rect 1487 414 1527 560
rect 2091 4510 2131 4840
rect 2091 4470 2131 4510
rect 2091 4324 2131 4470
rect 2091 3464 2131 4324
rect 2091 3356 2131 3464
rect 2091 2496 2131 3356
rect 2091 2388 2131 2496
rect 2091 1528 2131 2388
rect 2091 1420 2131 1528
rect 2091 560 2131 1420
rect 1487 374 1527 414
rect 1487 44 1527 374
rect 2091 414 2131 560
rect 2695 4510 2735 4840
rect 2695 4470 2735 4510
rect 2695 4324 2735 4470
rect 2695 3464 2735 4324
rect 2695 3356 2735 3464
rect 2695 2496 2735 3356
rect 2695 2388 2735 2496
rect 2695 1528 2735 2388
rect 2695 1420 2735 1528
rect 2695 560 2735 1420
rect 2091 374 2131 414
rect 2091 44 2131 374
rect 2695 414 2735 560
rect 3299 4510 3339 4840
rect 3299 4470 3339 4510
rect 3299 4324 3339 4470
rect 3299 3464 3339 4324
rect 3299 3356 3339 3464
rect 3299 2496 3339 3356
rect 3299 2388 3339 2496
rect 3299 1528 3339 2388
rect 3299 1420 3339 1528
rect 3299 560 3339 1420
rect 2695 374 2735 414
rect 2695 44 2735 374
rect 3299 414 3339 560
rect 3903 4510 3943 4840
rect 3903 4470 3943 4510
rect 3903 4324 3943 4470
rect 3903 3464 3943 4324
rect 3903 3356 3943 3464
rect 3903 2496 3943 3356
rect 3903 2388 3943 2496
rect 3903 1528 3943 2388
rect 3903 1420 3943 1528
rect 3903 560 3943 1420
rect 3299 374 3339 414
rect 3299 44 3339 374
rect 3903 414 3943 560
rect 4507 4510 4547 4840
rect 4507 4470 4547 4510
rect 4507 4324 4547 4470
rect 4507 3464 4547 4324
rect 4507 3356 4547 3464
rect 4507 2496 4547 3356
rect 4507 2388 4547 2496
rect 4507 1528 4547 2388
rect 4507 1420 4547 1528
rect 4507 560 4547 1420
rect 3903 374 3943 414
rect 3903 44 3943 374
rect 4507 414 4547 560
rect 5111 4510 5151 4840
rect 5111 4470 5151 4510
rect 5111 4324 5151 4470
rect 5111 3464 5151 4324
rect 5111 3356 5151 3464
rect 5111 2496 5151 3356
rect 5111 2388 5151 2496
rect 5111 1528 5151 2388
rect 5111 1420 5151 1528
rect 5111 560 5151 1420
rect 4507 374 4547 414
rect 4507 44 4547 374
rect 5111 414 5151 560
rect 5715 4510 5755 4840
rect 5715 4470 5755 4510
rect 5715 4324 5755 4470
rect 5715 3464 5755 4324
rect 5715 3356 5755 3464
rect 5715 2496 5755 3356
rect 5715 2388 5755 2496
rect 5715 1528 5755 2388
rect 5715 1420 5755 1528
rect 5715 560 5755 1420
rect 5111 374 5151 414
rect 5111 44 5151 374
rect 5715 414 5755 560
rect 6319 4510 6359 4840
rect 6319 4470 6359 4510
rect 6319 4324 6359 4470
rect 6319 3464 6359 4324
rect 6319 3356 6359 3464
rect 6319 2496 6359 3356
rect 6319 2388 6359 2496
rect 6319 1528 6359 2388
rect 6319 1420 6359 1528
rect 6319 560 6359 1420
rect 5715 374 5755 414
rect 5715 44 5755 374
rect 6319 414 6359 560
rect 6923 4510 6963 4840
rect 6923 4470 6963 4510
rect 6923 4324 6963 4470
rect 6923 3464 6963 4324
rect 6923 3356 6963 3464
rect 6923 2496 6963 3356
rect 6923 2388 6963 2496
rect 6923 1528 6963 2388
rect 6923 1420 6963 1528
rect 6923 560 6963 1420
rect 6319 374 6359 414
rect 6319 44 6359 374
rect 6923 414 6963 560
rect 7527 4510 7567 4840
rect 7527 4470 7567 4510
rect 7527 4324 7567 4470
rect 7527 3464 7567 4324
rect 7527 3356 7567 3464
rect 7527 2496 7567 3356
rect 7527 2388 7567 2496
rect 7527 1528 7567 2388
rect 7527 1420 7567 1528
rect 7527 560 7567 1420
rect 6923 374 6963 414
rect 6923 44 6963 374
rect 7527 414 7567 560
rect 8131 4510 8171 4840
rect 8131 4470 8171 4510
rect 8131 4324 8171 4470
rect 8131 3464 8171 4324
rect 8131 3356 8171 3464
rect 8131 2496 8171 3356
rect 8131 2388 8171 2496
rect 8131 1528 8171 2388
rect 8131 1420 8171 1528
rect 8131 560 8171 1420
rect 7527 374 7567 414
rect 7527 44 7567 374
rect 8131 414 8171 560
rect 8735 4510 8775 4840
rect 8735 4470 8775 4510
rect 8735 4324 8775 4470
rect 8735 3464 8775 4324
rect 8735 3356 8775 3464
rect 8735 2496 8775 3356
rect 8735 2388 8775 2496
rect 8735 1528 8775 2388
rect 8735 1420 8775 1528
rect 8735 560 8775 1420
rect 8131 374 8171 414
rect 8131 44 8171 374
rect 8735 414 8775 560
rect 9339 4510 9379 4840
rect 9339 4470 9379 4510
rect 9339 4324 9379 4470
rect 9339 3464 9379 4324
rect 9339 3356 9379 3464
rect 9339 2496 9379 3356
rect 9339 2388 9379 2496
rect 9339 1528 9379 2388
rect 9339 1420 9379 1528
rect 9339 560 9379 1420
rect 8735 374 8775 414
rect 8735 44 8775 374
rect 9339 414 9379 560
rect 9943 4510 9983 4840
rect 9943 4470 9983 4510
rect 9943 4324 9983 4470
rect 9943 3464 9983 4324
rect 9943 3356 9983 3464
rect 9943 2496 9983 3356
rect 9943 2388 9983 2496
rect 9943 1528 9983 2388
rect 9943 1420 9983 1528
rect 9943 560 9983 1420
rect 9339 374 9379 414
rect 9339 44 9379 374
rect 9943 414 9983 560
rect 10547 4510 10587 4840
rect 10547 4470 10587 4510
rect 10547 4324 10587 4470
rect 10547 3464 10587 4324
rect 10547 3356 10587 3464
rect 10547 2496 10587 3356
rect 10547 2388 10587 2496
rect 10547 1528 10587 2388
rect 10547 1420 10587 1528
rect 10547 560 10587 1420
rect 9943 374 9983 414
rect 9943 44 9983 374
rect 10547 414 10587 560
rect 11151 4510 11191 4840
rect 11151 4470 11191 4510
rect 11151 4324 11191 4470
rect 11151 3464 11191 4324
rect 11151 3356 11191 3464
rect 11151 2496 11191 3356
rect 11151 2388 11191 2496
rect 11151 1528 11191 2388
rect 11151 1420 11191 1528
rect 11151 560 11191 1420
rect 10547 374 10587 414
rect 10547 44 10587 374
rect 11151 414 11191 560
rect 11755 4510 11795 4840
rect 11755 4470 11795 4510
rect 11755 4324 11795 4470
rect 11755 3464 11795 4324
rect 11755 3356 11795 3464
rect 11755 2496 11795 3356
rect 11755 2388 11795 2496
rect 11755 1528 11795 2388
rect 11755 1420 11795 1528
rect 11755 560 11795 1420
rect 11151 374 11191 414
rect 11151 44 11191 374
rect 11755 414 11795 560
rect 12359 4510 12399 4840
rect 12359 4470 12399 4510
rect 12359 4324 12399 4470
rect 12359 3464 12399 4324
rect 12359 3356 12399 3464
rect 12359 2496 12399 3356
rect 12359 2388 12399 2496
rect 12359 1528 12399 2388
rect 12359 1420 12399 1528
rect 12359 560 12399 1420
rect 11755 374 11795 414
rect 11755 44 11795 374
rect 12359 414 12399 560
rect 12963 4510 13003 4840
rect 12963 4470 13003 4510
rect 12963 4324 13003 4470
rect 12963 3464 13003 4324
rect 12963 3356 13003 3464
rect 12963 2496 13003 3356
rect 12963 2388 13003 2496
rect 12963 1528 13003 2388
rect 12963 1420 13003 1528
rect 12963 560 13003 1420
rect 12359 374 12399 414
rect 12359 44 12399 374
rect 12963 414 13003 560
rect 13567 4510 13607 4840
rect 13567 4470 13607 4510
rect 13567 4324 13607 4470
rect 13567 3464 13607 4324
rect 13567 3356 13607 3464
rect 13567 2496 13607 3356
rect 13567 2388 13607 2496
rect 13567 1528 13607 2388
rect 13567 1420 13607 1528
rect 13567 560 13607 1420
rect 12963 374 13003 414
rect 12963 44 13003 374
rect 13567 414 13607 560
rect 14171 4510 14211 4840
rect 14171 4470 14211 4510
rect 14171 4324 14211 4470
rect 14171 3464 14211 4324
rect 14171 3356 14211 3464
rect 14171 2496 14211 3356
rect 14171 2388 14211 2496
rect 14171 1528 14211 2388
rect 14171 1420 14211 1528
rect 14171 560 14211 1420
rect 13567 374 13607 414
rect 13567 44 13607 374
rect 14171 414 14211 560
rect 14171 374 14211 414
rect 14171 44 14211 374
<< metal3 >>
rect 1487 4840 1527 4849
rect 1487 35 1527 44
rect 2091 4840 2131 4849
rect 2091 35 2131 44
rect 2695 4840 2735 4849
rect 2695 35 2735 44
rect 3299 4840 3339 4849
rect 3299 35 3339 44
rect 3903 4840 3943 4849
rect 3903 35 3943 44
rect 4507 4840 4547 4849
rect 4507 35 4547 44
rect 5111 4840 5151 4849
rect 5111 35 5151 44
rect 5715 4840 5755 4849
rect 5715 35 5755 44
rect 6319 4840 6359 4849
rect 6319 35 6359 44
rect 6923 4840 6963 4849
rect 6923 35 6963 44
rect 7527 4840 7567 4849
rect 7527 35 7567 44
rect 8131 4840 8171 4849
rect 8131 35 8171 44
rect 8735 4840 8775 4849
rect 8735 35 8775 44
rect 9339 4840 9379 4849
rect 9339 35 9379 44
rect 9943 4840 9983 4849
rect 9943 35 9983 44
rect 10547 4840 10587 4849
rect 10547 35 10587 44
rect 11151 4840 11191 4849
rect 11151 35 11191 44
rect 11755 4840 11795 4849
rect 11755 35 11795 44
rect 12359 4840 12399 4849
rect 12359 35 12399 44
rect 12963 4840 13003 4849
rect 12963 35 13003 44
rect 13567 4840 13607 4849
rect 13567 35 13607 44
rect 14171 4840 14211 4849
rect 14171 35 14211 44
<< labels >>
rlabel metal2 s 933 4237 973 4884 4 gate
port 3 nsew
rlabel metal2 s 2956 551 3078 4884 4 pad
port 2 nsew
rlabel metal2 s 3560 551 3682 4884 4 pad
port 2 nsew
rlabel metal2 s 11412 551 11534 4884 4 pad
port 2 nsew
rlabel metal2 s 12016 551 12138 4884 4 pad
port 2 nsew
rlabel metal2 s 8392 551 8514 4884 4 pad
port 2 nsew
rlabel metal2 s 8996 551 9118 4884 4 pad
port 2 nsew
rlabel metal2 s 12620 551 12742 4884 4 pad
port 2 nsew
rlabel metal2 s 9600 551 9722 4884 4 pad
port 2 nsew
rlabel metal2 s 10808 551 10930 4884 4 pad
port 2 nsew
rlabel metal2 s 4164 551 4286 4884 4 pad
port 2 nsew
rlabel metal2 s 14432 551 14554 4884 4 pad
port 2 nsew
rlabel metal2 s 7184 551 7306 4884 4 pad
port 2 nsew
rlabel metal2 s 5976 551 6098 4884 4 pad
port 2 nsew
rlabel metal2 s 13224 551 13346 4884 4 pad
port 2 nsew
rlabel metal2 s 7788 551 7910 4884 4 pad
port 2 nsew
rlabel metal2 s 4768 551 4890 4884 4 pad
port 2 nsew
rlabel metal2 s 10204 551 10326 4884 4 pad
port 2 nsew
rlabel metal2 s 5372 551 5494 4884 4 pad
port 2 nsew
rlabel metal2 s 2352 551 2474 4884 4 pad
port 2 nsew
rlabel metal2 s 1748 551 1870 4884 4 pad
port 2 nsew
rlabel metal2 s 13828 551 13950 4884 4 pad
port 2 nsew
rlabel metal2 s 6580 551 6702 4884 4 pad
port 2 nsew
rlabel comment s 394 394 394 394 4 sub!
flabel comment s 954 4196 954 4196 0 FreeSans 400 0 0 0 dant
flabel metal1 s 448 366 938 424 0 FreeSans 51 0 0 0 iovss
port 1 nsew
<< properties >>
string device primitive
string GDS_END 533726
string GDS_FILE sg13g2_io.gds
string GDS_START 122
<< end >>
