magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2026 -2026 18026 5878
<< nwell >>
rect 236 236 15764 3616
<< pwell >>
rect -26 3758 16026 3878
rect -26 94 94 3758
rect 15906 94 16026 3758
rect -26 -26 16026 94
<< hvpmos >>
rect 5799 1970 5919 3302
rect 6155 1970 6275 3302
rect 6403 1970 6523 3302
rect 6759 1970 6879 3302
rect 7007 1970 7127 3302
rect 7363 1970 7483 3302
rect 7611 1970 7731 3302
rect 7967 1970 8087 3302
rect 8215 1970 8335 3302
rect 8571 1970 8691 3302
rect 8819 1970 8939 3302
rect 9175 1970 9295 3302
rect 9423 1970 9543 3302
rect 9779 1970 9899 3302
rect 10027 1970 10147 3302
rect 5799 550 5919 1882
rect 6155 550 6275 1882
rect 6403 550 6523 1882
rect 6759 550 6879 1882
rect 7007 550 7127 1882
rect 7363 550 7483 1882
rect 7611 550 7731 1882
rect 7967 550 8087 1882
rect 8215 550 8335 1882
rect 8571 550 8691 1882
rect 8819 550 8939 1882
rect 9175 550 9295 1882
rect 9423 550 9543 1882
rect 9779 550 9899 1882
rect 10027 550 10147 1882
<< hvpdiff >>
rect 5705 3264 5799 3302
rect 5705 3232 5719 3264
rect 5751 3232 5799 3264
rect 5705 3196 5799 3232
rect 5705 3164 5719 3196
rect 5751 3164 5799 3196
rect 5705 3128 5799 3164
rect 5705 3096 5719 3128
rect 5751 3096 5799 3128
rect 5705 3060 5799 3096
rect 5705 3028 5719 3060
rect 5751 3028 5799 3060
rect 5705 2992 5799 3028
rect 5705 2960 5719 2992
rect 5751 2960 5799 2992
rect 5705 2924 5799 2960
rect 5705 2892 5719 2924
rect 5751 2892 5799 2924
rect 5705 2856 5799 2892
rect 5705 2824 5719 2856
rect 5751 2824 5799 2856
rect 5705 2788 5799 2824
rect 5705 2756 5719 2788
rect 5751 2756 5799 2788
rect 5705 2720 5799 2756
rect 5705 2688 5719 2720
rect 5751 2688 5799 2720
rect 5705 2652 5799 2688
rect 5705 2620 5719 2652
rect 5751 2620 5799 2652
rect 5705 2584 5799 2620
rect 5705 2552 5719 2584
rect 5751 2552 5799 2584
rect 5705 2516 5799 2552
rect 5705 2484 5719 2516
rect 5751 2484 5799 2516
rect 5705 2448 5799 2484
rect 5705 2416 5719 2448
rect 5751 2416 5799 2448
rect 5705 2380 5799 2416
rect 5705 2348 5719 2380
rect 5751 2348 5799 2380
rect 5705 2312 5799 2348
rect 5705 2280 5719 2312
rect 5751 2280 5799 2312
rect 5705 2244 5799 2280
rect 5705 2212 5719 2244
rect 5751 2212 5799 2244
rect 5705 2176 5799 2212
rect 5705 2144 5719 2176
rect 5751 2144 5799 2176
rect 5705 2108 5799 2144
rect 5705 2076 5719 2108
rect 5751 2076 5799 2108
rect 5705 2040 5799 2076
rect 5705 2008 5719 2040
rect 5751 2008 5799 2040
rect 5705 1970 5799 2008
rect 5919 3264 6155 3302
rect 5919 3232 6021 3264
rect 6053 3232 6155 3264
rect 5919 3196 6155 3232
rect 5919 3164 6021 3196
rect 6053 3164 6155 3196
rect 5919 3128 6155 3164
rect 5919 3096 6021 3128
rect 6053 3096 6155 3128
rect 5919 3060 6155 3096
rect 5919 3028 6021 3060
rect 6053 3028 6155 3060
rect 5919 2992 6155 3028
rect 5919 2960 6021 2992
rect 6053 2960 6155 2992
rect 5919 2924 6155 2960
rect 5919 2892 6021 2924
rect 6053 2892 6155 2924
rect 5919 2856 6155 2892
rect 5919 2824 6021 2856
rect 6053 2824 6155 2856
rect 5919 2788 6155 2824
rect 5919 2756 6021 2788
rect 6053 2756 6155 2788
rect 5919 2720 6155 2756
rect 5919 2688 6021 2720
rect 6053 2688 6155 2720
rect 5919 2652 6155 2688
rect 5919 2620 6021 2652
rect 6053 2620 6155 2652
rect 5919 2584 6155 2620
rect 5919 2552 6021 2584
rect 6053 2552 6155 2584
rect 5919 2516 6155 2552
rect 5919 2484 6021 2516
rect 6053 2484 6155 2516
rect 5919 2448 6155 2484
rect 5919 2416 6021 2448
rect 6053 2416 6155 2448
rect 5919 2380 6155 2416
rect 5919 2348 6021 2380
rect 6053 2348 6155 2380
rect 5919 2312 6155 2348
rect 5919 2280 6021 2312
rect 6053 2280 6155 2312
rect 5919 2244 6155 2280
rect 5919 2212 6021 2244
rect 6053 2212 6155 2244
rect 5919 2176 6155 2212
rect 5919 2144 6021 2176
rect 6053 2144 6155 2176
rect 5919 2108 6155 2144
rect 5919 2076 6021 2108
rect 6053 2076 6155 2108
rect 5919 2040 6155 2076
rect 5919 2008 6021 2040
rect 6053 2008 6155 2040
rect 5919 1970 6155 2008
rect 6275 3264 6403 3302
rect 6275 3232 6323 3264
rect 6355 3232 6403 3264
rect 6275 3196 6403 3232
rect 6275 3164 6323 3196
rect 6355 3164 6403 3196
rect 6275 3128 6403 3164
rect 6275 3096 6323 3128
rect 6355 3096 6403 3128
rect 6275 3060 6403 3096
rect 6275 3028 6323 3060
rect 6355 3028 6403 3060
rect 6275 2992 6403 3028
rect 6275 2960 6323 2992
rect 6355 2960 6403 2992
rect 6275 2924 6403 2960
rect 6275 2892 6323 2924
rect 6355 2892 6403 2924
rect 6275 2856 6403 2892
rect 6275 2824 6323 2856
rect 6355 2824 6403 2856
rect 6275 2788 6403 2824
rect 6275 2756 6323 2788
rect 6355 2756 6403 2788
rect 6275 2720 6403 2756
rect 6275 2688 6323 2720
rect 6355 2688 6403 2720
rect 6275 2652 6403 2688
rect 6275 2620 6323 2652
rect 6355 2620 6403 2652
rect 6275 2584 6403 2620
rect 6275 2552 6323 2584
rect 6355 2552 6403 2584
rect 6275 2516 6403 2552
rect 6275 2484 6323 2516
rect 6355 2484 6403 2516
rect 6275 2448 6403 2484
rect 6275 2416 6323 2448
rect 6355 2416 6403 2448
rect 6275 2380 6403 2416
rect 6275 2348 6323 2380
rect 6355 2348 6403 2380
rect 6275 2312 6403 2348
rect 6275 2280 6323 2312
rect 6355 2280 6403 2312
rect 6275 2244 6403 2280
rect 6275 2212 6323 2244
rect 6355 2212 6403 2244
rect 6275 2176 6403 2212
rect 6275 2144 6323 2176
rect 6355 2144 6403 2176
rect 6275 2108 6403 2144
rect 6275 2076 6323 2108
rect 6355 2076 6403 2108
rect 6275 2040 6403 2076
rect 6275 2008 6323 2040
rect 6355 2008 6403 2040
rect 6275 1970 6403 2008
rect 6523 3264 6759 3302
rect 6523 3232 6625 3264
rect 6657 3232 6759 3264
rect 6523 3196 6759 3232
rect 6523 3164 6625 3196
rect 6657 3164 6759 3196
rect 6523 3128 6759 3164
rect 6523 3096 6625 3128
rect 6657 3096 6759 3128
rect 6523 3060 6759 3096
rect 6523 3028 6625 3060
rect 6657 3028 6759 3060
rect 6523 2992 6759 3028
rect 6523 2960 6625 2992
rect 6657 2960 6759 2992
rect 6523 2924 6759 2960
rect 6523 2892 6625 2924
rect 6657 2892 6759 2924
rect 6523 2856 6759 2892
rect 6523 2824 6625 2856
rect 6657 2824 6759 2856
rect 6523 2788 6759 2824
rect 6523 2756 6625 2788
rect 6657 2756 6759 2788
rect 6523 2720 6759 2756
rect 6523 2688 6625 2720
rect 6657 2688 6759 2720
rect 6523 2652 6759 2688
rect 6523 2620 6625 2652
rect 6657 2620 6759 2652
rect 6523 2584 6759 2620
rect 6523 2552 6625 2584
rect 6657 2552 6759 2584
rect 6523 2516 6759 2552
rect 6523 2484 6625 2516
rect 6657 2484 6759 2516
rect 6523 2448 6759 2484
rect 6523 2416 6625 2448
rect 6657 2416 6759 2448
rect 6523 2380 6759 2416
rect 6523 2348 6625 2380
rect 6657 2348 6759 2380
rect 6523 2312 6759 2348
rect 6523 2280 6625 2312
rect 6657 2280 6759 2312
rect 6523 2244 6759 2280
rect 6523 2212 6625 2244
rect 6657 2212 6759 2244
rect 6523 2176 6759 2212
rect 6523 2144 6625 2176
rect 6657 2144 6759 2176
rect 6523 2108 6759 2144
rect 6523 2076 6625 2108
rect 6657 2076 6759 2108
rect 6523 2040 6759 2076
rect 6523 2008 6625 2040
rect 6657 2008 6759 2040
rect 6523 1970 6759 2008
rect 6879 3264 7007 3302
rect 6879 3232 6927 3264
rect 6959 3232 7007 3264
rect 6879 3196 7007 3232
rect 6879 3164 6927 3196
rect 6959 3164 7007 3196
rect 6879 3128 7007 3164
rect 6879 3096 6927 3128
rect 6959 3096 7007 3128
rect 6879 3060 7007 3096
rect 6879 3028 6927 3060
rect 6959 3028 7007 3060
rect 6879 2992 7007 3028
rect 6879 2960 6927 2992
rect 6959 2960 7007 2992
rect 6879 2924 7007 2960
rect 6879 2892 6927 2924
rect 6959 2892 7007 2924
rect 6879 2856 7007 2892
rect 6879 2824 6927 2856
rect 6959 2824 7007 2856
rect 6879 2788 7007 2824
rect 6879 2756 6927 2788
rect 6959 2756 7007 2788
rect 6879 2720 7007 2756
rect 6879 2688 6927 2720
rect 6959 2688 7007 2720
rect 6879 2652 7007 2688
rect 6879 2620 6927 2652
rect 6959 2620 7007 2652
rect 6879 2584 7007 2620
rect 6879 2552 6927 2584
rect 6959 2552 7007 2584
rect 6879 2516 7007 2552
rect 6879 2484 6927 2516
rect 6959 2484 7007 2516
rect 6879 2448 7007 2484
rect 6879 2416 6927 2448
rect 6959 2416 7007 2448
rect 6879 2380 7007 2416
rect 6879 2348 6927 2380
rect 6959 2348 7007 2380
rect 6879 2312 7007 2348
rect 6879 2280 6927 2312
rect 6959 2280 7007 2312
rect 6879 2244 7007 2280
rect 6879 2212 6927 2244
rect 6959 2212 7007 2244
rect 6879 2176 7007 2212
rect 6879 2144 6927 2176
rect 6959 2144 7007 2176
rect 6879 2108 7007 2144
rect 6879 2076 6927 2108
rect 6959 2076 7007 2108
rect 6879 2040 7007 2076
rect 6879 2008 6927 2040
rect 6959 2008 7007 2040
rect 6879 1970 7007 2008
rect 7127 3264 7363 3302
rect 7127 3232 7229 3264
rect 7261 3232 7363 3264
rect 7127 3196 7363 3232
rect 7127 3164 7229 3196
rect 7261 3164 7363 3196
rect 7127 3128 7363 3164
rect 7127 3096 7229 3128
rect 7261 3096 7363 3128
rect 7127 3060 7363 3096
rect 7127 3028 7229 3060
rect 7261 3028 7363 3060
rect 7127 2992 7363 3028
rect 7127 2960 7229 2992
rect 7261 2960 7363 2992
rect 7127 2924 7363 2960
rect 7127 2892 7229 2924
rect 7261 2892 7363 2924
rect 7127 2856 7363 2892
rect 7127 2824 7229 2856
rect 7261 2824 7363 2856
rect 7127 2788 7363 2824
rect 7127 2756 7229 2788
rect 7261 2756 7363 2788
rect 7127 2720 7363 2756
rect 7127 2688 7229 2720
rect 7261 2688 7363 2720
rect 7127 2652 7363 2688
rect 7127 2620 7229 2652
rect 7261 2620 7363 2652
rect 7127 2584 7363 2620
rect 7127 2552 7229 2584
rect 7261 2552 7363 2584
rect 7127 2516 7363 2552
rect 7127 2484 7229 2516
rect 7261 2484 7363 2516
rect 7127 2448 7363 2484
rect 7127 2416 7229 2448
rect 7261 2416 7363 2448
rect 7127 2380 7363 2416
rect 7127 2348 7229 2380
rect 7261 2348 7363 2380
rect 7127 2312 7363 2348
rect 7127 2280 7229 2312
rect 7261 2280 7363 2312
rect 7127 2244 7363 2280
rect 7127 2212 7229 2244
rect 7261 2212 7363 2244
rect 7127 2176 7363 2212
rect 7127 2144 7229 2176
rect 7261 2144 7363 2176
rect 7127 2108 7363 2144
rect 7127 2076 7229 2108
rect 7261 2076 7363 2108
rect 7127 2040 7363 2076
rect 7127 2008 7229 2040
rect 7261 2008 7363 2040
rect 7127 1970 7363 2008
rect 7483 3264 7611 3302
rect 7483 3232 7531 3264
rect 7563 3232 7611 3264
rect 7483 3196 7611 3232
rect 7483 3164 7531 3196
rect 7563 3164 7611 3196
rect 7483 3128 7611 3164
rect 7483 3096 7531 3128
rect 7563 3096 7611 3128
rect 7483 3060 7611 3096
rect 7483 3028 7531 3060
rect 7563 3028 7611 3060
rect 7483 2992 7611 3028
rect 7483 2960 7531 2992
rect 7563 2960 7611 2992
rect 7483 2924 7611 2960
rect 7483 2892 7531 2924
rect 7563 2892 7611 2924
rect 7483 2856 7611 2892
rect 7483 2824 7531 2856
rect 7563 2824 7611 2856
rect 7483 2788 7611 2824
rect 7483 2756 7531 2788
rect 7563 2756 7611 2788
rect 7483 2720 7611 2756
rect 7483 2688 7531 2720
rect 7563 2688 7611 2720
rect 7483 2652 7611 2688
rect 7483 2620 7531 2652
rect 7563 2620 7611 2652
rect 7483 2584 7611 2620
rect 7483 2552 7531 2584
rect 7563 2552 7611 2584
rect 7483 2516 7611 2552
rect 7483 2484 7531 2516
rect 7563 2484 7611 2516
rect 7483 2448 7611 2484
rect 7483 2416 7531 2448
rect 7563 2416 7611 2448
rect 7483 2380 7611 2416
rect 7483 2348 7531 2380
rect 7563 2348 7611 2380
rect 7483 2312 7611 2348
rect 7483 2280 7531 2312
rect 7563 2280 7611 2312
rect 7483 2244 7611 2280
rect 7483 2212 7531 2244
rect 7563 2212 7611 2244
rect 7483 2176 7611 2212
rect 7483 2144 7531 2176
rect 7563 2144 7611 2176
rect 7483 2108 7611 2144
rect 7483 2076 7531 2108
rect 7563 2076 7611 2108
rect 7483 2040 7611 2076
rect 7483 2008 7531 2040
rect 7563 2008 7611 2040
rect 7483 1970 7611 2008
rect 7731 3264 7967 3302
rect 7731 3232 7833 3264
rect 7865 3232 7967 3264
rect 7731 3196 7967 3232
rect 7731 3164 7833 3196
rect 7865 3164 7967 3196
rect 7731 3128 7967 3164
rect 7731 3096 7833 3128
rect 7865 3096 7967 3128
rect 7731 3060 7967 3096
rect 7731 3028 7833 3060
rect 7865 3028 7967 3060
rect 7731 2992 7967 3028
rect 7731 2960 7833 2992
rect 7865 2960 7967 2992
rect 7731 2924 7967 2960
rect 7731 2892 7833 2924
rect 7865 2892 7967 2924
rect 7731 2856 7967 2892
rect 7731 2824 7833 2856
rect 7865 2824 7967 2856
rect 7731 2788 7967 2824
rect 7731 2756 7833 2788
rect 7865 2756 7967 2788
rect 7731 2720 7967 2756
rect 7731 2688 7833 2720
rect 7865 2688 7967 2720
rect 7731 2652 7967 2688
rect 7731 2620 7833 2652
rect 7865 2620 7967 2652
rect 7731 2584 7967 2620
rect 7731 2552 7833 2584
rect 7865 2552 7967 2584
rect 7731 2516 7967 2552
rect 7731 2484 7833 2516
rect 7865 2484 7967 2516
rect 7731 2448 7967 2484
rect 7731 2416 7833 2448
rect 7865 2416 7967 2448
rect 7731 2380 7967 2416
rect 7731 2348 7833 2380
rect 7865 2348 7967 2380
rect 7731 2312 7967 2348
rect 7731 2280 7833 2312
rect 7865 2280 7967 2312
rect 7731 2244 7967 2280
rect 7731 2212 7833 2244
rect 7865 2212 7967 2244
rect 7731 2176 7967 2212
rect 7731 2144 7833 2176
rect 7865 2144 7967 2176
rect 7731 2108 7967 2144
rect 7731 2076 7833 2108
rect 7865 2076 7967 2108
rect 7731 2040 7967 2076
rect 7731 2008 7833 2040
rect 7865 2008 7967 2040
rect 7731 1970 7967 2008
rect 8087 3264 8215 3302
rect 8087 3232 8135 3264
rect 8167 3232 8215 3264
rect 8087 3196 8215 3232
rect 8087 3164 8135 3196
rect 8167 3164 8215 3196
rect 8087 3128 8215 3164
rect 8087 3096 8135 3128
rect 8167 3096 8215 3128
rect 8087 3060 8215 3096
rect 8087 3028 8135 3060
rect 8167 3028 8215 3060
rect 8087 2992 8215 3028
rect 8087 2960 8135 2992
rect 8167 2960 8215 2992
rect 8087 2924 8215 2960
rect 8087 2892 8135 2924
rect 8167 2892 8215 2924
rect 8087 2856 8215 2892
rect 8087 2824 8135 2856
rect 8167 2824 8215 2856
rect 8087 2788 8215 2824
rect 8087 2756 8135 2788
rect 8167 2756 8215 2788
rect 8087 2720 8215 2756
rect 8087 2688 8135 2720
rect 8167 2688 8215 2720
rect 8087 2652 8215 2688
rect 8087 2620 8135 2652
rect 8167 2620 8215 2652
rect 8087 2584 8215 2620
rect 8087 2552 8135 2584
rect 8167 2552 8215 2584
rect 8087 2516 8215 2552
rect 8087 2484 8135 2516
rect 8167 2484 8215 2516
rect 8087 2448 8215 2484
rect 8087 2416 8135 2448
rect 8167 2416 8215 2448
rect 8087 2380 8215 2416
rect 8087 2348 8135 2380
rect 8167 2348 8215 2380
rect 8087 2312 8215 2348
rect 8087 2280 8135 2312
rect 8167 2280 8215 2312
rect 8087 2244 8215 2280
rect 8087 2212 8135 2244
rect 8167 2212 8215 2244
rect 8087 2176 8215 2212
rect 8087 2144 8135 2176
rect 8167 2144 8215 2176
rect 8087 2108 8215 2144
rect 8087 2076 8135 2108
rect 8167 2076 8215 2108
rect 8087 2040 8215 2076
rect 8087 2008 8135 2040
rect 8167 2008 8215 2040
rect 8087 1970 8215 2008
rect 8335 3264 8571 3302
rect 8335 3232 8437 3264
rect 8469 3232 8571 3264
rect 8335 3196 8571 3232
rect 8335 3164 8437 3196
rect 8469 3164 8571 3196
rect 8335 3128 8571 3164
rect 8335 3096 8437 3128
rect 8469 3096 8571 3128
rect 8335 3060 8571 3096
rect 8335 3028 8437 3060
rect 8469 3028 8571 3060
rect 8335 2992 8571 3028
rect 8335 2960 8437 2992
rect 8469 2960 8571 2992
rect 8335 2924 8571 2960
rect 8335 2892 8437 2924
rect 8469 2892 8571 2924
rect 8335 2856 8571 2892
rect 8335 2824 8437 2856
rect 8469 2824 8571 2856
rect 8335 2788 8571 2824
rect 8335 2756 8437 2788
rect 8469 2756 8571 2788
rect 8335 2720 8571 2756
rect 8335 2688 8437 2720
rect 8469 2688 8571 2720
rect 8335 2652 8571 2688
rect 8335 2620 8437 2652
rect 8469 2620 8571 2652
rect 8335 2584 8571 2620
rect 8335 2552 8437 2584
rect 8469 2552 8571 2584
rect 8335 2516 8571 2552
rect 8335 2484 8437 2516
rect 8469 2484 8571 2516
rect 8335 2448 8571 2484
rect 8335 2416 8437 2448
rect 8469 2416 8571 2448
rect 8335 2380 8571 2416
rect 8335 2348 8437 2380
rect 8469 2348 8571 2380
rect 8335 2312 8571 2348
rect 8335 2280 8437 2312
rect 8469 2280 8571 2312
rect 8335 2244 8571 2280
rect 8335 2212 8437 2244
rect 8469 2212 8571 2244
rect 8335 2176 8571 2212
rect 8335 2144 8437 2176
rect 8469 2144 8571 2176
rect 8335 2108 8571 2144
rect 8335 2076 8437 2108
rect 8469 2076 8571 2108
rect 8335 2040 8571 2076
rect 8335 2008 8437 2040
rect 8469 2008 8571 2040
rect 8335 1970 8571 2008
rect 8691 3264 8819 3302
rect 8691 3232 8739 3264
rect 8771 3232 8819 3264
rect 8691 3196 8819 3232
rect 8691 3164 8739 3196
rect 8771 3164 8819 3196
rect 8691 3128 8819 3164
rect 8691 3096 8739 3128
rect 8771 3096 8819 3128
rect 8691 3060 8819 3096
rect 8691 3028 8739 3060
rect 8771 3028 8819 3060
rect 8691 2992 8819 3028
rect 8691 2960 8739 2992
rect 8771 2960 8819 2992
rect 8691 2924 8819 2960
rect 8691 2892 8739 2924
rect 8771 2892 8819 2924
rect 8691 2856 8819 2892
rect 8691 2824 8739 2856
rect 8771 2824 8819 2856
rect 8691 2788 8819 2824
rect 8691 2756 8739 2788
rect 8771 2756 8819 2788
rect 8691 2720 8819 2756
rect 8691 2688 8739 2720
rect 8771 2688 8819 2720
rect 8691 2652 8819 2688
rect 8691 2620 8739 2652
rect 8771 2620 8819 2652
rect 8691 2584 8819 2620
rect 8691 2552 8739 2584
rect 8771 2552 8819 2584
rect 8691 2516 8819 2552
rect 8691 2484 8739 2516
rect 8771 2484 8819 2516
rect 8691 2448 8819 2484
rect 8691 2416 8739 2448
rect 8771 2416 8819 2448
rect 8691 2380 8819 2416
rect 8691 2348 8739 2380
rect 8771 2348 8819 2380
rect 8691 2312 8819 2348
rect 8691 2280 8739 2312
rect 8771 2280 8819 2312
rect 8691 2244 8819 2280
rect 8691 2212 8739 2244
rect 8771 2212 8819 2244
rect 8691 2176 8819 2212
rect 8691 2144 8739 2176
rect 8771 2144 8819 2176
rect 8691 2108 8819 2144
rect 8691 2076 8739 2108
rect 8771 2076 8819 2108
rect 8691 2040 8819 2076
rect 8691 2008 8739 2040
rect 8771 2008 8819 2040
rect 8691 1970 8819 2008
rect 8939 3264 9175 3302
rect 8939 3232 9041 3264
rect 9073 3232 9175 3264
rect 8939 3196 9175 3232
rect 8939 3164 9041 3196
rect 9073 3164 9175 3196
rect 8939 3128 9175 3164
rect 8939 3096 9041 3128
rect 9073 3096 9175 3128
rect 8939 3060 9175 3096
rect 8939 3028 9041 3060
rect 9073 3028 9175 3060
rect 8939 2992 9175 3028
rect 8939 2960 9041 2992
rect 9073 2960 9175 2992
rect 8939 2924 9175 2960
rect 8939 2892 9041 2924
rect 9073 2892 9175 2924
rect 8939 2856 9175 2892
rect 8939 2824 9041 2856
rect 9073 2824 9175 2856
rect 8939 2788 9175 2824
rect 8939 2756 9041 2788
rect 9073 2756 9175 2788
rect 8939 2720 9175 2756
rect 8939 2688 9041 2720
rect 9073 2688 9175 2720
rect 8939 2652 9175 2688
rect 8939 2620 9041 2652
rect 9073 2620 9175 2652
rect 8939 2584 9175 2620
rect 8939 2552 9041 2584
rect 9073 2552 9175 2584
rect 8939 2516 9175 2552
rect 8939 2484 9041 2516
rect 9073 2484 9175 2516
rect 8939 2448 9175 2484
rect 8939 2416 9041 2448
rect 9073 2416 9175 2448
rect 8939 2380 9175 2416
rect 8939 2348 9041 2380
rect 9073 2348 9175 2380
rect 8939 2312 9175 2348
rect 8939 2280 9041 2312
rect 9073 2280 9175 2312
rect 8939 2244 9175 2280
rect 8939 2212 9041 2244
rect 9073 2212 9175 2244
rect 8939 2176 9175 2212
rect 8939 2144 9041 2176
rect 9073 2144 9175 2176
rect 8939 2108 9175 2144
rect 8939 2076 9041 2108
rect 9073 2076 9175 2108
rect 8939 2040 9175 2076
rect 8939 2008 9041 2040
rect 9073 2008 9175 2040
rect 8939 1970 9175 2008
rect 9295 3264 9423 3302
rect 9295 3232 9343 3264
rect 9375 3232 9423 3264
rect 9295 3196 9423 3232
rect 9295 3164 9343 3196
rect 9375 3164 9423 3196
rect 9295 3128 9423 3164
rect 9295 3096 9343 3128
rect 9375 3096 9423 3128
rect 9295 3060 9423 3096
rect 9295 3028 9343 3060
rect 9375 3028 9423 3060
rect 9295 2992 9423 3028
rect 9295 2960 9343 2992
rect 9375 2960 9423 2992
rect 9295 2924 9423 2960
rect 9295 2892 9343 2924
rect 9375 2892 9423 2924
rect 9295 2856 9423 2892
rect 9295 2824 9343 2856
rect 9375 2824 9423 2856
rect 9295 2788 9423 2824
rect 9295 2756 9343 2788
rect 9375 2756 9423 2788
rect 9295 2720 9423 2756
rect 9295 2688 9343 2720
rect 9375 2688 9423 2720
rect 9295 2652 9423 2688
rect 9295 2620 9343 2652
rect 9375 2620 9423 2652
rect 9295 2584 9423 2620
rect 9295 2552 9343 2584
rect 9375 2552 9423 2584
rect 9295 2516 9423 2552
rect 9295 2484 9343 2516
rect 9375 2484 9423 2516
rect 9295 2448 9423 2484
rect 9295 2416 9343 2448
rect 9375 2416 9423 2448
rect 9295 2380 9423 2416
rect 9295 2348 9343 2380
rect 9375 2348 9423 2380
rect 9295 2312 9423 2348
rect 9295 2280 9343 2312
rect 9375 2280 9423 2312
rect 9295 2244 9423 2280
rect 9295 2212 9343 2244
rect 9375 2212 9423 2244
rect 9295 2176 9423 2212
rect 9295 2144 9343 2176
rect 9375 2144 9423 2176
rect 9295 2108 9423 2144
rect 9295 2076 9343 2108
rect 9375 2076 9423 2108
rect 9295 2040 9423 2076
rect 9295 2008 9343 2040
rect 9375 2008 9423 2040
rect 9295 1970 9423 2008
rect 9543 3264 9779 3302
rect 9543 3232 9645 3264
rect 9677 3232 9779 3264
rect 9543 3196 9779 3232
rect 9543 3164 9645 3196
rect 9677 3164 9779 3196
rect 9543 3128 9779 3164
rect 9543 3096 9645 3128
rect 9677 3096 9779 3128
rect 9543 3060 9779 3096
rect 9543 3028 9645 3060
rect 9677 3028 9779 3060
rect 9543 2992 9779 3028
rect 9543 2960 9645 2992
rect 9677 2960 9779 2992
rect 9543 2924 9779 2960
rect 9543 2892 9645 2924
rect 9677 2892 9779 2924
rect 9543 2856 9779 2892
rect 9543 2824 9645 2856
rect 9677 2824 9779 2856
rect 9543 2788 9779 2824
rect 9543 2756 9645 2788
rect 9677 2756 9779 2788
rect 9543 2720 9779 2756
rect 9543 2688 9645 2720
rect 9677 2688 9779 2720
rect 9543 2652 9779 2688
rect 9543 2620 9645 2652
rect 9677 2620 9779 2652
rect 9543 2584 9779 2620
rect 9543 2552 9645 2584
rect 9677 2552 9779 2584
rect 9543 2516 9779 2552
rect 9543 2484 9645 2516
rect 9677 2484 9779 2516
rect 9543 2448 9779 2484
rect 9543 2416 9645 2448
rect 9677 2416 9779 2448
rect 9543 2380 9779 2416
rect 9543 2348 9645 2380
rect 9677 2348 9779 2380
rect 9543 2312 9779 2348
rect 9543 2280 9645 2312
rect 9677 2280 9779 2312
rect 9543 2244 9779 2280
rect 9543 2212 9645 2244
rect 9677 2212 9779 2244
rect 9543 2176 9779 2212
rect 9543 2144 9645 2176
rect 9677 2144 9779 2176
rect 9543 2108 9779 2144
rect 9543 2076 9645 2108
rect 9677 2076 9779 2108
rect 9543 2040 9779 2076
rect 9543 2008 9645 2040
rect 9677 2008 9779 2040
rect 9543 1970 9779 2008
rect 9899 3264 10027 3302
rect 9899 3232 9947 3264
rect 9979 3232 10027 3264
rect 9899 3196 10027 3232
rect 9899 3164 9947 3196
rect 9979 3164 10027 3196
rect 9899 3128 10027 3164
rect 9899 3096 9947 3128
rect 9979 3096 10027 3128
rect 9899 3060 10027 3096
rect 9899 3028 9947 3060
rect 9979 3028 10027 3060
rect 9899 2992 10027 3028
rect 9899 2960 9947 2992
rect 9979 2960 10027 2992
rect 9899 2924 10027 2960
rect 9899 2892 9947 2924
rect 9979 2892 10027 2924
rect 9899 2856 10027 2892
rect 9899 2824 9947 2856
rect 9979 2824 10027 2856
rect 9899 2788 10027 2824
rect 9899 2756 9947 2788
rect 9979 2756 10027 2788
rect 9899 2720 10027 2756
rect 9899 2688 9947 2720
rect 9979 2688 10027 2720
rect 9899 2652 10027 2688
rect 9899 2620 9947 2652
rect 9979 2620 10027 2652
rect 9899 2584 10027 2620
rect 9899 2552 9947 2584
rect 9979 2552 10027 2584
rect 9899 2516 10027 2552
rect 9899 2484 9947 2516
rect 9979 2484 10027 2516
rect 9899 2448 10027 2484
rect 9899 2416 9947 2448
rect 9979 2416 10027 2448
rect 9899 2380 10027 2416
rect 9899 2348 9947 2380
rect 9979 2348 10027 2380
rect 9899 2312 10027 2348
rect 9899 2280 9947 2312
rect 9979 2280 10027 2312
rect 9899 2244 10027 2280
rect 9899 2212 9947 2244
rect 9979 2212 10027 2244
rect 9899 2176 10027 2212
rect 9899 2144 9947 2176
rect 9979 2144 10027 2176
rect 9899 2108 10027 2144
rect 9899 2076 9947 2108
rect 9979 2076 10027 2108
rect 9899 2040 10027 2076
rect 9899 2008 9947 2040
rect 9979 2008 10027 2040
rect 9899 1970 10027 2008
rect 10147 3264 10295 3302
rect 10147 3232 10249 3264
rect 10281 3232 10295 3264
rect 10147 3196 10295 3232
rect 10147 3164 10249 3196
rect 10281 3164 10295 3196
rect 10147 3128 10295 3164
rect 10147 3096 10249 3128
rect 10281 3096 10295 3128
rect 10147 3060 10295 3096
rect 10147 3028 10249 3060
rect 10281 3028 10295 3060
rect 10147 2992 10295 3028
rect 10147 2960 10249 2992
rect 10281 2960 10295 2992
rect 10147 2924 10295 2960
rect 10147 2892 10249 2924
rect 10281 2892 10295 2924
rect 10147 2856 10295 2892
rect 10147 2824 10249 2856
rect 10281 2824 10295 2856
rect 10147 2788 10295 2824
rect 10147 2756 10249 2788
rect 10281 2756 10295 2788
rect 10147 2720 10295 2756
rect 10147 2688 10249 2720
rect 10281 2688 10295 2720
rect 10147 2652 10295 2688
rect 10147 2620 10249 2652
rect 10281 2620 10295 2652
rect 10147 2584 10295 2620
rect 10147 2552 10249 2584
rect 10281 2552 10295 2584
rect 10147 2516 10295 2552
rect 10147 2484 10249 2516
rect 10281 2484 10295 2516
rect 10147 2448 10295 2484
rect 10147 2416 10249 2448
rect 10281 2416 10295 2448
rect 10147 2380 10295 2416
rect 10147 2348 10249 2380
rect 10281 2348 10295 2380
rect 10147 2312 10295 2348
rect 10147 2280 10249 2312
rect 10281 2280 10295 2312
rect 10147 2244 10295 2280
rect 10147 2212 10249 2244
rect 10281 2212 10295 2244
rect 10147 2176 10295 2212
rect 10147 2144 10249 2176
rect 10281 2144 10295 2176
rect 10147 2108 10295 2144
rect 10147 2076 10249 2108
rect 10281 2076 10295 2108
rect 10147 2040 10295 2076
rect 10147 2008 10249 2040
rect 10281 2008 10295 2040
rect 10147 1970 10295 2008
rect 5705 1844 5799 1882
rect 5705 1812 5719 1844
rect 5751 1812 5799 1844
rect 5705 1776 5799 1812
rect 5705 1744 5719 1776
rect 5751 1744 5799 1776
rect 5705 1708 5799 1744
rect 5705 1676 5719 1708
rect 5751 1676 5799 1708
rect 5705 1640 5799 1676
rect 5705 1608 5719 1640
rect 5751 1608 5799 1640
rect 5705 1572 5799 1608
rect 5705 1540 5719 1572
rect 5751 1540 5799 1572
rect 5705 1504 5799 1540
rect 5705 1472 5719 1504
rect 5751 1472 5799 1504
rect 5705 1436 5799 1472
rect 5705 1404 5719 1436
rect 5751 1404 5799 1436
rect 5705 1368 5799 1404
rect 5705 1336 5719 1368
rect 5751 1336 5799 1368
rect 5705 1300 5799 1336
rect 5705 1268 5719 1300
rect 5751 1268 5799 1300
rect 5705 1232 5799 1268
rect 5705 1200 5719 1232
rect 5751 1200 5799 1232
rect 5705 1164 5799 1200
rect 5705 1132 5719 1164
rect 5751 1132 5799 1164
rect 5705 1096 5799 1132
rect 5705 1064 5719 1096
rect 5751 1064 5799 1096
rect 5705 1028 5799 1064
rect 5705 996 5719 1028
rect 5751 996 5799 1028
rect 5705 960 5799 996
rect 5705 928 5719 960
rect 5751 928 5799 960
rect 5705 892 5799 928
rect 5705 860 5719 892
rect 5751 860 5799 892
rect 5705 824 5799 860
rect 5705 792 5719 824
rect 5751 792 5799 824
rect 5705 756 5799 792
rect 5705 724 5719 756
rect 5751 724 5799 756
rect 5705 688 5799 724
rect 5705 656 5719 688
rect 5751 656 5799 688
rect 5705 620 5799 656
rect 5705 588 5719 620
rect 5751 588 5799 620
rect 5705 550 5799 588
rect 5919 1844 6155 1882
rect 5919 1812 6021 1844
rect 6053 1812 6155 1844
rect 5919 1776 6155 1812
rect 5919 1744 6021 1776
rect 6053 1744 6155 1776
rect 5919 1708 6155 1744
rect 5919 1676 6021 1708
rect 6053 1676 6155 1708
rect 5919 1640 6155 1676
rect 5919 1608 6021 1640
rect 6053 1608 6155 1640
rect 5919 1572 6155 1608
rect 5919 1540 6021 1572
rect 6053 1540 6155 1572
rect 5919 1504 6155 1540
rect 5919 1472 6021 1504
rect 6053 1472 6155 1504
rect 5919 1436 6155 1472
rect 5919 1404 6021 1436
rect 6053 1404 6155 1436
rect 5919 1368 6155 1404
rect 5919 1336 6021 1368
rect 6053 1336 6155 1368
rect 5919 1300 6155 1336
rect 5919 1268 6021 1300
rect 6053 1268 6155 1300
rect 5919 1232 6155 1268
rect 5919 1200 6021 1232
rect 6053 1200 6155 1232
rect 5919 1164 6155 1200
rect 5919 1132 6021 1164
rect 6053 1132 6155 1164
rect 5919 1096 6155 1132
rect 5919 1064 6021 1096
rect 6053 1064 6155 1096
rect 5919 1028 6155 1064
rect 5919 996 6021 1028
rect 6053 996 6155 1028
rect 5919 960 6155 996
rect 5919 928 6021 960
rect 6053 928 6155 960
rect 5919 892 6155 928
rect 5919 860 6021 892
rect 6053 860 6155 892
rect 5919 824 6155 860
rect 5919 792 6021 824
rect 6053 792 6155 824
rect 5919 756 6155 792
rect 5919 724 6021 756
rect 6053 724 6155 756
rect 5919 688 6155 724
rect 5919 656 6021 688
rect 6053 656 6155 688
rect 5919 620 6155 656
rect 5919 588 6021 620
rect 6053 588 6155 620
rect 5919 550 6155 588
rect 6275 1844 6403 1882
rect 6275 1812 6323 1844
rect 6355 1812 6403 1844
rect 6275 1776 6403 1812
rect 6275 1744 6323 1776
rect 6355 1744 6403 1776
rect 6275 1708 6403 1744
rect 6275 1676 6323 1708
rect 6355 1676 6403 1708
rect 6275 1640 6403 1676
rect 6275 1608 6323 1640
rect 6355 1608 6403 1640
rect 6275 1572 6403 1608
rect 6275 1540 6323 1572
rect 6355 1540 6403 1572
rect 6275 1504 6403 1540
rect 6275 1472 6323 1504
rect 6355 1472 6403 1504
rect 6275 1436 6403 1472
rect 6275 1404 6323 1436
rect 6355 1404 6403 1436
rect 6275 1368 6403 1404
rect 6275 1336 6323 1368
rect 6355 1336 6403 1368
rect 6275 1300 6403 1336
rect 6275 1268 6323 1300
rect 6355 1268 6403 1300
rect 6275 1232 6403 1268
rect 6275 1200 6323 1232
rect 6355 1200 6403 1232
rect 6275 1164 6403 1200
rect 6275 1132 6323 1164
rect 6355 1132 6403 1164
rect 6275 1096 6403 1132
rect 6275 1064 6323 1096
rect 6355 1064 6403 1096
rect 6275 1028 6403 1064
rect 6275 996 6323 1028
rect 6355 996 6403 1028
rect 6275 960 6403 996
rect 6275 928 6323 960
rect 6355 928 6403 960
rect 6275 892 6403 928
rect 6275 860 6323 892
rect 6355 860 6403 892
rect 6275 824 6403 860
rect 6275 792 6323 824
rect 6355 792 6403 824
rect 6275 756 6403 792
rect 6275 724 6323 756
rect 6355 724 6403 756
rect 6275 688 6403 724
rect 6275 656 6323 688
rect 6355 656 6403 688
rect 6275 620 6403 656
rect 6275 588 6323 620
rect 6355 588 6403 620
rect 6275 550 6403 588
rect 6523 1844 6759 1882
rect 6523 1812 6625 1844
rect 6657 1812 6759 1844
rect 6523 1776 6759 1812
rect 6523 1744 6625 1776
rect 6657 1744 6759 1776
rect 6523 1708 6759 1744
rect 6523 1676 6625 1708
rect 6657 1676 6759 1708
rect 6523 1640 6759 1676
rect 6523 1608 6625 1640
rect 6657 1608 6759 1640
rect 6523 1572 6759 1608
rect 6523 1540 6625 1572
rect 6657 1540 6759 1572
rect 6523 1504 6759 1540
rect 6523 1472 6625 1504
rect 6657 1472 6759 1504
rect 6523 1436 6759 1472
rect 6523 1404 6625 1436
rect 6657 1404 6759 1436
rect 6523 1368 6759 1404
rect 6523 1336 6625 1368
rect 6657 1336 6759 1368
rect 6523 1300 6759 1336
rect 6523 1268 6625 1300
rect 6657 1268 6759 1300
rect 6523 1232 6759 1268
rect 6523 1200 6625 1232
rect 6657 1200 6759 1232
rect 6523 1164 6759 1200
rect 6523 1132 6625 1164
rect 6657 1132 6759 1164
rect 6523 1096 6759 1132
rect 6523 1064 6625 1096
rect 6657 1064 6759 1096
rect 6523 1028 6759 1064
rect 6523 996 6625 1028
rect 6657 996 6759 1028
rect 6523 960 6759 996
rect 6523 928 6625 960
rect 6657 928 6759 960
rect 6523 892 6759 928
rect 6523 860 6625 892
rect 6657 860 6759 892
rect 6523 824 6759 860
rect 6523 792 6625 824
rect 6657 792 6759 824
rect 6523 756 6759 792
rect 6523 724 6625 756
rect 6657 724 6759 756
rect 6523 688 6759 724
rect 6523 656 6625 688
rect 6657 656 6759 688
rect 6523 620 6759 656
rect 6523 588 6625 620
rect 6657 588 6759 620
rect 6523 550 6759 588
rect 6879 1844 7007 1882
rect 6879 1812 6927 1844
rect 6959 1812 7007 1844
rect 6879 1776 7007 1812
rect 6879 1744 6927 1776
rect 6959 1744 7007 1776
rect 6879 1708 7007 1744
rect 6879 1676 6927 1708
rect 6959 1676 7007 1708
rect 6879 1640 7007 1676
rect 6879 1608 6927 1640
rect 6959 1608 7007 1640
rect 6879 1572 7007 1608
rect 6879 1540 6927 1572
rect 6959 1540 7007 1572
rect 6879 1504 7007 1540
rect 6879 1472 6927 1504
rect 6959 1472 7007 1504
rect 6879 1436 7007 1472
rect 6879 1404 6927 1436
rect 6959 1404 7007 1436
rect 6879 1368 7007 1404
rect 6879 1336 6927 1368
rect 6959 1336 7007 1368
rect 6879 1300 7007 1336
rect 6879 1268 6927 1300
rect 6959 1268 7007 1300
rect 6879 1232 7007 1268
rect 6879 1200 6927 1232
rect 6959 1200 7007 1232
rect 6879 1164 7007 1200
rect 6879 1132 6927 1164
rect 6959 1132 7007 1164
rect 6879 1096 7007 1132
rect 6879 1064 6927 1096
rect 6959 1064 7007 1096
rect 6879 1028 7007 1064
rect 6879 996 6927 1028
rect 6959 996 7007 1028
rect 6879 960 7007 996
rect 6879 928 6927 960
rect 6959 928 7007 960
rect 6879 892 7007 928
rect 6879 860 6927 892
rect 6959 860 7007 892
rect 6879 824 7007 860
rect 6879 792 6927 824
rect 6959 792 7007 824
rect 6879 756 7007 792
rect 6879 724 6927 756
rect 6959 724 7007 756
rect 6879 688 7007 724
rect 6879 656 6927 688
rect 6959 656 7007 688
rect 6879 620 7007 656
rect 6879 588 6927 620
rect 6959 588 7007 620
rect 6879 550 7007 588
rect 7127 1844 7363 1882
rect 7127 1812 7229 1844
rect 7261 1812 7363 1844
rect 7127 1776 7363 1812
rect 7127 1744 7229 1776
rect 7261 1744 7363 1776
rect 7127 1708 7363 1744
rect 7127 1676 7229 1708
rect 7261 1676 7363 1708
rect 7127 1640 7363 1676
rect 7127 1608 7229 1640
rect 7261 1608 7363 1640
rect 7127 1572 7363 1608
rect 7127 1540 7229 1572
rect 7261 1540 7363 1572
rect 7127 1504 7363 1540
rect 7127 1472 7229 1504
rect 7261 1472 7363 1504
rect 7127 1436 7363 1472
rect 7127 1404 7229 1436
rect 7261 1404 7363 1436
rect 7127 1368 7363 1404
rect 7127 1336 7229 1368
rect 7261 1336 7363 1368
rect 7127 1300 7363 1336
rect 7127 1268 7229 1300
rect 7261 1268 7363 1300
rect 7127 1232 7363 1268
rect 7127 1200 7229 1232
rect 7261 1200 7363 1232
rect 7127 1164 7363 1200
rect 7127 1132 7229 1164
rect 7261 1132 7363 1164
rect 7127 1096 7363 1132
rect 7127 1064 7229 1096
rect 7261 1064 7363 1096
rect 7127 1028 7363 1064
rect 7127 996 7229 1028
rect 7261 996 7363 1028
rect 7127 960 7363 996
rect 7127 928 7229 960
rect 7261 928 7363 960
rect 7127 892 7363 928
rect 7127 860 7229 892
rect 7261 860 7363 892
rect 7127 824 7363 860
rect 7127 792 7229 824
rect 7261 792 7363 824
rect 7127 756 7363 792
rect 7127 724 7229 756
rect 7261 724 7363 756
rect 7127 688 7363 724
rect 7127 656 7229 688
rect 7261 656 7363 688
rect 7127 620 7363 656
rect 7127 588 7229 620
rect 7261 588 7363 620
rect 7127 550 7363 588
rect 7483 1844 7611 1882
rect 7483 1812 7531 1844
rect 7563 1812 7611 1844
rect 7483 1776 7611 1812
rect 7483 1744 7531 1776
rect 7563 1744 7611 1776
rect 7483 1708 7611 1744
rect 7483 1676 7531 1708
rect 7563 1676 7611 1708
rect 7483 1640 7611 1676
rect 7483 1608 7531 1640
rect 7563 1608 7611 1640
rect 7483 1572 7611 1608
rect 7483 1540 7531 1572
rect 7563 1540 7611 1572
rect 7483 1504 7611 1540
rect 7483 1472 7531 1504
rect 7563 1472 7611 1504
rect 7483 1436 7611 1472
rect 7483 1404 7531 1436
rect 7563 1404 7611 1436
rect 7483 1368 7611 1404
rect 7483 1336 7531 1368
rect 7563 1336 7611 1368
rect 7483 1300 7611 1336
rect 7483 1268 7531 1300
rect 7563 1268 7611 1300
rect 7483 1232 7611 1268
rect 7483 1200 7531 1232
rect 7563 1200 7611 1232
rect 7483 1164 7611 1200
rect 7483 1132 7531 1164
rect 7563 1132 7611 1164
rect 7483 1096 7611 1132
rect 7483 1064 7531 1096
rect 7563 1064 7611 1096
rect 7483 1028 7611 1064
rect 7483 996 7531 1028
rect 7563 996 7611 1028
rect 7483 960 7611 996
rect 7483 928 7531 960
rect 7563 928 7611 960
rect 7483 892 7611 928
rect 7483 860 7531 892
rect 7563 860 7611 892
rect 7483 824 7611 860
rect 7483 792 7531 824
rect 7563 792 7611 824
rect 7483 756 7611 792
rect 7483 724 7531 756
rect 7563 724 7611 756
rect 7483 688 7611 724
rect 7483 656 7531 688
rect 7563 656 7611 688
rect 7483 620 7611 656
rect 7483 588 7531 620
rect 7563 588 7611 620
rect 7483 550 7611 588
rect 7731 1844 7967 1882
rect 7731 1812 7833 1844
rect 7865 1812 7967 1844
rect 7731 1776 7967 1812
rect 7731 1744 7833 1776
rect 7865 1744 7967 1776
rect 7731 1708 7967 1744
rect 7731 1676 7833 1708
rect 7865 1676 7967 1708
rect 7731 1640 7967 1676
rect 7731 1608 7833 1640
rect 7865 1608 7967 1640
rect 7731 1572 7967 1608
rect 7731 1540 7833 1572
rect 7865 1540 7967 1572
rect 7731 1504 7967 1540
rect 7731 1472 7833 1504
rect 7865 1472 7967 1504
rect 7731 1436 7967 1472
rect 7731 1404 7833 1436
rect 7865 1404 7967 1436
rect 7731 1368 7967 1404
rect 7731 1336 7833 1368
rect 7865 1336 7967 1368
rect 7731 1300 7967 1336
rect 7731 1268 7833 1300
rect 7865 1268 7967 1300
rect 7731 1232 7967 1268
rect 7731 1200 7833 1232
rect 7865 1200 7967 1232
rect 7731 1164 7967 1200
rect 7731 1132 7833 1164
rect 7865 1132 7967 1164
rect 7731 1096 7967 1132
rect 7731 1064 7833 1096
rect 7865 1064 7967 1096
rect 7731 1028 7967 1064
rect 7731 996 7833 1028
rect 7865 996 7967 1028
rect 7731 960 7967 996
rect 7731 928 7833 960
rect 7865 928 7967 960
rect 7731 892 7967 928
rect 7731 860 7833 892
rect 7865 860 7967 892
rect 7731 824 7967 860
rect 7731 792 7833 824
rect 7865 792 7967 824
rect 7731 756 7967 792
rect 7731 724 7833 756
rect 7865 724 7967 756
rect 7731 688 7967 724
rect 7731 656 7833 688
rect 7865 656 7967 688
rect 7731 620 7967 656
rect 7731 588 7833 620
rect 7865 588 7967 620
rect 7731 550 7967 588
rect 8087 1844 8215 1882
rect 8087 1812 8135 1844
rect 8167 1812 8215 1844
rect 8087 1776 8215 1812
rect 8087 1744 8135 1776
rect 8167 1744 8215 1776
rect 8087 1708 8215 1744
rect 8087 1676 8135 1708
rect 8167 1676 8215 1708
rect 8087 1640 8215 1676
rect 8087 1608 8135 1640
rect 8167 1608 8215 1640
rect 8087 1572 8215 1608
rect 8087 1540 8135 1572
rect 8167 1540 8215 1572
rect 8087 1504 8215 1540
rect 8087 1472 8135 1504
rect 8167 1472 8215 1504
rect 8087 1436 8215 1472
rect 8087 1404 8135 1436
rect 8167 1404 8215 1436
rect 8087 1368 8215 1404
rect 8087 1336 8135 1368
rect 8167 1336 8215 1368
rect 8087 1300 8215 1336
rect 8087 1268 8135 1300
rect 8167 1268 8215 1300
rect 8087 1232 8215 1268
rect 8087 1200 8135 1232
rect 8167 1200 8215 1232
rect 8087 1164 8215 1200
rect 8087 1132 8135 1164
rect 8167 1132 8215 1164
rect 8087 1096 8215 1132
rect 8087 1064 8135 1096
rect 8167 1064 8215 1096
rect 8087 1028 8215 1064
rect 8087 996 8135 1028
rect 8167 996 8215 1028
rect 8087 960 8215 996
rect 8087 928 8135 960
rect 8167 928 8215 960
rect 8087 892 8215 928
rect 8087 860 8135 892
rect 8167 860 8215 892
rect 8087 824 8215 860
rect 8087 792 8135 824
rect 8167 792 8215 824
rect 8087 756 8215 792
rect 8087 724 8135 756
rect 8167 724 8215 756
rect 8087 688 8215 724
rect 8087 656 8135 688
rect 8167 656 8215 688
rect 8087 620 8215 656
rect 8087 588 8135 620
rect 8167 588 8215 620
rect 8087 550 8215 588
rect 8335 1844 8571 1882
rect 8335 1812 8437 1844
rect 8469 1812 8571 1844
rect 8335 1776 8571 1812
rect 8335 1744 8437 1776
rect 8469 1744 8571 1776
rect 8335 1708 8571 1744
rect 8335 1676 8437 1708
rect 8469 1676 8571 1708
rect 8335 1640 8571 1676
rect 8335 1608 8437 1640
rect 8469 1608 8571 1640
rect 8335 1572 8571 1608
rect 8335 1540 8437 1572
rect 8469 1540 8571 1572
rect 8335 1504 8571 1540
rect 8335 1472 8437 1504
rect 8469 1472 8571 1504
rect 8335 1436 8571 1472
rect 8335 1404 8437 1436
rect 8469 1404 8571 1436
rect 8335 1368 8571 1404
rect 8335 1336 8437 1368
rect 8469 1336 8571 1368
rect 8335 1300 8571 1336
rect 8335 1268 8437 1300
rect 8469 1268 8571 1300
rect 8335 1232 8571 1268
rect 8335 1200 8437 1232
rect 8469 1200 8571 1232
rect 8335 1164 8571 1200
rect 8335 1132 8437 1164
rect 8469 1132 8571 1164
rect 8335 1096 8571 1132
rect 8335 1064 8437 1096
rect 8469 1064 8571 1096
rect 8335 1028 8571 1064
rect 8335 996 8437 1028
rect 8469 996 8571 1028
rect 8335 960 8571 996
rect 8335 928 8437 960
rect 8469 928 8571 960
rect 8335 892 8571 928
rect 8335 860 8437 892
rect 8469 860 8571 892
rect 8335 824 8571 860
rect 8335 792 8437 824
rect 8469 792 8571 824
rect 8335 756 8571 792
rect 8335 724 8437 756
rect 8469 724 8571 756
rect 8335 688 8571 724
rect 8335 656 8437 688
rect 8469 656 8571 688
rect 8335 620 8571 656
rect 8335 588 8437 620
rect 8469 588 8571 620
rect 8335 550 8571 588
rect 8691 1844 8819 1882
rect 8691 1812 8739 1844
rect 8771 1812 8819 1844
rect 8691 1776 8819 1812
rect 8691 1744 8739 1776
rect 8771 1744 8819 1776
rect 8691 1708 8819 1744
rect 8691 1676 8739 1708
rect 8771 1676 8819 1708
rect 8691 1640 8819 1676
rect 8691 1608 8739 1640
rect 8771 1608 8819 1640
rect 8691 1572 8819 1608
rect 8691 1540 8739 1572
rect 8771 1540 8819 1572
rect 8691 1504 8819 1540
rect 8691 1472 8739 1504
rect 8771 1472 8819 1504
rect 8691 1436 8819 1472
rect 8691 1404 8739 1436
rect 8771 1404 8819 1436
rect 8691 1368 8819 1404
rect 8691 1336 8739 1368
rect 8771 1336 8819 1368
rect 8691 1300 8819 1336
rect 8691 1268 8739 1300
rect 8771 1268 8819 1300
rect 8691 1232 8819 1268
rect 8691 1200 8739 1232
rect 8771 1200 8819 1232
rect 8691 1164 8819 1200
rect 8691 1132 8739 1164
rect 8771 1132 8819 1164
rect 8691 1096 8819 1132
rect 8691 1064 8739 1096
rect 8771 1064 8819 1096
rect 8691 1028 8819 1064
rect 8691 996 8739 1028
rect 8771 996 8819 1028
rect 8691 960 8819 996
rect 8691 928 8739 960
rect 8771 928 8819 960
rect 8691 892 8819 928
rect 8691 860 8739 892
rect 8771 860 8819 892
rect 8691 824 8819 860
rect 8691 792 8739 824
rect 8771 792 8819 824
rect 8691 756 8819 792
rect 8691 724 8739 756
rect 8771 724 8819 756
rect 8691 688 8819 724
rect 8691 656 8739 688
rect 8771 656 8819 688
rect 8691 620 8819 656
rect 8691 588 8739 620
rect 8771 588 8819 620
rect 8691 550 8819 588
rect 8939 1844 9175 1882
rect 8939 1812 9041 1844
rect 9073 1812 9175 1844
rect 8939 1776 9175 1812
rect 8939 1744 9041 1776
rect 9073 1744 9175 1776
rect 8939 1708 9175 1744
rect 8939 1676 9041 1708
rect 9073 1676 9175 1708
rect 8939 1640 9175 1676
rect 8939 1608 9041 1640
rect 9073 1608 9175 1640
rect 8939 1572 9175 1608
rect 8939 1540 9041 1572
rect 9073 1540 9175 1572
rect 8939 1504 9175 1540
rect 8939 1472 9041 1504
rect 9073 1472 9175 1504
rect 8939 1436 9175 1472
rect 8939 1404 9041 1436
rect 9073 1404 9175 1436
rect 8939 1368 9175 1404
rect 8939 1336 9041 1368
rect 9073 1336 9175 1368
rect 8939 1300 9175 1336
rect 8939 1268 9041 1300
rect 9073 1268 9175 1300
rect 8939 1232 9175 1268
rect 8939 1200 9041 1232
rect 9073 1200 9175 1232
rect 8939 1164 9175 1200
rect 8939 1132 9041 1164
rect 9073 1132 9175 1164
rect 8939 1096 9175 1132
rect 8939 1064 9041 1096
rect 9073 1064 9175 1096
rect 8939 1028 9175 1064
rect 8939 996 9041 1028
rect 9073 996 9175 1028
rect 8939 960 9175 996
rect 8939 928 9041 960
rect 9073 928 9175 960
rect 8939 892 9175 928
rect 8939 860 9041 892
rect 9073 860 9175 892
rect 8939 824 9175 860
rect 8939 792 9041 824
rect 9073 792 9175 824
rect 8939 756 9175 792
rect 8939 724 9041 756
rect 9073 724 9175 756
rect 8939 688 9175 724
rect 8939 656 9041 688
rect 9073 656 9175 688
rect 8939 620 9175 656
rect 8939 588 9041 620
rect 9073 588 9175 620
rect 8939 550 9175 588
rect 9295 1844 9423 1882
rect 9295 1812 9343 1844
rect 9375 1812 9423 1844
rect 9295 1776 9423 1812
rect 9295 1744 9343 1776
rect 9375 1744 9423 1776
rect 9295 1708 9423 1744
rect 9295 1676 9343 1708
rect 9375 1676 9423 1708
rect 9295 1640 9423 1676
rect 9295 1608 9343 1640
rect 9375 1608 9423 1640
rect 9295 1572 9423 1608
rect 9295 1540 9343 1572
rect 9375 1540 9423 1572
rect 9295 1504 9423 1540
rect 9295 1472 9343 1504
rect 9375 1472 9423 1504
rect 9295 1436 9423 1472
rect 9295 1404 9343 1436
rect 9375 1404 9423 1436
rect 9295 1368 9423 1404
rect 9295 1336 9343 1368
rect 9375 1336 9423 1368
rect 9295 1300 9423 1336
rect 9295 1268 9343 1300
rect 9375 1268 9423 1300
rect 9295 1232 9423 1268
rect 9295 1200 9343 1232
rect 9375 1200 9423 1232
rect 9295 1164 9423 1200
rect 9295 1132 9343 1164
rect 9375 1132 9423 1164
rect 9295 1096 9423 1132
rect 9295 1064 9343 1096
rect 9375 1064 9423 1096
rect 9295 1028 9423 1064
rect 9295 996 9343 1028
rect 9375 996 9423 1028
rect 9295 960 9423 996
rect 9295 928 9343 960
rect 9375 928 9423 960
rect 9295 892 9423 928
rect 9295 860 9343 892
rect 9375 860 9423 892
rect 9295 824 9423 860
rect 9295 792 9343 824
rect 9375 792 9423 824
rect 9295 756 9423 792
rect 9295 724 9343 756
rect 9375 724 9423 756
rect 9295 688 9423 724
rect 9295 656 9343 688
rect 9375 656 9423 688
rect 9295 620 9423 656
rect 9295 588 9343 620
rect 9375 588 9423 620
rect 9295 550 9423 588
rect 9543 1844 9779 1882
rect 9543 1812 9645 1844
rect 9677 1812 9779 1844
rect 9543 1776 9779 1812
rect 9543 1744 9645 1776
rect 9677 1744 9779 1776
rect 9543 1708 9779 1744
rect 9543 1676 9645 1708
rect 9677 1676 9779 1708
rect 9543 1640 9779 1676
rect 9543 1608 9645 1640
rect 9677 1608 9779 1640
rect 9543 1572 9779 1608
rect 9543 1540 9645 1572
rect 9677 1540 9779 1572
rect 9543 1504 9779 1540
rect 9543 1472 9645 1504
rect 9677 1472 9779 1504
rect 9543 1436 9779 1472
rect 9543 1404 9645 1436
rect 9677 1404 9779 1436
rect 9543 1368 9779 1404
rect 9543 1336 9645 1368
rect 9677 1336 9779 1368
rect 9543 1300 9779 1336
rect 9543 1268 9645 1300
rect 9677 1268 9779 1300
rect 9543 1232 9779 1268
rect 9543 1200 9645 1232
rect 9677 1200 9779 1232
rect 9543 1164 9779 1200
rect 9543 1132 9645 1164
rect 9677 1132 9779 1164
rect 9543 1096 9779 1132
rect 9543 1064 9645 1096
rect 9677 1064 9779 1096
rect 9543 1028 9779 1064
rect 9543 996 9645 1028
rect 9677 996 9779 1028
rect 9543 960 9779 996
rect 9543 928 9645 960
rect 9677 928 9779 960
rect 9543 892 9779 928
rect 9543 860 9645 892
rect 9677 860 9779 892
rect 9543 824 9779 860
rect 9543 792 9645 824
rect 9677 792 9779 824
rect 9543 756 9779 792
rect 9543 724 9645 756
rect 9677 724 9779 756
rect 9543 688 9779 724
rect 9543 656 9645 688
rect 9677 656 9779 688
rect 9543 620 9779 656
rect 9543 588 9645 620
rect 9677 588 9779 620
rect 9543 550 9779 588
rect 9899 1844 10027 1882
rect 9899 1812 9947 1844
rect 9979 1812 10027 1844
rect 9899 1776 10027 1812
rect 9899 1744 9947 1776
rect 9979 1744 10027 1776
rect 9899 1708 10027 1744
rect 9899 1676 9947 1708
rect 9979 1676 10027 1708
rect 9899 1640 10027 1676
rect 9899 1608 9947 1640
rect 9979 1608 10027 1640
rect 9899 1572 10027 1608
rect 9899 1540 9947 1572
rect 9979 1540 10027 1572
rect 9899 1504 10027 1540
rect 9899 1472 9947 1504
rect 9979 1472 10027 1504
rect 9899 1436 10027 1472
rect 9899 1404 9947 1436
rect 9979 1404 10027 1436
rect 9899 1368 10027 1404
rect 9899 1336 9947 1368
rect 9979 1336 10027 1368
rect 9899 1300 10027 1336
rect 9899 1268 9947 1300
rect 9979 1268 10027 1300
rect 9899 1232 10027 1268
rect 9899 1200 9947 1232
rect 9979 1200 10027 1232
rect 9899 1164 10027 1200
rect 9899 1132 9947 1164
rect 9979 1132 10027 1164
rect 9899 1096 10027 1132
rect 9899 1064 9947 1096
rect 9979 1064 10027 1096
rect 9899 1028 10027 1064
rect 9899 996 9947 1028
rect 9979 996 10027 1028
rect 9899 960 10027 996
rect 9899 928 9947 960
rect 9979 928 10027 960
rect 9899 892 10027 928
rect 9899 860 9947 892
rect 9979 860 10027 892
rect 9899 824 10027 860
rect 9899 792 9947 824
rect 9979 792 10027 824
rect 9899 756 10027 792
rect 9899 724 9947 756
rect 9979 724 10027 756
rect 9899 688 10027 724
rect 9899 656 9947 688
rect 9979 656 10027 688
rect 9899 620 10027 656
rect 9899 588 9947 620
rect 9979 588 10027 620
rect 9899 550 10027 588
rect 10147 1844 10295 1882
rect 10147 1812 10249 1844
rect 10281 1812 10295 1844
rect 10147 1776 10295 1812
rect 10147 1744 10249 1776
rect 10281 1744 10295 1776
rect 10147 1708 10295 1744
rect 10147 1676 10249 1708
rect 10281 1676 10295 1708
rect 10147 1640 10295 1676
rect 10147 1608 10249 1640
rect 10281 1608 10295 1640
rect 10147 1572 10295 1608
rect 10147 1540 10249 1572
rect 10281 1540 10295 1572
rect 10147 1504 10295 1540
rect 10147 1472 10249 1504
rect 10281 1472 10295 1504
rect 10147 1436 10295 1472
rect 10147 1404 10249 1436
rect 10281 1404 10295 1436
rect 10147 1368 10295 1404
rect 10147 1336 10249 1368
rect 10281 1336 10295 1368
rect 10147 1300 10295 1336
rect 10147 1268 10249 1300
rect 10281 1268 10295 1300
rect 10147 1232 10295 1268
rect 10147 1200 10249 1232
rect 10281 1200 10295 1232
rect 10147 1164 10295 1200
rect 10147 1132 10249 1164
rect 10281 1132 10295 1164
rect 10147 1096 10295 1132
rect 10147 1064 10249 1096
rect 10281 1064 10295 1096
rect 10147 1028 10295 1064
rect 10147 996 10249 1028
rect 10281 996 10295 1028
rect 10147 960 10295 996
rect 10147 928 10249 960
rect 10281 928 10295 960
rect 10147 892 10295 928
rect 10147 860 10249 892
rect 10281 860 10295 892
rect 10147 824 10295 860
rect 10147 792 10249 824
rect 10281 792 10295 824
rect 10147 756 10295 792
rect 10147 724 10249 756
rect 10281 724 10295 756
rect 10147 688 10295 724
rect 10147 656 10249 688
rect 10281 656 10295 688
rect 10147 620 10295 656
rect 10147 588 10249 620
rect 10281 588 10295 620
rect 10147 550 10295 588
<< hvpdiffc >>
rect 5719 3232 5751 3264
rect 5719 3164 5751 3196
rect 5719 3096 5751 3128
rect 5719 3028 5751 3060
rect 5719 2960 5751 2992
rect 5719 2892 5751 2924
rect 5719 2824 5751 2856
rect 5719 2756 5751 2788
rect 5719 2688 5751 2720
rect 5719 2620 5751 2652
rect 5719 2552 5751 2584
rect 5719 2484 5751 2516
rect 5719 2416 5751 2448
rect 5719 2348 5751 2380
rect 5719 2280 5751 2312
rect 5719 2212 5751 2244
rect 5719 2144 5751 2176
rect 5719 2076 5751 2108
rect 5719 2008 5751 2040
rect 6021 3232 6053 3264
rect 6021 3164 6053 3196
rect 6021 3096 6053 3128
rect 6021 3028 6053 3060
rect 6021 2960 6053 2992
rect 6021 2892 6053 2924
rect 6021 2824 6053 2856
rect 6021 2756 6053 2788
rect 6021 2688 6053 2720
rect 6021 2620 6053 2652
rect 6021 2552 6053 2584
rect 6021 2484 6053 2516
rect 6021 2416 6053 2448
rect 6021 2348 6053 2380
rect 6021 2280 6053 2312
rect 6021 2212 6053 2244
rect 6021 2144 6053 2176
rect 6021 2076 6053 2108
rect 6021 2008 6053 2040
rect 6323 3232 6355 3264
rect 6323 3164 6355 3196
rect 6323 3096 6355 3128
rect 6323 3028 6355 3060
rect 6323 2960 6355 2992
rect 6323 2892 6355 2924
rect 6323 2824 6355 2856
rect 6323 2756 6355 2788
rect 6323 2688 6355 2720
rect 6323 2620 6355 2652
rect 6323 2552 6355 2584
rect 6323 2484 6355 2516
rect 6323 2416 6355 2448
rect 6323 2348 6355 2380
rect 6323 2280 6355 2312
rect 6323 2212 6355 2244
rect 6323 2144 6355 2176
rect 6323 2076 6355 2108
rect 6323 2008 6355 2040
rect 6625 3232 6657 3264
rect 6625 3164 6657 3196
rect 6625 3096 6657 3128
rect 6625 3028 6657 3060
rect 6625 2960 6657 2992
rect 6625 2892 6657 2924
rect 6625 2824 6657 2856
rect 6625 2756 6657 2788
rect 6625 2688 6657 2720
rect 6625 2620 6657 2652
rect 6625 2552 6657 2584
rect 6625 2484 6657 2516
rect 6625 2416 6657 2448
rect 6625 2348 6657 2380
rect 6625 2280 6657 2312
rect 6625 2212 6657 2244
rect 6625 2144 6657 2176
rect 6625 2076 6657 2108
rect 6625 2008 6657 2040
rect 6927 3232 6959 3264
rect 6927 3164 6959 3196
rect 6927 3096 6959 3128
rect 6927 3028 6959 3060
rect 6927 2960 6959 2992
rect 6927 2892 6959 2924
rect 6927 2824 6959 2856
rect 6927 2756 6959 2788
rect 6927 2688 6959 2720
rect 6927 2620 6959 2652
rect 6927 2552 6959 2584
rect 6927 2484 6959 2516
rect 6927 2416 6959 2448
rect 6927 2348 6959 2380
rect 6927 2280 6959 2312
rect 6927 2212 6959 2244
rect 6927 2144 6959 2176
rect 6927 2076 6959 2108
rect 6927 2008 6959 2040
rect 7229 3232 7261 3264
rect 7229 3164 7261 3196
rect 7229 3096 7261 3128
rect 7229 3028 7261 3060
rect 7229 2960 7261 2992
rect 7229 2892 7261 2924
rect 7229 2824 7261 2856
rect 7229 2756 7261 2788
rect 7229 2688 7261 2720
rect 7229 2620 7261 2652
rect 7229 2552 7261 2584
rect 7229 2484 7261 2516
rect 7229 2416 7261 2448
rect 7229 2348 7261 2380
rect 7229 2280 7261 2312
rect 7229 2212 7261 2244
rect 7229 2144 7261 2176
rect 7229 2076 7261 2108
rect 7229 2008 7261 2040
rect 7531 3232 7563 3264
rect 7531 3164 7563 3196
rect 7531 3096 7563 3128
rect 7531 3028 7563 3060
rect 7531 2960 7563 2992
rect 7531 2892 7563 2924
rect 7531 2824 7563 2856
rect 7531 2756 7563 2788
rect 7531 2688 7563 2720
rect 7531 2620 7563 2652
rect 7531 2552 7563 2584
rect 7531 2484 7563 2516
rect 7531 2416 7563 2448
rect 7531 2348 7563 2380
rect 7531 2280 7563 2312
rect 7531 2212 7563 2244
rect 7531 2144 7563 2176
rect 7531 2076 7563 2108
rect 7531 2008 7563 2040
rect 7833 3232 7865 3264
rect 7833 3164 7865 3196
rect 7833 3096 7865 3128
rect 7833 3028 7865 3060
rect 7833 2960 7865 2992
rect 7833 2892 7865 2924
rect 7833 2824 7865 2856
rect 7833 2756 7865 2788
rect 7833 2688 7865 2720
rect 7833 2620 7865 2652
rect 7833 2552 7865 2584
rect 7833 2484 7865 2516
rect 7833 2416 7865 2448
rect 7833 2348 7865 2380
rect 7833 2280 7865 2312
rect 7833 2212 7865 2244
rect 7833 2144 7865 2176
rect 7833 2076 7865 2108
rect 7833 2008 7865 2040
rect 8135 3232 8167 3264
rect 8135 3164 8167 3196
rect 8135 3096 8167 3128
rect 8135 3028 8167 3060
rect 8135 2960 8167 2992
rect 8135 2892 8167 2924
rect 8135 2824 8167 2856
rect 8135 2756 8167 2788
rect 8135 2688 8167 2720
rect 8135 2620 8167 2652
rect 8135 2552 8167 2584
rect 8135 2484 8167 2516
rect 8135 2416 8167 2448
rect 8135 2348 8167 2380
rect 8135 2280 8167 2312
rect 8135 2212 8167 2244
rect 8135 2144 8167 2176
rect 8135 2076 8167 2108
rect 8135 2008 8167 2040
rect 8437 3232 8469 3264
rect 8437 3164 8469 3196
rect 8437 3096 8469 3128
rect 8437 3028 8469 3060
rect 8437 2960 8469 2992
rect 8437 2892 8469 2924
rect 8437 2824 8469 2856
rect 8437 2756 8469 2788
rect 8437 2688 8469 2720
rect 8437 2620 8469 2652
rect 8437 2552 8469 2584
rect 8437 2484 8469 2516
rect 8437 2416 8469 2448
rect 8437 2348 8469 2380
rect 8437 2280 8469 2312
rect 8437 2212 8469 2244
rect 8437 2144 8469 2176
rect 8437 2076 8469 2108
rect 8437 2008 8469 2040
rect 8739 3232 8771 3264
rect 8739 3164 8771 3196
rect 8739 3096 8771 3128
rect 8739 3028 8771 3060
rect 8739 2960 8771 2992
rect 8739 2892 8771 2924
rect 8739 2824 8771 2856
rect 8739 2756 8771 2788
rect 8739 2688 8771 2720
rect 8739 2620 8771 2652
rect 8739 2552 8771 2584
rect 8739 2484 8771 2516
rect 8739 2416 8771 2448
rect 8739 2348 8771 2380
rect 8739 2280 8771 2312
rect 8739 2212 8771 2244
rect 8739 2144 8771 2176
rect 8739 2076 8771 2108
rect 8739 2008 8771 2040
rect 9041 3232 9073 3264
rect 9041 3164 9073 3196
rect 9041 3096 9073 3128
rect 9041 3028 9073 3060
rect 9041 2960 9073 2992
rect 9041 2892 9073 2924
rect 9041 2824 9073 2856
rect 9041 2756 9073 2788
rect 9041 2688 9073 2720
rect 9041 2620 9073 2652
rect 9041 2552 9073 2584
rect 9041 2484 9073 2516
rect 9041 2416 9073 2448
rect 9041 2348 9073 2380
rect 9041 2280 9073 2312
rect 9041 2212 9073 2244
rect 9041 2144 9073 2176
rect 9041 2076 9073 2108
rect 9041 2008 9073 2040
rect 9343 3232 9375 3264
rect 9343 3164 9375 3196
rect 9343 3096 9375 3128
rect 9343 3028 9375 3060
rect 9343 2960 9375 2992
rect 9343 2892 9375 2924
rect 9343 2824 9375 2856
rect 9343 2756 9375 2788
rect 9343 2688 9375 2720
rect 9343 2620 9375 2652
rect 9343 2552 9375 2584
rect 9343 2484 9375 2516
rect 9343 2416 9375 2448
rect 9343 2348 9375 2380
rect 9343 2280 9375 2312
rect 9343 2212 9375 2244
rect 9343 2144 9375 2176
rect 9343 2076 9375 2108
rect 9343 2008 9375 2040
rect 9645 3232 9677 3264
rect 9645 3164 9677 3196
rect 9645 3096 9677 3128
rect 9645 3028 9677 3060
rect 9645 2960 9677 2992
rect 9645 2892 9677 2924
rect 9645 2824 9677 2856
rect 9645 2756 9677 2788
rect 9645 2688 9677 2720
rect 9645 2620 9677 2652
rect 9645 2552 9677 2584
rect 9645 2484 9677 2516
rect 9645 2416 9677 2448
rect 9645 2348 9677 2380
rect 9645 2280 9677 2312
rect 9645 2212 9677 2244
rect 9645 2144 9677 2176
rect 9645 2076 9677 2108
rect 9645 2008 9677 2040
rect 9947 3232 9979 3264
rect 9947 3164 9979 3196
rect 9947 3096 9979 3128
rect 9947 3028 9979 3060
rect 9947 2960 9979 2992
rect 9947 2892 9979 2924
rect 9947 2824 9979 2856
rect 9947 2756 9979 2788
rect 9947 2688 9979 2720
rect 9947 2620 9979 2652
rect 9947 2552 9979 2584
rect 9947 2484 9979 2516
rect 9947 2416 9979 2448
rect 9947 2348 9979 2380
rect 9947 2280 9979 2312
rect 9947 2212 9979 2244
rect 9947 2144 9979 2176
rect 9947 2076 9979 2108
rect 9947 2008 9979 2040
rect 10249 3232 10281 3264
rect 10249 3164 10281 3196
rect 10249 3096 10281 3128
rect 10249 3028 10281 3060
rect 10249 2960 10281 2992
rect 10249 2892 10281 2924
rect 10249 2824 10281 2856
rect 10249 2756 10281 2788
rect 10249 2688 10281 2720
rect 10249 2620 10281 2652
rect 10249 2552 10281 2584
rect 10249 2484 10281 2516
rect 10249 2416 10281 2448
rect 10249 2348 10281 2380
rect 10249 2280 10281 2312
rect 10249 2212 10281 2244
rect 10249 2144 10281 2176
rect 10249 2076 10281 2108
rect 10249 2008 10281 2040
rect 5719 1812 5751 1844
rect 5719 1744 5751 1776
rect 5719 1676 5751 1708
rect 5719 1608 5751 1640
rect 5719 1540 5751 1572
rect 5719 1472 5751 1504
rect 5719 1404 5751 1436
rect 5719 1336 5751 1368
rect 5719 1268 5751 1300
rect 5719 1200 5751 1232
rect 5719 1132 5751 1164
rect 5719 1064 5751 1096
rect 5719 996 5751 1028
rect 5719 928 5751 960
rect 5719 860 5751 892
rect 5719 792 5751 824
rect 5719 724 5751 756
rect 5719 656 5751 688
rect 5719 588 5751 620
rect 6021 1812 6053 1844
rect 6021 1744 6053 1776
rect 6021 1676 6053 1708
rect 6021 1608 6053 1640
rect 6021 1540 6053 1572
rect 6021 1472 6053 1504
rect 6021 1404 6053 1436
rect 6021 1336 6053 1368
rect 6021 1268 6053 1300
rect 6021 1200 6053 1232
rect 6021 1132 6053 1164
rect 6021 1064 6053 1096
rect 6021 996 6053 1028
rect 6021 928 6053 960
rect 6021 860 6053 892
rect 6021 792 6053 824
rect 6021 724 6053 756
rect 6021 656 6053 688
rect 6021 588 6053 620
rect 6323 1812 6355 1844
rect 6323 1744 6355 1776
rect 6323 1676 6355 1708
rect 6323 1608 6355 1640
rect 6323 1540 6355 1572
rect 6323 1472 6355 1504
rect 6323 1404 6355 1436
rect 6323 1336 6355 1368
rect 6323 1268 6355 1300
rect 6323 1200 6355 1232
rect 6323 1132 6355 1164
rect 6323 1064 6355 1096
rect 6323 996 6355 1028
rect 6323 928 6355 960
rect 6323 860 6355 892
rect 6323 792 6355 824
rect 6323 724 6355 756
rect 6323 656 6355 688
rect 6323 588 6355 620
rect 6625 1812 6657 1844
rect 6625 1744 6657 1776
rect 6625 1676 6657 1708
rect 6625 1608 6657 1640
rect 6625 1540 6657 1572
rect 6625 1472 6657 1504
rect 6625 1404 6657 1436
rect 6625 1336 6657 1368
rect 6625 1268 6657 1300
rect 6625 1200 6657 1232
rect 6625 1132 6657 1164
rect 6625 1064 6657 1096
rect 6625 996 6657 1028
rect 6625 928 6657 960
rect 6625 860 6657 892
rect 6625 792 6657 824
rect 6625 724 6657 756
rect 6625 656 6657 688
rect 6625 588 6657 620
rect 6927 1812 6959 1844
rect 6927 1744 6959 1776
rect 6927 1676 6959 1708
rect 6927 1608 6959 1640
rect 6927 1540 6959 1572
rect 6927 1472 6959 1504
rect 6927 1404 6959 1436
rect 6927 1336 6959 1368
rect 6927 1268 6959 1300
rect 6927 1200 6959 1232
rect 6927 1132 6959 1164
rect 6927 1064 6959 1096
rect 6927 996 6959 1028
rect 6927 928 6959 960
rect 6927 860 6959 892
rect 6927 792 6959 824
rect 6927 724 6959 756
rect 6927 656 6959 688
rect 6927 588 6959 620
rect 7229 1812 7261 1844
rect 7229 1744 7261 1776
rect 7229 1676 7261 1708
rect 7229 1608 7261 1640
rect 7229 1540 7261 1572
rect 7229 1472 7261 1504
rect 7229 1404 7261 1436
rect 7229 1336 7261 1368
rect 7229 1268 7261 1300
rect 7229 1200 7261 1232
rect 7229 1132 7261 1164
rect 7229 1064 7261 1096
rect 7229 996 7261 1028
rect 7229 928 7261 960
rect 7229 860 7261 892
rect 7229 792 7261 824
rect 7229 724 7261 756
rect 7229 656 7261 688
rect 7229 588 7261 620
rect 7531 1812 7563 1844
rect 7531 1744 7563 1776
rect 7531 1676 7563 1708
rect 7531 1608 7563 1640
rect 7531 1540 7563 1572
rect 7531 1472 7563 1504
rect 7531 1404 7563 1436
rect 7531 1336 7563 1368
rect 7531 1268 7563 1300
rect 7531 1200 7563 1232
rect 7531 1132 7563 1164
rect 7531 1064 7563 1096
rect 7531 996 7563 1028
rect 7531 928 7563 960
rect 7531 860 7563 892
rect 7531 792 7563 824
rect 7531 724 7563 756
rect 7531 656 7563 688
rect 7531 588 7563 620
rect 7833 1812 7865 1844
rect 7833 1744 7865 1776
rect 7833 1676 7865 1708
rect 7833 1608 7865 1640
rect 7833 1540 7865 1572
rect 7833 1472 7865 1504
rect 7833 1404 7865 1436
rect 7833 1336 7865 1368
rect 7833 1268 7865 1300
rect 7833 1200 7865 1232
rect 7833 1132 7865 1164
rect 7833 1064 7865 1096
rect 7833 996 7865 1028
rect 7833 928 7865 960
rect 7833 860 7865 892
rect 7833 792 7865 824
rect 7833 724 7865 756
rect 7833 656 7865 688
rect 7833 588 7865 620
rect 8135 1812 8167 1844
rect 8135 1744 8167 1776
rect 8135 1676 8167 1708
rect 8135 1608 8167 1640
rect 8135 1540 8167 1572
rect 8135 1472 8167 1504
rect 8135 1404 8167 1436
rect 8135 1336 8167 1368
rect 8135 1268 8167 1300
rect 8135 1200 8167 1232
rect 8135 1132 8167 1164
rect 8135 1064 8167 1096
rect 8135 996 8167 1028
rect 8135 928 8167 960
rect 8135 860 8167 892
rect 8135 792 8167 824
rect 8135 724 8167 756
rect 8135 656 8167 688
rect 8135 588 8167 620
rect 8437 1812 8469 1844
rect 8437 1744 8469 1776
rect 8437 1676 8469 1708
rect 8437 1608 8469 1640
rect 8437 1540 8469 1572
rect 8437 1472 8469 1504
rect 8437 1404 8469 1436
rect 8437 1336 8469 1368
rect 8437 1268 8469 1300
rect 8437 1200 8469 1232
rect 8437 1132 8469 1164
rect 8437 1064 8469 1096
rect 8437 996 8469 1028
rect 8437 928 8469 960
rect 8437 860 8469 892
rect 8437 792 8469 824
rect 8437 724 8469 756
rect 8437 656 8469 688
rect 8437 588 8469 620
rect 8739 1812 8771 1844
rect 8739 1744 8771 1776
rect 8739 1676 8771 1708
rect 8739 1608 8771 1640
rect 8739 1540 8771 1572
rect 8739 1472 8771 1504
rect 8739 1404 8771 1436
rect 8739 1336 8771 1368
rect 8739 1268 8771 1300
rect 8739 1200 8771 1232
rect 8739 1132 8771 1164
rect 8739 1064 8771 1096
rect 8739 996 8771 1028
rect 8739 928 8771 960
rect 8739 860 8771 892
rect 8739 792 8771 824
rect 8739 724 8771 756
rect 8739 656 8771 688
rect 8739 588 8771 620
rect 9041 1812 9073 1844
rect 9041 1744 9073 1776
rect 9041 1676 9073 1708
rect 9041 1608 9073 1640
rect 9041 1540 9073 1572
rect 9041 1472 9073 1504
rect 9041 1404 9073 1436
rect 9041 1336 9073 1368
rect 9041 1268 9073 1300
rect 9041 1200 9073 1232
rect 9041 1132 9073 1164
rect 9041 1064 9073 1096
rect 9041 996 9073 1028
rect 9041 928 9073 960
rect 9041 860 9073 892
rect 9041 792 9073 824
rect 9041 724 9073 756
rect 9041 656 9073 688
rect 9041 588 9073 620
rect 9343 1812 9375 1844
rect 9343 1744 9375 1776
rect 9343 1676 9375 1708
rect 9343 1608 9375 1640
rect 9343 1540 9375 1572
rect 9343 1472 9375 1504
rect 9343 1404 9375 1436
rect 9343 1336 9375 1368
rect 9343 1268 9375 1300
rect 9343 1200 9375 1232
rect 9343 1132 9375 1164
rect 9343 1064 9375 1096
rect 9343 996 9375 1028
rect 9343 928 9375 960
rect 9343 860 9375 892
rect 9343 792 9375 824
rect 9343 724 9375 756
rect 9343 656 9375 688
rect 9343 588 9375 620
rect 9645 1812 9677 1844
rect 9645 1744 9677 1776
rect 9645 1676 9677 1708
rect 9645 1608 9677 1640
rect 9645 1540 9677 1572
rect 9645 1472 9677 1504
rect 9645 1404 9677 1436
rect 9645 1336 9677 1368
rect 9645 1268 9677 1300
rect 9645 1200 9677 1232
rect 9645 1132 9677 1164
rect 9645 1064 9677 1096
rect 9645 996 9677 1028
rect 9645 928 9677 960
rect 9645 860 9677 892
rect 9645 792 9677 824
rect 9645 724 9677 756
rect 9645 656 9677 688
rect 9645 588 9677 620
rect 9947 1812 9979 1844
rect 9947 1744 9979 1776
rect 9947 1676 9979 1708
rect 9947 1608 9979 1640
rect 9947 1540 9979 1572
rect 9947 1472 9979 1504
rect 9947 1404 9979 1436
rect 9947 1336 9979 1368
rect 9947 1268 9979 1300
rect 9947 1200 9979 1232
rect 9947 1132 9979 1164
rect 9947 1064 9979 1096
rect 9947 996 9979 1028
rect 9947 928 9979 960
rect 9947 860 9979 892
rect 9947 792 9979 824
rect 9947 724 9979 756
rect 9947 656 9979 688
rect 9947 588 9979 620
rect 10249 1812 10281 1844
rect 10249 1744 10281 1776
rect 10249 1676 10281 1708
rect 10249 1608 10281 1640
rect 10249 1540 10281 1572
rect 10249 1472 10281 1504
rect 10249 1404 10281 1436
rect 10249 1336 10281 1368
rect 10249 1268 10281 1300
rect 10249 1200 10281 1232
rect 10249 1132 10281 1164
rect 10249 1064 10281 1096
rect 10249 996 10281 1028
rect 10249 928 10281 960
rect 10249 860 10281 892
rect 10249 792 10281 824
rect 10249 724 10281 756
rect 10249 656 10281 688
rect 10249 588 10281 620
<< psubdiff >>
rect 0 3834 16000 3852
rect 0 3802 28 3834
rect 60 3802 96 3834
rect 128 3802 164 3834
rect 196 3802 232 3834
rect 264 3802 300 3834
rect 332 3802 368 3834
rect 400 3802 436 3834
rect 468 3802 504 3834
rect 536 3802 572 3834
rect 604 3802 640 3834
rect 672 3802 708 3834
rect 740 3802 776 3834
rect 808 3802 844 3834
rect 876 3802 912 3834
rect 944 3802 980 3834
rect 1012 3802 1048 3834
rect 1080 3802 1116 3834
rect 1148 3802 1184 3834
rect 1216 3802 1252 3834
rect 1284 3802 1320 3834
rect 1352 3802 1388 3834
rect 1420 3802 1456 3834
rect 1488 3802 1524 3834
rect 1556 3802 1592 3834
rect 1624 3802 1660 3834
rect 1692 3802 1728 3834
rect 1760 3802 1796 3834
rect 1828 3802 1864 3834
rect 1896 3802 1932 3834
rect 1964 3802 2000 3834
rect 2032 3802 2068 3834
rect 2100 3802 2136 3834
rect 2168 3802 2204 3834
rect 2236 3802 2272 3834
rect 2304 3802 2340 3834
rect 2372 3802 2408 3834
rect 2440 3802 2476 3834
rect 2508 3802 2544 3834
rect 2576 3802 2612 3834
rect 2644 3802 2680 3834
rect 2712 3802 2748 3834
rect 2780 3802 2816 3834
rect 2848 3802 2884 3834
rect 2916 3802 2952 3834
rect 2984 3802 3020 3834
rect 3052 3802 3088 3834
rect 3120 3802 3156 3834
rect 3188 3802 3224 3834
rect 3256 3802 3292 3834
rect 3324 3802 3360 3834
rect 3392 3802 3428 3834
rect 3460 3802 3496 3834
rect 3528 3802 3564 3834
rect 3596 3802 3632 3834
rect 3664 3802 3700 3834
rect 3732 3802 3768 3834
rect 3800 3802 3836 3834
rect 3868 3802 3904 3834
rect 3936 3802 3972 3834
rect 4004 3802 4040 3834
rect 4072 3802 4108 3834
rect 4140 3802 4176 3834
rect 4208 3802 4244 3834
rect 4276 3802 4312 3834
rect 4344 3802 4380 3834
rect 4412 3802 4448 3834
rect 4480 3802 4516 3834
rect 4548 3802 4584 3834
rect 4616 3802 4652 3834
rect 4684 3802 4720 3834
rect 4752 3802 4788 3834
rect 4820 3802 4856 3834
rect 4888 3802 4924 3834
rect 4956 3802 4992 3834
rect 5024 3802 5060 3834
rect 5092 3802 5128 3834
rect 5160 3802 5196 3834
rect 5228 3802 5264 3834
rect 5296 3802 5332 3834
rect 5364 3802 5400 3834
rect 5432 3802 5468 3834
rect 5500 3802 5536 3834
rect 5568 3802 5604 3834
rect 5636 3802 5672 3834
rect 5704 3802 5740 3834
rect 5772 3802 5808 3834
rect 5840 3802 5876 3834
rect 5908 3802 5944 3834
rect 5976 3802 6012 3834
rect 6044 3802 6080 3834
rect 6112 3802 6148 3834
rect 6180 3802 6216 3834
rect 6248 3802 6284 3834
rect 6316 3802 6352 3834
rect 6384 3802 6420 3834
rect 6452 3802 6488 3834
rect 6520 3802 6556 3834
rect 6588 3802 6624 3834
rect 6656 3802 6692 3834
rect 6724 3802 6760 3834
rect 6792 3802 6828 3834
rect 6860 3802 6896 3834
rect 6928 3802 6964 3834
rect 6996 3802 7032 3834
rect 7064 3802 7100 3834
rect 7132 3802 7168 3834
rect 7200 3802 7236 3834
rect 7268 3802 7304 3834
rect 7336 3802 7372 3834
rect 7404 3802 7440 3834
rect 7472 3802 7508 3834
rect 7540 3802 7576 3834
rect 7608 3802 7644 3834
rect 7676 3802 7712 3834
rect 7744 3802 7780 3834
rect 7812 3802 7848 3834
rect 7880 3802 7916 3834
rect 7948 3802 7984 3834
rect 8016 3802 8052 3834
rect 8084 3802 8120 3834
rect 8152 3802 8188 3834
rect 8220 3802 8256 3834
rect 8288 3802 8324 3834
rect 8356 3802 8392 3834
rect 8424 3802 8460 3834
rect 8492 3802 8528 3834
rect 8560 3802 8596 3834
rect 8628 3802 8664 3834
rect 8696 3802 8732 3834
rect 8764 3802 8800 3834
rect 8832 3802 8868 3834
rect 8900 3802 8936 3834
rect 8968 3802 9004 3834
rect 9036 3802 9072 3834
rect 9104 3802 9140 3834
rect 9172 3802 9208 3834
rect 9240 3802 9276 3834
rect 9308 3802 9344 3834
rect 9376 3802 9412 3834
rect 9444 3802 9480 3834
rect 9512 3802 9548 3834
rect 9580 3802 9616 3834
rect 9648 3802 9684 3834
rect 9716 3802 9752 3834
rect 9784 3802 9820 3834
rect 9852 3802 9888 3834
rect 9920 3802 9956 3834
rect 9988 3802 10024 3834
rect 10056 3802 10092 3834
rect 10124 3802 10160 3834
rect 10192 3802 10228 3834
rect 10260 3802 10296 3834
rect 10328 3802 10364 3834
rect 10396 3802 10432 3834
rect 10464 3802 10500 3834
rect 10532 3802 10568 3834
rect 10600 3802 10636 3834
rect 10668 3802 10704 3834
rect 10736 3802 10772 3834
rect 10804 3802 10840 3834
rect 10872 3802 10908 3834
rect 10940 3802 10976 3834
rect 11008 3802 11044 3834
rect 11076 3802 11112 3834
rect 11144 3802 11180 3834
rect 11212 3802 11248 3834
rect 11280 3802 11316 3834
rect 11348 3802 11384 3834
rect 11416 3802 11452 3834
rect 11484 3802 11520 3834
rect 11552 3802 11588 3834
rect 11620 3802 11656 3834
rect 11688 3802 11724 3834
rect 11756 3802 11792 3834
rect 11824 3802 11860 3834
rect 11892 3802 11928 3834
rect 11960 3802 11996 3834
rect 12028 3802 12064 3834
rect 12096 3802 12132 3834
rect 12164 3802 12200 3834
rect 12232 3802 12268 3834
rect 12300 3802 12336 3834
rect 12368 3802 12404 3834
rect 12436 3802 12472 3834
rect 12504 3802 12540 3834
rect 12572 3802 12608 3834
rect 12640 3802 12676 3834
rect 12708 3802 12744 3834
rect 12776 3802 12812 3834
rect 12844 3802 12880 3834
rect 12912 3802 12948 3834
rect 12980 3802 13016 3834
rect 13048 3802 13084 3834
rect 13116 3802 13152 3834
rect 13184 3802 13220 3834
rect 13252 3802 13288 3834
rect 13320 3802 13356 3834
rect 13388 3802 13424 3834
rect 13456 3802 13492 3834
rect 13524 3802 13560 3834
rect 13592 3802 13628 3834
rect 13660 3802 13696 3834
rect 13728 3802 13764 3834
rect 13796 3802 13832 3834
rect 13864 3802 13900 3834
rect 13932 3802 13968 3834
rect 14000 3802 14036 3834
rect 14068 3802 14104 3834
rect 14136 3802 14172 3834
rect 14204 3802 14240 3834
rect 14272 3802 14308 3834
rect 14340 3802 14376 3834
rect 14408 3802 14444 3834
rect 14476 3802 14512 3834
rect 14544 3802 14580 3834
rect 14612 3802 14648 3834
rect 14680 3802 14716 3834
rect 14748 3802 14784 3834
rect 14816 3802 14852 3834
rect 14884 3802 14920 3834
rect 14952 3802 14988 3834
rect 15020 3802 15056 3834
rect 15088 3802 15124 3834
rect 15156 3802 15192 3834
rect 15224 3802 15260 3834
rect 15292 3802 15328 3834
rect 15360 3802 15396 3834
rect 15428 3802 15464 3834
rect 15496 3802 15532 3834
rect 15564 3802 15600 3834
rect 15632 3802 15668 3834
rect 15700 3802 15736 3834
rect 15768 3802 15804 3834
rect 15836 3802 15872 3834
rect 15904 3802 15940 3834
rect 15972 3802 16000 3834
rect 0 3784 16000 3802
rect 0 3744 68 3784
rect 0 3712 18 3744
rect 50 3712 68 3744
rect 0 3676 68 3712
rect 0 3644 18 3676
rect 50 3644 68 3676
rect 0 3608 68 3644
rect 0 3576 18 3608
rect 50 3576 68 3608
rect 0 3540 68 3576
rect 0 3508 18 3540
rect 50 3508 68 3540
rect 0 3472 68 3508
rect 15932 3744 16000 3784
rect 15932 3712 15950 3744
rect 15982 3712 16000 3744
rect 15932 3676 16000 3712
rect 15932 3644 15950 3676
rect 15982 3644 16000 3676
rect 15932 3608 16000 3644
rect 15932 3576 15950 3608
rect 15982 3576 16000 3608
rect 15932 3540 16000 3576
rect 15932 3508 15950 3540
rect 15982 3508 16000 3540
rect 0 3440 18 3472
rect 50 3440 68 3472
rect 0 3404 68 3440
rect 0 3372 18 3404
rect 50 3372 68 3404
rect 0 3336 68 3372
rect 0 3304 18 3336
rect 50 3304 68 3336
rect 0 3268 68 3304
rect 0 3236 18 3268
rect 50 3236 68 3268
rect 0 3200 68 3236
rect 0 3168 18 3200
rect 50 3168 68 3200
rect 0 3132 68 3168
rect 0 3100 18 3132
rect 50 3100 68 3132
rect 0 3064 68 3100
rect 0 3032 18 3064
rect 50 3032 68 3064
rect 0 2996 68 3032
rect 0 2964 18 2996
rect 50 2964 68 2996
rect 0 2928 68 2964
rect 0 2896 18 2928
rect 50 2896 68 2928
rect 0 2860 68 2896
rect 0 2828 18 2860
rect 50 2828 68 2860
rect 0 2792 68 2828
rect 0 2760 18 2792
rect 50 2760 68 2792
rect 0 2724 68 2760
rect 0 2692 18 2724
rect 50 2692 68 2724
rect 0 2656 68 2692
rect 0 2624 18 2656
rect 50 2624 68 2656
rect 0 2588 68 2624
rect 0 2556 18 2588
rect 50 2556 68 2588
rect 0 2520 68 2556
rect 0 2488 18 2520
rect 50 2488 68 2520
rect 0 2452 68 2488
rect 0 2420 18 2452
rect 50 2420 68 2452
rect 0 2384 68 2420
rect 0 2352 18 2384
rect 50 2352 68 2384
rect 0 2316 68 2352
rect 0 2284 18 2316
rect 50 2284 68 2316
rect 0 2248 68 2284
rect 0 2216 18 2248
rect 50 2216 68 2248
rect 0 2180 68 2216
rect 0 2148 18 2180
rect 50 2148 68 2180
rect 0 2112 68 2148
rect 0 2080 18 2112
rect 50 2080 68 2112
rect 0 2044 68 2080
rect 0 2012 18 2044
rect 50 2012 68 2044
rect 0 1976 68 2012
rect 0 1944 18 1976
rect 50 1944 68 1976
rect 0 1908 68 1944
rect 0 1876 18 1908
rect 50 1876 68 1908
rect 0 1840 68 1876
rect 0 1808 18 1840
rect 50 1808 68 1840
rect 0 1772 68 1808
rect 0 1740 18 1772
rect 50 1740 68 1772
rect 0 1704 68 1740
rect 0 1672 18 1704
rect 50 1672 68 1704
rect 0 1636 68 1672
rect 0 1604 18 1636
rect 50 1604 68 1636
rect 0 1568 68 1604
rect 0 1536 18 1568
rect 50 1536 68 1568
rect 0 1500 68 1536
rect 0 1468 18 1500
rect 50 1468 68 1500
rect 0 1432 68 1468
rect 0 1400 18 1432
rect 50 1400 68 1432
rect 0 1364 68 1400
rect 0 1332 18 1364
rect 50 1332 68 1364
rect 0 1296 68 1332
rect 0 1264 18 1296
rect 50 1264 68 1296
rect 0 1228 68 1264
rect 0 1196 18 1228
rect 50 1196 68 1228
rect 0 1160 68 1196
rect 0 1128 18 1160
rect 50 1128 68 1160
rect 0 1092 68 1128
rect 0 1060 18 1092
rect 50 1060 68 1092
rect 0 1024 68 1060
rect 0 992 18 1024
rect 50 992 68 1024
rect 0 956 68 992
rect 0 924 18 956
rect 50 924 68 956
rect 0 888 68 924
rect 0 856 18 888
rect 50 856 68 888
rect 0 820 68 856
rect 0 788 18 820
rect 50 788 68 820
rect 0 752 68 788
rect 0 720 18 752
rect 50 720 68 752
rect 0 684 68 720
rect 0 652 18 684
rect 50 652 68 684
rect 0 616 68 652
rect 0 584 18 616
rect 50 584 68 616
rect 0 548 68 584
rect 0 516 18 548
rect 50 516 68 548
rect 0 480 68 516
rect 0 448 18 480
rect 50 448 68 480
rect 0 412 68 448
rect 0 380 18 412
rect 50 380 68 412
rect 0 344 68 380
rect 15932 3472 16000 3508
rect 15932 3440 15950 3472
rect 15982 3440 16000 3472
rect 15932 3404 16000 3440
rect 15932 3372 15950 3404
rect 15982 3372 16000 3404
rect 15932 3336 16000 3372
rect 15932 3304 15950 3336
rect 15982 3304 16000 3336
rect 15932 3268 16000 3304
rect 15932 3236 15950 3268
rect 15982 3236 16000 3268
rect 15932 3200 16000 3236
rect 15932 3168 15950 3200
rect 15982 3168 16000 3200
rect 15932 3132 16000 3168
rect 15932 3100 15950 3132
rect 15982 3100 16000 3132
rect 15932 3064 16000 3100
rect 15932 3032 15950 3064
rect 15982 3032 16000 3064
rect 15932 2996 16000 3032
rect 15932 2964 15950 2996
rect 15982 2964 16000 2996
rect 15932 2928 16000 2964
rect 15932 2896 15950 2928
rect 15982 2896 16000 2928
rect 15932 2860 16000 2896
rect 15932 2828 15950 2860
rect 15982 2828 16000 2860
rect 15932 2792 16000 2828
rect 15932 2760 15950 2792
rect 15982 2760 16000 2792
rect 15932 2724 16000 2760
rect 15932 2692 15950 2724
rect 15982 2692 16000 2724
rect 15932 2656 16000 2692
rect 15932 2624 15950 2656
rect 15982 2624 16000 2656
rect 15932 2588 16000 2624
rect 15932 2556 15950 2588
rect 15982 2556 16000 2588
rect 15932 2520 16000 2556
rect 15932 2488 15950 2520
rect 15982 2488 16000 2520
rect 15932 2452 16000 2488
rect 15932 2420 15950 2452
rect 15982 2420 16000 2452
rect 15932 2384 16000 2420
rect 15932 2352 15950 2384
rect 15982 2352 16000 2384
rect 15932 2316 16000 2352
rect 15932 2284 15950 2316
rect 15982 2284 16000 2316
rect 15932 2248 16000 2284
rect 15932 2216 15950 2248
rect 15982 2216 16000 2248
rect 15932 2180 16000 2216
rect 15932 2148 15950 2180
rect 15982 2148 16000 2180
rect 15932 2112 16000 2148
rect 15932 2080 15950 2112
rect 15982 2080 16000 2112
rect 15932 2044 16000 2080
rect 15932 2012 15950 2044
rect 15982 2012 16000 2044
rect 15932 1976 16000 2012
rect 15932 1944 15950 1976
rect 15982 1944 16000 1976
rect 15932 1908 16000 1944
rect 15932 1876 15950 1908
rect 15982 1876 16000 1908
rect 15932 1840 16000 1876
rect 15932 1808 15950 1840
rect 15982 1808 16000 1840
rect 15932 1772 16000 1808
rect 15932 1740 15950 1772
rect 15982 1740 16000 1772
rect 15932 1704 16000 1740
rect 15932 1672 15950 1704
rect 15982 1672 16000 1704
rect 15932 1636 16000 1672
rect 15932 1604 15950 1636
rect 15982 1604 16000 1636
rect 15932 1568 16000 1604
rect 15932 1536 15950 1568
rect 15982 1536 16000 1568
rect 15932 1500 16000 1536
rect 15932 1468 15950 1500
rect 15982 1468 16000 1500
rect 15932 1432 16000 1468
rect 15932 1400 15950 1432
rect 15982 1400 16000 1432
rect 15932 1364 16000 1400
rect 15932 1332 15950 1364
rect 15982 1332 16000 1364
rect 15932 1296 16000 1332
rect 15932 1264 15950 1296
rect 15982 1264 16000 1296
rect 15932 1228 16000 1264
rect 15932 1196 15950 1228
rect 15982 1196 16000 1228
rect 15932 1160 16000 1196
rect 15932 1128 15950 1160
rect 15982 1128 16000 1160
rect 15932 1092 16000 1128
rect 15932 1060 15950 1092
rect 15982 1060 16000 1092
rect 15932 1024 16000 1060
rect 15932 992 15950 1024
rect 15982 992 16000 1024
rect 15932 956 16000 992
rect 15932 924 15950 956
rect 15982 924 16000 956
rect 15932 888 16000 924
rect 15932 856 15950 888
rect 15982 856 16000 888
rect 15932 820 16000 856
rect 15932 788 15950 820
rect 15982 788 16000 820
rect 15932 752 16000 788
rect 15932 720 15950 752
rect 15982 720 16000 752
rect 15932 684 16000 720
rect 15932 652 15950 684
rect 15982 652 16000 684
rect 15932 616 16000 652
rect 15932 584 15950 616
rect 15982 584 16000 616
rect 15932 548 16000 584
rect 15932 516 15950 548
rect 15982 516 16000 548
rect 15932 480 16000 516
rect 15932 448 15950 480
rect 15982 448 16000 480
rect 15932 412 16000 448
rect 15932 380 15950 412
rect 15982 380 16000 412
rect 0 312 18 344
rect 50 312 68 344
rect 0 276 68 312
rect 0 244 18 276
rect 50 244 68 276
rect 0 208 68 244
rect 0 176 18 208
rect 50 176 68 208
rect 0 140 68 176
rect 0 108 18 140
rect 50 108 68 140
rect 0 68 68 108
rect 15932 344 16000 380
rect 15932 312 15950 344
rect 15982 312 16000 344
rect 15932 276 16000 312
rect 15932 244 15950 276
rect 15982 244 16000 276
rect 15932 208 16000 244
rect 15932 176 15950 208
rect 15982 176 16000 208
rect 15932 140 16000 176
rect 15932 108 15950 140
rect 15982 108 16000 140
rect 15932 68 16000 108
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< nsubdiff >>
rect 360 3474 15640 3492
rect 360 3442 402 3474
rect 434 3442 470 3474
rect 502 3442 538 3474
rect 570 3442 606 3474
rect 638 3442 674 3474
rect 706 3442 742 3474
rect 774 3442 810 3474
rect 842 3442 878 3474
rect 910 3442 946 3474
rect 978 3442 1014 3474
rect 1046 3442 1082 3474
rect 1114 3442 1150 3474
rect 1182 3442 1218 3474
rect 1250 3442 1286 3474
rect 1318 3442 1354 3474
rect 1386 3442 1422 3474
rect 1454 3442 1490 3474
rect 1522 3442 1558 3474
rect 1590 3442 1626 3474
rect 1658 3442 1694 3474
rect 1726 3442 1762 3474
rect 1794 3442 1830 3474
rect 1862 3442 1898 3474
rect 1930 3442 1966 3474
rect 1998 3442 2034 3474
rect 2066 3442 2102 3474
rect 2134 3442 2170 3474
rect 2202 3442 2238 3474
rect 2270 3442 2306 3474
rect 2338 3442 2374 3474
rect 2406 3442 2442 3474
rect 2474 3442 2510 3474
rect 2542 3442 2578 3474
rect 2610 3442 2646 3474
rect 2678 3442 2714 3474
rect 2746 3442 2782 3474
rect 2814 3442 2850 3474
rect 2882 3442 2918 3474
rect 2950 3442 2986 3474
rect 3018 3442 3054 3474
rect 3086 3442 3122 3474
rect 3154 3442 3190 3474
rect 3222 3442 3258 3474
rect 3290 3442 3326 3474
rect 3358 3442 3394 3474
rect 3426 3442 3462 3474
rect 3494 3442 3530 3474
rect 3562 3442 3598 3474
rect 3630 3442 3666 3474
rect 3698 3442 3734 3474
rect 3766 3442 3802 3474
rect 3834 3442 3870 3474
rect 3902 3442 3938 3474
rect 3970 3442 4006 3474
rect 4038 3442 4074 3474
rect 4106 3442 4142 3474
rect 4174 3442 4210 3474
rect 4242 3442 4278 3474
rect 4310 3442 4346 3474
rect 4378 3442 4414 3474
rect 4446 3442 4482 3474
rect 4514 3442 4550 3474
rect 4582 3442 4618 3474
rect 4650 3442 4686 3474
rect 4718 3442 4754 3474
rect 4786 3442 4822 3474
rect 4854 3442 4890 3474
rect 4922 3442 4958 3474
rect 4990 3442 5026 3474
rect 5058 3442 5094 3474
rect 5126 3442 5162 3474
rect 5194 3442 5230 3474
rect 5262 3442 5298 3474
rect 5330 3442 5366 3474
rect 5398 3442 5434 3474
rect 5466 3442 5502 3474
rect 5534 3442 5570 3474
rect 5602 3442 5638 3474
rect 5670 3442 5706 3474
rect 5738 3442 5774 3474
rect 5806 3442 5842 3474
rect 5874 3442 5910 3474
rect 5942 3442 5978 3474
rect 6010 3442 6046 3474
rect 6078 3442 6114 3474
rect 6146 3442 6182 3474
rect 6214 3442 6250 3474
rect 6282 3442 6318 3474
rect 6350 3442 6386 3474
rect 6418 3442 6454 3474
rect 6486 3442 6522 3474
rect 6554 3442 6590 3474
rect 6622 3442 6658 3474
rect 6690 3442 6726 3474
rect 6758 3442 6794 3474
rect 6826 3442 6862 3474
rect 6894 3442 6930 3474
rect 6962 3442 6998 3474
rect 7030 3442 7066 3474
rect 7098 3442 7134 3474
rect 7166 3442 7202 3474
rect 7234 3442 7270 3474
rect 7302 3442 7338 3474
rect 7370 3442 7406 3474
rect 7438 3442 7474 3474
rect 7506 3442 7542 3474
rect 7574 3442 7610 3474
rect 7642 3442 7678 3474
rect 7710 3442 7746 3474
rect 7778 3442 7814 3474
rect 7846 3442 7882 3474
rect 7914 3442 7950 3474
rect 7982 3442 8018 3474
rect 8050 3442 8086 3474
rect 8118 3442 8154 3474
rect 8186 3442 8222 3474
rect 8254 3442 8290 3474
rect 8322 3442 8358 3474
rect 8390 3442 8426 3474
rect 8458 3442 8494 3474
rect 8526 3442 8562 3474
rect 8594 3442 8630 3474
rect 8662 3442 8698 3474
rect 8730 3442 8766 3474
rect 8798 3442 8834 3474
rect 8866 3442 8902 3474
rect 8934 3442 8970 3474
rect 9002 3442 9038 3474
rect 9070 3442 9106 3474
rect 9138 3442 9174 3474
rect 9206 3442 9242 3474
rect 9274 3442 9310 3474
rect 9342 3442 9378 3474
rect 9410 3442 9446 3474
rect 9478 3442 9514 3474
rect 9546 3442 9582 3474
rect 9614 3442 9650 3474
rect 9682 3442 9718 3474
rect 9750 3442 9786 3474
rect 9818 3442 9854 3474
rect 9886 3442 9922 3474
rect 9954 3442 9990 3474
rect 10022 3442 10058 3474
rect 10090 3442 10126 3474
rect 10158 3442 10194 3474
rect 10226 3442 10262 3474
rect 10294 3442 10330 3474
rect 10362 3442 10398 3474
rect 10430 3442 10466 3474
rect 10498 3442 10534 3474
rect 10566 3442 10602 3474
rect 10634 3442 10670 3474
rect 10702 3442 10738 3474
rect 10770 3442 10806 3474
rect 10838 3442 10874 3474
rect 10906 3442 10942 3474
rect 10974 3442 11010 3474
rect 11042 3442 11078 3474
rect 11110 3442 11146 3474
rect 11178 3442 11214 3474
rect 11246 3442 11282 3474
rect 11314 3442 11350 3474
rect 11382 3442 11418 3474
rect 11450 3442 11486 3474
rect 11518 3442 11554 3474
rect 11586 3442 11622 3474
rect 11654 3442 11690 3474
rect 11722 3442 11758 3474
rect 11790 3442 11826 3474
rect 11858 3442 11894 3474
rect 11926 3442 11962 3474
rect 11994 3442 12030 3474
rect 12062 3442 12098 3474
rect 12130 3442 12166 3474
rect 12198 3442 12234 3474
rect 12266 3442 12302 3474
rect 12334 3442 12370 3474
rect 12402 3442 12438 3474
rect 12470 3442 12506 3474
rect 12538 3442 12574 3474
rect 12606 3442 12642 3474
rect 12674 3442 12710 3474
rect 12742 3442 12778 3474
rect 12810 3442 12846 3474
rect 12878 3442 12914 3474
rect 12946 3442 12982 3474
rect 13014 3442 13050 3474
rect 13082 3442 13118 3474
rect 13150 3442 13186 3474
rect 13218 3442 13254 3474
rect 13286 3442 13322 3474
rect 13354 3442 13390 3474
rect 13422 3442 13458 3474
rect 13490 3442 13526 3474
rect 13558 3442 13594 3474
rect 13626 3442 13662 3474
rect 13694 3442 13730 3474
rect 13762 3442 13798 3474
rect 13830 3442 13866 3474
rect 13898 3442 13934 3474
rect 13966 3442 14002 3474
rect 14034 3442 14070 3474
rect 14102 3442 14138 3474
rect 14170 3442 14206 3474
rect 14238 3442 14274 3474
rect 14306 3442 14342 3474
rect 14374 3442 14410 3474
rect 14442 3442 14478 3474
rect 14510 3442 14546 3474
rect 14578 3442 14614 3474
rect 14646 3442 14682 3474
rect 14714 3442 14750 3474
rect 14782 3442 14818 3474
rect 14850 3442 14886 3474
rect 14918 3442 14954 3474
rect 14986 3442 15022 3474
rect 15054 3442 15090 3474
rect 15122 3442 15158 3474
rect 15190 3442 15226 3474
rect 15258 3442 15294 3474
rect 15326 3442 15362 3474
rect 15394 3442 15430 3474
rect 15462 3442 15498 3474
rect 15530 3442 15566 3474
rect 15598 3442 15640 3474
rect 360 3424 15640 3442
rect 360 3370 428 3424
rect 360 3338 378 3370
rect 410 3338 428 3370
rect 360 3302 428 3338
rect 15572 3370 15640 3424
rect 15572 3338 15590 3370
rect 15622 3338 15640 3370
rect 15572 3302 15640 3338
rect 360 3270 378 3302
rect 410 3270 428 3302
rect 360 3234 428 3270
rect 360 3202 378 3234
rect 410 3202 428 3234
rect 360 3166 428 3202
rect 360 3134 378 3166
rect 410 3134 428 3166
rect 360 3098 428 3134
rect 360 3066 378 3098
rect 410 3066 428 3098
rect 360 3030 428 3066
rect 360 2998 378 3030
rect 410 2998 428 3030
rect 360 2962 428 2998
rect 360 2930 378 2962
rect 410 2930 428 2962
rect 360 2894 428 2930
rect 360 2862 378 2894
rect 410 2862 428 2894
rect 360 2826 428 2862
rect 360 2794 378 2826
rect 410 2794 428 2826
rect 360 2758 428 2794
rect 360 2726 378 2758
rect 410 2726 428 2758
rect 360 2690 428 2726
rect 360 2658 378 2690
rect 410 2658 428 2690
rect 360 2622 428 2658
rect 360 2590 378 2622
rect 410 2590 428 2622
rect 360 2554 428 2590
rect 360 2522 378 2554
rect 410 2522 428 2554
rect 360 2486 428 2522
rect 360 2454 378 2486
rect 410 2454 428 2486
rect 360 2418 428 2454
rect 360 2386 378 2418
rect 410 2386 428 2418
rect 360 2350 428 2386
rect 360 2318 378 2350
rect 410 2318 428 2350
rect 360 2282 428 2318
rect 360 2250 378 2282
rect 410 2250 428 2282
rect 360 2214 428 2250
rect 360 2182 378 2214
rect 410 2182 428 2214
rect 360 2146 428 2182
rect 360 2114 378 2146
rect 410 2114 428 2146
rect 360 2078 428 2114
rect 360 2046 378 2078
rect 410 2046 428 2078
rect 360 2010 428 2046
rect 360 1978 378 2010
rect 410 1978 428 2010
rect 360 1942 428 1978
rect 15572 3270 15590 3302
rect 15622 3270 15640 3302
rect 15572 3234 15640 3270
rect 15572 3202 15590 3234
rect 15622 3202 15640 3234
rect 15572 3166 15640 3202
rect 15572 3134 15590 3166
rect 15622 3134 15640 3166
rect 15572 3098 15640 3134
rect 15572 3066 15590 3098
rect 15622 3066 15640 3098
rect 15572 3030 15640 3066
rect 15572 2998 15590 3030
rect 15622 2998 15640 3030
rect 15572 2962 15640 2998
rect 15572 2930 15590 2962
rect 15622 2930 15640 2962
rect 15572 2894 15640 2930
rect 15572 2862 15590 2894
rect 15622 2862 15640 2894
rect 15572 2826 15640 2862
rect 15572 2794 15590 2826
rect 15622 2794 15640 2826
rect 15572 2758 15640 2794
rect 15572 2726 15590 2758
rect 15622 2726 15640 2758
rect 15572 2690 15640 2726
rect 15572 2658 15590 2690
rect 15622 2658 15640 2690
rect 15572 2622 15640 2658
rect 15572 2590 15590 2622
rect 15622 2590 15640 2622
rect 15572 2554 15640 2590
rect 15572 2522 15590 2554
rect 15622 2522 15640 2554
rect 15572 2486 15640 2522
rect 15572 2454 15590 2486
rect 15622 2454 15640 2486
rect 15572 2418 15640 2454
rect 15572 2386 15590 2418
rect 15622 2386 15640 2418
rect 15572 2350 15640 2386
rect 15572 2318 15590 2350
rect 15622 2318 15640 2350
rect 15572 2282 15640 2318
rect 15572 2250 15590 2282
rect 15622 2250 15640 2282
rect 15572 2214 15640 2250
rect 15572 2182 15590 2214
rect 15622 2182 15640 2214
rect 15572 2146 15640 2182
rect 15572 2114 15590 2146
rect 15622 2114 15640 2146
rect 15572 2078 15640 2114
rect 15572 2046 15590 2078
rect 15622 2046 15640 2078
rect 15572 2010 15640 2046
rect 15572 1978 15590 2010
rect 15622 1978 15640 2010
rect 360 1910 378 1942
rect 410 1910 428 1942
rect 360 1874 428 1910
rect 15572 1942 15640 1978
rect 15572 1910 15590 1942
rect 15622 1910 15640 1942
rect 360 1842 378 1874
rect 410 1842 428 1874
rect 360 1806 428 1842
rect 360 1774 378 1806
rect 410 1774 428 1806
rect 360 1738 428 1774
rect 360 1706 378 1738
rect 410 1706 428 1738
rect 360 1670 428 1706
rect 360 1638 378 1670
rect 410 1638 428 1670
rect 360 1602 428 1638
rect 360 1570 378 1602
rect 410 1570 428 1602
rect 360 1534 428 1570
rect 360 1502 378 1534
rect 410 1502 428 1534
rect 360 1466 428 1502
rect 360 1434 378 1466
rect 410 1434 428 1466
rect 360 1398 428 1434
rect 360 1366 378 1398
rect 410 1366 428 1398
rect 360 1330 428 1366
rect 360 1298 378 1330
rect 410 1298 428 1330
rect 360 1262 428 1298
rect 360 1230 378 1262
rect 410 1230 428 1262
rect 360 1194 428 1230
rect 360 1162 378 1194
rect 410 1162 428 1194
rect 360 1126 428 1162
rect 360 1094 378 1126
rect 410 1094 428 1126
rect 360 1058 428 1094
rect 360 1026 378 1058
rect 410 1026 428 1058
rect 360 990 428 1026
rect 360 958 378 990
rect 410 958 428 990
rect 360 922 428 958
rect 360 890 378 922
rect 410 890 428 922
rect 360 854 428 890
rect 360 822 378 854
rect 410 822 428 854
rect 360 786 428 822
rect 360 754 378 786
rect 410 754 428 786
rect 360 718 428 754
rect 360 686 378 718
rect 410 686 428 718
rect 360 650 428 686
rect 360 618 378 650
rect 410 618 428 650
rect 360 582 428 618
rect 360 550 378 582
rect 410 550 428 582
rect 15572 1874 15640 1910
rect 15572 1842 15590 1874
rect 15622 1842 15640 1874
rect 15572 1806 15640 1842
rect 15572 1774 15590 1806
rect 15622 1774 15640 1806
rect 15572 1738 15640 1774
rect 15572 1706 15590 1738
rect 15622 1706 15640 1738
rect 15572 1670 15640 1706
rect 15572 1638 15590 1670
rect 15622 1638 15640 1670
rect 15572 1602 15640 1638
rect 15572 1570 15590 1602
rect 15622 1570 15640 1602
rect 15572 1534 15640 1570
rect 15572 1502 15590 1534
rect 15622 1502 15640 1534
rect 15572 1466 15640 1502
rect 15572 1434 15590 1466
rect 15622 1434 15640 1466
rect 15572 1398 15640 1434
rect 15572 1366 15590 1398
rect 15622 1366 15640 1398
rect 15572 1330 15640 1366
rect 15572 1298 15590 1330
rect 15622 1298 15640 1330
rect 15572 1262 15640 1298
rect 15572 1230 15590 1262
rect 15622 1230 15640 1262
rect 15572 1194 15640 1230
rect 15572 1162 15590 1194
rect 15622 1162 15640 1194
rect 15572 1126 15640 1162
rect 15572 1094 15590 1126
rect 15622 1094 15640 1126
rect 15572 1058 15640 1094
rect 15572 1026 15590 1058
rect 15622 1026 15640 1058
rect 15572 990 15640 1026
rect 15572 958 15590 990
rect 15622 958 15640 990
rect 15572 922 15640 958
rect 15572 890 15590 922
rect 15622 890 15640 922
rect 15572 854 15640 890
rect 15572 822 15590 854
rect 15622 822 15640 854
rect 15572 786 15640 822
rect 15572 754 15590 786
rect 15622 754 15640 786
rect 15572 718 15640 754
rect 15572 686 15590 718
rect 15622 686 15640 718
rect 15572 650 15640 686
rect 15572 618 15590 650
rect 15622 618 15640 650
rect 15572 582 15640 618
rect 15572 550 15590 582
rect 15622 550 15640 582
rect 360 514 428 550
rect 360 482 378 514
rect 410 482 428 514
rect 360 428 428 482
rect 15572 514 15640 550
rect 15572 482 15590 514
rect 15622 482 15640 514
rect 15572 428 15640 482
rect 360 410 15640 428
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 360 15640 378
<< psubdiffcont >>
rect 28 3802 60 3834
rect 96 3802 128 3834
rect 164 3802 196 3834
rect 232 3802 264 3834
rect 300 3802 332 3834
rect 368 3802 400 3834
rect 436 3802 468 3834
rect 504 3802 536 3834
rect 572 3802 604 3834
rect 640 3802 672 3834
rect 708 3802 740 3834
rect 776 3802 808 3834
rect 844 3802 876 3834
rect 912 3802 944 3834
rect 980 3802 1012 3834
rect 1048 3802 1080 3834
rect 1116 3802 1148 3834
rect 1184 3802 1216 3834
rect 1252 3802 1284 3834
rect 1320 3802 1352 3834
rect 1388 3802 1420 3834
rect 1456 3802 1488 3834
rect 1524 3802 1556 3834
rect 1592 3802 1624 3834
rect 1660 3802 1692 3834
rect 1728 3802 1760 3834
rect 1796 3802 1828 3834
rect 1864 3802 1896 3834
rect 1932 3802 1964 3834
rect 2000 3802 2032 3834
rect 2068 3802 2100 3834
rect 2136 3802 2168 3834
rect 2204 3802 2236 3834
rect 2272 3802 2304 3834
rect 2340 3802 2372 3834
rect 2408 3802 2440 3834
rect 2476 3802 2508 3834
rect 2544 3802 2576 3834
rect 2612 3802 2644 3834
rect 2680 3802 2712 3834
rect 2748 3802 2780 3834
rect 2816 3802 2848 3834
rect 2884 3802 2916 3834
rect 2952 3802 2984 3834
rect 3020 3802 3052 3834
rect 3088 3802 3120 3834
rect 3156 3802 3188 3834
rect 3224 3802 3256 3834
rect 3292 3802 3324 3834
rect 3360 3802 3392 3834
rect 3428 3802 3460 3834
rect 3496 3802 3528 3834
rect 3564 3802 3596 3834
rect 3632 3802 3664 3834
rect 3700 3802 3732 3834
rect 3768 3802 3800 3834
rect 3836 3802 3868 3834
rect 3904 3802 3936 3834
rect 3972 3802 4004 3834
rect 4040 3802 4072 3834
rect 4108 3802 4140 3834
rect 4176 3802 4208 3834
rect 4244 3802 4276 3834
rect 4312 3802 4344 3834
rect 4380 3802 4412 3834
rect 4448 3802 4480 3834
rect 4516 3802 4548 3834
rect 4584 3802 4616 3834
rect 4652 3802 4684 3834
rect 4720 3802 4752 3834
rect 4788 3802 4820 3834
rect 4856 3802 4888 3834
rect 4924 3802 4956 3834
rect 4992 3802 5024 3834
rect 5060 3802 5092 3834
rect 5128 3802 5160 3834
rect 5196 3802 5228 3834
rect 5264 3802 5296 3834
rect 5332 3802 5364 3834
rect 5400 3802 5432 3834
rect 5468 3802 5500 3834
rect 5536 3802 5568 3834
rect 5604 3802 5636 3834
rect 5672 3802 5704 3834
rect 5740 3802 5772 3834
rect 5808 3802 5840 3834
rect 5876 3802 5908 3834
rect 5944 3802 5976 3834
rect 6012 3802 6044 3834
rect 6080 3802 6112 3834
rect 6148 3802 6180 3834
rect 6216 3802 6248 3834
rect 6284 3802 6316 3834
rect 6352 3802 6384 3834
rect 6420 3802 6452 3834
rect 6488 3802 6520 3834
rect 6556 3802 6588 3834
rect 6624 3802 6656 3834
rect 6692 3802 6724 3834
rect 6760 3802 6792 3834
rect 6828 3802 6860 3834
rect 6896 3802 6928 3834
rect 6964 3802 6996 3834
rect 7032 3802 7064 3834
rect 7100 3802 7132 3834
rect 7168 3802 7200 3834
rect 7236 3802 7268 3834
rect 7304 3802 7336 3834
rect 7372 3802 7404 3834
rect 7440 3802 7472 3834
rect 7508 3802 7540 3834
rect 7576 3802 7608 3834
rect 7644 3802 7676 3834
rect 7712 3802 7744 3834
rect 7780 3802 7812 3834
rect 7848 3802 7880 3834
rect 7916 3802 7948 3834
rect 7984 3802 8016 3834
rect 8052 3802 8084 3834
rect 8120 3802 8152 3834
rect 8188 3802 8220 3834
rect 8256 3802 8288 3834
rect 8324 3802 8356 3834
rect 8392 3802 8424 3834
rect 8460 3802 8492 3834
rect 8528 3802 8560 3834
rect 8596 3802 8628 3834
rect 8664 3802 8696 3834
rect 8732 3802 8764 3834
rect 8800 3802 8832 3834
rect 8868 3802 8900 3834
rect 8936 3802 8968 3834
rect 9004 3802 9036 3834
rect 9072 3802 9104 3834
rect 9140 3802 9172 3834
rect 9208 3802 9240 3834
rect 9276 3802 9308 3834
rect 9344 3802 9376 3834
rect 9412 3802 9444 3834
rect 9480 3802 9512 3834
rect 9548 3802 9580 3834
rect 9616 3802 9648 3834
rect 9684 3802 9716 3834
rect 9752 3802 9784 3834
rect 9820 3802 9852 3834
rect 9888 3802 9920 3834
rect 9956 3802 9988 3834
rect 10024 3802 10056 3834
rect 10092 3802 10124 3834
rect 10160 3802 10192 3834
rect 10228 3802 10260 3834
rect 10296 3802 10328 3834
rect 10364 3802 10396 3834
rect 10432 3802 10464 3834
rect 10500 3802 10532 3834
rect 10568 3802 10600 3834
rect 10636 3802 10668 3834
rect 10704 3802 10736 3834
rect 10772 3802 10804 3834
rect 10840 3802 10872 3834
rect 10908 3802 10940 3834
rect 10976 3802 11008 3834
rect 11044 3802 11076 3834
rect 11112 3802 11144 3834
rect 11180 3802 11212 3834
rect 11248 3802 11280 3834
rect 11316 3802 11348 3834
rect 11384 3802 11416 3834
rect 11452 3802 11484 3834
rect 11520 3802 11552 3834
rect 11588 3802 11620 3834
rect 11656 3802 11688 3834
rect 11724 3802 11756 3834
rect 11792 3802 11824 3834
rect 11860 3802 11892 3834
rect 11928 3802 11960 3834
rect 11996 3802 12028 3834
rect 12064 3802 12096 3834
rect 12132 3802 12164 3834
rect 12200 3802 12232 3834
rect 12268 3802 12300 3834
rect 12336 3802 12368 3834
rect 12404 3802 12436 3834
rect 12472 3802 12504 3834
rect 12540 3802 12572 3834
rect 12608 3802 12640 3834
rect 12676 3802 12708 3834
rect 12744 3802 12776 3834
rect 12812 3802 12844 3834
rect 12880 3802 12912 3834
rect 12948 3802 12980 3834
rect 13016 3802 13048 3834
rect 13084 3802 13116 3834
rect 13152 3802 13184 3834
rect 13220 3802 13252 3834
rect 13288 3802 13320 3834
rect 13356 3802 13388 3834
rect 13424 3802 13456 3834
rect 13492 3802 13524 3834
rect 13560 3802 13592 3834
rect 13628 3802 13660 3834
rect 13696 3802 13728 3834
rect 13764 3802 13796 3834
rect 13832 3802 13864 3834
rect 13900 3802 13932 3834
rect 13968 3802 14000 3834
rect 14036 3802 14068 3834
rect 14104 3802 14136 3834
rect 14172 3802 14204 3834
rect 14240 3802 14272 3834
rect 14308 3802 14340 3834
rect 14376 3802 14408 3834
rect 14444 3802 14476 3834
rect 14512 3802 14544 3834
rect 14580 3802 14612 3834
rect 14648 3802 14680 3834
rect 14716 3802 14748 3834
rect 14784 3802 14816 3834
rect 14852 3802 14884 3834
rect 14920 3802 14952 3834
rect 14988 3802 15020 3834
rect 15056 3802 15088 3834
rect 15124 3802 15156 3834
rect 15192 3802 15224 3834
rect 15260 3802 15292 3834
rect 15328 3802 15360 3834
rect 15396 3802 15428 3834
rect 15464 3802 15496 3834
rect 15532 3802 15564 3834
rect 15600 3802 15632 3834
rect 15668 3802 15700 3834
rect 15736 3802 15768 3834
rect 15804 3802 15836 3834
rect 15872 3802 15904 3834
rect 15940 3802 15972 3834
rect 18 3712 50 3744
rect 18 3644 50 3676
rect 18 3576 50 3608
rect 18 3508 50 3540
rect 15950 3712 15982 3744
rect 15950 3644 15982 3676
rect 15950 3576 15982 3608
rect 15950 3508 15982 3540
rect 18 3440 50 3472
rect 18 3372 50 3404
rect 18 3304 50 3336
rect 18 3236 50 3268
rect 18 3168 50 3200
rect 18 3100 50 3132
rect 18 3032 50 3064
rect 18 2964 50 2996
rect 18 2896 50 2928
rect 18 2828 50 2860
rect 18 2760 50 2792
rect 18 2692 50 2724
rect 18 2624 50 2656
rect 18 2556 50 2588
rect 18 2488 50 2520
rect 18 2420 50 2452
rect 18 2352 50 2384
rect 18 2284 50 2316
rect 18 2216 50 2248
rect 18 2148 50 2180
rect 18 2080 50 2112
rect 18 2012 50 2044
rect 18 1944 50 1976
rect 18 1876 50 1908
rect 18 1808 50 1840
rect 18 1740 50 1772
rect 18 1672 50 1704
rect 18 1604 50 1636
rect 18 1536 50 1568
rect 18 1468 50 1500
rect 18 1400 50 1432
rect 18 1332 50 1364
rect 18 1264 50 1296
rect 18 1196 50 1228
rect 18 1128 50 1160
rect 18 1060 50 1092
rect 18 992 50 1024
rect 18 924 50 956
rect 18 856 50 888
rect 18 788 50 820
rect 18 720 50 752
rect 18 652 50 684
rect 18 584 50 616
rect 18 516 50 548
rect 18 448 50 480
rect 18 380 50 412
rect 15950 3440 15982 3472
rect 15950 3372 15982 3404
rect 15950 3304 15982 3336
rect 15950 3236 15982 3268
rect 15950 3168 15982 3200
rect 15950 3100 15982 3132
rect 15950 3032 15982 3064
rect 15950 2964 15982 2996
rect 15950 2896 15982 2928
rect 15950 2828 15982 2860
rect 15950 2760 15982 2792
rect 15950 2692 15982 2724
rect 15950 2624 15982 2656
rect 15950 2556 15982 2588
rect 15950 2488 15982 2520
rect 15950 2420 15982 2452
rect 15950 2352 15982 2384
rect 15950 2284 15982 2316
rect 15950 2216 15982 2248
rect 15950 2148 15982 2180
rect 15950 2080 15982 2112
rect 15950 2012 15982 2044
rect 15950 1944 15982 1976
rect 15950 1876 15982 1908
rect 15950 1808 15982 1840
rect 15950 1740 15982 1772
rect 15950 1672 15982 1704
rect 15950 1604 15982 1636
rect 15950 1536 15982 1568
rect 15950 1468 15982 1500
rect 15950 1400 15982 1432
rect 15950 1332 15982 1364
rect 15950 1264 15982 1296
rect 15950 1196 15982 1228
rect 15950 1128 15982 1160
rect 15950 1060 15982 1092
rect 15950 992 15982 1024
rect 15950 924 15982 956
rect 15950 856 15982 888
rect 15950 788 15982 820
rect 15950 720 15982 752
rect 15950 652 15982 684
rect 15950 584 15982 616
rect 15950 516 15982 548
rect 15950 448 15982 480
rect 15950 380 15982 412
rect 18 312 50 344
rect 18 244 50 276
rect 18 176 50 208
rect 18 108 50 140
rect 15950 312 15982 344
rect 15950 244 15982 276
rect 15950 176 15982 208
rect 15950 108 15982 140
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< nsubdiffcont >>
rect 402 3442 434 3474
rect 470 3442 502 3474
rect 538 3442 570 3474
rect 606 3442 638 3474
rect 674 3442 706 3474
rect 742 3442 774 3474
rect 810 3442 842 3474
rect 878 3442 910 3474
rect 946 3442 978 3474
rect 1014 3442 1046 3474
rect 1082 3442 1114 3474
rect 1150 3442 1182 3474
rect 1218 3442 1250 3474
rect 1286 3442 1318 3474
rect 1354 3442 1386 3474
rect 1422 3442 1454 3474
rect 1490 3442 1522 3474
rect 1558 3442 1590 3474
rect 1626 3442 1658 3474
rect 1694 3442 1726 3474
rect 1762 3442 1794 3474
rect 1830 3442 1862 3474
rect 1898 3442 1930 3474
rect 1966 3442 1998 3474
rect 2034 3442 2066 3474
rect 2102 3442 2134 3474
rect 2170 3442 2202 3474
rect 2238 3442 2270 3474
rect 2306 3442 2338 3474
rect 2374 3442 2406 3474
rect 2442 3442 2474 3474
rect 2510 3442 2542 3474
rect 2578 3442 2610 3474
rect 2646 3442 2678 3474
rect 2714 3442 2746 3474
rect 2782 3442 2814 3474
rect 2850 3442 2882 3474
rect 2918 3442 2950 3474
rect 2986 3442 3018 3474
rect 3054 3442 3086 3474
rect 3122 3442 3154 3474
rect 3190 3442 3222 3474
rect 3258 3442 3290 3474
rect 3326 3442 3358 3474
rect 3394 3442 3426 3474
rect 3462 3442 3494 3474
rect 3530 3442 3562 3474
rect 3598 3442 3630 3474
rect 3666 3442 3698 3474
rect 3734 3442 3766 3474
rect 3802 3442 3834 3474
rect 3870 3442 3902 3474
rect 3938 3442 3970 3474
rect 4006 3442 4038 3474
rect 4074 3442 4106 3474
rect 4142 3442 4174 3474
rect 4210 3442 4242 3474
rect 4278 3442 4310 3474
rect 4346 3442 4378 3474
rect 4414 3442 4446 3474
rect 4482 3442 4514 3474
rect 4550 3442 4582 3474
rect 4618 3442 4650 3474
rect 4686 3442 4718 3474
rect 4754 3442 4786 3474
rect 4822 3442 4854 3474
rect 4890 3442 4922 3474
rect 4958 3442 4990 3474
rect 5026 3442 5058 3474
rect 5094 3442 5126 3474
rect 5162 3442 5194 3474
rect 5230 3442 5262 3474
rect 5298 3442 5330 3474
rect 5366 3442 5398 3474
rect 5434 3442 5466 3474
rect 5502 3442 5534 3474
rect 5570 3442 5602 3474
rect 5638 3442 5670 3474
rect 5706 3442 5738 3474
rect 5774 3442 5806 3474
rect 5842 3442 5874 3474
rect 5910 3442 5942 3474
rect 5978 3442 6010 3474
rect 6046 3442 6078 3474
rect 6114 3442 6146 3474
rect 6182 3442 6214 3474
rect 6250 3442 6282 3474
rect 6318 3442 6350 3474
rect 6386 3442 6418 3474
rect 6454 3442 6486 3474
rect 6522 3442 6554 3474
rect 6590 3442 6622 3474
rect 6658 3442 6690 3474
rect 6726 3442 6758 3474
rect 6794 3442 6826 3474
rect 6862 3442 6894 3474
rect 6930 3442 6962 3474
rect 6998 3442 7030 3474
rect 7066 3442 7098 3474
rect 7134 3442 7166 3474
rect 7202 3442 7234 3474
rect 7270 3442 7302 3474
rect 7338 3442 7370 3474
rect 7406 3442 7438 3474
rect 7474 3442 7506 3474
rect 7542 3442 7574 3474
rect 7610 3442 7642 3474
rect 7678 3442 7710 3474
rect 7746 3442 7778 3474
rect 7814 3442 7846 3474
rect 7882 3442 7914 3474
rect 7950 3442 7982 3474
rect 8018 3442 8050 3474
rect 8086 3442 8118 3474
rect 8154 3442 8186 3474
rect 8222 3442 8254 3474
rect 8290 3442 8322 3474
rect 8358 3442 8390 3474
rect 8426 3442 8458 3474
rect 8494 3442 8526 3474
rect 8562 3442 8594 3474
rect 8630 3442 8662 3474
rect 8698 3442 8730 3474
rect 8766 3442 8798 3474
rect 8834 3442 8866 3474
rect 8902 3442 8934 3474
rect 8970 3442 9002 3474
rect 9038 3442 9070 3474
rect 9106 3442 9138 3474
rect 9174 3442 9206 3474
rect 9242 3442 9274 3474
rect 9310 3442 9342 3474
rect 9378 3442 9410 3474
rect 9446 3442 9478 3474
rect 9514 3442 9546 3474
rect 9582 3442 9614 3474
rect 9650 3442 9682 3474
rect 9718 3442 9750 3474
rect 9786 3442 9818 3474
rect 9854 3442 9886 3474
rect 9922 3442 9954 3474
rect 9990 3442 10022 3474
rect 10058 3442 10090 3474
rect 10126 3442 10158 3474
rect 10194 3442 10226 3474
rect 10262 3442 10294 3474
rect 10330 3442 10362 3474
rect 10398 3442 10430 3474
rect 10466 3442 10498 3474
rect 10534 3442 10566 3474
rect 10602 3442 10634 3474
rect 10670 3442 10702 3474
rect 10738 3442 10770 3474
rect 10806 3442 10838 3474
rect 10874 3442 10906 3474
rect 10942 3442 10974 3474
rect 11010 3442 11042 3474
rect 11078 3442 11110 3474
rect 11146 3442 11178 3474
rect 11214 3442 11246 3474
rect 11282 3442 11314 3474
rect 11350 3442 11382 3474
rect 11418 3442 11450 3474
rect 11486 3442 11518 3474
rect 11554 3442 11586 3474
rect 11622 3442 11654 3474
rect 11690 3442 11722 3474
rect 11758 3442 11790 3474
rect 11826 3442 11858 3474
rect 11894 3442 11926 3474
rect 11962 3442 11994 3474
rect 12030 3442 12062 3474
rect 12098 3442 12130 3474
rect 12166 3442 12198 3474
rect 12234 3442 12266 3474
rect 12302 3442 12334 3474
rect 12370 3442 12402 3474
rect 12438 3442 12470 3474
rect 12506 3442 12538 3474
rect 12574 3442 12606 3474
rect 12642 3442 12674 3474
rect 12710 3442 12742 3474
rect 12778 3442 12810 3474
rect 12846 3442 12878 3474
rect 12914 3442 12946 3474
rect 12982 3442 13014 3474
rect 13050 3442 13082 3474
rect 13118 3442 13150 3474
rect 13186 3442 13218 3474
rect 13254 3442 13286 3474
rect 13322 3442 13354 3474
rect 13390 3442 13422 3474
rect 13458 3442 13490 3474
rect 13526 3442 13558 3474
rect 13594 3442 13626 3474
rect 13662 3442 13694 3474
rect 13730 3442 13762 3474
rect 13798 3442 13830 3474
rect 13866 3442 13898 3474
rect 13934 3442 13966 3474
rect 14002 3442 14034 3474
rect 14070 3442 14102 3474
rect 14138 3442 14170 3474
rect 14206 3442 14238 3474
rect 14274 3442 14306 3474
rect 14342 3442 14374 3474
rect 14410 3442 14442 3474
rect 14478 3442 14510 3474
rect 14546 3442 14578 3474
rect 14614 3442 14646 3474
rect 14682 3442 14714 3474
rect 14750 3442 14782 3474
rect 14818 3442 14850 3474
rect 14886 3442 14918 3474
rect 14954 3442 14986 3474
rect 15022 3442 15054 3474
rect 15090 3442 15122 3474
rect 15158 3442 15190 3474
rect 15226 3442 15258 3474
rect 15294 3442 15326 3474
rect 15362 3442 15394 3474
rect 15430 3442 15462 3474
rect 15498 3442 15530 3474
rect 15566 3442 15598 3474
rect 378 3338 410 3370
rect 15590 3338 15622 3370
rect 378 3270 410 3302
rect 378 3202 410 3234
rect 378 3134 410 3166
rect 378 3066 410 3098
rect 378 2998 410 3030
rect 378 2930 410 2962
rect 378 2862 410 2894
rect 378 2794 410 2826
rect 378 2726 410 2758
rect 378 2658 410 2690
rect 378 2590 410 2622
rect 378 2522 410 2554
rect 378 2454 410 2486
rect 378 2386 410 2418
rect 378 2318 410 2350
rect 378 2250 410 2282
rect 378 2182 410 2214
rect 378 2114 410 2146
rect 378 2046 410 2078
rect 378 1978 410 2010
rect 15590 3270 15622 3302
rect 15590 3202 15622 3234
rect 15590 3134 15622 3166
rect 15590 3066 15622 3098
rect 15590 2998 15622 3030
rect 15590 2930 15622 2962
rect 15590 2862 15622 2894
rect 15590 2794 15622 2826
rect 15590 2726 15622 2758
rect 15590 2658 15622 2690
rect 15590 2590 15622 2622
rect 15590 2522 15622 2554
rect 15590 2454 15622 2486
rect 15590 2386 15622 2418
rect 15590 2318 15622 2350
rect 15590 2250 15622 2282
rect 15590 2182 15622 2214
rect 15590 2114 15622 2146
rect 15590 2046 15622 2078
rect 15590 1978 15622 2010
rect 378 1910 410 1942
rect 15590 1910 15622 1942
rect 378 1842 410 1874
rect 378 1774 410 1806
rect 378 1706 410 1738
rect 378 1638 410 1670
rect 378 1570 410 1602
rect 378 1502 410 1534
rect 378 1434 410 1466
rect 378 1366 410 1398
rect 378 1298 410 1330
rect 378 1230 410 1262
rect 378 1162 410 1194
rect 378 1094 410 1126
rect 378 1026 410 1058
rect 378 958 410 990
rect 378 890 410 922
rect 378 822 410 854
rect 378 754 410 786
rect 378 686 410 718
rect 378 618 410 650
rect 378 550 410 582
rect 15590 1842 15622 1874
rect 15590 1774 15622 1806
rect 15590 1706 15622 1738
rect 15590 1638 15622 1670
rect 15590 1570 15622 1602
rect 15590 1502 15622 1534
rect 15590 1434 15622 1466
rect 15590 1366 15622 1398
rect 15590 1298 15622 1330
rect 15590 1230 15622 1262
rect 15590 1162 15622 1194
rect 15590 1094 15622 1126
rect 15590 1026 15622 1058
rect 15590 958 15622 990
rect 15590 890 15622 922
rect 15590 822 15622 854
rect 15590 754 15622 786
rect 15590 686 15622 718
rect 15590 618 15622 650
rect 15590 550 15622 582
rect 378 482 410 514
rect 15590 482 15622 514
rect 402 378 434 410
rect 470 378 502 410
rect 538 378 570 410
rect 606 378 638 410
rect 674 378 706 410
rect 742 378 774 410
rect 810 378 842 410
rect 878 378 910 410
rect 946 378 978 410
rect 1014 378 1046 410
rect 1082 378 1114 410
rect 1150 378 1182 410
rect 1218 378 1250 410
rect 1286 378 1318 410
rect 1354 378 1386 410
rect 1422 378 1454 410
rect 1490 378 1522 410
rect 1558 378 1590 410
rect 1626 378 1658 410
rect 1694 378 1726 410
rect 1762 378 1794 410
rect 1830 378 1862 410
rect 1898 378 1930 410
rect 1966 378 1998 410
rect 2034 378 2066 410
rect 2102 378 2134 410
rect 2170 378 2202 410
rect 2238 378 2270 410
rect 2306 378 2338 410
rect 2374 378 2406 410
rect 2442 378 2474 410
rect 2510 378 2542 410
rect 2578 378 2610 410
rect 2646 378 2678 410
rect 2714 378 2746 410
rect 2782 378 2814 410
rect 2850 378 2882 410
rect 2918 378 2950 410
rect 2986 378 3018 410
rect 3054 378 3086 410
rect 3122 378 3154 410
rect 3190 378 3222 410
rect 3258 378 3290 410
rect 3326 378 3358 410
rect 3394 378 3426 410
rect 3462 378 3494 410
rect 3530 378 3562 410
rect 3598 378 3630 410
rect 3666 378 3698 410
rect 3734 378 3766 410
rect 3802 378 3834 410
rect 3870 378 3902 410
rect 3938 378 3970 410
rect 4006 378 4038 410
rect 4074 378 4106 410
rect 4142 378 4174 410
rect 4210 378 4242 410
rect 4278 378 4310 410
rect 4346 378 4378 410
rect 4414 378 4446 410
rect 4482 378 4514 410
rect 4550 378 4582 410
rect 4618 378 4650 410
rect 4686 378 4718 410
rect 4754 378 4786 410
rect 4822 378 4854 410
rect 4890 378 4922 410
rect 4958 378 4990 410
rect 5026 378 5058 410
rect 5094 378 5126 410
rect 5162 378 5194 410
rect 5230 378 5262 410
rect 5298 378 5330 410
rect 5366 378 5398 410
rect 5434 378 5466 410
rect 5502 378 5534 410
rect 5570 378 5602 410
rect 5638 378 5670 410
rect 5706 378 5738 410
rect 5774 378 5806 410
rect 5842 378 5874 410
rect 5910 378 5942 410
rect 5978 378 6010 410
rect 6046 378 6078 410
rect 6114 378 6146 410
rect 6182 378 6214 410
rect 6250 378 6282 410
rect 6318 378 6350 410
rect 6386 378 6418 410
rect 6454 378 6486 410
rect 6522 378 6554 410
rect 6590 378 6622 410
rect 6658 378 6690 410
rect 6726 378 6758 410
rect 6794 378 6826 410
rect 6862 378 6894 410
rect 6930 378 6962 410
rect 6998 378 7030 410
rect 7066 378 7098 410
rect 7134 378 7166 410
rect 7202 378 7234 410
rect 7270 378 7302 410
rect 7338 378 7370 410
rect 7406 378 7438 410
rect 7474 378 7506 410
rect 7542 378 7574 410
rect 7610 378 7642 410
rect 7678 378 7710 410
rect 7746 378 7778 410
rect 7814 378 7846 410
rect 7882 378 7914 410
rect 7950 378 7982 410
rect 8018 378 8050 410
rect 8086 378 8118 410
rect 8154 378 8186 410
rect 8222 378 8254 410
rect 8290 378 8322 410
rect 8358 378 8390 410
rect 8426 378 8458 410
rect 8494 378 8526 410
rect 8562 378 8594 410
rect 8630 378 8662 410
rect 8698 378 8730 410
rect 8766 378 8798 410
rect 8834 378 8866 410
rect 8902 378 8934 410
rect 8970 378 9002 410
rect 9038 378 9070 410
rect 9106 378 9138 410
rect 9174 378 9206 410
rect 9242 378 9274 410
rect 9310 378 9342 410
rect 9378 378 9410 410
rect 9446 378 9478 410
rect 9514 378 9546 410
rect 9582 378 9614 410
rect 9650 378 9682 410
rect 9718 378 9750 410
rect 9786 378 9818 410
rect 9854 378 9886 410
rect 9922 378 9954 410
rect 9990 378 10022 410
rect 10058 378 10090 410
rect 10126 378 10158 410
rect 10194 378 10226 410
rect 10262 378 10294 410
rect 10330 378 10362 410
rect 10398 378 10430 410
rect 10466 378 10498 410
rect 10534 378 10566 410
rect 10602 378 10634 410
rect 10670 378 10702 410
rect 10738 378 10770 410
rect 10806 378 10838 410
rect 10874 378 10906 410
rect 10942 378 10974 410
rect 11010 378 11042 410
rect 11078 378 11110 410
rect 11146 378 11178 410
rect 11214 378 11246 410
rect 11282 378 11314 410
rect 11350 378 11382 410
rect 11418 378 11450 410
rect 11486 378 11518 410
rect 11554 378 11586 410
rect 11622 378 11654 410
rect 11690 378 11722 410
rect 11758 378 11790 410
rect 11826 378 11858 410
rect 11894 378 11926 410
rect 11962 378 11994 410
rect 12030 378 12062 410
rect 12098 378 12130 410
rect 12166 378 12198 410
rect 12234 378 12266 410
rect 12302 378 12334 410
rect 12370 378 12402 410
rect 12438 378 12470 410
rect 12506 378 12538 410
rect 12574 378 12606 410
rect 12642 378 12674 410
rect 12710 378 12742 410
rect 12778 378 12810 410
rect 12846 378 12878 410
rect 12914 378 12946 410
rect 12982 378 13014 410
rect 13050 378 13082 410
rect 13118 378 13150 410
rect 13186 378 13218 410
rect 13254 378 13286 410
rect 13322 378 13354 410
rect 13390 378 13422 410
rect 13458 378 13490 410
rect 13526 378 13558 410
rect 13594 378 13626 410
rect 13662 378 13694 410
rect 13730 378 13762 410
rect 13798 378 13830 410
rect 13866 378 13898 410
rect 13934 378 13966 410
rect 14002 378 14034 410
rect 14070 378 14102 410
rect 14138 378 14170 410
rect 14206 378 14238 410
rect 14274 378 14306 410
rect 14342 378 14374 410
rect 14410 378 14442 410
rect 14478 378 14510 410
rect 14546 378 14578 410
rect 14614 378 14646 410
rect 14682 378 14714 410
rect 14750 378 14782 410
rect 14818 378 14850 410
rect 14886 378 14918 410
rect 14954 378 14986 410
rect 15022 378 15054 410
rect 15090 378 15122 410
rect 15158 378 15190 410
rect 15226 378 15258 410
rect 15294 378 15326 410
rect 15362 378 15394 410
rect 15430 378 15462 410
rect 15498 378 15530 410
rect 15566 378 15598 410
<< poly >>
rect 5799 3362 5919 3376
rect 5799 3330 5843 3362
rect 5875 3330 5919 3362
rect 5799 3302 5919 3330
rect 6155 3362 6275 3376
rect 6155 3330 6199 3362
rect 6231 3330 6275 3362
rect 6155 3302 6275 3330
rect 6403 3362 6523 3376
rect 6403 3330 6447 3362
rect 6479 3330 6523 3362
rect 6403 3302 6523 3330
rect 6759 3362 6879 3376
rect 6759 3330 6803 3362
rect 6835 3330 6879 3362
rect 6759 3302 6879 3330
rect 7007 3362 7127 3376
rect 7007 3330 7051 3362
rect 7083 3330 7127 3362
rect 7007 3302 7127 3330
rect 7363 3362 7483 3376
rect 7363 3330 7407 3362
rect 7439 3330 7483 3362
rect 7363 3302 7483 3330
rect 7611 3362 7731 3376
rect 7611 3330 7655 3362
rect 7687 3330 7731 3362
rect 7611 3302 7731 3330
rect 7967 3362 8087 3376
rect 7967 3330 8011 3362
rect 8043 3330 8087 3362
rect 7967 3302 8087 3330
rect 8215 3362 8335 3376
rect 8215 3330 8259 3362
rect 8291 3330 8335 3362
rect 8215 3302 8335 3330
rect 8571 3362 8691 3376
rect 8571 3330 8615 3362
rect 8647 3330 8691 3362
rect 8571 3302 8691 3330
rect 8819 3362 8939 3376
rect 8819 3330 8863 3362
rect 8895 3330 8939 3362
rect 8819 3302 8939 3330
rect 9175 3362 9295 3376
rect 9175 3330 9219 3362
rect 9251 3330 9295 3362
rect 9175 3302 9295 3330
rect 9423 3362 9543 3376
rect 9423 3330 9467 3362
rect 9499 3330 9543 3362
rect 9423 3302 9543 3330
rect 9779 3362 9899 3376
rect 9779 3330 9823 3362
rect 9855 3330 9899 3362
rect 9779 3302 9899 3330
rect 10027 3362 10147 3376
rect 10027 3330 10071 3362
rect 10103 3330 10147 3362
rect 10027 3302 10147 3330
rect 5799 1942 5919 1970
rect 5799 1910 5843 1942
rect 5875 1910 5919 1942
rect 5799 1882 5919 1910
rect 6155 1942 6275 1970
rect 6155 1910 6199 1942
rect 6231 1910 6275 1942
rect 6155 1882 6275 1910
rect 6403 1942 6523 1970
rect 6403 1910 6447 1942
rect 6479 1910 6523 1942
rect 6403 1882 6523 1910
rect 6759 1942 6879 1970
rect 6759 1910 6803 1942
rect 6835 1910 6879 1942
rect 6759 1882 6879 1910
rect 7007 1942 7127 1970
rect 7007 1910 7051 1942
rect 7083 1910 7127 1942
rect 7007 1882 7127 1910
rect 7363 1942 7483 1970
rect 7363 1910 7407 1942
rect 7439 1910 7483 1942
rect 7363 1882 7483 1910
rect 7611 1942 7731 1970
rect 7611 1910 7655 1942
rect 7687 1910 7731 1942
rect 7611 1882 7731 1910
rect 7967 1942 8087 1970
rect 7967 1910 8011 1942
rect 8043 1910 8087 1942
rect 7967 1882 8087 1910
rect 8215 1942 8335 1970
rect 8215 1910 8259 1942
rect 8291 1910 8335 1942
rect 8215 1882 8335 1910
rect 8571 1942 8691 1970
rect 8571 1910 8615 1942
rect 8647 1910 8691 1942
rect 8571 1882 8691 1910
rect 8819 1942 8939 1970
rect 8819 1910 8863 1942
rect 8895 1910 8939 1942
rect 8819 1882 8939 1910
rect 9175 1942 9295 1970
rect 9175 1910 9219 1942
rect 9251 1910 9295 1942
rect 9175 1882 9295 1910
rect 9423 1942 9543 1970
rect 9423 1910 9467 1942
rect 9499 1910 9543 1942
rect 9423 1882 9543 1910
rect 9779 1942 9899 1970
rect 9779 1910 9823 1942
rect 9855 1910 9899 1942
rect 9779 1882 9899 1910
rect 10027 1942 10147 1970
rect 10027 1910 10071 1942
rect 10103 1910 10147 1942
rect 10027 1882 10147 1910
rect 5799 522 5919 550
rect 5799 490 5843 522
rect 5875 490 5919 522
rect 5799 476 5919 490
rect 6155 522 6275 550
rect 6155 490 6199 522
rect 6231 490 6275 522
rect 6155 476 6275 490
rect 6403 522 6523 550
rect 6403 490 6447 522
rect 6479 490 6523 522
rect 6403 476 6523 490
rect 6759 522 6879 550
rect 6759 490 6803 522
rect 6835 490 6879 522
rect 6759 476 6879 490
rect 7007 522 7127 550
rect 7007 490 7051 522
rect 7083 490 7127 522
rect 7007 476 7127 490
rect 7363 522 7483 550
rect 7363 490 7407 522
rect 7439 490 7483 522
rect 7363 476 7483 490
rect 7611 522 7731 550
rect 7611 490 7655 522
rect 7687 490 7731 522
rect 7611 476 7731 490
rect 7967 522 8087 550
rect 7967 490 8011 522
rect 8043 490 8087 522
rect 7967 476 8087 490
rect 8215 522 8335 550
rect 8215 490 8259 522
rect 8291 490 8335 522
rect 8215 476 8335 490
rect 8571 522 8691 550
rect 8571 490 8615 522
rect 8647 490 8691 522
rect 8571 476 8691 490
rect 8819 522 8939 550
rect 8819 490 8863 522
rect 8895 490 8939 522
rect 8819 476 8939 490
rect 9175 522 9295 550
rect 9175 490 9219 522
rect 9251 490 9295 522
rect 9175 476 9295 490
rect 9423 522 9543 550
rect 9423 490 9467 522
rect 9499 490 9543 522
rect 9423 476 9543 490
rect 9779 522 9899 550
rect 9779 490 9823 522
rect 9855 490 9899 522
rect 9779 476 9899 490
rect 10027 522 10147 550
rect 10027 490 10071 522
rect 10103 490 10147 522
rect 10027 476 10147 490
<< polycont >>
rect 5843 3330 5875 3362
rect 6199 3330 6231 3362
rect 6447 3330 6479 3362
rect 6803 3330 6835 3362
rect 7051 3330 7083 3362
rect 7407 3330 7439 3362
rect 7655 3330 7687 3362
rect 8011 3330 8043 3362
rect 8259 3330 8291 3362
rect 8615 3330 8647 3362
rect 8863 3330 8895 3362
rect 9219 3330 9251 3362
rect 9467 3330 9499 3362
rect 9823 3330 9855 3362
rect 10071 3330 10103 3362
rect 5843 1910 5875 1942
rect 6199 1910 6231 1942
rect 6447 1910 6479 1942
rect 6803 1910 6835 1942
rect 7051 1910 7083 1942
rect 7407 1910 7439 1942
rect 7655 1910 7687 1942
rect 8011 1910 8043 1942
rect 8259 1910 8291 1942
rect 8615 1910 8647 1942
rect 8863 1910 8895 1942
rect 9219 1910 9251 1942
rect 9467 1910 9499 1942
rect 9823 1910 9855 1942
rect 10071 1910 10103 1942
rect 5843 490 5875 522
rect 6199 490 6231 522
rect 6447 490 6479 522
rect 6803 490 6835 522
rect 7051 490 7083 522
rect 7407 490 7439 522
rect 7655 490 7687 522
rect 8011 490 8043 522
rect 8259 490 8291 522
rect 8615 490 8647 522
rect 8863 490 8895 522
rect 9219 490 9251 522
rect 9467 490 9499 522
rect 9823 490 9855 522
rect 10071 490 10103 522
<< pdiode >>
rect 2992 3270 3148 3298
rect 2992 3238 3020 3270
rect 3052 3238 3088 3270
rect 3120 3238 3148 3270
rect 2992 3202 3148 3238
rect 2992 3170 3020 3202
rect 3052 3170 3088 3202
rect 3120 3170 3148 3202
rect 2992 3142 3148 3170
<< pdiodecont >>
rect 3020 3238 3052 3270
rect 3088 3238 3120 3270
rect 3020 3170 3052 3202
rect 3088 3170 3120 3202
<< metal1 >>
rect 0 3834 16000 3852
rect 0 3802 28 3834
rect 60 3802 96 3834
rect 128 3802 164 3834
rect 196 3802 232 3834
rect 264 3802 300 3834
rect 332 3802 368 3834
rect 400 3802 436 3834
rect 468 3802 504 3834
rect 536 3802 572 3834
rect 604 3802 640 3834
rect 672 3802 708 3834
rect 740 3802 776 3834
rect 808 3802 844 3834
rect 876 3802 912 3834
rect 944 3802 980 3834
rect 1012 3802 1048 3834
rect 1080 3802 1116 3834
rect 1148 3802 1184 3834
rect 1216 3802 1252 3834
rect 1284 3802 1320 3834
rect 1352 3802 1388 3834
rect 1420 3802 1456 3834
rect 1488 3802 1524 3834
rect 1556 3802 1592 3834
rect 1624 3802 1660 3834
rect 1692 3802 1728 3834
rect 1760 3802 1796 3834
rect 1828 3802 1864 3834
rect 1896 3802 1932 3834
rect 1964 3802 2000 3834
rect 2032 3802 2068 3834
rect 2100 3802 2136 3834
rect 2168 3802 2204 3834
rect 2236 3802 2272 3834
rect 2304 3802 2340 3834
rect 2372 3802 2408 3834
rect 2440 3802 2476 3834
rect 2508 3802 2544 3834
rect 2576 3802 2612 3834
rect 2644 3802 2680 3834
rect 2712 3802 2748 3834
rect 2780 3802 2816 3834
rect 2848 3802 2884 3834
rect 2916 3802 2952 3834
rect 2984 3802 3020 3834
rect 3052 3802 3088 3834
rect 3120 3802 3156 3834
rect 3188 3802 3224 3834
rect 3256 3802 3292 3834
rect 3324 3802 3360 3834
rect 3392 3802 3428 3834
rect 3460 3802 3496 3834
rect 3528 3802 3564 3834
rect 3596 3802 3632 3834
rect 3664 3802 3700 3834
rect 3732 3802 3768 3834
rect 3800 3802 3836 3834
rect 3868 3802 3904 3834
rect 3936 3802 3972 3834
rect 4004 3802 4040 3834
rect 4072 3802 4108 3834
rect 4140 3802 4176 3834
rect 4208 3802 4244 3834
rect 4276 3802 4312 3834
rect 4344 3802 4380 3834
rect 4412 3802 4448 3834
rect 4480 3802 4516 3834
rect 4548 3802 4584 3834
rect 4616 3802 4652 3834
rect 4684 3802 4720 3834
rect 4752 3802 4788 3834
rect 4820 3802 4856 3834
rect 4888 3802 4924 3834
rect 4956 3802 4992 3834
rect 5024 3802 5060 3834
rect 5092 3802 5128 3834
rect 5160 3802 5196 3834
rect 5228 3802 5264 3834
rect 5296 3802 5332 3834
rect 5364 3802 5400 3834
rect 5432 3802 5468 3834
rect 5500 3802 5536 3834
rect 5568 3802 5604 3834
rect 5636 3802 5672 3834
rect 5704 3802 5740 3834
rect 5772 3802 5808 3834
rect 5840 3802 5876 3834
rect 5908 3802 5944 3834
rect 5976 3802 6012 3834
rect 6044 3802 6080 3834
rect 6112 3802 6148 3834
rect 6180 3802 6216 3834
rect 6248 3802 6284 3834
rect 6316 3802 6352 3834
rect 6384 3802 6420 3834
rect 6452 3802 6488 3834
rect 6520 3802 6556 3834
rect 6588 3802 6624 3834
rect 6656 3802 6692 3834
rect 6724 3802 6760 3834
rect 6792 3802 6828 3834
rect 6860 3802 6896 3834
rect 6928 3802 6964 3834
rect 6996 3802 7032 3834
rect 7064 3802 7100 3834
rect 7132 3802 7168 3834
rect 7200 3802 7236 3834
rect 7268 3802 7304 3834
rect 7336 3802 7372 3834
rect 7404 3802 7440 3834
rect 7472 3802 7508 3834
rect 7540 3802 7576 3834
rect 7608 3802 7644 3834
rect 7676 3802 7712 3834
rect 7744 3802 7780 3834
rect 7812 3802 7848 3834
rect 7880 3802 7916 3834
rect 7948 3802 7984 3834
rect 8016 3802 8052 3834
rect 8084 3802 8120 3834
rect 8152 3802 8188 3834
rect 8220 3802 8256 3834
rect 8288 3802 8324 3834
rect 8356 3802 8392 3834
rect 8424 3802 8460 3834
rect 8492 3802 8528 3834
rect 8560 3802 8596 3834
rect 8628 3802 8664 3834
rect 8696 3802 8732 3834
rect 8764 3802 8800 3834
rect 8832 3802 8868 3834
rect 8900 3802 8936 3834
rect 8968 3802 9004 3834
rect 9036 3802 9072 3834
rect 9104 3802 9140 3834
rect 9172 3802 9208 3834
rect 9240 3802 9276 3834
rect 9308 3802 9344 3834
rect 9376 3802 9412 3834
rect 9444 3802 9480 3834
rect 9512 3802 9548 3834
rect 9580 3802 9616 3834
rect 9648 3802 9684 3834
rect 9716 3802 9752 3834
rect 9784 3802 9820 3834
rect 9852 3802 9888 3834
rect 9920 3802 9956 3834
rect 9988 3802 10024 3834
rect 10056 3802 10092 3834
rect 10124 3802 10160 3834
rect 10192 3802 10228 3834
rect 10260 3802 10296 3834
rect 10328 3802 10364 3834
rect 10396 3802 10432 3834
rect 10464 3802 10500 3834
rect 10532 3802 10568 3834
rect 10600 3802 10636 3834
rect 10668 3802 10704 3834
rect 10736 3802 10772 3834
rect 10804 3802 10840 3834
rect 10872 3802 10908 3834
rect 10940 3802 10976 3834
rect 11008 3802 11044 3834
rect 11076 3802 11112 3834
rect 11144 3802 11180 3834
rect 11212 3802 11248 3834
rect 11280 3802 11316 3834
rect 11348 3802 11384 3834
rect 11416 3802 11452 3834
rect 11484 3802 11520 3834
rect 11552 3802 11588 3834
rect 11620 3802 11656 3834
rect 11688 3802 11724 3834
rect 11756 3802 11792 3834
rect 11824 3802 11860 3834
rect 11892 3802 11928 3834
rect 11960 3802 11996 3834
rect 12028 3802 12064 3834
rect 12096 3802 12132 3834
rect 12164 3802 12200 3834
rect 12232 3802 12268 3834
rect 12300 3802 12336 3834
rect 12368 3802 12404 3834
rect 12436 3802 12472 3834
rect 12504 3802 12540 3834
rect 12572 3802 12608 3834
rect 12640 3802 12676 3834
rect 12708 3802 12744 3834
rect 12776 3802 12812 3834
rect 12844 3802 12880 3834
rect 12912 3802 12948 3834
rect 12980 3802 13016 3834
rect 13048 3802 13084 3834
rect 13116 3802 13152 3834
rect 13184 3802 13220 3834
rect 13252 3802 13288 3834
rect 13320 3802 13356 3834
rect 13388 3802 13424 3834
rect 13456 3802 13492 3834
rect 13524 3802 13560 3834
rect 13592 3802 13628 3834
rect 13660 3802 13696 3834
rect 13728 3802 13764 3834
rect 13796 3802 13832 3834
rect 13864 3802 13900 3834
rect 13932 3802 13968 3834
rect 14000 3802 14036 3834
rect 14068 3802 14104 3834
rect 14136 3802 14172 3834
rect 14204 3802 14240 3834
rect 14272 3802 14308 3834
rect 14340 3802 14376 3834
rect 14408 3802 14444 3834
rect 14476 3802 14512 3834
rect 14544 3802 14580 3834
rect 14612 3802 14648 3834
rect 14680 3802 14716 3834
rect 14748 3802 14784 3834
rect 14816 3802 14852 3834
rect 14884 3802 14920 3834
rect 14952 3802 14988 3834
rect 15020 3802 15056 3834
rect 15088 3802 15124 3834
rect 15156 3802 15192 3834
rect 15224 3802 15260 3834
rect 15292 3802 15328 3834
rect 15360 3802 15396 3834
rect 15428 3802 15464 3834
rect 15496 3802 15532 3834
rect 15564 3802 15600 3834
rect 15632 3802 15668 3834
rect 15700 3802 15736 3834
rect 15768 3802 15804 3834
rect 15836 3802 15872 3834
rect 15904 3802 15940 3834
rect 15972 3802 16000 3834
rect 0 3784 16000 3802
rect 0 3744 68 3784
rect 0 3712 18 3744
rect 50 3712 68 3744
rect 0 3676 68 3712
rect 0 3644 18 3676
rect 50 3644 68 3676
rect 0 3608 68 3644
rect 0 3576 18 3608
rect 50 3576 68 3608
rect 0 3540 68 3576
rect 0 3508 18 3540
rect 50 3508 68 3540
rect 0 3472 68 3508
rect 15932 3744 16000 3784
rect 15932 3712 15950 3744
rect 15982 3712 16000 3744
rect 15932 3676 16000 3712
rect 15932 3644 15950 3676
rect 15982 3644 16000 3676
rect 15932 3608 16000 3644
rect 15932 3576 15950 3608
rect 15982 3576 16000 3608
rect 15932 3540 16000 3576
rect 15932 3508 15950 3540
rect 15982 3508 16000 3540
rect 0 3440 18 3472
rect 50 3440 68 3472
rect 0 3404 68 3440
rect 0 3372 18 3404
rect 50 3372 68 3404
rect 0 3336 68 3372
rect 0 3304 18 3336
rect 50 3304 68 3336
rect 0 3268 68 3304
rect 0 3236 18 3268
rect 50 3236 68 3268
rect 0 3200 68 3236
rect 0 3168 18 3200
rect 50 3168 68 3200
rect 0 3132 68 3168
rect 0 3100 18 3132
rect 50 3100 68 3132
rect 0 3064 68 3100
rect 0 3032 18 3064
rect 50 3032 68 3064
rect 0 2996 68 3032
rect 0 2964 18 2996
rect 50 2964 68 2996
rect 0 2928 68 2964
rect 0 2896 18 2928
rect 50 2896 68 2928
rect 0 2860 68 2896
rect 0 2828 18 2860
rect 50 2828 68 2860
rect 0 2792 68 2828
rect 0 2760 18 2792
rect 50 2760 68 2792
rect 0 2724 68 2760
rect 0 2692 18 2724
rect 50 2692 68 2724
rect 0 2656 68 2692
rect 0 2624 18 2656
rect 50 2624 68 2656
rect 0 2588 68 2624
rect 0 2556 18 2588
rect 50 2556 68 2588
rect 0 2520 68 2556
rect 0 2488 18 2520
rect 50 2488 68 2520
rect 0 2452 68 2488
rect 0 2420 18 2452
rect 50 2420 68 2452
rect 0 2384 68 2420
rect 0 2352 18 2384
rect 50 2352 68 2384
rect 0 2316 68 2352
rect 0 2284 18 2316
rect 50 2284 68 2316
rect 0 2248 68 2284
rect 0 2216 18 2248
rect 50 2216 68 2248
rect 0 2180 68 2216
rect 0 2148 18 2180
rect 50 2148 68 2180
rect 0 2112 68 2148
rect 0 2080 18 2112
rect 50 2080 68 2112
rect 0 2044 68 2080
rect 0 2012 18 2044
rect 50 2012 68 2044
rect 0 1976 68 2012
rect 0 1944 18 1976
rect 50 1944 68 1976
rect 0 1908 68 1944
rect 0 1876 18 1908
rect 50 1876 68 1908
rect 0 1840 68 1876
rect 0 1808 18 1840
rect 50 1808 68 1840
rect 0 1772 68 1808
rect 0 1740 18 1772
rect 50 1740 68 1772
rect 0 1704 68 1740
rect 0 1672 18 1704
rect 50 1672 68 1704
rect 0 1636 68 1672
rect 0 1604 18 1636
rect 50 1604 68 1636
rect 0 1568 68 1604
rect 0 1536 18 1568
rect 50 1536 68 1568
rect 0 1500 68 1536
rect 0 1468 18 1500
rect 50 1468 68 1500
rect 0 1432 68 1468
rect 0 1400 18 1432
rect 50 1400 68 1432
rect 0 1364 68 1400
rect 0 1332 18 1364
rect 50 1332 68 1364
rect 0 1296 68 1332
rect 0 1264 18 1296
rect 50 1264 68 1296
rect 0 1228 68 1264
rect 0 1196 18 1228
rect 50 1196 68 1228
rect 0 1160 68 1196
rect 0 1128 18 1160
rect 50 1128 68 1160
rect 0 1092 68 1128
rect 0 1060 18 1092
rect 50 1060 68 1092
rect 0 1024 68 1060
rect 0 992 18 1024
rect 50 992 68 1024
rect 0 956 68 992
rect 0 924 18 956
rect 50 924 68 956
rect 0 888 68 924
rect 0 856 18 888
rect 50 856 68 888
rect 0 820 68 856
rect 0 788 18 820
rect 50 788 68 820
rect 0 752 68 788
rect 0 720 18 752
rect 50 720 68 752
rect 0 684 68 720
rect 0 652 18 684
rect 50 652 68 684
rect 0 616 68 652
rect 0 584 18 616
rect 50 584 68 616
rect 0 548 68 584
rect 0 516 18 548
rect 50 516 68 548
rect 0 480 68 516
rect 0 448 18 480
rect 50 448 68 480
rect 0 412 68 448
rect 0 380 18 412
rect 50 380 68 412
rect 0 344 68 380
rect 360 3478 15640 3492
rect 360 3474 5715 3478
rect 5755 3474 6319 3478
rect 6359 3474 6923 3478
rect 6963 3474 7527 3478
rect 7567 3474 8131 3478
rect 8171 3474 8735 3478
rect 8775 3474 9339 3478
rect 9379 3474 9943 3478
rect 9983 3474 15640 3478
rect 360 3442 402 3474
rect 434 3442 470 3474
rect 502 3442 538 3474
rect 570 3442 606 3474
rect 638 3442 674 3474
rect 706 3442 742 3474
rect 774 3442 810 3474
rect 842 3442 878 3474
rect 910 3442 946 3474
rect 978 3442 1014 3474
rect 1046 3442 1082 3474
rect 1114 3442 1150 3474
rect 1182 3442 1218 3474
rect 1250 3442 1286 3474
rect 1318 3442 1354 3474
rect 1386 3442 1422 3474
rect 1454 3442 1490 3474
rect 1522 3442 1558 3474
rect 1590 3442 1626 3474
rect 1658 3442 1694 3474
rect 1726 3442 1762 3474
rect 1794 3442 1830 3474
rect 1862 3442 1898 3474
rect 1930 3442 1966 3474
rect 1998 3442 2034 3474
rect 2066 3442 2102 3474
rect 2134 3442 2170 3474
rect 2202 3442 2238 3474
rect 2270 3442 2306 3474
rect 2338 3442 2374 3474
rect 2406 3442 2442 3474
rect 2474 3442 2510 3474
rect 2542 3442 2578 3474
rect 2610 3442 2646 3474
rect 2678 3442 2714 3474
rect 2746 3442 2782 3474
rect 2814 3442 2850 3474
rect 2882 3442 2918 3474
rect 2950 3442 2986 3474
rect 3018 3442 3054 3474
rect 3086 3442 3122 3474
rect 3154 3442 3190 3474
rect 3222 3442 3258 3474
rect 3290 3442 3326 3474
rect 3358 3442 3394 3474
rect 3426 3442 3462 3474
rect 3494 3442 3530 3474
rect 3562 3442 3598 3474
rect 3630 3442 3666 3474
rect 3698 3442 3734 3474
rect 3766 3442 3802 3474
rect 3834 3442 3870 3474
rect 3902 3442 3938 3474
rect 3970 3442 4006 3474
rect 4038 3442 4074 3474
rect 4106 3442 4142 3474
rect 4174 3442 4210 3474
rect 4242 3442 4278 3474
rect 4310 3442 4346 3474
rect 4378 3442 4414 3474
rect 4446 3442 4482 3474
rect 4514 3442 4550 3474
rect 4582 3442 4618 3474
rect 4650 3442 4686 3474
rect 4718 3442 4754 3474
rect 4786 3442 4822 3474
rect 4854 3442 4890 3474
rect 4922 3442 4958 3474
rect 4990 3442 5026 3474
rect 5058 3442 5094 3474
rect 5126 3442 5162 3474
rect 5194 3442 5230 3474
rect 5262 3442 5298 3474
rect 5330 3442 5366 3474
rect 5398 3442 5434 3474
rect 5466 3442 5502 3474
rect 5534 3442 5570 3474
rect 5602 3442 5638 3474
rect 5670 3442 5706 3474
rect 5755 3442 5774 3474
rect 5806 3442 5842 3474
rect 5874 3442 5910 3474
rect 5942 3442 5978 3474
rect 6010 3442 6046 3474
rect 6078 3442 6114 3474
rect 6146 3442 6182 3474
rect 6214 3442 6250 3474
rect 6282 3442 6318 3474
rect 6359 3442 6386 3474
rect 6418 3442 6454 3474
rect 6486 3442 6522 3474
rect 6554 3442 6590 3474
rect 6622 3442 6658 3474
rect 6690 3442 6726 3474
rect 6758 3442 6794 3474
rect 6826 3442 6862 3474
rect 6894 3442 6923 3474
rect 6963 3442 6998 3474
rect 7030 3442 7066 3474
rect 7098 3442 7134 3474
rect 7166 3442 7202 3474
rect 7234 3442 7270 3474
rect 7302 3442 7338 3474
rect 7370 3442 7406 3474
rect 7438 3442 7474 3474
rect 7506 3442 7527 3474
rect 7574 3442 7610 3474
rect 7642 3442 7678 3474
rect 7710 3442 7746 3474
rect 7778 3442 7814 3474
rect 7846 3442 7882 3474
rect 7914 3442 7950 3474
rect 7982 3442 8018 3474
rect 8050 3442 8086 3474
rect 8118 3442 8131 3474
rect 8186 3442 8222 3474
rect 8254 3442 8290 3474
rect 8322 3442 8358 3474
rect 8390 3442 8426 3474
rect 8458 3442 8494 3474
rect 8526 3442 8562 3474
rect 8594 3442 8630 3474
rect 8662 3442 8698 3474
rect 8730 3442 8735 3474
rect 8798 3442 8834 3474
rect 8866 3442 8902 3474
rect 8934 3442 8970 3474
rect 9002 3442 9038 3474
rect 9070 3442 9106 3474
rect 9138 3442 9174 3474
rect 9206 3442 9242 3474
rect 9274 3442 9310 3474
rect 9410 3442 9446 3474
rect 9478 3442 9514 3474
rect 9546 3442 9582 3474
rect 9614 3442 9650 3474
rect 9682 3442 9718 3474
rect 9750 3442 9786 3474
rect 9818 3442 9854 3474
rect 9886 3442 9922 3474
rect 9983 3442 9990 3474
rect 10022 3442 10058 3474
rect 10090 3442 10126 3474
rect 10158 3442 10194 3474
rect 10226 3442 10262 3474
rect 10294 3442 10330 3474
rect 10362 3442 10398 3474
rect 10430 3442 10466 3474
rect 10498 3442 10534 3474
rect 10566 3442 10602 3474
rect 10634 3442 10670 3474
rect 10702 3442 10738 3474
rect 10770 3442 10806 3474
rect 10838 3442 10874 3474
rect 10906 3442 10942 3474
rect 10974 3442 11010 3474
rect 11042 3442 11078 3474
rect 11110 3442 11146 3474
rect 11178 3442 11214 3474
rect 11246 3442 11282 3474
rect 11314 3442 11350 3474
rect 11382 3442 11418 3474
rect 11450 3442 11486 3474
rect 11518 3442 11554 3474
rect 11586 3442 11622 3474
rect 11654 3442 11690 3474
rect 11722 3442 11758 3474
rect 11790 3442 11826 3474
rect 11858 3442 11894 3474
rect 11926 3442 11962 3474
rect 11994 3442 12030 3474
rect 12062 3442 12098 3474
rect 12130 3442 12166 3474
rect 12198 3442 12234 3474
rect 12266 3442 12302 3474
rect 12334 3442 12370 3474
rect 12402 3442 12438 3474
rect 12470 3442 12506 3474
rect 12538 3442 12574 3474
rect 12606 3442 12642 3474
rect 12674 3442 12710 3474
rect 12742 3442 12778 3474
rect 12810 3442 12846 3474
rect 12878 3442 12914 3474
rect 12946 3442 12982 3474
rect 13014 3442 13050 3474
rect 13082 3442 13118 3474
rect 13150 3442 13186 3474
rect 13218 3442 13254 3474
rect 13286 3442 13322 3474
rect 13354 3442 13390 3474
rect 13422 3442 13458 3474
rect 13490 3442 13526 3474
rect 13558 3442 13594 3474
rect 13626 3442 13662 3474
rect 13694 3442 13730 3474
rect 13762 3442 13798 3474
rect 13830 3442 13866 3474
rect 13898 3442 13934 3474
rect 13966 3442 14002 3474
rect 14034 3442 14070 3474
rect 14102 3442 14138 3474
rect 14170 3442 14206 3474
rect 14238 3442 14274 3474
rect 14306 3442 14342 3474
rect 14374 3442 14410 3474
rect 14442 3442 14478 3474
rect 14510 3442 14546 3474
rect 14578 3442 14614 3474
rect 14646 3442 14682 3474
rect 14714 3442 14750 3474
rect 14782 3442 14818 3474
rect 14850 3442 14886 3474
rect 14918 3442 14954 3474
rect 14986 3442 15022 3474
rect 15054 3442 15090 3474
rect 15122 3442 15158 3474
rect 15190 3442 15226 3474
rect 15258 3442 15294 3474
rect 15326 3442 15362 3474
rect 15394 3442 15430 3474
rect 15462 3442 15498 3474
rect 15530 3442 15566 3474
rect 15598 3442 15640 3474
rect 360 3438 5715 3442
rect 5755 3438 6319 3442
rect 6359 3438 6923 3442
rect 6963 3438 7527 3442
rect 7567 3438 8131 3442
rect 8171 3438 8735 3442
rect 8775 3438 9339 3442
rect 9379 3438 9943 3442
rect 9983 3438 15640 3442
rect 360 3424 15640 3438
rect 360 3370 428 3424
rect 360 3338 378 3370
rect 410 3338 428 3370
rect 360 3302 428 3338
rect 360 3270 378 3302
rect 410 3270 428 3302
rect 3045 3362 10103 3378
rect 3045 3359 5843 3362
rect 3045 3319 3046 3359
rect 3086 3346 5843 3359
rect 3086 3319 3087 3346
rect 3045 3270 3087 3319
rect 5875 3346 6199 3362
rect 360 3234 428 3270
rect 360 3202 378 3234
rect 410 3202 428 3234
rect 360 3166 428 3202
rect 3010 3263 3130 3270
rect 3010 3223 3046 3263
rect 3086 3223 3130 3263
rect 3010 3170 3130 3223
rect 5714 3264 5756 3280
rect 5714 3232 5719 3264
rect 5751 3232 5756 3264
rect 5714 3230 5756 3232
rect 360 3134 378 3166
rect 410 3134 428 3166
rect 360 3098 428 3134
rect 360 3066 378 3098
rect 410 3066 428 3098
rect 360 3030 428 3066
rect 360 2998 378 3030
rect 410 2998 428 3030
rect 360 2962 428 2998
rect 360 2930 378 2962
rect 410 2930 428 2962
rect 360 2894 428 2930
rect 360 2862 378 2894
rect 410 2862 428 2894
rect 360 2826 428 2862
rect 360 2794 378 2826
rect 410 2794 428 2826
rect 360 2758 428 2794
rect 360 2726 378 2758
rect 410 2726 428 2758
rect 360 2690 428 2726
rect 360 2658 378 2690
rect 410 2658 428 2690
rect 360 2622 428 2658
rect 360 2590 378 2622
rect 410 2590 428 2622
rect 360 2554 428 2590
rect 360 2522 378 2554
rect 410 2522 428 2554
rect 360 2486 428 2522
rect 360 2454 378 2486
rect 410 2454 428 2486
rect 360 2418 428 2454
rect 360 2386 378 2418
rect 410 2386 428 2418
rect 360 2350 428 2386
rect 360 2318 378 2350
rect 410 2318 428 2350
rect 360 2282 428 2318
rect 360 2250 378 2282
rect 410 2250 428 2282
rect 360 2214 428 2250
rect 360 2182 378 2214
rect 410 2182 428 2214
rect 360 2146 428 2182
rect 360 2114 378 2146
rect 410 2114 428 2146
rect 360 2078 428 2114
rect 360 2046 378 2078
rect 410 2046 428 2078
rect 360 2010 428 2046
rect 360 1978 378 2010
rect 410 1978 428 2010
rect 5714 2042 5715 3230
rect 5755 2042 5756 3230
rect 5714 2040 5756 2042
rect 5714 2008 5719 2040
rect 5751 2008 5756 2040
rect 5714 1992 5756 2008
rect 360 1942 428 1978
rect 360 1910 378 1942
rect 410 1910 428 1942
rect 360 1874 428 1910
rect 360 1842 378 1874
rect 410 1842 428 1874
rect 5843 1942 5875 3330
rect 6231 3346 6447 3362
rect 5975 3264 6099 3280
rect 5975 3232 6021 3264
rect 6053 3232 6099 3264
rect 5975 3230 6099 3232
rect 5975 2042 5976 3230
rect 6098 2042 6099 3230
rect 5975 2040 6099 2042
rect 5975 2008 6021 2040
rect 6053 2008 6099 2040
rect 5975 1992 6099 2008
rect 360 1806 428 1842
rect 360 1774 378 1806
rect 410 1774 428 1806
rect 360 1738 428 1774
rect 360 1706 378 1738
rect 410 1706 428 1738
rect 360 1670 428 1706
rect 360 1638 378 1670
rect 410 1638 428 1670
rect 360 1602 428 1638
rect 360 1570 378 1602
rect 410 1570 428 1602
rect 360 1534 428 1570
rect 360 1502 378 1534
rect 410 1502 428 1534
rect 360 1466 428 1502
rect 360 1434 378 1466
rect 410 1434 428 1466
rect 360 1398 428 1434
rect 360 1366 378 1398
rect 410 1366 428 1398
rect 360 1330 428 1366
rect 360 1298 378 1330
rect 410 1298 428 1330
rect 360 1262 428 1298
rect 360 1230 378 1262
rect 410 1230 428 1262
rect 360 1194 428 1230
rect 360 1162 378 1194
rect 410 1162 428 1194
rect 360 1126 428 1162
rect 360 1094 378 1126
rect 410 1094 428 1126
rect 360 1058 428 1094
rect 360 1026 378 1058
rect 410 1026 428 1058
rect 360 990 428 1026
rect 360 958 378 990
rect 410 958 428 990
rect 360 922 428 958
rect 360 890 378 922
rect 410 890 428 922
rect 360 854 428 890
rect 360 822 378 854
rect 410 822 428 854
rect 360 786 428 822
rect 360 754 378 786
rect 410 754 428 786
rect 360 718 428 754
rect 360 686 378 718
rect 410 686 428 718
rect 360 650 428 686
rect 360 618 378 650
rect 410 618 428 650
rect 360 582 428 618
rect 360 550 378 582
rect 410 550 428 582
rect 5714 1844 5756 1860
rect 5714 1812 5719 1844
rect 5751 1812 5756 1844
rect 5714 1810 5756 1812
rect 5714 622 5715 1810
rect 5755 622 5756 1810
rect 5714 620 5756 622
rect 5714 588 5719 620
rect 5751 588 5756 620
rect 5714 572 5756 588
rect 360 514 428 550
rect 360 482 378 514
rect 410 482 428 514
rect 360 428 428 482
rect 5843 522 5875 1910
rect 6199 1942 6231 3330
rect 6479 3346 6803 3362
rect 6318 3264 6360 3280
rect 6318 3232 6323 3264
rect 6355 3232 6360 3264
rect 6318 3230 6360 3232
rect 6318 2042 6319 3230
rect 6359 2042 6360 3230
rect 6318 2040 6360 2042
rect 6318 2008 6323 2040
rect 6355 2008 6360 2040
rect 6318 1992 6360 2008
rect 5975 1844 6099 1860
rect 5975 1812 6021 1844
rect 6053 1812 6099 1844
rect 5975 1810 6099 1812
rect 5975 622 5976 1810
rect 6098 622 6099 1810
rect 5975 620 6099 622
rect 5975 588 6021 620
rect 6053 588 6099 620
rect 5975 572 6099 588
rect 5843 474 5875 490
rect 6199 522 6231 1910
rect 6447 1942 6479 3330
rect 6835 3346 7051 3362
rect 6579 3264 6703 3280
rect 6579 3232 6625 3264
rect 6657 3232 6703 3264
rect 6579 3230 6703 3232
rect 6579 2042 6580 3230
rect 6702 2042 6703 3230
rect 6579 2040 6703 2042
rect 6579 2008 6625 2040
rect 6657 2008 6703 2040
rect 6579 1992 6703 2008
rect 6318 1844 6360 1860
rect 6318 1812 6323 1844
rect 6355 1812 6360 1844
rect 6318 1810 6360 1812
rect 6318 622 6319 1810
rect 6359 622 6360 1810
rect 6318 620 6360 622
rect 6318 588 6323 620
rect 6355 588 6360 620
rect 6318 572 6360 588
rect 6199 474 6231 490
rect 6447 522 6479 1910
rect 6803 1942 6835 3330
rect 7083 3346 7407 3362
rect 6922 3264 6964 3280
rect 6922 3232 6927 3264
rect 6959 3232 6964 3264
rect 6922 3230 6964 3232
rect 6922 2042 6923 3230
rect 6963 2042 6964 3230
rect 6922 2040 6964 2042
rect 6922 2008 6927 2040
rect 6959 2008 6964 2040
rect 6922 1992 6964 2008
rect 6579 1844 6703 1860
rect 6579 1812 6625 1844
rect 6657 1812 6703 1844
rect 6579 1810 6703 1812
rect 6579 622 6580 1810
rect 6702 622 6703 1810
rect 6579 620 6703 622
rect 6579 588 6625 620
rect 6657 588 6703 620
rect 6579 572 6703 588
rect 6447 474 6479 490
rect 6803 522 6835 1910
rect 7051 1942 7083 3330
rect 7439 3346 7655 3362
rect 7183 3264 7307 3280
rect 7183 3232 7229 3264
rect 7261 3232 7307 3264
rect 7183 3230 7307 3232
rect 7183 2042 7184 3230
rect 7306 2042 7307 3230
rect 7183 2040 7307 2042
rect 7183 2008 7229 2040
rect 7261 2008 7307 2040
rect 7183 1992 7307 2008
rect 6922 1844 6964 1860
rect 6922 1812 6927 1844
rect 6959 1812 6964 1844
rect 6922 1810 6964 1812
rect 6922 622 6923 1810
rect 6963 622 6964 1810
rect 6922 620 6964 622
rect 6922 588 6927 620
rect 6959 588 6964 620
rect 6922 572 6964 588
rect 6803 474 6835 490
rect 7051 522 7083 1910
rect 7407 1942 7439 3330
rect 7687 3346 8011 3362
rect 7526 3264 7568 3280
rect 7526 3232 7531 3264
rect 7563 3232 7568 3264
rect 7526 3230 7568 3232
rect 7526 2042 7527 3230
rect 7567 2042 7568 3230
rect 7526 2040 7568 2042
rect 7526 2008 7531 2040
rect 7563 2008 7568 2040
rect 7526 1992 7568 2008
rect 7183 1844 7307 1860
rect 7183 1812 7229 1844
rect 7261 1812 7307 1844
rect 7183 1810 7307 1812
rect 7183 622 7184 1810
rect 7306 622 7307 1810
rect 7183 620 7307 622
rect 7183 588 7229 620
rect 7261 588 7307 620
rect 7183 572 7307 588
rect 7051 474 7083 490
rect 7407 522 7439 1910
rect 7655 1942 7687 3330
rect 8043 3346 8259 3362
rect 7787 3264 7911 3280
rect 7787 3232 7833 3264
rect 7865 3232 7911 3264
rect 7787 3230 7911 3232
rect 7787 2042 7788 3230
rect 7910 2042 7911 3230
rect 7787 2040 7911 2042
rect 7787 2008 7833 2040
rect 7865 2008 7911 2040
rect 7787 1992 7911 2008
rect 7526 1844 7568 1860
rect 7526 1812 7531 1844
rect 7563 1812 7568 1844
rect 7526 1810 7568 1812
rect 7526 622 7527 1810
rect 7567 622 7568 1810
rect 7526 620 7568 622
rect 7526 588 7531 620
rect 7563 588 7568 620
rect 7526 572 7568 588
rect 7407 474 7439 490
rect 7655 522 7687 1910
rect 8011 1942 8043 3330
rect 8291 3346 8615 3362
rect 8130 3264 8172 3280
rect 8130 3232 8135 3264
rect 8167 3232 8172 3264
rect 8130 3230 8172 3232
rect 8130 2042 8131 3230
rect 8171 2042 8172 3230
rect 8130 2040 8172 2042
rect 8130 2008 8135 2040
rect 8167 2008 8172 2040
rect 8130 1992 8172 2008
rect 7787 1844 7911 1860
rect 7787 1812 7833 1844
rect 7865 1812 7911 1844
rect 7787 1810 7911 1812
rect 7787 622 7788 1810
rect 7910 622 7911 1810
rect 7787 620 7911 622
rect 7787 588 7833 620
rect 7865 588 7911 620
rect 7787 572 7911 588
rect 7655 474 7687 490
rect 8011 522 8043 1910
rect 8259 1942 8291 3330
rect 8647 3346 8863 3362
rect 8391 3264 8515 3280
rect 8391 3232 8437 3264
rect 8469 3232 8515 3264
rect 8391 3230 8515 3232
rect 8391 2042 8392 3230
rect 8514 2042 8515 3230
rect 8391 2040 8515 2042
rect 8391 2008 8437 2040
rect 8469 2008 8515 2040
rect 8391 1992 8515 2008
rect 8130 1844 8172 1860
rect 8130 1812 8135 1844
rect 8167 1812 8172 1844
rect 8130 1810 8172 1812
rect 8130 622 8131 1810
rect 8171 622 8172 1810
rect 8130 620 8172 622
rect 8130 588 8135 620
rect 8167 588 8172 620
rect 8130 572 8172 588
rect 8011 474 8043 490
rect 8259 522 8291 1910
rect 8615 1942 8647 3330
rect 8895 3346 9219 3362
rect 8734 3264 8776 3280
rect 8734 3232 8739 3264
rect 8771 3232 8776 3264
rect 8734 3230 8776 3232
rect 8734 2042 8735 3230
rect 8775 2042 8776 3230
rect 8734 2040 8776 2042
rect 8734 2008 8739 2040
rect 8771 2008 8776 2040
rect 8734 1992 8776 2008
rect 8391 1844 8515 1860
rect 8391 1812 8437 1844
rect 8469 1812 8515 1844
rect 8391 1810 8515 1812
rect 8391 622 8392 1810
rect 8514 622 8515 1810
rect 8391 620 8515 622
rect 8391 588 8437 620
rect 8469 588 8515 620
rect 8391 572 8515 588
rect 8259 474 8291 490
rect 8615 522 8647 1910
rect 8863 1942 8895 3330
rect 9251 3346 9467 3362
rect 8995 3264 9119 3280
rect 8995 3232 9041 3264
rect 9073 3232 9119 3264
rect 8995 3230 9119 3232
rect 8995 2042 8996 3230
rect 9118 2042 9119 3230
rect 8995 2040 9119 2042
rect 8995 2008 9041 2040
rect 9073 2008 9119 2040
rect 8995 1992 9119 2008
rect 8734 1844 8776 1860
rect 8734 1812 8739 1844
rect 8771 1812 8776 1844
rect 8734 1810 8776 1812
rect 8734 622 8735 1810
rect 8775 622 8776 1810
rect 8734 620 8776 622
rect 8734 588 8739 620
rect 8771 588 8776 620
rect 8734 572 8776 588
rect 8615 474 8647 490
rect 8863 522 8895 1910
rect 9219 1942 9251 3330
rect 9499 3346 9823 3362
rect 9338 3264 9380 3280
rect 9338 3232 9343 3264
rect 9375 3232 9380 3264
rect 9338 3230 9380 3232
rect 9338 2042 9339 3230
rect 9379 2042 9380 3230
rect 9338 2040 9380 2042
rect 9338 2008 9343 2040
rect 9375 2008 9380 2040
rect 9338 1992 9380 2008
rect 8995 1844 9119 1860
rect 8995 1812 9041 1844
rect 9073 1812 9119 1844
rect 8995 1810 9119 1812
rect 8995 622 8996 1810
rect 9118 622 9119 1810
rect 8995 620 9119 622
rect 8995 588 9041 620
rect 9073 588 9119 620
rect 8995 572 9119 588
rect 8863 474 8895 490
rect 9219 522 9251 1910
rect 9467 1942 9499 3330
rect 9855 3346 10071 3362
rect 9599 3264 9723 3280
rect 9599 3232 9645 3264
rect 9677 3232 9723 3264
rect 9599 3230 9723 3232
rect 9599 2042 9600 3230
rect 9722 2042 9723 3230
rect 9599 2040 9723 2042
rect 9599 2008 9645 2040
rect 9677 2008 9723 2040
rect 9599 1992 9723 2008
rect 9338 1844 9380 1860
rect 9338 1812 9343 1844
rect 9375 1812 9380 1844
rect 9338 1810 9380 1812
rect 9338 622 9339 1810
rect 9379 622 9380 1810
rect 9338 620 9380 622
rect 9338 588 9343 620
rect 9375 588 9380 620
rect 9338 572 9380 588
rect 9219 474 9251 490
rect 9467 522 9499 1910
rect 9823 1942 9855 3330
rect 9942 3264 9984 3280
rect 9942 3232 9947 3264
rect 9979 3232 9984 3264
rect 9942 3230 9984 3232
rect 9942 2042 9943 3230
rect 9983 2042 9984 3230
rect 9942 2040 9984 2042
rect 9942 2008 9947 2040
rect 9979 2008 9984 2040
rect 9942 1992 9984 2008
rect 9599 1844 9723 1860
rect 9599 1812 9645 1844
rect 9677 1812 9723 1844
rect 9599 1810 9723 1812
rect 9599 622 9600 1810
rect 9722 622 9723 1810
rect 9599 620 9723 622
rect 9599 588 9645 620
rect 9677 588 9723 620
rect 9599 572 9723 588
rect 9467 474 9499 490
rect 9823 522 9855 1910
rect 10071 1942 10103 3330
rect 15572 3370 15640 3424
rect 15572 3338 15590 3370
rect 15622 3338 15640 3370
rect 15572 3302 15640 3338
rect 10203 3264 10327 3280
rect 10203 3232 10249 3264
rect 10281 3232 10327 3264
rect 10203 3230 10327 3232
rect 10203 2042 10204 3230
rect 10326 2042 10327 3230
rect 10203 2040 10327 2042
rect 10203 2008 10249 2040
rect 10281 2008 10327 2040
rect 10203 1992 10327 2008
rect 15572 3270 15590 3302
rect 15622 3270 15640 3302
rect 15572 3234 15640 3270
rect 15572 3202 15590 3234
rect 15622 3202 15640 3234
rect 15572 3166 15640 3202
rect 15572 3134 15590 3166
rect 15622 3134 15640 3166
rect 15572 3098 15640 3134
rect 15572 3066 15590 3098
rect 15622 3066 15640 3098
rect 15572 3030 15640 3066
rect 15572 2998 15590 3030
rect 15622 2998 15640 3030
rect 15572 2962 15640 2998
rect 15572 2930 15590 2962
rect 15622 2930 15640 2962
rect 15572 2894 15640 2930
rect 15572 2862 15590 2894
rect 15622 2862 15640 2894
rect 15572 2826 15640 2862
rect 15572 2794 15590 2826
rect 15622 2794 15640 2826
rect 15572 2758 15640 2794
rect 15572 2726 15590 2758
rect 15622 2726 15640 2758
rect 15572 2690 15640 2726
rect 15572 2658 15590 2690
rect 15622 2658 15640 2690
rect 15572 2622 15640 2658
rect 15572 2590 15590 2622
rect 15622 2590 15640 2622
rect 15572 2554 15640 2590
rect 15572 2522 15590 2554
rect 15622 2522 15640 2554
rect 15572 2486 15640 2522
rect 15572 2454 15590 2486
rect 15622 2454 15640 2486
rect 15572 2418 15640 2454
rect 15572 2386 15590 2418
rect 15622 2386 15640 2418
rect 15572 2350 15640 2386
rect 15572 2318 15590 2350
rect 15622 2318 15640 2350
rect 15572 2282 15640 2318
rect 15572 2250 15590 2282
rect 15622 2250 15640 2282
rect 15572 2214 15640 2250
rect 15572 2182 15590 2214
rect 15622 2182 15640 2214
rect 15572 2146 15640 2182
rect 15572 2114 15590 2146
rect 15622 2114 15640 2146
rect 15572 2078 15640 2114
rect 15572 2046 15590 2078
rect 15622 2046 15640 2078
rect 15572 2010 15640 2046
rect 9942 1844 9984 1860
rect 9942 1812 9947 1844
rect 9979 1812 9984 1844
rect 9942 1810 9984 1812
rect 9942 622 9943 1810
rect 9983 622 9984 1810
rect 9942 620 9984 622
rect 9942 588 9947 620
rect 9979 588 9984 620
rect 9942 572 9984 588
rect 9823 474 9855 490
rect 10071 522 10103 1910
rect 15572 1978 15590 2010
rect 15622 1978 15640 2010
rect 15572 1942 15640 1978
rect 15572 1910 15590 1942
rect 15622 1910 15640 1942
rect 15572 1874 15640 1910
rect 10203 1844 10327 1860
rect 10203 1812 10249 1844
rect 10281 1812 10327 1844
rect 10203 1810 10327 1812
rect 10203 622 10204 1810
rect 10326 622 10327 1810
rect 10203 620 10327 622
rect 10203 588 10249 620
rect 10281 588 10327 620
rect 10203 572 10327 588
rect 15572 1842 15590 1874
rect 15622 1842 15640 1874
rect 15572 1806 15640 1842
rect 15572 1774 15590 1806
rect 15622 1774 15640 1806
rect 15572 1738 15640 1774
rect 15572 1706 15590 1738
rect 15622 1706 15640 1738
rect 15572 1670 15640 1706
rect 15572 1638 15590 1670
rect 15622 1638 15640 1670
rect 15572 1602 15640 1638
rect 15572 1570 15590 1602
rect 15622 1570 15640 1602
rect 15572 1534 15640 1570
rect 15572 1502 15590 1534
rect 15622 1502 15640 1534
rect 15572 1466 15640 1502
rect 15572 1434 15590 1466
rect 15622 1434 15640 1466
rect 15572 1398 15640 1434
rect 15572 1366 15590 1398
rect 15622 1366 15640 1398
rect 15572 1330 15640 1366
rect 15572 1298 15590 1330
rect 15622 1298 15640 1330
rect 15572 1262 15640 1298
rect 15572 1230 15590 1262
rect 15622 1230 15640 1262
rect 15572 1194 15640 1230
rect 15572 1162 15590 1194
rect 15622 1162 15640 1194
rect 15572 1126 15640 1162
rect 15572 1094 15590 1126
rect 15622 1094 15640 1126
rect 15572 1058 15640 1094
rect 15572 1026 15590 1058
rect 15622 1026 15640 1058
rect 15572 990 15640 1026
rect 15572 958 15590 990
rect 15622 958 15640 990
rect 15572 922 15640 958
rect 15572 890 15590 922
rect 15622 890 15640 922
rect 15572 854 15640 890
rect 15572 822 15590 854
rect 15622 822 15640 854
rect 15572 786 15640 822
rect 15572 754 15590 786
rect 15622 754 15640 786
rect 15572 718 15640 754
rect 15572 686 15590 718
rect 15622 686 15640 718
rect 15572 650 15640 686
rect 15572 618 15590 650
rect 15622 618 15640 650
rect 15572 582 15640 618
rect 10071 474 10103 490
rect 15572 550 15590 582
rect 15622 550 15640 582
rect 15572 514 15640 550
rect 15572 482 15590 514
rect 15622 482 15640 514
rect 15572 428 15640 482
rect 360 414 15640 428
rect 360 410 5715 414
rect 5755 410 6319 414
rect 6359 410 6923 414
rect 6963 410 7527 414
rect 7567 410 8131 414
rect 8171 410 8735 414
rect 8775 410 9339 414
rect 9379 410 9943 414
rect 9983 410 15640 414
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5755 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6359 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6923 410
rect 6963 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7527 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8131 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8735 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9983 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 374 5715 378
rect 5755 374 6319 378
rect 6359 374 6923 378
rect 6963 374 7527 378
rect 7567 374 8131 378
rect 8171 374 8735 378
rect 8775 374 9339 378
rect 9379 374 9943 378
rect 9983 374 15640 378
rect 360 360 15640 374
rect 15932 3472 16000 3508
rect 15932 3440 15950 3472
rect 15982 3440 16000 3472
rect 15932 3404 16000 3440
rect 15932 3372 15950 3404
rect 15982 3372 16000 3404
rect 15932 3336 16000 3372
rect 15932 3304 15950 3336
rect 15982 3304 16000 3336
rect 15932 3268 16000 3304
rect 15932 3236 15950 3268
rect 15982 3236 16000 3268
rect 15932 3200 16000 3236
rect 15932 3168 15950 3200
rect 15982 3168 16000 3200
rect 15932 3132 16000 3168
rect 15932 3100 15950 3132
rect 15982 3100 16000 3132
rect 15932 3064 16000 3100
rect 15932 3032 15950 3064
rect 15982 3032 16000 3064
rect 15932 2996 16000 3032
rect 15932 2964 15950 2996
rect 15982 2964 16000 2996
rect 15932 2928 16000 2964
rect 15932 2896 15950 2928
rect 15982 2896 16000 2928
rect 15932 2860 16000 2896
rect 15932 2828 15950 2860
rect 15982 2828 16000 2860
rect 15932 2792 16000 2828
rect 15932 2760 15950 2792
rect 15982 2760 16000 2792
rect 15932 2724 16000 2760
rect 15932 2692 15950 2724
rect 15982 2692 16000 2724
rect 15932 2656 16000 2692
rect 15932 2624 15950 2656
rect 15982 2624 16000 2656
rect 15932 2588 16000 2624
rect 15932 2556 15950 2588
rect 15982 2556 16000 2588
rect 15932 2520 16000 2556
rect 15932 2488 15950 2520
rect 15982 2488 16000 2520
rect 15932 2452 16000 2488
rect 15932 2420 15950 2452
rect 15982 2420 16000 2452
rect 15932 2384 16000 2420
rect 15932 2352 15950 2384
rect 15982 2352 16000 2384
rect 15932 2316 16000 2352
rect 15932 2284 15950 2316
rect 15982 2284 16000 2316
rect 15932 2248 16000 2284
rect 15932 2216 15950 2248
rect 15982 2216 16000 2248
rect 15932 2180 16000 2216
rect 15932 2148 15950 2180
rect 15982 2148 16000 2180
rect 15932 2112 16000 2148
rect 15932 2080 15950 2112
rect 15982 2080 16000 2112
rect 15932 2044 16000 2080
rect 15932 2012 15950 2044
rect 15982 2012 16000 2044
rect 15932 1976 16000 2012
rect 15932 1944 15950 1976
rect 15982 1944 16000 1976
rect 15932 1908 16000 1944
rect 15932 1876 15950 1908
rect 15982 1876 16000 1908
rect 15932 1840 16000 1876
rect 15932 1808 15950 1840
rect 15982 1808 16000 1840
rect 15932 1772 16000 1808
rect 15932 1740 15950 1772
rect 15982 1740 16000 1772
rect 15932 1704 16000 1740
rect 15932 1672 15950 1704
rect 15982 1672 16000 1704
rect 15932 1636 16000 1672
rect 15932 1604 15950 1636
rect 15982 1604 16000 1636
rect 15932 1568 16000 1604
rect 15932 1536 15950 1568
rect 15982 1536 16000 1568
rect 15932 1500 16000 1536
rect 15932 1468 15950 1500
rect 15982 1468 16000 1500
rect 15932 1432 16000 1468
rect 15932 1400 15950 1432
rect 15982 1400 16000 1432
rect 15932 1364 16000 1400
rect 15932 1332 15950 1364
rect 15982 1332 16000 1364
rect 15932 1296 16000 1332
rect 15932 1264 15950 1296
rect 15982 1264 16000 1296
rect 15932 1228 16000 1264
rect 15932 1196 15950 1228
rect 15982 1196 16000 1228
rect 15932 1160 16000 1196
rect 15932 1128 15950 1160
rect 15982 1128 16000 1160
rect 15932 1092 16000 1128
rect 15932 1060 15950 1092
rect 15982 1060 16000 1092
rect 15932 1024 16000 1060
rect 15932 992 15950 1024
rect 15982 992 16000 1024
rect 15932 956 16000 992
rect 15932 924 15950 956
rect 15982 924 16000 956
rect 15932 888 16000 924
rect 15932 856 15950 888
rect 15982 856 16000 888
rect 15932 820 16000 856
rect 15932 788 15950 820
rect 15982 788 16000 820
rect 15932 752 16000 788
rect 15932 720 15950 752
rect 15982 720 16000 752
rect 15932 684 16000 720
rect 15932 652 15950 684
rect 15982 652 16000 684
rect 15932 616 16000 652
rect 15932 584 15950 616
rect 15982 584 16000 616
rect 15932 548 16000 584
rect 15932 516 15950 548
rect 15982 516 16000 548
rect 15932 480 16000 516
rect 15932 448 15950 480
rect 15982 448 16000 480
rect 15932 412 16000 448
rect 15932 380 15950 412
rect 15982 380 16000 412
rect 0 312 18 344
rect 50 312 68 344
rect 0 276 68 312
rect 0 244 18 276
rect 50 244 68 276
rect 0 208 68 244
rect 0 176 18 208
rect 50 176 68 208
rect 0 140 68 176
rect 0 108 18 140
rect 50 108 68 140
rect 0 68 68 108
rect 15932 344 16000 380
rect 15932 312 15950 344
rect 15982 312 16000 344
rect 15932 276 16000 312
rect 15932 244 15950 276
rect 15982 244 16000 276
rect 15932 208 16000 244
rect 15932 176 15950 208
rect 15982 176 16000 208
rect 15932 140 16000 176
rect 15932 108 15950 140
rect 15982 108 16000 140
rect 15932 68 16000 108
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 5715 3474 5755 3478
rect 6319 3474 6359 3478
rect 6923 3474 6963 3478
rect 7527 3474 7567 3478
rect 8131 3474 8171 3478
rect 8735 3474 8775 3478
rect 9339 3474 9379 3478
rect 9943 3474 9983 3478
rect 5715 3442 5738 3474
rect 5738 3442 5755 3474
rect 6319 3442 6350 3474
rect 6350 3442 6359 3474
rect 6923 3442 6930 3474
rect 6930 3442 6962 3474
rect 6962 3442 6963 3474
rect 7527 3442 7542 3474
rect 7542 3442 7567 3474
rect 8131 3442 8154 3474
rect 8154 3442 8171 3474
rect 8735 3442 8766 3474
rect 8766 3442 8775 3474
rect 9339 3442 9342 3474
rect 9342 3442 9378 3474
rect 9378 3442 9379 3474
rect 9943 3442 9954 3474
rect 9954 3442 9983 3474
rect 5715 3438 5755 3442
rect 6319 3438 6359 3442
rect 6923 3438 6963 3442
rect 7527 3438 7567 3442
rect 8131 3438 8171 3442
rect 8735 3438 8775 3442
rect 9339 3438 9379 3442
rect 9943 3438 9983 3442
rect 3046 3319 3086 3359
rect 3046 3223 3086 3263
rect 5715 3196 5755 3230
rect 5715 3164 5719 3196
rect 5719 3164 5751 3196
rect 5751 3164 5755 3196
rect 5715 3128 5755 3164
rect 5715 3096 5719 3128
rect 5719 3096 5751 3128
rect 5751 3096 5755 3128
rect 5715 3060 5755 3096
rect 5715 3028 5719 3060
rect 5719 3028 5751 3060
rect 5751 3028 5755 3060
rect 5715 2992 5755 3028
rect 5715 2960 5719 2992
rect 5719 2960 5751 2992
rect 5751 2960 5755 2992
rect 5715 2924 5755 2960
rect 5715 2892 5719 2924
rect 5719 2892 5751 2924
rect 5751 2892 5755 2924
rect 5715 2856 5755 2892
rect 5715 2824 5719 2856
rect 5719 2824 5751 2856
rect 5751 2824 5755 2856
rect 5715 2788 5755 2824
rect 5715 2756 5719 2788
rect 5719 2756 5751 2788
rect 5751 2756 5755 2788
rect 5715 2720 5755 2756
rect 5715 2688 5719 2720
rect 5719 2688 5751 2720
rect 5751 2688 5755 2720
rect 5715 2652 5755 2688
rect 5715 2620 5719 2652
rect 5719 2620 5751 2652
rect 5751 2620 5755 2652
rect 5715 2584 5755 2620
rect 5715 2552 5719 2584
rect 5719 2552 5751 2584
rect 5751 2552 5755 2584
rect 5715 2516 5755 2552
rect 5715 2484 5719 2516
rect 5719 2484 5751 2516
rect 5751 2484 5755 2516
rect 5715 2448 5755 2484
rect 5715 2416 5719 2448
rect 5719 2416 5751 2448
rect 5751 2416 5755 2448
rect 5715 2380 5755 2416
rect 5715 2348 5719 2380
rect 5719 2348 5751 2380
rect 5751 2348 5755 2380
rect 5715 2312 5755 2348
rect 5715 2280 5719 2312
rect 5719 2280 5751 2312
rect 5751 2280 5755 2312
rect 5715 2244 5755 2280
rect 5715 2212 5719 2244
rect 5719 2212 5751 2244
rect 5751 2212 5755 2244
rect 5715 2176 5755 2212
rect 5715 2144 5719 2176
rect 5719 2144 5751 2176
rect 5751 2144 5755 2176
rect 5715 2108 5755 2144
rect 5715 2076 5719 2108
rect 5719 2076 5751 2108
rect 5751 2076 5755 2108
rect 5715 2042 5755 2076
rect 5976 3196 6098 3230
rect 5976 3164 6021 3196
rect 6021 3164 6053 3196
rect 6053 3164 6098 3196
rect 5976 3128 6098 3164
rect 5976 3096 6021 3128
rect 6021 3096 6053 3128
rect 6053 3096 6098 3128
rect 5976 3060 6098 3096
rect 5976 3028 6021 3060
rect 6021 3028 6053 3060
rect 6053 3028 6098 3060
rect 5976 2992 6098 3028
rect 5976 2960 6021 2992
rect 6021 2960 6053 2992
rect 6053 2960 6098 2992
rect 5976 2924 6098 2960
rect 5976 2892 6021 2924
rect 6021 2892 6053 2924
rect 6053 2892 6098 2924
rect 5976 2856 6098 2892
rect 5976 2824 6021 2856
rect 6021 2824 6053 2856
rect 6053 2824 6098 2856
rect 5976 2788 6098 2824
rect 5976 2756 6021 2788
rect 6021 2756 6053 2788
rect 6053 2756 6098 2788
rect 5976 2720 6098 2756
rect 5976 2688 6021 2720
rect 6021 2688 6053 2720
rect 6053 2688 6098 2720
rect 5976 2652 6098 2688
rect 5976 2620 6021 2652
rect 6021 2620 6053 2652
rect 6053 2620 6098 2652
rect 5976 2584 6098 2620
rect 5976 2552 6021 2584
rect 6021 2552 6053 2584
rect 6053 2552 6098 2584
rect 5976 2516 6098 2552
rect 5976 2484 6021 2516
rect 6021 2484 6053 2516
rect 6053 2484 6098 2516
rect 5976 2448 6098 2484
rect 5976 2416 6021 2448
rect 6021 2416 6053 2448
rect 6053 2416 6098 2448
rect 5976 2380 6098 2416
rect 5976 2348 6021 2380
rect 6021 2348 6053 2380
rect 6053 2348 6098 2380
rect 5976 2312 6098 2348
rect 5976 2280 6021 2312
rect 6021 2280 6053 2312
rect 6053 2280 6098 2312
rect 5976 2244 6098 2280
rect 5976 2212 6021 2244
rect 6021 2212 6053 2244
rect 6053 2212 6098 2244
rect 5976 2176 6098 2212
rect 5976 2144 6021 2176
rect 6021 2144 6053 2176
rect 6053 2144 6098 2176
rect 5976 2108 6098 2144
rect 5976 2076 6021 2108
rect 6021 2076 6053 2108
rect 6053 2076 6098 2108
rect 5976 2042 6098 2076
rect 5715 1776 5755 1810
rect 5715 1744 5719 1776
rect 5719 1744 5751 1776
rect 5751 1744 5755 1776
rect 5715 1708 5755 1744
rect 5715 1676 5719 1708
rect 5719 1676 5751 1708
rect 5751 1676 5755 1708
rect 5715 1640 5755 1676
rect 5715 1608 5719 1640
rect 5719 1608 5751 1640
rect 5751 1608 5755 1640
rect 5715 1572 5755 1608
rect 5715 1540 5719 1572
rect 5719 1540 5751 1572
rect 5751 1540 5755 1572
rect 5715 1504 5755 1540
rect 5715 1472 5719 1504
rect 5719 1472 5751 1504
rect 5751 1472 5755 1504
rect 5715 1436 5755 1472
rect 5715 1404 5719 1436
rect 5719 1404 5751 1436
rect 5751 1404 5755 1436
rect 5715 1368 5755 1404
rect 5715 1336 5719 1368
rect 5719 1336 5751 1368
rect 5751 1336 5755 1368
rect 5715 1300 5755 1336
rect 5715 1268 5719 1300
rect 5719 1268 5751 1300
rect 5751 1268 5755 1300
rect 5715 1232 5755 1268
rect 5715 1200 5719 1232
rect 5719 1200 5751 1232
rect 5751 1200 5755 1232
rect 5715 1164 5755 1200
rect 5715 1132 5719 1164
rect 5719 1132 5751 1164
rect 5751 1132 5755 1164
rect 5715 1096 5755 1132
rect 5715 1064 5719 1096
rect 5719 1064 5751 1096
rect 5751 1064 5755 1096
rect 5715 1028 5755 1064
rect 5715 996 5719 1028
rect 5719 996 5751 1028
rect 5751 996 5755 1028
rect 5715 960 5755 996
rect 5715 928 5719 960
rect 5719 928 5751 960
rect 5751 928 5755 960
rect 5715 892 5755 928
rect 5715 860 5719 892
rect 5719 860 5751 892
rect 5751 860 5755 892
rect 5715 824 5755 860
rect 5715 792 5719 824
rect 5719 792 5751 824
rect 5751 792 5755 824
rect 5715 756 5755 792
rect 5715 724 5719 756
rect 5719 724 5751 756
rect 5751 724 5755 756
rect 5715 688 5755 724
rect 5715 656 5719 688
rect 5719 656 5751 688
rect 5751 656 5755 688
rect 5715 622 5755 656
rect 6319 3196 6359 3230
rect 6319 3164 6323 3196
rect 6323 3164 6355 3196
rect 6355 3164 6359 3196
rect 6319 3128 6359 3164
rect 6319 3096 6323 3128
rect 6323 3096 6355 3128
rect 6355 3096 6359 3128
rect 6319 3060 6359 3096
rect 6319 3028 6323 3060
rect 6323 3028 6355 3060
rect 6355 3028 6359 3060
rect 6319 2992 6359 3028
rect 6319 2960 6323 2992
rect 6323 2960 6355 2992
rect 6355 2960 6359 2992
rect 6319 2924 6359 2960
rect 6319 2892 6323 2924
rect 6323 2892 6355 2924
rect 6355 2892 6359 2924
rect 6319 2856 6359 2892
rect 6319 2824 6323 2856
rect 6323 2824 6355 2856
rect 6355 2824 6359 2856
rect 6319 2788 6359 2824
rect 6319 2756 6323 2788
rect 6323 2756 6355 2788
rect 6355 2756 6359 2788
rect 6319 2720 6359 2756
rect 6319 2688 6323 2720
rect 6323 2688 6355 2720
rect 6355 2688 6359 2720
rect 6319 2652 6359 2688
rect 6319 2620 6323 2652
rect 6323 2620 6355 2652
rect 6355 2620 6359 2652
rect 6319 2584 6359 2620
rect 6319 2552 6323 2584
rect 6323 2552 6355 2584
rect 6355 2552 6359 2584
rect 6319 2516 6359 2552
rect 6319 2484 6323 2516
rect 6323 2484 6355 2516
rect 6355 2484 6359 2516
rect 6319 2448 6359 2484
rect 6319 2416 6323 2448
rect 6323 2416 6355 2448
rect 6355 2416 6359 2448
rect 6319 2380 6359 2416
rect 6319 2348 6323 2380
rect 6323 2348 6355 2380
rect 6355 2348 6359 2380
rect 6319 2312 6359 2348
rect 6319 2280 6323 2312
rect 6323 2280 6355 2312
rect 6355 2280 6359 2312
rect 6319 2244 6359 2280
rect 6319 2212 6323 2244
rect 6323 2212 6355 2244
rect 6355 2212 6359 2244
rect 6319 2176 6359 2212
rect 6319 2144 6323 2176
rect 6323 2144 6355 2176
rect 6355 2144 6359 2176
rect 6319 2108 6359 2144
rect 6319 2076 6323 2108
rect 6323 2076 6355 2108
rect 6355 2076 6359 2108
rect 6319 2042 6359 2076
rect 5976 1776 6098 1810
rect 5976 1744 6021 1776
rect 6021 1744 6053 1776
rect 6053 1744 6098 1776
rect 5976 1708 6098 1744
rect 5976 1676 6021 1708
rect 6021 1676 6053 1708
rect 6053 1676 6098 1708
rect 5976 1640 6098 1676
rect 5976 1608 6021 1640
rect 6021 1608 6053 1640
rect 6053 1608 6098 1640
rect 5976 1572 6098 1608
rect 5976 1540 6021 1572
rect 6021 1540 6053 1572
rect 6053 1540 6098 1572
rect 5976 1504 6098 1540
rect 5976 1472 6021 1504
rect 6021 1472 6053 1504
rect 6053 1472 6098 1504
rect 5976 1436 6098 1472
rect 5976 1404 6021 1436
rect 6021 1404 6053 1436
rect 6053 1404 6098 1436
rect 5976 1368 6098 1404
rect 5976 1336 6021 1368
rect 6021 1336 6053 1368
rect 6053 1336 6098 1368
rect 5976 1300 6098 1336
rect 5976 1268 6021 1300
rect 6021 1268 6053 1300
rect 6053 1268 6098 1300
rect 5976 1232 6098 1268
rect 5976 1200 6021 1232
rect 6021 1200 6053 1232
rect 6053 1200 6098 1232
rect 5976 1164 6098 1200
rect 5976 1132 6021 1164
rect 6021 1132 6053 1164
rect 6053 1132 6098 1164
rect 5976 1096 6098 1132
rect 5976 1064 6021 1096
rect 6021 1064 6053 1096
rect 6053 1064 6098 1096
rect 5976 1028 6098 1064
rect 5976 996 6021 1028
rect 6021 996 6053 1028
rect 6053 996 6098 1028
rect 5976 960 6098 996
rect 5976 928 6021 960
rect 6021 928 6053 960
rect 6053 928 6098 960
rect 5976 892 6098 928
rect 5976 860 6021 892
rect 6021 860 6053 892
rect 6053 860 6098 892
rect 5976 824 6098 860
rect 5976 792 6021 824
rect 6021 792 6053 824
rect 6053 792 6098 824
rect 5976 756 6098 792
rect 5976 724 6021 756
rect 6021 724 6053 756
rect 6053 724 6098 756
rect 5976 688 6098 724
rect 5976 656 6021 688
rect 6021 656 6053 688
rect 6053 656 6098 688
rect 5976 622 6098 656
rect 6580 3196 6702 3230
rect 6580 3164 6625 3196
rect 6625 3164 6657 3196
rect 6657 3164 6702 3196
rect 6580 3128 6702 3164
rect 6580 3096 6625 3128
rect 6625 3096 6657 3128
rect 6657 3096 6702 3128
rect 6580 3060 6702 3096
rect 6580 3028 6625 3060
rect 6625 3028 6657 3060
rect 6657 3028 6702 3060
rect 6580 2992 6702 3028
rect 6580 2960 6625 2992
rect 6625 2960 6657 2992
rect 6657 2960 6702 2992
rect 6580 2924 6702 2960
rect 6580 2892 6625 2924
rect 6625 2892 6657 2924
rect 6657 2892 6702 2924
rect 6580 2856 6702 2892
rect 6580 2824 6625 2856
rect 6625 2824 6657 2856
rect 6657 2824 6702 2856
rect 6580 2788 6702 2824
rect 6580 2756 6625 2788
rect 6625 2756 6657 2788
rect 6657 2756 6702 2788
rect 6580 2720 6702 2756
rect 6580 2688 6625 2720
rect 6625 2688 6657 2720
rect 6657 2688 6702 2720
rect 6580 2652 6702 2688
rect 6580 2620 6625 2652
rect 6625 2620 6657 2652
rect 6657 2620 6702 2652
rect 6580 2584 6702 2620
rect 6580 2552 6625 2584
rect 6625 2552 6657 2584
rect 6657 2552 6702 2584
rect 6580 2516 6702 2552
rect 6580 2484 6625 2516
rect 6625 2484 6657 2516
rect 6657 2484 6702 2516
rect 6580 2448 6702 2484
rect 6580 2416 6625 2448
rect 6625 2416 6657 2448
rect 6657 2416 6702 2448
rect 6580 2380 6702 2416
rect 6580 2348 6625 2380
rect 6625 2348 6657 2380
rect 6657 2348 6702 2380
rect 6580 2312 6702 2348
rect 6580 2280 6625 2312
rect 6625 2280 6657 2312
rect 6657 2280 6702 2312
rect 6580 2244 6702 2280
rect 6580 2212 6625 2244
rect 6625 2212 6657 2244
rect 6657 2212 6702 2244
rect 6580 2176 6702 2212
rect 6580 2144 6625 2176
rect 6625 2144 6657 2176
rect 6657 2144 6702 2176
rect 6580 2108 6702 2144
rect 6580 2076 6625 2108
rect 6625 2076 6657 2108
rect 6657 2076 6702 2108
rect 6580 2042 6702 2076
rect 6319 1776 6359 1810
rect 6319 1744 6323 1776
rect 6323 1744 6355 1776
rect 6355 1744 6359 1776
rect 6319 1708 6359 1744
rect 6319 1676 6323 1708
rect 6323 1676 6355 1708
rect 6355 1676 6359 1708
rect 6319 1640 6359 1676
rect 6319 1608 6323 1640
rect 6323 1608 6355 1640
rect 6355 1608 6359 1640
rect 6319 1572 6359 1608
rect 6319 1540 6323 1572
rect 6323 1540 6355 1572
rect 6355 1540 6359 1572
rect 6319 1504 6359 1540
rect 6319 1472 6323 1504
rect 6323 1472 6355 1504
rect 6355 1472 6359 1504
rect 6319 1436 6359 1472
rect 6319 1404 6323 1436
rect 6323 1404 6355 1436
rect 6355 1404 6359 1436
rect 6319 1368 6359 1404
rect 6319 1336 6323 1368
rect 6323 1336 6355 1368
rect 6355 1336 6359 1368
rect 6319 1300 6359 1336
rect 6319 1268 6323 1300
rect 6323 1268 6355 1300
rect 6355 1268 6359 1300
rect 6319 1232 6359 1268
rect 6319 1200 6323 1232
rect 6323 1200 6355 1232
rect 6355 1200 6359 1232
rect 6319 1164 6359 1200
rect 6319 1132 6323 1164
rect 6323 1132 6355 1164
rect 6355 1132 6359 1164
rect 6319 1096 6359 1132
rect 6319 1064 6323 1096
rect 6323 1064 6355 1096
rect 6355 1064 6359 1096
rect 6319 1028 6359 1064
rect 6319 996 6323 1028
rect 6323 996 6355 1028
rect 6355 996 6359 1028
rect 6319 960 6359 996
rect 6319 928 6323 960
rect 6323 928 6355 960
rect 6355 928 6359 960
rect 6319 892 6359 928
rect 6319 860 6323 892
rect 6323 860 6355 892
rect 6355 860 6359 892
rect 6319 824 6359 860
rect 6319 792 6323 824
rect 6323 792 6355 824
rect 6355 792 6359 824
rect 6319 756 6359 792
rect 6319 724 6323 756
rect 6323 724 6355 756
rect 6355 724 6359 756
rect 6319 688 6359 724
rect 6319 656 6323 688
rect 6323 656 6355 688
rect 6355 656 6359 688
rect 6319 622 6359 656
rect 6923 3196 6963 3230
rect 6923 3164 6927 3196
rect 6927 3164 6959 3196
rect 6959 3164 6963 3196
rect 6923 3128 6963 3164
rect 6923 3096 6927 3128
rect 6927 3096 6959 3128
rect 6959 3096 6963 3128
rect 6923 3060 6963 3096
rect 6923 3028 6927 3060
rect 6927 3028 6959 3060
rect 6959 3028 6963 3060
rect 6923 2992 6963 3028
rect 6923 2960 6927 2992
rect 6927 2960 6959 2992
rect 6959 2960 6963 2992
rect 6923 2924 6963 2960
rect 6923 2892 6927 2924
rect 6927 2892 6959 2924
rect 6959 2892 6963 2924
rect 6923 2856 6963 2892
rect 6923 2824 6927 2856
rect 6927 2824 6959 2856
rect 6959 2824 6963 2856
rect 6923 2788 6963 2824
rect 6923 2756 6927 2788
rect 6927 2756 6959 2788
rect 6959 2756 6963 2788
rect 6923 2720 6963 2756
rect 6923 2688 6927 2720
rect 6927 2688 6959 2720
rect 6959 2688 6963 2720
rect 6923 2652 6963 2688
rect 6923 2620 6927 2652
rect 6927 2620 6959 2652
rect 6959 2620 6963 2652
rect 6923 2584 6963 2620
rect 6923 2552 6927 2584
rect 6927 2552 6959 2584
rect 6959 2552 6963 2584
rect 6923 2516 6963 2552
rect 6923 2484 6927 2516
rect 6927 2484 6959 2516
rect 6959 2484 6963 2516
rect 6923 2448 6963 2484
rect 6923 2416 6927 2448
rect 6927 2416 6959 2448
rect 6959 2416 6963 2448
rect 6923 2380 6963 2416
rect 6923 2348 6927 2380
rect 6927 2348 6959 2380
rect 6959 2348 6963 2380
rect 6923 2312 6963 2348
rect 6923 2280 6927 2312
rect 6927 2280 6959 2312
rect 6959 2280 6963 2312
rect 6923 2244 6963 2280
rect 6923 2212 6927 2244
rect 6927 2212 6959 2244
rect 6959 2212 6963 2244
rect 6923 2176 6963 2212
rect 6923 2144 6927 2176
rect 6927 2144 6959 2176
rect 6959 2144 6963 2176
rect 6923 2108 6963 2144
rect 6923 2076 6927 2108
rect 6927 2076 6959 2108
rect 6959 2076 6963 2108
rect 6923 2042 6963 2076
rect 6580 1776 6702 1810
rect 6580 1744 6625 1776
rect 6625 1744 6657 1776
rect 6657 1744 6702 1776
rect 6580 1708 6702 1744
rect 6580 1676 6625 1708
rect 6625 1676 6657 1708
rect 6657 1676 6702 1708
rect 6580 1640 6702 1676
rect 6580 1608 6625 1640
rect 6625 1608 6657 1640
rect 6657 1608 6702 1640
rect 6580 1572 6702 1608
rect 6580 1540 6625 1572
rect 6625 1540 6657 1572
rect 6657 1540 6702 1572
rect 6580 1504 6702 1540
rect 6580 1472 6625 1504
rect 6625 1472 6657 1504
rect 6657 1472 6702 1504
rect 6580 1436 6702 1472
rect 6580 1404 6625 1436
rect 6625 1404 6657 1436
rect 6657 1404 6702 1436
rect 6580 1368 6702 1404
rect 6580 1336 6625 1368
rect 6625 1336 6657 1368
rect 6657 1336 6702 1368
rect 6580 1300 6702 1336
rect 6580 1268 6625 1300
rect 6625 1268 6657 1300
rect 6657 1268 6702 1300
rect 6580 1232 6702 1268
rect 6580 1200 6625 1232
rect 6625 1200 6657 1232
rect 6657 1200 6702 1232
rect 6580 1164 6702 1200
rect 6580 1132 6625 1164
rect 6625 1132 6657 1164
rect 6657 1132 6702 1164
rect 6580 1096 6702 1132
rect 6580 1064 6625 1096
rect 6625 1064 6657 1096
rect 6657 1064 6702 1096
rect 6580 1028 6702 1064
rect 6580 996 6625 1028
rect 6625 996 6657 1028
rect 6657 996 6702 1028
rect 6580 960 6702 996
rect 6580 928 6625 960
rect 6625 928 6657 960
rect 6657 928 6702 960
rect 6580 892 6702 928
rect 6580 860 6625 892
rect 6625 860 6657 892
rect 6657 860 6702 892
rect 6580 824 6702 860
rect 6580 792 6625 824
rect 6625 792 6657 824
rect 6657 792 6702 824
rect 6580 756 6702 792
rect 6580 724 6625 756
rect 6625 724 6657 756
rect 6657 724 6702 756
rect 6580 688 6702 724
rect 6580 656 6625 688
rect 6625 656 6657 688
rect 6657 656 6702 688
rect 6580 622 6702 656
rect 7184 3196 7306 3230
rect 7184 3164 7229 3196
rect 7229 3164 7261 3196
rect 7261 3164 7306 3196
rect 7184 3128 7306 3164
rect 7184 3096 7229 3128
rect 7229 3096 7261 3128
rect 7261 3096 7306 3128
rect 7184 3060 7306 3096
rect 7184 3028 7229 3060
rect 7229 3028 7261 3060
rect 7261 3028 7306 3060
rect 7184 2992 7306 3028
rect 7184 2960 7229 2992
rect 7229 2960 7261 2992
rect 7261 2960 7306 2992
rect 7184 2924 7306 2960
rect 7184 2892 7229 2924
rect 7229 2892 7261 2924
rect 7261 2892 7306 2924
rect 7184 2856 7306 2892
rect 7184 2824 7229 2856
rect 7229 2824 7261 2856
rect 7261 2824 7306 2856
rect 7184 2788 7306 2824
rect 7184 2756 7229 2788
rect 7229 2756 7261 2788
rect 7261 2756 7306 2788
rect 7184 2720 7306 2756
rect 7184 2688 7229 2720
rect 7229 2688 7261 2720
rect 7261 2688 7306 2720
rect 7184 2652 7306 2688
rect 7184 2620 7229 2652
rect 7229 2620 7261 2652
rect 7261 2620 7306 2652
rect 7184 2584 7306 2620
rect 7184 2552 7229 2584
rect 7229 2552 7261 2584
rect 7261 2552 7306 2584
rect 7184 2516 7306 2552
rect 7184 2484 7229 2516
rect 7229 2484 7261 2516
rect 7261 2484 7306 2516
rect 7184 2448 7306 2484
rect 7184 2416 7229 2448
rect 7229 2416 7261 2448
rect 7261 2416 7306 2448
rect 7184 2380 7306 2416
rect 7184 2348 7229 2380
rect 7229 2348 7261 2380
rect 7261 2348 7306 2380
rect 7184 2312 7306 2348
rect 7184 2280 7229 2312
rect 7229 2280 7261 2312
rect 7261 2280 7306 2312
rect 7184 2244 7306 2280
rect 7184 2212 7229 2244
rect 7229 2212 7261 2244
rect 7261 2212 7306 2244
rect 7184 2176 7306 2212
rect 7184 2144 7229 2176
rect 7229 2144 7261 2176
rect 7261 2144 7306 2176
rect 7184 2108 7306 2144
rect 7184 2076 7229 2108
rect 7229 2076 7261 2108
rect 7261 2076 7306 2108
rect 7184 2042 7306 2076
rect 6923 1776 6963 1810
rect 6923 1744 6927 1776
rect 6927 1744 6959 1776
rect 6959 1744 6963 1776
rect 6923 1708 6963 1744
rect 6923 1676 6927 1708
rect 6927 1676 6959 1708
rect 6959 1676 6963 1708
rect 6923 1640 6963 1676
rect 6923 1608 6927 1640
rect 6927 1608 6959 1640
rect 6959 1608 6963 1640
rect 6923 1572 6963 1608
rect 6923 1540 6927 1572
rect 6927 1540 6959 1572
rect 6959 1540 6963 1572
rect 6923 1504 6963 1540
rect 6923 1472 6927 1504
rect 6927 1472 6959 1504
rect 6959 1472 6963 1504
rect 6923 1436 6963 1472
rect 6923 1404 6927 1436
rect 6927 1404 6959 1436
rect 6959 1404 6963 1436
rect 6923 1368 6963 1404
rect 6923 1336 6927 1368
rect 6927 1336 6959 1368
rect 6959 1336 6963 1368
rect 6923 1300 6963 1336
rect 6923 1268 6927 1300
rect 6927 1268 6959 1300
rect 6959 1268 6963 1300
rect 6923 1232 6963 1268
rect 6923 1200 6927 1232
rect 6927 1200 6959 1232
rect 6959 1200 6963 1232
rect 6923 1164 6963 1200
rect 6923 1132 6927 1164
rect 6927 1132 6959 1164
rect 6959 1132 6963 1164
rect 6923 1096 6963 1132
rect 6923 1064 6927 1096
rect 6927 1064 6959 1096
rect 6959 1064 6963 1096
rect 6923 1028 6963 1064
rect 6923 996 6927 1028
rect 6927 996 6959 1028
rect 6959 996 6963 1028
rect 6923 960 6963 996
rect 6923 928 6927 960
rect 6927 928 6959 960
rect 6959 928 6963 960
rect 6923 892 6963 928
rect 6923 860 6927 892
rect 6927 860 6959 892
rect 6959 860 6963 892
rect 6923 824 6963 860
rect 6923 792 6927 824
rect 6927 792 6959 824
rect 6959 792 6963 824
rect 6923 756 6963 792
rect 6923 724 6927 756
rect 6927 724 6959 756
rect 6959 724 6963 756
rect 6923 688 6963 724
rect 6923 656 6927 688
rect 6927 656 6959 688
rect 6959 656 6963 688
rect 6923 622 6963 656
rect 7527 3196 7567 3230
rect 7527 3164 7531 3196
rect 7531 3164 7563 3196
rect 7563 3164 7567 3196
rect 7527 3128 7567 3164
rect 7527 3096 7531 3128
rect 7531 3096 7563 3128
rect 7563 3096 7567 3128
rect 7527 3060 7567 3096
rect 7527 3028 7531 3060
rect 7531 3028 7563 3060
rect 7563 3028 7567 3060
rect 7527 2992 7567 3028
rect 7527 2960 7531 2992
rect 7531 2960 7563 2992
rect 7563 2960 7567 2992
rect 7527 2924 7567 2960
rect 7527 2892 7531 2924
rect 7531 2892 7563 2924
rect 7563 2892 7567 2924
rect 7527 2856 7567 2892
rect 7527 2824 7531 2856
rect 7531 2824 7563 2856
rect 7563 2824 7567 2856
rect 7527 2788 7567 2824
rect 7527 2756 7531 2788
rect 7531 2756 7563 2788
rect 7563 2756 7567 2788
rect 7527 2720 7567 2756
rect 7527 2688 7531 2720
rect 7531 2688 7563 2720
rect 7563 2688 7567 2720
rect 7527 2652 7567 2688
rect 7527 2620 7531 2652
rect 7531 2620 7563 2652
rect 7563 2620 7567 2652
rect 7527 2584 7567 2620
rect 7527 2552 7531 2584
rect 7531 2552 7563 2584
rect 7563 2552 7567 2584
rect 7527 2516 7567 2552
rect 7527 2484 7531 2516
rect 7531 2484 7563 2516
rect 7563 2484 7567 2516
rect 7527 2448 7567 2484
rect 7527 2416 7531 2448
rect 7531 2416 7563 2448
rect 7563 2416 7567 2448
rect 7527 2380 7567 2416
rect 7527 2348 7531 2380
rect 7531 2348 7563 2380
rect 7563 2348 7567 2380
rect 7527 2312 7567 2348
rect 7527 2280 7531 2312
rect 7531 2280 7563 2312
rect 7563 2280 7567 2312
rect 7527 2244 7567 2280
rect 7527 2212 7531 2244
rect 7531 2212 7563 2244
rect 7563 2212 7567 2244
rect 7527 2176 7567 2212
rect 7527 2144 7531 2176
rect 7531 2144 7563 2176
rect 7563 2144 7567 2176
rect 7527 2108 7567 2144
rect 7527 2076 7531 2108
rect 7531 2076 7563 2108
rect 7563 2076 7567 2108
rect 7527 2042 7567 2076
rect 7184 1776 7306 1810
rect 7184 1744 7229 1776
rect 7229 1744 7261 1776
rect 7261 1744 7306 1776
rect 7184 1708 7306 1744
rect 7184 1676 7229 1708
rect 7229 1676 7261 1708
rect 7261 1676 7306 1708
rect 7184 1640 7306 1676
rect 7184 1608 7229 1640
rect 7229 1608 7261 1640
rect 7261 1608 7306 1640
rect 7184 1572 7306 1608
rect 7184 1540 7229 1572
rect 7229 1540 7261 1572
rect 7261 1540 7306 1572
rect 7184 1504 7306 1540
rect 7184 1472 7229 1504
rect 7229 1472 7261 1504
rect 7261 1472 7306 1504
rect 7184 1436 7306 1472
rect 7184 1404 7229 1436
rect 7229 1404 7261 1436
rect 7261 1404 7306 1436
rect 7184 1368 7306 1404
rect 7184 1336 7229 1368
rect 7229 1336 7261 1368
rect 7261 1336 7306 1368
rect 7184 1300 7306 1336
rect 7184 1268 7229 1300
rect 7229 1268 7261 1300
rect 7261 1268 7306 1300
rect 7184 1232 7306 1268
rect 7184 1200 7229 1232
rect 7229 1200 7261 1232
rect 7261 1200 7306 1232
rect 7184 1164 7306 1200
rect 7184 1132 7229 1164
rect 7229 1132 7261 1164
rect 7261 1132 7306 1164
rect 7184 1096 7306 1132
rect 7184 1064 7229 1096
rect 7229 1064 7261 1096
rect 7261 1064 7306 1096
rect 7184 1028 7306 1064
rect 7184 996 7229 1028
rect 7229 996 7261 1028
rect 7261 996 7306 1028
rect 7184 960 7306 996
rect 7184 928 7229 960
rect 7229 928 7261 960
rect 7261 928 7306 960
rect 7184 892 7306 928
rect 7184 860 7229 892
rect 7229 860 7261 892
rect 7261 860 7306 892
rect 7184 824 7306 860
rect 7184 792 7229 824
rect 7229 792 7261 824
rect 7261 792 7306 824
rect 7184 756 7306 792
rect 7184 724 7229 756
rect 7229 724 7261 756
rect 7261 724 7306 756
rect 7184 688 7306 724
rect 7184 656 7229 688
rect 7229 656 7261 688
rect 7261 656 7306 688
rect 7184 622 7306 656
rect 7788 3196 7910 3230
rect 7788 3164 7833 3196
rect 7833 3164 7865 3196
rect 7865 3164 7910 3196
rect 7788 3128 7910 3164
rect 7788 3096 7833 3128
rect 7833 3096 7865 3128
rect 7865 3096 7910 3128
rect 7788 3060 7910 3096
rect 7788 3028 7833 3060
rect 7833 3028 7865 3060
rect 7865 3028 7910 3060
rect 7788 2992 7910 3028
rect 7788 2960 7833 2992
rect 7833 2960 7865 2992
rect 7865 2960 7910 2992
rect 7788 2924 7910 2960
rect 7788 2892 7833 2924
rect 7833 2892 7865 2924
rect 7865 2892 7910 2924
rect 7788 2856 7910 2892
rect 7788 2824 7833 2856
rect 7833 2824 7865 2856
rect 7865 2824 7910 2856
rect 7788 2788 7910 2824
rect 7788 2756 7833 2788
rect 7833 2756 7865 2788
rect 7865 2756 7910 2788
rect 7788 2720 7910 2756
rect 7788 2688 7833 2720
rect 7833 2688 7865 2720
rect 7865 2688 7910 2720
rect 7788 2652 7910 2688
rect 7788 2620 7833 2652
rect 7833 2620 7865 2652
rect 7865 2620 7910 2652
rect 7788 2584 7910 2620
rect 7788 2552 7833 2584
rect 7833 2552 7865 2584
rect 7865 2552 7910 2584
rect 7788 2516 7910 2552
rect 7788 2484 7833 2516
rect 7833 2484 7865 2516
rect 7865 2484 7910 2516
rect 7788 2448 7910 2484
rect 7788 2416 7833 2448
rect 7833 2416 7865 2448
rect 7865 2416 7910 2448
rect 7788 2380 7910 2416
rect 7788 2348 7833 2380
rect 7833 2348 7865 2380
rect 7865 2348 7910 2380
rect 7788 2312 7910 2348
rect 7788 2280 7833 2312
rect 7833 2280 7865 2312
rect 7865 2280 7910 2312
rect 7788 2244 7910 2280
rect 7788 2212 7833 2244
rect 7833 2212 7865 2244
rect 7865 2212 7910 2244
rect 7788 2176 7910 2212
rect 7788 2144 7833 2176
rect 7833 2144 7865 2176
rect 7865 2144 7910 2176
rect 7788 2108 7910 2144
rect 7788 2076 7833 2108
rect 7833 2076 7865 2108
rect 7865 2076 7910 2108
rect 7788 2042 7910 2076
rect 7527 1776 7567 1810
rect 7527 1744 7531 1776
rect 7531 1744 7563 1776
rect 7563 1744 7567 1776
rect 7527 1708 7567 1744
rect 7527 1676 7531 1708
rect 7531 1676 7563 1708
rect 7563 1676 7567 1708
rect 7527 1640 7567 1676
rect 7527 1608 7531 1640
rect 7531 1608 7563 1640
rect 7563 1608 7567 1640
rect 7527 1572 7567 1608
rect 7527 1540 7531 1572
rect 7531 1540 7563 1572
rect 7563 1540 7567 1572
rect 7527 1504 7567 1540
rect 7527 1472 7531 1504
rect 7531 1472 7563 1504
rect 7563 1472 7567 1504
rect 7527 1436 7567 1472
rect 7527 1404 7531 1436
rect 7531 1404 7563 1436
rect 7563 1404 7567 1436
rect 7527 1368 7567 1404
rect 7527 1336 7531 1368
rect 7531 1336 7563 1368
rect 7563 1336 7567 1368
rect 7527 1300 7567 1336
rect 7527 1268 7531 1300
rect 7531 1268 7563 1300
rect 7563 1268 7567 1300
rect 7527 1232 7567 1268
rect 7527 1200 7531 1232
rect 7531 1200 7563 1232
rect 7563 1200 7567 1232
rect 7527 1164 7567 1200
rect 7527 1132 7531 1164
rect 7531 1132 7563 1164
rect 7563 1132 7567 1164
rect 7527 1096 7567 1132
rect 7527 1064 7531 1096
rect 7531 1064 7563 1096
rect 7563 1064 7567 1096
rect 7527 1028 7567 1064
rect 7527 996 7531 1028
rect 7531 996 7563 1028
rect 7563 996 7567 1028
rect 7527 960 7567 996
rect 7527 928 7531 960
rect 7531 928 7563 960
rect 7563 928 7567 960
rect 7527 892 7567 928
rect 7527 860 7531 892
rect 7531 860 7563 892
rect 7563 860 7567 892
rect 7527 824 7567 860
rect 7527 792 7531 824
rect 7531 792 7563 824
rect 7563 792 7567 824
rect 7527 756 7567 792
rect 7527 724 7531 756
rect 7531 724 7563 756
rect 7563 724 7567 756
rect 7527 688 7567 724
rect 7527 656 7531 688
rect 7531 656 7563 688
rect 7563 656 7567 688
rect 7527 622 7567 656
rect 8131 3196 8171 3230
rect 8131 3164 8135 3196
rect 8135 3164 8167 3196
rect 8167 3164 8171 3196
rect 8131 3128 8171 3164
rect 8131 3096 8135 3128
rect 8135 3096 8167 3128
rect 8167 3096 8171 3128
rect 8131 3060 8171 3096
rect 8131 3028 8135 3060
rect 8135 3028 8167 3060
rect 8167 3028 8171 3060
rect 8131 2992 8171 3028
rect 8131 2960 8135 2992
rect 8135 2960 8167 2992
rect 8167 2960 8171 2992
rect 8131 2924 8171 2960
rect 8131 2892 8135 2924
rect 8135 2892 8167 2924
rect 8167 2892 8171 2924
rect 8131 2856 8171 2892
rect 8131 2824 8135 2856
rect 8135 2824 8167 2856
rect 8167 2824 8171 2856
rect 8131 2788 8171 2824
rect 8131 2756 8135 2788
rect 8135 2756 8167 2788
rect 8167 2756 8171 2788
rect 8131 2720 8171 2756
rect 8131 2688 8135 2720
rect 8135 2688 8167 2720
rect 8167 2688 8171 2720
rect 8131 2652 8171 2688
rect 8131 2620 8135 2652
rect 8135 2620 8167 2652
rect 8167 2620 8171 2652
rect 8131 2584 8171 2620
rect 8131 2552 8135 2584
rect 8135 2552 8167 2584
rect 8167 2552 8171 2584
rect 8131 2516 8171 2552
rect 8131 2484 8135 2516
rect 8135 2484 8167 2516
rect 8167 2484 8171 2516
rect 8131 2448 8171 2484
rect 8131 2416 8135 2448
rect 8135 2416 8167 2448
rect 8167 2416 8171 2448
rect 8131 2380 8171 2416
rect 8131 2348 8135 2380
rect 8135 2348 8167 2380
rect 8167 2348 8171 2380
rect 8131 2312 8171 2348
rect 8131 2280 8135 2312
rect 8135 2280 8167 2312
rect 8167 2280 8171 2312
rect 8131 2244 8171 2280
rect 8131 2212 8135 2244
rect 8135 2212 8167 2244
rect 8167 2212 8171 2244
rect 8131 2176 8171 2212
rect 8131 2144 8135 2176
rect 8135 2144 8167 2176
rect 8167 2144 8171 2176
rect 8131 2108 8171 2144
rect 8131 2076 8135 2108
rect 8135 2076 8167 2108
rect 8167 2076 8171 2108
rect 8131 2042 8171 2076
rect 7788 1776 7910 1810
rect 7788 1744 7833 1776
rect 7833 1744 7865 1776
rect 7865 1744 7910 1776
rect 7788 1708 7910 1744
rect 7788 1676 7833 1708
rect 7833 1676 7865 1708
rect 7865 1676 7910 1708
rect 7788 1640 7910 1676
rect 7788 1608 7833 1640
rect 7833 1608 7865 1640
rect 7865 1608 7910 1640
rect 7788 1572 7910 1608
rect 7788 1540 7833 1572
rect 7833 1540 7865 1572
rect 7865 1540 7910 1572
rect 7788 1504 7910 1540
rect 7788 1472 7833 1504
rect 7833 1472 7865 1504
rect 7865 1472 7910 1504
rect 7788 1436 7910 1472
rect 7788 1404 7833 1436
rect 7833 1404 7865 1436
rect 7865 1404 7910 1436
rect 7788 1368 7910 1404
rect 7788 1336 7833 1368
rect 7833 1336 7865 1368
rect 7865 1336 7910 1368
rect 7788 1300 7910 1336
rect 7788 1268 7833 1300
rect 7833 1268 7865 1300
rect 7865 1268 7910 1300
rect 7788 1232 7910 1268
rect 7788 1200 7833 1232
rect 7833 1200 7865 1232
rect 7865 1200 7910 1232
rect 7788 1164 7910 1200
rect 7788 1132 7833 1164
rect 7833 1132 7865 1164
rect 7865 1132 7910 1164
rect 7788 1096 7910 1132
rect 7788 1064 7833 1096
rect 7833 1064 7865 1096
rect 7865 1064 7910 1096
rect 7788 1028 7910 1064
rect 7788 996 7833 1028
rect 7833 996 7865 1028
rect 7865 996 7910 1028
rect 7788 960 7910 996
rect 7788 928 7833 960
rect 7833 928 7865 960
rect 7865 928 7910 960
rect 7788 892 7910 928
rect 7788 860 7833 892
rect 7833 860 7865 892
rect 7865 860 7910 892
rect 7788 824 7910 860
rect 7788 792 7833 824
rect 7833 792 7865 824
rect 7865 792 7910 824
rect 7788 756 7910 792
rect 7788 724 7833 756
rect 7833 724 7865 756
rect 7865 724 7910 756
rect 7788 688 7910 724
rect 7788 656 7833 688
rect 7833 656 7865 688
rect 7865 656 7910 688
rect 7788 622 7910 656
rect 8392 3196 8514 3230
rect 8392 3164 8437 3196
rect 8437 3164 8469 3196
rect 8469 3164 8514 3196
rect 8392 3128 8514 3164
rect 8392 3096 8437 3128
rect 8437 3096 8469 3128
rect 8469 3096 8514 3128
rect 8392 3060 8514 3096
rect 8392 3028 8437 3060
rect 8437 3028 8469 3060
rect 8469 3028 8514 3060
rect 8392 2992 8514 3028
rect 8392 2960 8437 2992
rect 8437 2960 8469 2992
rect 8469 2960 8514 2992
rect 8392 2924 8514 2960
rect 8392 2892 8437 2924
rect 8437 2892 8469 2924
rect 8469 2892 8514 2924
rect 8392 2856 8514 2892
rect 8392 2824 8437 2856
rect 8437 2824 8469 2856
rect 8469 2824 8514 2856
rect 8392 2788 8514 2824
rect 8392 2756 8437 2788
rect 8437 2756 8469 2788
rect 8469 2756 8514 2788
rect 8392 2720 8514 2756
rect 8392 2688 8437 2720
rect 8437 2688 8469 2720
rect 8469 2688 8514 2720
rect 8392 2652 8514 2688
rect 8392 2620 8437 2652
rect 8437 2620 8469 2652
rect 8469 2620 8514 2652
rect 8392 2584 8514 2620
rect 8392 2552 8437 2584
rect 8437 2552 8469 2584
rect 8469 2552 8514 2584
rect 8392 2516 8514 2552
rect 8392 2484 8437 2516
rect 8437 2484 8469 2516
rect 8469 2484 8514 2516
rect 8392 2448 8514 2484
rect 8392 2416 8437 2448
rect 8437 2416 8469 2448
rect 8469 2416 8514 2448
rect 8392 2380 8514 2416
rect 8392 2348 8437 2380
rect 8437 2348 8469 2380
rect 8469 2348 8514 2380
rect 8392 2312 8514 2348
rect 8392 2280 8437 2312
rect 8437 2280 8469 2312
rect 8469 2280 8514 2312
rect 8392 2244 8514 2280
rect 8392 2212 8437 2244
rect 8437 2212 8469 2244
rect 8469 2212 8514 2244
rect 8392 2176 8514 2212
rect 8392 2144 8437 2176
rect 8437 2144 8469 2176
rect 8469 2144 8514 2176
rect 8392 2108 8514 2144
rect 8392 2076 8437 2108
rect 8437 2076 8469 2108
rect 8469 2076 8514 2108
rect 8392 2042 8514 2076
rect 8131 1776 8171 1810
rect 8131 1744 8135 1776
rect 8135 1744 8167 1776
rect 8167 1744 8171 1776
rect 8131 1708 8171 1744
rect 8131 1676 8135 1708
rect 8135 1676 8167 1708
rect 8167 1676 8171 1708
rect 8131 1640 8171 1676
rect 8131 1608 8135 1640
rect 8135 1608 8167 1640
rect 8167 1608 8171 1640
rect 8131 1572 8171 1608
rect 8131 1540 8135 1572
rect 8135 1540 8167 1572
rect 8167 1540 8171 1572
rect 8131 1504 8171 1540
rect 8131 1472 8135 1504
rect 8135 1472 8167 1504
rect 8167 1472 8171 1504
rect 8131 1436 8171 1472
rect 8131 1404 8135 1436
rect 8135 1404 8167 1436
rect 8167 1404 8171 1436
rect 8131 1368 8171 1404
rect 8131 1336 8135 1368
rect 8135 1336 8167 1368
rect 8167 1336 8171 1368
rect 8131 1300 8171 1336
rect 8131 1268 8135 1300
rect 8135 1268 8167 1300
rect 8167 1268 8171 1300
rect 8131 1232 8171 1268
rect 8131 1200 8135 1232
rect 8135 1200 8167 1232
rect 8167 1200 8171 1232
rect 8131 1164 8171 1200
rect 8131 1132 8135 1164
rect 8135 1132 8167 1164
rect 8167 1132 8171 1164
rect 8131 1096 8171 1132
rect 8131 1064 8135 1096
rect 8135 1064 8167 1096
rect 8167 1064 8171 1096
rect 8131 1028 8171 1064
rect 8131 996 8135 1028
rect 8135 996 8167 1028
rect 8167 996 8171 1028
rect 8131 960 8171 996
rect 8131 928 8135 960
rect 8135 928 8167 960
rect 8167 928 8171 960
rect 8131 892 8171 928
rect 8131 860 8135 892
rect 8135 860 8167 892
rect 8167 860 8171 892
rect 8131 824 8171 860
rect 8131 792 8135 824
rect 8135 792 8167 824
rect 8167 792 8171 824
rect 8131 756 8171 792
rect 8131 724 8135 756
rect 8135 724 8167 756
rect 8167 724 8171 756
rect 8131 688 8171 724
rect 8131 656 8135 688
rect 8135 656 8167 688
rect 8167 656 8171 688
rect 8131 622 8171 656
rect 8735 3196 8775 3230
rect 8735 3164 8739 3196
rect 8739 3164 8771 3196
rect 8771 3164 8775 3196
rect 8735 3128 8775 3164
rect 8735 3096 8739 3128
rect 8739 3096 8771 3128
rect 8771 3096 8775 3128
rect 8735 3060 8775 3096
rect 8735 3028 8739 3060
rect 8739 3028 8771 3060
rect 8771 3028 8775 3060
rect 8735 2992 8775 3028
rect 8735 2960 8739 2992
rect 8739 2960 8771 2992
rect 8771 2960 8775 2992
rect 8735 2924 8775 2960
rect 8735 2892 8739 2924
rect 8739 2892 8771 2924
rect 8771 2892 8775 2924
rect 8735 2856 8775 2892
rect 8735 2824 8739 2856
rect 8739 2824 8771 2856
rect 8771 2824 8775 2856
rect 8735 2788 8775 2824
rect 8735 2756 8739 2788
rect 8739 2756 8771 2788
rect 8771 2756 8775 2788
rect 8735 2720 8775 2756
rect 8735 2688 8739 2720
rect 8739 2688 8771 2720
rect 8771 2688 8775 2720
rect 8735 2652 8775 2688
rect 8735 2620 8739 2652
rect 8739 2620 8771 2652
rect 8771 2620 8775 2652
rect 8735 2584 8775 2620
rect 8735 2552 8739 2584
rect 8739 2552 8771 2584
rect 8771 2552 8775 2584
rect 8735 2516 8775 2552
rect 8735 2484 8739 2516
rect 8739 2484 8771 2516
rect 8771 2484 8775 2516
rect 8735 2448 8775 2484
rect 8735 2416 8739 2448
rect 8739 2416 8771 2448
rect 8771 2416 8775 2448
rect 8735 2380 8775 2416
rect 8735 2348 8739 2380
rect 8739 2348 8771 2380
rect 8771 2348 8775 2380
rect 8735 2312 8775 2348
rect 8735 2280 8739 2312
rect 8739 2280 8771 2312
rect 8771 2280 8775 2312
rect 8735 2244 8775 2280
rect 8735 2212 8739 2244
rect 8739 2212 8771 2244
rect 8771 2212 8775 2244
rect 8735 2176 8775 2212
rect 8735 2144 8739 2176
rect 8739 2144 8771 2176
rect 8771 2144 8775 2176
rect 8735 2108 8775 2144
rect 8735 2076 8739 2108
rect 8739 2076 8771 2108
rect 8771 2076 8775 2108
rect 8735 2042 8775 2076
rect 8392 1776 8514 1810
rect 8392 1744 8437 1776
rect 8437 1744 8469 1776
rect 8469 1744 8514 1776
rect 8392 1708 8514 1744
rect 8392 1676 8437 1708
rect 8437 1676 8469 1708
rect 8469 1676 8514 1708
rect 8392 1640 8514 1676
rect 8392 1608 8437 1640
rect 8437 1608 8469 1640
rect 8469 1608 8514 1640
rect 8392 1572 8514 1608
rect 8392 1540 8437 1572
rect 8437 1540 8469 1572
rect 8469 1540 8514 1572
rect 8392 1504 8514 1540
rect 8392 1472 8437 1504
rect 8437 1472 8469 1504
rect 8469 1472 8514 1504
rect 8392 1436 8514 1472
rect 8392 1404 8437 1436
rect 8437 1404 8469 1436
rect 8469 1404 8514 1436
rect 8392 1368 8514 1404
rect 8392 1336 8437 1368
rect 8437 1336 8469 1368
rect 8469 1336 8514 1368
rect 8392 1300 8514 1336
rect 8392 1268 8437 1300
rect 8437 1268 8469 1300
rect 8469 1268 8514 1300
rect 8392 1232 8514 1268
rect 8392 1200 8437 1232
rect 8437 1200 8469 1232
rect 8469 1200 8514 1232
rect 8392 1164 8514 1200
rect 8392 1132 8437 1164
rect 8437 1132 8469 1164
rect 8469 1132 8514 1164
rect 8392 1096 8514 1132
rect 8392 1064 8437 1096
rect 8437 1064 8469 1096
rect 8469 1064 8514 1096
rect 8392 1028 8514 1064
rect 8392 996 8437 1028
rect 8437 996 8469 1028
rect 8469 996 8514 1028
rect 8392 960 8514 996
rect 8392 928 8437 960
rect 8437 928 8469 960
rect 8469 928 8514 960
rect 8392 892 8514 928
rect 8392 860 8437 892
rect 8437 860 8469 892
rect 8469 860 8514 892
rect 8392 824 8514 860
rect 8392 792 8437 824
rect 8437 792 8469 824
rect 8469 792 8514 824
rect 8392 756 8514 792
rect 8392 724 8437 756
rect 8437 724 8469 756
rect 8469 724 8514 756
rect 8392 688 8514 724
rect 8392 656 8437 688
rect 8437 656 8469 688
rect 8469 656 8514 688
rect 8392 622 8514 656
rect 8996 3196 9118 3230
rect 8996 3164 9041 3196
rect 9041 3164 9073 3196
rect 9073 3164 9118 3196
rect 8996 3128 9118 3164
rect 8996 3096 9041 3128
rect 9041 3096 9073 3128
rect 9073 3096 9118 3128
rect 8996 3060 9118 3096
rect 8996 3028 9041 3060
rect 9041 3028 9073 3060
rect 9073 3028 9118 3060
rect 8996 2992 9118 3028
rect 8996 2960 9041 2992
rect 9041 2960 9073 2992
rect 9073 2960 9118 2992
rect 8996 2924 9118 2960
rect 8996 2892 9041 2924
rect 9041 2892 9073 2924
rect 9073 2892 9118 2924
rect 8996 2856 9118 2892
rect 8996 2824 9041 2856
rect 9041 2824 9073 2856
rect 9073 2824 9118 2856
rect 8996 2788 9118 2824
rect 8996 2756 9041 2788
rect 9041 2756 9073 2788
rect 9073 2756 9118 2788
rect 8996 2720 9118 2756
rect 8996 2688 9041 2720
rect 9041 2688 9073 2720
rect 9073 2688 9118 2720
rect 8996 2652 9118 2688
rect 8996 2620 9041 2652
rect 9041 2620 9073 2652
rect 9073 2620 9118 2652
rect 8996 2584 9118 2620
rect 8996 2552 9041 2584
rect 9041 2552 9073 2584
rect 9073 2552 9118 2584
rect 8996 2516 9118 2552
rect 8996 2484 9041 2516
rect 9041 2484 9073 2516
rect 9073 2484 9118 2516
rect 8996 2448 9118 2484
rect 8996 2416 9041 2448
rect 9041 2416 9073 2448
rect 9073 2416 9118 2448
rect 8996 2380 9118 2416
rect 8996 2348 9041 2380
rect 9041 2348 9073 2380
rect 9073 2348 9118 2380
rect 8996 2312 9118 2348
rect 8996 2280 9041 2312
rect 9041 2280 9073 2312
rect 9073 2280 9118 2312
rect 8996 2244 9118 2280
rect 8996 2212 9041 2244
rect 9041 2212 9073 2244
rect 9073 2212 9118 2244
rect 8996 2176 9118 2212
rect 8996 2144 9041 2176
rect 9041 2144 9073 2176
rect 9073 2144 9118 2176
rect 8996 2108 9118 2144
rect 8996 2076 9041 2108
rect 9041 2076 9073 2108
rect 9073 2076 9118 2108
rect 8996 2042 9118 2076
rect 8735 1776 8775 1810
rect 8735 1744 8739 1776
rect 8739 1744 8771 1776
rect 8771 1744 8775 1776
rect 8735 1708 8775 1744
rect 8735 1676 8739 1708
rect 8739 1676 8771 1708
rect 8771 1676 8775 1708
rect 8735 1640 8775 1676
rect 8735 1608 8739 1640
rect 8739 1608 8771 1640
rect 8771 1608 8775 1640
rect 8735 1572 8775 1608
rect 8735 1540 8739 1572
rect 8739 1540 8771 1572
rect 8771 1540 8775 1572
rect 8735 1504 8775 1540
rect 8735 1472 8739 1504
rect 8739 1472 8771 1504
rect 8771 1472 8775 1504
rect 8735 1436 8775 1472
rect 8735 1404 8739 1436
rect 8739 1404 8771 1436
rect 8771 1404 8775 1436
rect 8735 1368 8775 1404
rect 8735 1336 8739 1368
rect 8739 1336 8771 1368
rect 8771 1336 8775 1368
rect 8735 1300 8775 1336
rect 8735 1268 8739 1300
rect 8739 1268 8771 1300
rect 8771 1268 8775 1300
rect 8735 1232 8775 1268
rect 8735 1200 8739 1232
rect 8739 1200 8771 1232
rect 8771 1200 8775 1232
rect 8735 1164 8775 1200
rect 8735 1132 8739 1164
rect 8739 1132 8771 1164
rect 8771 1132 8775 1164
rect 8735 1096 8775 1132
rect 8735 1064 8739 1096
rect 8739 1064 8771 1096
rect 8771 1064 8775 1096
rect 8735 1028 8775 1064
rect 8735 996 8739 1028
rect 8739 996 8771 1028
rect 8771 996 8775 1028
rect 8735 960 8775 996
rect 8735 928 8739 960
rect 8739 928 8771 960
rect 8771 928 8775 960
rect 8735 892 8775 928
rect 8735 860 8739 892
rect 8739 860 8771 892
rect 8771 860 8775 892
rect 8735 824 8775 860
rect 8735 792 8739 824
rect 8739 792 8771 824
rect 8771 792 8775 824
rect 8735 756 8775 792
rect 8735 724 8739 756
rect 8739 724 8771 756
rect 8771 724 8775 756
rect 8735 688 8775 724
rect 8735 656 8739 688
rect 8739 656 8771 688
rect 8771 656 8775 688
rect 8735 622 8775 656
rect 9339 3196 9379 3230
rect 9339 3164 9343 3196
rect 9343 3164 9375 3196
rect 9375 3164 9379 3196
rect 9339 3128 9379 3164
rect 9339 3096 9343 3128
rect 9343 3096 9375 3128
rect 9375 3096 9379 3128
rect 9339 3060 9379 3096
rect 9339 3028 9343 3060
rect 9343 3028 9375 3060
rect 9375 3028 9379 3060
rect 9339 2992 9379 3028
rect 9339 2960 9343 2992
rect 9343 2960 9375 2992
rect 9375 2960 9379 2992
rect 9339 2924 9379 2960
rect 9339 2892 9343 2924
rect 9343 2892 9375 2924
rect 9375 2892 9379 2924
rect 9339 2856 9379 2892
rect 9339 2824 9343 2856
rect 9343 2824 9375 2856
rect 9375 2824 9379 2856
rect 9339 2788 9379 2824
rect 9339 2756 9343 2788
rect 9343 2756 9375 2788
rect 9375 2756 9379 2788
rect 9339 2720 9379 2756
rect 9339 2688 9343 2720
rect 9343 2688 9375 2720
rect 9375 2688 9379 2720
rect 9339 2652 9379 2688
rect 9339 2620 9343 2652
rect 9343 2620 9375 2652
rect 9375 2620 9379 2652
rect 9339 2584 9379 2620
rect 9339 2552 9343 2584
rect 9343 2552 9375 2584
rect 9375 2552 9379 2584
rect 9339 2516 9379 2552
rect 9339 2484 9343 2516
rect 9343 2484 9375 2516
rect 9375 2484 9379 2516
rect 9339 2448 9379 2484
rect 9339 2416 9343 2448
rect 9343 2416 9375 2448
rect 9375 2416 9379 2448
rect 9339 2380 9379 2416
rect 9339 2348 9343 2380
rect 9343 2348 9375 2380
rect 9375 2348 9379 2380
rect 9339 2312 9379 2348
rect 9339 2280 9343 2312
rect 9343 2280 9375 2312
rect 9375 2280 9379 2312
rect 9339 2244 9379 2280
rect 9339 2212 9343 2244
rect 9343 2212 9375 2244
rect 9375 2212 9379 2244
rect 9339 2176 9379 2212
rect 9339 2144 9343 2176
rect 9343 2144 9375 2176
rect 9375 2144 9379 2176
rect 9339 2108 9379 2144
rect 9339 2076 9343 2108
rect 9343 2076 9375 2108
rect 9375 2076 9379 2108
rect 9339 2042 9379 2076
rect 8996 1776 9118 1810
rect 8996 1744 9041 1776
rect 9041 1744 9073 1776
rect 9073 1744 9118 1776
rect 8996 1708 9118 1744
rect 8996 1676 9041 1708
rect 9041 1676 9073 1708
rect 9073 1676 9118 1708
rect 8996 1640 9118 1676
rect 8996 1608 9041 1640
rect 9041 1608 9073 1640
rect 9073 1608 9118 1640
rect 8996 1572 9118 1608
rect 8996 1540 9041 1572
rect 9041 1540 9073 1572
rect 9073 1540 9118 1572
rect 8996 1504 9118 1540
rect 8996 1472 9041 1504
rect 9041 1472 9073 1504
rect 9073 1472 9118 1504
rect 8996 1436 9118 1472
rect 8996 1404 9041 1436
rect 9041 1404 9073 1436
rect 9073 1404 9118 1436
rect 8996 1368 9118 1404
rect 8996 1336 9041 1368
rect 9041 1336 9073 1368
rect 9073 1336 9118 1368
rect 8996 1300 9118 1336
rect 8996 1268 9041 1300
rect 9041 1268 9073 1300
rect 9073 1268 9118 1300
rect 8996 1232 9118 1268
rect 8996 1200 9041 1232
rect 9041 1200 9073 1232
rect 9073 1200 9118 1232
rect 8996 1164 9118 1200
rect 8996 1132 9041 1164
rect 9041 1132 9073 1164
rect 9073 1132 9118 1164
rect 8996 1096 9118 1132
rect 8996 1064 9041 1096
rect 9041 1064 9073 1096
rect 9073 1064 9118 1096
rect 8996 1028 9118 1064
rect 8996 996 9041 1028
rect 9041 996 9073 1028
rect 9073 996 9118 1028
rect 8996 960 9118 996
rect 8996 928 9041 960
rect 9041 928 9073 960
rect 9073 928 9118 960
rect 8996 892 9118 928
rect 8996 860 9041 892
rect 9041 860 9073 892
rect 9073 860 9118 892
rect 8996 824 9118 860
rect 8996 792 9041 824
rect 9041 792 9073 824
rect 9073 792 9118 824
rect 8996 756 9118 792
rect 8996 724 9041 756
rect 9041 724 9073 756
rect 9073 724 9118 756
rect 8996 688 9118 724
rect 8996 656 9041 688
rect 9041 656 9073 688
rect 9073 656 9118 688
rect 8996 622 9118 656
rect 9600 3196 9722 3230
rect 9600 3164 9645 3196
rect 9645 3164 9677 3196
rect 9677 3164 9722 3196
rect 9600 3128 9722 3164
rect 9600 3096 9645 3128
rect 9645 3096 9677 3128
rect 9677 3096 9722 3128
rect 9600 3060 9722 3096
rect 9600 3028 9645 3060
rect 9645 3028 9677 3060
rect 9677 3028 9722 3060
rect 9600 2992 9722 3028
rect 9600 2960 9645 2992
rect 9645 2960 9677 2992
rect 9677 2960 9722 2992
rect 9600 2924 9722 2960
rect 9600 2892 9645 2924
rect 9645 2892 9677 2924
rect 9677 2892 9722 2924
rect 9600 2856 9722 2892
rect 9600 2824 9645 2856
rect 9645 2824 9677 2856
rect 9677 2824 9722 2856
rect 9600 2788 9722 2824
rect 9600 2756 9645 2788
rect 9645 2756 9677 2788
rect 9677 2756 9722 2788
rect 9600 2720 9722 2756
rect 9600 2688 9645 2720
rect 9645 2688 9677 2720
rect 9677 2688 9722 2720
rect 9600 2652 9722 2688
rect 9600 2620 9645 2652
rect 9645 2620 9677 2652
rect 9677 2620 9722 2652
rect 9600 2584 9722 2620
rect 9600 2552 9645 2584
rect 9645 2552 9677 2584
rect 9677 2552 9722 2584
rect 9600 2516 9722 2552
rect 9600 2484 9645 2516
rect 9645 2484 9677 2516
rect 9677 2484 9722 2516
rect 9600 2448 9722 2484
rect 9600 2416 9645 2448
rect 9645 2416 9677 2448
rect 9677 2416 9722 2448
rect 9600 2380 9722 2416
rect 9600 2348 9645 2380
rect 9645 2348 9677 2380
rect 9677 2348 9722 2380
rect 9600 2312 9722 2348
rect 9600 2280 9645 2312
rect 9645 2280 9677 2312
rect 9677 2280 9722 2312
rect 9600 2244 9722 2280
rect 9600 2212 9645 2244
rect 9645 2212 9677 2244
rect 9677 2212 9722 2244
rect 9600 2176 9722 2212
rect 9600 2144 9645 2176
rect 9645 2144 9677 2176
rect 9677 2144 9722 2176
rect 9600 2108 9722 2144
rect 9600 2076 9645 2108
rect 9645 2076 9677 2108
rect 9677 2076 9722 2108
rect 9600 2042 9722 2076
rect 9339 1776 9379 1810
rect 9339 1744 9343 1776
rect 9343 1744 9375 1776
rect 9375 1744 9379 1776
rect 9339 1708 9379 1744
rect 9339 1676 9343 1708
rect 9343 1676 9375 1708
rect 9375 1676 9379 1708
rect 9339 1640 9379 1676
rect 9339 1608 9343 1640
rect 9343 1608 9375 1640
rect 9375 1608 9379 1640
rect 9339 1572 9379 1608
rect 9339 1540 9343 1572
rect 9343 1540 9375 1572
rect 9375 1540 9379 1572
rect 9339 1504 9379 1540
rect 9339 1472 9343 1504
rect 9343 1472 9375 1504
rect 9375 1472 9379 1504
rect 9339 1436 9379 1472
rect 9339 1404 9343 1436
rect 9343 1404 9375 1436
rect 9375 1404 9379 1436
rect 9339 1368 9379 1404
rect 9339 1336 9343 1368
rect 9343 1336 9375 1368
rect 9375 1336 9379 1368
rect 9339 1300 9379 1336
rect 9339 1268 9343 1300
rect 9343 1268 9375 1300
rect 9375 1268 9379 1300
rect 9339 1232 9379 1268
rect 9339 1200 9343 1232
rect 9343 1200 9375 1232
rect 9375 1200 9379 1232
rect 9339 1164 9379 1200
rect 9339 1132 9343 1164
rect 9343 1132 9375 1164
rect 9375 1132 9379 1164
rect 9339 1096 9379 1132
rect 9339 1064 9343 1096
rect 9343 1064 9375 1096
rect 9375 1064 9379 1096
rect 9339 1028 9379 1064
rect 9339 996 9343 1028
rect 9343 996 9375 1028
rect 9375 996 9379 1028
rect 9339 960 9379 996
rect 9339 928 9343 960
rect 9343 928 9375 960
rect 9375 928 9379 960
rect 9339 892 9379 928
rect 9339 860 9343 892
rect 9343 860 9375 892
rect 9375 860 9379 892
rect 9339 824 9379 860
rect 9339 792 9343 824
rect 9343 792 9375 824
rect 9375 792 9379 824
rect 9339 756 9379 792
rect 9339 724 9343 756
rect 9343 724 9375 756
rect 9375 724 9379 756
rect 9339 688 9379 724
rect 9339 656 9343 688
rect 9343 656 9375 688
rect 9375 656 9379 688
rect 9339 622 9379 656
rect 9943 3196 9983 3230
rect 9943 3164 9947 3196
rect 9947 3164 9979 3196
rect 9979 3164 9983 3196
rect 9943 3128 9983 3164
rect 9943 3096 9947 3128
rect 9947 3096 9979 3128
rect 9979 3096 9983 3128
rect 9943 3060 9983 3096
rect 9943 3028 9947 3060
rect 9947 3028 9979 3060
rect 9979 3028 9983 3060
rect 9943 2992 9983 3028
rect 9943 2960 9947 2992
rect 9947 2960 9979 2992
rect 9979 2960 9983 2992
rect 9943 2924 9983 2960
rect 9943 2892 9947 2924
rect 9947 2892 9979 2924
rect 9979 2892 9983 2924
rect 9943 2856 9983 2892
rect 9943 2824 9947 2856
rect 9947 2824 9979 2856
rect 9979 2824 9983 2856
rect 9943 2788 9983 2824
rect 9943 2756 9947 2788
rect 9947 2756 9979 2788
rect 9979 2756 9983 2788
rect 9943 2720 9983 2756
rect 9943 2688 9947 2720
rect 9947 2688 9979 2720
rect 9979 2688 9983 2720
rect 9943 2652 9983 2688
rect 9943 2620 9947 2652
rect 9947 2620 9979 2652
rect 9979 2620 9983 2652
rect 9943 2584 9983 2620
rect 9943 2552 9947 2584
rect 9947 2552 9979 2584
rect 9979 2552 9983 2584
rect 9943 2516 9983 2552
rect 9943 2484 9947 2516
rect 9947 2484 9979 2516
rect 9979 2484 9983 2516
rect 9943 2448 9983 2484
rect 9943 2416 9947 2448
rect 9947 2416 9979 2448
rect 9979 2416 9983 2448
rect 9943 2380 9983 2416
rect 9943 2348 9947 2380
rect 9947 2348 9979 2380
rect 9979 2348 9983 2380
rect 9943 2312 9983 2348
rect 9943 2280 9947 2312
rect 9947 2280 9979 2312
rect 9979 2280 9983 2312
rect 9943 2244 9983 2280
rect 9943 2212 9947 2244
rect 9947 2212 9979 2244
rect 9979 2212 9983 2244
rect 9943 2176 9983 2212
rect 9943 2144 9947 2176
rect 9947 2144 9979 2176
rect 9979 2144 9983 2176
rect 9943 2108 9983 2144
rect 9943 2076 9947 2108
rect 9947 2076 9979 2108
rect 9979 2076 9983 2108
rect 9943 2042 9983 2076
rect 9600 1776 9722 1810
rect 9600 1744 9645 1776
rect 9645 1744 9677 1776
rect 9677 1744 9722 1776
rect 9600 1708 9722 1744
rect 9600 1676 9645 1708
rect 9645 1676 9677 1708
rect 9677 1676 9722 1708
rect 9600 1640 9722 1676
rect 9600 1608 9645 1640
rect 9645 1608 9677 1640
rect 9677 1608 9722 1640
rect 9600 1572 9722 1608
rect 9600 1540 9645 1572
rect 9645 1540 9677 1572
rect 9677 1540 9722 1572
rect 9600 1504 9722 1540
rect 9600 1472 9645 1504
rect 9645 1472 9677 1504
rect 9677 1472 9722 1504
rect 9600 1436 9722 1472
rect 9600 1404 9645 1436
rect 9645 1404 9677 1436
rect 9677 1404 9722 1436
rect 9600 1368 9722 1404
rect 9600 1336 9645 1368
rect 9645 1336 9677 1368
rect 9677 1336 9722 1368
rect 9600 1300 9722 1336
rect 9600 1268 9645 1300
rect 9645 1268 9677 1300
rect 9677 1268 9722 1300
rect 9600 1232 9722 1268
rect 9600 1200 9645 1232
rect 9645 1200 9677 1232
rect 9677 1200 9722 1232
rect 9600 1164 9722 1200
rect 9600 1132 9645 1164
rect 9645 1132 9677 1164
rect 9677 1132 9722 1164
rect 9600 1096 9722 1132
rect 9600 1064 9645 1096
rect 9645 1064 9677 1096
rect 9677 1064 9722 1096
rect 9600 1028 9722 1064
rect 9600 996 9645 1028
rect 9645 996 9677 1028
rect 9677 996 9722 1028
rect 9600 960 9722 996
rect 9600 928 9645 960
rect 9645 928 9677 960
rect 9677 928 9722 960
rect 9600 892 9722 928
rect 9600 860 9645 892
rect 9645 860 9677 892
rect 9677 860 9722 892
rect 9600 824 9722 860
rect 9600 792 9645 824
rect 9645 792 9677 824
rect 9677 792 9722 824
rect 9600 756 9722 792
rect 9600 724 9645 756
rect 9645 724 9677 756
rect 9677 724 9722 756
rect 9600 688 9722 724
rect 9600 656 9645 688
rect 9645 656 9677 688
rect 9677 656 9722 688
rect 9600 622 9722 656
rect 10204 3196 10326 3230
rect 10204 3164 10249 3196
rect 10249 3164 10281 3196
rect 10281 3164 10326 3196
rect 10204 3128 10326 3164
rect 10204 3096 10249 3128
rect 10249 3096 10281 3128
rect 10281 3096 10326 3128
rect 10204 3060 10326 3096
rect 10204 3028 10249 3060
rect 10249 3028 10281 3060
rect 10281 3028 10326 3060
rect 10204 2992 10326 3028
rect 10204 2960 10249 2992
rect 10249 2960 10281 2992
rect 10281 2960 10326 2992
rect 10204 2924 10326 2960
rect 10204 2892 10249 2924
rect 10249 2892 10281 2924
rect 10281 2892 10326 2924
rect 10204 2856 10326 2892
rect 10204 2824 10249 2856
rect 10249 2824 10281 2856
rect 10281 2824 10326 2856
rect 10204 2788 10326 2824
rect 10204 2756 10249 2788
rect 10249 2756 10281 2788
rect 10281 2756 10326 2788
rect 10204 2720 10326 2756
rect 10204 2688 10249 2720
rect 10249 2688 10281 2720
rect 10281 2688 10326 2720
rect 10204 2652 10326 2688
rect 10204 2620 10249 2652
rect 10249 2620 10281 2652
rect 10281 2620 10326 2652
rect 10204 2584 10326 2620
rect 10204 2552 10249 2584
rect 10249 2552 10281 2584
rect 10281 2552 10326 2584
rect 10204 2516 10326 2552
rect 10204 2484 10249 2516
rect 10249 2484 10281 2516
rect 10281 2484 10326 2516
rect 10204 2448 10326 2484
rect 10204 2416 10249 2448
rect 10249 2416 10281 2448
rect 10281 2416 10326 2448
rect 10204 2380 10326 2416
rect 10204 2348 10249 2380
rect 10249 2348 10281 2380
rect 10281 2348 10326 2380
rect 10204 2312 10326 2348
rect 10204 2280 10249 2312
rect 10249 2280 10281 2312
rect 10281 2280 10326 2312
rect 10204 2244 10326 2280
rect 10204 2212 10249 2244
rect 10249 2212 10281 2244
rect 10281 2212 10326 2244
rect 10204 2176 10326 2212
rect 10204 2144 10249 2176
rect 10249 2144 10281 2176
rect 10281 2144 10326 2176
rect 10204 2108 10326 2144
rect 10204 2076 10249 2108
rect 10249 2076 10281 2108
rect 10281 2076 10326 2108
rect 10204 2042 10326 2076
rect 9943 1776 9983 1810
rect 9943 1744 9947 1776
rect 9947 1744 9979 1776
rect 9979 1744 9983 1776
rect 9943 1708 9983 1744
rect 9943 1676 9947 1708
rect 9947 1676 9979 1708
rect 9979 1676 9983 1708
rect 9943 1640 9983 1676
rect 9943 1608 9947 1640
rect 9947 1608 9979 1640
rect 9979 1608 9983 1640
rect 9943 1572 9983 1608
rect 9943 1540 9947 1572
rect 9947 1540 9979 1572
rect 9979 1540 9983 1572
rect 9943 1504 9983 1540
rect 9943 1472 9947 1504
rect 9947 1472 9979 1504
rect 9979 1472 9983 1504
rect 9943 1436 9983 1472
rect 9943 1404 9947 1436
rect 9947 1404 9979 1436
rect 9979 1404 9983 1436
rect 9943 1368 9983 1404
rect 9943 1336 9947 1368
rect 9947 1336 9979 1368
rect 9979 1336 9983 1368
rect 9943 1300 9983 1336
rect 9943 1268 9947 1300
rect 9947 1268 9979 1300
rect 9979 1268 9983 1300
rect 9943 1232 9983 1268
rect 9943 1200 9947 1232
rect 9947 1200 9979 1232
rect 9979 1200 9983 1232
rect 9943 1164 9983 1200
rect 9943 1132 9947 1164
rect 9947 1132 9979 1164
rect 9979 1132 9983 1164
rect 9943 1096 9983 1132
rect 9943 1064 9947 1096
rect 9947 1064 9979 1096
rect 9979 1064 9983 1096
rect 9943 1028 9983 1064
rect 9943 996 9947 1028
rect 9947 996 9979 1028
rect 9979 996 9983 1028
rect 9943 960 9983 996
rect 9943 928 9947 960
rect 9947 928 9979 960
rect 9979 928 9983 960
rect 9943 892 9983 928
rect 9943 860 9947 892
rect 9947 860 9979 892
rect 9979 860 9983 892
rect 9943 824 9983 860
rect 9943 792 9947 824
rect 9947 792 9979 824
rect 9979 792 9983 824
rect 9943 756 9983 792
rect 9943 724 9947 756
rect 9947 724 9979 756
rect 9979 724 9983 756
rect 9943 688 9983 724
rect 9943 656 9947 688
rect 9947 656 9979 688
rect 9979 656 9983 688
rect 9943 622 9983 656
rect 10204 1776 10326 1810
rect 10204 1744 10249 1776
rect 10249 1744 10281 1776
rect 10281 1744 10326 1776
rect 10204 1708 10326 1744
rect 10204 1676 10249 1708
rect 10249 1676 10281 1708
rect 10281 1676 10326 1708
rect 10204 1640 10326 1676
rect 10204 1608 10249 1640
rect 10249 1608 10281 1640
rect 10281 1608 10326 1640
rect 10204 1572 10326 1608
rect 10204 1540 10249 1572
rect 10249 1540 10281 1572
rect 10281 1540 10326 1572
rect 10204 1504 10326 1540
rect 10204 1472 10249 1504
rect 10249 1472 10281 1504
rect 10281 1472 10326 1504
rect 10204 1436 10326 1472
rect 10204 1404 10249 1436
rect 10249 1404 10281 1436
rect 10281 1404 10326 1436
rect 10204 1368 10326 1404
rect 10204 1336 10249 1368
rect 10249 1336 10281 1368
rect 10281 1336 10326 1368
rect 10204 1300 10326 1336
rect 10204 1268 10249 1300
rect 10249 1268 10281 1300
rect 10281 1268 10326 1300
rect 10204 1232 10326 1268
rect 10204 1200 10249 1232
rect 10249 1200 10281 1232
rect 10281 1200 10326 1232
rect 10204 1164 10326 1200
rect 10204 1132 10249 1164
rect 10249 1132 10281 1164
rect 10281 1132 10326 1164
rect 10204 1096 10326 1132
rect 10204 1064 10249 1096
rect 10249 1064 10281 1096
rect 10281 1064 10326 1096
rect 10204 1028 10326 1064
rect 10204 996 10249 1028
rect 10249 996 10281 1028
rect 10281 996 10326 1028
rect 10204 960 10326 996
rect 10204 928 10249 960
rect 10249 928 10281 960
rect 10281 928 10326 960
rect 10204 892 10326 928
rect 10204 860 10249 892
rect 10249 860 10281 892
rect 10281 860 10326 892
rect 10204 824 10326 860
rect 10204 792 10249 824
rect 10249 792 10281 824
rect 10281 792 10326 824
rect 10204 756 10326 792
rect 10204 724 10249 756
rect 10249 724 10281 756
rect 10281 724 10326 756
rect 10204 688 10326 724
rect 10204 656 10249 688
rect 10249 656 10281 688
rect 10281 656 10326 688
rect 10204 622 10326 656
rect 5715 410 5755 414
rect 6319 410 6359 414
rect 6923 410 6963 414
rect 7527 410 7567 414
rect 8131 410 8171 414
rect 8735 410 8775 414
rect 9339 410 9379 414
rect 9943 410 9983 414
rect 5715 378 5738 410
rect 5738 378 5755 410
rect 6319 378 6350 410
rect 6350 378 6359 410
rect 6923 378 6930 410
rect 6930 378 6962 410
rect 6962 378 6963 410
rect 7527 378 7542 410
rect 7542 378 7567 410
rect 8131 378 8154 410
rect 8154 378 8171 410
rect 8735 378 8766 410
rect 8766 378 8775 410
rect 9339 378 9342 410
rect 9342 378 9378 410
rect 9378 378 9379 410
rect 9943 378 9954 410
rect 9954 378 9983 410
rect 5715 374 5755 378
rect 6319 374 6359 378
rect 6923 374 6963 378
rect 7527 374 7567 378
rect 8131 374 8171 378
rect 8735 374 8775 378
rect 9339 374 9379 378
rect 9943 374 9983 378
<< metal2 >>
rect 3046 3359 3086 3852
rect 3046 3263 3086 3319
rect 3046 3205 3086 3223
rect 5715 3832 5755 3852
rect 5976 3230 6098 3852
rect 5976 1810 6098 2042
rect 5976 613 6098 622
rect 6319 3832 6359 3852
rect 5715 0 5755 20
rect 6580 3230 6702 3852
rect 6580 1810 6702 2042
rect 6580 613 6702 622
rect 6923 3832 6963 3852
rect 6319 0 6359 20
rect 7184 3230 7306 3852
rect 7184 1810 7306 2042
rect 7184 613 7306 622
rect 7527 3832 7567 3852
rect 6923 0 6963 20
rect 7788 3230 7910 3852
rect 7788 1810 7910 2042
rect 7788 613 7910 622
rect 8131 3832 8171 3852
rect 7527 0 7567 20
rect 8392 3230 8514 3852
rect 8392 1810 8514 2042
rect 8392 613 8514 622
rect 8735 3832 8775 3852
rect 8131 0 8171 20
rect 8996 3230 9118 3852
rect 8996 1810 9118 2042
rect 8996 613 9118 622
rect 9339 3832 9379 3852
rect 8735 0 8775 20
rect 9600 3230 9722 3852
rect 9600 1810 9722 2042
rect 9600 613 9722 622
rect 9943 3832 9983 3852
rect 9339 0 9379 20
rect 10204 3230 10326 3852
rect 10204 1810 10326 2042
rect 10204 613 10326 622
rect 9943 0 9983 20
<< via2 >>
rect 5715 3478 5755 3832
rect 5715 3438 5755 3478
rect 5715 3230 5755 3438
rect 5715 2042 5755 3230
rect 5715 1810 5755 2042
rect 5715 622 5755 1810
rect 5715 414 5755 622
rect 6319 3478 6359 3832
rect 6319 3438 6359 3478
rect 6319 3230 6359 3438
rect 6319 2042 6359 3230
rect 6319 1810 6359 2042
rect 6319 622 6359 1810
rect 5715 374 5755 414
rect 5715 20 5755 374
rect 6319 414 6359 622
rect 6923 3478 6963 3832
rect 6923 3438 6963 3478
rect 6923 3230 6963 3438
rect 6923 2042 6963 3230
rect 6923 1810 6963 2042
rect 6923 622 6963 1810
rect 6319 374 6359 414
rect 6319 20 6359 374
rect 6923 414 6963 622
rect 7527 3478 7567 3832
rect 7527 3438 7567 3478
rect 7527 3230 7567 3438
rect 7527 2042 7567 3230
rect 7527 1810 7567 2042
rect 7527 622 7567 1810
rect 6923 374 6963 414
rect 6923 20 6963 374
rect 7527 414 7567 622
rect 8131 3478 8171 3832
rect 8131 3438 8171 3478
rect 8131 3230 8171 3438
rect 8131 2042 8171 3230
rect 8131 1810 8171 2042
rect 8131 622 8171 1810
rect 7527 374 7567 414
rect 7527 20 7567 374
rect 8131 414 8171 622
rect 8735 3478 8775 3832
rect 8735 3438 8775 3478
rect 8735 3230 8775 3438
rect 8735 2042 8775 3230
rect 8735 1810 8775 2042
rect 8735 622 8775 1810
rect 8131 374 8171 414
rect 8131 20 8171 374
rect 8735 414 8775 622
rect 9339 3478 9379 3832
rect 9339 3438 9379 3478
rect 9339 3230 9379 3438
rect 9339 2042 9379 3230
rect 9339 1810 9379 2042
rect 9339 622 9379 1810
rect 8735 374 8775 414
rect 8735 20 8775 374
rect 9339 414 9379 622
rect 9943 3478 9983 3832
rect 9943 3438 9983 3478
rect 9943 3230 9983 3438
rect 9943 2042 9983 3230
rect 9943 1810 9983 2042
rect 9943 622 9983 1810
rect 9339 374 9379 414
rect 9339 20 9379 374
rect 9943 414 9983 622
rect 9943 374 9983 414
rect 9943 20 9983 374
<< metal3 >>
rect 5715 3832 5755 3841
rect 5715 11 5755 20
rect 6319 3832 6359 3841
rect 6319 11 6359 20
rect 6923 3832 6963 3841
rect 6923 11 6963 20
rect 7527 3832 7567 3841
rect 7527 11 7567 20
rect 8131 3832 8171 3841
rect 8131 11 8171 20
rect 8735 3832 8775 3841
rect 8735 11 8775 20
rect 9339 3832 9379 3841
rect 9339 11 9379 20
rect 9943 3832 9983 3841
rect 9943 11 9983 20
<< labels >>
flabel metal2 s 9600 613 9722 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 8996 613 9118 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 8392 613 8514 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 7788 613 7910 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 7184 613 7306 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 6580 613 6702 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 5976 613 6098 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
rlabel metal2 s 3046 3205 3086 3852 4 gate
port 4 nsew
flabel metal2 s 10204 613 10326 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
rlabel comment s 34 34 34 34 4 sub!
flabel comment s 3070 3220 3070 3220 0 FreeSans 400 0 0 0 dpant
flabel metal1 s 173 3791 440 3839 0 FreeSans 51 0 0 0 iovss
port 1 nsew
flabel metal1 s 521 3436 763 3479 0 FreeSans 51 0 0 0 iovdd
port 2 nsew
<< properties >>
string device primitive
string GDS_END 26313672
string GDS_FILE sg13g2_io.gds
string GDS_START 26119954
<< end >>
