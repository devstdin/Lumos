magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< m2fill >>
rect 3360 19837 3760 20837
rect 4000 19837 4400 20837
rect 4640 19837 5040 20837
rect 5597 20641 5997 21641
rect 3360 18597 3760 19597
rect 4000 18597 4400 19597
rect 4640 18597 5040 19597
rect 5596 19129 5996 20129
rect 3360 17357 3760 18357
rect 4000 17357 4400 18357
rect 20380 17797 20780 18797
rect 3360 16117 3760 17117
rect 4000 16117 4400 17117
rect 3360 14877 3760 15877
rect 3360 13637 3760 14637
rect 3360 12397 3760 13397
rect 3360 11157 3760 12157
rect 21584 11077 21984 12077
rect 3360 9917 3760 10917
rect 3360 8677 3760 9677
rect 6016 7033 6416 8033
rect 17440 7500 17840 8500
rect 19360 7500 19760 8500
rect 20000 7500 20400 8500
rect 14240 6260 14640 7260
rect 14880 6260 15280 7260
rect 15520 6260 15920 7260
rect 16160 6260 16560 7260
rect 16800 6260 17200 7260
rect 17440 6260 17840 7260
rect 18080 6260 18480 7260
rect 18720 6260 19120 7260
rect 19360 6260 19760 7260
rect 20000 6260 20400 7260
rect 3360 5020 3760 6020
rect 4000 5020 4400 6020
rect 4640 5020 5040 6020
rect 5280 5020 5680 6020
rect 6560 5020 6960 6020
rect 7840 5020 8240 6020
rect 8480 5020 8880 6020
rect 9120 5020 9520 6020
rect 9760 5020 10160 6020
rect 10400 5020 10800 6020
rect 11040 5020 11440 6020
rect 11680 5020 12080 6020
rect 12320 5020 12720 6020
rect 14240 5020 14640 6020
rect 14880 5020 15280 6020
rect 15520 5020 15920 6020
rect 16160 5020 16560 6020
rect 16800 5020 17200 6020
rect 17440 5020 17840 6020
rect 18080 5020 18480 6020
rect 18720 5020 19120 6020
rect 19360 5020 19760 6020
rect 20000 5020 20400 6020
rect 3360 3780 3760 4780
rect 4000 3780 4400 4780
rect 4640 3780 5040 4780
rect 5280 3780 5680 4780
rect 6560 3780 6960 4780
rect 7200 3780 7600 4780
rect 7840 3780 8240 4780
rect 8480 3780 8880 4780
rect 9120 3780 9520 4780
rect 9760 3780 10160 4780
rect 10400 3780 10800 4780
rect 11040 3780 11440 4780
rect 11680 3780 12080 4780
rect 12320 3780 12720 4780
rect 14240 3780 14640 4780
rect 14880 3780 15280 4780
rect 15520 3780 15920 4780
rect 16160 3780 16560 4780
rect 16800 3780 17200 4780
rect 17440 3780 17840 4780
rect 18080 3780 18480 4780
rect 18720 3780 19120 4780
rect 19360 3780 19760 4780
rect 20000 3780 20400 4780
<< m3fill >>
rect 3360 21436 4360 21836
rect 3360 20796 4360 21196
rect 4600 20796 5600 21196
rect 18921 20732 19921 21132
rect 20161 20732 21161 21132
rect 3360 20156 4360 20556
rect 4600 20156 5600 20556
rect 16441 20092 17441 20492
rect 3360 19516 4360 19916
rect 4600 19516 5600 19916
rect 19465 19516 20465 19916
rect 20705 19516 21705 19916
rect 3360 18876 4360 19276
rect 3360 18236 4360 18636
rect 20769 18140 21769 18540
rect 3360 17596 4360 17996
rect 18289 17500 19289 17900
rect 19529 17500 20529 17900
rect 3360 16956 4360 17356
rect 3360 16316 4360 16716
rect 3360 15676 4360 16076
rect 3360 14556 4360 14956
rect 12053 14524 13053 14924
rect 17113 14716 18113 15116
rect 20473 14584 21473 14984
rect 3360 13916 4360 14316
rect 8001 13756 9001 14156
rect 3360 13276 4360 13676
rect 15937 13276 16937 13676
rect 20641 13072 21641 13472
rect 3360 12220 4360 12620
rect 17449 11740 18449 12140
rect 20557 11932 21557 12332
rect 3360 10940 4360 11340
rect 3360 10300 4360 10700
rect 4600 10300 5600 10700
rect 5840 10300 6840 10700
rect 20221 10396 21221 10796
rect 3360 9308 4360 9708
rect 3360 8668 4360 9068
rect 19213 8860 20213 9260
rect 20453 8860 21453 9260
rect 15760 7620 16760 8020
rect 17000 7620 18000 8020
rect 18240 7620 19240 8020
rect 19480 7620 20480 8020
rect 20720 7620 21720 8020
rect 3360 7132 4360 7532
rect 14520 6980 15520 7380
rect 15760 6980 16760 7380
rect 17000 6980 18000 7380
rect 18240 6980 19240 7380
rect 19480 6980 20480 7380
rect 10800 6340 11800 6740
rect 12040 6340 13040 6740
rect 13280 6340 14280 6740
rect 14520 6340 15520 6740
rect 15760 6340 16760 6740
rect 17000 6340 18000 6740
rect 18240 6340 19240 6740
rect 19480 6340 20480 6740
rect 3360 5700 4360 6100
rect 4600 5700 5600 6100
rect 5840 5700 6840 6100
rect 7080 5700 8080 6100
rect 8320 5700 9320 6100
rect 9560 5700 10560 6100
rect 10800 5700 11800 6100
rect 12040 5700 13040 6100
rect 14520 5700 15520 6100
rect 15760 5700 16760 6100
rect 17000 5700 18000 6100
rect 18240 5700 19240 6100
rect 19480 5700 20480 6100
rect 20720 5700 21720 6100
rect 3360 5060 4360 5460
rect 4600 5060 5600 5460
rect 7080 5060 8080 5460
rect 8320 5060 9320 5460
rect 9560 5060 10560 5460
rect 10800 5060 11800 5460
rect 12040 5060 13040 5460
rect 13280 5060 14280 5460
rect 14520 5060 15520 5460
rect 15760 5060 16760 5460
rect 17000 5060 18000 5460
rect 18240 5060 19240 5460
rect 19480 5060 20480 5460
rect 3360 4420 4360 4820
rect 4600 4420 5600 4820
rect 5840 4420 6840 4820
rect 7080 4420 8080 4820
rect 8320 4420 9320 4820
rect 9560 4420 10560 4820
rect 10800 4420 11800 4820
rect 12040 4420 13040 4820
rect 14520 4420 15520 4820
rect 15760 4420 16760 4820
rect 17000 4420 18000 4820
rect 18240 4420 19240 4820
rect 19480 4420 20480 4820
rect 20720 4420 21720 4820
rect 3360 3780 4360 4180
rect 4600 3780 5600 4180
rect 7080 3780 8080 4180
rect 8320 3780 9320 4180
rect 9560 3780 10560 4180
rect 10800 3780 11800 4180
rect 12040 3780 13040 4180
rect 13280 3780 14280 4180
rect 14520 3780 15520 4180
rect 15760 3780 16760 4180
rect 17000 3780 18000 4180
rect 18240 3780 19240 4180
rect 19480 3780 20480 4180
<< m4fill >>
rect 3360 19900 3760 20900
rect 4000 19900 4400 20900
rect 4640 19900 5040 20900
rect 5280 19900 5680 20900
rect 6560 19900 6960 20900
rect 7200 19900 7600 20900
rect 7840 19900 8240 20900
rect 8480 19900 8880 20900
rect 9120 19900 9520 20900
rect 9760 19900 10160 20900
rect 10400 19900 10800 20900
rect 11040 19900 11440 20900
rect 11680 19900 12080 20900
rect 12320 19900 12720 20900
rect 12960 19900 13360 20900
rect 13600 19900 14000 20900
rect 14240 19900 14640 20900
rect 14880 19900 15280 20900
rect 15520 19900 15920 20900
rect 16160 19900 16560 20900
rect 16800 19900 17200 20900
rect 17440 19900 17840 20900
rect 18080 19900 18480 20900
rect 18720 19900 19120 20900
rect 19360 19900 19760 20900
rect 20000 19900 20400 20900
rect 3360 18660 3760 19660
rect 4000 18660 4400 19660
rect 4640 18660 5040 19660
rect 7200 18660 7600 19660
rect 7840 18660 8240 19660
rect 8480 18660 8880 19660
rect 9120 18660 9520 19660
rect 9760 18660 10160 19660
rect 11040 18660 11440 19660
rect 11680 18660 12080 19660
rect 12320 18660 12720 19660
rect 14240 18660 14640 19660
rect 14880 18660 15280 19660
rect 15520 18660 15920 19660
rect 16160 18660 16560 19660
rect 16800 18660 17200 19660
rect 17440 18660 17840 19660
rect 18080 18660 18480 19660
rect 18720 18660 19120 19660
rect 19360 18660 19760 19660
rect 20000 18660 20400 19660
rect 3360 17420 3760 18420
rect 4000 17420 4400 18420
rect 4640 17420 5040 18420
rect 6016 17617 6416 18617
rect 7200 17420 7600 18420
rect 7840 17420 8240 18420
rect 8480 17420 8880 18420
rect 9120 17420 9520 18420
rect 9760 17420 10160 18420
rect 11040 17420 11440 18420
rect 11680 17420 12080 18420
rect 12320 17420 12720 18420
rect 14240 17420 14640 18420
rect 14880 17420 15280 18420
rect 15520 17420 15920 18420
rect 16160 17420 16560 18420
rect 16800 17420 17200 18420
rect 17440 17420 17840 18420
rect 18080 17420 18480 18420
rect 18720 17420 19120 18420
rect 19360 17420 19760 18420
rect 20000 17420 20400 18420
rect 3360 16180 3760 17180
rect 4000 16180 4400 17180
rect 4640 16180 5040 17180
rect 6016 16105 6416 17105
rect 7200 16180 7600 17180
rect 7840 16180 8240 17180
rect 8480 16180 8880 17180
rect 9120 16180 9520 17180
rect 9760 16180 10160 17180
rect 11040 16180 11440 17180
rect 11680 16180 12080 17180
rect 12320 16180 12720 17180
rect 14240 16180 14640 17180
rect 14880 16180 15280 17180
rect 15520 16180 15920 17180
rect 16160 16180 16560 17180
rect 16800 16180 17200 17180
rect 17440 16180 17840 17180
rect 18080 16180 18480 17180
rect 18720 16180 19120 17180
rect 19360 16180 19760 17180
rect 20000 16180 20400 17180
rect 3360 14940 3760 15940
rect 4000 14940 4400 15940
rect 4640 14940 5040 15940
rect 3360 13700 3760 14700
rect 4000 13700 4400 14700
rect 4640 13700 5040 14700
rect 6016 14593 6416 15593
rect 7200 14940 7600 15940
rect 7840 14940 8240 15940
rect 8480 14940 8880 15940
rect 9120 14940 9520 15940
rect 9760 14940 10160 15940
rect 11040 14940 11440 15940
rect 11680 14940 12080 15940
rect 12320 14940 12720 15940
rect 14240 14940 14640 15940
rect 14880 14940 15280 15940
rect 15520 14940 15920 15940
rect 16160 14940 16560 15940
rect 16800 14940 17200 15940
rect 17440 14940 17840 15940
rect 18080 14940 18480 15940
rect 18720 14940 19120 15940
rect 19360 14940 19760 15940
rect 20000 14940 20400 15940
rect 3360 12460 3760 13460
rect 4000 12460 4400 13460
rect 4640 12460 5040 13460
rect 6016 13081 6416 14081
rect 7200 13700 7600 14700
rect 7840 13700 8240 14700
rect 8480 13700 8880 14700
rect 9120 13700 9520 14700
rect 11040 13700 11440 14700
rect 11680 13700 12080 14700
rect 12320 13700 12720 14700
rect 14240 13700 14640 14700
rect 14880 13700 15280 14700
rect 15520 13700 15920 14700
rect 16160 13700 16560 14700
rect 16800 13700 17200 14700
rect 18080 13700 18480 14700
rect 18720 13700 19120 14700
rect 19360 13700 19760 14700
rect 20000 13700 20400 14700
rect 7200 12460 7600 13460
rect 7840 12460 8240 13460
rect 8480 12460 8880 13460
rect 9120 12460 9520 13460
rect 11040 12460 11440 13460
rect 11680 12460 12080 13460
rect 12320 12460 12720 13460
rect 14240 12460 14640 13460
rect 14880 12460 15280 13460
rect 15520 12460 15920 13460
rect 16160 12460 16560 13460
rect 16800 12460 17200 13460
rect 18080 12460 18480 13460
rect 18720 12460 19120 13460
rect 19360 12460 19760 13460
rect 20000 12460 20400 13460
rect 3360 11220 3760 12220
rect 4000 11220 4400 12220
rect 4640 11220 5040 12220
rect 5280 11220 5680 12220
rect 7200 11220 7600 12220
rect 7840 11220 8240 12220
rect 8480 11220 8880 12220
rect 9120 11220 9520 12220
rect 9760 11220 10160 12220
rect 10400 11220 10800 12220
rect 11040 11220 11440 12220
rect 11680 11220 12080 12220
rect 14240 11220 14640 12220
rect 14880 11220 15280 12220
rect 15520 11220 15920 12220
rect 16160 11220 16560 12220
rect 16800 11220 17200 12220
rect 18080 11220 18480 12220
rect 18720 11220 19120 12220
rect 19360 11220 19760 12220
rect 20000 11220 20400 12220
rect 3360 9980 3760 10980
rect 4000 9980 4400 10980
rect 4640 9980 5040 10980
rect 6560 9980 6960 10980
rect 7200 9980 7600 10980
rect 7840 9980 8240 10980
rect 8480 9980 8880 10980
rect 9120 9980 9520 10980
rect 9760 9980 10160 10980
rect 10400 9980 10800 10980
rect 11040 9980 11440 10980
rect 11680 9980 12080 10980
rect 14240 9980 14640 10980
rect 14880 9980 15280 10980
rect 15520 9980 15920 10980
rect 16160 9980 16560 10980
rect 16800 9980 17200 10980
rect 18080 9980 18480 10980
rect 18720 9980 19120 10980
rect 19360 9980 19760 10980
rect 20000 9980 20400 10980
rect 3360 8740 3760 9740
rect 4000 8740 4400 9740
rect 4640 8740 5040 9740
rect 6560 8740 6960 9740
rect 7200 8740 7600 9740
rect 7840 8740 8240 9740
rect 8480 8740 8880 9740
rect 9120 8740 9520 9740
rect 9760 8740 10160 9740
rect 10400 8740 10800 9740
rect 11040 8740 11440 9740
rect 11680 8740 12080 9740
rect 12320 8740 12720 9740
rect 14240 8740 14640 9740
rect 14880 8740 15280 9740
rect 15520 8740 15920 9740
rect 16160 8740 16560 9740
rect 16800 8740 17200 9740
rect 17440 8740 17840 9740
rect 18080 8740 18480 9740
rect 18720 8740 19120 9740
rect 19360 8740 19760 9740
rect 20000 8740 20400 9740
rect 3360 7500 3760 8500
rect 4000 7500 4400 8500
rect 4640 7500 5040 8500
rect 5280 7500 5680 8500
rect 6560 7500 6960 8500
rect 7200 7500 7600 8500
rect 7840 7500 8240 8500
rect 8480 7500 8880 8500
rect 9120 7500 9520 8500
rect 9760 7500 10160 8500
rect 10400 7500 10800 8500
rect 11040 7500 11440 8500
rect 11680 7500 12080 8500
rect 12320 7500 12720 8500
rect 14240 7500 14640 8500
rect 14880 7500 15280 8500
rect 15520 7500 15920 8500
rect 16160 7500 16560 8500
rect 16800 7500 17200 8500
rect 17440 7500 17840 8500
rect 18080 7500 18480 8500
rect 18720 7500 19120 8500
rect 19360 7500 19760 8500
rect 20000 7500 20400 8500
rect 3360 6260 3760 7260
rect 4000 6260 4400 7260
rect 4640 6260 5040 7260
rect 5280 6260 5680 7260
rect 6560 6260 6960 7260
rect 7200 6260 7600 7260
rect 7840 6260 8240 7260
rect 8480 6260 8880 7260
rect 9120 6260 9520 7260
rect 9760 6260 10160 7260
rect 10400 6260 10800 7260
rect 11040 6260 11440 7260
rect 11680 6260 12080 7260
rect 12320 6260 12720 7260
rect 14240 6260 14640 7260
rect 14880 6260 15280 7260
rect 15520 6260 15920 7260
rect 16160 6260 16560 7260
rect 16800 6260 17200 7260
rect 17440 6260 17840 7260
rect 18080 6260 18480 7260
rect 18720 6260 19120 7260
rect 19360 6260 19760 7260
rect 20000 6260 20400 7260
rect 3360 5020 3760 6020
rect 4000 5020 4400 6020
rect 4640 5020 5040 6020
rect 5280 5020 5680 6020
rect 6560 5020 6960 6020
rect 7200 5020 7600 6020
rect 7840 5020 8240 6020
rect 8480 5020 8880 6020
rect 9120 5020 9520 6020
rect 9760 5020 10160 6020
rect 10400 5020 10800 6020
rect 11040 5020 11440 6020
rect 11680 5020 12080 6020
rect 12320 5020 12720 6020
rect 14240 5020 14640 6020
rect 14880 5020 15280 6020
rect 15520 5020 15920 6020
rect 16160 5020 16560 6020
rect 16800 5020 17200 6020
rect 17440 5020 17840 6020
rect 18080 5020 18480 6020
rect 18720 5020 19120 6020
rect 19360 5020 19760 6020
rect 20000 5020 20400 6020
rect 3360 3780 3760 4780
rect 4000 3780 4400 4780
rect 4640 3780 5040 4780
rect 5280 3780 5680 4780
rect 6560 3780 6960 4780
rect 7200 3780 7600 4780
rect 7840 3780 8240 4780
rect 8480 3780 8880 4780
rect 9120 3780 9520 4780
rect 9760 3780 10160 4780
rect 10400 3780 10800 4780
rect 11040 3780 11440 4780
rect 11680 3780 12080 4780
rect 12320 3780 12720 4780
rect 14240 3780 14640 4780
rect 14880 3780 15280 4780
rect 15520 3780 15920 4780
rect 16160 3780 16560 4780
rect 16800 3780 17200 4780
rect 17440 3780 17840 4780
rect 18080 3780 18480 4780
rect 18720 3780 19120 4780
rect 19360 3780 19760 4780
rect 20000 3780 20400 4780
<< m5fill >>
rect 3360 21060 4360 21460
rect 4600 21060 5600 21460
rect 5840 21060 6840 21460
rect 7080 21060 8080 21460
rect 8320 21060 9320 21460
rect 9560 21060 10560 21460
rect 10800 21060 11800 21460
rect 12040 21060 13040 21460
rect 14520 21060 15520 21460
rect 15760 21060 16760 21460
rect 17000 21060 18000 21460
rect 18240 21060 19240 21460
rect 19480 21060 20480 21460
rect 20720 21060 21720 21460
rect 3360 20420 4360 20820
rect 4600 20420 5600 20820
rect 7080 20420 8080 20820
rect 8320 20420 9320 20820
rect 9560 20420 10560 20820
rect 10800 20420 11800 20820
rect 12040 20420 13040 20820
rect 13280 20420 14280 20820
rect 14520 20420 15520 20820
rect 15760 20420 16760 20820
rect 17000 20420 18000 20820
rect 18240 20420 19240 20820
rect 19480 20420 20480 20820
rect 3360 19780 4360 20180
rect 4600 19780 5600 20180
rect 7080 19780 8080 20180
rect 8320 19780 9320 20180
rect 9560 19780 10560 20180
rect 10800 19780 11800 20180
rect 12040 19780 13040 20180
rect 14520 19780 15520 20180
rect 15760 19780 16760 20180
rect 17000 19780 18000 20180
rect 18240 19780 19240 20180
rect 19480 19780 20480 20180
rect 3360 19140 4360 19540
rect 4600 19140 5600 19540
rect 7080 19140 8080 19540
rect 8320 19140 9320 19540
rect 9560 19140 10560 19540
rect 10800 19140 11800 19540
rect 12040 19140 13040 19540
rect 14520 19140 15520 19540
rect 15760 19140 16760 19540
rect 17000 19140 18000 19540
rect 18240 19140 19240 19540
rect 19480 19140 20480 19540
rect 3360 18500 4360 18900
rect 4600 18500 5600 18900
rect 7080 18500 8080 18900
rect 8320 18500 9320 18900
rect 9560 18500 10560 18900
rect 10800 18500 11800 18900
rect 12040 18500 13040 18900
rect 13280 18500 14280 18900
rect 14520 18500 15520 18900
rect 15760 18500 16760 18900
rect 17000 18500 18000 18900
rect 18240 18500 19240 18900
rect 19480 18500 20480 18900
rect 3360 17860 4360 18260
rect 4600 17860 5600 18260
rect 5840 17860 6840 18260
rect 7080 17860 8080 18260
rect 8320 17860 9320 18260
rect 9560 17860 10560 18260
rect 10800 17860 11800 18260
rect 12040 17860 13040 18260
rect 14520 17860 15520 18260
rect 15760 17860 16760 18260
rect 17000 17860 18000 18260
rect 18240 17860 19240 18260
rect 19480 17860 20480 18260
rect 20720 17860 21720 18260
rect 3360 17220 4360 17620
rect 4600 17220 5600 17620
rect 7080 17220 8080 17620
rect 8320 17220 9320 17620
rect 9560 17220 10560 17620
rect 10800 17220 11800 17620
rect 12040 17220 13040 17620
rect 13280 17220 14280 17620
rect 14520 17220 15520 17620
rect 15760 17220 16760 17620
rect 17000 17220 18000 17620
rect 18240 17220 19240 17620
rect 19480 17220 20480 17620
rect 3360 16580 4360 16980
rect 4600 16580 5600 16980
rect 5840 16580 6840 16980
rect 7080 16580 8080 16980
rect 8320 16580 9320 16980
rect 9560 16580 10560 16980
rect 10800 16580 11800 16980
rect 12040 16580 13040 16980
rect 14520 16580 15520 16980
rect 15760 16580 16760 16980
rect 17000 16580 18000 16980
rect 18240 16580 19240 16980
rect 19480 16580 20480 16980
rect 20720 16580 21720 16980
rect 3360 15940 4360 16340
rect 4600 15940 5600 16340
rect 7080 15940 8080 16340
rect 8320 15940 9320 16340
rect 9560 15940 10560 16340
rect 10800 15940 11800 16340
rect 12040 15940 13040 16340
rect 13280 15940 14280 16340
rect 14520 15940 15520 16340
rect 15760 15940 16760 16340
rect 17000 15940 18000 16340
rect 18240 15940 19240 16340
rect 19480 15940 20480 16340
rect 3360 15300 4360 15700
rect 4600 15300 5600 15700
rect 7080 15300 8080 15700
rect 8320 15300 9320 15700
rect 9560 15300 10560 15700
rect 10800 15300 11800 15700
rect 12040 15300 13040 15700
rect 14520 15300 15520 15700
rect 15760 15300 16760 15700
rect 17000 15300 18000 15700
rect 18240 15300 19240 15700
rect 19480 15300 20480 15700
rect 3360 14660 4360 15060
rect 4600 14660 5600 15060
rect 5840 14660 6840 15060
rect 7080 14660 8080 15060
rect 8320 14660 9320 15060
rect 9560 14660 10560 15060
rect 10800 14660 11800 15060
rect 12040 14660 13040 15060
rect 14520 14660 15520 15060
rect 15760 14660 16760 15060
rect 17000 14660 18000 15060
rect 18240 14660 19240 15060
rect 19480 14660 20480 15060
rect 20720 14660 21720 15060
rect 3360 14020 4360 14420
rect 4600 14020 5600 14420
rect 7080 14020 8080 14420
rect 8320 14020 9320 14420
rect 9560 14020 10560 14420
rect 10800 14020 11800 14420
rect 12040 14020 13040 14420
rect 13280 14020 14280 14420
rect 14520 14020 15520 14420
rect 15760 14020 16760 14420
rect 17000 14020 18000 14420
rect 18240 14020 19240 14420
rect 19480 14020 20480 14420
rect 3360 13380 4360 13780
rect 4600 13380 5600 13780
rect 5840 13380 6840 13780
rect 7080 13380 8080 13780
rect 8320 13380 9320 13780
rect 9560 13380 10560 13780
rect 10800 13380 11800 13780
rect 12040 13380 13040 13780
rect 14520 13380 15520 13780
rect 15760 13380 16760 13780
rect 17000 13380 18000 13780
rect 18240 13380 19240 13780
rect 19480 13380 20480 13780
rect 20720 13380 21720 13780
rect 3360 12740 4360 13140
rect 4600 12740 5600 13140
rect 7080 12740 8080 13140
rect 8320 12740 9320 13140
rect 9560 12740 10560 13140
rect 10800 12740 11800 13140
rect 12040 12740 13040 13140
rect 13280 12740 14280 13140
rect 14520 12740 15520 13140
rect 15760 12740 16760 13140
rect 17000 12740 18000 13140
rect 18240 12740 19240 13140
rect 19480 12740 20480 13140
rect 3360 12100 4360 12500
rect 4600 12100 5600 12500
rect 5840 12100 6840 12500
rect 7080 12100 8080 12500
rect 8320 12100 9320 12500
rect 9560 12100 10560 12500
rect 10800 12100 11800 12500
rect 12040 12100 13040 12500
rect 14520 12100 15520 12500
rect 15760 12100 16760 12500
rect 17000 12100 18000 12500
rect 18240 12100 19240 12500
rect 19480 12100 20480 12500
rect 20720 12100 21720 12500
rect 3360 11460 4360 11860
rect 4600 11460 5600 11860
rect 7080 11460 8080 11860
rect 8320 11460 9320 11860
rect 9560 11460 10560 11860
rect 10800 11460 11800 11860
rect 12040 11460 13040 11860
rect 14520 11460 15520 11860
rect 15760 11460 16760 11860
rect 17000 11460 18000 11860
rect 18240 11460 19240 11860
rect 19480 11460 20480 11860
rect 3360 10820 4360 11220
rect 4600 10820 5600 11220
rect 7080 10820 8080 11220
rect 8320 10820 9320 11220
rect 9560 10820 10560 11220
rect 10800 10820 11800 11220
rect 12040 10820 13040 11220
rect 14520 10820 15520 11220
rect 15760 10820 16760 11220
rect 17000 10820 18000 11220
rect 18240 10820 19240 11220
rect 19480 10820 20480 11220
rect 3360 10180 4360 10580
rect 4600 10180 5600 10580
rect 5840 10180 6840 10580
rect 7080 10180 8080 10580
rect 8320 10180 9320 10580
rect 9560 10180 10560 10580
rect 10800 10180 11800 10580
rect 12040 10180 13040 10580
rect 14520 10180 15520 10580
rect 15760 10180 16760 10580
rect 17000 10180 18000 10580
rect 18240 10180 19240 10580
rect 19480 10180 20480 10580
rect 20720 10180 21720 10580
rect 3360 9540 4360 9940
rect 4600 9540 5600 9940
rect 7080 9540 8080 9940
rect 8320 9540 9320 9940
rect 9560 9540 10560 9940
rect 10800 9540 11800 9940
rect 12040 9540 13040 9940
rect 13280 9540 14280 9940
rect 14520 9540 15520 9940
rect 15760 9540 16760 9940
rect 17000 9540 18000 9940
rect 18240 9540 19240 9940
rect 19480 9540 20480 9940
rect 3360 8900 4360 9300
rect 4600 8900 5600 9300
rect 5840 8900 6840 9300
rect 7080 8900 8080 9300
rect 8320 8900 9320 9300
rect 9560 8900 10560 9300
rect 10800 8900 11800 9300
rect 12040 8900 13040 9300
rect 14520 8900 15520 9300
rect 15760 8900 16760 9300
rect 17000 8900 18000 9300
rect 18240 8900 19240 9300
rect 19480 8900 20480 9300
rect 20720 8900 21720 9300
rect 3360 8260 4360 8660
rect 4600 8260 5600 8660
rect 7080 8260 8080 8660
rect 8320 8260 9320 8660
rect 9560 8260 10560 8660
rect 10800 8260 11800 8660
rect 12040 8260 13040 8660
rect 13280 8260 14280 8660
rect 14520 8260 15520 8660
rect 15760 8260 16760 8660
rect 17000 8260 18000 8660
rect 18240 8260 19240 8660
rect 19480 8260 20480 8660
rect 3360 7620 4360 8020
rect 4600 7620 5600 8020
rect 5840 7620 6840 8020
rect 7080 7620 8080 8020
rect 8320 7620 9320 8020
rect 9560 7620 10560 8020
rect 10800 7620 11800 8020
rect 12040 7620 13040 8020
rect 14520 7620 15520 8020
rect 15760 7620 16760 8020
rect 17000 7620 18000 8020
rect 18240 7620 19240 8020
rect 19480 7620 20480 8020
rect 20720 7620 21720 8020
rect 3360 6980 4360 7380
rect 4600 6980 5600 7380
rect 7080 6980 8080 7380
rect 8320 6980 9320 7380
rect 9560 6980 10560 7380
rect 10800 6980 11800 7380
rect 12040 6980 13040 7380
rect 14520 6980 15520 7380
rect 15760 6980 16760 7380
rect 17000 6980 18000 7380
rect 18240 6980 19240 7380
rect 19480 6980 20480 7380
rect 3360 6340 4360 6740
rect 4600 6340 5600 6740
rect 7080 6340 8080 6740
rect 8320 6340 9320 6740
rect 9560 6340 10560 6740
rect 10800 6340 11800 6740
rect 12040 6340 13040 6740
rect 13280 6340 14280 6740
rect 14520 6340 15520 6740
rect 15760 6340 16760 6740
rect 17000 6340 18000 6740
rect 18240 6340 19240 6740
rect 19480 6340 20480 6740
rect 3360 5700 4360 6100
rect 4600 5700 5600 6100
rect 5840 5700 6840 6100
rect 7080 5700 8080 6100
rect 8320 5700 9320 6100
rect 9560 5700 10560 6100
rect 10800 5700 11800 6100
rect 12040 5700 13040 6100
rect 14520 5700 15520 6100
rect 15760 5700 16760 6100
rect 17000 5700 18000 6100
rect 18240 5700 19240 6100
rect 19480 5700 20480 6100
rect 20720 5700 21720 6100
rect 3360 5060 4360 5460
rect 4600 5060 5600 5460
rect 7080 5060 8080 5460
rect 8320 5060 9320 5460
rect 9560 5060 10560 5460
rect 10800 5060 11800 5460
rect 12040 5060 13040 5460
rect 13280 5060 14280 5460
rect 14520 5060 15520 5460
rect 15760 5060 16760 5460
rect 17000 5060 18000 5460
rect 18240 5060 19240 5460
rect 19480 5060 20480 5460
rect 3360 4420 4360 4820
rect 4600 4420 5600 4820
rect 5840 4420 6840 4820
rect 7080 4420 8080 4820
rect 8320 4420 9320 4820
rect 9560 4420 10560 4820
rect 10800 4420 11800 4820
rect 12040 4420 13040 4820
rect 14520 4420 15520 4820
rect 15760 4420 16760 4820
rect 17000 4420 18000 4820
rect 18240 4420 19240 4820
rect 19480 4420 20480 4820
rect 20720 4420 21720 4820
rect 3360 3780 4360 4180
rect 4600 3780 5600 4180
rect 7080 3780 8080 4180
rect 8320 3780 9320 4180
rect 9560 3780 10560 4180
rect 10800 3780 11800 4180
rect 12040 3780 13040 4180
rect 13280 3780 14280 4180
rect 14520 3780 15520 4180
rect 15760 3780 16760 4180
rect 17000 3780 18000 4180
rect 18240 3780 19240 4180
rect 19480 3780 20480 4180
<< m6fill >>
rect 3440 19380 4440 21380
rect 7280 19380 8280 21380
rect 8880 19380 9880 21380
rect 10480 19380 11480 21380
rect 14840 19380 15840 21380
rect 16440 19380 17440 21380
rect 18040 19380 19040 21380
rect 3440 16780 4440 18780
rect 7280 16780 8280 18780
rect 8880 16780 9880 18780
rect 10480 16780 11480 18780
rect 14840 16780 15840 18780
rect 16440 16780 17440 18780
rect 18040 16780 19040 18780
rect 3440 14180 4440 16180
rect 7280 14180 8280 16180
rect 8880 14180 9880 16180
rect 10480 14180 11480 16180
rect 14840 14180 15840 16180
rect 16440 14180 17440 16180
rect 18040 14180 19040 16180
rect 3440 11580 4440 13580
rect 7280 11580 8280 13580
rect 8880 11580 9880 13580
rect 10480 11580 11480 13580
rect 14840 11580 15840 13580
rect 16440 11580 17440 13580
rect 18040 11580 19040 13580
rect 3440 8980 4440 10980
rect 7280 8980 8280 10980
rect 8880 8980 9880 10980
rect 10480 8980 11480 10980
rect 14840 8980 15840 10980
rect 16440 8980 17440 10980
rect 18040 8980 19040 10980
rect 3440 6380 4440 8380
rect 7280 6380 8280 8380
rect 8880 6380 9880 8380
rect 10480 6380 11480 8380
rect 14840 6380 15840 8380
rect 16440 6380 17440 8380
rect 18040 6380 19040 8380
rect 3440 3780 4440 5780
rect 7280 3780 8280 5780
rect 8880 3780 9880 5780
rect 10480 3780 11480 5780
rect 14840 3780 15840 5780
rect 16440 3780 17440 5780
rect 18040 3780 19040 5780
<< m7fill >>
rect 3360 18454 5360 19454
rect 5960 18454 7960 19454
rect 8560 18454 10560 19454
rect 11160 18454 13160 19454
rect 13760 18454 15760 19454
rect 16360 18454 18360 19454
rect 18960 18454 20960 19454
rect 3360 16854 5360 17854
rect 5960 16854 7960 17854
rect 8560 16854 10560 17854
rect 11160 16854 13160 17854
rect 13760 16854 15760 17854
rect 16360 16854 18360 17854
rect 18960 16854 20960 17854
rect 3360 15254 5360 16254
rect 5960 15254 7960 16254
rect 8560 15254 10560 16254
rect 11160 15254 13160 16254
rect 13760 15254 15760 16254
rect 16360 15254 18360 16254
rect 18960 15254 20960 16254
rect 3360 10894 5360 11894
rect 5960 10894 7960 11894
rect 8560 10894 10560 11894
rect 11160 10894 13160 11894
rect 13760 10894 15760 11894
rect 16360 10894 18360 11894
rect 18960 10894 20960 11894
rect 3360 9294 5360 10294
rect 5960 9294 7960 10294
rect 8560 9294 10560 10294
rect 11160 9294 13160 10294
rect 13760 9294 15760 10294
rect 16360 9294 18360 10294
rect 18960 9294 20960 10294
rect 3360 7694 5360 8694
rect 5960 7694 7960 8694
rect 8560 7694 10560 8694
rect 11160 7694 13160 8694
rect 13760 7694 15760 8694
rect 16360 7694 18360 8694
rect 18960 7694 20960 8694
rect 3360 3860 5360 4860
rect 5960 3860 7960 4860
rect 8560 3860 10560 4860
rect 11160 3860 13160 4860
rect 13760 3860 15760 4860
rect 16360 3860 18360 4860
rect 18960 3860 20960 4860
<< properties >>
string GDS_END 71662
string GDS_FILE 6_final.gds
string GDS_START 9194
<< end >>
