magic
tech ihp-sg13g2
timestamp 1752522241
<< error_p >>
rect -18 3030 -13 3035
rect 13 3030 18 3035
rect 121 3030 126 3035
rect 152 3030 157 3035
rect 260 3030 265 3035
rect 291 3030 296 3035
rect 399 3030 404 3035
rect 430 3030 435 3035
rect 538 3030 543 3035
rect 569 3030 574 3035
rect 677 3030 682 3035
rect 708 3030 713 3035
rect 816 3030 821 3035
rect 847 3030 852 3035
rect 955 3030 960 3035
rect 986 3030 991 3035
rect 1094 3030 1099 3035
rect 1125 3030 1130 3035
rect 1233 3030 1238 3035
rect 1264 3030 1269 3035
rect 1372 3030 1377 3035
rect 1403 3030 1408 3035
rect 1511 3030 1516 3035
rect 1542 3030 1547 3035
rect 1650 3030 1655 3035
rect 1681 3030 1686 3035
rect 1789 3030 1794 3035
rect 1820 3030 1825 3035
rect 1928 3030 1933 3035
rect 1959 3030 1964 3035
rect 2067 3030 2072 3035
rect 2098 3030 2103 3035
rect 2206 3030 2211 3035
rect 2237 3030 2242 3035
rect 2345 3030 2350 3035
rect 2376 3030 2381 3035
rect 2484 3030 2489 3035
rect 2515 3030 2520 3035
rect 2623 3030 2628 3035
rect 2654 3030 2659 3035
rect 2762 3030 2767 3035
rect 2793 3030 2798 3035
rect 2901 3030 2906 3035
rect 2932 3030 2937 3035
rect 3040 3030 3045 3035
rect 3071 3030 3076 3035
rect 3179 3030 3184 3035
rect 3210 3030 3215 3035
rect 3318 3030 3323 3035
rect 3349 3030 3354 3035
rect 3457 3030 3462 3035
rect 3488 3030 3493 3035
rect 3596 3030 3601 3035
rect 3627 3030 3632 3035
rect 3735 3030 3740 3035
rect 3766 3030 3771 3035
rect 3874 3030 3879 3035
rect 3905 3030 3910 3035
rect 4013 3030 4018 3035
rect 4044 3030 4049 3035
rect -23 3025 23 3030
rect 116 3025 162 3030
rect 255 3025 301 3030
rect 394 3025 440 3030
rect 533 3025 579 3030
rect 672 3025 718 3030
rect 811 3025 857 3030
rect 950 3025 996 3030
rect 1089 3025 1135 3030
rect 1228 3025 1274 3030
rect 1367 3025 1413 3030
rect 1506 3025 1552 3030
rect 1645 3025 1691 3030
rect 1784 3025 1830 3030
rect 1923 3025 1969 3030
rect 2062 3025 2108 3030
rect 2201 3025 2247 3030
rect 2340 3025 2386 3030
rect 2479 3025 2525 3030
rect 2618 3025 2664 3030
rect 2757 3025 2803 3030
rect 2896 3025 2942 3030
rect 3035 3025 3081 3030
rect 3174 3025 3220 3030
rect 3313 3025 3359 3030
rect 3452 3025 3498 3030
rect 3591 3025 3637 3030
rect 3730 3025 3776 3030
rect 3869 3025 3915 3030
rect 4008 3025 4054 3030
rect -18 3019 18 3025
rect 121 3019 157 3025
rect 260 3019 296 3025
rect 399 3019 435 3025
rect 538 3019 574 3025
rect 677 3019 713 3025
rect 816 3019 852 3025
rect 955 3019 991 3025
rect 1094 3019 1130 3025
rect 1233 3019 1269 3025
rect 1372 3019 1408 3025
rect 1511 3019 1547 3025
rect 1650 3019 1686 3025
rect 1789 3019 1825 3025
rect 1928 3019 1964 3025
rect 2067 3019 2103 3025
rect 2206 3019 2242 3025
rect 2345 3019 2381 3025
rect 2484 3019 2520 3025
rect 2623 3019 2659 3025
rect 2762 3019 2798 3025
rect 2901 3019 2937 3025
rect 3040 3019 3076 3025
rect 3179 3019 3215 3025
rect 3318 3019 3354 3025
rect 3457 3019 3493 3025
rect 3596 3019 3632 3025
rect 3735 3019 3771 3025
rect 3874 3019 3910 3025
rect 4013 3019 4049 3025
rect -23 3014 23 3019
rect 116 3014 162 3019
rect 255 3014 301 3019
rect 394 3014 440 3019
rect 533 3014 579 3019
rect 672 3014 718 3019
rect 811 3014 857 3019
rect 950 3014 996 3019
rect 1089 3014 1135 3019
rect 1228 3014 1274 3019
rect 1367 3014 1413 3019
rect 1506 3014 1552 3019
rect 1645 3014 1691 3019
rect 1784 3014 1830 3019
rect 1923 3014 1969 3019
rect 2062 3014 2108 3019
rect 2201 3014 2247 3019
rect 2340 3014 2386 3019
rect 2479 3014 2525 3019
rect 2618 3014 2664 3019
rect 2757 3014 2803 3019
rect 2896 3014 2942 3019
rect 3035 3014 3081 3019
rect 3174 3014 3220 3019
rect 3313 3014 3359 3019
rect 3452 3014 3498 3019
rect 3591 3014 3637 3019
rect 3730 3014 3776 3019
rect 3869 3014 3915 3019
rect 4008 3014 4054 3019
rect -18 3009 -13 3014
rect 13 3009 18 3014
rect 121 3009 126 3014
rect 152 3009 157 3014
rect 260 3009 265 3014
rect 291 3009 296 3014
rect 399 3009 404 3014
rect 430 3009 435 3014
rect 538 3009 543 3014
rect 569 3009 574 3014
rect 677 3009 682 3014
rect 708 3009 713 3014
rect 816 3009 821 3014
rect 847 3009 852 3014
rect 955 3009 960 3014
rect 986 3009 991 3014
rect 1094 3009 1099 3014
rect 1125 3009 1130 3014
rect 1233 3009 1238 3014
rect 1264 3009 1269 3014
rect 1372 3009 1377 3014
rect 1403 3009 1408 3014
rect 1511 3009 1516 3014
rect 1542 3009 1547 3014
rect 1650 3009 1655 3014
rect 1681 3009 1686 3014
rect 1789 3009 1794 3014
rect 1820 3009 1825 3014
rect 1928 3009 1933 3014
rect 1959 3009 1964 3014
rect 2067 3009 2072 3014
rect 2098 3009 2103 3014
rect 2206 3009 2211 3014
rect 2237 3009 2242 3014
rect 2345 3009 2350 3014
rect 2376 3009 2381 3014
rect 2484 3009 2489 3014
rect 2515 3009 2520 3014
rect 2623 3009 2628 3014
rect 2654 3009 2659 3014
rect 2762 3009 2767 3014
rect 2793 3009 2798 3014
rect 2901 3009 2906 3014
rect 2932 3009 2937 3014
rect 3040 3009 3045 3014
rect 3071 3009 3076 3014
rect 3179 3009 3184 3014
rect 3210 3009 3215 3014
rect 3318 3009 3323 3014
rect 3349 3009 3354 3014
rect 3457 3009 3462 3014
rect 3488 3009 3493 3014
rect 3596 3009 3601 3014
rect 3627 3009 3632 3014
rect 3735 3009 3740 3014
rect 3766 3009 3771 3014
rect 3874 3009 3879 3014
rect 3905 3009 3910 3014
rect 4013 3009 4018 3014
rect 4044 3009 4049 3014
rect -52 2993 -47 2998
rect -41 2993 -36 2998
rect 36 2993 41 2998
rect 47 2993 52 2998
rect 87 2993 92 2998
rect 98 2993 103 2998
rect 175 2993 180 2998
rect 186 2993 191 2998
rect 226 2993 231 2998
rect 237 2993 242 2998
rect 314 2993 319 2998
rect 325 2993 330 2998
rect 365 2993 370 2998
rect 376 2993 381 2998
rect 453 2993 458 2998
rect 464 2993 469 2998
rect 504 2993 509 2998
rect 515 2993 520 2998
rect 592 2993 597 2998
rect 603 2993 608 2998
rect 643 2993 648 2998
rect 654 2993 659 2998
rect 731 2993 736 2998
rect 742 2993 747 2998
rect 782 2993 787 2998
rect 793 2993 798 2998
rect 870 2993 875 2998
rect 881 2993 886 2998
rect 921 2993 926 2998
rect 932 2993 937 2998
rect 1009 2993 1014 2998
rect 1020 2993 1025 2998
rect 1060 2993 1065 2998
rect 1071 2993 1076 2998
rect 1148 2993 1153 2998
rect 1159 2993 1164 2998
rect 1199 2993 1204 2998
rect 1210 2993 1215 2998
rect 1287 2993 1292 2998
rect 1298 2993 1303 2998
rect 1338 2993 1343 2998
rect 1349 2993 1354 2998
rect 1426 2993 1431 2998
rect 1437 2993 1442 2998
rect 1477 2993 1482 2998
rect 1488 2993 1493 2998
rect 1565 2993 1570 2998
rect 1576 2993 1581 2998
rect 1616 2993 1621 2998
rect 1627 2993 1632 2998
rect 1704 2993 1709 2998
rect 1715 2993 1720 2998
rect 1755 2993 1760 2998
rect 1766 2993 1771 2998
rect 1843 2993 1848 2998
rect 1854 2993 1859 2998
rect 1894 2993 1899 2998
rect 1905 2993 1910 2998
rect 1982 2993 1987 2998
rect 1993 2993 1998 2998
rect 2033 2993 2038 2998
rect 2044 2993 2049 2998
rect 2121 2993 2126 2998
rect 2132 2993 2137 2998
rect 2172 2993 2177 2998
rect 2183 2993 2188 2998
rect 2260 2993 2265 2998
rect 2271 2993 2276 2998
rect 2311 2993 2316 2998
rect 2322 2993 2327 2998
rect 2399 2993 2404 2998
rect 2410 2993 2415 2998
rect 2450 2993 2455 2998
rect 2461 2993 2466 2998
rect 2538 2993 2543 2998
rect 2549 2993 2554 2998
rect 2589 2993 2594 2998
rect 2600 2993 2605 2998
rect 2677 2993 2682 2998
rect 2688 2993 2693 2998
rect 2728 2993 2733 2998
rect 2739 2993 2744 2998
rect 2816 2993 2821 2998
rect 2827 2993 2832 2998
rect 2867 2993 2872 2998
rect 2878 2993 2883 2998
rect 2955 2993 2960 2998
rect 2966 2993 2971 2998
rect 3006 2993 3011 2998
rect 3017 2993 3022 2998
rect 3094 2993 3099 2998
rect 3105 2993 3110 2998
rect 3145 2993 3150 2998
rect 3156 2993 3161 2998
rect 3233 2993 3238 2998
rect 3244 2993 3249 2998
rect 3284 2993 3289 2998
rect 3295 2993 3300 2998
rect 3372 2993 3377 2998
rect 3383 2993 3388 2998
rect 3423 2993 3428 2998
rect 3434 2993 3439 2998
rect 3511 2993 3516 2998
rect 3522 2993 3527 2998
rect 3562 2993 3567 2998
rect 3573 2993 3578 2998
rect 3650 2993 3655 2998
rect 3661 2993 3666 2998
rect 3701 2993 3706 2998
rect 3712 2993 3717 2998
rect 3789 2993 3794 2998
rect 3800 2993 3805 2998
rect 3840 2993 3845 2998
rect 3851 2993 3856 2998
rect 3928 2993 3933 2998
rect 3939 2993 3944 2998
rect 3979 2993 3984 2998
rect 3990 2993 3995 2998
rect 4067 2993 4072 2998
rect 4078 2993 4083 2998
rect -57 2988 -52 2993
rect -36 2988 -31 2993
rect 31 2988 36 2993
rect 52 2988 57 2993
rect 82 2988 87 2993
rect 103 2988 108 2993
rect 170 2988 175 2993
rect 191 2988 196 2993
rect 221 2988 226 2993
rect 242 2988 247 2993
rect 309 2988 314 2993
rect 330 2988 335 2993
rect 360 2988 365 2993
rect 381 2988 386 2993
rect 448 2988 453 2993
rect 469 2988 474 2993
rect 499 2988 504 2993
rect 520 2988 525 2993
rect 587 2988 592 2993
rect 608 2988 613 2993
rect 638 2988 643 2993
rect 659 2988 664 2993
rect 726 2988 731 2993
rect 747 2988 752 2993
rect 777 2988 782 2993
rect 798 2988 803 2993
rect 865 2988 870 2993
rect 886 2988 891 2993
rect 916 2988 921 2993
rect 937 2988 942 2993
rect 1004 2988 1009 2993
rect 1025 2988 1030 2993
rect 1055 2988 1060 2993
rect 1076 2988 1081 2993
rect 1143 2988 1148 2993
rect 1164 2988 1169 2993
rect 1194 2988 1199 2993
rect 1215 2988 1220 2993
rect 1282 2988 1287 2993
rect 1303 2988 1308 2993
rect 1333 2988 1338 2993
rect 1354 2988 1359 2993
rect 1421 2988 1426 2993
rect 1442 2988 1447 2993
rect 1472 2988 1477 2993
rect 1493 2988 1498 2993
rect 1560 2988 1565 2993
rect 1581 2988 1586 2993
rect 1611 2988 1616 2993
rect 1632 2988 1637 2993
rect 1699 2988 1704 2993
rect 1720 2988 1725 2993
rect 1750 2988 1755 2993
rect 1771 2988 1776 2993
rect 1838 2988 1843 2993
rect 1859 2988 1864 2993
rect 1889 2988 1894 2993
rect 1910 2988 1915 2993
rect 1977 2988 1982 2993
rect 1998 2988 2003 2993
rect 2028 2988 2033 2993
rect 2049 2988 2054 2993
rect 2116 2988 2121 2993
rect 2137 2988 2142 2993
rect 2167 2988 2172 2993
rect 2188 2988 2193 2993
rect 2255 2988 2260 2993
rect 2276 2988 2281 2993
rect 2306 2988 2311 2993
rect 2327 2988 2332 2993
rect 2394 2988 2399 2993
rect 2415 2988 2420 2993
rect 2445 2988 2450 2993
rect 2466 2988 2471 2993
rect 2533 2988 2538 2993
rect 2554 2988 2559 2993
rect 2584 2988 2589 2993
rect 2605 2988 2610 2993
rect 2672 2988 2677 2993
rect 2693 2988 2698 2993
rect 2723 2988 2728 2993
rect 2744 2988 2749 2993
rect 2811 2988 2816 2993
rect 2832 2988 2837 2993
rect 2862 2988 2867 2993
rect 2883 2988 2888 2993
rect 2950 2988 2955 2993
rect 2971 2988 2976 2993
rect 3001 2988 3006 2993
rect 3022 2988 3027 2993
rect 3089 2988 3094 2993
rect 3110 2988 3115 2993
rect 3140 2988 3145 2993
rect 3161 2988 3166 2993
rect 3228 2988 3233 2993
rect 3249 2988 3254 2993
rect 3279 2988 3284 2993
rect 3300 2988 3305 2993
rect 3367 2988 3372 2993
rect 3388 2988 3393 2993
rect 3418 2988 3423 2993
rect 3439 2988 3444 2993
rect 3506 2988 3511 2993
rect 3527 2988 3532 2993
rect 3557 2988 3562 2993
rect 3578 2988 3583 2993
rect 3645 2988 3650 2993
rect 3666 2988 3671 2993
rect 3696 2988 3701 2993
rect 3717 2988 3722 2993
rect 3784 2988 3789 2993
rect 3805 2988 3810 2993
rect 3835 2988 3840 2993
rect 3856 2988 3861 2993
rect 3923 2988 3928 2993
rect 3944 2988 3949 2993
rect 3974 2988 3979 2993
rect 3995 2988 4000 2993
rect 4062 2988 4067 2993
rect 4083 2988 4088 2993
rect -57 -2993 -52 -2988
rect -36 -2993 -31 -2988
rect 31 -2993 36 -2988
rect 52 -2993 57 -2988
rect 82 -2993 87 -2988
rect 103 -2993 108 -2988
rect 170 -2993 175 -2988
rect 191 -2993 196 -2988
rect 221 -2993 226 -2988
rect 242 -2993 247 -2988
rect 309 -2993 314 -2988
rect 330 -2993 335 -2988
rect 360 -2993 365 -2988
rect 381 -2993 386 -2988
rect 448 -2993 453 -2988
rect 469 -2993 474 -2988
rect 499 -2993 504 -2988
rect 520 -2993 525 -2988
rect 587 -2993 592 -2988
rect 608 -2993 613 -2988
rect 638 -2993 643 -2988
rect 659 -2993 664 -2988
rect 726 -2993 731 -2988
rect 747 -2993 752 -2988
rect 777 -2993 782 -2988
rect 798 -2993 803 -2988
rect 865 -2993 870 -2988
rect 886 -2993 891 -2988
rect 916 -2993 921 -2988
rect 937 -2993 942 -2988
rect 1004 -2993 1009 -2988
rect 1025 -2993 1030 -2988
rect 1055 -2993 1060 -2988
rect 1076 -2993 1081 -2988
rect 1143 -2993 1148 -2988
rect 1164 -2993 1169 -2988
rect 1194 -2993 1199 -2988
rect 1215 -2993 1220 -2988
rect 1282 -2993 1287 -2988
rect 1303 -2993 1308 -2988
rect 1333 -2993 1338 -2988
rect 1354 -2993 1359 -2988
rect 1421 -2993 1426 -2988
rect 1442 -2993 1447 -2988
rect 1472 -2993 1477 -2988
rect 1493 -2993 1498 -2988
rect 1560 -2993 1565 -2988
rect 1581 -2993 1586 -2988
rect 1611 -2993 1616 -2988
rect 1632 -2993 1637 -2988
rect 1699 -2993 1704 -2988
rect 1720 -2993 1725 -2988
rect 1750 -2993 1755 -2988
rect 1771 -2993 1776 -2988
rect 1838 -2993 1843 -2988
rect 1859 -2993 1864 -2988
rect 1889 -2993 1894 -2988
rect 1910 -2993 1915 -2988
rect 1977 -2993 1982 -2988
rect 1998 -2993 2003 -2988
rect 2028 -2993 2033 -2988
rect 2049 -2993 2054 -2988
rect 2116 -2993 2121 -2988
rect 2137 -2993 2142 -2988
rect 2167 -2993 2172 -2988
rect 2188 -2993 2193 -2988
rect 2255 -2993 2260 -2988
rect 2276 -2993 2281 -2988
rect 2306 -2993 2311 -2988
rect 2327 -2993 2332 -2988
rect 2394 -2993 2399 -2988
rect 2415 -2993 2420 -2988
rect 2445 -2993 2450 -2988
rect 2466 -2993 2471 -2988
rect 2533 -2993 2538 -2988
rect 2554 -2993 2559 -2988
rect 2584 -2993 2589 -2988
rect 2605 -2993 2610 -2988
rect 2672 -2993 2677 -2988
rect 2693 -2993 2698 -2988
rect 2723 -2993 2728 -2988
rect 2744 -2993 2749 -2988
rect 2811 -2993 2816 -2988
rect 2832 -2993 2837 -2988
rect 2862 -2993 2867 -2988
rect 2883 -2993 2888 -2988
rect 2950 -2993 2955 -2988
rect 2971 -2993 2976 -2988
rect 3001 -2993 3006 -2988
rect 3022 -2993 3027 -2988
rect 3089 -2993 3094 -2988
rect 3110 -2993 3115 -2988
rect 3140 -2993 3145 -2988
rect 3161 -2993 3166 -2988
rect 3228 -2993 3233 -2988
rect 3249 -2993 3254 -2988
rect 3279 -2993 3284 -2988
rect 3300 -2993 3305 -2988
rect 3367 -2993 3372 -2988
rect 3388 -2993 3393 -2988
rect 3418 -2993 3423 -2988
rect 3439 -2993 3444 -2988
rect 3506 -2993 3511 -2988
rect 3527 -2993 3532 -2988
rect 3557 -2993 3562 -2988
rect 3578 -2993 3583 -2988
rect 3645 -2993 3650 -2988
rect 3666 -2993 3671 -2988
rect 3696 -2993 3701 -2988
rect 3717 -2993 3722 -2988
rect 3784 -2993 3789 -2988
rect 3805 -2993 3810 -2988
rect 3835 -2993 3840 -2988
rect 3856 -2993 3861 -2988
rect 3923 -2993 3928 -2988
rect 3944 -2993 3949 -2988
rect 3974 -2993 3979 -2988
rect 3995 -2993 4000 -2988
rect 4062 -2993 4067 -2988
rect 4083 -2993 4088 -2988
rect -52 -2998 -47 -2993
rect -41 -2998 -36 -2993
rect 36 -2998 41 -2993
rect 47 -2998 52 -2993
rect 87 -2998 92 -2993
rect 98 -2998 103 -2993
rect 175 -2998 180 -2993
rect 186 -2998 191 -2993
rect 226 -2998 231 -2993
rect 237 -2998 242 -2993
rect 314 -2998 319 -2993
rect 325 -2998 330 -2993
rect 365 -2998 370 -2993
rect 376 -2998 381 -2993
rect 453 -2998 458 -2993
rect 464 -2998 469 -2993
rect 504 -2998 509 -2993
rect 515 -2998 520 -2993
rect 592 -2998 597 -2993
rect 603 -2998 608 -2993
rect 643 -2998 648 -2993
rect 654 -2998 659 -2993
rect 731 -2998 736 -2993
rect 742 -2998 747 -2993
rect 782 -2998 787 -2993
rect 793 -2998 798 -2993
rect 870 -2998 875 -2993
rect 881 -2998 886 -2993
rect 921 -2998 926 -2993
rect 932 -2998 937 -2993
rect 1009 -2998 1014 -2993
rect 1020 -2998 1025 -2993
rect 1060 -2998 1065 -2993
rect 1071 -2998 1076 -2993
rect 1148 -2998 1153 -2993
rect 1159 -2998 1164 -2993
rect 1199 -2998 1204 -2993
rect 1210 -2998 1215 -2993
rect 1287 -2998 1292 -2993
rect 1298 -2998 1303 -2993
rect 1338 -2998 1343 -2993
rect 1349 -2998 1354 -2993
rect 1426 -2998 1431 -2993
rect 1437 -2998 1442 -2993
rect 1477 -2998 1482 -2993
rect 1488 -2998 1493 -2993
rect 1565 -2998 1570 -2993
rect 1576 -2998 1581 -2993
rect 1616 -2998 1621 -2993
rect 1627 -2998 1632 -2993
rect 1704 -2998 1709 -2993
rect 1715 -2998 1720 -2993
rect 1755 -2998 1760 -2993
rect 1766 -2998 1771 -2993
rect 1843 -2998 1848 -2993
rect 1854 -2998 1859 -2993
rect 1894 -2998 1899 -2993
rect 1905 -2998 1910 -2993
rect 1982 -2998 1987 -2993
rect 1993 -2998 1998 -2993
rect 2033 -2998 2038 -2993
rect 2044 -2998 2049 -2993
rect 2121 -2998 2126 -2993
rect 2132 -2998 2137 -2993
rect 2172 -2998 2177 -2993
rect 2183 -2998 2188 -2993
rect 2260 -2998 2265 -2993
rect 2271 -2998 2276 -2993
rect 2311 -2998 2316 -2993
rect 2322 -2998 2327 -2993
rect 2399 -2998 2404 -2993
rect 2410 -2998 2415 -2993
rect 2450 -2998 2455 -2993
rect 2461 -2998 2466 -2993
rect 2538 -2998 2543 -2993
rect 2549 -2998 2554 -2993
rect 2589 -2998 2594 -2993
rect 2600 -2998 2605 -2993
rect 2677 -2998 2682 -2993
rect 2688 -2998 2693 -2993
rect 2728 -2998 2733 -2993
rect 2739 -2998 2744 -2993
rect 2816 -2998 2821 -2993
rect 2827 -2998 2832 -2993
rect 2867 -2998 2872 -2993
rect 2878 -2998 2883 -2993
rect 2955 -2998 2960 -2993
rect 2966 -2998 2971 -2993
rect 3006 -2998 3011 -2993
rect 3017 -2998 3022 -2993
rect 3094 -2998 3099 -2993
rect 3105 -2998 3110 -2993
rect 3145 -2998 3150 -2993
rect 3156 -2998 3161 -2993
rect 3233 -2998 3238 -2993
rect 3244 -2998 3249 -2993
rect 3284 -2998 3289 -2993
rect 3295 -2998 3300 -2993
rect 3372 -2998 3377 -2993
rect 3383 -2998 3388 -2993
rect 3423 -2998 3428 -2993
rect 3434 -2998 3439 -2993
rect 3511 -2998 3516 -2993
rect 3522 -2998 3527 -2993
rect 3562 -2998 3567 -2993
rect 3573 -2998 3578 -2993
rect 3650 -2998 3655 -2993
rect 3661 -2998 3666 -2993
rect 3701 -2998 3706 -2993
rect 3712 -2998 3717 -2993
rect 3789 -2998 3794 -2993
rect 3800 -2998 3805 -2993
rect 3840 -2998 3845 -2993
rect 3851 -2998 3856 -2993
rect 3928 -2998 3933 -2993
rect 3939 -2998 3944 -2993
rect 3979 -2998 3984 -2993
rect 3990 -2998 3995 -2993
rect 4067 -2998 4072 -2993
rect 4078 -2998 4083 -2993
rect -18 -3014 -13 -3009
rect 13 -3014 18 -3009
rect 121 -3014 126 -3009
rect 152 -3014 157 -3009
rect 260 -3014 265 -3009
rect 291 -3014 296 -3009
rect 399 -3014 404 -3009
rect 430 -3014 435 -3009
rect 538 -3014 543 -3009
rect 569 -3014 574 -3009
rect 677 -3014 682 -3009
rect 708 -3014 713 -3009
rect 816 -3014 821 -3009
rect 847 -3014 852 -3009
rect 955 -3014 960 -3009
rect 986 -3014 991 -3009
rect 1094 -3014 1099 -3009
rect 1125 -3014 1130 -3009
rect 1233 -3014 1238 -3009
rect 1264 -3014 1269 -3009
rect 1372 -3014 1377 -3009
rect 1403 -3014 1408 -3009
rect 1511 -3014 1516 -3009
rect 1542 -3014 1547 -3009
rect 1650 -3014 1655 -3009
rect 1681 -3014 1686 -3009
rect 1789 -3014 1794 -3009
rect 1820 -3014 1825 -3009
rect 1928 -3014 1933 -3009
rect 1959 -3014 1964 -3009
rect 2067 -3014 2072 -3009
rect 2098 -3014 2103 -3009
rect 2206 -3014 2211 -3009
rect 2237 -3014 2242 -3009
rect 2345 -3014 2350 -3009
rect 2376 -3014 2381 -3009
rect 2484 -3014 2489 -3009
rect 2515 -3014 2520 -3009
rect 2623 -3014 2628 -3009
rect 2654 -3014 2659 -3009
rect 2762 -3014 2767 -3009
rect 2793 -3014 2798 -3009
rect 2901 -3014 2906 -3009
rect 2932 -3014 2937 -3009
rect 3040 -3014 3045 -3009
rect 3071 -3014 3076 -3009
rect 3179 -3014 3184 -3009
rect 3210 -3014 3215 -3009
rect 3318 -3014 3323 -3009
rect 3349 -3014 3354 -3009
rect 3457 -3014 3462 -3009
rect 3488 -3014 3493 -3009
rect 3596 -3014 3601 -3009
rect 3627 -3014 3632 -3009
rect 3735 -3014 3740 -3009
rect 3766 -3014 3771 -3009
rect 3874 -3014 3879 -3009
rect 3905 -3014 3910 -3009
rect 4013 -3014 4018 -3009
rect 4044 -3014 4049 -3009
rect -23 -3019 23 -3014
rect 116 -3019 162 -3014
rect 255 -3019 301 -3014
rect 394 -3019 440 -3014
rect 533 -3019 579 -3014
rect 672 -3019 718 -3014
rect 811 -3019 857 -3014
rect 950 -3019 996 -3014
rect 1089 -3019 1135 -3014
rect 1228 -3019 1274 -3014
rect 1367 -3019 1413 -3014
rect 1506 -3019 1552 -3014
rect 1645 -3019 1691 -3014
rect 1784 -3019 1830 -3014
rect 1923 -3019 1969 -3014
rect 2062 -3019 2108 -3014
rect 2201 -3019 2247 -3014
rect 2340 -3019 2386 -3014
rect 2479 -3019 2525 -3014
rect 2618 -3019 2664 -3014
rect 2757 -3019 2803 -3014
rect 2896 -3019 2942 -3014
rect 3035 -3019 3081 -3014
rect 3174 -3019 3220 -3014
rect 3313 -3019 3359 -3014
rect 3452 -3019 3498 -3014
rect 3591 -3019 3637 -3014
rect 3730 -3019 3776 -3014
rect 3869 -3019 3915 -3014
rect 4008 -3019 4054 -3014
rect -18 -3025 18 -3019
rect 121 -3025 157 -3019
rect 260 -3025 296 -3019
rect 399 -3025 435 -3019
rect 538 -3025 574 -3019
rect 677 -3025 713 -3019
rect 816 -3025 852 -3019
rect 955 -3025 991 -3019
rect 1094 -3025 1130 -3019
rect 1233 -3025 1269 -3019
rect 1372 -3025 1408 -3019
rect 1511 -3025 1547 -3019
rect 1650 -3025 1686 -3019
rect 1789 -3025 1825 -3019
rect 1928 -3025 1964 -3019
rect 2067 -3025 2103 -3019
rect 2206 -3025 2242 -3019
rect 2345 -3025 2381 -3019
rect 2484 -3025 2520 -3019
rect 2623 -3025 2659 -3019
rect 2762 -3025 2798 -3019
rect 2901 -3025 2937 -3019
rect 3040 -3025 3076 -3019
rect 3179 -3025 3215 -3019
rect 3318 -3025 3354 -3019
rect 3457 -3025 3493 -3019
rect 3596 -3025 3632 -3019
rect 3735 -3025 3771 -3019
rect 3874 -3025 3910 -3019
rect 4013 -3025 4049 -3019
rect -23 -3030 23 -3025
rect 116 -3030 162 -3025
rect 255 -3030 301 -3025
rect 394 -3030 440 -3025
rect 533 -3030 579 -3025
rect 672 -3030 718 -3025
rect 811 -3030 857 -3025
rect 950 -3030 996 -3025
rect 1089 -3030 1135 -3025
rect 1228 -3030 1274 -3025
rect 1367 -3030 1413 -3025
rect 1506 -3030 1552 -3025
rect 1645 -3030 1691 -3025
rect 1784 -3030 1830 -3025
rect 1923 -3030 1969 -3025
rect 2062 -3030 2108 -3025
rect 2201 -3030 2247 -3025
rect 2340 -3030 2386 -3025
rect 2479 -3030 2525 -3025
rect 2618 -3030 2664 -3025
rect 2757 -3030 2803 -3025
rect 2896 -3030 2942 -3025
rect 3035 -3030 3081 -3025
rect 3174 -3030 3220 -3025
rect 3313 -3030 3359 -3025
rect 3452 -3030 3498 -3025
rect 3591 -3030 3637 -3025
rect 3730 -3030 3776 -3025
rect 3869 -3030 3915 -3025
rect 4008 -3030 4054 -3025
rect -18 -3035 -13 -3030
rect 13 -3035 18 -3030
rect 121 -3035 126 -3030
rect 152 -3035 157 -3030
rect 260 -3035 265 -3030
rect 291 -3035 296 -3030
rect 399 -3035 404 -3030
rect 430 -3035 435 -3030
rect 538 -3035 543 -3030
rect 569 -3035 574 -3030
rect 677 -3035 682 -3030
rect 708 -3035 713 -3030
rect 816 -3035 821 -3030
rect 847 -3035 852 -3030
rect 955 -3035 960 -3030
rect 986 -3035 991 -3030
rect 1094 -3035 1099 -3030
rect 1125 -3035 1130 -3030
rect 1233 -3035 1238 -3030
rect 1264 -3035 1269 -3030
rect 1372 -3035 1377 -3030
rect 1403 -3035 1408 -3030
rect 1511 -3035 1516 -3030
rect 1542 -3035 1547 -3030
rect 1650 -3035 1655 -3030
rect 1681 -3035 1686 -3030
rect 1789 -3035 1794 -3030
rect 1820 -3035 1825 -3030
rect 1928 -3035 1933 -3030
rect 1959 -3035 1964 -3030
rect 2067 -3035 2072 -3030
rect 2098 -3035 2103 -3030
rect 2206 -3035 2211 -3030
rect 2237 -3035 2242 -3030
rect 2345 -3035 2350 -3030
rect 2376 -3035 2381 -3030
rect 2484 -3035 2489 -3030
rect 2515 -3035 2520 -3030
rect 2623 -3035 2628 -3030
rect 2654 -3035 2659 -3030
rect 2762 -3035 2767 -3030
rect 2793 -3035 2798 -3030
rect 2901 -3035 2906 -3030
rect 2932 -3035 2937 -3030
rect 3040 -3035 3045 -3030
rect 3071 -3035 3076 -3030
rect 3179 -3035 3184 -3030
rect 3210 -3035 3215 -3030
rect 3318 -3035 3323 -3030
rect 3349 -3035 3354 -3030
rect 3457 -3035 3462 -3030
rect 3488 -3035 3493 -3030
rect 3596 -3035 3601 -3030
rect 3627 -3035 3632 -3030
rect 3735 -3035 3740 -3030
rect 3766 -3035 3771 -3030
rect 3874 -3035 3879 -3030
rect 3905 -3035 3910 -3030
rect 4013 -3035 4018 -3030
rect 4044 -3035 4049 -3030
<< nwell >>
rect -259 -3173 4290 3173
<< hvpmos >>
rect -25 -3000 25 3000
rect 114 -3000 164 3000
rect 253 -3000 303 3000
rect 392 -3000 442 3000
rect 531 -3000 581 3000
rect 670 -3000 720 3000
rect 809 -3000 859 3000
rect 948 -3000 998 3000
rect 1087 -3000 1137 3000
rect 1226 -3000 1276 3000
rect 1365 -3000 1415 3000
rect 1504 -3000 1554 3000
rect 1643 -3000 1693 3000
rect 1782 -3000 1832 3000
rect 1921 -3000 1971 3000
rect 2060 -3000 2110 3000
rect 2199 -3000 2249 3000
rect 2338 -3000 2388 3000
rect 2477 -3000 2527 3000
rect 2616 -3000 2666 3000
rect 2755 -3000 2805 3000
rect 2894 -3000 2944 3000
rect 3033 -3000 3083 3000
rect 3172 -3000 3222 3000
rect 3311 -3000 3361 3000
rect 3450 -3000 3500 3000
rect 3589 -3000 3639 3000
rect 3728 -3000 3778 3000
rect 3867 -3000 3917 3000
rect 4006 -3000 4056 3000
<< hvpdiff >>
rect -59 2993 -25 3000
rect -59 -2993 -52 2993
rect -36 -2993 -25 2993
rect -59 -3000 -25 -2993
rect 25 2993 59 3000
rect 25 -2993 36 2993
rect 52 -2993 59 2993
rect 25 -3000 59 -2993
rect 80 2993 114 3000
rect 80 -2993 87 2993
rect 103 -2993 114 2993
rect 80 -3000 114 -2993
rect 164 2993 198 3000
rect 164 -2993 175 2993
rect 191 -2993 198 2993
rect 164 -3000 198 -2993
rect 219 2993 253 3000
rect 219 -2993 226 2993
rect 242 -2993 253 2993
rect 219 -3000 253 -2993
rect 303 2993 337 3000
rect 303 -2993 314 2993
rect 330 -2993 337 2993
rect 303 -3000 337 -2993
rect 358 2993 392 3000
rect 358 -2993 365 2993
rect 381 -2993 392 2993
rect 358 -3000 392 -2993
rect 442 2993 476 3000
rect 442 -2993 453 2993
rect 469 -2993 476 2993
rect 442 -3000 476 -2993
rect 497 2993 531 3000
rect 497 -2993 504 2993
rect 520 -2993 531 2993
rect 497 -3000 531 -2993
rect 581 2993 615 3000
rect 581 -2993 592 2993
rect 608 -2993 615 2993
rect 581 -3000 615 -2993
rect 636 2993 670 3000
rect 636 -2993 643 2993
rect 659 -2993 670 2993
rect 636 -3000 670 -2993
rect 720 2993 754 3000
rect 720 -2993 731 2993
rect 747 -2993 754 2993
rect 720 -3000 754 -2993
rect 775 2993 809 3000
rect 775 -2993 782 2993
rect 798 -2993 809 2993
rect 775 -3000 809 -2993
rect 859 2993 893 3000
rect 859 -2993 870 2993
rect 886 -2993 893 2993
rect 859 -3000 893 -2993
rect 914 2993 948 3000
rect 914 -2993 921 2993
rect 937 -2993 948 2993
rect 914 -3000 948 -2993
rect 998 2993 1032 3000
rect 998 -2993 1009 2993
rect 1025 -2993 1032 2993
rect 998 -3000 1032 -2993
rect 1053 2993 1087 3000
rect 1053 -2993 1060 2993
rect 1076 -2993 1087 2993
rect 1053 -3000 1087 -2993
rect 1137 2993 1171 3000
rect 1137 -2993 1148 2993
rect 1164 -2993 1171 2993
rect 1137 -3000 1171 -2993
rect 1192 2993 1226 3000
rect 1192 -2993 1199 2993
rect 1215 -2993 1226 2993
rect 1192 -3000 1226 -2993
rect 1276 2993 1310 3000
rect 1276 -2993 1287 2993
rect 1303 -2993 1310 2993
rect 1276 -3000 1310 -2993
rect 1331 2993 1365 3000
rect 1331 -2993 1338 2993
rect 1354 -2993 1365 2993
rect 1331 -3000 1365 -2993
rect 1415 2993 1449 3000
rect 1415 -2993 1426 2993
rect 1442 -2993 1449 2993
rect 1415 -3000 1449 -2993
rect 1470 2993 1504 3000
rect 1470 -2993 1477 2993
rect 1493 -2993 1504 2993
rect 1470 -3000 1504 -2993
rect 1554 2993 1588 3000
rect 1554 -2993 1565 2993
rect 1581 -2993 1588 2993
rect 1554 -3000 1588 -2993
rect 1609 2993 1643 3000
rect 1609 -2993 1616 2993
rect 1632 -2993 1643 2993
rect 1609 -3000 1643 -2993
rect 1693 2993 1727 3000
rect 1693 -2993 1704 2993
rect 1720 -2993 1727 2993
rect 1693 -3000 1727 -2993
rect 1748 2993 1782 3000
rect 1748 -2993 1755 2993
rect 1771 -2993 1782 2993
rect 1748 -3000 1782 -2993
rect 1832 2993 1866 3000
rect 1832 -2993 1843 2993
rect 1859 -2993 1866 2993
rect 1832 -3000 1866 -2993
rect 1887 2993 1921 3000
rect 1887 -2993 1894 2993
rect 1910 -2993 1921 2993
rect 1887 -3000 1921 -2993
rect 1971 2993 2005 3000
rect 1971 -2993 1982 2993
rect 1998 -2993 2005 2993
rect 1971 -3000 2005 -2993
rect 2026 2993 2060 3000
rect 2026 -2993 2033 2993
rect 2049 -2993 2060 2993
rect 2026 -3000 2060 -2993
rect 2110 2993 2144 3000
rect 2110 -2993 2121 2993
rect 2137 -2993 2144 2993
rect 2110 -3000 2144 -2993
rect 2165 2993 2199 3000
rect 2165 -2993 2172 2993
rect 2188 -2993 2199 2993
rect 2165 -3000 2199 -2993
rect 2249 2993 2283 3000
rect 2249 -2993 2260 2993
rect 2276 -2993 2283 2993
rect 2249 -3000 2283 -2993
rect 2304 2993 2338 3000
rect 2304 -2993 2311 2993
rect 2327 -2993 2338 2993
rect 2304 -3000 2338 -2993
rect 2388 2993 2422 3000
rect 2388 -2993 2399 2993
rect 2415 -2993 2422 2993
rect 2388 -3000 2422 -2993
rect 2443 2993 2477 3000
rect 2443 -2993 2450 2993
rect 2466 -2993 2477 2993
rect 2443 -3000 2477 -2993
rect 2527 2993 2561 3000
rect 2527 -2993 2538 2993
rect 2554 -2993 2561 2993
rect 2527 -3000 2561 -2993
rect 2582 2993 2616 3000
rect 2582 -2993 2589 2993
rect 2605 -2993 2616 2993
rect 2582 -3000 2616 -2993
rect 2666 2993 2700 3000
rect 2666 -2993 2677 2993
rect 2693 -2993 2700 2993
rect 2666 -3000 2700 -2993
rect 2721 2993 2755 3000
rect 2721 -2993 2728 2993
rect 2744 -2993 2755 2993
rect 2721 -3000 2755 -2993
rect 2805 2993 2839 3000
rect 2805 -2993 2816 2993
rect 2832 -2993 2839 2993
rect 2805 -3000 2839 -2993
rect 2860 2993 2894 3000
rect 2860 -2993 2867 2993
rect 2883 -2993 2894 2993
rect 2860 -3000 2894 -2993
rect 2944 2993 2978 3000
rect 2944 -2993 2955 2993
rect 2971 -2993 2978 2993
rect 2944 -3000 2978 -2993
rect 2999 2993 3033 3000
rect 2999 -2993 3006 2993
rect 3022 -2993 3033 2993
rect 2999 -3000 3033 -2993
rect 3083 2993 3117 3000
rect 3083 -2993 3094 2993
rect 3110 -2993 3117 2993
rect 3083 -3000 3117 -2993
rect 3138 2993 3172 3000
rect 3138 -2993 3145 2993
rect 3161 -2993 3172 2993
rect 3138 -3000 3172 -2993
rect 3222 2993 3256 3000
rect 3222 -2993 3233 2993
rect 3249 -2993 3256 2993
rect 3222 -3000 3256 -2993
rect 3277 2993 3311 3000
rect 3277 -2993 3284 2993
rect 3300 -2993 3311 2993
rect 3277 -3000 3311 -2993
rect 3361 2993 3395 3000
rect 3361 -2993 3372 2993
rect 3388 -2993 3395 2993
rect 3361 -3000 3395 -2993
rect 3416 2993 3450 3000
rect 3416 -2993 3423 2993
rect 3439 -2993 3450 2993
rect 3416 -3000 3450 -2993
rect 3500 2993 3534 3000
rect 3500 -2993 3511 2993
rect 3527 -2993 3534 2993
rect 3500 -3000 3534 -2993
rect 3555 2993 3589 3000
rect 3555 -2993 3562 2993
rect 3578 -2993 3589 2993
rect 3555 -3000 3589 -2993
rect 3639 2993 3673 3000
rect 3639 -2993 3650 2993
rect 3666 -2993 3673 2993
rect 3639 -3000 3673 -2993
rect 3694 2993 3728 3000
rect 3694 -2993 3701 2993
rect 3717 -2993 3728 2993
rect 3694 -3000 3728 -2993
rect 3778 2993 3812 3000
rect 3778 -2993 3789 2993
rect 3805 -2993 3812 2993
rect 3778 -3000 3812 -2993
rect 3833 2993 3867 3000
rect 3833 -2993 3840 2993
rect 3856 -2993 3867 2993
rect 3833 -3000 3867 -2993
rect 3917 2993 3951 3000
rect 3917 -2993 3928 2993
rect 3944 -2993 3951 2993
rect 3917 -3000 3951 -2993
rect 3972 2993 4006 3000
rect 3972 -2993 3979 2993
rect 3995 -2993 4006 2993
rect 3972 -3000 4006 -2993
rect 4056 2993 4090 3000
rect 4056 -2993 4067 2993
rect 4083 -2993 4090 2993
rect 4056 -3000 4090 -2993
<< hvpdiffc >>
rect -52 -2993 -36 2993
rect 36 -2993 52 2993
rect 87 -2993 103 2993
rect 175 -2993 191 2993
rect 226 -2993 242 2993
rect 314 -2993 330 2993
rect 365 -2993 381 2993
rect 453 -2993 469 2993
rect 504 -2993 520 2993
rect 592 -2993 608 2993
rect 643 -2993 659 2993
rect 731 -2993 747 2993
rect 782 -2993 798 2993
rect 870 -2993 886 2993
rect 921 -2993 937 2993
rect 1009 -2993 1025 2993
rect 1060 -2993 1076 2993
rect 1148 -2993 1164 2993
rect 1199 -2993 1215 2993
rect 1287 -2993 1303 2993
rect 1338 -2993 1354 2993
rect 1426 -2993 1442 2993
rect 1477 -2993 1493 2993
rect 1565 -2993 1581 2993
rect 1616 -2993 1632 2993
rect 1704 -2993 1720 2993
rect 1755 -2993 1771 2993
rect 1843 -2993 1859 2993
rect 1894 -2993 1910 2993
rect 1982 -2993 1998 2993
rect 2033 -2993 2049 2993
rect 2121 -2993 2137 2993
rect 2172 -2993 2188 2993
rect 2260 -2993 2276 2993
rect 2311 -2993 2327 2993
rect 2399 -2993 2415 2993
rect 2450 -2993 2466 2993
rect 2538 -2993 2554 2993
rect 2589 -2993 2605 2993
rect 2677 -2993 2693 2993
rect 2728 -2993 2744 2993
rect 2816 -2993 2832 2993
rect 2867 -2993 2883 2993
rect 2955 -2993 2971 2993
rect 3006 -2993 3022 2993
rect 3094 -2993 3110 2993
rect 3145 -2993 3161 2993
rect 3233 -2993 3249 2993
rect 3284 -2993 3300 2993
rect 3372 -2993 3388 2993
rect 3423 -2993 3439 2993
rect 3511 -2993 3527 2993
rect 3562 -2993 3578 2993
rect 3650 -2993 3666 2993
rect 3701 -2993 3717 2993
rect 3789 -2993 3805 2993
rect 3840 -2993 3856 2993
rect 3928 -2993 3944 2993
rect 3979 -2993 3995 2993
rect 4067 -2993 4083 2993
<< nsubdiff >>
rect -197 3104 4228 3111
rect -197 3088 -160 3104
rect 4191 3088 4228 3104
rect -197 3081 4228 3088
rect -197 3074 -167 3081
rect -197 -3074 -190 3074
rect -174 -3074 -167 3074
rect 4198 3074 4228 3081
rect -197 -3081 -167 -3074
rect 4198 -3074 4205 3074
rect 4221 -3074 4228 3074
rect 4198 -3081 4228 -3074
rect -197 -3088 4228 -3081
rect -197 -3104 -160 -3088
rect 4191 -3104 4228 -3088
rect -197 -3111 4228 -3104
<< nsubdiffcont >>
rect -160 3088 4191 3104
rect -190 -3074 -174 3074
rect 4205 -3074 4221 3074
rect -160 -3104 4191 -3088
<< poly >>
rect -25 3030 25 3037
rect -25 3014 -18 3030
rect 18 3014 25 3030
rect -25 3000 25 3014
rect 114 3030 164 3037
rect 114 3014 121 3030
rect 157 3014 164 3030
rect 114 3000 164 3014
rect 253 3030 303 3037
rect 253 3014 260 3030
rect 296 3014 303 3030
rect 253 3000 303 3014
rect 392 3030 442 3037
rect 392 3014 399 3030
rect 435 3014 442 3030
rect 392 3000 442 3014
rect 531 3030 581 3037
rect 531 3014 538 3030
rect 574 3014 581 3030
rect 531 3000 581 3014
rect 670 3030 720 3037
rect 670 3014 677 3030
rect 713 3014 720 3030
rect 670 3000 720 3014
rect 809 3030 859 3037
rect 809 3014 816 3030
rect 852 3014 859 3030
rect 809 3000 859 3014
rect 948 3030 998 3037
rect 948 3014 955 3030
rect 991 3014 998 3030
rect 948 3000 998 3014
rect 1087 3030 1137 3037
rect 1087 3014 1094 3030
rect 1130 3014 1137 3030
rect 1087 3000 1137 3014
rect 1226 3030 1276 3037
rect 1226 3014 1233 3030
rect 1269 3014 1276 3030
rect 1226 3000 1276 3014
rect 1365 3030 1415 3037
rect 1365 3014 1372 3030
rect 1408 3014 1415 3030
rect 1365 3000 1415 3014
rect 1504 3030 1554 3037
rect 1504 3014 1511 3030
rect 1547 3014 1554 3030
rect 1504 3000 1554 3014
rect 1643 3030 1693 3037
rect 1643 3014 1650 3030
rect 1686 3014 1693 3030
rect 1643 3000 1693 3014
rect 1782 3030 1832 3037
rect 1782 3014 1789 3030
rect 1825 3014 1832 3030
rect 1782 3000 1832 3014
rect 1921 3030 1971 3037
rect 1921 3014 1928 3030
rect 1964 3014 1971 3030
rect 1921 3000 1971 3014
rect 2060 3030 2110 3037
rect 2060 3014 2067 3030
rect 2103 3014 2110 3030
rect 2060 3000 2110 3014
rect 2199 3030 2249 3037
rect 2199 3014 2206 3030
rect 2242 3014 2249 3030
rect 2199 3000 2249 3014
rect 2338 3030 2388 3037
rect 2338 3014 2345 3030
rect 2381 3014 2388 3030
rect 2338 3000 2388 3014
rect 2477 3030 2527 3037
rect 2477 3014 2484 3030
rect 2520 3014 2527 3030
rect 2477 3000 2527 3014
rect 2616 3030 2666 3037
rect 2616 3014 2623 3030
rect 2659 3014 2666 3030
rect 2616 3000 2666 3014
rect 2755 3030 2805 3037
rect 2755 3014 2762 3030
rect 2798 3014 2805 3030
rect 2755 3000 2805 3014
rect 2894 3030 2944 3037
rect 2894 3014 2901 3030
rect 2937 3014 2944 3030
rect 2894 3000 2944 3014
rect 3033 3030 3083 3037
rect 3033 3014 3040 3030
rect 3076 3014 3083 3030
rect 3033 3000 3083 3014
rect 3172 3030 3222 3037
rect 3172 3014 3179 3030
rect 3215 3014 3222 3030
rect 3172 3000 3222 3014
rect 3311 3030 3361 3037
rect 3311 3014 3318 3030
rect 3354 3014 3361 3030
rect 3311 3000 3361 3014
rect 3450 3030 3500 3037
rect 3450 3014 3457 3030
rect 3493 3014 3500 3030
rect 3450 3000 3500 3014
rect 3589 3030 3639 3037
rect 3589 3014 3596 3030
rect 3632 3014 3639 3030
rect 3589 3000 3639 3014
rect 3728 3030 3778 3037
rect 3728 3014 3735 3030
rect 3771 3014 3778 3030
rect 3728 3000 3778 3014
rect 3867 3030 3917 3037
rect 3867 3014 3874 3030
rect 3910 3014 3917 3030
rect 3867 3000 3917 3014
rect 4006 3030 4056 3037
rect 4006 3014 4013 3030
rect 4049 3014 4056 3030
rect 4006 3000 4056 3014
rect -25 -3014 25 -3000
rect -25 -3030 -18 -3014
rect 18 -3030 25 -3014
rect -25 -3037 25 -3030
rect 114 -3014 164 -3000
rect 114 -3030 121 -3014
rect 157 -3030 164 -3014
rect 114 -3037 164 -3030
rect 253 -3014 303 -3000
rect 253 -3030 260 -3014
rect 296 -3030 303 -3014
rect 253 -3037 303 -3030
rect 392 -3014 442 -3000
rect 392 -3030 399 -3014
rect 435 -3030 442 -3014
rect 392 -3037 442 -3030
rect 531 -3014 581 -3000
rect 531 -3030 538 -3014
rect 574 -3030 581 -3014
rect 531 -3037 581 -3030
rect 670 -3014 720 -3000
rect 670 -3030 677 -3014
rect 713 -3030 720 -3014
rect 670 -3037 720 -3030
rect 809 -3014 859 -3000
rect 809 -3030 816 -3014
rect 852 -3030 859 -3014
rect 809 -3037 859 -3030
rect 948 -3014 998 -3000
rect 948 -3030 955 -3014
rect 991 -3030 998 -3014
rect 948 -3037 998 -3030
rect 1087 -3014 1137 -3000
rect 1087 -3030 1094 -3014
rect 1130 -3030 1137 -3014
rect 1087 -3037 1137 -3030
rect 1226 -3014 1276 -3000
rect 1226 -3030 1233 -3014
rect 1269 -3030 1276 -3014
rect 1226 -3037 1276 -3030
rect 1365 -3014 1415 -3000
rect 1365 -3030 1372 -3014
rect 1408 -3030 1415 -3014
rect 1365 -3037 1415 -3030
rect 1504 -3014 1554 -3000
rect 1504 -3030 1511 -3014
rect 1547 -3030 1554 -3014
rect 1504 -3037 1554 -3030
rect 1643 -3014 1693 -3000
rect 1643 -3030 1650 -3014
rect 1686 -3030 1693 -3014
rect 1643 -3037 1693 -3030
rect 1782 -3014 1832 -3000
rect 1782 -3030 1789 -3014
rect 1825 -3030 1832 -3014
rect 1782 -3037 1832 -3030
rect 1921 -3014 1971 -3000
rect 1921 -3030 1928 -3014
rect 1964 -3030 1971 -3014
rect 1921 -3037 1971 -3030
rect 2060 -3014 2110 -3000
rect 2060 -3030 2067 -3014
rect 2103 -3030 2110 -3014
rect 2060 -3037 2110 -3030
rect 2199 -3014 2249 -3000
rect 2199 -3030 2206 -3014
rect 2242 -3030 2249 -3014
rect 2199 -3037 2249 -3030
rect 2338 -3014 2388 -3000
rect 2338 -3030 2345 -3014
rect 2381 -3030 2388 -3014
rect 2338 -3037 2388 -3030
rect 2477 -3014 2527 -3000
rect 2477 -3030 2484 -3014
rect 2520 -3030 2527 -3014
rect 2477 -3037 2527 -3030
rect 2616 -3014 2666 -3000
rect 2616 -3030 2623 -3014
rect 2659 -3030 2666 -3014
rect 2616 -3037 2666 -3030
rect 2755 -3014 2805 -3000
rect 2755 -3030 2762 -3014
rect 2798 -3030 2805 -3014
rect 2755 -3037 2805 -3030
rect 2894 -3014 2944 -3000
rect 2894 -3030 2901 -3014
rect 2937 -3030 2944 -3014
rect 2894 -3037 2944 -3030
rect 3033 -3014 3083 -3000
rect 3033 -3030 3040 -3014
rect 3076 -3030 3083 -3014
rect 3033 -3037 3083 -3030
rect 3172 -3014 3222 -3000
rect 3172 -3030 3179 -3014
rect 3215 -3030 3222 -3014
rect 3172 -3037 3222 -3030
rect 3311 -3014 3361 -3000
rect 3311 -3030 3318 -3014
rect 3354 -3030 3361 -3014
rect 3311 -3037 3361 -3030
rect 3450 -3014 3500 -3000
rect 3450 -3030 3457 -3014
rect 3493 -3030 3500 -3014
rect 3450 -3037 3500 -3030
rect 3589 -3014 3639 -3000
rect 3589 -3030 3596 -3014
rect 3632 -3030 3639 -3014
rect 3589 -3037 3639 -3030
rect 3728 -3014 3778 -3000
rect 3728 -3030 3735 -3014
rect 3771 -3030 3778 -3014
rect 3728 -3037 3778 -3030
rect 3867 -3014 3917 -3000
rect 3867 -3030 3874 -3014
rect 3910 -3030 3917 -3014
rect 3867 -3037 3917 -3030
rect 4006 -3014 4056 -3000
rect 4006 -3030 4013 -3014
rect 4049 -3030 4056 -3014
rect 4006 -3037 4056 -3030
<< polycont >>
rect -18 3014 18 3030
rect 121 3014 157 3030
rect 260 3014 296 3030
rect 399 3014 435 3030
rect 538 3014 574 3030
rect 677 3014 713 3030
rect 816 3014 852 3030
rect 955 3014 991 3030
rect 1094 3014 1130 3030
rect 1233 3014 1269 3030
rect 1372 3014 1408 3030
rect 1511 3014 1547 3030
rect 1650 3014 1686 3030
rect 1789 3014 1825 3030
rect 1928 3014 1964 3030
rect 2067 3014 2103 3030
rect 2206 3014 2242 3030
rect 2345 3014 2381 3030
rect 2484 3014 2520 3030
rect 2623 3014 2659 3030
rect 2762 3014 2798 3030
rect 2901 3014 2937 3030
rect 3040 3014 3076 3030
rect 3179 3014 3215 3030
rect 3318 3014 3354 3030
rect 3457 3014 3493 3030
rect 3596 3014 3632 3030
rect 3735 3014 3771 3030
rect 3874 3014 3910 3030
rect 4013 3014 4049 3030
rect -18 -3030 18 -3014
rect 121 -3030 157 -3014
rect 260 -3030 296 -3014
rect 399 -3030 435 -3014
rect 538 -3030 574 -3014
rect 677 -3030 713 -3014
rect 816 -3030 852 -3014
rect 955 -3030 991 -3014
rect 1094 -3030 1130 -3014
rect 1233 -3030 1269 -3014
rect 1372 -3030 1408 -3014
rect 1511 -3030 1547 -3014
rect 1650 -3030 1686 -3014
rect 1789 -3030 1825 -3014
rect 1928 -3030 1964 -3014
rect 2067 -3030 2103 -3014
rect 2206 -3030 2242 -3014
rect 2345 -3030 2381 -3014
rect 2484 -3030 2520 -3014
rect 2623 -3030 2659 -3014
rect 2762 -3030 2798 -3014
rect 2901 -3030 2937 -3014
rect 3040 -3030 3076 -3014
rect 3179 -3030 3215 -3014
rect 3318 -3030 3354 -3014
rect 3457 -3030 3493 -3014
rect 3596 -3030 3632 -3014
rect 3735 -3030 3771 -3014
rect 3874 -3030 3910 -3014
rect 4013 -3030 4049 -3014
<< metal1 >>
rect -195 3104 4226 3109
rect -195 3088 -160 3104
rect 4191 3088 4226 3104
rect -195 3083 4226 3088
rect -195 3074 -169 3083
rect -195 -3074 -190 3074
rect -174 -3074 -169 3074
rect 4200 3074 4226 3083
rect -195 -3083 -169 -3074
rect 4200 -3074 4205 3074
rect 4221 -3074 4226 3074
rect 4200 -3083 4226 -3074
rect -195 -3088 4226 -3083
rect -195 -3104 -160 -3088
rect 4191 -3104 4226 -3088
rect -195 -3109 4226 -3104
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 60 l 0.5 nf 1 nx 30 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 2 glc 1 grc 1 gtc 1 gbc 1
<< end >>
