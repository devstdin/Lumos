magic
tech ihp-sg13g2
magscale 1 2
timestamp 1748629122
<< nwell >>
rect -803 776 -712 883
rect -3434 775 -712 776
rect -3456 725 -712 775
<< metal1 >>
rect -6389 2975 1480 3287
rect -6389 1678 -6186 2975
rect -5935 2855 -4935 2921
rect -5935 2845 -5863 2855
rect -5579 2845 -5507 2855
rect -5223 2845 -5151 2855
rect -6041 1841 -5961 2813
rect -6075 1796 -6003 1841
rect -5915 1809 -5883 2845
rect -5837 1841 -5757 2813
rect -5685 1841 -5605 2813
rect -6075 1747 -6065 1796
rect -6013 1747 -6003 1796
rect -5935 1757 -5863 1809
rect -6075 1737 -6003 1747
rect -5795 1678 -5757 1841
rect -5719 1796 -5647 1841
rect -5559 1809 -5527 2845
rect -5481 1841 -5401 2813
rect -5329 1841 -5249 2813
rect -5719 1747 -5709 1796
rect -5657 1747 -5647 1796
rect -5579 1757 -5507 1809
rect -5719 1737 -5647 1747
rect -5439 1678 -5401 1841
rect -5363 1796 -5291 1841
rect -5203 1809 -5171 2845
rect -4973 2813 -4935 2855
rect -4867 2845 -4795 2897
rect -4511 2845 -4439 2897
rect -4155 2845 -4083 2897
rect -3799 2845 -3727 2897
rect -5125 1841 -5045 2813
rect -4973 2545 -4893 2813
rect -4973 2465 -4963 2545
rect -4903 2465 -4893 2545
rect -4973 1841 -4893 2465
rect -5363 1747 -5353 1796
rect -5301 1747 -5291 1796
rect -5223 1757 -5151 1809
rect -5363 1737 -5291 1747
rect -5083 1678 -5045 1841
rect -4847 1809 -4815 2845
rect -4769 2188 -4689 2813
rect -4769 2108 -4759 2188
rect -4699 2108 -4689 2188
rect -4769 1841 -4689 2108
rect -4617 2545 -4537 2813
rect -4617 2465 -4607 2545
rect -4547 2465 -4537 2545
rect -4617 1841 -4537 2465
rect -4491 1809 -4459 2845
rect -4413 2188 -4333 2813
rect -4413 2108 -4403 2188
rect -4343 2108 -4333 2188
rect -4413 1841 -4333 2108
rect -4261 2545 -4181 2813
rect -4261 2465 -4251 2545
rect -4191 2465 -4181 2545
rect -4261 1841 -4181 2465
rect -4135 1809 -4103 2845
rect -4057 2188 -3977 2813
rect -4057 2108 -4047 2188
rect -3987 2108 -3977 2188
rect -4057 1841 -3977 2108
rect -3905 2545 -3825 2813
rect -3905 2465 -3895 2545
rect -3835 2465 -3825 2545
rect -3905 1841 -3825 2465
rect -3779 1809 -3747 2845
rect -3701 2188 -3621 2813
rect -3701 2108 -3691 2188
rect -3631 2108 -3621 2188
rect -3701 1841 -3621 2108
rect -4867 1796 -4795 1809
rect -4867 1731 -4857 1796
rect -4805 1731 -4795 1796
rect -4867 1721 -4795 1731
rect -4511 1796 -4439 1809
rect -4511 1731 -4501 1796
rect -4449 1731 -4439 1796
rect -4511 1721 -4439 1731
rect -4155 1796 -4083 1809
rect -4155 1731 -4145 1796
rect -4093 1731 -4083 1796
rect -4155 1721 -4083 1731
rect -3799 1796 -3727 1809
rect -3799 1731 -3789 1796
rect -3737 1731 -3727 1796
rect -3799 1721 -3727 1731
rect -3479 1683 -3281 2975
rect -3082 2867 -2710 2919
rect -4378 1678 -3281 1683
rect -6389 1556 -3281 1678
rect -6389 1447 -4139 1457
rect -6389 1367 -4229 1447
rect -4149 1367 -4139 1447
rect -6389 1357 -4139 1367
rect -6389 1333 -4239 1357
rect -6389 482 -5979 1333
rect -5845 1271 -5753 1281
rect -5845 1158 -5835 1271
rect -5763 1158 -5753 1271
rect -5845 1148 -5753 1158
rect -5709 1148 -5481 1200
rect -5437 1148 -5209 1200
rect -5165 1148 -4937 1200
rect -4893 1148 -4665 1200
rect -4621 1148 -4529 1333
rect -6389 -96 -5973 482
rect -5845 36 -5617 88
rect -5573 36 -5345 88
rect -5301 36 -5073 88
rect -5029 36 -4801 88
rect -4757 36 -4529 88
rect -4397 -96 -4239 1333
rect -3434 773 -3281 1556
rect -3228 863 -3108 2835
rect -2966 1939 -2826 2867
rect -2642 2835 -2564 2975
rect -2270 2867 -1898 2919
rect -2966 1759 -2956 1939
rect -2836 1759 -2826 1939
rect -3228 725 -3150 863
rect -2966 831 -2826 1759
rect -2684 863 -2564 2835
rect -2416 863 -2296 2835
rect -2154 1939 -2014 2867
rect -1830 2835 -1752 2975
rect -1141 2971 1480 2975
rect -1458 2867 -1086 2919
rect -2154 1759 -2144 1939
rect -2024 1759 -2014 1939
rect -3082 779 -2710 831
rect -2416 725 -2338 863
rect -2154 831 -2014 1759
rect -1872 863 -1752 2835
rect -1604 863 -1484 2835
rect -1342 1939 -1202 2867
rect -1018 2835 -940 2971
rect -1342 1759 -1332 1939
rect -1212 1759 -1202 1939
rect -2270 779 -1898 831
rect -1604 725 -1526 863
rect -1342 831 -1202 1759
rect -1060 863 -940 2835
rect -1458 779 -1086 831
rect -887 773 -799 2971
rect -705 2301 -34 2777
rect -3228 715 -3061 725
rect -3228 342 -3218 715
rect -3071 342 -3061 715
rect -3228 332 -3061 342
rect -2416 715 -2249 725
rect -2416 342 -2406 715
rect -2259 342 -2249 715
rect -2416 332 -2249 342
rect -1604 715 -1437 725
rect -1604 342 -1594 715
rect -1447 489 -1437 715
rect -705 489 -548 2301
rect 213 1487 1480 2971
rect 1580 3263 2969 3273
rect 1580 3087 2773 3263
rect 2959 3087 2969 3263
rect 1580 3077 2969 3087
rect 1580 2291 1776 3077
rect 1580 2098 1590 2291
rect 1766 2098 1776 2291
rect 1580 2088 1776 2098
rect -1447 342 -548 489
rect -1604 332 -548 342
rect -6389 -279 -4239 -96
rect -6389 -443 -1045 -279
rect -6389 -4870 -5973 -443
rect -5845 -505 -5653 -495
rect -5845 -617 -5835 -505
rect -5663 -617 -5653 -505
rect -5137 -505 -4945 -495
rect -5845 -627 -5653 -617
rect -5609 -627 -5181 -575
rect -5137 -617 -5127 -505
rect -4955 -617 -4945 -505
rect -5137 -627 -4945 -617
rect -5845 -4739 -5417 -4687
rect -5373 -4739 -4945 -4687
rect -4814 -4870 -4560 -443
rect -4426 -505 -4234 -495
rect -4426 -617 -4416 -505
rect -4244 -617 -4234 -505
rect -3718 -505 -3526 -495
rect -4426 -627 -4234 -617
rect -4190 -627 -3762 -575
rect -3718 -617 -3708 -505
rect -3536 -617 -3526 -505
rect -3718 -627 -3526 -617
rect -4426 -4739 -3998 -4687
rect -3954 -4739 -3526 -4687
rect -3392 -4870 -3134 -443
rect -2999 -505 -2807 -495
rect -2999 -617 -2989 -505
rect -2817 -617 -2807 -505
rect -2999 -627 -2807 -617
rect -2999 -2837 -2807 -2827
rect -2999 -2961 -2989 -2837
rect -2817 -2961 -2807 -2837
rect -2999 -2971 -2807 -2961
rect -6389 -4919 -3134 -4870
rect -2674 -4919 -2413 -443
rect -2279 -505 -2087 -495
rect -2279 -617 -2269 -505
rect -2097 -617 -2087 -505
rect -1571 -505 -1379 -495
rect -2279 -627 -2087 -617
rect -2043 -627 -1615 -575
rect -1571 -617 -1561 -505
rect -1389 -617 -1379 -505
rect -1571 -627 -1379 -617
rect -2279 -4739 -1851 -4687
rect -1807 -4739 -1379 -4687
rect -1246 -4919 -1045 -443
rect -942 -537 -782 -527
rect -942 -677 -932 -537
rect -792 -677 -782 -537
rect -6389 -4923 -3135 -4919
rect -6389 -5199 -3417 -4923
rect -942 -5022 -782 -677
rect -3339 -5032 -782 -5022
rect -3339 -5190 -3329 -5032
rect -3198 -5190 -782 -5032
rect -6389 -5573 -5973 -5199
rect -3339 -5200 -782 -5190
rect -682 -765 -522 -527
rect -682 -905 -672 -765
rect -532 -905 -522 -765
rect -682 -5300 -522 -905
rect -4760 -5310 -522 -5300
rect -4760 -5468 -4750 -5310
rect -4621 -5468 -522 -5310
rect -4760 -5478 -522 -5468
rect -418 -5007 -121 -3396
rect -6389 -5900 -2485 -5573
rect -418 -5854 30 -5007
rect -6389 -6475 -5706 -5900
rect -5619 -6102 -5219 -5989
rect -5619 -6274 -5503 -6102
rect -5331 -6274 -5219 -6102
rect -5619 -6389 -5219 -6274
rect -5135 -6475 -4545 -5900
rect -4459 -6102 -4059 -5989
rect -4459 -6274 -4346 -6102
rect -4174 -6274 -4059 -6102
rect -4459 -6389 -4059 -6274
rect -3971 -6475 -3381 -5900
rect -3299 -6102 -2899 -5989
rect -3299 -6274 -3183 -6102
rect -3011 -6274 -2899 -6102
rect -3299 -6389 -2899 -6274
rect -2814 -6475 -2485 -5900
rect -6389 -7065 -2485 -6475
rect -6389 -7635 -5706 -7065
rect -5619 -7264 -5219 -7149
rect -5619 -7436 -5503 -7264
rect -5331 -7436 -5219 -7264
rect -5619 -7549 -5219 -7436
rect -5135 -7635 -4545 -7065
rect -4459 -7285 -4059 -7149
rect -4459 -7414 -4322 -7285
rect -4193 -7414 -4059 -7285
rect -4459 -7549 -4059 -7414
rect -3971 -7635 -3381 -7065
rect -3299 -7261 -2899 -7149
rect -3299 -7433 -3183 -7261
rect -3011 -7433 -2899 -7261
rect -3299 -7549 -2899 -7433
rect -2814 -7635 -2485 -7065
rect -6389 -7888 -2485 -7635
rect -1382 -6320 30 -5854
rect -1382 -7888 -916 -6320
rect -6389 -8225 -916 -7888
rect -6389 -8792 -5706 -8225
rect -5619 -8424 -5219 -8309
rect -5619 -8596 -5503 -8424
rect -5331 -8596 -5219 -8424
rect -5619 -8709 -5219 -8596
rect -5135 -8792 -4545 -8225
rect -4459 -8424 -4059 -8309
rect -4459 -8596 -4345 -8424
rect -4173 -8596 -4059 -8424
rect -4459 -8709 -4059 -8596
rect -3971 -8792 -3381 -8225
rect -3299 -8424 -2899 -8309
rect -3299 -8596 -3183 -8424
rect -3011 -8596 -2899 -8424
rect -3299 -8709 -2899 -8596
rect -2814 -8792 -2224 -8225
rect -2139 -8446 -1739 -8309
rect -2139 -8571 -2006 -8446
rect -1877 -8571 -1739 -8446
rect -2139 -8709 -1739 -8571
rect -1658 -8792 -916 -8225
rect -6389 -9452 -916 -8792
<< via1 >>
rect -6065 1747 -6013 1796
rect -5709 1747 -5657 1796
rect -4963 2465 -4903 2545
rect -5353 1747 -5301 1796
rect -4759 2108 -4699 2188
rect -4607 2465 -4547 2545
rect -4403 2108 -4343 2188
rect -4251 2465 -4191 2545
rect -4047 2108 -3987 2188
rect -3895 2465 -3835 2545
rect -3691 2108 -3631 2188
rect -4857 1731 -4805 1796
rect -4501 1731 -4449 1796
rect -4145 1731 -4093 1796
rect -3789 1731 -3737 1796
rect -4229 1367 -4149 1447
rect -5835 1158 -5763 1271
rect -2956 1759 -2836 1939
rect -2144 1759 -2024 1939
rect -1332 1759 -1212 1939
rect -3218 342 -3071 715
rect -2406 342 -2259 715
rect -1594 342 -1447 715
rect 2773 3087 2959 3263
rect 1590 2098 1766 2291
rect -5835 -617 -5663 -505
rect -5127 -617 -4955 -505
rect -4416 -617 -4244 -505
rect -3708 -617 -3536 -505
rect -2989 -617 -2817 -505
rect -2989 -2961 -2817 -2837
rect -2269 -617 -2097 -505
rect -1561 -617 -1389 -505
rect -932 -677 -792 -537
rect -3329 -5190 -3198 -5032
rect -672 -905 -532 -765
rect -4750 -5468 -4621 -5310
rect -5503 -6274 -5331 -6102
rect -4346 -6274 -4174 -6102
rect -3183 -6274 -3011 -6102
rect -5503 -7436 -5331 -7264
rect -4322 -7414 -4193 -7285
rect -3183 -7433 -3011 -7261
rect -5503 -8596 -5331 -8424
rect -4345 -8596 -4173 -8424
rect -3183 -8596 -3011 -8424
rect -2006 -8571 -1877 -8446
<< metal2 >>
rect 2763 3263 7678 3273
rect 2763 3087 2773 3263
rect 2959 3087 7678 3263
rect 2763 3077 7678 3087
rect -4973 2545 -3322 2555
rect -4973 2465 -4963 2545
rect -4903 2465 -4607 2545
rect -4547 2465 -4251 2545
rect -4191 2465 -3895 2545
rect -3835 2465 -3322 2545
rect -4973 2455 -3322 2465
rect -4973 2188 -3501 2198
rect -4973 2108 -4759 2188
rect -4699 2108 -4403 2188
rect -4343 2108 -4047 2188
rect -3987 2108 -3691 2188
rect -3631 2108 -3501 2188
rect -4973 2098 -3501 2108
rect -6075 1796 -3651 1806
rect -6075 1747 -6065 1796
rect -6013 1747 -5709 1796
rect -5657 1747 -5353 1796
rect -5301 1747 -4857 1796
rect -6075 1731 -4857 1747
rect -4805 1731 -4501 1796
rect -4449 1731 -4145 1796
rect -4093 1731 -3789 1796
rect -3737 1731 -3651 1796
rect -6075 1714 -3651 1731
rect -5866 1271 -5753 1714
rect -3601 1457 -3501 2098
rect -3422 1949 -3322 2455
rect 2307 2331 2902 2743
rect 1580 2291 1776 2301
rect 1580 2098 1590 2291
rect 1766 2098 1776 2291
rect 1580 1949 1776 2098
rect 7482 2023 7678 3077
rect -3422 1939 1776 1949
rect -3422 1759 -2956 1939
rect -2836 1759 -2144 1939
rect -2024 1759 -1332 1939
rect -1212 1759 1776 1939
rect -3422 1749 1776 1759
rect -4239 1447 -3501 1457
rect -4239 1367 -4229 1447
rect -4149 1367 -3501 1447
rect -4239 1357 -3501 1367
rect -5866 1158 -5835 1271
rect -5763 1158 -5753 1271
rect -5866 1148 -5753 1158
rect -3228 715 -3061 725
rect -3228 342 -3218 715
rect -3071 342 -3061 715
rect -3228 -65 -3061 342
rect -2416 715 -2249 725
rect -2416 342 -2406 715
rect -2259 342 -2249 715
rect -2416 288 -2249 342
rect -5845 -187 -3061 -65
rect -2924 121 -2249 288
rect -1604 715 -1437 725
rect -1604 342 -1594 715
rect -1447 342 -1437 715
rect -5845 -505 -5653 -187
rect -2924 -263 -2757 121
rect -1604 -39 -1437 342
rect -4426 -385 -2757 -263
rect -2279 -206 -1437 -39
rect -5845 -617 -5835 -505
rect -5663 -617 -5653 -505
rect -5845 -627 -5653 -617
rect -5137 -505 -4611 -495
rect -5137 -617 -5127 -505
rect -4955 -617 -4611 -505
rect -5137 -627 -4611 -617
rect -4426 -505 -4234 -385
rect -4426 -617 -4416 -505
rect -4244 -617 -4234 -505
rect -4426 -627 -4234 -617
rect -3718 -505 -2807 -495
rect -3718 -617 -3708 -505
rect -3536 -617 -2989 -505
rect -2817 -617 -2807 -505
rect -3718 -627 -2807 -617
rect -2279 -505 -2087 -206
rect -2279 -617 -2269 -505
rect -2097 -617 -2087 -505
rect -2279 -627 -2087 -617
rect -1571 -505 -1045 -495
rect -1571 -617 -1561 -505
rect -1389 -617 -1045 -505
rect -1571 -627 -1045 -617
rect -4760 -5310 -4611 -627
rect -3339 -5032 -3188 -627
rect -3339 -5190 -3329 -5032
rect -3198 -5190 -3188 -5032
rect -3339 -5200 -3188 -5190
rect -2999 -2837 -2807 -2827
rect -2999 -2961 -2989 -2837
rect -2817 -2961 -2807 -2837
rect -4760 -5468 -4750 -5310
rect -4621 -5468 -4611 -5310
rect -5513 -6102 -5321 -6092
rect -5513 -6274 -5503 -6102
rect -5331 -6274 -5321 -6102
rect -5513 -7264 -5321 -6274
rect -5513 -7436 -5503 -7264
rect -5331 -7436 -5321 -7264
rect -4760 -7275 -4611 -5468
rect -2999 -6092 -2807 -2961
rect -1194 -5598 -1045 -627
rect -942 -537 -346 -527
rect -942 -677 -932 -537
rect -792 -677 -346 -537
rect -942 -687 -346 -677
rect -942 -765 -350 -755
rect -942 -905 -672 -765
rect -532 -905 -350 -765
rect -942 -915 -350 -905
rect -4356 -6102 -2807 -6092
rect -4356 -6274 -4346 -6102
rect -4174 -6274 -3183 -6102
rect -3011 -6274 -2807 -6102
rect -4356 -6284 -2807 -6274
rect -2016 -5747 -1045 -5598
rect -3193 -7261 -3001 -6284
rect -4760 -7285 -4183 -7275
rect -4760 -7414 -4322 -7285
rect -4193 -7414 -4183 -7285
rect -4760 -7424 -4183 -7414
rect -5513 -8414 -5321 -7436
rect -3193 -7433 -3183 -7261
rect -3011 -7433 -3001 -7261
rect -3193 -8414 -3001 -7433
rect -5513 -8424 -3001 -8414
rect -5513 -8596 -5503 -8424
rect -5331 -8596 -4345 -8424
rect -4173 -8596 -3183 -8424
rect -3011 -8596 -3001 -8424
rect -2016 -8446 -1867 -5747
rect -2016 -8571 -2006 -8446
rect -1877 -8571 -1867 -8446
rect -2016 -8581 -1867 -8571
rect -5513 -8606 -3001 -8596
use bmbgota  bmbgota_0
timestamp 1748514987
transform 1 0 4 0 1 0
box -422 -9462 7674 3284
use hvpmos_5L3PPQ  hvpmos_5L3PPQ_0
timestamp 1748546292
transform 1 0 -2896 0 1 1849
box -560 -1124 560 1302
use hvpmos_5L3PPQ  hvpmos_5L3PPQ_1
timestamp 1748546292
transform 1 0 -2084 0 1 1849
box -560 -1124 560 1302
use hvpmos_5L3PPQ  hvpmos_5L3PPQ_2
timestamp 1748546292
transform 1 0 -1272 0 1 1849
box -560 -1124 560 1302
use hvpmos_UB3TJ6  hvpmos_UB3TJ6_0
timestamp 1748595295
transform 1 0 -5899 0 1 2327
box -464 -824 2600 824
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_0
timestamp 1748598742
transform 1 0 -5419 0 1 -6189
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_1
timestamp 1748598742
transform 1 0 -4259 0 1 -6189
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_2
timestamp 1748598742
transform 1 0 -3099 0 1 -6189
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_3
timestamp 1748598742
transform 1 0 -5419 0 1 -7349
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_4
timestamp 1748598742
transform 1 0 -4259 0 1 -7349
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_5
timestamp 1748598742
transform 1 0 -3099 0 1 -7349
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_6
timestamp 1748598742
transform 1 0 -5419 0 1 -8509
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_7
timestamp 1748598742
transform 1 0 -4259 0 1 -8509
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_8
timestamp 1748598742
transform 1 0 -3099 0 1 -8509
box -508 -508 508 508
use pnpmpa_KGYYW3  pnpmpa_KGYYW3_9
timestamp 1748598742
transform 1 0 -1939 0 1 -8509
box -508 -508 508 508
use rhigh_2665BW  rhigh_2665BW_0
timestamp 1748543940
transform 1 0 -5799 0 1 618
box -230 -766 1454 766
use rppd_7BUPFW  rppd_7BUPFW_0
timestamp 1748556962
transform 1 0 -2903 0 1 -1727
box -280 -1336 280 1336
use rppd_R9R9UC  rppd_R9R9UC_0
timestamp 1748556962
transform 1 0 -4330 0 1 -2657
box -280 -2266 988 2266
use rppd_R9R9UC  rppd_R9R9UC_1
timestamp 1748556962
transform 1 0 -5749 0 1 -2657
box -280 -2266 988 2266
use rppd_R9R9UC  rppd_R9R9UC_2
timestamp 1748556962
transform 1 0 -2183 0 1 -2657
box -280 -2266 988 2266
<< labels >>
flabel metal1 -6389 430 -6156 1457 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal2 2307 2331 2902 2743 0 FreeSans 800 0 0 0 IB
port 3 nsew
flabel metal1 -705 2301 -34 2777 0 FreeSans 800 0 0 0 VREF
port 2 nsew
flabel metal1 -6389 3037 -5550 3287 0 FreeSans 800 0 0 0 VDD
port 4 nsew
<< end >>
