magic
tech ihp-sg13g2
timestamp 1749416725
<< error_p >>
rect -93 530 -88 535
rect 88 530 93 535
rect 225 530 230 535
rect 406 530 411 535
rect 543 530 548 535
rect 724 530 729 535
rect 861 530 866 535
rect 1042 530 1047 535
rect 1179 530 1184 535
rect 1360 530 1365 535
rect 1497 530 1502 535
rect 1678 530 1683 535
rect 1815 530 1820 535
rect 1996 530 2001 535
rect 2133 530 2138 535
rect 2314 530 2319 535
rect 2451 530 2456 535
rect 2632 530 2637 535
rect 2769 530 2774 535
rect 2950 530 2955 535
rect -98 525 -93 530
rect 93 525 98 530
rect 220 525 225 530
rect 411 525 416 530
rect 538 525 543 530
rect 729 525 734 530
rect 856 525 861 530
rect 1047 525 1052 530
rect 1174 525 1179 530
rect 1365 525 1370 530
rect 1492 525 1497 530
rect 1683 525 1688 530
rect 1810 525 1815 530
rect 2001 525 2006 530
rect 2128 525 2133 530
rect 2319 525 2324 530
rect 2446 525 2451 530
rect 2637 525 2642 530
rect 2764 525 2769 530
rect 2955 525 2960 530
rect -98 514 -93 519
rect 93 514 98 519
rect 220 514 225 519
rect 411 514 416 519
rect 538 514 543 519
rect 729 514 734 519
rect 856 514 861 519
rect 1047 514 1052 519
rect 1174 514 1179 519
rect 1365 514 1370 519
rect 1492 514 1497 519
rect 1683 514 1688 519
rect 1810 514 1815 519
rect 2001 514 2006 519
rect 2128 514 2133 519
rect 2319 514 2324 519
rect 2446 514 2451 519
rect 2637 514 2642 519
rect 2764 514 2769 519
rect 2955 514 2960 519
rect -93 509 -88 514
rect 88 509 93 514
rect 225 509 230 514
rect 406 509 411 514
rect 543 509 548 514
rect 724 509 729 514
rect 861 509 866 514
rect 1042 509 1047 514
rect 1179 509 1184 514
rect 1360 509 1365 514
rect 1497 509 1502 514
rect 1678 509 1683 514
rect 1815 509 1820 514
rect 1996 509 2001 514
rect 2133 509 2138 514
rect 2314 509 2319 514
rect 2451 509 2456 514
rect 2632 509 2637 514
rect 2769 509 2774 514
rect 2950 509 2955 514
rect -127 493 -122 498
rect -116 493 -111 498
rect 111 493 116 498
rect 122 493 127 498
rect 191 493 196 498
rect 202 493 207 498
rect 429 493 434 498
rect 440 493 445 498
rect 509 493 514 498
rect 520 493 525 498
rect 747 493 752 498
rect 758 493 763 498
rect 827 493 832 498
rect 838 493 843 498
rect 1065 493 1070 498
rect 1076 493 1081 498
rect 1145 493 1150 498
rect 1156 493 1161 498
rect 1383 493 1388 498
rect 1394 493 1399 498
rect 1463 493 1468 498
rect 1474 493 1479 498
rect 1701 493 1706 498
rect 1712 493 1717 498
rect 1781 493 1786 498
rect 1792 493 1797 498
rect 2019 493 2024 498
rect 2030 493 2035 498
rect 2099 493 2104 498
rect 2110 493 2115 498
rect 2337 493 2342 498
rect 2348 493 2353 498
rect 2417 493 2422 498
rect 2428 493 2433 498
rect 2655 493 2660 498
rect 2666 493 2671 498
rect 2735 493 2740 498
rect 2746 493 2751 498
rect 2973 493 2978 498
rect 2984 493 2989 498
rect -132 488 -127 493
rect -111 488 -106 493
rect 106 488 111 493
rect 127 488 132 493
rect 186 488 191 493
rect 207 488 212 493
rect 424 488 429 493
rect 445 488 450 493
rect 504 488 509 493
rect 525 488 530 493
rect 742 488 747 493
rect 763 488 768 493
rect 822 488 827 493
rect 843 488 848 493
rect 1060 488 1065 493
rect 1081 488 1086 493
rect 1140 488 1145 493
rect 1161 488 1166 493
rect 1378 488 1383 493
rect 1399 488 1404 493
rect 1458 488 1463 493
rect 1479 488 1484 493
rect 1696 488 1701 493
rect 1717 488 1722 493
rect 1776 488 1781 493
rect 1797 488 1802 493
rect 2014 488 2019 493
rect 2035 488 2040 493
rect 2094 488 2099 493
rect 2115 488 2120 493
rect 2332 488 2337 493
rect 2353 488 2358 493
rect 2412 488 2417 493
rect 2433 488 2438 493
rect 2650 488 2655 493
rect 2671 488 2676 493
rect 2730 488 2735 493
rect 2751 488 2756 493
rect 2968 488 2973 493
rect 2989 488 2994 493
rect -132 -493 -127 -488
rect -111 -493 -106 -488
rect 106 -493 111 -488
rect 127 -493 132 -488
rect 186 -493 191 -488
rect 207 -493 212 -488
rect 424 -493 429 -488
rect 445 -493 450 -488
rect 504 -493 509 -488
rect 525 -493 530 -488
rect 742 -493 747 -488
rect 763 -493 768 -488
rect 822 -493 827 -488
rect 843 -493 848 -488
rect 1060 -493 1065 -488
rect 1081 -493 1086 -488
rect 1140 -493 1145 -488
rect 1161 -493 1166 -488
rect 1378 -493 1383 -488
rect 1399 -493 1404 -488
rect 1458 -493 1463 -488
rect 1479 -493 1484 -488
rect 1696 -493 1701 -488
rect 1717 -493 1722 -488
rect 1776 -493 1781 -488
rect 1797 -493 1802 -488
rect 2014 -493 2019 -488
rect 2035 -493 2040 -488
rect 2094 -493 2099 -488
rect 2115 -493 2120 -488
rect 2332 -493 2337 -488
rect 2353 -493 2358 -488
rect 2412 -493 2417 -488
rect 2433 -493 2438 -488
rect 2650 -493 2655 -488
rect 2671 -493 2676 -488
rect 2730 -493 2735 -488
rect 2751 -493 2756 -488
rect 2968 -493 2973 -488
rect 2989 -493 2994 -488
rect -127 -498 -122 -493
rect -116 -498 -111 -493
rect 111 -498 116 -493
rect 122 -498 127 -493
rect 191 -498 196 -493
rect 202 -498 207 -493
rect 429 -498 434 -493
rect 440 -498 445 -493
rect 509 -498 514 -493
rect 520 -498 525 -493
rect 747 -498 752 -493
rect 758 -498 763 -493
rect 827 -498 832 -493
rect 838 -498 843 -493
rect 1065 -498 1070 -493
rect 1076 -498 1081 -493
rect 1145 -498 1150 -493
rect 1156 -498 1161 -493
rect 1383 -498 1388 -493
rect 1394 -498 1399 -493
rect 1463 -498 1468 -493
rect 1474 -498 1479 -493
rect 1701 -498 1706 -493
rect 1712 -498 1717 -493
rect 1781 -498 1786 -493
rect 1792 -498 1797 -493
rect 2019 -498 2024 -493
rect 2030 -498 2035 -493
rect 2099 -498 2104 -493
rect 2110 -498 2115 -493
rect 2337 -498 2342 -493
rect 2348 -498 2353 -493
rect 2417 -498 2422 -493
rect 2428 -498 2433 -493
rect 2655 -498 2660 -493
rect 2666 -498 2671 -493
rect 2735 -498 2740 -493
rect 2746 -498 2751 -493
rect 2973 -498 2978 -493
rect 2984 -498 2989 -493
rect -93 -514 -88 -509
rect 88 -514 93 -509
rect 225 -514 230 -509
rect 406 -514 411 -509
rect 543 -514 548 -509
rect 724 -514 729 -509
rect 861 -514 866 -509
rect 1042 -514 1047 -509
rect 1179 -514 1184 -509
rect 1360 -514 1365 -509
rect 1497 -514 1502 -509
rect 1678 -514 1683 -509
rect 1815 -514 1820 -509
rect 1996 -514 2001 -509
rect 2133 -514 2138 -509
rect 2314 -514 2319 -509
rect 2451 -514 2456 -509
rect 2632 -514 2637 -509
rect 2769 -514 2774 -509
rect 2950 -514 2955 -509
rect -98 -519 -93 -514
rect 93 -519 98 -514
rect 220 -519 225 -514
rect 411 -519 416 -514
rect 538 -519 543 -514
rect 729 -519 734 -514
rect 856 -519 861 -514
rect 1047 -519 1052 -514
rect 1174 -519 1179 -514
rect 1365 -519 1370 -514
rect 1492 -519 1497 -514
rect 1683 -519 1688 -514
rect 1810 -519 1815 -514
rect 2001 -519 2006 -514
rect 2128 -519 2133 -514
rect 2319 -519 2324 -514
rect 2446 -519 2451 -514
rect 2637 -519 2642 -514
rect 2764 -519 2769 -514
rect 2955 -519 2960 -514
rect -98 -530 -93 -525
rect 93 -530 98 -525
rect 220 -530 225 -525
rect 411 -530 416 -525
rect 538 -530 543 -525
rect 729 -530 734 -525
rect 856 -530 861 -525
rect 1047 -530 1052 -525
rect 1174 -530 1179 -525
rect 1365 -530 1370 -525
rect 1492 -530 1497 -525
rect 1683 -530 1688 -525
rect 1810 -530 1815 -525
rect 2001 -530 2006 -525
rect 2128 -530 2133 -525
rect 2319 -530 2324 -525
rect 2446 -530 2451 -525
rect 2637 -530 2642 -525
rect 2764 -530 2769 -525
rect 2955 -530 2960 -525
rect -93 -535 -88 -530
rect 88 -535 93 -530
rect 225 -535 230 -530
rect 406 -535 411 -530
rect 543 -535 548 -530
rect 724 -535 729 -530
rect 861 -535 866 -530
rect 1042 -535 1047 -530
rect 1179 -535 1184 -530
rect 1360 -535 1365 -530
rect 1497 -535 1502 -530
rect 1678 -535 1683 -530
rect 1815 -535 1820 -530
rect 1996 -535 2001 -530
rect 2133 -535 2138 -530
rect 2314 -535 2319 -530
rect 2451 -535 2456 -530
rect 2632 -535 2637 -530
rect 2769 -535 2774 -530
rect 2950 -535 2955 -530
<< hvnmos >>
rect -100 -500 100 500
rect 218 -500 418 500
rect 536 -500 736 500
rect 854 -500 1054 500
rect 1172 -500 1372 500
rect 1490 -500 1690 500
rect 1808 -500 2008 500
rect 2126 -500 2326 500
rect 2444 -500 2644 500
rect 2762 -500 2962 500
<< hvndiff >>
rect -134 493 -100 500
rect -134 -493 -127 493
rect -111 -493 -100 493
rect -134 -500 -100 -493
rect 100 493 134 500
rect 100 -493 111 493
rect 127 -493 134 493
rect 100 -500 134 -493
rect 184 493 218 500
rect 184 -493 191 493
rect 207 -493 218 493
rect 184 -500 218 -493
rect 418 493 452 500
rect 418 -493 429 493
rect 445 -493 452 493
rect 418 -500 452 -493
rect 502 493 536 500
rect 502 -493 509 493
rect 525 -493 536 493
rect 502 -500 536 -493
rect 736 493 770 500
rect 736 -493 747 493
rect 763 -493 770 493
rect 736 -500 770 -493
rect 820 493 854 500
rect 820 -493 827 493
rect 843 -493 854 493
rect 820 -500 854 -493
rect 1054 493 1088 500
rect 1054 -493 1065 493
rect 1081 -493 1088 493
rect 1054 -500 1088 -493
rect 1138 493 1172 500
rect 1138 -493 1145 493
rect 1161 -493 1172 493
rect 1138 -500 1172 -493
rect 1372 493 1406 500
rect 1372 -493 1383 493
rect 1399 -493 1406 493
rect 1372 -500 1406 -493
rect 1456 493 1490 500
rect 1456 -493 1463 493
rect 1479 -493 1490 493
rect 1456 -500 1490 -493
rect 1690 493 1724 500
rect 1690 -493 1701 493
rect 1717 -493 1724 493
rect 1690 -500 1724 -493
rect 1774 493 1808 500
rect 1774 -493 1781 493
rect 1797 -493 1808 493
rect 1774 -500 1808 -493
rect 2008 493 2042 500
rect 2008 -493 2019 493
rect 2035 -493 2042 493
rect 2008 -500 2042 -493
rect 2092 493 2126 500
rect 2092 -493 2099 493
rect 2115 -493 2126 493
rect 2092 -500 2126 -493
rect 2326 493 2360 500
rect 2326 -493 2337 493
rect 2353 -493 2360 493
rect 2326 -500 2360 -493
rect 2410 493 2444 500
rect 2410 -493 2417 493
rect 2433 -493 2444 493
rect 2410 -500 2444 -493
rect 2644 493 2678 500
rect 2644 -493 2655 493
rect 2671 -493 2678 493
rect 2644 -500 2678 -493
rect 2728 493 2762 500
rect 2728 -493 2735 493
rect 2751 -493 2762 493
rect 2728 -500 2762 -493
rect 2962 493 2996 500
rect 2962 -493 2973 493
rect 2989 -493 2996 493
rect 2962 -500 2996 -493
<< hvndiffc >>
rect -127 -493 -111 493
rect 111 -493 127 493
rect 191 -493 207 493
rect 429 -493 445 493
rect 509 -493 525 493
rect 747 -493 763 493
rect 827 -493 843 493
rect 1065 -493 1081 493
rect 1145 -493 1161 493
rect 1383 -493 1399 493
rect 1463 -493 1479 493
rect 1701 -493 1717 493
rect 1781 -493 1797 493
rect 2019 -493 2035 493
rect 2099 -493 2115 493
rect 2337 -493 2353 493
rect 2417 -493 2433 493
rect 2655 -493 2671 493
rect 2735 -493 2751 493
rect 2973 -493 2989 493
<< psubdiff >>
rect -218 582 3080 589
rect -218 566 -181 582
rect 3043 566 3080 582
rect -218 559 3080 566
rect -218 552 -188 559
rect -218 -552 -211 552
rect -195 -552 -188 552
rect 3050 552 3080 559
rect -218 -559 -188 -552
rect 3050 -552 3057 552
rect 3073 -552 3080 552
rect 3050 -559 3080 -552
rect -218 -566 3080 -559
rect -218 -582 -181 -566
rect 3043 -582 3080 -566
rect -218 -589 3080 -582
<< psubdiffcont >>
rect -181 566 3043 582
rect -211 -552 -195 552
rect 3057 -552 3073 552
rect -181 -582 3043 -566
<< poly >>
rect -100 530 100 537
rect -100 514 -93 530
rect 93 514 100 530
rect -100 500 100 514
rect 218 530 418 537
rect 218 514 225 530
rect 411 514 418 530
rect 218 500 418 514
rect 536 530 736 537
rect 536 514 543 530
rect 729 514 736 530
rect 536 500 736 514
rect 854 530 1054 537
rect 854 514 861 530
rect 1047 514 1054 530
rect 854 500 1054 514
rect 1172 530 1372 537
rect 1172 514 1179 530
rect 1365 514 1372 530
rect 1172 500 1372 514
rect 1490 530 1690 537
rect 1490 514 1497 530
rect 1683 514 1690 530
rect 1490 500 1690 514
rect 1808 530 2008 537
rect 1808 514 1815 530
rect 2001 514 2008 530
rect 1808 500 2008 514
rect 2126 530 2326 537
rect 2126 514 2133 530
rect 2319 514 2326 530
rect 2126 500 2326 514
rect 2444 530 2644 537
rect 2444 514 2451 530
rect 2637 514 2644 530
rect 2444 500 2644 514
rect 2762 530 2962 537
rect 2762 514 2769 530
rect 2955 514 2962 530
rect 2762 500 2962 514
rect -100 -514 100 -500
rect -100 -530 -93 -514
rect 93 -530 100 -514
rect -100 -537 100 -530
rect 218 -514 418 -500
rect 218 -530 225 -514
rect 411 -530 418 -514
rect 218 -537 418 -530
rect 536 -514 736 -500
rect 536 -530 543 -514
rect 729 -530 736 -514
rect 536 -537 736 -530
rect 854 -514 1054 -500
rect 854 -530 861 -514
rect 1047 -530 1054 -514
rect 854 -537 1054 -530
rect 1172 -514 1372 -500
rect 1172 -530 1179 -514
rect 1365 -530 1372 -514
rect 1172 -537 1372 -530
rect 1490 -514 1690 -500
rect 1490 -530 1497 -514
rect 1683 -530 1690 -514
rect 1490 -537 1690 -530
rect 1808 -514 2008 -500
rect 1808 -530 1815 -514
rect 2001 -530 2008 -514
rect 1808 -537 2008 -530
rect 2126 -514 2326 -500
rect 2126 -530 2133 -514
rect 2319 -530 2326 -514
rect 2126 -537 2326 -530
rect 2444 -514 2644 -500
rect 2444 -530 2451 -514
rect 2637 -530 2644 -514
rect 2444 -537 2644 -530
rect 2762 -514 2962 -500
rect 2762 -530 2769 -514
rect 2955 -530 2962 -514
rect 2762 -537 2962 -530
<< polycont >>
rect -93 514 93 530
rect 225 514 411 530
rect 543 514 729 530
rect 861 514 1047 530
rect 1179 514 1365 530
rect 1497 514 1683 530
rect 1815 514 2001 530
rect 2133 514 2319 530
rect 2451 514 2637 530
rect 2769 514 2955 530
rect -93 -530 93 -514
rect 225 -530 411 -514
rect 543 -530 729 -514
rect 861 -530 1047 -514
rect 1179 -530 1365 -514
rect 1497 -530 1683 -514
rect 1815 -530 2001 -514
rect 2133 -530 2319 -514
rect 2451 -530 2637 -514
rect 2769 -530 2955 -514
<< metal1 >>
rect -216 582 3078 587
rect -216 566 -181 582
rect 3043 566 3078 582
rect -216 561 3078 566
rect -216 552 -190 561
rect -216 -552 -211 552
rect -195 -552 -190 552
rect 3052 552 3078 561
rect -216 -561 -190 -552
rect 3052 -552 3057 552
rect 3073 -552 3078 552
rect 3052 -561 3078 -552
rect -216 -566 3078 -561
rect -216 -582 -181 -566
rect 3043 -582 3078 -566
rect -216 -587 3078 -582
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 10 l 2 nf 1 nx 10 dx 0.5 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
