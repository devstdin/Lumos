magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757367233
<< poly >>
rect -224 342 56 362
rect -224 6 -204 342
rect -25 188 56 342
rect 256 342 536 362
rect 256 188 337 342
rect -25 160 337 188
rect -25 6 56 160
rect -224 -14 56 6
rect 256 6 337 160
rect 516 6 536 342
rect 256 -14 536 6
<< polycont >>
rect -204 6 -25 342
rect 337 6 516 342
<< metal1 >>
rect -586 1421 -5 1441
rect -586 -1055 -566 1421
rect -25 -1055 -5 1421
rect 317 612 657 622
rect 317 -248 327 612
rect 647 -248 657 612
rect 317 -258 657 -248
rect -586 -1075 -5 -1055
<< via1 >>
rect -566 342 -25 1421
rect -566 6 -204 342
rect -204 6 -25 342
rect -566 -1055 -25 6
rect 327 342 647 612
rect 327 6 337 342
rect 337 6 516 342
rect 516 6 647 342
rect 327 -248 647 6
<< metal2 >>
rect -586 1421 -5 1441
rect -586 -1055 -566 1421
rect -25 -1055 -5 1421
rect 317 612 657 622
rect 317 -248 327 612
rect 647 -248 657 612
rect 317 -258 657 -248
rect -586 -1075 -5 -1055
<< via2 >>
rect -566 -1055 -25 1421
rect 337 -238 637 602
<< metal3 >>
rect -586 1421 -5 1441
rect -586 -1055 -566 1421
rect -25 -1055 -5 1421
rect 317 602 657 622
rect 317 -238 337 602
rect 637 -238 657 602
rect 317 -258 657 -238
rect -586 -1075 -5 -1055
<< fillblock >>
rect -284 -194 596 542
<< labels >>
flabel metal3 -586 -1075 -427 1441 0 FreeSans 800 0 0 0 T1
port 1 nsew
flabel metal3 527 -258 657 622 0 FreeSans 800 0 0 0 T2
port 3 nsew
<< properties >>
string device primitive
<< end >>
