magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757447377
<< psubdiff >>
rect 750 1232 810 1246
rect 750 -866 764 1232
rect 796 -866 810 1232
rect 12184 1097 12244 1111
rect 12184 -731 12198 1097
rect 12230 -731 12244 1097
rect 12184 -745 12244 -731
rect 750 -880 810 -866
<< psubdiffcont >>
rect 764 -866 796 1232
rect 12198 -731 12230 1097
<< metal1 >>
rect -586 -1075 -546 1441
rect 754 1349 962 1401
rect 754 1232 806 1349
rect 754 -866 764 1232
rect 796 -866 806 1232
rect 1035 1211 12571 1302
rect 1035 1201 1107 1211
rect 1313 1201 1385 1211
rect 1591 1201 1663 1211
rect 1869 1201 1941 1211
rect 2147 1201 2219 1211
rect 2425 1201 2497 1211
rect 2703 1201 2775 1211
rect 2981 1201 3053 1211
rect 3259 1201 3331 1211
rect 3537 1201 3609 1211
rect 3815 1201 3887 1211
rect 4093 1201 4165 1211
rect 4371 1201 4443 1211
rect 4649 1201 4721 1211
rect 4927 1201 4999 1211
rect 5205 1201 5277 1211
rect 5483 1201 5555 1211
rect 5761 1201 5833 1211
rect 6039 1201 6111 1211
rect 6317 1201 6389 1211
rect 6595 1201 6667 1211
rect 6873 1201 6945 1211
rect 7151 1201 7223 1211
rect 7429 1201 7501 1211
rect 7707 1201 7779 1211
rect 7985 1201 8057 1211
rect 8263 1201 8335 1211
rect 8541 1201 8613 1211
rect 8819 1201 8891 1211
rect 9097 1201 9169 1211
rect 9375 1201 9447 1211
rect 9653 1201 9725 1211
rect 9931 1201 10003 1211
rect 10209 1201 10281 1211
rect 10487 1201 10559 1211
rect 10765 1201 10837 1211
rect 11043 1201 11115 1211
rect 11321 1201 11393 1211
rect 11599 1201 11671 1211
rect 11877 1201 11949 1211
rect 953 612 1009 1169
rect 953 -248 959 612
rect 1003 -248 1009 612
rect 953 -803 1009 -248
rect 1055 -835 1087 1201
rect 1133 1159 1189 1169
rect 1133 732 1139 1159
rect 1183 732 1189 1159
rect 1133 -368 1189 732
rect 1133 -793 1139 -368
rect 1183 -793 1189 -368
rect 1133 -803 1189 -793
rect 1231 612 1287 1169
rect 1231 -248 1237 612
rect 1281 -248 1287 612
rect 1231 -803 1287 -248
rect 1333 -835 1365 1201
rect 1411 1159 1467 1169
rect 1411 732 1417 1159
rect 1461 732 1467 1159
rect 1411 -368 1467 732
rect 1411 -793 1417 -368
rect 1461 -793 1467 -368
rect 1411 -803 1467 -793
rect 1509 612 1565 1169
rect 1509 -248 1515 612
rect 1559 -248 1565 612
rect 1509 -803 1565 -248
rect 1611 -835 1643 1201
rect 1689 1159 1745 1169
rect 1689 732 1695 1159
rect 1739 732 1745 1159
rect 1689 -368 1745 732
rect 1689 -793 1695 -368
rect 1739 -793 1745 -368
rect 1689 -803 1745 -793
rect 1787 612 1843 1169
rect 1787 -248 1793 612
rect 1837 -248 1843 612
rect 1787 -803 1843 -248
rect 1889 -835 1921 1201
rect 1967 1159 2023 1169
rect 1967 732 1973 1159
rect 2017 732 2023 1159
rect 1967 -368 2023 732
rect 1967 -793 1973 -368
rect 2017 -793 2023 -368
rect 1967 -803 2023 -793
rect 2065 612 2121 1169
rect 2065 -248 2071 612
rect 2115 -248 2121 612
rect 2065 -803 2121 -248
rect 2167 -835 2199 1201
rect 2245 1159 2301 1169
rect 2245 732 2251 1159
rect 2295 732 2301 1159
rect 2245 -368 2301 732
rect 2245 -793 2251 -368
rect 2295 -793 2301 -368
rect 2245 -803 2301 -793
rect 2343 612 2399 1169
rect 2343 -248 2349 612
rect 2393 -248 2399 612
rect 2343 -803 2399 -248
rect 2445 -835 2477 1201
rect 2523 1159 2579 1169
rect 2523 732 2529 1159
rect 2573 732 2579 1159
rect 2523 -368 2579 732
rect 2523 -793 2529 -368
rect 2573 -793 2579 -368
rect 2523 -803 2579 -793
rect 2621 612 2677 1169
rect 2621 -248 2627 612
rect 2671 -248 2677 612
rect 2621 -803 2677 -248
rect 2723 -835 2755 1201
rect 2801 1159 2857 1169
rect 2801 732 2807 1159
rect 2851 732 2857 1159
rect 2801 -368 2857 732
rect 2801 -793 2807 -368
rect 2851 -793 2857 -368
rect 2801 -803 2857 -793
rect 2899 612 2955 1169
rect 2899 -248 2905 612
rect 2949 -248 2955 612
rect 2899 -803 2955 -248
rect 3001 -835 3033 1201
rect 3079 1159 3135 1169
rect 3079 732 3085 1159
rect 3129 732 3135 1159
rect 3079 -368 3135 732
rect 3079 -793 3085 -368
rect 3129 -793 3135 -368
rect 3079 -803 3135 -793
rect 3177 612 3233 1169
rect 3177 -248 3183 612
rect 3227 -248 3233 612
rect 3177 -803 3233 -248
rect 3279 -835 3311 1201
rect 3357 1159 3413 1169
rect 3357 732 3363 1159
rect 3407 732 3413 1159
rect 3357 -368 3413 732
rect 3357 -793 3363 -368
rect 3407 -793 3413 -368
rect 3357 -803 3413 -793
rect 3455 612 3511 1169
rect 3455 -248 3461 612
rect 3505 -248 3511 612
rect 3455 -803 3511 -248
rect 3557 -835 3589 1201
rect 3635 1159 3691 1169
rect 3635 732 3641 1159
rect 3685 732 3691 1159
rect 3635 -368 3691 732
rect 3635 -793 3641 -368
rect 3685 -793 3691 -368
rect 3635 -803 3691 -793
rect 3733 612 3789 1169
rect 3733 -248 3739 612
rect 3783 -248 3789 612
rect 3733 -803 3789 -248
rect 3835 -835 3867 1201
rect 3913 1159 3969 1169
rect 3913 732 3919 1159
rect 3963 732 3969 1159
rect 3913 -368 3969 732
rect 3913 -793 3919 -368
rect 3963 -793 3969 -368
rect 3913 -803 3969 -793
rect 4011 612 4067 1169
rect 4011 -248 4017 612
rect 4061 -248 4067 612
rect 4011 -803 4067 -248
rect 4113 -835 4145 1201
rect 4191 1159 4247 1169
rect 4191 732 4197 1159
rect 4241 732 4247 1159
rect 4191 -368 4247 732
rect 4191 -793 4197 -368
rect 4241 -793 4247 -368
rect 4191 -803 4247 -793
rect 4289 612 4345 1169
rect 4289 -248 4295 612
rect 4339 -248 4345 612
rect 4289 -803 4345 -248
rect 4391 -835 4423 1201
rect 4469 1159 4525 1169
rect 4469 732 4475 1159
rect 4519 732 4525 1159
rect 4469 -368 4525 732
rect 4469 -793 4475 -368
rect 4519 -793 4525 -368
rect 4469 -803 4525 -793
rect 4567 612 4623 1169
rect 4567 -248 4573 612
rect 4617 -248 4623 612
rect 4567 -803 4623 -248
rect 4669 -835 4701 1201
rect 4747 1159 4803 1169
rect 4747 732 4753 1159
rect 4797 732 4803 1159
rect 4747 -368 4803 732
rect 4747 -793 4753 -368
rect 4797 -793 4803 -368
rect 4747 -803 4803 -793
rect 4845 612 4901 1169
rect 4845 -248 4851 612
rect 4895 -248 4901 612
rect 4845 -803 4901 -248
rect 4947 -835 4979 1201
rect 5025 1159 5081 1169
rect 5025 732 5031 1159
rect 5075 732 5081 1159
rect 5025 -368 5081 732
rect 5025 -793 5031 -368
rect 5075 -793 5081 -368
rect 5025 -803 5081 -793
rect 5123 612 5179 1169
rect 5123 -248 5129 612
rect 5173 -248 5179 612
rect 5123 -803 5179 -248
rect 5225 -835 5257 1201
rect 5303 1159 5359 1169
rect 5303 732 5309 1159
rect 5353 732 5359 1159
rect 5303 -368 5359 732
rect 5303 -793 5309 -368
rect 5353 -793 5359 -368
rect 5303 -803 5359 -793
rect 5401 612 5457 1169
rect 5401 -248 5407 612
rect 5451 -248 5457 612
rect 5401 -803 5457 -248
rect 5503 -835 5535 1201
rect 5581 1159 5637 1169
rect 5581 732 5587 1159
rect 5631 732 5637 1159
rect 5581 -368 5637 732
rect 5581 -793 5587 -368
rect 5631 -793 5637 -368
rect 5581 -803 5637 -793
rect 5679 612 5735 1169
rect 5679 -248 5685 612
rect 5729 -248 5735 612
rect 5679 -803 5735 -248
rect 5781 -835 5813 1201
rect 5859 1159 5915 1169
rect 5859 732 5865 1159
rect 5909 732 5915 1159
rect 5859 -368 5915 732
rect 5859 -793 5865 -368
rect 5909 -793 5915 -368
rect 5859 -803 5915 -793
rect 5957 612 6013 1169
rect 5957 -248 5963 612
rect 6007 -248 6013 612
rect 5957 -803 6013 -248
rect 6059 -835 6091 1201
rect 6137 1159 6193 1169
rect 6137 732 6143 1159
rect 6187 732 6193 1159
rect 6137 -368 6193 732
rect 6137 -793 6143 -368
rect 6187 -793 6193 -368
rect 6137 -803 6193 -793
rect 6235 612 6291 1169
rect 6235 -248 6241 612
rect 6285 -248 6291 612
rect 6235 -803 6291 -248
rect 6337 -835 6369 1201
rect 6415 1159 6471 1169
rect 6415 732 6421 1159
rect 6465 732 6471 1159
rect 6415 -368 6471 732
rect 6415 -793 6421 -368
rect 6465 -793 6471 -368
rect 6415 -803 6471 -793
rect 6513 612 6569 1169
rect 6513 -248 6519 612
rect 6563 -248 6569 612
rect 6513 -803 6569 -248
rect 6615 -835 6647 1201
rect 6693 1159 6749 1169
rect 6693 732 6699 1159
rect 6743 732 6749 1159
rect 6693 -368 6749 732
rect 6693 -793 6699 -368
rect 6743 -793 6749 -368
rect 6693 -803 6749 -793
rect 6791 612 6847 1169
rect 6791 -248 6797 612
rect 6841 -248 6847 612
rect 6791 -803 6847 -248
rect 6893 -835 6925 1201
rect 6971 1159 7027 1169
rect 6971 732 6977 1159
rect 7021 732 7027 1159
rect 6971 -368 7027 732
rect 6971 -793 6977 -368
rect 7021 -793 7027 -368
rect 6971 -803 7027 -793
rect 7069 612 7125 1169
rect 7069 -248 7075 612
rect 7119 -248 7125 612
rect 7069 -803 7125 -248
rect 7171 -835 7203 1201
rect 7249 1159 7305 1169
rect 7249 732 7255 1159
rect 7299 732 7305 1159
rect 7249 -368 7305 732
rect 7249 -793 7255 -368
rect 7299 -793 7305 -368
rect 7249 -803 7305 -793
rect 7347 612 7403 1169
rect 7347 -248 7353 612
rect 7397 -248 7403 612
rect 7347 -803 7403 -248
rect 7449 -835 7481 1201
rect 7527 1159 7583 1169
rect 7527 732 7533 1159
rect 7577 732 7583 1159
rect 7527 -368 7583 732
rect 7527 -793 7533 -368
rect 7577 -793 7583 -368
rect 7527 -803 7583 -793
rect 7625 612 7681 1169
rect 7625 -248 7631 612
rect 7675 -248 7681 612
rect 7625 -803 7681 -248
rect 7727 -835 7759 1201
rect 7805 1159 7861 1169
rect 7805 732 7811 1159
rect 7855 732 7861 1159
rect 7805 -368 7861 732
rect 7805 -793 7811 -368
rect 7855 -793 7861 -368
rect 7805 -803 7861 -793
rect 7903 612 7959 1169
rect 7903 -248 7909 612
rect 7953 -248 7959 612
rect 7903 -803 7959 -248
rect 8005 -835 8037 1201
rect 8083 1159 8139 1169
rect 8083 732 8089 1159
rect 8133 732 8139 1159
rect 8083 -368 8139 732
rect 8083 -793 8089 -368
rect 8133 -793 8139 -368
rect 8083 -803 8139 -793
rect 8181 612 8237 1169
rect 8181 -248 8187 612
rect 8231 -248 8237 612
rect 8181 -803 8237 -248
rect 8283 -835 8315 1201
rect 8361 1159 8417 1169
rect 8361 732 8367 1159
rect 8411 732 8417 1159
rect 8361 -368 8417 732
rect 8361 -793 8367 -368
rect 8411 -793 8417 -368
rect 8361 -803 8417 -793
rect 8459 612 8515 1169
rect 8459 -248 8465 612
rect 8509 -248 8515 612
rect 8459 -803 8515 -248
rect 8561 -835 8593 1201
rect 8639 1159 8695 1169
rect 8639 732 8645 1159
rect 8689 732 8695 1159
rect 8639 -368 8695 732
rect 8639 -793 8645 -368
rect 8689 -793 8695 -368
rect 8639 -803 8695 -793
rect 8737 612 8793 1169
rect 8737 -248 8743 612
rect 8787 -248 8793 612
rect 8737 -803 8793 -248
rect 8839 -835 8871 1201
rect 8917 1159 8973 1169
rect 8917 732 8923 1159
rect 8967 732 8973 1159
rect 8917 -368 8973 732
rect 8917 -793 8923 -368
rect 8967 -793 8973 -368
rect 8917 -803 8973 -793
rect 9015 612 9071 1169
rect 9015 -248 9021 612
rect 9065 -248 9071 612
rect 9015 -803 9071 -248
rect 9117 -835 9149 1201
rect 9195 1159 9251 1169
rect 9195 732 9201 1159
rect 9245 732 9251 1159
rect 9195 -368 9251 732
rect 9195 -793 9201 -368
rect 9245 -793 9251 -368
rect 9195 -803 9251 -793
rect 9293 612 9349 1169
rect 9293 -248 9299 612
rect 9343 -248 9349 612
rect 9293 -803 9349 -248
rect 9395 -835 9427 1201
rect 9473 1159 9529 1169
rect 9473 732 9479 1159
rect 9523 732 9529 1159
rect 9473 -368 9529 732
rect 9473 -793 9479 -368
rect 9523 -793 9529 -368
rect 9473 -803 9529 -793
rect 9571 612 9627 1169
rect 9571 -248 9577 612
rect 9621 -248 9627 612
rect 9571 -803 9627 -248
rect 9673 -835 9705 1201
rect 9751 1159 9807 1169
rect 9751 732 9757 1159
rect 9801 732 9807 1159
rect 9751 -368 9807 732
rect 9751 -793 9757 -368
rect 9801 -793 9807 -368
rect 9751 -803 9807 -793
rect 9849 612 9905 1169
rect 9849 -248 9855 612
rect 9899 -248 9905 612
rect 9849 -803 9905 -248
rect 9951 -835 9983 1201
rect 10029 1159 10085 1169
rect 10029 732 10035 1159
rect 10079 732 10085 1159
rect 10029 -368 10085 732
rect 10029 -793 10035 -368
rect 10079 -793 10085 -368
rect 10029 -803 10085 -793
rect 10127 612 10183 1169
rect 10127 -248 10133 612
rect 10177 -248 10183 612
rect 10127 -803 10183 -248
rect 10229 -835 10261 1201
rect 10307 1159 10363 1169
rect 10307 732 10313 1159
rect 10357 732 10363 1159
rect 10307 -368 10363 732
rect 10307 -793 10313 -368
rect 10357 -793 10363 -368
rect 10307 -803 10363 -793
rect 10405 612 10461 1169
rect 10405 -248 10411 612
rect 10455 -248 10461 612
rect 10405 -803 10461 -248
rect 10507 -835 10539 1201
rect 10585 1159 10641 1169
rect 10585 732 10591 1159
rect 10635 732 10641 1159
rect 10585 -368 10641 732
rect 10585 -793 10591 -368
rect 10635 -793 10641 -368
rect 10585 -803 10641 -793
rect 10683 612 10739 1169
rect 10683 -248 10689 612
rect 10733 -248 10739 612
rect 10683 -803 10739 -248
rect 10785 -835 10817 1201
rect 10863 1159 10919 1169
rect 10863 732 10869 1159
rect 10913 732 10919 1159
rect 10863 -368 10919 732
rect 10863 -793 10869 -368
rect 10913 -793 10919 -368
rect 10863 -803 10919 -793
rect 10961 612 11017 1169
rect 10961 -248 10967 612
rect 11011 -248 11017 612
rect 10961 -803 11017 -248
rect 11063 -835 11095 1201
rect 11141 1159 11197 1169
rect 11141 732 11147 1159
rect 11191 732 11197 1159
rect 11141 -368 11197 732
rect 11141 -793 11147 -368
rect 11191 -793 11197 -368
rect 11141 -803 11197 -793
rect 11239 612 11295 1169
rect 11239 -248 11245 612
rect 11289 -248 11295 612
rect 11239 -803 11295 -248
rect 11341 -835 11373 1201
rect 11419 1159 11475 1169
rect 11419 732 11425 1159
rect 11469 732 11475 1159
rect 11419 -368 11475 732
rect 11419 -793 11425 -368
rect 11469 -793 11475 -368
rect 11419 -803 11475 -793
rect 11517 612 11573 1169
rect 11517 -248 11523 612
rect 11567 -248 11573 612
rect 11517 -803 11573 -248
rect 11619 -835 11651 1201
rect 11697 1159 11753 1169
rect 11697 732 11703 1159
rect 11747 732 11753 1159
rect 11697 -368 11753 732
rect 11697 -793 11703 -368
rect 11747 -793 11753 -368
rect 11697 -803 11753 -793
rect 11795 612 11851 1169
rect 11795 -248 11801 612
rect 11845 -248 11851 612
rect 11795 -803 11851 -248
rect 11897 -835 11929 1201
rect 11975 1159 12031 1169
rect 11975 732 11981 1159
rect 12025 732 12031 1159
rect 11975 -368 12031 732
rect 11975 -793 11981 -368
rect 12025 -793 12031 -368
rect 12188 1097 12240 1107
rect 12188 -731 12190 1097
rect 12238 -731 12240 1097
rect 12188 -741 12240 -731
rect 11975 -803 12031 -793
rect 754 -983 806 -866
rect 1035 -845 1107 -835
rect 1313 -845 1385 -835
rect 1591 -845 1663 -835
rect 1869 -845 1941 -835
rect 2147 -845 2219 -835
rect 2425 -845 2497 -835
rect 2703 -845 2775 -835
rect 2981 -845 3053 -835
rect 3259 -845 3331 -835
rect 3537 -845 3609 -835
rect 3815 -845 3887 -835
rect 4093 -845 4165 -835
rect 4371 -845 4443 -835
rect 4649 -845 4721 -835
rect 4927 -845 4999 -835
rect 5205 -845 5277 -835
rect 5483 -845 5555 -835
rect 5761 -845 5833 -835
rect 6039 -845 6111 -835
rect 6317 -845 6389 -835
rect 6595 -845 6667 -835
rect 6873 -845 6945 -835
rect 7151 -845 7223 -835
rect 7429 -845 7501 -835
rect 7707 -845 7779 -835
rect 7985 -845 8057 -835
rect 8263 -845 8335 -835
rect 8541 -845 8613 -835
rect 8819 -845 8891 -835
rect 9097 -845 9169 -835
rect 9375 -845 9447 -835
rect 9653 -845 9725 -835
rect 9931 -845 10003 -835
rect 10209 -845 10281 -835
rect 10487 -845 10559 -835
rect 10765 -845 10837 -835
rect 11043 -845 11115 -835
rect 11321 -845 11393 -835
rect 11599 -845 11671 -835
rect 11877 -845 11949 -835
rect 12499 -845 12571 1211
rect 1035 -936 12571 -845
rect 754 -1035 962 -983
<< via1 >>
rect 967 1351 12017 1399
rect 959 -248 1003 612
rect 1139 732 1183 1159
rect 1139 -793 1183 -368
rect 1237 -248 1281 612
rect 1417 732 1461 1159
rect 1417 -793 1461 -368
rect 1515 -248 1559 612
rect 1695 732 1739 1159
rect 1695 -793 1739 -368
rect 1793 -248 1837 612
rect 1973 732 2017 1159
rect 1973 -793 2017 -368
rect 2071 -248 2115 612
rect 2251 732 2295 1159
rect 2251 -793 2295 -368
rect 2349 -248 2393 612
rect 2529 732 2573 1159
rect 2529 -793 2573 -368
rect 2627 -248 2671 612
rect 2807 732 2851 1159
rect 2807 -793 2851 -368
rect 2905 -248 2949 612
rect 3085 732 3129 1159
rect 3085 -793 3129 -368
rect 3183 -248 3227 612
rect 3363 732 3407 1159
rect 3363 -793 3407 -368
rect 3461 -248 3505 612
rect 3641 732 3685 1159
rect 3641 -793 3685 -368
rect 3739 -248 3783 612
rect 3919 732 3963 1159
rect 3919 -793 3963 -368
rect 4017 -248 4061 612
rect 4197 732 4241 1159
rect 4197 -793 4241 -368
rect 4295 -248 4339 612
rect 4475 732 4519 1159
rect 4475 -793 4519 -368
rect 4573 -248 4617 612
rect 4753 732 4797 1159
rect 4753 -793 4797 -368
rect 4851 -248 4895 612
rect 5031 732 5075 1159
rect 5031 -793 5075 -368
rect 5129 -248 5173 612
rect 5309 732 5353 1159
rect 5309 -793 5353 -368
rect 5407 -248 5451 612
rect 5587 732 5631 1159
rect 5587 -793 5631 -368
rect 5685 -248 5729 612
rect 5865 732 5909 1159
rect 5865 -793 5909 -368
rect 5963 -248 6007 612
rect 6143 732 6187 1159
rect 6143 -793 6187 -368
rect 6241 -248 6285 612
rect 6421 732 6465 1159
rect 6421 -793 6465 -368
rect 6519 -248 6563 612
rect 6699 732 6743 1159
rect 6699 -793 6743 -368
rect 6797 -248 6841 612
rect 6977 732 7021 1159
rect 6977 -793 7021 -368
rect 7075 -248 7119 612
rect 7255 732 7299 1159
rect 7255 -793 7299 -368
rect 7353 -248 7397 612
rect 7533 732 7577 1159
rect 7533 -793 7577 -368
rect 7631 -248 7675 612
rect 7811 732 7855 1159
rect 7811 -793 7855 -368
rect 7909 -248 7953 612
rect 8089 732 8133 1159
rect 8089 -793 8133 -368
rect 8187 -248 8231 612
rect 8367 732 8411 1159
rect 8367 -793 8411 -368
rect 8465 -248 8509 612
rect 8645 732 8689 1159
rect 8645 -793 8689 -368
rect 8743 -248 8787 612
rect 8923 732 8967 1159
rect 8923 -793 8967 -368
rect 9021 -248 9065 612
rect 9201 732 9245 1159
rect 9201 -793 9245 -368
rect 9299 -248 9343 612
rect 9479 732 9523 1159
rect 9479 -793 9523 -368
rect 9577 -248 9621 612
rect 9757 732 9801 1159
rect 9757 -793 9801 -368
rect 9855 -248 9899 612
rect 10035 732 10079 1159
rect 10035 -793 10079 -368
rect 10133 -248 10177 612
rect 10313 732 10357 1159
rect 10313 -793 10357 -368
rect 10411 -248 10455 612
rect 10591 732 10635 1159
rect 10591 -793 10635 -368
rect 10689 -248 10733 612
rect 10869 732 10913 1159
rect 10869 -793 10913 -368
rect 10967 -248 11011 612
rect 11147 732 11191 1159
rect 11147 -793 11191 -368
rect 11245 -248 11289 612
rect 11425 732 11469 1159
rect 11425 -793 11469 -368
rect 11523 -248 11567 612
rect 11703 732 11747 1159
rect 11703 -793 11747 -368
rect 11801 -248 11845 612
rect 11981 732 12025 1159
rect 11981 -793 12025 -368
rect 12190 -731 12198 1097
rect 12198 -731 12230 1097
rect 12230 -731 12238 1097
rect 967 -1033 12017 -985
<< metal2 >>
rect -586 -1075 -546 1441
rect 914 1421 12499 1441
rect 914 742 934 1421
rect 12479 742 12499 1421
rect 914 732 1139 742
rect 1183 732 1417 742
rect 1461 732 1695 742
rect 1739 732 1973 742
rect 2017 732 2251 742
rect 2295 732 2529 742
rect 2573 732 2807 742
rect 2851 732 3085 742
rect 3129 732 3363 742
rect 3407 732 3641 742
rect 3685 732 3919 742
rect 3963 732 4197 742
rect 4241 732 4475 742
rect 4519 732 4753 742
rect 4797 732 5031 742
rect 5075 732 5309 742
rect 5353 732 5587 742
rect 5631 732 5865 742
rect 5909 732 6143 742
rect 6187 732 6421 742
rect 6465 732 6699 742
rect 6743 732 6977 742
rect 7021 732 7255 742
rect 7299 732 7533 742
rect 7577 732 7811 742
rect 7855 732 8089 742
rect 8133 732 8367 742
rect 8411 732 8645 742
rect 8689 732 8923 742
rect 8967 732 9201 742
rect 9245 732 9479 742
rect 9523 732 9757 742
rect 9801 732 10035 742
rect 10079 732 10313 742
rect 10357 732 10591 742
rect 10635 732 10869 742
rect 10913 732 11147 742
rect 11191 732 11425 742
rect 11469 732 11703 742
rect 11747 732 11981 742
rect 12025 732 12190 742
rect 914 722 12190 732
rect 657 612 12031 622
rect 657 602 959 612
rect 1003 602 1237 612
rect 1281 602 1515 612
rect 1559 602 1793 612
rect 1837 602 2071 612
rect 2115 602 2349 612
rect 2393 602 2627 612
rect 2671 602 2905 612
rect 2949 602 3183 612
rect 3227 602 3461 612
rect 3505 602 3739 612
rect 3783 602 4017 612
rect 4061 602 4295 612
rect 4339 602 4573 612
rect 4617 602 4851 612
rect 4895 602 5129 612
rect 5173 602 5407 612
rect 5451 602 5685 612
rect 5729 602 5963 612
rect 6007 602 6241 612
rect 6285 602 6519 612
rect 6563 602 6797 612
rect 6841 602 7075 612
rect 7119 602 7353 612
rect 7397 602 7631 612
rect 7675 602 7909 612
rect 7953 602 8187 612
rect 8231 602 8465 612
rect 8509 602 8743 612
rect 8787 602 9021 612
rect 9065 602 9299 612
rect 9343 602 9577 612
rect 9621 602 9855 612
rect 9899 602 10133 612
rect 10177 602 10411 612
rect 10455 602 10689 612
rect 10733 602 10967 612
rect 11011 602 11245 612
rect 11289 602 11523 612
rect 11567 602 11801 612
rect 11845 602 12031 612
rect 657 -238 679 602
rect 12011 -238 12031 602
rect 657 -248 959 -238
rect 1003 -248 1237 -238
rect 1281 -248 1515 -238
rect 1559 -248 1793 -238
rect 1837 -248 2071 -238
rect 2115 -248 2349 -238
rect 2393 -248 2627 -238
rect 2671 -248 2905 -238
rect 2949 -248 3183 -238
rect 3227 -248 3461 -238
rect 3505 -248 3739 -238
rect 3783 -248 4017 -238
rect 4061 -248 4295 -238
rect 4339 -248 4573 -238
rect 4617 -248 4851 -238
rect 4895 -248 5129 -238
rect 5173 -248 5407 -238
rect 5451 -248 5685 -238
rect 5729 -248 5963 -238
rect 6007 -248 6241 -238
rect 6285 -248 6519 -238
rect 6563 -248 6797 -238
rect 6841 -248 7075 -238
rect 7119 -248 7353 -238
rect 7397 -248 7631 -238
rect 7675 -248 7909 -238
rect 7953 -248 8187 -238
rect 8231 -248 8465 -238
rect 8509 -248 8743 -238
rect 8787 -248 9021 -238
rect 9065 -248 9299 -238
rect 9343 -248 9577 -238
rect 9621 -248 9855 -238
rect 9899 -248 10133 -238
rect 10177 -248 10411 -238
rect 10455 -248 10689 -238
rect 10733 -248 10967 -238
rect 11011 -248 11245 -238
rect 11289 -248 11523 -238
rect 11567 -248 11801 -238
rect 11845 -248 12031 -238
rect 657 -258 12031 -248
rect 12108 -358 12190 722
rect 914 -368 12190 -358
rect 914 -378 1139 -368
rect 1183 -378 1417 -368
rect 1461 -378 1695 -368
rect 1739 -378 1973 -368
rect 2017 -378 2251 -368
rect 2295 -378 2529 -368
rect 2573 -378 2807 -368
rect 2851 -378 3085 -368
rect 3129 -378 3363 -368
rect 3407 -378 3641 -368
rect 3685 -378 3919 -368
rect 3963 -378 4197 -368
rect 4241 -378 4475 -368
rect 4519 -378 4753 -368
rect 4797 -378 5031 -368
rect 5075 -378 5309 -368
rect 5353 -378 5587 -368
rect 5631 -378 5865 -368
rect 5909 -378 6143 -368
rect 6187 -378 6421 -368
rect 6465 -378 6699 -368
rect 6743 -378 6977 -368
rect 7021 -378 7255 -368
rect 7299 -378 7533 -368
rect 7577 -378 7811 -368
rect 7855 -378 8089 -368
rect 8133 -378 8367 -368
rect 8411 -378 8645 -368
rect 8689 -378 8923 -368
rect 8967 -378 9201 -368
rect 9245 -378 9479 -368
rect 9523 -378 9757 -368
rect 9801 -378 10035 -368
rect 10079 -378 10313 -368
rect 10357 -378 10591 -368
rect 10635 -378 10869 -368
rect 10913 -378 11147 -368
rect 11191 -378 11425 -368
rect 11469 -378 11703 -368
rect 11747 -378 11981 -368
rect 12025 -378 12190 -368
rect 12238 -378 12499 742
rect 914 -1055 934 -378
rect 12479 -1055 12499 -378
rect 914 -1075 12499 -1055
<< via2 >>
rect 934 1399 12479 1421
rect 934 1351 967 1399
rect 967 1351 12017 1399
rect 12017 1351 12479 1399
rect 934 1159 12479 1351
rect 934 742 1139 1159
rect 1139 742 1183 1159
rect 1183 742 1417 1159
rect 1417 742 1461 1159
rect 1461 742 1695 1159
rect 1695 742 1739 1159
rect 1739 742 1973 1159
rect 1973 742 2017 1159
rect 2017 742 2251 1159
rect 2251 742 2295 1159
rect 2295 742 2529 1159
rect 2529 742 2573 1159
rect 2573 742 2807 1159
rect 2807 742 2851 1159
rect 2851 742 3085 1159
rect 3085 742 3129 1159
rect 3129 742 3363 1159
rect 3363 742 3407 1159
rect 3407 742 3641 1159
rect 3641 742 3685 1159
rect 3685 742 3919 1159
rect 3919 742 3963 1159
rect 3963 742 4197 1159
rect 4197 742 4241 1159
rect 4241 742 4475 1159
rect 4475 742 4519 1159
rect 4519 742 4753 1159
rect 4753 742 4797 1159
rect 4797 742 5031 1159
rect 5031 742 5075 1159
rect 5075 742 5309 1159
rect 5309 742 5353 1159
rect 5353 742 5587 1159
rect 5587 742 5631 1159
rect 5631 742 5865 1159
rect 5865 742 5909 1159
rect 5909 742 6143 1159
rect 6143 742 6187 1159
rect 6187 742 6421 1159
rect 6421 742 6465 1159
rect 6465 742 6699 1159
rect 6699 742 6743 1159
rect 6743 742 6977 1159
rect 6977 742 7021 1159
rect 7021 742 7255 1159
rect 7255 742 7299 1159
rect 7299 742 7533 1159
rect 7533 742 7577 1159
rect 7577 742 7811 1159
rect 7811 742 7855 1159
rect 7855 742 8089 1159
rect 8089 742 8133 1159
rect 8133 742 8367 1159
rect 8367 742 8411 1159
rect 8411 742 8645 1159
rect 8645 742 8689 1159
rect 8689 742 8923 1159
rect 8923 742 8967 1159
rect 8967 742 9201 1159
rect 9201 742 9245 1159
rect 9245 742 9479 1159
rect 9479 742 9523 1159
rect 9523 742 9757 1159
rect 9757 742 9801 1159
rect 9801 742 10035 1159
rect 10035 742 10079 1159
rect 10079 742 10313 1159
rect 10313 742 10357 1159
rect 10357 742 10591 1159
rect 10591 742 10635 1159
rect 10635 742 10869 1159
rect 10869 742 10913 1159
rect 10913 742 11147 1159
rect 11147 742 11191 1159
rect 11191 742 11425 1159
rect 11425 742 11469 1159
rect 11469 742 11703 1159
rect 11703 742 11747 1159
rect 11747 742 11981 1159
rect 11981 742 12025 1159
rect 12025 1097 12479 1159
rect 12025 742 12190 1097
rect 12190 742 12238 1097
rect 12238 742 12479 1097
rect 679 -238 959 602
rect 959 -238 1003 602
rect 1003 -238 1237 602
rect 1237 -238 1281 602
rect 1281 -238 1515 602
rect 1515 -238 1559 602
rect 1559 -238 1793 602
rect 1793 -238 1837 602
rect 1837 -238 2071 602
rect 2071 -238 2115 602
rect 2115 -238 2349 602
rect 2349 -238 2393 602
rect 2393 -238 2627 602
rect 2627 -238 2671 602
rect 2671 -238 2905 602
rect 2905 -238 2949 602
rect 2949 -238 3183 602
rect 3183 -238 3227 602
rect 3227 -238 3461 602
rect 3461 -238 3505 602
rect 3505 -238 3739 602
rect 3739 -238 3783 602
rect 3783 -238 4017 602
rect 4017 -238 4061 602
rect 4061 -238 4295 602
rect 4295 -238 4339 602
rect 4339 -238 4573 602
rect 4573 -238 4617 602
rect 4617 -238 4851 602
rect 4851 -238 4895 602
rect 4895 -238 5129 602
rect 5129 -238 5173 602
rect 5173 -238 5407 602
rect 5407 -238 5451 602
rect 5451 -238 5685 602
rect 5685 -238 5729 602
rect 5729 -238 5963 602
rect 5963 -238 6007 602
rect 6007 -238 6241 602
rect 6241 -238 6285 602
rect 6285 -238 6519 602
rect 6519 -238 6563 602
rect 6563 -238 6797 602
rect 6797 -238 6841 602
rect 6841 -238 7075 602
rect 7075 -238 7119 602
rect 7119 -238 7353 602
rect 7353 -238 7397 602
rect 7397 -238 7631 602
rect 7631 -238 7675 602
rect 7675 -238 7909 602
rect 7909 -238 7953 602
rect 7953 -238 8187 602
rect 8187 -238 8231 602
rect 8231 -238 8465 602
rect 8465 -238 8509 602
rect 8509 -238 8743 602
rect 8743 -238 8787 602
rect 8787 -238 9021 602
rect 9021 -238 9065 602
rect 9065 -238 9299 602
rect 9299 -238 9343 602
rect 9343 -238 9577 602
rect 9577 -238 9621 602
rect 9621 -238 9855 602
rect 9855 -238 9899 602
rect 9899 -238 10133 602
rect 10133 -238 10177 602
rect 10177 -238 10411 602
rect 10411 -238 10455 602
rect 10455 -238 10689 602
rect 10689 -238 10733 602
rect 10733 -238 10967 602
rect 10967 -238 11011 602
rect 11011 -238 11245 602
rect 11245 -238 11289 602
rect 11289 -238 11523 602
rect 11523 -238 11567 602
rect 11567 -238 11801 602
rect 11801 -238 11845 602
rect 11845 -238 12011 602
rect 934 -793 1139 -378
rect 1139 -793 1183 -378
rect 1183 -793 1417 -378
rect 1417 -793 1461 -378
rect 1461 -793 1695 -378
rect 1695 -793 1739 -378
rect 1739 -793 1973 -378
rect 1973 -793 2017 -378
rect 2017 -793 2251 -378
rect 2251 -793 2295 -378
rect 2295 -793 2529 -378
rect 2529 -793 2573 -378
rect 2573 -793 2807 -378
rect 2807 -793 2851 -378
rect 2851 -793 3085 -378
rect 3085 -793 3129 -378
rect 3129 -793 3363 -378
rect 3363 -793 3407 -378
rect 3407 -793 3641 -378
rect 3641 -793 3685 -378
rect 3685 -793 3919 -378
rect 3919 -793 3963 -378
rect 3963 -793 4197 -378
rect 4197 -793 4241 -378
rect 4241 -793 4475 -378
rect 4475 -793 4519 -378
rect 4519 -793 4753 -378
rect 4753 -793 4797 -378
rect 4797 -793 5031 -378
rect 5031 -793 5075 -378
rect 5075 -793 5309 -378
rect 5309 -793 5353 -378
rect 5353 -793 5587 -378
rect 5587 -793 5631 -378
rect 5631 -793 5865 -378
rect 5865 -793 5909 -378
rect 5909 -793 6143 -378
rect 6143 -793 6187 -378
rect 6187 -793 6421 -378
rect 6421 -793 6465 -378
rect 6465 -793 6699 -378
rect 6699 -793 6743 -378
rect 6743 -793 6977 -378
rect 6977 -793 7021 -378
rect 7021 -793 7255 -378
rect 7255 -793 7299 -378
rect 7299 -793 7533 -378
rect 7533 -793 7577 -378
rect 7577 -793 7811 -378
rect 7811 -793 7855 -378
rect 7855 -793 8089 -378
rect 8089 -793 8133 -378
rect 8133 -793 8367 -378
rect 8367 -793 8411 -378
rect 8411 -793 8645 -378
rect 8645 -793 8689 -378
rect 8689 -793 8923 -378
rect 8923 -793 8967 -378
rect 8967 -793 9201 -378
rect 9201 -793 9245 -378
rect 9245 -793 9479 -378
rect 9479 -793 9523 -378
rect 9523 -793 9757 -378
rect 9757 -793 9801 -378
rect 9801 -793 10035 -378
rect 10035 -793 10079 -378
rect 10079 -793 10313 -378
rect 10313 -793 10357 -378
rect 10357 -793 10591 -378
rect 10591 -793 10635 -378
rect 10635 -793 10869 -378
rect 10869 -793 10913 -378
rect 10913 -793 11147 -378
rect 11147 -793 11191 -378
rect 11191 -793 11425 -378
rect 11425 -793 11469 -378
rect 11469 -793 11703 -378
rect 11703 -793 11747 -378
rect 11747 -793 11981 -378
rect 11981 -793 12025 -378
rect 12025 -731 12190 -378
rect 12190 -731 12238 -378
rect 12238 -731 12479 -378
rect 12025 -793 12479 -731
rect 934 -985 12479 -793
rect 934 -1033 967 -985
rect 967 -1033 12017 -985
rect 12017 -1033 12479 -985
rect 934 -1055 12479 -1033
<< metal3 >>
rect -586 -1075 -546 1441
rect 914 1421 12499 1441
rect 914 742 934 1421
rect 12479 742 12499 1421
rect 914 722 12499 742
rect 657 602 12031 622
rect 657 -238 679 602
rect 12011 -238 12031 602
rect 657 -258 12031 -238
rect 12108 -358 12499 722
rect 914 -378 12499 -358
rect 914 -1055 934 -378
rect 12479 -1055 12499 -378
rect 914 -1075 12499 -1055
use fuse_prim  fuse_prim_0
timestamp 1757368577
transform 1 0 0 0 1 0
box -586 -1075 657 1441
use hvnmos_LATSBM  hvnmos_LATSBM_0
timestamp 1757367233
transform 1 0 1071 0 1 183
box -118 -1222 10960 1222
<< labels >>
flabel metal3 12340 -1075 12499 1441 0 FreeSans 800 0 0 0 VSS
port 0 nsew
flabel metal1 12512 -936 12571 1302 0 FreeSans 800 0 0 0 SEL
port 2 nsew
flabel metal3 -586 -1075 -566 1441 0 FreeSans 800 0 0 0 VDD
port 1 nsew
<< end >>
