magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752864670
<< error_p >>
rect -36 160 -26 170
rect 26 160 36 170
rect -46 150 46 160
rect -36 138 36 150
rect -46 128 46 138
rect -36 118 -26 128
rect 26 118 36 128
rect -104 86 -94 96
rect -82 86 -72 96
rect 72 86 82 96
rect 94 86 104 96
rect -114 76 -104 86
rect -72 76 -62 86
rect 62 76 72 86
rect 104 76 114 86
rect -114 -86 -104 -76
rect -72 -86 -62 -76
rect 62 -86 72 -76
rect 104 -86 114 -76
rect -104 -96 -94 -86
rect -82 -96 -72 -86
rect 72 -96 82 -86
rect 94 -96 104 -86
rect -36 -128 -26 -118
rect 26 -128 36 -118
rect -46 -138 46 -128
rect -36 -150 36 -138
rect -46 -160 46 -150
rect -36 -170 -26 -160
rect 26 -170 36 -160
<< nmos >>
rect -50 -100 50 100
<< ndiff >>
rect -118 86 -50 100
rect -118 -86 -104 86
rect -72 -86 -50 86
rect -118 -100 -50 -86
rect 50 86 118 100
rect 50 -86 72 86
rect 104 -86 118 86
rect 50 -100 118 -86
<< ndiffc >>
rect -104 -86 -72 86
rect 72 -86 104 86
<< psubdiff >>
rect -241 262 241 276
rect -241 230 -167 262
rect 167 230 241 262
rect -241 216 241 230
rect -241 202 -181 216
rect -241 -202 -227 202
rect -195 -202 -181 202
rect 181 202 241 216
rect -241 -216 -181 -202
rect 181 -202 195 202
rect 227 -202 241 202
rect 181 -216 241 -202
rect -241 -230 241 -216
rect -241 -262 -167 -230
rect 167 -262 241 -230
rect -241 -276 241 -262
<< psubdiffcont >>
rect -167 230 167 262
rect -227 -202 -195 202
rect 195 -202 227 202
rect -167 -262 167 -230
<< poly >>
rect -50 160 50 174
rect -50 128 -36 160
rect 36 128 50 160
rect -50 100 50 128
rect -50 -128 50 -100
rect -50 -160 -36 -128
rect 36 -160 50 -128
rect -50 -174 50 -160
<< polycont >>
rect -36 128 36 160
rect -36 -160 36 -128
<< metal1 >>
rect -237 262 237 272
rect -237 230 -167 262
rect 167 230 237 262
rect -237 220 237 230
rect -237 202 -185 220
rect -237 -202 -227 202
rect -195 -202 -185 202
rect 185 202 237 220
rect -237 -220 -185 -202
rect 185 -202 195 202
rect 227 -202 237 202
rect 185 -220 237 -202
rect -237 -230 237 -220
rect -237 -262 -167 -230
rect 167 -262 237 -230
rect -237 -272 237 -262
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 1 l 0.5 nf 1 nx 1 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 1
<< end >>
