magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 443 2640 834
rect -48 370 454 443
rect -48 350 187 370
rect 1044 367 2640 443
rect 1044 348 1463 367
rect 2131 350 2640 367
<< pwell >>
rect 669 358 1008 382
rect 223 237 426 333
rect 647 309 1008 358
rect 647 301 1435 309
rect 647 246 1790 301
rect 647 237 706 246
rect 223 224 706 237
rect 12 56 706 224
rect 1081 224 1790 246
rect 2225 224 2541 288
rect 1081 56 2541 224
rect -26 -56 2618 56
<< nmos >>
rect 106 114 132 198
rect 190 114 216 198
rect 306 159 332 307
rect 741 272 767 356
rect 843 272 869 356
rect 524 127 550 211
rect 586 127 612 211
rect 1175 135 1201 283
rect 1315 135 1341 283
rect 1557 191 1583 275
rect 1664 127 1690 275
rect 1874 114 1900 198
rect 1976 114 2002 198
rect 2038 114 2064 198
rect 2319 114 2345 262
rect 2421 114 2447 262
<< pmos >>
rect 106 432 132 516
rect 208 432 234 516
rect 298 432 324 632
rect 508 505 534 589
rect 655 505 681 589
rect 741 505 767 589
rect 843 505 869 589
rect 1175 410 1201 634
rect 1315 410 1341 634
rect 1607 429 1633 629
rect 1759 429 1785 513
rect 1874 429 1900 513
rect 1976 429 2002 513
rect 2078 429 2104 513
rect 2319 412 2345 636
rect 2421 412 2447 636
<< ndiff >>
rect 249 198 306 307
rect 38 160 106 198
rect 38 128 52 160
rect 84 128 106 160
rect 38 114 106 128
rect 132 114 190 198
rect 216 160 306 198
rect 216 128 238 160
rect 270 159 306 160
rect 332 208 400 307
rect 695 332 741 356
rect 673 318 741 332
rect 673 286 687 318
rect 719 286 741 318
rect 673 272 741 286
rect 767 342 843 356
rect 767 310 789 342
rect 821 310 843 342
rect 767 272 843 310
rect 869 330 982 356
rect 869 298 936 330
rect 968 298 982 330
rect 869 272 982 298
rect 332 176 354 208
rect 386 176 400 208
rect 332 159 400 176
rect 443 173 524 211
rect 270 128 289 159
rect 216 114 289 128
rect 443 141 457 173
rect 489 141 524 173
rect 443 127 524 141
rect 550 127 586 211
rect 612 191 680 211
rect 612 159 634 191
rect 666 159 680 191
rect 612 127 680 159
rect 1107 226 1175 283
rect 1107 194 1121 226
rect 1153 194 1175 226
rect 1107 135 1175 194
rect 1201 135 1315 283
rect 1341 226 1409 283
rect 1341 194 1363 226
rect 1395 194 1409 226
rect 1341 135 1409 194
rect 1489 247 1557 275
rect 1489 215 1503 247
rect 1535 215 1557 247
rect 1489 191 1557 215
rect 1583 261 1664 275
rect 1583 229 1605 261
rect 1637 229 1664 261
rect 1583 191 1664 229
rect 1215 36 1301 135
rect 1612 127 1664 191
rect 1690 127 1764 275
rect 2251 228 2319 262
rect 1704 125 1764 127
rect 1704 93 1718 125
rect 1750 93 1764 125
rect 1806 160 1874 198
rect 1806 128 1820 160
rect 1852 128 1874 160
rect 1806 114 1874 128
rect 1900 160 1976 198
rect 1900 128 1922 160
rect 1954 128 1976 160
rect 1900 114 1976 128
rect 2002 114 2038 198
rect 2064 160 2132 198
rect 2064 128 2086 160
rect 2118 128 2132 160
rect 2064 114 2132 128
rect 2251 196 2265 228
rect 2297 196 2319 228
rect 2251 160 2319 196
rect 2251 128 2265 160
rect 2297 128 2319 160
rect 2251 114 2319 128
rect 2345 228 2421 262
rect 2345 196 2367 228
rect 2399 196 2421 228
rect 2345 160 2421 196
rect 2345 128 2367 160
rect 2399 128 2421 160
rect 2345 114 2421 128
rect 2447 228 2515 262
rect 2447 196 2469 228
rect 2501 196 2515 228
rect 2447 160 2515 196
rect 2447 128 2469 160
rect 2501 128 2515 160
rect 2447 114 2515 128
rect 1704 78 1764 93
<< pdiff >>
rect 38 656 283 679
rect 38 624 53 656
rect 85 632 283 656
rect 85 624 298 632
rect 38 602 298 624
rect 248 516 298 602
rect 38 490 106 516
rect 38 458 52 490
rect 84 458 106 490
rect 38 432 106 458
rect 132 490 208 516
rect 132 458 154 490
rect 186 458 208 490
rect 132 432 208 458
rect 234 432 298 516
rect 324 542 392 632
rect 576 614 636 628
rect 576 589 590 614
rect 324 510 346 542
rect 378 510 392 542
rect 324 432 392 510
rect 438 570 508 589
rect 438 538 452 570
rect 484 538 508 570
rect 438 505 508 538
rect 534 582 590 589
rect 622 589 636 614
rect 1215 634 1301 720
rect 622 582 655 589
rect 534 505 655 582
rect 681 505 741 589
rect 767 551 843 589
rect 767 519 789 551
rect 821 519 843 551
rect 767 505 843 519
rect 869 573 937 589
rect 869 541 891 573
rect 923 541 937 573
rect 869 505 937 541
rect 1106 540 1175 634
rect 1106 508 1120 540
rect 1152 508 1175 540
rect 1106 456 1175 508
rect 1106 424 1120 456
rect 1152 424 1175 456
rect 1106 410 1175 424
rect 1201 410 1315 634
rect 1341 456 1414 634
rect 1539 475 1607 629
rect 1341 424 1368 456
rect 1400 424 1414 456
rect 1341 410 1414 424
rect 1539 443 1553 475
rect 1585 443 1607 475
rect 1539 429 1607 443
rect 1633 513 1683 629
rect 1914 513 1962 720
rect 2118 623 2178 720
rect 2118 591 2132 623
rect 2164 591 2178 623
rect 2118 555 2178 591
rect 2118 523 2132 555
rect 2164 523 2178 555
rect 2118 513 2178 523
rect 1633 487 1759 513
rect 1633 455 1705 487
rect 1737 455 1759 487
rect 1633 429 1759 455
rect 1785 429 1874 513
rect 1900 429 1976 513
rect 2002 487 2078 513
rect 2002 455 2024 487
rect 2056 455 2078 487
rect 2002 429 2078 455
rect 2104 487 2178 513
rect 2104 455 2132 487
rect 2164 455 2178 487
rect 2104 429 2178 455
rect 2250 621 2319 636
rect 2250 589 2264 621
rect 2296 589 2319 621
rect 2250 540 2319 589
rect 2250 508 2264 540
rect 2296 508 2319 540
rect 2250 459 2319 508
rect 2250 427 2264 459
rect 2296 427 2319 459
rect 2250 412 2319 427
rect 2345 621 2421 636
rect 2345 589 2367 621
rect 2399 589 2421 621
rect 2345 540 2421 589
rect 2345 508 2367 540
rect 2399 508 2421 540
rect 2345 459 2421 508
rect 2345 427 2367 459
rect 2399 427 2421 459
rect 2345 412 2421 427
rect 2447 621 2515 636
rect 2447 589 2469 621
rect 2501 589 2515 621
rect 2447 540 2515 589
rect 2447 508 2469 540
rect 2501 508 2515 540
rect 2447 459 2515 508
rect 2447 427 2469 459
rect 2501 427 2515 459
rect 2447 412 2515 427
<< ndiffc >>
rect 52 128 84 160
rect 238 128 270 160
rect 687 286 719 318
rect 789 310 821 342
rect 936 298 968 330
rect 354 176 386 208
rect 457 141 489 173
rect 634 159 666 191
rect 1121 194 1153 226
rect 1363 194 1395 226
rect 1503 215 1535 247
rect 1605 229 1637 261
rect 1718 93 1750 125
rect 1820 128 1852 160
rect 1922 128 1954 160
rect 2086 128 2118 160
rect 2265 196 2297 228
rect 2265 128 2297 160
rect 2367 196 2399 228
rect 2367 128 2399 160
rect 2469 196 2501 228
rect 2469 128 2501 160
<< pdiffc >>
rect 53 624 85 656
rect 52 458 84 490
rect 154 458 186 490
rect 346 510 378 542
rect 452 538 484 570
rect 590 582 622 614
rect 789 519 821 551
rect 891 541 923 573
rect 1120 508 1152 540
rect 1120 424 1152 456
rect 1368 424 1400 456
rect 1553 443 1585 475
rect 2132 591 2164 623
rect 2132 523 2164 555
rect 1705 455 1737 487
rect 2024 455 2056 487
rect 2132 455 2164 487
rect 2264 589 2296 621
rect 2264 508 2296 540
rect 2264 427 2296 459
rect 2367 589 2399 621
rect 2367 508 2399 540
rect 2367 427 2399 459
rect 2469 589 2501 621
rect 2469 508 2501 540
rect 2469 427 2501 459
<< psubdiff >>
rect 1215 30 1301 36
rect 0 16 2592 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2528 16
rect 2560 -16 2592 16
rect 0 -30 2592 -16
<< nsubdiff >>
rect 0 772 2592 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2528 772
rect 2560 740 2592 772
rect 0 726 2592 740
rect 1215 720 1301 726
rect 1914 720 1962 726
rect 2118 720 2178 726
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
rect 1280 -16 1312 16
rect 1376 -16 1408 16
rect 1472 -16 1504 16
rect 1568 -16 1600 16
rect 1664 -16 1696 16
rect 1760 -16 1792 16
rect 1856 -16 1888 16
rect 1952 -16 1984 16
rect 2048 -16 2080 16
rect 2144 -16 2176 16
rect 2240 -16 2272 16
rect 2336 -16 2368 16
rect 2432 -16 2464 16
rect 2528 -16 2560 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
rect 1280 740 1312 772
rect 1376 740 1408 772
rect 1472 740 1504 772
rect 1568 740 1600 772
rect 1664 740 1696 772
rect 1760 740 1792 772
rect 1856 740 1888 772
rect 1952 740 1984 772
rect 2048 740 2080 772
rect 2144 740 2176 772
rect 2240 740 2272 772
rect 2336 740 2368 772
rect 2432 740 2464 772
rect 2528 740 2560 772
<< poly >>
rect 298 632 324 668
rect 508 661 1027 687
rect 106 516 132 552
rect 208 516 234 552
rect 508 589 534 661
rect 967 647 1027 661
rect 655 589 681 625
rect 741 589 767 625
rect 843 589 869 625
rect 967 615 981 647
rect 1013 615 1027 647
rect 1175 634 1201 670
rect 1315 634 1341 670
rect 967 601 1027 615
rect 106 351 132 432
rect 208 396 234 432
rect 47 337 132 351
rect 47 305 61 337
rect 93 305 132 337
rect 47 291 132 305
rect 106 198 132 291
rect 190 337 234 396
rect 298 397 324 432
rect 508 397 534 505
rect 655 397 681 505
rect 298 383 373 397
rect 298 351 327 383
rect 359 351 373 383
rect 298 337 373 351
rect 490 383 550 397
rect 490 351 504 383
rect 536 351 550 383
rect 490 337 550 351
rect 190 198 216 337
rect 306 307 332 337
rect 524 211 550 337
rect 586 383 681 397
rect 586 351 600 383
rect 632 371 681 383
rect 632 351 646 371
rect 741 356 767 505
rect 843 488 869 505
rect 843 474 1027 488
rect 843 458 981 474
rect 843 356 869 458
rect 967 442 981 458
rect 1013 442 1027 474
rect 967 428 1027 442
rect 1607 629 1633 665
rect 1449 456 1509 470
rect 1449 424 1463 456
rect 1495 424 1509 456
rect 1759 513 1785 549
rect 1874 513 1900 549
rect 1976 647 2036 661
rect 1976 615 1990 647
rect 2022 615 2036 647
rect 1976 601 2036 615
rect 2319 636 2345 672
rect 2421 636 2447 672
rect 1976 513 2002 601
rect 2078 513 2104 549
rect 1449 414 1509 424
rect 1607 414 1633 429
rect 1175 371 1201 410
rect 1141 357 1201 371
rect 586 337 646 351
rect 586 211 612 337
rect 1141 325 1155 357
rect 1187 325 1201 357
rect 1141 311 1201 325
rect 1175 283 1201 311
rect 1315 371 1341 410
rect 1449 384 1633 414
rect 1315 357 1375 371
rect 1315 325 1329 357
rect 1361 325 1375 357
rect 1315 311 1375 325
rect 1315 283 1341 311
rect 306 123 332 159
rect 106 78 132 114
rect 190 86 216 114
rect 524 86 550 127
rect 190 59 550 86
rect 586 85 612 127
rect 741 121 767 272
rect 843 236 869 272
rect 1557 275 1583 384
rect 1759 361 1785 429
rect 1874 394 1900 429
rect 1664 347 1785 361
rect 1664 315 1678 347
rect 1710 332 1785 347
rect 1840 380 1900 394
rect 1840 348 1854 380
rect 1886 348 1900 380
rect 1840 334 1900 348
rect 1710 315 1724 332
rect 1664 301 1724 315
rect 1664 275 1690 301
rect 1557 153 1583 191
rect 1175 121 1201 135
rect 741 93 1201 121
rect 1315 99 1341 135
rect 1874 198 1900 334
rect 1976 198 2002 429
rect 2078 327 2104 429
rect 2319 327 2345 412
rect 2421 349 2447 412
rect 2038 313 2345 327
rect 2038 281 2052 313
rect 2084 290 2345 313
rect 2084 281 2098 290
rect 2038 267 2098 281
rect 2038 198 2064 267
rect 2319 262 2345 290
rect 2404 335 2464 349
rect 2404 303 2418 335
rect 2450 303 2464 335
rect 2404 289 2464 303
rect 2421 262 2447 289
rect 1664 89 1690 127
rect 1874 78 1900 114
rect 1976 78 2002 114
rect 2038 78 2064 114
rect 2319 78 2345 114
rect 2421 78 2447 114
<< polycont >>
rect 981 615 1013 647
rect 61 305 93 337
rect 327 351 359 383
rect 504 351 536 383
rect 600 351 632 383
rect 981 442 1013 474
rect 1463 424 1495 456
rect 1990 615 2022 647
rect 1155 325 1187 357
rect 1329 325 1361 357
rect 1678 315 1710 347
rect 1854 348 1886 380
rect 2052 281 2084 313
rect 2418 303 2450 335
<< metal1 >>
rect 0 772 2592 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2528 772
rect 2560 740 2592 772
rect 0 712 2592 740
rect 43 656 95 712
rect 43 624 53 656
rect 85 624 95 656
rect 43 490 95 624
rect 157 616 553 648
rect 157 500 190 616
rect 449 570 485 580
rect 240 542 388 552
rect 240 510 346 542
rect 378 510 388 542
rect 240 500 388 510
rect 449 538 452 570
rect 484 538 485 570
rect 43 458 52 490
rect 84 458 95 490
rect 43 448 95 458
rect 144 490 196 500
rect 144 458 154 490
rect 186 458 196 490
rect 144 448 196 458
rect 51 337 120 378
rect 51 305 61 337
rect 93 305 120 337
rect 51 214 120 305
rect 157 170 190 448
rect 240 262 272 500
rect 449 463 485 538
rect 521 536 553 616
rect 589 614 623 712
rect 589 582 590 614
rect 622 582 623 614
rect 589 572 623 582
rect 673 616 901 648
rect 673 536 707 616
rect 864 583 901 616
rect 971 647 1023 657
rect 1982 647 2032 657
rect 971 615 981 647
rect 1013 615 1990 647
rect 2022 615 2032 647
rect 971 605 1023 615
rect 1982 605 2032 615
rect 2122 623 2175 712
rect 2122 591 2132 623
rect 2164 591 2175 623
rect 864 573 933 583
rect 521 504 707 536
rect 779 551 823 561
rect 779 519 789 551
rect 821 519 823 551
rect 779 463 823 519
rect 449 461 823 463
rect 317 429 823 461
rect 317 383 369 429
rect 317 351 327 383
rect 359 351 369 383
rect 317 341 369 351
rect 429 383 550 393
rect 429 351 504 383
rect 536 351 550 383
rect 429 302 550 351
rect 590 383 642 393
rect 590 351 600 383
rect 632 351 642 383
rect 590 341 642 351
rect 779 342 823 429
rect 590 262 622 341
rect 240 230 622 262
rect 677 318 729 328
rect 677 286 687 318
rect 719 286 729 318
rect 779 310 789 342
rect 821 310 823 342
rect 779 300 823 310
rect 864 541 891 573
rect 923 541 933 573
rect 864 531 933 541
rect 1110 540 1655 560
rect 677 264 729 286
rect 864 264 896 531
rect 1110 508 1120 540
rect 1152 526 1655 540
rect 1152 508 1162 526
rect 1110 484 1162 508
rect 971 474 1162 484
rect 971 442 981 474
rect 1013 456 1162 474
rect 1549 475 1587 485
rect 1013 442 1120 456
rect 971 432 1120 442
rect 1029 424 1120 432
rect 1152 424 1162 456
rect 1029 414 1162 424
rect 1204 456 1505 466
rect 1204 424 1368 456
rect 1400 424 1463 456
rect 1495 424 1505 456
rect 1204 414 1505 424
rect 1549 443 1553 475
rect 1585 443 1587 475
rect 932 330 981 340
rect 932 298 936 330
rect 968 298 981 330
rect 932 288 981 298
rect 677 232 896 264
rect 344 208 396 230
rect 344 176 354 208
rect 386 176 396 208
rect 42 160 190 170
rect 42 128 52 160
rect 84 128 190 160
rect 42 118 190 128
rect 228 160 282 170
rect 344 163 396 176
rect 447 173 499 183
rect 228 128 238 160
rect 270 128 282 160
rect 228 44 282 128
rect 447 141 457 173
rect 489 141 499 173
rect 447 44 499 141
rect 541 121 575 230
rect 945 192 981 288
rect 624 191 981 192
rect 624 159 634 191
rect 666 159 981 191
rect 1029 236 1084 414
rect 1204 367 1236 414
rect 1145 357 1236 367
rect 1145 325 1155 357
rect 1187 325 1236 357
rect 1145 315 1236 325
rect 1029 226 1163 236
rect 1029 194 1121 226
rect 1153 194 1163 226
rect 1204 228 1236 315
rect 1290 357 1398 368
rect 1290 325 1329 357
rect 1361 325 1398 357
rect 1549 345 1587 443
rect 1290 304 1398 325
rect 1434 311 1587 345
rect 1623 357 1655 526
rect 2122 555 2175 591
rect 2122 523 2132 555
rect 2164 523 2175 555
rect 1695 487 1790 497
rect 1695 455 1705 487
rect 1737 455 1790 487
rect 1695 445 1790 455
rect 1623 347 1720 357
rect 1623 315 1678 347
rect 1710 315 1720 347
rect 1351 228 1398 236
rect 1204 226 1398 228
rect 1204 196 1363 226
rect 1029 184 1163 194
rect 1351 194 1363 196
rect 1395 194 1398 226
rect 1351 184 1398 194
rect 624 157 981 159
rect 1434 121 1466 311
rect 1623 305 1720 315
rect 1758 302 1790 445
rect 2014 487 2066 499
rect 2014 455 2024 487
rect 2056 455 2066 487
rect 2014 404 2066 455
rect 2122 487 2175 523
rect 2122 455 2132 487
rect 2164 455 2175 487
rect 2122 445 2175 455
rect 2255 621 2307 631
rect 2255 589 2264 621
rect 2296 589 2307 621
rect 2255 540 2307 589
rect 2255 508 2264 540
rect 2296 508 2307 540
rect 2255 459 2307 508
rect 2255 427 2264 459
rect 2296 427 2307 459
rect 1844 380 2167 404
rect 1844 348 1854 380
rect 1886 372 2167 380
rect 1886 348 1896 372
rect 1844 338 1896 348
rect 2033 313 2094 325
rect 2033 302 2052 313
rect 1758 281 2052 302
rect 2084 281 2094 313
rect 1758 270 2094 281
rect 1758 263 1794 270
rect 1502 247 1545 262
rect 1502 215 1503 247
rect 1535 215 1545 247
rect 1592 261 1794 263
rect 1592 229 1605 261
rect 1637 229 1794 261
rect 2135 238 2167 372
rect 1502 193 1545 215
rect 2114 206 2167 238
rect 2255 342 2307 427
rect 2357 621 2409 712
rect 2357 589 2367 621
rect 2399 589 2409 621
rect 2357 540 2409 589
rect 2357 508 2367 540
rect 2399 508 2409 540
rect 2357 459 2409 508
rect 2357 427 2367 459
rect 2399 427 2409 459
rect 2357 420 2409 427
rect 2459 621 2542 631
rect 2459 589 2469 621
rect 2501 589 2542 621
rect 2459 540 2542 589
rect 2459 508 2469 540
rect 2501 508 2542 540
rect 2459 459 2542 508
rect 2459 427 2469 459
rect 2501 427 2542 459
rect 2459 419 2542 427
rect 2404 342 2464 349
rect 2255 335 2464 342
rect 2255 303 2418 335
rect 2450 303 2464 335
rect 2255 297 2464 303
rect 2255 228 2307 297
rect 2404 289 2464 297
rect 2500 238 2542 419
rect 1502 161 1862 193
rect 2114 177 2146 206
rect 1810 160 1862 161
rect 1810 128 1820 160
rect 1852 128 1862 160
rect 1708 121 1718 125
rect 541 93 1718 121
rect 1750 93 1760 125
rect 1810 118 1862 128
rect 1912 160 1964 170
rect 1912 128 1922 160
rect 1954 128 1964 160
rect 541 88 1760 93
rect 1912 44 1964 128
rect 2076 160 2146 177
rect 2076 128 2086 160
rect 2118 128 2146 160
rect 2076 125 2146 128
rect 2255 196 2265 228
rect 2297 196 2307 228
rect 2255 160 2307 196
rect 2255 128 2265 160
rect 2297 128 2307 160
rect 2255 118 2307 128
rect 2357 228 2409 238
rect 2357 196 2367 228
rect 2399 196 2409 228
rect 2357 160 2409 196
rect 2357 128 2367 160
rect 2399 128 2409 160
rect 2357 44 2409 128
rect 2455 228 2542 238
rect 2455 196 2469 228
rect 2501 196 2542 228
rect 2455 160 2542 196
rect 2455 128 2469 160
rect 2501 128 2542 160
rect 2455 118 2542 128
rect 0 16 2592 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2528 16
rect 2560 -16 2592 16
rect 0 -44 2592 -16
<< labels >>
flabel metal1 s 1290 304 1398 368 0 FreeSans 400 0 0 0 CLK
port 2 nsew
flabel metal1 s 0 -44 2592 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 51 214 120 378 0 FreeSans 340 0 0 0 D
port 4 nsew
flabel metal1 s 2459 419 2542 631 0 FreeSans 340 0 0 0 Q
port 5 nsew
flabel metal1 s 0 712 2592 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s 429 302 550 393 0 FreeSans 400 0 0 0 RESET_B
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 756
string GDS_END 108338
string GDS_FILE 6_final.gds
string GDS_START 94454
<< end >>
