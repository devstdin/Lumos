magic
tech ihp-sg13g2
timestamp 1748556962
<< error_p >>
rect -48 1036 48 1041
rect -48 1020 -43 1036
rect 43 1020 48 1036
rect -48 1015 48 1020
rect 70 1036 166 1041
rect 70 1020 75 1036
rect 161 1020 166 1036
rect 70 1015 166 1020
rect 188 1036 284 1041
rect 188 1020 193 1036
rect 279 1020 284 1036
rect 188 1015 284 1020
rect 306 1036 402 1041
rect 306 1020 311 1036
rect 397 1020 402 1036
rect 306 1015 402 1020
rect -48 -1020 48 -1015
rect -48 -1036 -43 -1020
rect 43 -1036 48 -1020
rect -48 -1041 48 -1036
rect 70 -1020 166 -1015
rect 70 -1036 75 -1020
rect 161 -1036 166 -1020
rect 70 -1041 166 -1036
rect 188 -1020 284 -1015
rect 188 -1036 193 -1020
rect 279 -1036 284 -1020
rect 188 -1041 284 -1036
rect 306 -1020 402 -1015
rect 306 -1036 311 -1020
rect 397 -1036 402 -1020
rect 306 -1041 402 -1036
<< psubdiff >>
rect -140 1126 494 1133
rect -140 1110 -103 1126
rect 457 1110 494 1126
rect -140 1103 494 1110
rect -140 1096 -110 1103
rect -140 -1096 -133 1096
rect -117 -1096 -110 1096
rect 464 1096 494 1103
rect -140 -1103 -110 -1096
rect 464 -1096 471 1096
rect 487 -1096 494 1096
rect 464 -1103 494 -1096
rect -140 -1110 494 -1103
rect -140 -1126 -103 -1110
rect 457 -1126 494 -1110
rect -140 -1133 494 -1126
<< psubdiffcont >>
rect -103 1110 457 1126
rect -133 -1096 -117 1096
rect 471 -1096 487 1096
rect -103 -1126 457 -1110
<< poly >>
rect -50 1036 50 1043
rect -50 1020 -43 1036
rect 43 1020 50 1036
rect -50 1000 50 1020
rect -50 -1020 50 -1000
rect -50 -1036 -43 -1020
rect 43 -1036 50 -1020
rect -50 -1043 50 -1036
rect 68 1036 168 1043
rect 68 1020 75 1036
rect 161 1020 168 1036
rect 68 1000 168 1020
rect 68 -1020 168 -1000
rect 68 -1036 75 -1020
rect 161 -1036 168 -1020
rect 68 -1043 168 -1036
rect 186 1036 286 1043
rect 186 1020 193 1036
rect 279 1020 286 1036
rect 186 1000 286 1020
rect 186 -1020 286 -1000
rect 186 -1036 193 -1020
rect 279 -1036 286 -1020
rect 186 -1043 286 -1036
rect 304 1036 404 1043
rect 304 1020 311 1036
rect 397 1020 404 1036
rect 304 1000 404 1020
rect 304 -1020 404 -1000
rect 304 -1036 311 -1020
rect 397 -1036 404 -1020
rect 304 -1043 404 -1036
<< polycont >>
rect -43 1020 43 1036
rect -43 -1036 43 -1020
rect 75 1020 161 1036
rect 75 -1036 161 -1020
rect 193 1020 279 1036
rect 193 -1036 279 -1020
rect 311 1020 397 1036
rect 311 -1036 397 -1020
<< ppolyres >>
rect -50 -1000 50 1000
rect 68 -1000 168 1000
rect 186 -1000 286 1000
rect 304 -1000 404 1000
<< metal1 >>
rect -138 1126 492 1131
rect -138 1110 -103 1126
rect 457 1110 492 1126
rect -138 1105 492 1110
rect -138 1096 -112 1105
rect -138 -1096 -133 1096
rect -117 -1096 -112 1096
rect 466 1096 492 1105
rect -138 -1105 -112 -1096
rect 466 -1096 471 1096
rect 487 -1096 492 1096
rect 466 -1105 492 -1096
rect -138 -1110 492 -1105
rect -138 -1126 -103 -1110
rect 457 -1126 492 -1110
rect -138 -1131 492 -1126
<< properties >>
string gencell rppd
string library sg13g2_devstdin
string parameters w 1 l 20 nx 4 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class resistor endcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
