magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757454070
<< nwell >>
rect 19018 61711 19682 62359
rect 19018 59529 19682 59559
rect 17481 59451 19682 59529
rect 19018 58911 19682 59451
rect 19018 56729 19682 56759
rect 17481 56651 19682 56729
rect 19018 56111 19682 56651
rect 19018 53929 19682 53959
rect 17481 53851 19682 53929
rect 19018 53311 19682 53851
rect 19018 51129 19682 51159
rect 17481 51051 19682 51129
rect 19018 50511 19682 51051
rect 19018 48329 19682 48359
rect 17481 48251 19682 48329
rect 19018 47711 19682 48251
rect 19018 45529 19682 45559
rect 17481 45451 19682 45529
rect 19018 44911 19682 45451
rect 19018 42729 19682 42759
rect 17481 42651 19682 42729
rect 19018 42111 19682 42651
rect 19018 39929 19682 39959
rect 17481 39851 19682 39929
rect 19018 39311 19682 39851
rect 19018 37129 19682 37159
rect 17481 37051 19682 37129
rect 19018 36511 19682 37051
rect 19018 34329 19682 34359
rect 17481 34251 19682 34329
rect 19018 33711 19682 34251
rect 19018 31529 19682 31559
rect 17481 31451 19682 31529
rect 19018 30911 19682 31451
rect 19018 28729 19682 28759
rect 17481 28651 19682 28729
rect 19018 28111 19682 28651
rect 19018 25929 19682 25959
rect 17481 25851 19682 25929
rect 19018 25311 19682 25851
rect 19018 23129 19682 23159
rect 17481 23051 19682 23129
rect 19018 22511 19682 23051
rect 19018 20329 19682 20359
rect 17481 20251 19682 20329
rect 19018 19711 19682 20251
rect 17481 17451 19682 17529
<< metal1 >>
rect 16241 62963 18113 63063
rect 16241 62663 16341 62963
rect 18013 62663 18113 62963
rect 16241 62411 18113 62663
rect 26356 62963 27860 63063
rect -1354 61158 1738 62358
rect -1354 14839 -154 61158
rect 538 16731 1738 61158
rect 16241 62316 17324 62411
rect 16241 61929 16757 62316
rect 17163 61929 17324 62316
rect 20836 62312 26044 62426
rect 17432 62302 26044 62312
rect 17432 62236 17442 62302
rect 17508 62236 26044 62302
rect 17432 62226 26044 62236
rect 16241 61746 17324 61929
rect 17624 62109 20655 62129
rect 17624 61895 20244 62109
rect 16241 59825 16482 61746
rect 17624 61744 18894 61895
rect 20224 61778 20244 61895
rect 20635 61778 20655 62109
rect 19631 61739 20062 61759
rect 20224 61758 20655 61778
rect 19631 60252 19651 61739
rect 20042 60252 20062 61739
rect 19631 60232 20062 60252
rect 14699 59758 16401 59759
rect 14300 59749 16401 59758
rect 14300 59600 16251 59749
rect 16391 59600 16401 59749
rect 14300 59590 16401 59600
rect 14300 59589 15721 59590
rect 16467 59521 17324 59595
rect 16241 59516 17324 59521
rect 16241 59129 16757 59516
rect 17163 59129 17324 59516
rect 20836 59512 25572 59626
rect 17432 59502 25572 59512
rect 17432 59436 17442 59502
rect 17508 59436 25572 59502
rect 17432 59426 25572 59436
rect 16241 58946 17324 59129
rect 17624 59309 20655 59329
rect 17624 59095 20244 59309
rect 16241 57025 16482 58946
rect 17624 58944 18894 59095
rect 20224 58978 20244 59095
rect 20635 58978 20655 59309
rect 19631 58939 20062 58959
rect 20224 58958 20655 58978
rect 19631 57452 19651 58939
rect 20042 57452 20062 58939
rect 19631 57432 20062 57452
rect 14699 56958 16401 56959
rect 14300 56949 16401 56958
rect 14300 56800 16251 56949
rect 16391 56800 16401 56949
rect 14300 56790 16401 56800
rect 14300 56789 15721 56790
rect 16467 56721 17324 56795
rect 16241 56716 17324 56721
rect 16241 56329 16757 56716
rect 17163 56329 17324 56716
rect 20836 56712 25100 56826
rect 17432 56702 25100 56712
rect 17432 56636 17442 56702
rect 17508 56636 25100 56702
rect 17432 56626 25100 56636
rect 16241 56146 17324 56329
rect 17624 56509 20655 56529
rect 17624 56295 20244 56509
rect 16241 54225 16482 56146
rect 17624 56144 18894 56295
rect 20224 56178 20244 56295
rect 20635 56178 20655 56509
rect 19631 56139 20062 56159
rect 20224 56158 20655 56178
rect 19631 54652 19651 56139
rect 20042 54652 20062 56139
rect 19631 54632 20062 54652
rect 14699 54158 16401 54159
rect 14300 54149 16401 54158
rect 14300 54000 16251 54149
rect 16391 54000 16401 54149
rect 14300 53990 16401 54000
rect 14300 53989 15721 53990
rect 16467 53921 17324 53995
rect 16241 53916 17324 53921
rect 16241 53529 16757 53916
rect 17163 53529 17324 53916
rect 20836 53912 24628 54026
rect 17432 53902 24628 53912
rect 17432 53836 17442 53902
rect 17508 53836 24628 53902
rect 17432 53826 24628 53836
rect 16241 53346 17324 53529
rect 17624 53709 20655 53729
rect 17624 53495 20244 53709
rect 16241 51425 16482 53346
rect 17624 53344 18894 53495
rect 20224 53378 20244 53495
rect 20635 53378 20655 53709
rect 19631 53339 20062 53359
rect 20224 53358 20655 53378
rect 19631 51852 19651 53339
rect 20042 51852 20062 53339
rect 19631 51832 20062 51852
rect 14699 51358 16401 51359
rect 14300 51349 16401 51358
rect 14300 51200 16251 51349
rect 16391 51200 16401 51349
rect 14300 51190 16401 51200
rect 14300 51189 15721 51190
rect 16467 51121 17324 51195
rect 16241 51116 17324 51121
rect 16241 50729 16757 51116
rect 17163 50729 17324 51116
rect 20836 51112 24156 51226
rect 17432 51102 24156 51112
rect 17432 51036 17442 51102
rect 17508 51036 24156 51102
rect 17432 51026 24156 51036
rect 16241 50546 17324 50729
rect 17624 50909 20655 50929
rect 17624 50695 20244 50909
rect 16241 48625 16482 50546
rect 17624 50544 18894 50695
rect 20224 50578 20244 50695
rect 20635 50578 20655 50909
rect 19631 50539 20062 50559
rect 20224 50558 20655 50578
rect 19631 49052 19651 50539
rect 20042 49052 20062 50539
rect 19631 49032 20062 49052
rect 14699 48558 16401 48559
rect 14300 48549 16401 48558
rect 14300 48400 16251 48549
rect 16391 48400 16401 48549
rect 14300 48390 16401 48400
rect 14300 48389 15721 48390
rect 16467 48321 17324 48395
rect 16241 48316 17324 48321
rect 16241 47929 16757 48316
rect 17163 47929 17324 48316
rect 20836 48312 23684 48426
rect 17432 48302 23684 48312
rect 17432 48236 17442 48302
rect 17508 48236 23684 48302
rect 17432 48226 23684 48236
rect 16241 47746 17324 47929
rect 17624 48109 20655 48129
rect 17624 47895 20244 48109
rect 16241 45825 16482 47746
rect 17624 47744 18894 47895
rect 20224 47778 20244 47895
rect 20635 47778 20655 48109
rect 19631 47739 20062 47759
rect 20224 47758 20655 47778
rect 19631 46252 19651 47739
rect 20042 46252 20062 47739
rect 19631 46232 20062 46252
rect 14699 45758 16401 45759
rect 14300 45749 16401 45758
rect 14300 45600 16251 45749
rect 16391 45600 16401 45749
rect 14300 45590 16401 45600
rect 14300 45589 15721 45590
rect 16467 45521 17324 45595
rect 16241 45516 17324 45521
rect 16241 45129 16757 45516
rect 17163 45129 17324 45516
rect 20836 45512 23212 45626
rect 17432 45502 23212 45512
rect 17432 45436 17442 45502
rect 17508 45436 23212 45502
rect 17432 45426 23212 45436
rect 16241 44946 17324 45129
rect 17624 45309 20655 45329
rect 17624 45095 20244 45309
rect 16241 43025 16482 44946
rect 17624 44944 18894 45095
rect 20224 44978 20244 45095
rect 20635 44978 20655 45309
rect 19631 44939 20062 44959
rect 20224 44958 20655 44978
rect 19631 43452 19651 44939
rect 20042 43452 20062 44939
rect 19631 43432 20062 43452
rect 14699 42958 16401 42959
rect 14300 42949 16401 42958
rect 14300 42800 16251 42949
rect 16391 42800 16401 42949
rect 14300 42790 16401 42800
rect 14300 42789 15721 42790
rect 16467 42721 17324 42795
rect 16241 42716 17324 42721
rect 16241 42329 16757 42716
rect 17163 42329 17324 42716
rect 20836 42712 22740 42826
rect 17432 42702 22740 42712
rect 17432 42636 17442 42702
rect 17508 42636 22740 42702
rect 17432 42626 22740 42636
rect 16241 42146 17324 42329
rect 17624 42509 20655 42529
rect 17624 42295 20244 42509
rect 16241 40225 16482 42146
rect 17624 42144 18894 42295
rect 20224 42178 20244 42295
rect 20635 42178 20655 42509
rect 19631 42139 20062 42159
rect 20224 42158 20655 42178
rect 19631 40652 19651 42139
rect 20042 40652 20062 42139
rect 19631 40632 20062 40652
rect 14699 40158 16401 40159
rect 14300 40149 16401 40158
rect 14300 40000 16251 40149
rect 16391 40000 16401 40149
rect 14300 39990 16401 40000
rect 14300 39989 15721 39990
rect 16467 39921 17324 39995
rect 16241 39916 17324 39921
rect 16241 39529 16757 39916
rect 17163 39529 17324 39916
rect 20836 39912 22268 40026
rect 17432 39902 22268 39912
rect 17432 39836 17442 39902
rect 17508 39836 22268 39902
rect 17432 39826 22268 39836
rect 16241 39346 17324 39529
rect 17624 39709 20655 39729
rect 17624 39495 20244 39709
rect 16241 37425 16482 39346
rect 17624 39344 18894 39495
rect 20224 39378 20244 39495
rect 20635 39378 20655 39709
rect 19631 39339 20062 39359
rect 20224 39358 20655 39378
rect 19631 37852 19651 39339
rect 20042 37852 20062 39339
rect 19631 37832 20062 37852
rect 14699 37358 16401 37359
rect 14300 37349 16401 37358
rect 14300 37200 16251 37349
rect 16391 37200 16401 37349
rect 14300 37190 16401 37200
rect 14300 37189 15721 37190
rect 16467 37121 17324 37195
rect 16241 37116 17324 37121
rect 16241 36729 16757 37116
rect 17163 36729 17324 37116
rect 20836 37112 21796 37226
rect 17432 37102 21796 37112
rect 17432 37036 17442 37102
rect 17508 37036 21796 37102
rect 17432 37026 21796 37036
rect 16241 36546 17324 36729
rect 17624 36909 20655 36929
rect 17624 36695 20244 36909
rect 16241 34625 16482 36546
rect 17624 36544 18894 36695
rect 20224 36578 20244 36695
rect 20635 36578 20655 36909
rect 19631 36539 20062 36559
rect 20224 36558 20655 36578
rect 19631 35052 19651 36539
rect 20042 35052 20062 36539
rect 19631 35032 20062 35052
rect 14699 34558 16401 34559
rect 14300 34549 16401 34558
rect 14300 34400 16251 34549
rect 16391 34400 16401 34549
rect 14300 34390 16401 34400
rect 14300 34389 15721 34390
rect 16467 34321 17324 34395
rect 16241 34316 17324 34321
rect 16241 33929 16757 34316
rect 17163 33929 17324 34316
rect 20836 34312 21324 34426
rect 17432 34302 21324 34312
rect 17432 34236 17442 34302
rect 17508 34236 21324 34302
rect 17432 34226 21324 34236
rect 16241 33746 17324 33929
rect 17624 34109 20655 34129
rect 17624 33895 20244 34109
rect 16241 31825 16482 33746
rect 17624 33744 18894 33895
rect 20224 33778 20244 33895
rect 20635 33778 20655 34109
rect 19631 33739 20062 33759
rect 20224 33758 20655 33778
rect 19631 32252 19651 33739
rect 20042 32252 20062 33739
rect 21124 33508 21324 34226
rect 21124 33328 21134 33508
rect 21314 33328 21324 33508
rect 21124 33318 21324 33328
rect 19631 32232 20062 32252
rect 21124 33008 21324 33018
rect 21124 32828 21134 33008
rect 21314 32828 21324 33008
rect 14699 31758 16401 31759
rect 14300 31749 16401 31758
rect 14300 31600 16251 31749
rect 16391 31600 16401 31749
rect 21124 31626 21324 32828
rect 21596 32508 21796 37026
rect 21596 32328 21606 32508
rect 21786 32328 21796 32508
rect 21596 32318 21796 32328
rect 14300 31590 16401 31600
rect 14300 31589 15721 31590
rect 16467 31521 17324 31595
rect 16241 31516 17324 31521
rect 16241 31129 16757 31516
rect 17163 31129 17324 31516
rect 20836 31512 21324 31626
rect 17432 31502 21324 31512
rect 17432 31436 17442 31502
rect 17508 31436 21324 31502
rect 17432 31426 21324 31436
rect 21596 32008 21796 32018
rect 21596 31828 21606 32008
rect 21786 31828 21796 32008
rect 16241 30946 17324 31129
rect 17624 31309 20655 31329
rect 17624 31095 20244 31309
rect 16241 29025 16482 30946
rect 17624 30944 18894 31095
rect 20224 30978 20244 31095
rect 20635 30978 20655 31309
rect 19631 30939 20062 30959
rect 20224 30958 20655 30978
rect 19631 29452 19651 30939
rect 20042 29452 20062 30939
rect 19631 29432 20062 29452
rect 14699 28958 16401 28959
rect 14300 28949 16401 28958
rect 14300 28800 16251 28949
rect 16391 28800 16401 28949
rect 21596 28826 21796 31828
rect 22068 31508 22268 39826
rect 22068 31328 22078 31508
rect 22258 31328 22268 31508
rect 22068 31318 22268 31328
rect 14300 28790 16401 28800
rect 14300 28789 15721 28790
rect 16467 28721 17324 28795
rect 16241 28716 17324 28721
rect 16241 28329 16757 28716
rect 17163 28329 17324 28716
rect 20836 28712 21796 28826
rect 17432 28702 21796 28712
rect 17432 28636 17442 28702
rect 17508 28636 21796 28702
rect 17432 28626 21796 28636
rect 22068 31008 22268 31018
rect 22068 30828 22078 31008
rect 22258 30828 22268 31008
rect 16241 28146 17324 28329
rect 17624 28509 20655 28529
rect 17624 28295 20244 28509
rect 16241 26225 16482 28146
rect 17624 28144 18894 28295
rect 20224 28178 20244 28295
rect 20635 28178 20655 28509
rect 19631 28139 20062 28159
rect 20224 28158 20655 28178
rect 19631 26652 19651 28139
rect 20042 26652 20062 28139
rect 19631 26632 20062 26652
rect 14699 26158 16401 26159
rect 14300 26149 16401 26158
rect 14300 26000 16251 26149
rect 16391 26000 16401 26149
rect 22068 26026 22268 30828
rect 22540 30508 22740 42626
rect 22540 30328 22550 30508
rect 22730 30328 22740 30508
rect 22540 30318 22740 30328
rect 14300 25990 16401 26000
rect 14300 25989 15721 25990
rect 16467 25921 17324 25995
rect 16241 25916 17324 25921
rect 16241 25529 16757 25916
rect 17163 25529 17324 25916
rect 20836 25912 22268 26026
rect 17432 25902 22268 25912
rect 17432 25836 17442 25902
rect 17508 25836 22268 25902
rect 17432 25826 22268 25836
rect 22540 30008 22740 30018
rect 22540 29828 22550 30008
rect 22730 29828 22740 30008
rect 16241 25346 17324 25529
rect 17624 25709 20655 25729
rect 17624 25495 20244 25709
rect 16241 23425 16482 25346
rect 17624 25344 18894 25495
rect 20224 25378 20244 25495
rect 20635 25378 20655 25709
rect 19631 25339 20062 25359
rect 20224 25358 20655 25378
rect 19631 23852 19651 25339
rect 20042 23852 20062 25339
rect 19631 23832 20062 23852
rect 14699 23358 16401 23359
rect 14300 23349 16401 23358
rect 14300 23200 16251 23349
rect 16391 23200 16401 23349
rect 22540 23226 22740 29828
rect 23012 29508 23212 45426
rect 23012 29328 23022 29508
rect 23202 29328 23212 29508
rect 23012 29318 23212 29328
rect 14300 23190 16401 23200
rect 14300 23189 15721 23190
rect 16467 23121 17324 23195
rect 16241 23116 17324 23121
rect 16241 22729 16757 23116
rect 17163 22729 17324 23116
rect 20836 23112 22740 23226
rect 17432 23102 22740 23112
rect 17432 23036 17442 23102
rect 17508 23036 22740 23102
rect 17432 23026 22740 23036
rect 23012 29008 23212 29018
rect 23012 28828 23022 29008
rect 23202 28828 23212 29008
rect 16241 22546 17324 22729
rect 17624 22909 20655 22929
rect 17624 22695 20244 22909
rect 16241 20625 16482 22546
rect 17624 22544 18894 22695
rect 20224 22578 20244 22695
rect 20635 22578 20655 22909
rect 19631 22539 20062 22559
rect 20224 22558 20655 22578
rect 19631 21052 19651 22539
rect 20042 21052 20062 22539
rect 19631 21032 20062 21052
rect 14699 20558 16401 20559
rect 14300 20549 16401 20558
rect 14300 20400 16251 20549
rect 16391 20400 16401 20549
rect 23012 20426 23212 28828
rect 23484 28508 23684 48226
rect 23484 28328 23494 28508
rect 23674 28328 23684 28508
rect 23484 28318 23684 28328
rect 23956 28008 24156 51026
rect 23956 27828 23966 28008
rect 24146 27828 24156 28008
rect 23956 27818 24156 27828
rect 24428 27508 24628 53826
rect 24428 27328 24438 27508
rect 24618 27328 24628 27508
rect 24428 27318 24628 27328
rect 24900 27008 25100 56626
rect 24900 26828 24910 27008
rect 25090 26828 25100 27008
rect 24900 26818 25100 26828
rect 25372 26508 25572 59426
rect 25372 26328 25382 26508
rect 25562 26328 25572 26508
rect 25372 26318 25572 26328
rect 25844 26008 26044 62226
rect 26356 62263 26456 62963
rect 27760 62263 27860 62963
rect 26356 61969 27860 62263
rect 26356 34278 26556 61969
rect 27232 61960 27860 61969
rect 28404 62963 58632 63063
rect 28404 62263 28504 62963
rect 32937 62263 54100 62963
rect 58532 62263 58632 62963
rect 28404 62063 58632 62263
rect 27232 34278 27432 61960
rect 28404 61958 58110 62063
rect 41584 53264 58110 53536
rect 41416 41612 41779 42497
rect 58432 42279 58632 62063
rect 59036 62963 63078 63063
rect 59036 62263 59136 62963
rect 62978 62263 63078 62963
rect 59036 61915 63078 62263
rect 64909 62963 68168 63063
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 61926 68168 62363
rect 64765 61921 68168 61926
rect 71457 62970 75284 63070
rect 71457 62283 71557 62970
rect 75184 62283 75284 62970
rect 71457 62183 75284 62283
rect 59036 52413 59313 61915
rect 64765 60835 64916 61921
rect 71457 61790 72778 62183
rect 61697 59704 65212 60544
rect 61697 50746 62497 59704
rect 70717 56705 70907 56715
rect 70717 56505 70727 56705
rect 70897 56505 70907 56705
rect 70717 51441 70907 56505
rect 71137 56705 71327 56715
rect 71137 56505 71147 56705
rect 71317 56505 71327 56705
rect 71137 52141 71327 56505
rect 71457 55812 72097 61790
rect 76075 61705 76949 61805
rect 76075 52782 76199 61705
rect 76849 52782 76949 61705
rect 76075 52682 76949 52782
rect 71137 52131 81037 52141
rect 71137 51751 76319 52131
rect 76699 51751 81037 52131
rect 71137 51741 81037 51751
rect 70717 51041 81037 51441
rect 58196 42079 58632 42279
rect 41416 41602 71917 41612
rect 41416 41259 71546 41602
rect 71907 41259 71917 41602
rect 41416 41249 71917 41259
rect 41399 40607 59348 40617
rect 41399 40246 58977 40607
rect 59338 40246 59348 40607
rect 41399 40236 59348 40246
rect 62933 40509 63123 40519
rect 62933 40329 62943 40509
rect 63113 40329 63123 40509
rect 41399 38167 41780 40236
rect 60413 36515 60603 36525
rect 60413 36335 60423 36515
rect 60593 36335 60603 36515
rect 26356 34078 27432 34278
rect 41402 33270 41783 34584
rect 25844 25828 25854 26008
rect 26034 25828 26044 26008
rect 25844 25818 26044 25828
rect 27820 33068 41783 33270
rect 42570 34359 42951 34369
rect 42570 34068 42580 34359
rect 42941 34068 42951 34359
rect 14300 20390 16401 20400
rect 14300 20389 15721 20390
rect 16467 20321 17324 20395
rect 16241 20316 17324 20321
rect 16241 19929 16757 20316
rect 17163 19929 17324 20316
rect 20836 20312 23212 20426
rect 17432 20302 23212 20312
rect 17432 20236 17442 20302
rect 17508 20236 23212 20302
rect 17432 20226 23212 20236
rect 16241 19746 17324 19929
rect 17624 20109 20655 20129
rect 17624 19895 20244 20109
rect 16241 17825 16482 19746
rect 17624 19744 18894 19895
rect 20224 19778 20244 19895
rect 20635 19778 20655 20109
rect 19631 19739 20062 19759
rect 20224 19758 20655 19778
rect 19631 18252 19651 19739
rect 20042 18252 20062 19739
rect 19631 18232 20062 18252
rect 14699 17758 16401 17759
rect 14300 17749 16401 17758
rect 14300 17600 16251 17749
rect 16391 17600 16401 17749
rect 14300 17590 16401 17600
rect 14300 17589 15721 17590
rect 16467 17518 17324 17595
rect 16241 17451 17324 17518
rect 538 15531 12911 16731
rect -1354 13639 10705 14839
rect 9367 1041 10705 13639
rect 11397 1041 12911 15531
rect 27820 14620 28202 33068
rect 42570 32269 42951 34068
rect 27820 14290 27830 14620
rect 28192 14290 28202 14620
rect 27820 14280 28202 14290
rect 28847 32067 42951 32269
rect 28847 13602 29228 32067
rect 60413 24612 60603 36335
rect 60413 24431 60423 24612
rect 60593 24431 60603 24612
rect 60413 24421 60603 24431
rect 60833 36015 61023 36025
rect 60833 35835 60843 36015
rect 61013 35835 61023 36015
rect 60833 24612 61023 35835
rect 60833 24431 60843 24612
rect 61013 24431 61023 24612
rect 60833 24421 61023 24431
rect 61253 35515 61443 35525
rect 61253 35335 61263 35515
rect 61433 35335 61443 35515
rect 61253 24612 61443 35335
rect 61253 24431 61263 24612
rect 61433 24431 61443 24612
rect 61253 24421 61443 24431
rect 61673 35015 61863 35025
rect 61673 34835 61683 35015
rect 61853 34835 61863 35015
rect 61673 24612 61863 34835
rect 61673 24431 61683 24612
rect 61853 24431 61863 24612
rect 61673 24421 61863 24431
rect 62093 34515 62283 34525
rect 62093 34335 62103 34515
rect 62273 34335 62283 34515
rect 62093 24612 62283 34335
rect 62093 24431 62103 24612
rect 62273 24431 62283 24612
rect 62093 24421 62283 24431
rect 62513 34015 62703 34025
rect 62513 33835 62523 34015
rect 62693 33835 62703 34015
rect 62513 24612 62703 33835
rect 62513 24431 62523 24612
rect 62693 24431 62703 24612
rect 62513 24421 62703 24431
rect 62933 24612 63123 40329
rect 67969 40509 68159 40519
rect 67969 40329 67979 40509
rect 68149 40329 68159 40509
rect 62933 24431 62943 24612
rect 63113 24431 63123 24612
rect 62933 24421 63123 24431
rect 63353 40009 63543 40019
rect 63353 39829 63363 40009
rect 63533 39829 63543 40009
rect 63353 24612 63543 39829
rect 65873 39509 66063 39519
rect 65873 39329 65883 39509
rect 66053 39329 66063 39509
rect 65453 39009 65643 39019
rect 65453 38829 65463 39009
rect 65633 38829 65643 39009
rect 65033 38509 65223 38519
rect 65033 38329 65043 38509
rect 65213 38329 65223 38509
rect 64613 38009 64803 38019
rect 64613 37829 64623 38009
rect 64793 37829 64803 38009
rect 64193 37509 64383 37519
rect 64193 37329 64203 37509
rect 64373 37329 64383 37509
rect 63353 24431 63363 24612
rect 63533 24431 63543 24612
rect 63353 24421 63543 24431
rect 63773 37009 63963 37019
rect 63773 36829 63783 37009
rect 63953 36829 63963 37009
rect 63773 24612 63963 36829
rect 63773 24431 63783 24612
rect 63953 24431 63963 24612
rect 63773 24421 63963 24431
rect 64193 24612 64383 37329
rect 64193 24431 64203 24612
rect 64373 24431 64383 24612
rect 64193 24421 64383 24431
rect 64613 24612 64803 37829
rect 64613 24431 64623 24612
rect 64793 24431 64803 24612
rect 64613 24421 64803 24431
rect 65033 24612 65223 38329
rect 65033 24431 65043 24612
rect 65213 24431 65223 24612
rect 65033 24421 65223 24431
rect 65453 24612 65643 38829
rect 65453 24431 65463 24612
rect 65633 24431 65643 24612
rect 65453 24421 65643 24431
rect 65873 24612 66063 39329
rect 67133 33508 67323 33518
rect 67133 33328 67143 33508
rect 67313 33328 67323 33508
rect 66713 32508 66903 32518
rect 66713 32328 66723 32508
rect 66893 32328 66903 32508
rect 65873 24431 65883 24612
rect 66053 24431 66063 24612
rect 65873 24421 66063 24431
rect 66293 31508 66483 31518
rect 66293 31328 66303 31508
rect 66473 31328 66483 31508
rect 66293 24612 66483 31328
rect 66293 24431 66303 24612
rect 66473 24431 66483 24612
rect 66293 24421 66483 24431
rect 66713 24612 66903 32328
rect 66713 24431 66723 24612
rect 66893 24431 66903 24612
rect 66713 24421 66903 24431
rect 67133 24612 67323 33328
rect 67133 24431 67143 24612
rect 67313 24431 67323 24612
rect 67133 24421 67323 24431
rect 67553 33008 67743 33018
rect 67553 32828 67563 33008
rect 67733 32828 67743 33008
rect 67553 24612 67743 32828
rect 67969 32777 68159 40329
rect 68389 40009 68579 40019
rect 68389 39829 68399 40009
rect 68569 39829 68579 40009
rect 68389 33277 68579 39829
rect 68809 39509 68999 39519
rect 68809 39329 68819 39509
rect 68989 39329 68999 39509
rect 68809 33777 68999 39329
rect 69229 39009 69419 39019
rect 69229 38829 69239 39009
rect 69409 38829 69419 39009
rect 69229 34277 69419 38829
rect 69649 38509 69839 38519
rect 69649 38329 69659 38509
rect 69829 38329 69839 38509
rect 69649 34777 69839 38329
rect 70069 38009 70259 38019
rect 70069 37829 70079 38009
rect 70249 37829 70259 38009
rect 70069 35277 70259 37829
rect 70489 37509 70679 37519
rect 70489 37329 70499 37509
rect 70669 37329 70679 37509
rect 70489 35771 70679 37329
rect 70909 37009 71099 37019
rect 70909 36829 70919 37009
rect 71089 36829 71099 37009
rect 70909 36271 71099 36829
rect 70909 36071 76143 36271
rect 70489 35571 75723 35771
rect 70069 35077 75303 35277
rect 69649 34577 74883 34777
rect 69229 34077 74463 34277
rect 68809 33577 74043 33777
rect 68389 33077 73623 33277
rect 67969 32577 73203 32777
rect 67553 24431 67563 24612
rect 67733 24431 67743 24612
rect 67553 24421 67743 24431
rect 67973 32008 68163 32018
rect 67973 31828 67983 32008
rect 68153 31828 68163 32008
rect 67973 24612 68163 31828
rect 67973 24431 67983 24612
rect 68153 24431 68163 24612
rect 67973 24421 68163 24431
rect 68393 31008 68583 31018
rect 68393 30828 68403 31008
rect 68573 30828 68583 31008
rect 68393 24612 68583 30828
rect 72593 30508 72783 30518
rect 72593 30328 72603 30508
rect 72773 30328 72783 30508
rect 68393 24431 68403 24612
rect 68573 24431 68583 24612
rect 68393 24421 68583 24431
rect 68813 30008 69003 30018
rect 68813 29828 68823 30008
rect 68993 29828 69003 30008
rect 68813 24612 69003 29828
rect 72173 29508 72363 29518
rect 72173 29328 72183 29508
rect 72353 29328 72363 29508
rect 68813 24431 68823 24612
rect 68993 24431 69003 24612
rect 68813 24421 69003 24431
rect 69233 29008 69423 29018
rect 69233 28828 69243 29008
rect 69413 28828 69423 29008
rect 69233 24612 69423 28828
rect 71753 28508 71943 28518
rect 71753 28328 71763 28508
rect 71933 28328 71943 28508
rect 71333 28008 71523 28018
rect 71333 27828 71343 28008
rect 71513 27828 71523 28008
rect 70913 27508 71103 27518
rect 70913 27328 70923 27508
rect 71093 27328 71103 27508
rect 70493 27008 70683 27018
rect 70493 26828 70503 27008
rect 70673 26828 70683 27008
rect 70073 26508 70263 26518
rect 70073 26328 70083 26508
rect 70253 26328 70263 26508
rect 69233 24431 69243 24612
rect 69413 24431 69423 24612
rect 69233 24421 69423 24431
rect 69653 26008 69843 26018
rect 69653 25828 69663 26008
rect 69833 25828 69843 26008
rect 69653 24612 69843 25828
rect 69653 24431 69663 24612
rect 69833 24431 69843 24612
rect 69653 24421 69843 24431
rect 70073 24612 70263 26328
rect 70073 24431 70083 24612
rect 70253 24431 70263 24612
rect 70073 24421 70263 24431
rect 70493 24612 70683 26828
rect 70493 24431 70503 24612
rect 70673 24431 70683 24612
rect 70493 24421 70683 24431
rect 70913 24612 71103 27328
rect 70913 24431 70923 24612
rect 71093 24431 71103 24612
rect 70913 24421 71103 24431
rect 71333 24612 71523 27828
rect 71333 24431 71343 24612
rect 71513 24431 71523 24612
rect 71333 24421 71523 24431
rect 71753 24612 71943 28328
rect 71753 24431 71763 24612
rect 71933 24431 71943 24612
rect 71753 24421 71943 24431
rect 72173 24612 72363 29328
rect 72173 24431 72183 24612
rect 72353 24431 72363 24612
rect 72173 24421 72363 24431
rect 72593 24612 72783 30328
rect 72593 24431 72603 24612
rect 72773 24431 72783 24612
rect 72593 24421 72783 24431
rect 73013 24612 73203 32577
rect 73013 24431 73023 24612
rect 73193 24431 73203 24612
rect 73013 24421 73203 24431
rect 73433 24612 73623 33077
rect 73433 24431 73443 24612
rect 73613 24431 73623 24612
rect 73433 24421 73623 24431
rect 73853 24612 74043 33577
rect 73853 24431 73863 24612
rect 74033 24431 74043 24612
rect 73853 24421 74043 24431
rect 74273 24612 74463 34077
rect 74273 24431 74283 24612
rect 74453 24431 74463 24612
rect 74273 24421 74463 24431
rect 74693 24612 74883 34577
rect 74693 24431 74703 24612
rect 74873 24431 74883 24612
rect 74693 24421 74883 24431
rect 75113 24612 75303 35077
rect 75113 24431 75123 24612
rect 75293 24431 75303 24612
rect 75113 24421 75303 24431
rect 75533 24612 75723 35571
rect 75533 24431 75543 24612
rect 75713 24431 75723 24612
rect 75533 24421 75723 24431
rect 75953 24612 76143 36071
rect 75953 24431 75963 24612
rect 76133 24431 76143 24612
rect 75953 24421 76143 24431
rect 28847 13272 28857 13602
rect 29218 13272 29228 13602
rect 28847 13262 29228 13272
rect 28416 12447 30903 12658
rect 47878 12558 48289 12658
rect -1884 524 -787 725
rect 9367 585 12911 1041
rect 13048 7276 14456 9031
rect -1884 -5827 -1484 524
rect -912 -602 9370 -502
rect -912 -1416 -812 -602
rect 9270 -1416 9370 -602
rect -912 -1516 9370 -1416
rect 10344 -5827 11144 585
rect 13048 -56 14114 7276
rect 28416 4302 30569 12447
rect 28416 2423 30903 4302
rect 22075 1569 22746 1579
rect 22075 1113 22085 1569
rect 22736 1113 22746 1569
rect 22075 1103 22746 1113
rect 30354 777 30899 2423
rect 13048 -657 13148 -56
rect 14014 -657 14114 -56
rect 13048 -757 14114 -657
rect 14438 -57 18572 612
rect 14438 -657 14538 -57
rect 18472 -657 18572 -57
rect 14438 -757 18572 -657
rect 20819 298 21171 308
rect 20819 -34 20829 298
rect 21161 -34 21171 298
rect 20819 -959 21171 -34
rect 22953 -369 28430 636
rect 30354 622 33209 777
rect 48189 670 48289 12558
rect 30354 -166 30454 622
rect 33109 -166 33209 622
rect 47878 570 48289 670
rect 44588 470 48289 570
rect 33443 332 37478 342
rect 33443 -10 33453 332
rect 33786 -10 37135 332
rect 37468 -10 37478 332
rect 33443 -20 37478 -10
rect 30354 -266 33209 -166
rect 44588 -261 44688 470
rect 48189 -261 48289 470
rect 44588 -361 48289 -261
rect 22953 -669 23053 -369
rect 28330 -669 28430 -369
rect 22953 -769 28430 -669
rect 20819 -1291 20829 -959
rect 21161 -1291 21171 -959
rect 20819 -1301 21171 -1291
<< via1 >>
rect 16341 62663 18013 62963
rect -154 15531 538 61158
rect 16757 61929 17163 62316
rect 17442 62236 17508 62302
rect 20244 61778 20635 62109
rect 19651 60252 20042 61739
rect 16251 59600 16391 59749
rect 16757 59129 17163 59516
rect 17442 59436 17508 59502
rect 20244 58978 20635 59309
rect 19651 57452 20042 58939
rect 16251 56800 16391 56949
rect 16757 56329 17163 56716
rect 17442 56636 17508 56702
rect 20244 56178 20635 56509
rect 19651 54652 20042 56139
rect 16251 54000 16391 54149
rect 16757 53529 17163 53916
rect 17442 53836 17508 53902
rect 20244 53378 20635 53709
rect 19651 51852 20042 53339
rect 16251 51200 16391 51349
rect 16757 50729 17163 51116
rect 17442 51036 17508 51102
rect 20244 50578 20635 50909
rect 19651 49052 20042 50539
rect 16251 48400 16391 48549
rect 16757 47929 17163 48316
rect 17442 48236 17508 48302
rect 20244 47778 20635 48109
rect 19651 46252 20042 47739
rect 16251 45600 16391 45749
rect 16757 45129 17163 45516
rect 17442 45436 17508 45502
rect 20244 44978 20635 45309
rect 19651 43452 20042 44939
rect 16251 42800 16391 42949
rect 16757 42329 17163 42716
rect 17442 42636 17508 42702
rect 20244 42178 20635 42509
rect 19651 40652 20042 42139
rect 16251 40000 16391 40149
rect 16757 39529 17163 39916
rect 17442 39836 17508 39902
rect 20244 39378 20635 39709
rect 19651 37852 20042 39339
rect 16251 37200 16391 37349
rect 16757 36729 17163 37116
rect 17442 37036 17508 37102
rect 20244 36578 20635 36909
rect 19651 35052 20042 36539
rect 16251 34400 16391 34549
rect 16757 33929 17163 34316
rect 17442 34236 17508 34302
rect 20244 33778 20635 34109
rect 19651 32252 20042 33739
rect 21134 33328 21314 33508
rect 21134 32828 21314 33008
rect 16251 31600 16391 31749
rect 21606 32328 21786 32508
rect 16757 31129 17163 31516
rect 17442 31436 17508 31502
rect 21606 31828 21786 32008
rect 20244 30978 20635 31309
rect 19651 29452 20042 30939
rect 16251 28800 16391 28949
rect 22078 31328 22258 31508
rect 16757 28329 17163 28716
rect 17442 28636 17508 28702
rect 22078 30828 22258 31008
rect 20244 28178 20635 28509
rect 19651 26652 20042 28139
rect 16251 26000 16391 26149
rect 22550 30328 22730 30508
rect 16757 25529 17163 25916
rect 17442 25836 17508 25902
rect 22550 29828 22730 30008
rect 20244 25378 20635 25709
rect 19651 23852 20042 25339
rect 16251 23200 16391 23349
rect 23022 29328 23202 29508
rect 16757 22729 17163 23116
rect 17442 23036 17508 23102
rect 23022 28828 23202 29008
rect 20244 22578 20635 22909
rect 19651 21052 20042 22539
rect 16251 20400 16391 20549
rect 23494 28328 23674 28508
rect 23966 27828 24146 28008
rect 24438 27328 24618 27508
rect 24910 26828 25090 27008
rect 25382 26328 25562 26508
rect 26456 62263 27760 62963
rect 26556 34278 27232 61969
rect 28504 62263 32937 62963
rect 54100 62263 58532 62963
rect 58110 42279 58432 62063
rect 59136 62263 62978 62963
rect 65009 62363 68068 62963
rect 71557 62283 75184 62970
rect 70727 56505 70897 56705
rect 71147 56505 71317 56705
rect 76199 52782 76849 61705
rect 76319 51751 76699 52131
rect 71546 41259 71907 41602
rect 58977 40246 59338 40607
rect 62943 40329 63113 40509
rect 60423 36335 60593 36515
rect 25854 25828 26034 26008
rect 42580 34068 42941 34359
rect 16757 19929 17163 20316
rect 17442 20236 17508 20302
rect 20244 19778 20635 20109
rect 19651 18252 20042 19739
rect 16251 17600 16391 17749
rect -154 14839 11397 15531
rect 10705 1041 11397 14839
rect 27830 14290 28192 14620
rect 60423 24431 60593 24612
rect 60843 35835 61013 36015
rect 60843 24431 61013 24612
rect 61263 35335 61433 35515
rect 61263 24431 61433 24612
rect 61683 34835 61853 35015
rect 61683 24431 61853 24612
rect 62103 34335 62273 34515
rect 62103 24431 62273 24612
rect 62523 33835 62693 34015
rect 62523 24431 62693 24612
rect 67979 40329 68149 40509
rect 62943 24431 63113 24612
rect 63363 39829 63533 40009
rect 65883 39329 66053 39509
rect 65463 38829 65633 39009
rect 65043 38329 65213 38509
rect 64623 37829 64793 38009
rect 64203 37329 64373 37509
rect 63363 24431 63533 24612
rect 63783 36829 63953 37009
rect 63783 24431 63953 24612
rect 64203 24431 64373 24612
rect 64623 24431 64793 24612
rect 65043 24431 65213 24612
rect 65463 24431 65633 24612
rect 67143 33328 67313 33508
rect 66723 32328 66893 32508
rect 65883 24431 66053 24612
rect 66303 31328 66473 31508
rect 66303 24431 66473 24612
rect 66723 24431 66893 24612
rect 67143 24431 67313 24612
rect 67563 32828 67733 33008
rect 68399 39829 68569 40009
rect 68819 39329 68989 39509
rect 69239 38829 69409 39009
rect 69659 38329 69829 38509
rect 70079 37829 70249 38009
rect 70499 37329 70669 37509
rect 70919 36829 71089 37009
rect 67563 24431 67733 24612
rect 67983 31828 68153 32008
rect 67983 24431 68153 24612
rect 68403 30828 68573 31008
rect 72603 30328 72773 30508
rect 68403 24431 68573 24612
rect 68823 29828 68993 30008
rect 72183 29328 72353 29508
rect 68823 24431 68993 24612
rect 69243 28828 69413 29008
rect 71763 28328 71933 28508
rect 71343 27828 71513 28008
rect 70923 27328 71093 27508
rect 70503 26828 70673 27008
rect 70083 26328 70253 26508
rect 69243 24431 69413 24612
rect 69663 25828 69833 26008
rect 69663 24431 69833 24612
rect 70083 24431 70253 24612
rect 70503 24431 70673 24612
rect 70923 24431 71093 24612
rect 71343 24431 71513 24612
rect 71763 24431 71933 24612
rect 72183 24431 72353 24612
rect 72603 24431 72773 24612
rect 73023 24431 73193 24612
rect 73443 24431 73613 24612
rect 73863 24431 74033 24612
rect 74283 24431 74453 24612
rect 74703 24431 74873 24612
rect 75123 24431 75293 24612
rect 75543 24431 75713 24612
rect 75963 24431 76133 24612
rect 28857 13272 29218 13602
rect -812 -1416 9270 -602
rect 30569 4302 30920 12447
rect 22085 1113 22736 1569
rect 39602 1281 42582 1536
rect 13148 -657 14014 -56
rect 14538 -657 18472 -57
rect 20829 -34 21161 298
rect 47858 670 48189 12558
rect 30454 -166 33109 622
rect 33453 -10 33786 332
rect 37135 -10 37468 332
rect 44688 -261 48189 470
rect 23053 -669 28330 -369
rect 20829 -1291 21161 -959
<< metal2 >>
rect 2657 62966 15745 63066
rect 2657 62466 2757 62966
rect 15645 62466 15745 62966
rect 16241 62963 18113 63063
rect 16241 62663 16341 62963
rect 18013 62663 18113 62963
rect 16241 62563 18113 62663
rect 18444 62963 20062 63063
rect 2657 62358 15745 62466
rect 18444 62463 18544 62963
rect 19962 62463 20062 62963
rect 18444 62364 20062 62463
rect -1354 61158 1738 62358
rect 2657 62003 16178 62358
rect 2657 61956 15027 62003
rect -1354 14839 -154 61158
rect 538 16731 1738 61158
rect 14226 59558 15027 61956
rect 2657 59156 15027 59558
rect 14226 56758 15027 59156
rect 2657 56356 15027 56758
rect 14226 53958 15027 56356
rect 2657 53556 15027 53958
rect 14226 51158 15027 53556
rect 2657 50756 15027 51158
rect 14226 48358 15027 50756
rect 2657 47956 15027 48358
rect 14226 45558 15027 47956
rect 2657 45156 15027 45558
rect 14226 42758 15027 45156
rect 2657 42356 15027 42758
rect 14226 39958 15027 42356
rect 2657 39556 15027 39958
rect 14226 37158 15027 39556
rect 2657 36756 15027 37158
rect 14226 34358 15027 36756
rect 2657 33956 15027 34358
rect 14226 31558 15027 33956
rect 2657 31156 15027 31558
rect 14226 28758 15027 31156
rect 2657 28356 15027 28758
rect 14226 25958 15027 28356
rect 2657 25556 15027 25958
rect 14226 23158 15027 25556
rect 2657 22756 15027 23158
rect 14226 20358 15027 22756
rect 2657 19956 15027 20358
rect 14226 17576 15027 19956
rect 15499 17576 16178 62003
rect 16747 62316 17173 62326
rect 16747 61929 16757 62316
rect 17163 61929 17173 62316
rect 16747 61919 17173 61929
rect 17432 62302 17518 62312
rect 17432 62236 17442 62302
rect 17508 62236 17518 62302
rect 17432 61712 17518 62236
rect 19631 61739 20062 62364
rect 19631 60252 19651 61739
rect 20042 60252 20062 61739
rect 16241 59749 17523 59759
rect 16241 59600 16251 59749
rect 16391 59600 17523 59749
rect 16241 59590 17523 59600
rect 16747 59516 17173 59526
rect 16747 59129 16757 59516
rect 17163 59129 17173 59516
rect 16747 59119 17173 59129
rect 17432 59502 17518 59512
rect 17432 59436 17442 59502
rect 17508 59436 17518 59502
rect 17432 58912 17518 59436
rect 19631 58939 20062 60252
rect 19631 57452 19651 58939
rect 20042 57452 20062 58939
rect 16241 56949 17523 56959
rect 16241 56800 16251 56949
rect 16391 56800 17523 56949
rect 16241 56790 17523 56800
rect 16747 56716 17173 56726
rect 16747 56329 16757 56716
rect 17163 56329 17173 56716
rect 16747 56319 17173 56329
rect 17432 56702 17518 56712
rect 17432 56636 17442 56702
rect 17508 56636 17518 56702
rect 17432 56112 17518 56636
rect 19631 56139 20062 57452
rect 19631 54652 19651 56139
rect 20042 54652 20062 56139
rect 16241 54149 17523 54159
rect 16241 54000 16251 54149
rect 16391 54000 17523 54149
rect 16241 53990 17523 54000
rect 16747 53916 17173 53926
rect 16747 53529 16757 53916
rect 17163 53529 17173 53916
rect 16747 53519 17173 53529
rect 17432 53902 17518 53912
rect 17432 53836 17442 53902
rect 17508 53836 17518 53902
rect 17432 53312 17518 53836
rect 19631 53339 20062 54652
rect 19631 51852 19651 53339
rect 20042 51852 20062 53339
rect 16241 51349 17523 51359
rect 16241 51200 16251 51349
rect 16391 51200 17523 51349
rect 16241 51190 17523 51200
rect 16747 51116 17173 51126
rect 16747 50729 16757 51116
rect 17163 50729 17173 51116
rect 16747 50719 17173 50729
rect 17432 51102 17518 51112
rect 17432 51036 17442 51102
rect 17508 51036 17518 51102
rect 17432 50512 17518 51036
rect 19631 50539 20062 51852
rect 19631 49052 19651 50539
rect 20042 49052 20062 50539
rect 16241 48549 17523 48559
rect 16241 48400 16251 48549
rect 16391 48400 17523 48549
rect 16241 48390 17523 48400
rect 16747 48316 17173 48326
rect 16747 47929 16757 48316
rect 17163 47929 17173 48316
rect 16747 47919 17173 47929
rect 17432 48302 17518 48312
rect 17432 48236 17442 48302
rect 17508 48236 17518 48302
rect 17432 47712 17518 48236
rect 19631 47739 20062 49052
rect 19631 46252 19651 47739
rect 20042 46252 20062 47739
rect 16241 45749 17523 45759
rect 16241 45600 16251 45749
rect 16391 45600 17523 45749
rect 16241 45590 17523 45600
rect 16747 45516 17173 45526
rect 16747 45129 16757 45516
rect 17163 45129 17173 45516
rect 16747 45119 17173 45129
rect 17432 45502 17518 45512
rect 17432 45436 17442 45502
rect 17508 45436 17518 45502
rect 17432 44912 17518 45436
rect 19631 44939 20062 46252
rect 19631 43452 19651 44939
rect 20042 43452 20062 44939
rect 16241 42949 17523 42959
rect 16241 42800 16251 42949
rect 16391 42800 17523 42949
rect 16241 42790 17523 42800
rect 16747 42716 17173 42726
rect 16747 42329 16757 42716
rect 17163 42329 17173 42716
rect 16747 42319 17173 42329
rect 17432 42702 17518 42712
rect 17432 42636 17442 42702
rect 17508 42636 17518 42702
rect 17432 42112 17518 42636
rect 19631 42139 20062 43452
rect 19631 40652 19651 42139
rect 20042 40652 20062 42139
rect 16241 40149 17523 40159
rect 16241 40000 16251 40149
rect 16391 40000 17523 40149
rect 16241 39990 17523 40000
rect 16747 39916 17173 39926
rect 16747 39529 16757 39916
rect 17163 39529 17173 39916
rect 16747 39519 17173 39529
rect 17432 39902 17518 39912
rect 17432 39836 17442 39902
rect 17508 39836 17518 39902
rect 17432 39312 17518 39836
rect 19631 39339 20062 40652
rect 19631 37852 19651 39339
rect 20042 37852 20062 39339
rect 16241 37349 17523 37359
rect 16241 37200 16251 37349
rect 16391 37200 17523 37349
rect 16241 37190 17523 37200
rect 16747 37116 17173 37126
rect 16747 36729 16757 37116
rect 17163 36729 17173 37116
rect 16747 36719 17173 36729
rect 17432 37102 17518 37112
rect 17432 37036 17442 37102
rect 17508 37036 17518 37102
rect 17432 36512 17518 37036
rect 19631 36539 20062 37852
rect 19631 35052 19651 36539
rect 20042 35052 20062 36539
rect 16241 34549 17523 34559
rect 16241 34400 16251 34549
rect 16391 34400 17523 34549
rect 16241 34390 17523 34400
rect 16747 34316 17173 34326
rect 16747 33929 16757 34316
rect 17163 33929 17173 34316
rect 16747 33919 17173 33929
rect 17432 34302 17518 34312
rect 17432 34236 17442 34302
rect 17508 34236 17518 34302
rect 17432 33712 17518 34236
rect 19631 33739 20062 35052
rect 19631 32252 19651 33739
rect 20042 32252 20062 33739
rect 16241 31749 17523 31759
rect 16241 31600 16251 31749
rect 16391 31600 17523 31749
rect 16241 31590 17523 31600
rect 16747 31516 17173 31526
rect 16747 31129 16757 31516
rect 17163 31129 17173 31516
rect 16747 31119 17173 31129
rect 17432 31502 17518 31512
rect 17432 31436 17442 31502
rect 17508 31436 17518 31502
rect 17432 30912 17518 31436
rect 19631 30939 20062 32252
rect 19631 29452 19651 30939
rect 20042 29452 20062 30939
rect 16241 28949 17523 28959
rect 16241 28800 16251 28949
rect 16391 28800 17523 28949
rect 16241 28790 17523 28800
rect 16747 28716 17173 28726
rect 16747 28329 16757 28716
rect 17163 28329 17173 28716
rect 16747 28319 17173 28329
rect 17432 28702 17518 28712
rect 17432 28636 17442 28702
rect 17508 28636 17518 28702
rect 17432 28112 17518 28636
rect 19631 28139 20062 29452
rect 19631 26652 19651 28139
rect 20042 26652 20062 28139
rect 16241 26149 17523 26159
rect 16241 26000 16251 26149
rect 16391 26000 17523 26149
rect 16241 25990 17523 26000
rect 16747 25916 17173 25926
rect 16747 25529 16757 25916
rect 17163 25529 17173 25916
rect 16747 25519 17173 25529
rect 17432 25902 17518 25912
rect 17432 25836 17442 25902
rect 17508 25836 17518 25902
rect 17432 25312 17518 25836
rect 19631 25339 20062 26652
rect 19631 23852 19651 25339
rect 20042 23852 20062 25339
rect 16241 23349 17523 23359
rect 16241 23200 16251 23349
rect 16391 23200 17523 23349
rect 16241 23190 17523 23200
rect 16747 23116 17173 23126
rect 16747 22729 16757 23116
rect 17163 22729 17173 23116
rect 16747 22719 17173 22729
rect 17432 23102 17518 23112
rect 17432 23036 17442 23102
rect 17508 23036 17518 23102
rect 17432 22512 17518 23036
rect 19631 22539 20062 23852
rect 19631 21052 19651 22539
rect 20042 21052 20062 22539
rect 16241 20549 17523 20559
rect 16241 20400 16251 20549
rect 16391 20400 17523 20549
rect 16241 20390 17523 20400
rect 16747 20316 17173 20326
rect 16747 19929 16757 20316
rect 17163 19929 17173 20316
rect 16747 19919 17173 19929
rect 17432 20302 17518 20312
rect 17432 20236 17442 20302
rect 17508 20236 17518 20302
rect 17432 19712 17518 20236
rect 19631 19739 20062 21052
rect 19631 18252 19651 19739
rect 20042 18252 20062 19739
rect 16241 17749 17523 17759
rect 16241 17600 16251 17749
rect 16391 17600 17523 17749
rect 16241 17590 17523 17600
rect 14226 17450 16178 17576
rect 19631 17451 20062 18252
rect 20224 62963 21842 63063
rect 20224 62463 20324 62963
rect 21742 62463 21842 62963
rect 20224 62363 21842 62463
rect 26356 62963 27860 63063
rect 20224 62109 20655 62363
rect 20224 61778 20244 62109
rect 20635 61778 20655 62109
rect 20224 59309 20655 61778
rect 20224 58978 20244 59309
rect 20635 58978 20655 59309
rect 20224 56509 20655 58978
rect 20224 56178 20244 56509
rect 20635 56178 20655 56509
rect 20224 53709 20655 56178
rect 20224 53378 20244 53709
rect 20635 53378 20655 53709
rect 20224 50909 20655 53378
rect 20224 50578 20244 50909
rect 20635 50578 20655 50909
rect 20224 48109 20655 50578
rect 20224 47778 20244 48109
rect 20635 47778 20655 48109
rect 20224 45309 20655 47778
rect 20224 44978 20244 45309
rect 20635 44978 20655 45309
rect 20224 42509 20655 44978
rect 20224 42178 20244 42509
rect 20635 42178 20655 42509
rect 20224 39709 20655 42178
rect 20224 39378 20244 39709
rect 20635 39378 20655 39709
rect 20224 36909 20655 39378
rect 20224 36578 20244 36909
rect 20635 36578 20655 36909
rect 20224 34109 20655 36578
rect 20224 33778 20244 34109
rect 20635 33778 20655 34109
rect 26356 62263 26456 62963
rect 27760 62263 27860 62963
rect 26356 62163 27860 62263
rect 28404 62963 33037 63063
rect 28404 62263 28504 62963
rect 32937 62263 33037 62963
rect 28404 62163 33037 62263
rect 54000 62963 58632 63063
rect 54000 62263 54100 62963
rect 58532 62263 58632 62963
rect 54000 62163 58632 62263
rect 59036 62963 63078 63063
rect 59036 62263 59136 62963
rect 62978 62263 63078 62963
rect 64909 62963 68168 63063
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 62263 68168 62363
rect 71457 62970 75284 63070
rect 71457 62283 71557 62970
rect 75184 62283 75284 62970
rect 59036 62163 63078 62263
rect 71457 62183 75284 62283
rect 26356 61969 27432 62163
rect 26356 34278 26556 61969
rect 27232 34278 27432 61969
rect 57910 62063 58632 62163
rect 42109 41817 42490 42569
rect 57910 42279 58110 62063
rect 58432 42279 58632 62063
rect 64620 61928 70907 62139
rect 64620 61828 64840 61928
rect 70717 56705 70907 61928
rect 70717 56505 70727 56705
rect 70897 56505 70907 56705
rect 70717 56495 70907 56505
rect 71137 61688 73477 61899
rect 71137 56705 71327 61688
rect 73338 61659 73477 61688
rect 75508 61565 75908 67159
rect 76099 61705 76949 61805
rect 71137 56505 71147 56705
rect 71317 56505 71327 56705
rect 71137 56495 71327 56505
rect 70343 55335 72232 55532
rect 57910 42079 58632 42279
rect 58967 51939 59520 52132
rect 42109 41436 42951 41817
rect 26356 34078 27432 34278
rect 42570 34359 42951 41436
rect 58967 40607 59348 51939
rect 58967 40246 58977 40607
rect 59338 40246 59348 40607
rect 70343 40519 70540 55335
rect 71536 54947 72253 55144
rect 71536 41602 71917 54947
rect 71536 41259 71546 41602
rect 71907 41259 71917 41602
rect 71536 41249 71917 41259
rect 62933 40509 70540 40519
rect 62933 40329 62943 40509
rect 63113 40329 67979 40509
rect 68149 40329 70540 40509
rect 62933 40319 70540 40329
rect 58967 40236 59348 40246
rect 63353 40009 68579 40019
rect 63353 39829 63363 40009
rect 63533 39829 68399 40009
rect 68569 39829 68579 40009
rect 63353 39819 68579 39829
rect 72648 39519 72848 52817
rect 65873 39509 72848 39519
rect 65873 39329 65883 39509
rect 66053 39329 68819 39509
rect 68989 39329 72848 39509
rect 65873 39319 72848 39329
rect 73248 39019 73448 52817
rect 65453 39009 73448 39019
rect 65453 38829 65463 39009
rect 65633 38829 69239 39009
rect 69409 38829 73448 39009
rect 65453 38819 73448 38829
rect 73848 38519 74048 52817
rect 65033 38509 74048 38519
rect 65033 38329 65043 38509
rect 65213 38329 69659 38509
rect 69829 38329 74048 38509
rect 65033 38319 74048 38329
rect 74448 38019 74648 52817
rect 64613 38009 74648 38019
rect 64613 37829 64623 38009
rect 64793 37829 70079 38009
rect 70249 37829 74648 38009
rect 64613 37819 74648 37829
rect 75048 37519 75248 52817
rect 64193 37509 75248 37519
rect 64193 37329 64203 37509
rect 64373 37329 70499 37509
rect 70669 37329 75248 37509
rect 64193 37319 75248 37329
rect 75648 37019 75848 52817
rect 76099 52782 76199 61705
rect 76849 52782 76949 61705
rect 76099 52682 76949 52782
rect 63773 37009 75848 37019
rect 63773 36829 63783 37009
rect 63953 36829 70919 37009
rect 71089 36829 75848 37009
rect 63773 36819 75848 36829
rect 76309 52131 76709 52141
rect 76309 51751 76319 52131
rect 76699 51751 76709 52131
rect 76309 36525 76709 51751
rect 81212 37033 81612 37133
rect 60413 36515 76709 36525
rect 60413 36335 60423 36515
rect 60593 36335 76709 36515
rect 60413 36325 76709 36335
rect 80417 36833 81612 37033
rect 80417 36025 80617 36833
rect 81212 36733 81612 36833
rect 60833 36015 80617 36025
rect 81212 36022 81612 36122
rect 60833 35835 60843 36015
rect 61013 35835 80617 36015
rect 60833 35825 80617 35835
rect 80861 35822 81612 36022
rect 80861 35525 81061 35822
rect 81212 35722 81612 35822
rect 61253 35515 81061 35525
rect 61253 35335 61263 35515
rect 61433 35335 81061 35515
rect 61253 35325 81061 35335
rect 81212 35025 81612 35125
rect 61673 35015 81612 35025
rect 61673 34835 61683 35015
rect 61853 34835 81612 35015
rect 61673 34825 81612 34835
rect 81212 34725 81612 34825
rect 42570 34068 42580 34359
rect 42941 34068 42951 34359
rect 62093 34515 81061 34525
rect 62093 34335 62103 34515
rect 62273 34335 81061 34515
rect 62093 34325 81061 34335
rect 42570 34058 42951 34068
rect 62513 34015 80608 34025
rect 62513 33835 62523 34015
rect 62693 33835 80608 34015
rect 62513 33825 80608 33835
rect 20224 31309 20655 33778
rect 21124 33508 67323 33518
rect 21124 33328 21134 33508
rect 21314 33328 67143 33508
rect 67313 33328 67323 33508
rect 21124 33318 67323 33328
rect 21124 33008 67743 33018
rect 21124 32828 21134 33008
rect 21314 32828 67563 33008
rect 67733 32828 67743 33008
rect 21124 32818 67743 32828
rect 80408 33012 80608 33825
rect 80861 34023 81061 34325
rect 81212 34023 81612 34123
rect 80861 33823 81612 34023
rect 81212 33723 81612 33823
rect 81212 33012 81612 33112
rect 80408 32812 81612 33012
rect 81212 32712 81612 32812
rect 21596 32508 66903 32518
rect 21596 32328 21606 32508
rect 21786 32328 66723 32508
rect 66893 32328 66903 32508
rect 21596 32318 66903 32328
rect 21596 32008 68163 32018
rect 21596 31828 21606 32008
rect 21786 31828 67983 32008
rect 68153 31828 68163 32008
rect 21596 31818 68163 31828
rect 22068 31508 66483 31518
rect 22068 31328 22078 31508
rect 22258 31328 66303 31508
rect 66473 31328 66483 31508
rect 22068 31318 66483 31328
rect 20224 30978 20244 31309
rect 20635 30978 20655 31309
rect 20224 28509 20655 30978
rect 22068 31008 68583 31018
rect 22068 30828 22078 31008
rect 22258 30828 68403 31008
rect 68573 30828 68583 31008
rect 22068 30818 68583 30828
rect 22540 30508 72783 30518
rect 22540 30328 22550 30508
rect 22730 30328 72603 30508
rect 72773 30328 72783 30508
rect 22540 30318 72783 30328
rect 22540 30008 69003 30018
rect 22540 29828 22550 30008
rect 22730 29828 68823 30008
rect 68993 29828 69003 30008
rect 22540 29818 69003 29828
rect 23012 29508 72363 29518
rect 23012 29328 23022 29508
rect 23202 29328 72183 29508
rect 72353 29328 72363 29508
rect 23012 29318 72363 29328
rect 23012 29008 69423 29018
rect 23012 28828 23022 29008
rect 23202 28828 69243 29008
rect 69413 28828 69423 29008
rect 23012 28818 69423 28828
rect 20224 28178 20244 28509
rect 20635 28178 20655 28509
rect 23484 28508 71943 28518
rect 23484 28328 23494 28508
rect 23674 28328 71763 28508
rect 71933 28328 71943 28508
rect 23484 28318 71943 28328
rect 20224 25709 20655 28178
rect 23956 28008 71523 28018
rect 23956 27828 23966 28008
rect 24146 27828 71343 28008
rect 71513 27828 71523 28008
rect 23956 27818 71523 27828
rect 24428 27508 71103 27518
rect 24428 27328 24438 27508
rect 24618 27328 70923 27508
rect 71093 27328 71103 27508
rect 24428 27318 71103 27328
rect 24900 27008 70683 27018
rect 24900 26828 24910 27008
rect 25090 26828 70503 27008
rect 70673 26828 70683 27008
rect 24900 26818 70683 26828
rect 25372 26508 70263 26518
rect 25372 26328 25382 26508
rect 25562 26328 70083 26508
rect 70253 26328 70263 26508
rect 25372 26318 70263 26328
rect 25844 26008 69843 26018
rect 25844 25828 25854 26008
rect 26034 25828 69663 26008
rect 69833 25828 69843 26008
rect 25844 25818 69843 25828
rect 20224 25378 20244 25709
rect 20635 25378 20655 25709
rect 20224 22909 20655 25378
rect 60413 24612 60603 24622
rect 60413 24431 60423 24612
rect 60593 24431 60603 24612
rect 60413 24421 60603 24431
rect 60833 24612 61023 24622
rect 60833 24431 60843 24612
rect 61013 24431 61023 24612
rect 60833 24421 61023 24431
rect 61253 24612 61443 24622
rect 61253 24431 61263 24612
rect 61433 24431 61443 24612
rect 61253 24421 61443 24431
rect 61673 24612 61863 24622
rect 61673 24431 61683 24612
rect 61853 24431 61863 24612
rect 61673 24421 61863 24431
rect 62093 24612 62283 24622
rect 62093 24431 62103 24612
rect 62273 24431 62283 24612
rect 62093 24421 62283 24431
rect 62513 24612 62703 24622
rect 62513 24431 62523 24612
rect 62693 24431 62703 24612
rect 62513 24421 62703 24431
rect 62933 24612 63123 24622
rect 62933 24431 62943 24612
rect 63113 24431 63123 24612
rect 62933 24421 63123 24431
rect 63353 24612 63543 24622
rect 63353 24431 63363 24612
rect 63533 24431 63543 24612
rect 63353 24421 63543 24431
rect 63773 24612 63963 24622
rect 63773 24431 63783 24612
rect 63953 24431 63963 24612
rect 63773 24421 63963 24431
rect 64193 24612 64383 24622
rect 64193 24431 64203 24612
rect 64373 24431 64383 24612
rect 64193 24421 64383 24431
rect 64613 24612 64803 24622
rect 64613 24431 64623 24612
rect 64793 24431 64803 24612
rect 64613 24421 64803 24431
rect 65033 24612 65223 24622
rect 65033 24431 65043 24612
rect 65213 24431 65223 24612
rect 65033 24421 65223 24431
rect 65453 24612 65643 24622
rect 65453 24431 65463 24612
rect 65633 24431 65643 24612
rect 65453 24421 65643 24431
rect 65873 24612 66063 24622
rect 65873 24431 65883 24612
rect 66053 24431 66063 24612
rect 65873 24421 66063 24431
rect 66293 24612 66483 24622
rect 66293 24431 66303 24612
rect 66473 24431 66483 24612
rect 66293 24421 66483 24431
rect 66713 24612 66903 24622
rect 66713 24431 66723 24612
rect 66893 24431 66903 24612
rect 66713 24421 66903 24431
rect 67133 24612 67323 24622
rect 67133 24431 67143 24612
rect 67313 24431 67323 24612
rect 67133 24421 67323 24431
rect 67553 24612 67743 24622
rect 67553 24431 67563 24612
rect 67733 24431 67743 24612
rect 67553 24421 67743 24431
rect 67973 24612 68163 24622
rect 67973 24431 67983 24612
rect 68153 24431 68163 24612
rect 67973 24421 68163 24431
rect 68393 24612 68583 24622
rect 68393 24431 68403 24612
rect 68573 24431 68583 24612
rect 68393 24421 68583 24431
rect 68813 24612 69003 24622
rect 68813 24431 68823 24612
rect 68993 24431 69003 24612
rect 68813 24421 69003 24431
rect 69233 24612 69423 24622
rect 69233 24431 69243 24612
rect 69413 24431 69423 24612
rect 69233 24421 69423 24431
rect 69653 24612 69843 24622
rect 69653 24431 69663 24612
rect 69833 24431 69843 24612
rect 69653 24421 69843 24431
rect 70073 24612 70263 24622
rect 70073 24431 70083 24612
rect 70253 24431 70263 24612
rect 70073 24421 70263 24431
rect 70493 24612 70683 24622
rect 70493 24431 70503 24612
rect 70673 24431 70683 24612
rect 70493 24421 70683 24431
rect 70913 24612 71103 24622
rect 70913 24431 70923 24612
rect 71093 24431 71103 24612
rect 70913 24421 71103 24431
rect 71333 24612 71523 24622
rect 71333 24431 71343 24612
rect 71513 24431 71523 24612
rect 71333 24421 71523 24431
rect 71753 24612 71943 24622
rect 71753 24431 71763 24612
rect 71933 24431 71943 24612
rect 71753 24421 71943 24431
rect 72173 24612 72363 24622
rect 72173 24431 72183 24612
rect 72353 24431 72363 24612
rect 72173 24421 72363 24431
rect 72593 24612 72783 24622
rect 72593 24431 72603 24612
rect 72773 24431 72783 24612
rect 72593 24421 72783 24431
rect 73013 24612 73203 24622
rect 73013 24431 73023 24612
rect 73193 24431 73203 24612
rect 73013 24421 73203 24431
rect 73433 24612 73623 24622
rect 73433 24431 73443 24612
rect 73613 24431 73623 24612
rect 73433 24421 73623 24431
rect 73853 24612 74043 24622
rect 73853 24431 73863 24612
rect 74033 24431 74043 24612
rect 73853 24421 74043 24431
rect 74273 24612 74463 24622
rect 74273 24431 74283 24612
rect 74453 24431 74463 24612
rect 74273 24421 74463 24431
rect 74693 24612 74883 24622
rect 74693 24431 74703 24612
rect 74873 24431 74883 24612
rect 74693 24421 74883 24431
rect 75113 24612 75303 24622
rect 75113 24431 75123 24612
rect 75293 24431 75303 24612
rect 75113 24421 75303 24431
rect 75533 24612 75723 24622
rect 75533 24431 75543 24612
rect 75713 24431 75723 24612
rect 75533 24421 75723 24431
rect 75953 24612 76143 24622
rect 75953 24431 75963 24612
rect 76133 24431 76143 24612
rect 75953 24421 76143 24431
rect 20224 22578 20244 22909
rect 20635 22578 20655 22909
rect 20224 20109 20655 22578
rect 20224 19778 20244 20109
rect 20635 19778 20655 20109
rect 20224 17451 20655 19778
rect 538 15531 12911 16731
rect -1354 13639 10705 14839
rect -2014 12385 -1145 12485
rect -2014 1885 -1914 12385
rect -1245 1885 -1145 12385
rect -2014 1785 -1145 1885
rect 9367 1041 10705 13639
rect 11397 1041 12911 15531
rect 27820 14620 30223 14630
rect 27820 14290 27830 14620
rect 28192 14290 30223 14620
rect 27820 14280 30223 14290
rect 28847 13602 29228 13612
rect 28847 13272 28857 13602
rect 29218 13272 29228 13602
rect 22075 1569 22746 1579
rect 9367 585 12911 1041
rect 13048 -56 14114 44
rect -912 -602 9370 -502
rect -912 -1416 -812 -602
rect 9270 -1416 9370 -602
rect 13048 -657 13148 -56
rect 14014 -657 14114 -56
rect 13048 -757 14114 -657
rect 14438 -57 18572 43
rect 14438 -657 14538 -57
rect 18472 -657 18572 -57
rect 14438 -757 18572 -657
rect 19437 -271 19849 1549
rect 22075 1509 22085 1569
rect 20819 1157 22085 1509
rect 20819 298 21171 1157
rect 22075 1113 22085 1157
rect 22736 1113 22746 1569
rect 22075 1103 22746 1113
rect 28847 329 29228 13272
rect 20819 -34 20829 298
rect 21161 -34 21171 298
rect 20819 -44 21171 -34
rect 21577 -83 29228 329
rect 21577 -271 21989 -83
rect 19437 -683 21989 -271
rect 22953 -369 28430 -269
rect 22953 -669 23053 -369
rect 28330 -669 28430 -369
rect 22953 -769 28430 -669
rect 29841 -413 30223 14280
rect 47022 12800 50637 14090
rect 47349 12558 48289 12658
rect 30469 12447 31020 12547
rect 30469 4302 30569 12447
rect 30920 4302 31020 12447
rect 30469 4202 31020 4302
rect 39592 1536 42592 1546
rect 39592 1281 39602 1536
rect 42582 1281 42592 1536
rect 30354 622 33209 722
rect 30354 -166 30454 622
rect 33109 -166 33209 622
rect 33443 332 33796 982
rect 33443 -10 33453 332
rect 33786 -10 33796 332
rect 33443 -20 33796 -10
rect 30354 -266 33209 -166
rect 35935 -413 36317 981
rect 37125 332 37478 940
rect 37125 -10 37135 332
rect 37468 -10 37478 332
rect 37125 -20 37478 -10
rect 29841 -795 36317 -413
rect 37626 -949 37978 939
rect 39592 244 42592 1281
rect 47349 670 47858 12558
rect 48189 670 48289 12558
rect 47349 570 48289 670
rect 39592 -265 39692 244
rect 42492 -265 42592 244
rect 39592 -365 42592 -265
rect 44588 470 48289 570
rect 44588 -261 44688 470
rect 48189 -261 48289 470
rect 44588 -361 48289 -261
rect 20819 -959 37978 -949
rect 20819 -1291 20829 -959
rect 21161 -1291 37978 -959
rect 20819 -1301 37978 -1291
rect -912 -1516 9370 -1416
rect 48470 -5827 50637 12800
<< via2 >>
rect 2757 62466 15645 62966
rect 16341 62663 18013 62963
rect 18544 62463 19962 62963
rect -154 15531 538 61158
rect 15027 17576 15499 62003
rect 16757 61929 17163 62316
rect 19651 60252 20042 61739
rect 16757 59129 17163 59516
rect 19651 57452 20042 58939
rect 16757 56329 17163 56716
rect 19651 54652 20042 56139
rect 16757 53529 17163 53916
rect 19651 51852 20042 53339
rect 16757 50729 17163 51116
rect 19651 49052 20042 50539
rect 16757 47929 17163 48316
rect 19651 46252 20042 47739
rect 16757 45129 17163 45516
rect 19651 43452 20042 44939
rect 16757 42329 17163 42716
rect 19651 40652 20042 42139
rect 16757 39529 17163 39916
rect 19651 37852 20042 39339
rect 16757 36729 17163 37116
rect 19651 35052 20042 36539
rect 16757 33929 17163 34316
rect 19651 32252 20042 33739
rect 16757 31129 17163 31516
rect 19651 29452 20042 30939
rect 16757 28329 17163 28716
rect 19651 26652 20042 28139
rect 16757 25529 17163 25916
rect 19651 23852 20042 25339
rect 16757 22729 17163 23116
rect 19651 21052 20042 22539
rect 16757 19929 17163 20316
rect 19651 18252 20042 19739
rect 20324 62463 21742 62963
rect 20244 61778 20635 62109
rect 20244 58978 20635 59309
rect 20244 56178 20635 56509
rect 20244 53378 20635 53709
rect 20244 50578 20635 50909
rect 20244 47778 20635 48109
rect 20244 44978 20635 45309
rect 20244 42178 20635 42509
rect 20244 39378 20635 39709
rect 20244 36578 20635 36909
rect 20244 33778 20635 34109
rect 26456 62263 27760 62963
rect 28504 62263 32937 62963
rect 54100 62263 58532 62963
rect 59136 62263 62978 62963
rect 65009 62363 68068 62963
rect 71557 62283 75184 62970
rect 26556 34278 27232 61969
rect 58110 42279 58432 62063
rect 76199 52782 76849 61705
rect 20244 30978 20635 31309
rect 20244 28178 20635 28509
rect 20244 25378 20635 25709
rect 20244 22578 20635 22909
rect 20244 19778 20635 20109
rect -154 14839 11397 15531
rect -1914 1885 -1245 12385
rect 10705 1041 11397 14839
rect -812 -1416 9270 -602
rect 13148 -657 14014 -56
rect 14538 -657 18472 -57
rect 23053 -669 28330 -369
rect 30569 4302 30920 12447
rect 30454 -166 33109 622
rect 47858 670 48189 12558
rect 39692 -265 42492 244
rect 44688 -261 48189 470
<< metal3 >>
rect -5353 63359 80237 66359
rect -5353 12485 -2353 63359
rect 2657 62966 15745 63066
rect 2657 62466 2757 62966
rect 15645 62466 15745 62966
rect 16241 62963 18113 63063
rect 16241 62663 16341 62963
rect 18013 62663 18113 62963
rect 16241 62563 18113 62663
rect 18444 62963 20062 63359
rect 2657 62358 15745 62466
rect 18444 62463 18544 62963
rect 19962 62463 20062 62963
rect 18444 62364 20062 62463
rect -1354 61158 1738 62358
rect 2657 62003 16178 62358
rect 2657 61956 15027 62003
rect -1354 14839 -154 61158
rect 538 16731 1738 61158
rect 14226 59558 15027 61956
rect 2657 59156 15027 59558
rect 14226 56758 15027 59156
rect 2657 56356 15027 56758
rect 14226 53958 15027 56356
rect 2657 53556 15027 53958
rect 14226 51158 15027 53556
rect 2657 50756 15027 51158
rect 14226 48358 15027 50756
rect 2657 47956 15027 48358
rect 14226 45558 15027 47956
rect 2657 45156 15027 45558
rect 14226 42758 15027 45156
rect 2657 42356 15027 42758
rect 14226 39958 15027 42356
rect 2657 39556 15027 39958
rect 14226 37158 15027 39556
rect 2657 36756 15027 37158
rect 14226 34358 15027 36756
rect 2657 33956 15027 34358
rect 14226 31558 15027 33956
rect 2657 31156 15027 31558
rect 14226 28758 15027 31156
rect 2657 28356 15027 28758
rect 14226 25958 15027 28356
rect 2657 25556 15027 25958
rect 14226 23158 15027 25556
rect 2657 22756 15027 23158
rect 14226 20358 15027 22756
rect 2657 19956 15027 20358
rect 14226 17576 15027 19956
rect 15499 17576 16178 62003
rect 16747 62316 17173 62326
rect 16747 61929 16757 62316
rect 17163 61929 17173 62316
rect 16747 61919 17173 61929
rect 19631 61739 20062 62364
rect 19631 60252 19651 61739
rect 20042 60252 20062 61739
rect 16747 59516 17173 59526
rect 16747 59129 16757 59516
rect 17163 59129 17173 59516
rect 16747 59119 17173 59129
rect 19631 58939 20062 60252
rect 19631 57452 19651 58939
rect 20042 57452 20062 58939
rect 16747 56716 17173 56726
rect 16747 56329 16757 56716
rect 17163 56329 17173 56716
rect 16747 56319 17173 56329
rect 19631 56139 20062 57452
rect 19631 54652 19651 56139
rect 20042 54652 20062 56139
rect 16747 53916 17173 53926
rect 16747 53529 16757 53916
rect 17163 53529 17173 53916
rect 16747 53519 17173 53529
rect 19631 53339 20062 54652
rect 19631 51852 19651 53339
rect 20042 51852 20062 53339
rect 16747 51116 17173 51126
rect 16747 50729 16757 51116
rect 17163 50729 17173 51116
rect 16747 50719 17173 50729
rect 19631 50539 20062 51852
rect 19631 49052 19651 50539
rect 20042 49052 20062 50539
rect 16747 48316 17173 48326
rect 16747 47929 16757 48316
rect 17163 47929 17173 48316
rect 16747 47919 17173 47929
rect 19631 47739 20062 49052
rect 19631 46252 19651 47739
rect 20042 46252 20062 47739
rect 16747 45516 17173 45526
rect 16747 45129 16757 45516
rect 17163 45129 17173 45516
rect 16747 45119 17173 45129
rect 19631 44939 20062 46252
rect 19631 43452 19651 44939
rect 20042 43452 20062 44939
rect 16747 42716 17173 42726
rect 16747 42329 16757 42716
rect 17163 42329 17173 42716
rect 16747 42319 17173 42329
rect 19631 42139 20062 43452
rect 19631 40652 19651 42139
rect 20042 40652 20062 42139
rect 16747 39916 17173 39926
rect 16747 39529 16757 39916
rect 17163 39529 17173 39916
rect 16747 39519 17173 39529
rect 19631 39339 20062 40652
rect 19631 37852 19651 39339
rect 20042 37852 20062 39339
rect 16747 37116 17173 37126
rect 16747 36729 16757 37116
rect 17163 36729 17173 37116
rect 16747 36719 17173 36729
rect 19631 36539 20062 37852
rect 19631 35052 19651 36539
rect 20042 35052 20062 36539
rect 16747 34316 17173 34326
rect 16747 33929 16757 34316
rect 17163 33929 17173 34316
rect 16747 33919 17173 33929
rect 19631 33739 20062 35052
rect 19631 32252 19651 33739
rect 20042 32252 20062 33739
rect 16747 31516 17173 31526
rect 16747 31129 16757 31516
rect 17163 31129 17173 31516
rect 16747 31119 17173 31129
rect 19631 30939 20062 32252
rect 19631 29452 19651 30939
rect 20042 29452 20062 30939
rect 16747 28716 17173 28726
rect 16747 28329 16757 28716
rect 17163 28329 17173 28716
rect 16747 28319 17173 28329
rect 19631 28139 20062 29452
rect 19631 26652 19651 28139
rect 20042 26652 20062 28139
rect 16747 25916 17173 25926
rect 16747 25529 16757 25916
rect 17163 25529 17173 25916
rect 16747 25519 17173 25529
rect 19631 25339 20062 26652
rect 19631 23852 19651 25339
rect 20042 23852 20062 25339
rect 16747 23116 17173 23126
rect 16747 22729 16757 23116
rect 17163 22729 17173 23116
rect 16747 22719 17173 22729
rect 19631 22539 20062 23852
rect 19631 21052 19651 22539
rect 20042 21052 20062 22539
rect 16747 20316 17173 20326
rect 16747 19929 16757 20316
rect 17163 19929 17173 20316
rect 16747 19919 17173 19929
rect 14226 17450 16178 17576
rect 19631 19739 20062 21052
rect 19631 18252 19651 19739
rect 20042 18252 20062 19739
rect 19631 17451 20062 18252
rect 20224 62963 21842 63063
rect 20224 62463 20324 62963
rect 21742 62463 21842 62963
rect 20224 62363 21842 62463
rect 26356 62963 27860 63359
rect 20224 62109 20655 62363
rect 20224 61778 20244 62109
rect 20635 61778 20655 62109
rect 20224 59309 20655 61778
rect 20224 58978 20244 59309
rect 20635 58978 20655 59309
rect 20224 56509 20655 58978
rect 20224 56178 20244 56509
rect 20635 56178 20655 56509
rect 20224 53709 20655 56178
rect 20224 53378 20244 53709
rect 20635 53378 20655 53709
rect 20224 50909 20655 53378
rect 20224 50578 20244 50909
rect 20635 50578 20655 50909
rect 20224 48109 20655 50578
rect 20224 47778 20244 48109
rect 20635 47778 20655 48109
rect 20224 45309 20655 47778
rect 20224 44978 20244 45309
rect 20635 44978 20655 45309
rect 20224 42509 20655 44978
rect 20224 42178 20244 42509
rect 20635 42178 20655 42509
rect 20224 39709 20655 42178
rect 20224 39378 20244 39709
rect 20635 39378 20655 39709
rect 20224 36909 20655 39378
rect 20224 36578 20244 36909
rect 20635 36578 20655 36909
rect 20224 34109 20655 36578
rect 20224 33778 20244 34109
rect 20635 33778 20655 34109
rect 26356 62263 26456 62963
rect 27760 62263 27860 62963
rect 26356 62163 27860 62263
rect 28404 62963 33037 63063
rect 28404 62263 28504 62963
rect 32937 62263 33037 62963
rect 28404 62163 33037 62263
rect 54000 62963 58632 63063
rect 54000 62263 54100 62963
rect 58532 62263 58632 62963
rect 54000 62163 58632 62263
rect 59036 62963 63078 63063
rect 59036 62263 59136 62963
rect 62978 62263 63078 62963
rect 64909 62963 68168 63063
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 62263 68168 62363
rect 71457 62970 75284 63070
rect 71457 62283 71557 62970
rect 75184 62283 75284 62970
rect 59036 62163 63078 62263
rect 71457 62183 75284 62283
rect 26356 61969 27432 62163
rect 26356 34278 26556 61969
rect 27232 34278 27432 61969
rect 57910 62063 58632 62163
rect 57910 42279 58110 62063
rect 58432 42279 58632 62063
rect 76099 61705 76949 61805
rect 76099 52782 76199 61705
rect 76849 52782 76949 61705
rect 76099 52682 76949 52782
rect 57910 42079 58632 42279
rect 26356 34078 27432 34278
rect 20224 31309 20655 33778
rect 20224 30978 20244 31309
rect 20635 30978 20655 31309
rect 20224 28509 20655 30978
rect 20224 28178 20244 28509
rect 20635 28178 20655 28509
rect 20224 25709 20655 28178
rect 20224 25378 20244 25709
rect 20635 25378 20655 25709
rect 20224 22909 20655 25378
rect 20224 22578 20244 22909
rect 20635 22578 20655 22909
rect 20224 20109 20655 22578
rect 20224 19778 20244 20109
rect 20635 19778 20655 20109
rect 20224 17451 20655 19778
rect 538 15531 12911 16731
rect -1354 13639 10705 14839
rect -5353 12385 -1145 12485
rect -5353 1885 -1914 12385
rect -1245 1885 -1145 12385
rect -5353 1785 -1145 1885
rect -5353 -1027 -2353 1785
rect 9367 1041 10705 13639
rect 11397 1041 12911 15531
rect 9367 585 12911 1041
rect 30354 12447 31154 12658
rect 30354 4302 30569 12447
rect 30920 4302 31154 12447
rect 30354 722 31154 4302
rect 47349 12558 48289 12658
rect 30354 622 33209 722
rect 13048 -56 14114 44
rect -7353 -2027 -2353 -1027
rect -912 -602 9370 -502
rect -912 -1416 -812 -602
rect 9270 -1416 9370 -602
rect 13048 -657 13148 -56
rect 14014 -657 14114 -56
rect 13048 -757 14114 -657
rect 14438 -57 18572 43
rect 14438 -657 14538 -57
rect 18472 -657 18572 -57
rect 30354 -166 30454 622
rect 33109 -166 33209 622
rect 47349 670 47858 12558
rect 48189 670 48289 12558
rect 47349 570 48289 670
rect 44588 470 48289 570
rect 30354 -266 33209 -166
rect 39592 244 42592 344
rect 39592 -265 39692 244
rect 42492 -265 42592 244
rect -912 -1516 9370 -1416
rect -5353 -2028 -2353 -2027
rect 14438 -2028 18572 -657
rect 22953 -369 28430 -269
rect 39592 -365 42592 -265
rect 44588 -261 44688 470
rect 48189 -261 48289 470
rect 22953 -669 23053 -369
rect 28330 -669 28430 -369
rect 22953 -2028 28430 -669
rect 44588 -2028 48289 -261
rect 77237 -2028 80237 63359
rect -5353 -5027 80237 -2028
<< via3 >>
rect 2757 62466 15645 62966
rect 16341 62663 18013 62963
rect 16757 61929 17163 62316
rect 16757 59129 17163 59516
rect 16757 56329 17163 56716
rect 16757 53529 17163 53916
rect 16757 50729 17163 51116
rect 16757 47929 17163 48316
rect 16757 45129 17163 45516
rect 16757 42329 17163 42716
rect 16757 39529 17163 39916
rect 16757 36729 17163 37116
rect 16757 33929 17163 34316
rect 16757 31129 17163 31516
rect 16757 28329 17163 28716
rect 16757 25529 17163 25916
rect 16757 22729 17163 23116
rect 16757 19929 17163 20316
rect 20324 62463 21742 62963
rect 28504 62263 32937 62963
rect 54100 62263 58532 62963
rect 59136 62263 62978 62963
rect 65009 62363 68068 62963
rect 71557 62283 75184 62970
rect 76199 52782 76849 61705
rect -812 -1416 9270 -602
rect 13148 -657 14014 -56
rect 30454 -166 33109 622
rect 39692 -265 42492 244
<< metal4 >>
rect -5353 68259 26411 68359
rect -5353 67459 -5253 68259
rect 26311 67459 26411 68259
rect -5353 66359 26411 67459
rect -7353 66259 80237 66359
rect -7353 26725 -7253 66259
rect -6453 63359 80237 66259
rect -6453 26725 -2353 63359
rect 2657 62966 15745 63359
rect 2657 62466 2757 62966
rect 15645 62466 15745 62966
rect 2657 62366 15745 62466
rect 16241 62963 18113 63359
rect 16241 62663 16341 62963
rect 18013 62663 18113 62963
rect -7353 26625 -2353 26725
rect -5353 19004 -2353 26625
rect -7353 18004 -2353 19004
rect -5353 -2027 -2353 18004
rect 16241 62316 18113 62663
rect 20224 62963 21842 63063
rect 20224 62463 20324 62963
rect 21742 62463 21842 62963
rect 20224 62363 21842 62463
rect 28404 62963 33037 63359
rect 16241 61929 16757 62316
rect 17163 61929 18113 62316
rect 28404 62263 28504 62963
rect 32937 62263 33037 62963
rect 28404 62163 33037 62263
rect 54000 62963 58632 63359
rect 54000 62263 54100 62963
rect 58532 62263 58632 62963
rect 54000 62163 58632 62263
rect 59036 62963 63078 63063
rect 59036 62263 59136 62963
rect 62978 62263 63078 62963
rect 64909 62963 68168 63063
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 62263 68168 62363
rect 71457 62970 75284 63070
rect 71457 62283 71557 62970
rect 75184 62283 75284 62970
rect 59036 62163 63078 62263
rect 71457 62183 75284 62283
rect 16241 59516 18113 61929
rect 16241 59129 16757 59516
rect 17163 59129 18113 59516
rect 16241 56716 18113 59129
rect 16241 56329 16757 56716
rect 17163 56329 18113 56716
rect 16241 53916 18113 56329
rect 16241 53529 16757 53916
rect 17163 53529 18113 53916
rect 16241 51116 18113 53529
rect 76099 61705 76949 61805
rect 76099 52782 76199 61705
rect 76849 52782 76949 61705
rect 76099 52682 76949 52782
rect 16241 50729 16757 51116
rect 17163 50729 18113 51116
rect 16241 48316 18113 50729
rect 16241 47929 16757 48316
rect 17163 47929 18113 48316
rect 16241 45516 18113 47929
rect 16241 45129 16757 45516
rect 17163 45129 18113 45516
rect 16241 42716 18113 45129
rect 16241 42329 16757 42716
rect 17163 42329 18113 42716
rect 16241 39916 18113 42329
rect 16241 39529 16757 39916
rect 17163 39529 18113 39916
rect 16241 37116 18113 39529
rect 16241 36729 16757 37116
rect 17163 36729 18113 37116
rect 16241 34316 18113 36729
rect 16241 33929 16757 34316
rect 17163 33929 18113 34316
rect 16241 31516 18113 33929
rect 16241 31129 16757 31516
rect 17163 31129 18113 31516
rect 16241 28716 18113 31129
rect 16241 28329 16757 28716
rect 17163 28329 18113 28716
rect 16241 25916 18113 28329
rect 16241 25529 16757 25916
rect 17163 25529 18113 25916
rect 16241 23116 18113 25529
rect 16241 22729 16757 23116
rect 17163 22729 18113 23116
rect 16241 20316 18113 22729
rect 16241 19929 16757 20316
rect 17163 19929 18113 20316
rect 16241 17451 18113 19929
rect 30354 622 33209 722
rect 13048 -56 14114 44
rect -912 -602 9370 -502
rect -912 -1416 -812 -602
rect 9270 -1416 9370 -602
rect -912 -2027 9370 -1416
rect 13048 -657 13148 -56
rect 14014 -657 14114 -56
rect 13048 -2027 14114 -657
rect 30354 -166 30454 622
rect 33109 -166 33209 622
rect 30354 -2027 33209 -166
rect 39592 244 42592 344
rect 39592 -265 39692 244
rect 42492 -265 42592 244
rect 39592 -2027 42592 -265
rect 77237 -2027 80237 63359
rect -5353 -5027 80237 -2027
<< via4 >>
rect -5253 67459 26311 68259
rect -7253 26725 -6453 66259
rect 20324 62463 21742 62963
rect 59136 62263 62978 62963
rect 65009 62363 68068 62963
rect 71557 62283 75184 62970
rect 76199 52782 76849 61705
<< metal5 >>
rect -5353 68259 26411 68359
rect -5353 67459 -5253 68259
rect 26311 67459 26411 68259
rect -5353 67359 26411 67459
rect 56769 66359 57769 68359
rect -7353 66259 -6353 66359
rect -7353 26725 -7253 66259
rect -6453 26725 -6353 66259
rect -7353 26625 -6353 26725
rect -5353 63359 80237 66359
rect -5353 -2027 -2353 63359
rect 20224 62963 21842 63359
rect 20224 62463 20324 62963
rect 21742 62463 21842 62963
rect 20224 62363 21842 62463
rect 59036 62963 63078 63359
rect 59036 62263 59136 62963
rect 62978 62263 63078 62963
rect 64909 62963 68168 63063
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 62263 68168 62363
rect 71457 62970 75284 63359
rect 71457 62283 71557 62970
rect 75184 62283 75284 62970
rect 59036 62163 63078 62263
rect 71457 62183 75284 62283
rect 76099 61705 76949 61805
rect 76099 52782 76199 61705
rect 76849 52782 76949 61705
rect 76099 52682 76949 52782
rect 58893 392 61675 492
rect 58893 -408 58993 392
rect 61575 -408 61675 392
rect 58893 -2027 61675 -408
rect 67544 392 70326 492
rect 67544 -408 67644 392
rect 70226 -408 70326 392
rect 67544 -2027 70326 -408
rect 77237 -2027 80237 63359
rect -5353 -5027 80237 -2027
<< via5 >>
rect -5253 67459 26311 68259
rect -7253 26725 -6453 66259
rect 65009 62363 68068 62963
rect 76199 52782 76849 61705
rect 58993 -408 61575 392
rect 67644 -408 70226 392
<< metal6 >>
rect -5353 68259 26411 68359
rect -5353 67459 -5253 68259
rect 26311 67459 26411 68259
rect -5353 66359 26411 67459
rect 36394 66359 37394 68359
rect -7353 66259 80237 66359
rect -7353 26725 -7253 66259
rect -6453 63359 80237 66259
rect -6453 26725 -2353 63359
rect 64909 62963 68168 63359
rect 64909 62363 65009 62963
rect 68068 62363 68168 62963
rect 64909 62263 68168 62363
rect 77237 61805 80237 63359
rect 76099 61705 80237 61805
rect 76099 52782 76199 61705
rect 76849 52782 80237 61705
rect 76099 52682 80237 52782
rect -7353 26625 -2353 26725
rect -5353 -2027 -2353 26625
rect 52317 1792 57157 1892
rect 52317 992 53417 1792
rect 56617 992 57157 1792
rect 52317 -2027 57157 992
rect 71837 1792 74835 1892
rect 71837 992 72377 1792
rect 73737 992 74835 1792
rect 58893 392 61675 492
rect 58893 -408 58993 392
rect 61575 -408 61675 392
rect 58893 -508 61675 -408
rect 67544 392 70326 492
rect 67544 -408 67644 392
rect 70226 -408 70326 392
rect 67544 -508 70326 -408
rect 71837 -2027 74835 992
rect 77237 -2027 80237 52682
rect -5353 -5027 80237 -2027
<< via6 >>
rect 53417 992 56617 1792
rect 72377 992 73737 1792
rect 58993 -408 61575 392
rect 67644 -408 70226 392
use bmbg  bmbg_0 ../ip/bmbg/magic
timestamp 1748629122
transform -1 0 22041 0 -1 3880
box -6389 -9462 7678 3287
use fuse  fuse_0 ../ip/util/magic
timestamp 1757447377
transform 1 0 1743 0 1 18525
box -586 -1075 12571 1441
use fuse  fuse_1
timestamp 1757447377
transform 1 0 1743 0 1 21325
box -586 -1075 12571 1441
use fuse  fuse_2
timestamp 1757447377
transform 1 0 1743 0 1 24125
box -586 -1075 12571 1441
use fuse  fuse_3
timestamp 1757447377
transform 1 0 1743 0 1 26925
box -586 -1075 12571 1441
use fuse  fuse_4
timestamp 1757447377
transform 1 0 1743 0 1 29725
box -586 -1075 12571 1441
use fuse  fuse_5
timestamp 1757447377
transform 1 0 1743 0 1 32525
box -586 -1075 12571 1441
use fuse  fuse_6
timestamp 1757447377
transform 1 0 1743 0 1 35325
box -586 -1075 12571 1441
use fuse  fuse_7
timestamp 1757447377
transform 1 0 1743 0 1 38125
box -586 -1075 12571 1441
use fuse  fuse_8
timestamp 1757447377
transform 1 0 1743 0 1 40925
box -586 -1075 12571 1441
use fuse  fuse_9
timestamp 1757447377
transform 1 0 1743 0 1 43725
box -586 -1075 12571 1441
use fuse  fuse_10
timestamp 1757447377
transform 1 0 1743 0 1 46525
box -586 -1075 12571 1441
use fuse  fuse_11
timestamp 1757447377
transform 1 0 1743 0 1 49325
box -586 -1075 12571 1441
use fuse  fuse_12
timestamp 1757447377
transform 1 0 1743 0 1 52125
box -586 -1075 12571 1441
use fuse  fuse_13
timestamp 1757447377
transform 1 0 1743 0 1 54925
box -586 -1075 12571 1441
use fuse  fuse_14
timestamp 1757447377
transform 1 0 1743 0 1 57725
box -586 -1075 12571 1441
use fuse  fuse_15
timestamp 1757447377
transform 1 0 1743 0 1 60525
box -586 -1075 12571 1441
use ldo  ldo_0 ../ip/ldo/magic
timestamp 1749474908
transform 0 1 30839 1 0 552
box 0 -1 29931 17112
use levelup  levelup_0 ../ip/util/magic
timestamp 1752511086
transform 0 1 17510 -1 0 18891
box -868 -1043 1370 2172
use levelup  levelup_1
timestamp 1752511086
transform 0 1 17510 -1 0 21691
box -868 -1043 1370 2172
use levelup  levelup_2
timestamp 1752511086
transform 0 1 17510 -1 0 24491
box -868 -1043 1370 2172
use levelup  levelup_3
timestamp 1752511086
transform 0 1 17510 -1 0 27291
box -868 -1043 1370 2172
use levelup  levelup_4
timestamp 1752511086
transform 0 1 17510 -1 0 30091
box -868 -1043 1370 2172
use levelup  levelup_5
timestamp 1752511086
transform 0 1 17510 -1 0 32891
box -868 -1043 1370 2172
use levelup  levelup_6
timestamp 1752511086
transform 0 1 17510 -1 0 35691
box -868 -1043 1370 2172
use levelup  levelup_7
timestamp 1752511086
transform 0 1 17510 -1 0 38491
box -868 -1043 1370 2172
use levelup  levelup_8
timestamp 1752511086
transform 0 1 17510 -1 0 41291
box -868 -1043 1370 2172
use levelup  levelup_9
timestamp 1752511086
transform 0 1 17510 -1 0 44091
box -868 -1043 1370 2172
use levelup  levelup_10
timestamp 1752511086
transform 0 1 17510 -1 0 46891
box -868 -1043 1370 2172
use levelup  levelup_11
timestamp 1752511086
transform 0 1 17510 -1 0 49691
box -868 -1043 1370 2172
use levelup  levelup_12
timestamp 1752511086
transform 0 1 17510 -1 0 52491
box -868 -1043 1370 2172
use levelup  levelup_13
timestamp 1752511086
transform 0 1 17510 -1 0 55291
box -868 -1043 1370 2172
use levelup  levelup_14
timestamp 1752511086
transform 0 1 17510 -1 0 58091
box -868 -1043 1370 2172
use levelup  levelup_15
timestamp 1752511086
transform 0 1 17510 -1 0 60891
box -868 -1043 1370 2172
use por  por_0 ../ip/por/magic
timestamp 1757240632
transform 0 -1 60088 1 0 52673
box -9582 -10167 9253 801
use powersw  powersw_0 ../ip/util/magic
timestamp 1753301161
transform -1 0 9367 0 1 189
box -977 -713 10525 12692
use riosc  riosc_0 ../ip/riosc/magic
timestamp 1757364080
transform 0 -1 74685 1 0 57174
box -4492 -1414 4631 2905
use spi  spi_0 ../ip/spi/magic
timestamp 1757240632
transform 1 0 50857 0 1 -988
box 60 480 25380 25446
use vthref  vthref_0 ../ip/vthref/magic
timestamp 1757240632
transform 0 -1 41215 -1 0 60017
box -1948 -17053 17940 14105
use vthref_source  vthref_source_0 ../ip/vthref/magic
timestamp 1757240632
transform 0 -1 41215 -1 0 56015
box 13299 -637 17939 14105
use vthref_source  vthref_source_1
timestamp 1757240632
transform 0 -1 41215 -1 0 52017
box 13299 -637 17939 14105
<< labels >>
flabel metal1 80237 51741 81037 52141 0 FreeSans 1600 0 0 0 RESET
port 11 nsew
flabel metal1 80237 51041 81037 51441 0 FreeSans 1600 0 0 0 POR
port 13 nsew
flabel metal2 48470 -5827 50637 -5027 0 FreeSans 1600 0 0 0 VLDO
port 21 nsew
flabel metal1 10344 -5827 11144 -5027 0 FreeSans 1600 0 0 0 FTOP
port 23 nsew
flabel metal1 -1884 -5827 -1484 -5027 0 FreeSans 1600 0 0 0 FPROG
port 25 nsew
flabel metal2 81212 36733 81612 37133 0 FreeSans 1600 0 0 0 CS
port 14 nsew
flabel metal2 81212 35722 81612 36122 0 FreeSans 1600 0 0 0 SCLK
port 15 nsew
flabel metal2 81212 34725 81612 35125 0 FreeSans 1600 0 0 0 DIN
port 16 nsew
flabel metal2 81212 33723 81612 34123 0 FreeSans 1600 0 0 0 DOUT
port 17 nsew
flabel metal2 81212 32712 81612 33112 0 FreeSans 1600 0 0 0 DOUT_EN
port 19 nsew
flabel metal5 56769 66359 57769 68359 0 FreeSans 1600 0 0 0 DVDD
port 27 nsew
flabel metal3 -7353 -2027 -5353 -1027 0 FreeSans 1600 0 0 0 AVDD
port 33 nsew
flabel metal4 -7353 18004 -5353 19004 0 FreeSans 1600 0 0 0 VSS
port 31 nsew
flabel metal6 36394 66359 37394 68359 0 FreeSans 1600 0 0 0 VSS
port 29 nsew
flabel metal2 75508 66359 75908 67159 0 FreeSans 1600 0 0 0 OSC
port 9 nsew
<< end >>
