magic
tech ihp-sg13g2
timestamp 1757240632
<< error_p >>
rect -33 1622 -28 1627
rect 28 1622 33 1627
rect -38 1617 -33 1622
rect 33 1617 38 1622
rect -38 1606 -33 1611
rect 33 1606 38 1611
rect -33 1601 -28 1606
rect 28 1601 33 1606
rect -67 1585 -62 1590
rect -56 1585 -51 1590
rect 51 1585 56 1590
rect 62 1585 67 1590
rect -72 1580 -67 1585
rect -51 1580 -46 1585
rect 46 1580 51 1585
rect 67 1580 72 1585
rect -72 599 -67 604
rect -51 599 -46 604
rect 46 599 51 604
rect 67 599 72 604
rect -67 594 -62 599
rect -56 594 -51 599
rect 51 594 56 599
rect 62 594 67 599
rect -33 578 -28 583
rect 28 578 33 583
rect -38 573 -33 578
rect 33 573 38 578
rect -38 562 -33 567
rect 33 562 38 567
rect -33 557 -28 562
rect 28 557 33 562
rect -33 530 -28 535
rect 28 530 33 535
rect -38 525 -33 530
rect 33 525 38 530
rect -38 514 -33 519
rect 33 514 38 519
rect -33 509 -28 514
rect 28 509 33 514
rect -67 493 -62 498
rect -56 493 -51 498
rect 51 493 56 498
rect 62 493 67 498
rect -72 488 -67 493
rect -51 488 -46 493
rect 46 488 51 493
rect 67 488 72 493
rect -72 -493 -67 -488
rect -51 -493 -46 -488
rect 46 -493 51 -488
rect 67 -493 72 -488
rect -67 -498 -62 -493
rect -56 -498 -51 -493
rect 51 -498 56 -493
rect 62 -498 67 -493
rect -33 -514 -28 -509
rect 28 -514 33 -509
rect -38 -519 -33 -514
rect 33 -519 38 -514
rect -38 -530 -33 -525
rect 33 -530 38 -525
rect -33 -535 -28 -530
rect 28 -535 33 -530
<< hvnmos >>
rect -40 592 40 1592
rect -40 -500 40 500
<< hvndiff >>
rect -74 1585 -40 1592
rect -74 599 -67 1585
rect -51 599 -40 1585
rect -74 592 -40 599
rect 40 1585 74 1592
rect 40 599 51 1585
rect 67 599 74 1585
rect 40 592 74 599
rect -74 493 -40 500
rect -74 -493 -67 493
rect -51 -493 -40 493
rect -74 -500 -40 -493
rect 40 493 74 500
rect 40 -493 51 493
rect 67 -493 74 493
rect 40 -500 74 -493
<< hvndiffc >>
rect -67 599 -51 1585
rect 51 599 67 1585
rect -67 -493 -51 493
rect 51 -493 67 493
<< psubdiff >>
rect -185 1622 -155 1629
rect -185 -563 -178 1622
rect -162 -563 -155 1622
rect 155 1622 185 1629
rect -185 -570 -155 -563
rect 155 -563 162 1622
rect 178 -563 185 1622
rect 155 -570 185 -563
rect -185 -577 185 -570
rect -185 -593 -148 -577
rect 148 -593 185 -577
rect -185 -600 185 -593
<< psubdiffcont >>
rect -178 -563 -162 1622
rect 162 -563 178 1622
rect -148 -593 148 -577
<< poly >>
rect -40 1622 40 1629
rect -40 1606 -33 1622
rect 33 1606 40 1622
rect -40 1592 40 1606
rect -40 578 40 592
rect -40 562 -33 578
rect 33 562 40 578
rect -40 555 40 562
rect -40 530 40 537
rect -40 514 -33 530
rect 33 514 40 530
rect -40 500 40 514
rect -40 -514 40 -500
rect -40 -530 -33 -514
rect 33 -530 40 -514
rect -40 -537 40 -530
<< polycont >>
rect -33 1606 33 1622
rect -33 562 33 578
rect -33 514 33 530
rect -33 -530 33 -514
<< metal1 >>
rect -183 1622 -157 1627
rect 157 1622 183 1627
rect -183 -563 -178 1622
rect -162 -563 -157 1622
rect -183 -572 -157 -563
rect 157 -563 162 1622
rect 178 -563 183 1622
rect 157 -572 183 -563
rect -183 -577 183 -572
rect -183 -593 -148 -577
rect 148 -593 183 -577
rect -183 -598 183 -593
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 10 l 0.8 nf 1 nx 1 dx 0.21 ny 2 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 0 gbc 1
<< end >>
