magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2000 18124 37600
<< isosubstrate >>
rect 0 23124 16000 28034
<< nwell >>
rect -124 33246 16124 33554
rect -124 29546 16124 29854
rect -124 12516 16124 12832
rect -124 6276 192 12516
rect 15808 6276 16124 12516
rect -124 5960 16124 6276
rect -124 1076 154 5960
rect 15846 1076 16124 5960
<< pwell >>
rect -26 31344 16026 31456
rect -26 23098 16026 28060
rect -26 12974 94 23098
rect 15908 12974 16026 23098
<< psubdiff >>
rect 118 31384 150 31416
rect 186 31384 218 31416
rect 254 31384 286 31416
rect 322 31384 354 31416
rect 390 31384 422 31416
rect 458 31384 490 31416
rect 526 31384 558 31416
rect 594 31384 626 31416
rect 662 31384 694 31416
rect 730 31384 762 31416
rect 798 31384 830 31416
rect 866 31384 898 31416
rect 934 31384 966 31416
rect 1002 31384 1034 31416
rect 1070 31384 1102 31416
rect 1138 31384 1170 31416
rect 1206 31384 1238 31416
rect 1274 31384 1306 31416
rect 1342 31384 1374 31416
rect 1410 31384 1442 31416
rect 1478 31384 1510 31416
rect 1546 31384 1578 31416
rect 1614 31384 1646 31416
rect 1682 31384 1714 31416
rect 1750 31384 1782 31416
rect 1818 31384 1850 31416
rect 1886 31384 1918 31416
rect 1954 31384 1986 31416
rect 2022 31384 2054 31416
rect 2090 31384 2122 31416
rect 2158 31384 2190 31416
rect 2226 31384 2258 31416
rect 2294 31384 2326 31416
rect 2362 31384 2394 31416
rect 2430 31384 2462 31416
rect 2498 31384 2530 31416
rect 2566 31384 2598 31416
rect 2634 31384 2666 31416
rect 2702 31384 2734 31416
rect 2770 31384 2802 31416
rect 2838 31384 2870 31416
rect 2906 31384 2938 31416
rect 2974 31384 3006 31416
rect 3042 31384 3074 31416
rect 3110 31384 3142 31416
rect 3178 31384 3210 31416
rect 3246 31384 3278 31416
rect 3314 31384 3346 31416
rect 3382 31384 3414 31416
rect 3450 31384 3482 31416
rect 3518 31384 3550 31416
rect 3586 31384 3618 31416
rect 3654 31384 3686 31416
rect 3722 31384 3754 31416
rect 3790 31384 3822 31416
rect 3858 31384 3890 31416
rect 3926 31384 3958 31416
rect 3994 31384 4026 31416
rect 4062 31384 4094 31416
rect 4130 31384 4162 31416
rect 4198 31384 4230 31416
rect 4266 31384 4298 31416
rect 4334 31384 4366 31416
rect 4402 31384 4434 31416
rect 4470 31384 4502 31416
rect 4538 31384 4570 31416
rect 4606 31384 4638 31416
rect 4674 31384 4706 31416
rect 4742 31384 4774 31416
rect 4810 31384 4842 31416
rect 4878 31384 4910 31416
rect 4946 31384 4978 31416
rect 5014 31384 5046 31416
rect 5082 31384 5114 31416
rect 5150 31384 5182 31416
rect 5218 31384 5250 31416
rect 5286 31384 5318 31416
rect 5354 31384 5386 31416
rect 5422 31384 5454 31416
rect 5490 31384 5522 31416
rect 5558 31384 5590 31416
rect 5626 31384 5658 31416
rect 5694 31384 5726 31416
rect 5762 31384 5794 31416
rect 5830 31384 5862 31416
rect 5898 31384 5930 31416
rect 5966 31384 5998 31416
rect 6034 31384 6066 31416
rect 6102 31384 6134 31416
rect 6170 31384 6202 31416
rect 6238 31384 6270 31416
rect 6306 31384 6338 31416
rect 6374 31384 6406 31416
rect 6442 31384 6474 31416
rect 6510 31384 6542 31416
rect 6578 31384 6610 31416
rect 6646 31384 6678 31416
rect 6714 31384 6746 31416
rect 6782 31384 6814 31416
rect 6850 31384 6882 31416
rect 6918 31384 6950 31416
rect 6986 31384 7018 31416
rect 7054 31384 7086 31416
rect 7122 31384 7154 31416
rect 7190 31384 7222 31416
rect 7258 31384 7290 31416
rect 7326 31384 7358 31416
rect 7394 31384 7426 31416
rect 7462 31384 7494 31416
rect 7530 31384 7562 31416
rect 7598 31384 7630 31416
rect 7666 31384 7698 31416
rect 7734 31384 7766 31416
rect 7802 31384 7834 31416
rect 7870 31384 7902 31416
rect 7938 31384 7970 31416
rect 8006 31384 8038 31416
rect 8074 31384 8106 31416
rect 8142 31384 8174 31416
rect 8210 31384 8242 31416
rect 8278 31384 8310 31416
rect 8346 31384 8378 31416
rect 8414 31384 8446 31416
rect 8482 31384 8514 31416
rect 8550 31384 8582 31416
rect 8618 31384 8650 31416
rect 8686 31384 8718 31416
rect 8754 31384 8786 31416
rect 8822 31384 8854 31416
rect 8890 31384 8922 31416
rect 8958 31384 8990 31416
rect 9026 31384 9058 31416
rect 9094 31384 9126 31416
rect 9162 31384 9194 31416
rect 9230 31384 9262 31416
rect 9298 31384 9330 31416
rect 9366 31384 9398 31416
rect 9434 31384 9466 31416
rect 9502 31384 9534 31416
rect 9570 31384 9602 31416
rect 9638 31384 9670 31416
rect 9706 31384 9738 31416
rect 9774 31384 9806 31416
rect 9842 31384 9874 31416
rect 9910 31384 9942 31416
rect 9978 31384 10010 31416
rect 10046 31384 10078 31416
rect 10114 31384 10146 31416
rect 10182 31384 10214 31416
rect 10250 31384 10282 31416
rect 10318 31384 10350 31416
rect 10386 31384 10418 31416
rect 10454 31384 10486 31416
rect 10522 31384 10554 31416
rect 10590 31384 10622 31416
rect 10658 31384 10690 31416
rect 10726 31384 10758 31416
rect 10794 31384 10826 31416
rect 10862 31384 10894 31416
rect 10930 31384 10962 31416
rect 10998 31384 11030 31416
rect 11066 31384 11098 31416
rect 11134 31384 11166 31416
rect 11202 31384 11234 31416
rect 11270 31384 11302 31416
rect 11338 31384 11370 31416
rect 11406 31384 11438 31416
rect 11474 31384 11506 31416
rect 11542 31384 11574 31416
rect 11610 31384 11642 31416
rect 11678 31384 11710 31416
rect 11746 31384 11778 31416
rect 11814 31384 11846 31416
rect 11882 31384 11914 31416
rect 11950 31384 11982 31416
rect 12018 31384 12050 31416
rect 12086 31384 12118 31416
rect 12154 31384 12186 31416
rect 12222 31384 12254 31416
rect 12290 31384 12322 31416
rect 12358 31384 12390 31416
rect 12426 31384 12458 31416
rect 12494 31384 12526 31416
rect 12562 31384 12594 31416
rect 12630 31384 12662 31416
rect 12698 31384 12730 31416
rect 12766 31384 12798 31416
rect 12834 31384 12866 31416
rect 12902 31384 12934 31416
rect 12970 31384 13002 31416
rect 13038 31384 13070 31416
rect 13106 31384 13138 31416
rect 13174 31384 13206 31416
rect 13242 31384 13274 31416
rect 13310 31384 13342 31416
rect 13378 31384 13410 31416
rect 13446 31384 13478 31416
rect 13514 31384 13546 31416
rect 13582 31384 13614 31416
rect 13650 31384 13682 31416
rect 13718 31384 13750 31416
rect 13786 31384 13818 31416
rect 13854 31384 13886 31416
rect 13922 31384 13954 31416
rect 13990 31384 14022 31416
rect 14058 31384 14090 31416
rect 14126 31384 14158 31416
rect 14194 31384 14226 31416
rect 14262 31384 14294 31416
rect 14330 31384 14362 31416
rect 14398 31384 14430 31416
rect 14466 31384 14498 31416
rect 14534 31384 14566 31416
rect 14602 31384 14634 31416
rect 14670 31384 14702 31416
rect 14738 31384 14770 31416
rect 14806 31384 14838 31416
rect 14874 31384 14906 31416
rect 14942 31384 14974 31416
rect 15010 31384 15042 31416
rect 15078 31384 15110 31416
rect 15146 31384 15178 31416
rect 15214 31384 15246 31416
rect 15282 31384 15314 31416
rect 15350 31384 15382 31416
rect 15442 31384 15474 31416
rect 15510 31384 15542 31416
rect 15578 31384 15610 31416
rect 15646 31384 15678 31416
rect 15714 31384 15746 31416
rect 15782 31384 15814 31416
rect 15850 31384 15882 31416
rect 15918 31384 15950 31416
rect 136 27939 168 27971
rect 208 27939 240 27971
rect 280 27939 312 27971
rect 352 27939 384 27971
rect 424 27939 456 27971
rect 496 27939 528 27971
rect 568 27939 600 27971
rect 640 27939 672 27971
rect 712 27939 744 27971
rect 784 27939 816 27971
rect 856 27939 888 27971
rect 928 27939 960 27971
rect 1000 27939 1032 27971
rect 1072 27939 1104 27971
rect 1144 27939 1176 27971
rect 1216 27939 1248 27971
rect 1288 27939 1320 27971
rect 1360 27939 1392 27971
rect 1432 27939 1464 27971
rect 1504 27939 1536 27971
rect 1576 27939 1608 27971
rect 1648 27939 1680 27971
rect 1720 27939 1752 27971
rect 1792 27939 1824 27971
rect 1864 27939 1896 27971
rect 1936 27939 1968 27971
rect 2008 27939 2040 27971
rect 2080 27939 2112 27971
rect 2152 27939 2184 27971
rect 2224 27939 2256 27971
rect 2296 27939 2328 27971
rect 2368 27939 2400 27971
rect 2440 27939 2472 27971
rect 2512 27939 2544 27971
rect 2584 27939 2616 27971
rect 2656 27939 2688 27971
rect 2728 27939 2760 27971
rect 2800 27939 2832 27971
rect 2872 27939 2904 27971
rect 2944 27939 2976 27971
rect 3016 27939 3048 27971
rect 3088 27939 3120 27971
rect 3160 27939 3192 27971
rect 3232 27939 3264 27971
rect 3304 27939 3336 27971
rect 3376 27939 3408 27971
rect 3448 27939 3480 27971
rect 3520 27939 3552 27971
rect 3592 27939 3624 27971
rect 3664 27939 3696 27971
rect 3736 27939 3768 27971
rect 3808 27939 3840 27971
rect 3880 27939 3912 27971
rect 3952 27939 3984 27971
rect 4024 27939 4056 27971
rect 4096 27939 4128 27971
rect 4168 27939 4200 27971
rect 4240 27939 4272 27971
rect 4312 27939 4344 27971
rect 4384 27939 4416 27971
rect 4456 27939 4488 27971
rect 4528 27939 4560 27971
rect 4600 27939 4632 27971
rect 4672 27939 4704 27971
rect 4744 27939 4776 27971
rect 4816 27939 4848 27971
rect 4888 27939 4920 27971
rect 4960 27939 4992 27971
rect 5032 27939 5064 27971
rect 5104 27939 5136 27971
rect 5176 27939 5208 27971
rect 5248 27939 5280 27971
rect 5320 27939 5352 27971
rect 5392 27939 5424 27971
rect 5464 27939 5496 27971
rect 5536 27939 5568 27971
rect 5608 27939 5640 27971
rect 5680 27939 5712 27971
rect 5752 27939 5784 27971
rect 5824 27939 5856 27971
rect 5896 27939 5928 27971
rect 5968 27939 6000 27971
rect 6040 27939 6072 27971
rect 6112 27939 6144 27971
rect 6184 27939 6216 27971
rect 6256 27939 6288 27971
rect 6328 27939 6360 27971
rect 6400 27939 6432 27971
rect 6472 27939 6504 27971
rect 6544 27939 6576 27971
rect 6616 27939 6648 27971
rect 6688 27939 6720 27971
rect 6760 27939 6792 27971
rect 6832 27939 6864 27971
rect 6904 27939 6936 27971
rect 6976 27939 7008 27971
rect 7048 27939 7080 27971
rect 7120 27939 7152 27971
rect 7192 27939 7224 27971
rect 7264 27939 7296 27971
rect 7336 27939 7368 27971
rect 7408 27939 7440 27971
rect 7480 27939 7512 27971
rect 7552 27939 7584 27971
rect 7624 27939 7656 27971
rect 7696 27939 7728 27971
rect 7768 27939 7800 27971
rect 7840 27939 7872 27971
rect 7912 27939 7944 27971
rect 7984 27939 8016 27971
rect 8056 27939 8088 27971
rect 8128 27939 8160 27971
rect 8200 27939 8232 27971
rect 8272 27939 8304 27971
rect 8344 27939 8376 27971
rect 8416 27939 8448 27971
rect 8488 27939 8520 27971
rect 8560 27939 8592 27971
rect 8632 27939 8664 27971
rect 8704 27939 8736 27971
rect 8776 27939 8808 27971
rect 8848 27939 8880 27971
rect 8920 27939 8952 27971
rect 8992 27939 9024 27971
rect 9064 27939 9096 27971
rect 9136 27939 9168 27971
rect 9208 27939 9240 27971
rect 9280 27939 9312 27971
rect 9352 27939 9384 27971
rect 9424 27939 9456 27971
rect 9496 27939 9528 27971
rect 9568 27939 9600 27971
rect 9640 27939 9672 27971
rect 9712 27939 9744 27971
rect 9784 27939 9816 27971
rect 9856 27939 9888 27971
rect 9928 27939 9960 27971
rect 10000 27939 10032 27971
rect 10072 27939 10104 27971
rect 10144 27939 10176 27971
rect 10216 27939 10248 27971
rect 10288 27939 10320 27971
rect 10360 27939 10392 27971
rect 10432 27939 10464 27971
rect 10504 27939 10536 27971
rect 10576 27939 10608 27971
rect 10648 27939 10680 27971
rect 10720 27939 10752 27971
rect 10792 27939 10824 27971
rect 10864 27939 10896 27971
rect 10936 27939 10968 27971
rect 11008 27939 11040 27971
rect 11080 27939 11112 27971
rect 11152 27939 11184 27971
rect 11224 27939 11256 27971
rect 11296 27939 11328 27971
rect 11368 27939 11400 27971
rect 11440 27939 11472 27971
rect 11512 27939 11544 27971
rect 11584 27939 11616 27971
rect 11656 27939 11688 27971
rect 11728 27939 11760 27971
rect 11800 27939 11832 27971
rect 11872 27939 11904 27971
rect 11944 27939 11976 27971
rect 12016 27939 12048 27971
rect 12088 27939 12120 27971
rect 12160 27939 12192 27971
rect 12232 27939 12264 27971
rect 12304 27939 12336 27971
rect 12376 27939 12408 27971
rect 12448 27939 12480 27971
rect 12520 27939 12552 27971
rect 12592 27939 12624 27971
rect 12664 27939 12696 27971
rect 12736 27939 12768 27971
rect 12808 27939 12840 27971
rect 12880 27939 12912 27971
rect 12952 27939 12984 27971
rect 13024 27939 13056 27971
rect 13096 27939 13128 27971
rect 13168 27939 13200 27971
rect 13240 27939 13272 27971
rect 13312 27939 13344 27971
rect 13384 27939 13416 27971
rect 13456 27939 13488 27971
rect 13528 27939 13560 27971
rect 13600 27939 13632 27971
rect 13672 27939 13704 27971
rect 13744 27939 13776 27971
rect 13816 27939 13848 27971
rect 13888 27939 13920 27971
rect 13960 27939 13992 27971
rect 14032 27939 14064 27971
rect 14104 27939 14136 27971
rect 14176 27939 14208 27971
rect 14248 27939 14280 27971
rect 14320 27939 14352 27971
rect 14392 27939 14424 27971
rect 14464 27939 14496 27971
rect 14536 27939 14568 27971
rect 14608 27939 14640 27971
rect 14680 27939 14712 27971
rect 14752 27939 14784 27971
rect 14824 27939 14856 27971
rect 14896 27939 14928 27971
rect 14968 27939 15000 27971
rect 15040 27939 15072 27971
rect 15112 27939 15144 27971
rect 15184 27939 15216 27971
rect 15256 27939 15288 27971
rect 15328 27939 15360 27971
rect 15400 27939 15432 27971
rect 15472 27939 15504 27971
rect 15544 27939 15576 27971
rect 15616 27939 15648 27971
rect 15688 27939 15720 27971
rect 15760 27939 15792 27971
rect 15832 27939 15864 27971
rect 15904 27939 15936 27971
rect 64 27867 96 27899
rect 136 27867 168 27899
rect 208 27867 240 27899
rect 280 27867 312 27899
rect 352 27867 384 27899
rect 424 27867 456 27899
rect 496 27867 528 27899
rect 568 27867 600 27899
rect 640 27867 672 27899
rect 712 27867 744 27899
rect 784 27867 816 27899
rect 856 27867 888 27899
rect 928 27867 960 27899
rect 1000 27867 1032 27899
rect 1072 27867 1104 27899
rect 1144 27867 1176 27899
rect 1216 27867 1248 27899
rect 1288 27867 1320 27899
rect 1360 27867 1392 27899
rect 1432 27867 1464 27899
rect 1504 27867 1536 27899
rect 1576 27867 1608 27899
rect 1648 27867 1680 27899
rect 1720 27867 1752 27899
rect 1792 27867 1824 27899
rect 1864 27867 1896 27899
rect 1936 27867 1968 27899
rect 2008 27867 2040 27899
rect 2080 27867 2112 27899
rect 2152 27867 2184 27899
rect 2224 27867 2256 27899
rect 2296 27867 2328 27899
rect 2368 27867 2400 27899
rect 2440 27867 2472 27899
rect 2512 27867 2544 27899
rect 2584 27867 2616 27899
rect 2656 27867 2688 27899
rect 2728 27867 2760 27899
rect 2800 27867 2832 27899
rect 2872 27867 2904 27899
rect 2944 27867 2976 27899
rect 3016 27867 3048 27899
rect 3088 27867 3120 27899
rect 3160 27867 3192 27899
rect 3232 27867 3264 27899
rect 3304 27867 3336 27899
rect 3376 27867 3408 27899
rect 3448 27867 3480 27899
rect 3520 27867 3552 27899
rect 3592 27867 3624 27899
rect 3664 27867 3696 27899
rect 3736 27867 3768 27899
rect 3808 27867 3840 27899
rect 3880 27867 3912 27899
rect 3952 27867 3984 27899
rect 4024 27867 4056 27899
rect 4096 27867 4128 27899
rect 4168 27867 4200 27899
rect 4240 27867 4272 27899
rect 4312 27867 4344 27899
rect 4384 27867 4416 27899
rect 4456 27867 4488 27899
rect 4528 27867 4560 27899
rect 4600 27867 4632 27899
rect 4672 27867 4704 27899
rect 4744 27867 4776 27899
rect 4816 27867 4848 27899
rect 4888 27867 4920 27899
rect 4960 27867 4992 27899
rect 5032 27867 5064 27899
rect 5104 27867 5136 27899
rect 5176 27867 5208 27899
rect 5248 27867 5280 27899
rect 5320 27867 5352 27899
rect 5392 27867 5424 27899
rect 5464 27867 5496 27899
rect 5536 27867 5568 27899
rect 5608 27867 5640 27899
rect 5680 27867 5712 27899
rect 5752 27867 5784 27899
rect 5824 27867 5856 27899
rect 5896 27867 5928 27899
rect 5968 27867 6000 27899
rect 6040 27867 6072 27899
rect 6112 27867 6144 27899
rect 6184 27867 6216 27899
rect 6256 27867 6288 27899
rect 6328 27867 6360 27899
rect 6400 27867 6432 27899
rect 6472 27867 6504 27899
rect 6544 27867 6576 27899
rect 6616 27867 6648 27899
rect 6688 27867 6720 27899
rect 6760 27867 6792 27899
rect 6832 27867 6864 27899
rect 6904 27867 6936 27899
rect 6976 27867 7008 27899
rect 7048 27867 7080 27899
rect 7120 27867 7152 27899
rect 7192 27867 7224 27899
rect 7264 27867 7296 27899
rect 7336 27867 7368 27899
rect 7408 27867 7440 27899
rect 7480 27867 7512 27899
rect 7552 27867 7584 27899
rect 7624 27867 7656 27899
rect 7696 27867 7728 27899
rect 7768 27867 7800 27899
rect 7840 27867 7872 27899
rect 7912 27867 7944 27899
rect 7984 27867 8016 27899
rect 8056 27867 8088 27899
rect 8128 27867 8160 27899
rect 8200 27867 8232 27899
rect 8272 27867 8304 27899
rect 8344 27867 8376 27899
rect 8416 27867 8448 27899
rect 8488 27867 8520 27899
rect 8560 27867 8592 27899
rect 8632 27867 8664 27899
rect 8704 27867 8736 27899
rect 8776 27867 8808 27899
rect 8848 27867 8880 27899
rect 8920 27867 8952 27899
rect 8992 27867 9024 27899
rect 9064 27867 9096 27899
rect 9136 27867 9168 27899
rect 9208 27867 9240 27899
rect 9280 27867 9312 27899
rect 9352 27867 9384 27899
rect 9424 27867 9456 27899
rect 9496 27867 9528 27899
rect 9568 27867 9600 27899
rect 9640 27867 9672 27899
rect 9712 27867 9744 27899
rect 9784 27867 9816 27899
rect 9856 27867 9888 27899
rect 9928 27867 9960 27899
rect 10000 27867 10032 27899
rect 10072 27867 10104 27899
rect 10144 27867 10176 27899
rect 10216 27867 10248 27899
rect 10288 27867 10320 27899
rect 10360 27867 10392 27899
rect 10432 27867 10464 27899
rect 10504 27867 10536 27899
rect 10576 27867 10608 27899
rect 10648 27867 10680 27899
rect 10720 27867 10752 27899
rect 10792 27867 10824 27899
rect 10864 27867 10896 27899
rect 10936 27867 10968 27899
rect 11008 27867 11040 27899
rect 11080 27867 11112 27899
rect 11152 27867 11184 27899
rect 11224 27867 11256 27899
rect 11296 27867 11328 27899
rect 11368 27867 11400 27899
rect 11440 27867 11472 27899
rect 11512 27867 11544 27899
rect 11584 27867 11616 27899
rect 11656 27867 11688 27899
rect 11728 27867 11760 27899
rect 11800 27867 11832 27899
rect 11872 27867 11904 27899
rect 11944 27867 11976 27899
rect 12016 27867 12048 27899
rect 12088 27867 12120 27899
rect 12160 27867 12192 27899
rect 12232 27867 12264 27899
rect 12304 27867 12336 27899
rect 12376 27867 12408 27899
rect 12448 27867 12480 27899
rect 12520 27867 12552 27899
rect 12592 27867 12624 27899
rect 12664 27867 12696 27899
rect 12736 27867 12768 27899
rect 12808 27867 12840 27899
rect 12880 27867 12912 27899
rect 12952 27867 12984 27899
rect 13024 27867 13056 27899
rect 13096 27867 13128 27899
rect 13168 27867 13200 27899
rect 13240 27867 13272 27899
rect 13312 27867 13344 27899
rect 13384 27867 13416 27899
rect 13456 27867 13488 27899
rect 13528 27867 13560 27899
rect 13600 27867 13632 27899
rect 13672 27867 13704 27899
rect 13744 27867 13776 27899
rect 13816 27867 13848 27899
rect 13888 27867 13920 27899
rect 13960 27867 13992 27899
rect 14032 27867 14064 27899
rect 14104 27867 14136 27899
rect 14176 27867 14208 27899
rect 14248 27867 14280 27899
rect 14320 27867 14352 27899
rect 14392 27867 14424 27899
rect 14464 27867 14496 27899
rect 14536 27867 14568 27899
rect 14608 27867 14640 27899
rect 14680 27867 14712 27899
rect 14752 27867 14784 27899
rect 14824 27867 14856 27899
rect 14896 27867 14928 27899
rect 14968 27867 15000 27899
rect 15040 27867 15072 27899
rect 15112 27867 15144 27899
rect 15184 27867 15216 27899
rect 15256 27867 15288 27899
rect 15328 27867 15360 27899
rect 15400 27867 15432 27899
rect 15472 27867 15504 27899
rect 15544 27867 15576 27899
rect 15616 27867 15648 27899
rect 15688 27867 15720 27899
rect 15760 27867 15792 27899
rect 15832 27867 15864 27899
rect 15904 27867 15936 27899
rect 64 27795 96 27827
rect 136 27795 168 27827
rect 208 27795 240 27827
rect 280 27795 312 27827
rect 352 27795 384 27827
rect 424 27795 456 27827
rect 496 27795 528 27827
rect 568 27795 600 27827
rect 640 27795 672 27827
rect 712 27795 744 27827
rect 784 27795 816 27827
rect 856 27795 888 27827
rect 928 27795 960 27827
rect 1000 27795 1032 27827
rect 1072 27795 1104 27827
rect 1144 27795 1176 27827
rect 1216 27795 1248 27827
rect 1288 27795 1320 27827
rect 1360 27795 1392 27827
rect 1432 27795 1464 27827
rect 1504 27795 1536 27827
rect 1576 27795 1608 27827
rect 1648 27795 1680 27827
rect 1720 27795 1752 27827
rect 1792 27795 1824 27827
rect 1864 27795 1896 27827
rect 1936 27795 1968 27827
rect 2008 27795 2040 27827
rect 2080 27795 2112 27827
rect 2152 27795 2184 27827
rect 2224 27795 2256 27827
rect 2296 27795 2328 27827
rect 2368 27795 2400 27827
rect 2440 27795 2472 27827
rect 2512 27795 2544 27827
rect 2584 27795 2616 27827
rect 2656 27795 2688 27827
rect 2728 27795 2760 27827
rect 2800 27795 2832 27827
rect 2872 27795 2904 27827
rect 2944 27795 2976 27827
rect 3016 27795 3048 27827
rect 3088 27795 3120 27827
rect 3160 27795 3192 27827
rect 3232 27795 3264 27827
rect 3304 27795 3336 27827
rect 3376 27795 3408 27827
rect 3448 27795 3480 27827
rect 3520 27795 3552 27827
rect 3592 27795 3624 27827
rect 3664 27795 3696 27827
rect 3736 27795 3768 27827
rect 3808 27795 3840 27827
rect 3880 27795 3912 27827
rect 3952 27795 3984 27827
rect 4024 27795 4056 27827
rect 4096 27795 4128 27827
rect 4168 27795 4200 27827
rect 4240 27795 4272 27827
rect 4312 27795 4344 27827
rect 4384 27795 4416 27827
rect 4456 27795 4488 27827
rect 4528 27795 4560 27827
rect 4600 27795 4632 27827
rect 4672 27795 4704 27827
rect 4744 27795 4776 27827
rect 4816 27795 4848 27827
rect 4888 27795 4920 27827
rect 4960 27795 4992 27827
rect 5032 27795 5064 27827
rect 5104 27795 5136 27827
rect 5176 27795 5208 27827
rect 5248 27795 5280 27827
rect 5320 27795 5352 27827
rect 5392 27795 5424 27827
rect 5464 27795 5496 27827
rect 5536 27795 5568 27827
rect 5608 27795 5640 27827
rect 5680 27795 5712 27827
rect 5752 27795 5784 27827
rect 5824 27795 5856 27827
rect 5896 27795 5928 27827
rect 5968 27795 6000 27827
rect 6040 27795 6072 27827
rect 6112 27795 6144 27827
rect 6184 27795 6216 27827
rect 6256 27795 6288 27827
rect 6328 27795 6360 27827
rect 6400 27795 6432 27827
rect 6472 27795 6504 27827
rect 6544 27795 6576 27827
rect 6616 27795 6648 27827
rect 6688 27795 6720 27827
rect 6760 27795 6792 27827
rect 6832 27795 6864 27827
rect 6904 27795 6936 27827
rect 6976 27795 7008 27827
rect 7048 27795 7080 27827
rect 7120 27795 7152 27827
rect 7192 27795 7224 27827
rect 7264 27795 7296 27827
rect 7336 27795 7368 27827
rect 7408 27795 7440 27827
rect 7480 27795 7512 27827
rect 7552 27795 7584 27827
rect 7624 27795 7656 27827
rect 7696 27795 7728 27827
rect 7768 27795 7800 27827
rect 7840 27795 7872 27827
rect 7912 27795 7944 27827
rect 7984 27795 8016 27827
rect 8056 27795 8088 27827
rect 8128 27795 8160 27827
rect 8200 27795 8232 27827
rect 8272 27795 8304 27827
rect 8344 27795 8376 27827
rect 8416 27795 8448 27827
rect 8488 27795 8520 27827
rect 8560 27795 8592 27827
rect 8632 27795 8664 27827
rect 8704 27795 8736 27827
rect 8776 27795 8808 27827
rect 8848 27795 8880 27827
rect 8920 27795 8952 27827
rect 8992 27795 9024 27827
rect 9064 27795 9096 27827
rect 9136 27795 9168 27827
rect 9208 27795 9240 27827
rect 9280 27795 9312 27827
rect 9352 27795 9384 27827
rect 9424 27795 9456 27827
rect 9496 27795 9528 27827
rect 9568 27795 9600 27827
rect 9640 27795 9672 27827
rect 9712 27795 9744 27827
rect 9784 27795 9816 27827
rect 9856 27795 9888 27827
rect 9928 27795 9960 27827
rect 10000 27795 10032 27827
rect 10072 27795 10104 27827
rect 10144 27795 10176 27827
rect 10216 27795 10248 27827
rect 10288 27795 10320 27827
rect 10360 27795 10392 27827
rect 10432 27795 10464 27827
rect 10504 27795 10536 27827
rect 10576 27795 10608 27827
rect 10648 27795 10680 27827
rect 10720 27795 10752 27827
rect 10792 27795 10824 27827
rect 10864 27795 10896 27827
rect 10936 27795 10968 27827
rect 11008 27795 11040 27827
rect 11080 27795 11112 27827
rect 11152 27795 11184 27827
rect 11224 27795 11256 27827
rect 11296 27795 11328 27827
rect 11368 27795 11400 27827
rect 11440 27795 11472 27827
rect 11512 27795 11544 27827
rect 11584 27795 11616 27827
rect 11656 27795 11688 27827
rect 11728 27795 11760 27827
rect 11800 27795 11832 27827
rect 11872 27795 11904 27827
rect 11944 27795 11976 27827
rect 12016 27795 12048 27827
rect 12088 27795 12120 27827
rect 12160 27795 12192 27827
rect 12232 27795 12264 27827
rect 12304 27795 12336 27827
rect 12376 27795 12408 27827
rect 12448 27795 12480 27827
rect 12520 27795 12552 27827
rect 12592 27795 12624 27827
rect 12664 27795 12696 27827
rect 12736 27795 12768 27827
rect 12808 27795 12840 27827
rect 12880 27795 12912 27827
rect 12952 27795 12984 27827
rect 13024 27795 13056 27827
rect 13096 27795 13128 27827
rect 13168 27795 13200 27827
rect 13240 27795 13272 27827
rect 13312 27795 13344 27827
rect 13384 27795 13416 27827
rect 13456 27795 13488 27827
rect 13528 27795 13560 27827
rect 13600 27795 13632 27827
rect 13672 27795 13704 27827
rect 13744 27795 13776 27827
rect 13816 27795 13848 27827
rect 13888 27795 13920 27827
rect 13960 27795 13992 27827
rect 14032 27795 14064 27827
rect 14104 27795 14136 27827
rect 14176 27795 14208 27827
rect 14248 27795 14280 27827
rect 14320 27795 14352 27827
rect 14392 27795 14424 27827
rect 14464 27795 14496 27827
rect 14536 27795 14568 27827
rect 14608 27795 14640 27827
rect 14680 27795 14712 27827
rect 14752 27795 14784 27827
rect 14824 27795 14856 27827
rect 14896 27795 14928 27827
rect 14968 27795 15000 27827
rect 15040 27795 15072 27827
rect 15112 27795 15144 27827
rect 15184 27795 15216 27827
rect 15256 27795 15288 27827
rect 15328 27795 15360 27827
rect 15400 27795 15432 27827
rect 15472 27795 15504 27827
rect 15544 27795 15576 27827
rect 15616 27795 15648 27827
rect 15688 27795 15720 27827
rect 15760 27795 15792 27827
rect 15832 27795 15864 27827
rect 15904 27795 15936 27827
rect 64 27723 96 27755
rect 136 27723 168 27755
rect 208 27723 240 27755
rect 280 27723 312 27755
rect 352 27723 384 27755
rect 424 27723 456 27755
rect 496 27723 528 27755
rect 568 27723 600 27755
rect 640 27723 672 27755
rect 712 27723 744 27755
rect 784 27723 816 27755
rect 856 27723 888 27755
rect 928 27723 960 27755
rect 1000 27723 1032 27755
rect 1072 27723 1104 27755
rect 1144 27723 1176 27755
rect 1216 27723 1248 27755
rect 1288 27723 1320 27755
rect 1360 27723 1392 27755
rect 1432 27723 1464 27755
rect 1504 27723 1536 27755
rect 1576 27723 1608 27755
rect 1648 27723 1680 27755
rect 1720 27723 1752 27755
rect 1792 27723 1824 27755
rect 1864 27723 1896 27755
rect 1936 27723 1968 27755
rect 2008 27723 2040 27755
rect 2080 27723 2112 27755
rect 2152 27723 2184 27755
rect 2224 27723 2256 27755
rect 2296 27723 2328 27755
rect 2368 27723 2400 27755
rect 2440 27723 2472 27755
rect 2512 27723 2544 27755
rect 2584 27723 2616 27755
rect 2656 27723 2688 27755
rect 2728 27723 2760 27755
rect 2800 27723 2832 27755
rect 2872 27723 2904 27755
rect 2944 27723 2976 27755
rect 3016 27723 3048 27755
rect 3088 27723 3120 27755
rect 3160 27723 3192 27755
rect 3232 27723 3264 27755
rect 3304 27723 3336 27755
rect 3376 27723 3408 27755
rect 3448 27723 3480 27755
rect 3520 27723 3552 27755
rect 3592 27723 3624 27755
rect 3664 27723 3696 27755
rect 3736 27723 3768 27755
rect 3808 27723 3840 27755
rect 3880 27723 3912 27755
rect 3952 27723 3984 27755
rect 4024 27723 4056 27755
rect 4096 27723 4128 27755
rect 4168 27723 4200 27755
rect 4240 27723 4272 27755
rect 4312 27723 4344 27755
rect 4384 27723 4416 27755
rect 4456 27723 4488 27755
rect 4528 27723 4560 27755
rect 4600 27723 4632 27755
rect 4672 27723 4704 27755
rect 4744 27723 4776 27755
rect 4816 27723 4848 27755
rect 4888 27723 4920 27755
rect 4960 27723 4992 27755
rect 5032 27723 5064 27755
rect 5104 27723 5136 27755
rect 5176 27723 5208 27755
rect 5248 27723 5280 27755
rect 5320 27723 5352 27755
rect 5392 27723 5424 27755
rect 5464 27723 5496 27755
rect 5536 27723 5568 27755
rect 5608 27723 5640 27755
rect 5680 27723 5712 27755
rect 5752 27723 5784 27755
rect 5824 27723 5856 27755
rect 5896 27723 5928 27755
rect 5968 27723 6000 27755
rect 6040 27723 6072 27755
rect 6112 27723 6144 27755
rect 6184 27723 6216 27755
rect 6256 27723 6288 27755
rect 6328 27723 6360 27755
rect 6400 27723 6432 27755
rect 6472 27723 6504 27755
rect 6544 27723 6576 27755
rect 6616 27723 6648 27755
rect 6688 27723 6720 27755
rect 6760 27723 6792 27755
rect 6832 27723 6864 27755
rect 6904 27723 6936 27755
rect 6976 27723 7008 27755
rect 7048 27723 7080 27755
rect 7120 27723 7152 27755
rect 7192 27723 7224 27755
rect 7264 27723 7296 27755
rect 7336 27723 7368 27755
rect 7408 27723 7440 27755
rect 7480 27723 7512 27755
rect 7552 27723 7584 27755
rect 7624 27723 7656 27755
rect 7696 27723 7728 27755
rect 7768 27723 7800 27755
rect 7840 27723 7872 27755
rect 7912 27723 7944 27755
rect 7984 27723 8016 27755
rect 8056 27723 8088 27755
rect 8128 27723 8160 27755
rect 8200 27723 8232 27755
rect 8272 27723 8304 27755
rect 8344 27723 8376 27755
rect 8416 27723 8448 27755
rect 8488 27723 8520 27755
rect 8560 27723 8592 27755
rect 8632 27723 8664 27755
rect 8704 27723 8736 27755
rect 8776 27723 8808 27755
rect 8848 27723 8880 27755
rect 8920 27723 8952 27755
rect 8992 27723 9024 27755
rect 9064 27723 9096 27755
rect 9136 27723 9168 27755
rect 9208 27723 9240 27755
rect 9280 27723 9312 27755
rect 9352 27723 9384 27755
rect 9424 27723 9456 27755
rect 9496 27723 9528 27755
rect 9568 27723 9600 27755
rect 9640 27723 9672 27755
rect 9712 27723 9744 27755
rect 9784 27723 9816 27755
rect 9856 27723 9888 27755
rect 9928 27723 9960 27755
rect 10000 27723 10032 27755
rect 10072 27723 10104 27755
rect 10144 27723 10176 27755
rect 10216 27723 10248 27755
rect 10288 27723 10320 27755
rect 10360 27723 10392 27755
rect 10432 27723 10464 27755
rect 10504 27723 10536 27755
rect 10576 27723 10608 27755
rect 10648 27723 10680 27755
rect 10720 27723 10752 27755
rect 10792 27723 10824 27755
rect 10864 27723 10896 27755
rect 10936 27723 10968 27755
rect 11008 27723 11040 27755
rect 11080 27723 11112 27755
rect 11152 27723 11184 27755
rect 11224 27723 11256 27755
rect 11296 27723 11328 27755
rect 11368 27723 11400 27755
rect 11440 27723 11472 27755
rect 11512 27723 11544 27755
rect 11584 27723 11616 27755
rect 11656 27723 11688 27755
rect 11728 27723 11760 27755
rect 11800 27723 11832 27755
rect 11872 27723 11904 27755
rect 11944 27723 11976 27755
rect 12016 27723 12048 27755
rect 12088 27723 12120 27755
rect 12160 27723 12192 27755
rect 12232 27723 12264 27755
rect 12304 27723 12336 27755
rect 12376 27723 12408 27755
rect 12448 27723 12480 27755
rect 12520 27723 12552 27755
rect 12592 27723 12624 27755
rect 12664 27723 12696 27755
rect 12736 27723 12768 27755
rect 12808 27723 12840 27755
rect 12880 27723 12912 27755
rect 12952 27723 12984 27755
rect 13024 27723 13056 27755
rect 13096 27723 13128 27755
rect 13168 27723 13200 27755
rect 13240 27723 13272 27755
rect 13312 27723 13344 27755
rect 13384 27723 13416 27755
rect 13456 27723 13488 27755
rect 13528 27723 13560 27755
rect 13600 27723 13632 27755
rect 13672 27723 13704 27755
rect 13744 27723 13776 27755
rect 13816 27723 13848 27755
rect 13888 27723 13920 27755
rect 13960 27723 13992 27755
rect 14032 27723 14064 27755
rect 14104 27723 14136 27755
rect 14176 27723 14208 27755
rect 14248 27723 14280 27755
rect 14320 27723 14352 27755
rect 14392 27723 14424 27755
rect 14464 27723 14496 27755
rect 14536 27723 14568 27755
rect 14608 27723 14640 27755
rect 14680 27723 14712 27755
rect 14752 27723 14784 27755
rect 14824 27723 14856 27755
rect 14896 27723 14928 27755
rect 14968 27723 15000 27755
rect 15040 27723 15072 27755
rect 15112 27723 15144 27755
rect 15184 27723 15216 27755
rect 15256 27723 15288 27755
rect 15328 27723 15360 27755
rect 15400 27723 15432 27755
rect 15472 27723 15504 27755
rect 15544 27723 15576 27755
rect 15616 27723 15648 27755
rect 15688 27723 15720 27755
rect 15760 27723 15792 27755
rect 15832 27723 15864 27755
rect 15904 27723 15936 27755
rect 64 27651 96 27683
rect 136 27651 168 27683
rect 208 27651 240 27683
rect 280 27651 312 27683
rect 352 27651 384 27683
rect 424 27651 456 27683
rect 496 27651 528 27683
rect 568 27651 600 27683
rect 640 27651 672 27683
rect 712 27651 744 27683
rect 784 27651 816 27683
rect 856 27651 888 27683
rect 928 27651 960 27683
rect 1000 27651 1032 27683
rect 1072 27651 1104 27683
rect 1144 27651 1176 27683
rect 1216 27651 1248 27683
rect 1288 27651 1320 27683
rect 1360 27651 1392 27683
rect 1432 27651 1464 27683
rect 1504 27651 1536 27683
rect 1576 27651 1608 27683
rect 1648 27651 1680 27683
rect 1720 27651 1752 27683
rect 1792 27651 1824 27683
rect 1864 27651 1896 27683
rect 1936 27651 1968 27683
rect 2008 27651 2040 27683
rect 2080 27651 2112 27683
rect 2152 27651 2184 27683
rect 2224 27651 2256 27683
rect 2296 27651 2328 27683
rect 2368 27651 2400 27683
rect 2440 27651 2472 27683
rect 2512 27651 2544 27683
rect 2584 27651 2616 27683
rect 2656 27651 2688 27683
rect 2728 27651 2760 27683
rect 2800 27651 2832 27683
rect 2872 27651 2904 27683
rect 2944 27651 2976 27683
rect 3016 27651 3048 27683
rect 3088 27651 3120 27683
rect 3160 27651 3192 27683
rect 3232 27651 3264 27683
rect 3304 27651 3336 27683
rect 3376 27651 3408 27683
rect 3448 27651 3480 27683
rect 3520 27651 3552 27683
rect 3592 27651 3624 27683
rect 3664 27651 3696 27683
rect 3736 27651 3768 27683
rect 3808 27651 3840 27683
rect 3880 27651 3912 27683
rect 3952 27651 3984 27683
rect 4024 27651 4056 27683
rect 4096 27651 4128 27683
rect 4168 27651 4200 27683
rect 4240 27651 4272 27683
rect 4312 27651 4344 27683
rect 4384 27651 4416 27683
rect 4456 27651 4488 27683
rect 4528 27651 4560 27683
rect 4600 27651 4632 27683
rect 4672 27651 4704 27683
rect 4744 27651 4776 27683
rect 4816 27651 4848 27683
rect 4888 27651 4920 27683
rect 4960 27651 4992 27683
rect 5032 27651 5064 27683
rect 5104 27651 5136 27683
rect 5176 27651 5208 27683
rect 5248 27651 5280 27683
rect 5320 27651 5352 27683
rect 5392 27651 5424 27683
rect 5464 27651 5496 27683
rect 5536 27651 5568 27683
rect 5608 27651 5640 27683
rect 5680 27651 5712 27683
rect 5752 27651 5784 27683
rect 5824 27651 5856 27683
rect 5896 27651 5928 27683
rect 5968 27651 6000 27683
rect 6040 27651 6072 27683
rect 6112 27651 6144 27683
rect 6184 27651 6216 27683
rect 6256 27651 6288 27683
rect 6328 27651 6360 27683
rect 6400 27651 6432 27683
rect 6472 27651 6504 27683
rect 6544 27651 6576 27683
rect 6616 27651 6648 27683
rect 6688 27651 6720 27683
rect 6760 27651 6792 27683
rect 6832 27651 6864 27683
rect 6904 27651 6936 27683
rect 6976 27651 7008 27683
rect 7048 27651 7080 27683
rect 7120 27651 7152 27683
rect 7192 27651 7224 27683
rect 7264 27651 7296 27683
rect 7336 27651 7368 27683
rect 7408 27651 7440 27683
rect 7480 27651 7512 27683
rect 7552 27651 7584 27683
rect 7624 27651 7656 27683
rect 7696 27651 7728 27683
rect 7768 27651 7800 27683
rect 7840 27651 7872 27683
rect 7912 27651 7944 27683
rect 7984 27651 8016 27683
rect 8056 27651 8088 27683
rect 8128 27651 8160 27683
rect 8200 27651 8232 27683
rect 8272 27651 8304 27683
rect 8344 27651 8376 27683
rect 8416 27651 8448 27683
rect 8488 27651 8520 27683
rect 8560 27651 8592 27683
rect 8632 27651 8664 27683
rect 8704 27651 8736 27683
rect 8776 27651 8808 27683
rect 8848 27651 8880 27683
rect 8920 27651 8952 27683
rect 8992 27651 9024 27683
rect 9064 27651 9096 27683
rect 9136 27651 9168 27683
rect 9208 27651 9240 27683
rect 9280 27651 9312 27683
rect 9352 27651 9384 27683
rect 9424 27651 9456 27683
rect 9496 27651 9528 27683
rect 9568 27651 9600 27683
rect 9640 27651 9672 27683
rect 9712 27651 9744 27683
rect 9784 27651 9816 27683
rect 9856 27651 9888 27683
rect 9928 27651 9960 27683
rect 10000 27651 10032 27683
rect 10072 27651 10104 27683
rect 10144 27651 10176 27683
rect 10216 27651 10248 27683
rect 10288 27651 10320 27683
rect 10360 27651 10392 27683
rect 10432 27651 10464 27683
rect 10504 27651 10536 27683
rect 10576 27651 10608 27683
rect 10648 27651 10680 27683
rect 10720 27651 10752 27683
rect 10792 27651 10824 27683
rect 10864 27651 10896 27683
rect 10936 27651 10968 27683
rect 11008 27651 11040 27683
rect 11080 27651 11112 27683
rect 11152 27651 11184 27683
rect 11224 27651 11256 27683
rect 11296 27651 11328 27683
rect 11368 27651 11400 27683
rect 11440 27651 11472 27683
rect 11512 27651 11544 27683
rect 11584 27651 11616 27683
rect 11656 27651 11688 27683
rect 11728 27651 11760 27683
rect 11800 27651 11832 27683
rect 11872 27651 11904 27683
rect 11944 27651 11976 27683
rect 12016 27651 12048 27683
rect 12088 27651 12120 27683
rect 12160 27651 12192 27683
rect 12232 27651 12264 27683
rect 12304 27651 12336 27683
rect 12376 27651 12408 27683
rect 12448 27651 12480 27683
rect 12520 27651 12552 27683
rect 12592 27651 12624 27683
rect 12664 27651 12696 27683
rect 12736 27651 12768 27683
rect 12808 27651 12840 27683
rect 12880 27651 12912 27683
rect 12952 27651 12984 27683
rect 13024 27651 13056 27683
rect 13096 27651 13128 27683
rect 13168 27651 13200 27683
rect 13240 27651 13272 27683
rect 13312 27651 13344 27683
rect 13384 27651 13416 27683
rect 13456 27651 13488 27683
rect 13528 27651 13560 27683
rect 13600 27651 13632 27683
rect 13672 27651 13704 27683
rect 13744 27651 13776 27683
rect 13816 27651 13848 27683
rect 13888 27651 13920 27683
rect 13960 27651 13992 27683
rect 14032 27651 14064 27683
rect 14104 27651 14136 27683
rect 14176 27651 14208 27683
rect 14248 27651 14280 27683
rect 14320 27651 14352 27683
rect 14392 27651 14424 27683
rect 14464 27651 14496 27683
rect 14536 27651 14568 27683
rect 14608 27651 14640 27683
rect 14680 27651 14712 27683
rect 14752 27651 14784 27683
rect 14824 27651 14856 27683
rect 14896 27651 14928 27683
rect 14968 27651 15000 27683
rect 15040 27651 15072 27683
rect 15112 27651 15144 27683
rect 15184 27651 15216 27683
rect 15256 27651 15288 27683
rect 15328 27651 15360 27683
rect 15400 27651 15432 27683
rect 15472 27651 15504 27683
rect 15544 27651 15576 27683
rect 15616 27651 15648 27683
rect 15688 27651 15720 27683
rect 15760 27651 15792 27683
rect 15832 27651 15864 27683
rect 15904 27651 15936 27683
rect 64 27579 96 27611
rect 136 27579 168 27611
rect 208 27579 240 27611
rect 280 27579 312 27611
rect 352 27579 384 27611
rect 424 27579 456 27611
rect 496 27579 528 27611
rect 568 27579 600 27611
rect 640 27579 672 27611
rect 712 27579 744 27611
rect 784 27579 816 27611
rect 856 27579 888 27611
rect 928 27579 960 27611
rect 1000 27579 1032 27611
rect 1072 27579 1104 27611
rect 1144 27579 1176 27611
rect 1216 27579 1248 27611
rect 1288 27579 1320 27611
rect 1360 27579 1392 27611
rect 1432 27579 1464 27611
rect 1504 27579 1536 27611
rect 1576 27579 1608 27611
rect 1648 27579 1680 27611
rect 1720 27579 1752 27611
rect 1792 27579 1824 27611
rect 1864 27579 1896 27611
rect 1936 27579 1968 27611
rect 2008 27579 2040 27611
rect 2080 27579 2112 27611
rect 2152 27579 2184 27611
rect 2224 27579 2256 27611
rect 2296 27579 2328 27611
rect 2368 27579 2400 27611
rect 2440 27579 2472 27611
rect 2512 27579 2544 27611
rect 2584 27579 2616 27611
rect 2656 27579 2688 27611
rect 2728 27579 2760 27611
rect 2800 27579 2832 27611
rect 2872 27579 2904 27611
rect 2944 27579 2976 27611
rect 3016 27579 3048 27611
rect 3088 27579 3120 27611
rect 3160 27579 3192 27611
rect 3232 27579 3264 27611
rect 3304 27579 3336 27611
rect 3376 27579 3408 27611
rect 3448 27579 3480 27611
rect 3520 27579 3552 27611
rect 3592 27579 3624 27611
rect 3664 27579 3696 27611
rect 3736 27579 3768 27611
rect 3808 27579 3840 27611
rect 3880 27579 3912 27611
rect 3952 27579 3984 27611
rect 4024 27579 4056 27611
rect 4096 27579 4128 27611
rect 4168 27579 4200 27611
rect 4240 27579 4272 27611
rect 4312 27579 4344 27611
rect 4384 27579 4416 27611
rect 4456 27579 4488 27611
rect 4528 27579 4560 27611
rect 4600 27579 4632 27611
rect 4672 27579 4704 27611
rect 4744 27579 4776 27611
rect 4816 27579 4848 27611
rect 4888 27579 4920 27611
rect 4960 27579 4992 27611
rect 5032 27579 5064 27611
rect 5104 27579 5136 27611
rect 5176 27579 5208 27611
rect 5248 27579 5280 27611
rect 5320 27579 5352 27611
rect 5392 27579 5424 27611
rect 5464 27579 5496 27611
rect 5536 27579 5568 27611
rect 5608 27579 5640 27611
rect 5680 27579 5712 27611
rect 5752 27579 5784 27611
rect 5824 27579 5856 27611
rect 5896 27579 5928 27611
rect 5968 27579 6000 27611
rect 6040 27579 6072 27611
rect 6112 27579 6144 27611
rect 6184 27579 6216 27611
rect 6256 27579 6288 27611
rect 6328 27579 6360 27611
rect 6400 27579 6432 27611
rect 6472 27579 6504 27611
rect 6544 27579 6576 27611
rect 6616 27579 6648 27611
rect 6688 27579 6720 27611
rect 6760 27579 6792 27611
rect 6832 27579 6864 27611
rect 6904 27579 6936 27611
rect 6976 27579 7008 27611
rect 7048 27579 7080 27611
rect 7120 27579 7152 27611
rect 7192 27579 7224 27611
rect 7264 27579 7296 27611
rect 7336 27579 7368 27611
rect 7408 27579 7440 27611
rect 7480 27579 7512 27611
rect 7552 27579 7584 27611
rect 7624 27579 7656 27611
rect 7696 27579 7728 27611
rect 7768 27579 7800 27611
rect 7840 27579 7872 27611
rect 7912 27579 7944 27611
rect 7984 27579 8016 27611
rect 8056 27579 8088 27611
rect 8128 27579 8160 27611
rect 8200 27579 8232 27611
rect 8272 27579 8304 27611
rect 8344 27579 8376 27611
rect 8416 27579 8448 27611
rect 8488 27579 8520 27611
rect 8560 27579 8592 27611
rect 8632 27579 8664 27611
rect 8704 27579 8736 27611
rect 8776 27579 8808 27611
rect 8848 27579 8880 27611
rect 8920 27579 8952 27611
rect 8992 27579 9024 27611
rect 9064 27579 9096 27611
rect 9136 27579 9168 27611
rect 9208 27579 9240 27611
rect 9280 27579 9312 27611
rect 9352 27579 9384 27611
rect 9424 27579 9456 27611
rect 9496 27579 9528 27611
rect 9568 27579 9600 27611
rect 9640 27579 9672 27611
rect 9712 27579 9744 27611
rect 9784 27579 9816 27611
rect 9856 27579 9888 27611
rect 9928 27579 9960 27611
rect 10000 27579 10032 27611
rect 10072 27579 10104 27611
rect 10144 27579 10176 27611
rect 10216 27579 10248 27611
rect 10288 27579 10320 27611
rect 10360 27579 10392 27611
rect 10432 27579 10464 27611
rect 10504 27579 10536 27611
rect 10576 27579 10608 27611
rect 10648 27579 10680 27611
rect 10720 27579 10752 27611
rect 10792 27579 10824 27611
rect 10864 27579 10896 27611
rect 10936 27579 10968 27611
rect 11008 27579 11040 27611
rect 11080 27579 11112 27611
rect 11152 27579 11184 27611
rect 11224 27579 11256 27611
rect 11296 27579 11328 27611
rect 11368 27579 11400 27611
rect 11440 27579 11472 27611
rect 11512 27579 11544 27611
rect 11584 27579 11616 27611
rect 11656 27579 11688 27611
rect 11728 27579 11760 27611
rect 11800 27579 11832 27611
rect 11872 27579 11904 27611
rect 11944 27579 11976 27611
rect 12016 27579 12048 27611
rect 12088 27579 12120 27611
rect 12160 27579 12192 27611
rect 12232 27579 12264 27611
rect 12304 27579 12336 27611
rect 12376 27579 12408 27611
rect 12448 27579 12480 27611
rect 12520 27579 12552 27611
rect 12592 27579 12624 27611
rect 12664 27579 12696 27611
rect 12736 27579 12768 27611
rect 12808 27579 12840 27611
rect 12880 27579 12912 27611
rect 12952 27579 12984 27611
rect 13024 27579 13056 27611
rect 13096 27579 13128 27611
rect 13168 27579 13200 27611
rect 13240 27579 13272 27611
rect 13312 27579 13344 27611
rect 13384 27579 13416 27611
rect 13456 27579 13488 27611
rect 13528 27579 13560 27611
rect 13600 27579 13632 27611
rect 13672 27579 13704 27611
rect 13744 27579 13776 27611
rect 13816 27579 13848 27611
rect 13888 27579 13920 27611
rect 13960 27579 13992 27611
rect 14032 27579 14064 27611
rect 14104 27579 14136 27611
rect 14176 27579 14208 27611
rect 14248 27579 14280 27611
rect 14320 27579 14352 27611
rect 14392 27579 14424 27611
rect 14464 27579 14496 27611
rect 14536 27579 14568 27611
rect 14608 27579 14640 27611
rect 14680 27579 14712 27611
rect 14752 27579 14784 27611
rect 14824 27579 14856 27611
rect 14896 27579 14928 27611
rect 14968 27579 15000 27611
rect 15040 27579 15072 27611
rect 15112 27579 15144 27611
rect 15184 27579 15216 27611
rect 15256 27579 15288 27611
rect 15328 27579 15360 27611
rect 15400 27579 15432 27611
rect 15472 27579 15504 27611
rect 15544 27579 15576 27611
rect 15616 27579 15648 27611
rect 15688 27579 15720 27611
rect 15760 27579 15792 27611
rect 15832 27579 15864 27611
rect 15904 27579 15936 27611
rect 64 27507 96 27539
rect 136 27507 168 27539
rect 208 27507 240 27539
rect 280 27507 312 27539
rect 352 27507 384 27539
rect 424 27507 456 27539
rect 496 27507 528 27539
rect 568 27507 600 27539
rect 640 27507 672 27539
rect 712 27507 744 27539
rect 784 27507 816 27539
rect 856 27507 888 27539
rect 928 27507 960 27539
rect 1000 27507 1032 27539
rect 1072 27507 1104 27539
rect 1144 27507 1176 27539
rect 1216 27507 1248 27539
rect 1288 27507 1320 27539
rect 1360 27507 1392 27539
rect 1432 27507 1464 27539
rect 1504 27507 1536 27539
rect 1576 27507 1608 27539
rect 1648 27507 1680 27539
rect 1720 27507 1752 27539
rect 1792 27507 1824 27539
rect 1864 27507 1896 27539
rect 1936 27507 1968 27539
rect 2008 27507 2040 27539
rect 2080 27507 2112 27539
rect 2152 27507 2184 27539
rect 2224 27507 2256 27539
rect 2296 27507 2328 27539
rect 2368 27507 2400 27539
rect 2440 27507 2472 27539
rect 2512 27507 2544 27539
rect 2584 27507 2616 27539
rect 2656 27507 2688 27539
rect 2728 27507 2760 27539
rect 2800 27507 2832 27539
rect 2872 27507 2904 27539
rect 2944 27507 2976 27539
rect 3016 27507 3048 27539
rect 3088 27507 3120 27539
rect 3160 27507 3192 27539
rect 3232 27507 3264 27539
rect 3304 27507 3336 27539
rect 3376 27507 3408 27539
rect 3448 27507 3480 27539
rect 3520 27507 3552 27539
rect 3592 27507 3624 27539
rect 3664 27507 3696 27539
rect 3736 27507 3768 27539
rect 3808 27507 3840 27539
rect 3880 27507 3912 27539
rect 3952 27507 3984 27539
rect 4024 27507 4056 27539
rect 4096 27507 4128 27539
rect 4168 27507 4200 27539
rect 4240 27507 4272 27539
rect 4312 27507 4344 27539
rect 4384 27507 4416 27539
rect 4456 27507 4488 27539
rect 4528 27507 4560 27539
rect 4600 27507 4632 27539
rect 4672 27507 4704 27539
rect 4744 27507 4776 27539
rect 4816 27507 4848 27539
rect 4888 27507 4920 27539
rect 4960 27507 4992 27539
rect 5032 27507 5064 27539
rect 5104 27507 5136 27539
rect 5176 27507 5208 27539
rect 5248 27507 5280 27539
rect 5320 27507 5352 27539
rect 5392 27507 5424 27539
rect 5464 27507 5496 27539
rect 5536 27507 5568 27539
rect 5608 27507 5640 27539
rect 5680 27507 5712 27539
rect 5752 27507 5784 27539
rect 5824 27507 5856 27539
rect 5896 27507 5928 27539
rect 5968 27507 6000 27539
rect 6040 27507 6072 27539
rect 6112 27507 6144 27539
rect 6184 27507 6216 27539
rect 6256 27507 6288 27539
rect 6328 27507 6360 27539
rect 6400 27507 6432 27539
rect 6472 27507 6504 27539
rect 6544 27507 6576 27539
rect 6616 27507 6648 27539
rect 6688 27507 6720 27539
rect 6760 27507 6792 27539
rect 6832 27507 6864 27539
rect 6904 27507 6936 27539
rect 6976 27507 7008 27539
rect 7048 27507 7080 27539
rect 7120 27507 7152 27539
rect 7192 27507 7224 27539
rect 7264 27507 7296 27539
rect 7336 27507 7368 27539
rect 7408 27507 7440 27539
rect 7480 27507 7512 27539
rect 7552 27507 7584 27539
rect 7624 27507 7656 27539
rect 7696 27507 7728 27539
rect 7768 27507 7800 27539
rect 7840 27507 7872 27539
rect 7912 27507 7944 27539
rect 7984 27507 8016 27539
rect 8056 27507 8088 27539
rect 8128 27507 8160 27539
rect 8200 27507 8232 27539
rect 8272 27507 8304 27539
rect 8344 27507 8376 27539
rect 8416 27507 8448 27539
rect 8488 27507 8520 27539
rect 8560 27507 8592 27539
rect 8632 27507 8664 27539
rect 8704 27507 8736 27539
rect 8776 27507 8808 27539
rect 8848 27507 8880 27539
rect 8920 27507 8952 27539
rect 8992 27507 9024 27539
rect 9064 27507 9096 27539
rect 9136 27507 9168 27539
rect 9208 27507 9240 27539
rect 9280 27507 9312 27539
rect 9352 27507 9384 27539
rect 9424 27507 9456 27539
rect 9496 27507 9528 27539
rect 9568 27507 9600 27539
rect 9640 27507 9672 27539
rect 9712 27507 9744 27539
rect 9784 27507 9816 27539
rect 9856 27507 9888 27539
rect 9928 27507 9960 27539
rect 10000 27507 10032 27539
rect 10072 27507 10104 27539
rect 10144 27507 10176 27539
rect 10216 27507 10248 27539
rect 10288 27507 10320 27539
rect 10360 27507 10392 27539
rect 10432 27507 10464 27539
rect 10504 27507 10536 27539
rect 10576 27507 10608 27539
rect 10648 27507 10680 27539
rect 10720 27507 10752 27539
rect 10792 27507 10824 27539
rect 10864 27507 10896 27539
rect 10936 27507 10968 27539
rect 11008 27507 11040 27539
rect 11080 27507 11112 27539
rect 11152 27507 11184 27539
rect 11224 27507 11256 27539
rect 11296 27507 11328 27539
rect 11368 27507 11400 27539
rect 11440 27507 11472 27539
rect 11512 27507 11544 27539
rect 11584 27507 11616 27539
rect 11656 27507 11688 27539
rect 11728 27507 11760 27539
rect 11800 27507 11832 27539
rect 11872 27507 11904 27539
rect 11944 27507 11976 27539
rect 12016 27507 12048 27539
rect 12088 27507 12120 27539
rect 12160 27507 12192 27539
rect 12232 27507 12264 27539
rect 12304 27507 12336 27539
rect 12376 27507 12408 27539
rect 12448 27507 12480 27539
rect 12520 27507 12552 27539
rect 12592 27507 12624 27539
rect 12664 27507 12696 27539
rect 12736 27507 12768 27539
rect 12808 27507 12840 27539
rect 12880 27507 12912 27539
rect 12952 27507 12984 27539
rect 13024 27507 13056 27539
rect 13096 27507 13128 27539
rect 13168 27507 13200 27539
rect 13240 27507 13272 27539
rect 13312 27507 13344 27539
rect 13384 27507 13416 27539
rect 13456 27507 13488 27539
rect 13528 27507 13560 27539
rect 13600 27507 13632 27539
rect 13672 27507 13704 27539
rect 13744 27507 13776 27539
rect 13816 27507 13848 27539
rect 13888 27507 13920 27539
rect 13960 27507 13992 27539
rect 14032 27507 14064 27539
rect 14104 27507 14136 27539
rect 14176 27507 14208 27539
rect 14248 27507 14280 27539
rect 14320 27507 14352 27539
rect 14392 27507 14424 27539
rect 14464 27507 14496 27539
rect 14536 27507 14568 27539
rect 14608 27507 14640 27539
rect 14680 27507 14712 27539
rect 14752 27507 14784 27539
rect 14824 27507 14856 27539
rect 14896 27507 14928 27539
rect 14968 27507 15000 27539
rect 15040 27507 15072 27539
rect 15112 27507 15144 27539
rect 15184 27507 15216 27539
rect 15256 27507 15288 27539
rect 15328 27507 15360 27539
rect 15400 27507 15432 27539
rect 15472 27507 15504 27539
rect 15544 27507 15576 27539
rect 15616 27507 15648 27539
rect 15688 27507 15720 27539
rect 15760 27507 15792 27539
rect 15832 27507 15864 27539
rect 15904 27507 15936 27539
rect 64 27435 96 27467
rect 136 27435 168 27467
rect 208 27435 240 27467
rect 280 27435 312 27467
rect 352 27435 384 27467
rect 424 27435 456 27467
rect 496 27435 528 27467
rect 568 27435 600 27467
rect 640 27435 672 27467
rect 712 27435 744 27467
rect 784 27435 816 27467
rect 856 27435 888 27467
rect 928 27435 960 27467
rect 1000 27435 1032 27467
rect 1072 27435 1104 27467
rect 1144 27435 1176 27467
rect 1216 27435 1248 27467
rect 1288 27435 1320 27467
rect 1360 27435 1392 27467
rect 1432 27435 1464 27467
rect 1504 27435 1536 27467
rect 1576 27435 1608 27467
rect 1648 27435 1680 27467
rect 1720 27435 1752 27467
rect 1792 27435 1824 27467
rect 1864 27435 1896 27467
rect 1936 27435 1968 27467
rect 2008 27435 2040 27467
rect 2080 27435 2112 27467
rect 2152 27435 2184 27467
rect 2224 27435 2256 27467
rect 2296 27435 2328 27467
rect 2368 27435 2400 27467
rect 2440 27435 2472 27467
rect 2512 27435 2544 27467
rect 2584 27435 2616 27467
rect 2656 27435 2688 27467
rect 2728 27435 2760 27467
rect 2800 27435 2832 27467
rect 2872 27435 2904 27467
rect 2944 27435 2976 27467
rect 3016 27435 3048 27467
rect 3088 27435 3120 27467
rect 3160 27435 3192 27467
rect 3232 27435 3264 27467
rect 3304 27435 3336 27467
rect 3376 27435 3408 27467
rect 3448 27435 3480 27467
rect 3520 27435 3552 27467
rect 3592 27435 3624 27467
rect 3664 27435 3696 27467
rect 3736 27435 3768 27467
rect 3808 27435 3840 27467
rect 3880 27435 3912 27467
rect 3952 27435 3984 27467
rect 4024 27435 4056 27467
rect 4096 27435 4128 27467
rect 4168 27435 4200 27467
rect 4240 27435 4272 27467
rect 4312 27435 4344 27467
rect 4384 27435 4416 27467
rect 4456 27435 4488 27467
rect 4528 27435 4560 27467
rect 4600 27435 4632 27467
rect 4672 27435 4704 27467
rect 4744 27435 4776 27467
rect 4816 27435 4848 27467
rect 4888 27435 4920 27467
rect 4960 27435 4992 27467
rect 5032 27435 5064 27467
rect 5104 27435 5136 27467
rect 5176 27435 5208 27467
rect 5248 27435 5280 27467
rect 5320 27435 5352 27467
rect 5392 27435 5424 27467
rect 5464 27435 5496 27467
rect 5536 27435 5568 27467
rect 5608 27435 5640 27467
rect 5680 27435 5712 27467
rect 5752 27435 5784 27467
rect 5824 27435 5856 27467
rect 5896 27435 5928 27467
rect 5968 27435 6000 27467
rect 6040 27435 6072 27467
rect 6112 27435 6144 27467
rect 6184 27435 6216 27467
rect 6256 27435 6288 27467
rect 6328 27435 6360 27467
rect 6400 27435 6432 27467
rect 6472 27435 6504 27467
rect 6544 27435 6576 27467
rect 6616 27435 6648 27467
rect 6688 27435 6720 27467
rect 6760 27435 6792 27467
rect 6832 27435 6864 27467
rect 6904 27435 6936 27467
rect 6976 27435 7008 27467
rect 7048 27435 7080 27467
rect 7120 27435 7152 27467
rect 7192 27435 7224 27467
rect 7264 27435 7296 27467
rect 7336 27435 7368 27467
rect 7408 27435 7440 27467
rect 7480 27435 7512 27467
rect 7552 27435 7584 27467
rect 7624 27435 7656 27467
rect 7696 27435 7728 27467
rect 7768 27435 7800 27467
rect 7840 27435 7872 27467
rect 7912 27435 7944 27467
rect 7984 27435 8016 27467
rect 8056 27435 8088 27467
rect 8128 27435 8160 27467
rect 8200 27435 8232 27467
rect 8272 27435 8304 27467
rect 8344 27435 8376 27467
rect 8416 27435 8448 27467
rect 8488 27435 8520 27467
rect 8560 27435 8592 27467
rect 8632 27435 8664 27467
rect 8704 27435 8736 27467
rect 8776 27435 8808 27467
rect 8848 27435 8880 27467
rect 8920 27435 8952 27467
rect 8992 27435 9024 27467
rect 9064 27435 9096 27467
rect 9136 27435 9168 27467
rect 9208 27435 9240 27467
rect 9280 27435 9312 27467
rect 9352 27435 9384 27467
rect 9424 27435 9456 27467
rect 9496 27435 9528 27467
rect 9568 27435 9600 27467
rect 9640 27435 9672 27467
rect 9712 27435 9744 27467
rect 9784 27435 9816 27467
rect 9856 27435 9888 27467
rect 9928 27435 9960 27467
rect 10000 27435 10032 27467
rect 10072 27435 10104 27467
rect 10144 27435 10176 27467
rect 10216 27435 10248 27467
rect 10288 27435 10320 27467
rect 10360 27435 10392 27467
rect 10432 27435 10464 27467
rect 10504 27435 10536 27467
rect 10576 27435 10608 27467
rect 10648 27435 10680 27467
rect 10720 27435 10752 27467
rect 10792 27435 10824 27467
rect 10864 27435 10896 27467
rect 10936 27435 10968 27467
rect 11008 27435 11040 27467
rect 11080 27435 11112 27467
rect 11152 27435 11184 27467
rect 11224 27435 11256 27467
rect 11296 27435 11328 27467
rect 11368 27435 11400 27467
rect 11440 27435 11472 27467
rect 11512 27435 11544 27467
rect 11584 27435 11616 27467
rect 11656 27435 11688 27467
rect 11728 27435 11760 27467
rect 11800 27435 11832 27467
rect 11872 27435 11904 27467
rect 11944 27435 11976 27467
rect 12016 27435 12048 27467
rect 12088 27435 12120 27467
rect 12160 27435 12192 27467
rect 12232 27435 12264 27467
rect 12304 27435 12336 27467
rect 12376 27435 12408 27467
rect 12448 27435 12480 27467
rect 12520 27435 12552 27467
rect 12592 27435 12624 27467
rect 12664 27435 12696 27467
rect 12736 27435 12768 27467
rect 12808 27435 12840 27467
rect 12880 27435 12912 27467
rect 12952 27435 12984 27467
rect 13024 27435 13056 27467
rect 13096 27435 13128 27467
rect 13168 27435 13200 27467
rect 13240 27435 13272 27467
rect 13312 27435 13344 27467
rect 13384 27435 13416 27467
rect 13456 27435 13488 27467
rect 13528 27435 13560 27467
rect 13600 27435 13632 27467
rect 13672 27435 13704 27467
rect 13744 27435 13776 27467
rect 13816 27435 13848 27467
rect 13888 27435 13920 27467
rect 13960 27435 13992 27467
rect 14032 27435 14064 27467
rect 14104 27435 14136 27467
rect 14176 27435 14208 27467
rect 14248 27435 14280 27467
rect 14320 27435 14352 27467
rect 14392 27435 14424 27467
rect 14464 27435 14496 27467
rect 14536 27435 14568 27467
rect 14608 27435 14640 27467
rect 14680 27435 14712 27467
rect 14752 27435 14784 27467
rect 14824 27435 14856 27467
rect 14896 27435 14928 27467
rect 14968 27435 15000 27467
rect 15040 27435 15072 27467
rect 15112 27435 15144 27467
rect 15184 27435 15216 27467
rect 15256 27435 15288 27467
rect 15328 27435 15360 27467
rect 15400 27435 15432 27467
rect 15472 27435 15504 27467
rect 15544 27435 15576 27467
rect 15616 27435 15648 27467
rect 15688 27435 15720 27467
rect 15760 27435 15792 27467
rect 15832 27435 15864 27467
rect 15904 27435 15936 27467
rect 64 27363 96 27395
rect 136 27363 168 27395
rect 208 27363 240 27395
rect 280 27363 312 27395
rect 352 27363 384 27395
rect 424 27363 456 27395
rect 496 27363 528 27395
rect 568 27363 600 27395
rect 640 27363 672 27395
rect 712 27363 744 27395
rect 784 27363 816 27395
rect 856 27363 888 27395
rect 928 27363 960 27395
rect 1000 27363 1032 27395
rect 1072 27363 1104 27395
rect 1144 27363 1176 27395
rect 1216 27363 1248 27395
rect 1288 27363 1320 27395
rect 1360 27363 1392 27395
rect 1432 27363 1464 27395
rect 1504 27363 1536 27395
rect 1576 27363 1608 27395
rect 1648 27363 1680 27395
rect 1720 27363 1752 27395
rect 1792 27363 1824 27395
rect 1864 27363 1896 27395
rect 1936 27363 1968 27395
rect 2008 27363 2040 27395
rect 2080 27363 2112 27395
rect 2152 27363 2184 27395
rect 2224 27363 2256 27395
rect 2296 27363 2328 27395
rect 2368 27363 2400 27395
rect 2440 27363 2472 27395
rect 2512 27363 2544 27395
rect 2584 27363 2616 27395
rect 2656 27363 2688 27395
rect 2728 27363 2760 27395
rect 2800 27363 2832 27395
rect 2872 27363 2904 27395
rect 2944 27363 2976 27395
rect 3016 27363 3048 27395
rect 3088 27363 3120 27395
rect 3160 27363 3192 27395
rect 3232 27363 3264 27395
rect 3304 27363 3336 27395
rect 3376 27363 3408 27395
rect 3448 27363 3480 27395
rect 3520 27363 3552 27395
rect 3592 27363 3624 27395
rect 3664 27363 3696 27395
rect 3736 27363 3768 27395
rect 3808 27363 3840 27395
rect 3880 27363 3912 27395
rect 3952 27363 3984 27395
rect 4024 27363 4056 27395
rect 4096 27363 4128 27395
rect 4168 27363 4200 27395
rect 4240 27363 4272 27395
rect 4312 27363 4344 27395
rect 4384 27363 4416 27395
rect 4456 27363 4488 27395
rect 4528 27363 4560 27395
rect 4600 27363 4632 27395
rect 4672 27363 4704 27395
rect 4744 27363 4776 27395
rect 4816 27363 4848 27395
rect 4888 27363 4920 27395
rect 4960 27363 4992 27395
rect 5032 27363 5064 27395
rect 5104 27363 5136 27395
rect 5176 27363 5208 27395
rect 5248 27363 5280 27395
rect 5320 27363 5352 27395
rect 5392 27363 5424 27395
rect 5464 27363 5496 27395
rect 5536 27363 5568 27395
rect 5608 27363 5640 27395
rect 5680 27363 5712 27395
rect 5752 27363 5784 27395
rect 5824 27363 5856 27395
rect 5896 27363 5928 27395
rect 5968 27363 6000 27395
rect 6040 27363 6072 27395
rect 6112 27363 6144 27395
rect 6184 27363 6216 27395
rect 6256 27363 6288 27395
rect 6328 27363 6360 27395
rect 6400 27363 6432 27395
rect 6472 27363 6504 27395
rect 6544 27363 6576 27395
rect 6616 27363 6648 27395
rect 6688 27363 6720 27395
rect 6760 27363 6792 27395
rect 6832 27363 6864 27395
rect 6904 27363 6936 27395
rect 6976 27363 7008 27395
rect 7048 27363 7080 27395
rect 7120 27363 7152 27395
rect 7192 27363 7224 27395
rect 7264 27363 7296 27395
rect 7336 27363 7368 27395
rect 7408 27363 7440 27395
rect 7480 27363 7512 27395
rect 7552 27363 7584 27395
rect 7624 27363 7656 27395
rect 7696 27363 7728 27395
rect 7768 27363 7800 27395
rect 7840 27363 7872 27395
rect 7912 27363 7944 27395
rect 7984 27363 8016 27395
rect 8056 27363 8088 27395
rect 8128 27363 8160 27395
rect 8200 27363 8232 27395
rect 8272 27363 8304 27395
rect 8344 27363 8376 27395
rect 8416 27363 8448 27395
rect 8488 27363 8520 27395
rect 8560 27363 8592 27395
rect 8632 27363 8664 27395
rect 8704 27363 8736 27395
rect 8776 27363 8808 27395
rect 8848 27363 8880 27395
rect 8920 27363 8952 27395
rect 8992 27363 9024 27395
rect 9064 27363 9096 27395
rect 9136 27363 9168 27395
rect 9208 27363 9240 27395
rect 9280 27363 9312 27395
rect 9352 27363 9384 27395
rect 9424 27363 9456 27395
rect 9496 27363 9528 27395
rect 9568 27363 9600 27395
rect 9640 27363 9672 27395
rect 9712 27363 9744 27395
rect 9784 27363 9816 27395
rect 9856 27363 9888 27395
rect 9928 27363 9960 27395
rect 10000 27363 10032 27395
rect 10072 27363 10104 27395
rect 10144 27363 10176 27395
rect 10216 27363 10248 27395
rect 10288 27363 10320 27395
rect 10360 27363 10392 27395
rect 10432 27363 10464 27395
rect 10504 27363 10536 27395
rect 10576 27363 10608 27395
rect 10648 27363 10680 27395
rect 10720 27363 10752 27395
rect 10792 27363 10824 27395
rect 10864 27363 10896 27395
rect 10936 27363 10968 27395
rect 11008 27363 11040 27395
rect 11080 27363 11112 27395
rect 11152 27363 11184 27395
rect 11224 27363 11256 27395
rect 11296 27363 11328 27395
rect 11368 27363 11400 27395
rect 11440 27363 11472 27395
rect 11512 27363 11544 27395
rect 11584 27363 11616 27395
rect 11656 27363 11688 27395
rect 11728 27363 11760 27395
rect 11800 27363 11832 27395
rect 11872 27363 11904 27395
rect 11944 27363 11976 27395
rect 12016 27363 12048 27395
rect 12088 27363 12120 27395
rect 12160 27363 12192 27395
rect 12232 27363 12264 27395
rect 12304 27363 12336 27395
rect 12376 27363 12408 27395
rect 12448 27363 12480 27395
rect 12520 27363 12552 27395
rect 12592 27363 12624 27395
rect 12664 27363 12696 27395
rect 12736 27363 12768 27395
rect 12808 27363 12840 27395
rect 12880 27363 12912 27395
rect 12952 27363 12984 27395
rect 13024 27363 13056 27395
rect 13096 27363 13128 27395
rect 13168 27363 13200 27395
rect 13240 27363 13272 27395
rect 13312 27363 13344 27395
rect 13384 27363 13416 27395
rect 13456 27363 13488 27395
rect 13528 27363 13560 27395
rect 13600 27363 13632 27395
rect 13672 27363 13704 27395
rect 13744 27363 13776 27395
rect 13816 27363 13848 27395
rect 13888 27363 13920 27395
rect 13960 27363 13992 27395
rect 14032 27363 14064 27395
rect 14104 27363 14136 27395
rect 14176 27363 14208 27395
rect 14248 27363 14280 27395
rect 14320 27363 14352 27395
rect 14392 27363 14424 27395
rect 14464 27363 14496 27395
rect 14536 27363 14568 27395
rect 14608 27363 14640 27395
rect 14680 27363 14712 27395
rect 14752 27363 14784 27395
rect 14824 27363 14856 27395
rect 14896 27363 14928 27395
rect 14968 27363 15000 27395
rect 15040 27363 15072 27395
rect 15112 27363 15144 27395
rect 15184 27363 15216 27395
rect 15256 27363 15288 27395
rect 15328 27363 15360 27395
rect 15400 27363 15432 27395
rect 15472 27363 15504 27395
rect 15544 27363 15576 27395
rect 15616 27363 15648 27395
rect 15688 27363 15720 27395
rect 15760 27363 15792 27395
rect 15832 27363 15864 27395
rect 15904 27363 15936 27395
rect 64 27291 96 27323
rect 136 27291 168 27323
rect 208 27291 240 27323
rect 280 27291 312 27323
rect 352 27291 384 27323
rect 424 27291 456 27323
rect 496 27291 528 27323
rect 568 27291 600 27323
rect 640 27291 672 27323
rect 712 27291 744 27323
rect 784 27291 816 27323
rect 856 27291 888 27323
rect 928 27291 960 27323
rect 1000 27291 1032 27323
rect 1072 27291 1104 27323
rect 1144 27291 1176 27323
rect 1216 27291 1248 27323
rect 1288 27291 1320 27323
rect 1360 27291 1392 27323
rect 1432 27291 1464 27323
rect 1504 27291 1536 27323
rect 1576 27291 1608 27323
rect 1648 27291 1680 27323
rect 1720 27291 1752 27323
rect 1792 27291 1824 27323
rect 1864 27291 1896 27323
rect 1936 27291 1968 27323
rect 2008 27291 2040 27323
rect 2080 27291 2112 27323
rect 2152 27291 2184 27323
rect 2224 27291 2256 27323
rect 2296 27291 2328 27323
rect 2368 27291 2400 27323
rect 2440 27291 2472 27323
rect 2512 27291 2544 27323
rect 2584 27291 2616 27323
rect 2656 27291 2688 27323
rect 2728 27291 2760 27323
rect 2800 27291 2832 27323
rect 2872 27291 2904 27323
rect 2944 27291 2976 27323
rect 3016 27291 3048 27323
rect 3088 27291 3120 27323
rect 3160 27291 3192 27323
rect 3232 27291 3264 27323
rect 3304 27291 3336 27323
rect 3376 27291 3408 27323
rect 3448 27291 3480 27323
rect 3520 27291 3552 27323
rect 3592 27291 3624 27323
rect 3664 27291 3696 27323
rect 3736 27291 3768 27323
rect 3808 27291 3840 27323
rect 3880 27291 3912 27323
rect 3952 27291 3984 27323
rect 4024 27291 4056 27323
rect 4096 27291 4128 27323
rect 4168 27291 4200 27323
rect 4240 27291 4272 27323
rect 4312 27291 4344 27323
rect 4384 27291 4416 27323
rect 4456 27291 4488 27323
rect 4528 27291 4560 27323
rect 4600 27291 4632 27323
rect 4672 27291 4704 27323
rect 4744 27291 4776 27323
rect 4816 27291 4848 27323
rect 4888 27291 4920 27323
rect 4960 27291 4992 27323
rect 5032 27291 5064 27323
rect 5104 27291 5136 27323
rect 5176 27291 5208 27323
rect 5248 27291 5280 27323
rect 5320 27291 5352 27323
rect 5392 27291 5424 27323
rect 5464 27291 5496 27323
rect 5536 27291 5568 27323
rect 5608 27291 5640 27323
rect 5680 27291 5712 27323
rect 5752 27291 5784 27323
rect 5824 27291 5856 27323
rect 5896 27291 5928 27323
rect 5968 27291 6000 27323
rect 6040 27291 6072 27323
rect 6112 27291 6144 27323
rect 6184 27291 6216 27323
rect 6256 27291 6288 27323
rect 6328 27291 6360 27323
rect 6400 27291 6432 27323
rect 6472 27291 6504 27323
rect 6544 27291 6576 27323
rect 6616 27291 6648 27323
rect 6688 27291 6720 27323
rect 6760 27291 6792 27323
rect 6832 27291 6864 27323
rect 6904 27291 6936 27323
rect 6976 27291 7008 27323
rect 7048 27291 7080 27323
rect 7120 27291 7152 27323
rect 7192 27291 7224 27323
rect 7264 27291 7296 27323
rect 7336 27291 7368 27323
rect 7408 27291 7440 27323
rect 7480 27291 7512 27323
rect 7552 27291 7584 27323
rect 7624 27291 7656 27323
rect 7696 27291 7728 27323
rect 7768 27291 7800 27323
rect 7840 27291 7872 27323
rect 7912 27291 7944 27323
rect 7984 27291 8016 27323
rect 8056 27291 8088 27323
rect 8128 27291 8160 27323
rect 8200 27291 8232 27323
rect 8272 27291 8304 27323
rect 8344 27291 8376 27323
rect 8416 27291 8448 27323
rect 8488 27291 8520 27323
rect 8560 27291 8592 27323
rect 8632 27291 8664 27323
rect 8704 27291 8736 27323
rect 8776 27291 8808 27323
rect 8848 27291 8880 27323
rect 8920 27291 8952 27323
rect 8992 27291 9024 27323
rect 9064 27291 9096 27323
rect 9136 27291 9168 27323
rect 9208 27291 9240 27323
rect 9280 27291 9312 27323
rect 9352 27291 9384 27323
rect 9424 27291 9456 27323
rect 9496 27291 9528 27323
rect 9568 27291 9600 27323
rect 9640 27291 9672 27323
rect 9712 27291 9744 27323
rect 9784 27291 9816 27323
rect 9856 27291 9888 27323
rect 9928 27291 9960 27323
rect 10000 27291 10032 27323
rect 10072 27291 10104 27323
rect 10144 27291 10176 27323
rect 10216 27291 10248 27323
rect 10288 27291 10320 27323
rect 10360 27291 10392 27323
rect 10432 27291 10464 27323
rect 10504 27291 10536 27323
rect 10576 27291 10608 27323
rect 10648 27291 10680 27323
rect 10720 27291 10752 27323
rect 10792 27291 10824 27323
rect 10864 27291 10896 27323
rect 10936 27291 10968 27323
rect 11008 27291 11040 27323
rect 11080 27291 11112 27323
rect 11152 27291 11184 27323
rect 11224 27291 11256 27323
rect 11296 27291 11328 27323
rect 11368 27291 11400 27323
rect 11440 27291 11472 27323
rect 11512 27291 11544 27323
rect 11584 27291 11616 27323
rect 11656 27291 11688 27323
rect 11728 27291 11760 27323
rect 11800 27291 11832 27323
rect 11872 27291 11904 27323
rect 11944 27291 11976 27323
rect 12016 27291 12048 27323
rect 12088 27291 12120 27323
rect 12160 27291 12192 27323
rect 12232 27291 12264 27323
rect 12304 27291 12336 27323
rect 12376 27291 12408 27323
rect 12448 27291 12480 27323
rect 12520 27291 12552 27323
rect 12592 27291 12624 27323
rect 12664 27291 12696 27323
rect 12736 27291 12768 27323
rect 12808 27291 12840 27323
rect 12880 27291 12912 27323
rect 12952 27291 12984 27323
rect 13024 27291 13056 27323
rect 13096 27291 13128 27323
rect 13168 27291 13200 27323
rect 13240 27291 13272 27323
rect 13312 27291 13344 27323
rect 13384 27291 13416 27323
rect 13456 27291 13488 27323
rect 13528 27291 13560 27323
rect 13600 27291 13632 27323
rect 13672 27291 13704 27323
rect 13744 27291 13776 27323
rect 13816 27291 13848 27323
rect 13888 27291 13920 27323
rect 13960 27291 13992 27323
rect 14032 27291 14064 27323
rect 14104 27291 14136 27323
rect 14176 27291 14208 27323
rect 14248 27291 14280 27323
rect 14320 27291 14352 27323
rect 14392 27291 14424 27323
rect 14464 27291 14496 27323
rect 14536 27291 14568 27323
rect 14608 27291 14640 27323
rect 14680 27291 14712 27323
rect 14752 27291 14784 27323
rect 14824 27291 14856 27323
rect 14896 27291 14928 27323
rect 14968 27291 15000 27323
rect 15040 27291 15072 27323
rect 15112 27291 15144 27323
rect 15184 27291 15216 27323
rect 15256 27291 15288 27323
rect 15328 27291 15360 27323
rect 15400 27291 15432 27323
rect 15472 27291 15504 27323
rect 15544 27291 15576 27323
rect 15616 27291 15648 27323
rect 15688 27291 15720 27323
rect 15760 27291 15792 27323
rect 15832 27291 15864 27323
rect 15904 27291 15936 27323
rect 64 27219 96 27251
rect 136 27219 168 27251
rect 208 27219 240 27251
rect 280 27219 312 27251
rect 352 27219 384 27251
rect 424 27219 456 27251
rect 496 27219 528 27251
rect 568 27219 600 27251
rect 640 27219 672 27251
rect 712 27219 744 27251
rect 784 27219 816 27251
rect 856 27219 888 27251
rect 928 27219 960 27251
rect 1000 27219 1032 27251
rect 1072 27219 1104 27251
rect 1144 27219 1176 27251
rect 1216 27219 1248 27251
rect 1288 27219 1320 27251
rect 1360 27219 1392 27251
rect 1432 27219 1464 27251
rect 1504 27219 1536 27251
rect 1576 27219 1608 27251
rect 1648 27219 1680 27251
rect 1720 27219 1752 27251
rect 1792 27219 1824 27251
rect 1864 27219 1896 27251
rect 1936 27219 1968 27251
rect 2008 27219 2040 27251
rect 2080 27219 2112 27251
rect 2152 27219 2184 27251
rect 2224 27219 2256 27251
rect 2296 27219 2328 27251
rect 2368 27219 2400 27251
rect 2440 27219 2472 27251
rect 2512 27219 2544 27251
rect 2584 27219 2616 27251
rect 2656 27219 2688 27251
rect 2728 27219 2760 27251
rect 2800 27219 2832 27251
rect 2872 27219 2904 27251
rect 2944 27219 2976 27251
rect 3016 27219 3048 27251
rect 3088 27219 3120 27251
rect 3160 27219 3192 27251
rect 3232 27219 3264 27251
rect 3304 27219 3336 27251
rect 3376 27219 3408 27251
rect 3448 27219 3480 27251
rect 3520 27219 3552 27251
rect 3592 27219 3624 27251
rect 3664 27219 3696 27251
rect 3736 27219 3768 27251
rect 3808 27219 3840 27251
rect 3880 27219 3912 27251
rect 3952 27219 3984 27251
rect 4024 27219 4056 27251
rect 4096 27219 4128 27251
rect 4168 27219 4200 27251
rect 4240 27219 4272 27251
rect 4312 27219 4344 27251
rect 4384 27219 4416 27251
rect 4456 27219 4488 27251
rect 4528 27219 4560 27251
rect 4600 27219 4632 27251
rect 4672 27219 4704 27251
rect 4744 27219 4776 27251
rect 4816 27219 4848 27251
rect 4888 27219 4920 27251
rect 4960 27219 4992 27251
rect 5032 27219 5064 27251
rect 5104 27219 5136 27251
rect 5176 27219 5208 27251
rect 5248 27219 5280 27251
rect 5320 27219 5352 27251
rect 5392 27219 5424 27251
rect 5464 27219 5496 27251
rect 5536 27219 5568 27251
rect 5608 27219 5640 27251
rect 5680 27219 5712 27251
rect 5752 27219 5784 27251
rect 5824 27219 5856 27251
rect 5896 27219 5928 27251
rect 5968 27219 6000 27251
rect 6040 27219 6072 27251
rect 6112 27219 6144 27251
rect 6184 27219 6216 27251
rect 6256 27219 6288 27251
rect 6328 27219 6360 27251
rect 6400 27219 6432 27251
rect 6472 27219 6504 27251
rect 6544 27219 6576 27251
rect 6616 27219 6648 27251
rect 6688 27219 6720 27251
rect 6760 27219 6792 27251
rect 6832 27219 6864 27251
rect 6904 27219 6936 27251
rect 6976 27219 7008 27251
rect 7048 27219 7080 27251
rect 7120 27219 7152 27251
rect 7192 27219 7224 27251
rect 7264 27219 7296 27251
rect 7336 27219 7368 27251
rect 7408 27219 7440 27251
rect 7480 27219 7512 27251
rect 7552 27219 7584 27251
rect 7624 27219 7656 27251
rect 7696 27219 7728 27251
rect 7768 27219 7800 27251
rect 7840 27219 7872 27251
rect 7912 27219 7944 27251
rect 7984 27219 8016 27251
rect 8056 27219 8088 27251
rect 8128 27219 8160 27251
rect 8200 27219 8232 27251
rect 8272 27219 8304 27251
rect 8344 27219 8376 27251
rect 8416 27219 8448 27251
rect 8488 27219 8520 27251
rect 8560 27219 8592 27251
rect 8632 27219 8664 27251
rect 8704 27219 8736 27251
rect 8776 27219 8808 27251
rect 8848 27219 8880 27251
rect 8920 27219 8952 27251
rect 8992 27219 9024 27251
rect 9064 27219 9096 27251
rect 9136 27219 9168 27251
rect 9208 27219 9240 27251
rect 9280 27219 9312 27251
rect 9352 27219 9384 27251
rect 9424 27219 9456 27251
rect 9496 27219 9528 27251
rect 9568 27219 9600 27251
rect 9640 27219 9672 27251
rect 9712 27219 9744 27251
rect 9784 27219 9816 27251
rect 9856 27219 9888 27251
rect 9928 27219 9960 27251
rect 10000 27219 10032 27251
rect 10072 27219 10104 27251
rect 10144 27219 10176 27251
rect 10216 27219 10248 27251
rect 10288 27219 10320 27251
rect 10360 27219 10392 27251
rect 10432 27219 10464 27251
rect 10504 27219 10536 27251
rect 10576 27219 10608 27251
rect 10648 27219 10680 27251
rect 10720 27219 10752 27251
rect 10792 27219 10824 27251
rect 10864 27219 10896 27251
rect 10936 27219 10968 27251
rect 11008 27219 11040 27251
rect 11080 27219 11112 27251
rect 11152 27219 11184 27251
rect 11224 27219 11256 27251
rect 11296 27219 11328 27251
rect 11368 27219 11400 27251
rect 11440 27219 11472 27251
rect 11512 27219 11544 27251
rect 11584 27219 11616 27251
rect 11656 27219 11688 27251
rect 11728 27219 11760 27251
rect 11800 27219 11832 27251
rect 11872 27219 11904 27251
rect 11944 27219 11976 27251
rect 12016 27219 12048 27251
rect 12088 27219 12120 27251
rect 12160 27219 12192 27251
rect 12232 27219 12264 27251
rect 12304 27219 12336 27251
rect 12376 27219 12408 27251
rect 12448 27219 12480 27251
rect 12520 27219 12552 27251
rect 12592 27219 12624 27251
rect 12664 27219 12696 27251
rect 12736 27219 12768 27251
rect 12808 27219 12840 27251
rect 12880 27219 12912 27251
rect 12952 27219 12984 27251
rect 13024 27219 13056 27251
rect 13096 27219 13128 27251
rect 13168 27219 13200 27251
rect 13240 27219 13272 27251
rect 13312 27219 13344 27251
rect 13384 27219 13416 27251
rect 13456 27219 13488 27251
rect 13528 27219 13560 27251
rect 13600 27219 13632 27251
rect 13672 27219 13704 27251
rect 13744 27219 13776 27251
rect 13816 27219 13848 27251
rect 13888 27219 13920 27251
rect 13960 27219 13992 27251
rect 14032 27219 14064 27251
rect 14104 27219 14136 27251
rect 14176 27219 14208 27251
rect 14248 27219 14280 27251
rect 14320 27219 14352 27251
rect 14392 27219 14424 27251
rect 14464 27219 14496 27251
rect 14536 27219 14568 27251
rect 14608 27219 14640 27251
rect 14680 27219 14712 27251
rect 14752 27219 14784 27251
rect 14824 27219 14856 27251
rect 14896 27219 14928 27251
rect 14968 27219 15000 27251
rect 15040 27219 15072 27251
rect 15112 27219 15144 27251
rect 15184 27219 15216 27251
rect 15256 27219 15288 27251
rect 15328 27219 15360 27251
rect 15400 27219 15432 27251
rect 15472 27219 15504 27251
rect 15544 27219 15576 27251
rect 15616 27219 15648 27251
rect 15688 27219 15720 27251
rect 15760 27219 15792 27251
rect 15832 27219 15864 27251
rect 15904 27219 15936 27251
rect 64 27147 96 27179
rect 136 27147 168 27179
rect 208 27147 240 27179
rect 280 27147 312 27179
rect 352 27147 384 27179
rect 424 27147 456 27179
rect 496 27147 528 27179
rect 568 27147 600 27179
rect 640 27147 672 27179
rect 712 27147 744 27179
rect 784 27147 816 27179
rect 856 27147 888 27179
rect 928 27147 960 27179
rect 1000 27147 1032 27179
rect 1072 27147 1104 27179
rect 1144 27147 1176 27179
rect 1216 27147 1248 27179
rect 1288 27147 1320 27179
rect 1360 27147 1392 27179
rect 1432 27147 1464 27179
rect 1504 27147 1536 27179
rect 1576 27147 1608 27179
rect 1648 27147 1680 27179
rect 1720 27147 1752 27179
rect 1792 27147 1824 27179
rect 1864 27147 1896 27179
rect 1936 27147 1968 27179
rect 2008 27147 2040 27179
rect 2080 27147 2112 27179
rect 2152 27147 2184 27179
rect 2224 27147 2256 27179
rect 2296 27147 2328 27179
rect 2368 27147 2400 27179
rect 2440 27147 2472 27179
rect 2512 27147 2544 27179
rect 2584 27147 2616 27179
rect 2656 27147 2688 27179
rect 2728 27147 2760 27179
rect 2800 27147 2832 27179
rect 2872 27147 2904 27179
rect 2944 27147 2976 27179
rect 3016 27147 3048 27179
rect 3088 27147 3120 27179
rect 3160 27147 3192 27179
rect 3232 27147 3264 27179
rect 3304 27147 3336 27179
rect 3376 27147 3408 27179
rect 3448 27147 3480 27179
rect 3520 27147 3552 27179
rect 3592 27147 3624 27179
rect 3664 27147 3696 27179
rect 3736 27147 3768 27179
rect 3808 27147 3840 27179
rect 3880 27147 3912 27179
rect 3952 27147 3984 27179
rect 4024 27147 4056 27179
rect 4096 27147 4128 27179
rect 4168 27147 4200 27179
rect 4240 27147 4272 27179
rect 4312 27147 4344 27179
rect 4384 27147 4416 27179
rect 4456 27147 4488 27179
rect 4528 27147 4560 27179
rect 4600 27147 4632 27179
rect 4672 27147 4704 27179
rect 4744 27147 4776 27179
rect 4816 27147 4848 27179
rect 4888 27147 4920 27179
rect 4960 27147 4992 27179
rect 5032 27147 5064 27179
rect 5104 27147 5136 27179
rect 5176 27147 5208 27179
rect 5248 27147 5280 27179
rect 5320 27147 5352 27179
rect 5392 27147 5424 27179
rect 5464 27147 5496 27179
rect 5536 27147 5568 27179
rect 5608 27147 5640 27179
rect 5680 27147 5712 27179
rect 5752 27147 5784 27179
rect 5824 27147 5856 27179
rect 5896 27147 5928 27179
rect 5968 27147 6000 27179
rect 6040 27147 6072 27179
rect 6112 27147 6144 27179
rect 6184 27147 6216 27179
rect 6256 27147 6288 27179
rect 6328 27147 6360 27179
rect 6400 27147 6432 27179
rect 6472 27147 6504 27179
rect 6544 27147 6576 27179
rect 6616 27147 6648 27179
rect 6688 27147 6720 27179
rect 6760 27147 6792 27179
rect 6832 27147 6864 27179
rect 6904 27147 6936 27179
rect 6976 27147 7008 27179
rect 7048 27147 7080 27179
rect 7120 27147 7152 27179
rect 7192 27147 7224 27179
rect 7264 27147 7296 27179
rect 7336 27147 7368 27179
rect 7408 27147 7440 27179
rect 7480 27147 7512 27179
rect 7552 27147 7584 27179
rect 7624 27147 7656 27179
rect 7696 27147 7728 27179
rect 7768 27147 7800 27179
rect 7840 27147 7872 27179
rect 7912 27147 7944 27179
rect 7984 27147 8016 27179
rect 8056 27147 8088 27179
rect 8128 27147 8160 27179
rect 8200 27147 8232 27179
rect 8272 27147 8304 27179
rect 8344 27147 8376 27179
rect 8416 27147 8448 27179
rect 8488 27147 8520 27179
rect 8560 27147 8592 27179
rect 8632 27147 8664 27179
rect 8704 27147 8736 27179
rect 8776 27147 8808 27179
rect 8848 27147 8880 27179
rect 8920 27147 8952 27179
rect 8992 27147 9024 27179
rect 9064 27147 9096 27179
rect 9136 27147 9168 27179
rect 9208 27147 9240 27179
rect 9280 27147 9312 27179
rect 9352 27147 9384 27179
rect 9424 27147 9456 27179
rect 9496 27147 9528 27179
rect 9568 27147 9600 27179
rect 9640 27147 9672 27179
rect 9712 27147 9744 27179
rect 9784 27147 9816 27179
rect 9856 27147 9888 27179
rect 9928 27147 9960 27179
rect 10000 27147 10032 27179
rect 10072 27147 10104 27179
rect 10144 27147 10176 27179
rect 10216 27147 10248 27179
rect 10288 27147 10320 27179
rect 10360 27147 10392 27179
rect 10432 27147 10464 27179
rect 10504 27147 10536 27179
rect 10576 27147 10608 27179
rect 10648 27147 10680 27179
rect 10720 27147 10752 27179
rect 10792 27147 10824 27179
rect 10864 27147 10896 27179
rect 10936 27147 10968 27179
rect 11008 27147 11040 27179
rect 11080 27147 11112 27179
rect 11152 27147 11184 27179
rect 11224 27147 11256 27179
rect 11296 27147 11328 27179
rect 11368 27147 11400 27179
rect 11440 27147 11472 27179
rect 11512 27147 11544 27179
rect 11584 27147 11616 27179
rect 11656 27147 11688 27179
rect 11728 27147 11760 27179
rect 11800 27147 11832 27179
rect 11872 27147 11904 27179
rect 11944 27147 11976 27179
rect 12016 27147 12048 27179
rect 12088 27147 12120 27179
rect 12160 27147 12192 27179
rect 12232 27147 12264 27179
rect 12304 27147 12336 27179
rect 12376 27147 12408 27179
rect 12448 27147 12480 27179
rect 12520 27147 12552 27179
rect 12592 27147 12624 27179
rect 12664 27147 12696 27179
rect 12736 27147 12768 27179
rect 12808 27147 12840 27179
rect 12880 27147 12912 27179
rect 12952 27147 12984 27179
rect 13024 27147 13056 27179
rect 13096 27147 13128 27179
rect 13168 27147 13200 27179
rect 13240 27147 13272 27179
rect 13312 27147 13344 27179
rect 13384 27147 13416 27179
rect 13456 27147 13488 27179
rect 13528 27147 13560 27179
rect 13600 27147 13632 27179
rect 13672 27147 13704 27179
rect 13744 27147 13776 27179
rect 13816 27147 13848 27179
rect 13888 27147 13920 27179
rect 13960 27147 13992 27179
rect 14032 27147 14064 27179
rect 14104 27147 14136 27179
rect 14176 27147 14208 27179
rect 14248 27147 14280 27179
rect 14320 27147 14352 27179
rect 14392 27147 14424 27179
rect 14464 27147 14496 27179
rect 14536 27147 14568 27179
rect 14608 27147 14640 27179
rect 14680 27147 14712 27179
rect 14752 27147 14784 27179
rect 14824 27147 14856 27179
rect 14896 27147 14928 27179
rect 14968 27147 15000 27179
rect 15040 27147 15072 27179
rect 15112 27147 15144 27179
rect 15184 27147 15216 27179
rect 15256 27147 15288 27179
rect 15328 27147 15360 27179
rect 15400 27147 15432 27179
rect 15472 27147 15504 27179
rect 15544 27147 15576 27179
rect 15616 27147 15648 27179
rect 15688 27147 15720 27179
rect 15760 27147 15792 27179
rect 15832 27147 15864 27179
rect 15904 27147 15936 27179
rect 64 27075 96 27107
rect 136 27075 168 27107
rect 208 27075 240 27107
rect 280 27075 312 27107
rect 352 27075 384 27107
rect 424 27075 456 27107
rect 496 27075 528 27107
rect 568 27075 600 27107
rect 640 27075 672 27107
rect 712 27075 744 27107
rect 784 27075 816 27107
rect 856 27075 888 27107
rect 928 27075 960 27107
rect 1000 27075 1032 27107
rect 1072 27075 1104 27107
rect 1144 27075 1176 27107
rect 1216 27075 1248 27107
rect 1288 27075 1320 27107
rect 1360 27075 1392 27107
rect 1432 27075 1464 27107
rect 1504 27075 1536 27107
rect 1576 27075 1608 27107
rect 1648 27075 1680 27107
rect 1720 27075 1752 27107
rect 1792 27075 1824 27107
rect 1864 27075 1896 27107
rect 1936 27075 1968 27107
rect 2008 27075 2040 27107
rect 2080 27075 2112 27107
rect 2152 27075 2184 27107
rect 2224 27075 2256 27107
rect 2296 27075 2328 27107
rect 2368 27075 2400 27107
rect 2440 27075 2472 27107
rect 2512 27075 2544 27107
rect 2584 27075 2616 27107
rect 2656 27075 2688 27107
rect 2728 27075 2760 27107
rect 2800 27075 2832 27107
rect 2872 27075 2904 27107
rect 2944 27075 2976 27107
rect 3016 27075 3048 27107
rect 3088 27075 3120 27107
rect 3160 27075 3192 27107
rect 3232 27075 3264 27107
rect 3304 27075 3336 27107
rect 3376 27075 3408 27107
rect 3448 27075 3480 27107
rect 3520 27075 3552 27107
rect 3592 27075 3624 27107
rect 3664 27075 3696 27107
rect 3736 27075 3768 27107
rect 3808 27075 3840 27107
rect 3880 27075 3912 27107
rect 3952 27075 3984 27107
rect 4024 27075 4056 27107
rect 4096 27075 4128 27107
rect 4168 27075 4200 27107
rect 4240 27075 4272 27107
rect 4312 27075 4344 27107
rect 4384 27075 4416 27107
rect 4456 27075 4488 27107
rect 4528 27075 4560 27107
rect 4600 27075 4632 27107
rect 4672 27075 4704 27107
rect 4744 27075 4776 27107
rect 4816 27075 4848 27107
rect 4888 27075 4920 27107
rect 4960 27075 4992 27107
rect 5032 27075 5064 27107
rect 5104 27075 5136 27107
rect 5176 27075 5208 27107
rect 5248 27075 5280 27107
rect 5320 27075 5352 27107
rect 5392 27075 5424 27107
rect 5464 27075 5496 27107
rect 5536 27075 5568 27107
rect 5608 27075 5640 27107
rect 5680 27075 5712 27107
rect 5752 27075 5784 27107
rect 5824 27075 5856 27107
rect 5896 27075 5928 27107
rect 5968 27075 6000 27107
rect 6040 27075 6072 27107
rect 6112 27075 6144 27107
rect 6184 27075 6216 27107
rect 6256 27075 6288 27107
rect 6328 27075 6360 27107
rect 6400 27075 6432 27107
rect 6472 27075 6504 27107
rect 6544 27075 6576 27107
rect 6616 27075 6648 27107
rect 6688 27075 6720 27107
rect 6760 27075 6792 27107
rect 6832 27075 6864 27107
rect 6904 27075 6936 27107
rect 6976 27075 7008 27107
rect 7048 27075 7080 27107
rect 7120 27075 7152 27107
rect 7192 27075 7224 27107
rect 7264 27075 7296 27107
rect 7336 27075 7368 27107
rect 7408 27075 7440 27107
rect 7480 27075 7512 27107
rect 7552 27075 7584 27107
rect 7624 27075 7656 27107
rect 7696 27075 7728 27107
rect 7768 27075 7800 27107
rect 7840 27075 7872 27107
rect 7912 27075 7944 27107
rect 7984 27075 8016 27107
rect 8056 27075 8088 27107
rect 8128 27075 8160 27107
rect 8200 27075 8232 27107
rect 8272 27075 8304 27107
rect 8344 27075 8376 27107
rect 8416 27075 8448 27107
rect 8488 27075 8520 27107
rect 8560 27075 8592 27107
rect 8632 27075 8664 27107
rect 8704 27075 8736 27107
rect 8776 27075 8808 27107
rect 8848 27075 8880 27107
rect 8920 27075 8952 27107
rect 8992 27075 9024 27107
rect 9064 27075 9096 27107
rect 9136 27075 9168 27107
rect 9208 27075 9240 27107
rect 9280 27075 9312 27107
rect 9352 27075 9384 27107
rect 9424 27075 9456 27107
rect 9496 27075 9528 27107
rect 9568 27075 9600 27107
rect 9640 27075 9672 27107
rect 9712 27075 9744 27107
rect 9784 27075 9816 27107
rect 9856 27075 9888 27107
rect 9928 27075 9960 27107
rect 10000 27075 10032 27107
rect 10072 27075 10104 27107
rect 10144 27075 10176 27107
rect 10216 27075 10248 27107
rect 10288 27075 10320 27107
rect 10360 27075 10392 27107
rect 10432 27075 10464 27107
rect 10504 27075 10536 27107
rect 10576 27075 10608 27107
rect 10648 27075 10680 27107
rect 10720 27075 10752 27107
rect 10792 27075 10824 27107
rect 10864 27075 10896 27107
rect 10936 27075 10968 27107
rect 11008 27075 11040 27107
rect 11080 27075 11112 27107
rect 11152 27075 11184 27107
rect 11224 27075 11256 27107
rect 11296 27075 11328 27107
rect 11368 27075 11400 27107
rect 11440 27075 11472 27107
rect 11512 27075 11544 27107
rect 11584 27075 11616 27107
rect 11656 27075 11688 27107
rect 11728 27075 11760 27107
rect 11800 27075 11832 27107
rect 11872 27075 11904 27107
rect 11944 27075 11976 27107
rect 12016 27075 12048 27107
rect 12088 27075 12120 27107
rect 12160 27075 12192 27107
rect 12232 27075 12264 27107
rect 12304 27075 12336 27107
rect 12376 27075 12408 27107
rect 12448 27075 12480 27107
rect 12520 27075 12552 27107
rect 12592 27075 12624 27107
rect 12664 27075 12696 27107
rect 12736 27075 12768 27107
rect 12808 27075 12840 27107
rect 12880 27075 12912 27107
rect 12952 27075 12984 27107
rect 13024 27075 13056 27107
rect 13096 27075 13128 27107
rect 13168 27075 13200 27107
rect 13240 27075 13272 27107
rect 13312 27075 13344 27107
rect 13384 27075 13416 27107
rect 13456 27075 13488 27107
rect 13528 27075 13560 27107
rect 13600 27075 13632 27107
rect 13672 27075 13704 27107
rect 13744 27075 13776 27107
rect 13816 27075 13848 27107
rect 13888 27075 13920 27107
rect 13960 27075 13992 27107
rect 14032 27075 14064 27107
rect 14104 27075 14136 27107
rect 14176 27075 14208 27107
rect 14248 27075 14280 27107
rect 14320 27075 14352 27107
rect 14392 27075 14424 27107
rect 14464 27075 14496 27107
rect 14536 27075 14568 27107
rect 14608 27075 14640 27107
rect 14680 27075 14712 27107
rect 14752 27075 14784 27107
rect 14824 27075 14856 27107
rect 14896 27075 14928 27107
rect 14968 27075 15000 27107
rect 15040 27075 15072 27107
rect 15112 27075 15144 27107
rect 15184 27075 15216 27107
rect 15256 27075 15288 27107
rect 15328 27075 15360 27107
rect 15400 27075 15432 27107
rect 15472 27075 15504 27107
rect 15544 27075 15576 27107
rect 15616 27075 15648 27107
rect 15688 27075 15720 27107
rect 15760 27075 15792 27107
rect 15832 27075 15864 27107
rect 15904 27075 15936 27107
rect 64 27003 96 27035
rect 136 27003 168 27035
rect 208 27003 240 27035
rect 280 27003 312 27035
rect 352 27003 384 27035
rect 424 27003 456 27035
rect 496 27003 528 27035
rect 568 27003 600 27035
rect 640 27003 672 27035
rect 712 27003 744 27035
rect 784 27003 816 27035
rect 856 27003 888 27035
rect 928 27003 960 27035
rect 1000 27003 1032 27035
rect 1072 27003 1104 27035
rect 1144 27003 1176 27035
rect 1216 27003 1248 27035
rect 1288 27003 1320 27035
rect 1360 27003 1392 27035
rect 1432 27003 1464 27035
rect 1504 27003 1536 27035
rect 1576 27003 1608 27035
rect 1648 27003 1680 27035
rect 1720 27003 1752 27035
rect 1792 27003 1824 27035
rect 1864 27003 1896 27035
rect 1936 27003 1968 27035
rect 2008 27003 2040 27035
rect 2080 27003 2112 27035
rect 2152 27003 2184 27035
rect 2224 27003 2256 27035
rect 2296 27003 2328 27035
rect 2368 27003 2400 27035
rect 2440 27003 2472 27035
rect 2512 27003 2544 27035
rect 2584 27003 2616 27035
rect 2656 27003 2688 27035
rect 2728 27003 2760 27035
rect 2800 27003 2832 27035
rect 2872 27003 2904 27035
rect 2944 27003 2976 27035
rect 3016 27003 3048 27035
rect 3088 27003 3120 27035
rect 3160 27003 3192 27035
rect 3232 27003 3264 27035
rect 3304 27003 3336 27035
rect 3376 27003 3408 27035
rect 3448 27003 3480 27035
rect 3520 27003 3552 27035
rect 3592 27003 3624 27035
rect 3664 27003 3696 27035
rect 3736 27003 3768 27035
rect 3808 27003 3840 27035
rect 3880 27003 3912 27035
rect 3952 27003 3984 27035
rect 4024 27003 4056 27035
rect 4096 27003 4128 27035
rect 4168 27003 4200 27035
rect 4240 27003 4272 27035
rect 4312 27003 4344 27035
rect 4384 27003 4416 27035
rect 4456 27003 4488 27035
rect 4528 27003 4560 27035
rect 4600 27003 4632 27035
rect 4672 27003 4704 27035
rect 4744 27003 4776 27035
rect 4816 27003 4848 27035
rect 4888 27003 4920 27035
rect 4960 27003 4992 27035
rect 5032 27003 5064 27035
rect 5104 27003 5136 27035
rect 5176 27003 5208 27035
rect 5248 27003 5280 27035
rect 5320 27003 5352 27035
rect 5392 27003 5424 27035
rect 5464 27003 5496 27035
rect 5536 27003 5568 27035
rect 5608 27003 5640 27035
rect 5680 27003 5712 27035
rect 5752 27003 5784 27035
rect 5824 27003 5856 27035
rect 5896 27003 5928 27035
rect 5968 27003 6000 27035
rect 6040 27003 6072 27035
rect 6112 27003 6144 27035
rect 6184 27003 6216 27035
rect 6256 27003 6288 27035
rect 6328 27003 6360 27035
rect 6400 27003 6432 27035
rect 6472 27003 6504 27035
rect 6544 27003 6576 27035
rect 6616 27003 6648 27035
rect 6688 27003 6720 27035
rect 6760 27003 6792 27035
rect 6832 27003 6864 27035
rect 6904 27003 6936 27035
rect 6976 27003 7008 27035
rect 7048 27003 7080 27035
rect 7120 27003 7152 27035
rect 7192 27003 7224 27035
rect 7264 27003 7296 27035
rect 7336 27003 7368 27035
rect 7408 27003 7440 27035
rect 7480 27003 7512 27035
rect 7552 27003 7584 27035
rect 7624 27003 7656 27035
rect 7696 27003 7728 27035
rect 7768 27003 7800 27035
rect 7840 27003 7872 27035
rect 7912 27003 7944 27035
rect 7984 27003 8016 27035
rect 8056 27003 8088 27035
rect 8128 27003 8160 27035
rect 8200 27003 8232 27035
rect 8272 27003 8304 27035
rect 8344 27003 8376 27035
rect 8416 27003 8448 27035
rect 8488 27003 8520 27035
rect 8560 27003 8592 27035
rect 8632 27003 8664 27035
rect 8704 27003 8736 27035
rect 8776 27003 8808 27035
rect 8848 27003 8880 27035
rect 8920 27003 8952 27035
rect 8992 27003 9024 27035
rect 9064 27003 9096 27035
rect 9136 27003 9168 27035
rect 9208 27003 9240 27035
rect 9280 27003 9312 27035
rect 9352 27003 9384 27035
rect 9424 27003 9456 27035
rect 9496 27003 9528 27035
rect 9568 27003 9600 27035
rect 9640 27003 9672 27035
rect 9712 27003 9744 27035
rect 9784 27003 9816 27035
rect 9856 27003 9888 27035
rect 9928 27003 9960 27035
rect 10000 27003 10032 27035
rect 10072 27003 10104 27035
rect 10144 27003 10176 27035
rect 10216 27003 10248 27035
rect 10288 27003 10320 27035
rect 10360 27003 10392 27035
rect 10432 27003 10464 27035
rect 10504 27003 10536 27035
rect 10576 27003 10608 27035
rect 10648 27003 10680 27035
rect 10720 27003 10752 27035
rect 10792 27003 10824 27035
rect 10864 27003 10896 27035
rect 10936 27003 10968 27035
rect 11008 27003 11040 27035
rect 11080 27003 11112 27035
rect 11152 27003 11184 27035
rect 11224 27003 11256 27035
rect 11296 27003 11328 27035
rect 11368 27003 11400 27035
rect 11440 27003 11472 27035
rect 11512 27003 11544 27035
rect 11584 27003 11616 27035
rect 11656 27003 11688 27035
rect 11728 27003 11760 27035
rect 11800 27003 11832 27035
rect 11872 27003 11904 27035
rect 11944 27003 11976 27035
rect 12016 27003 12048 27035
rect 12088 27003 12120 27035
rect 12160 27003 12192 27035
rect 12232 27003 12264 27035
rect 12304 27003 12336 27035
rect 12376 27003 12408 27035
rect 12448 27003 12480 27035
rect 12520 27003 12552 27035
rect 12592 27003 12624 27035
rect 12664 27003 12696 27035
rect 12736 27003 12768 27035
rect 12808 27003 12840 27035
rect 12880 27003 12912 27035
rect 12952 27003 12984 27035
rect 13024 27003 13056 27035
rect 13096 27003 13128 27035
rect 13168 27003 13200 27035
rect 13240 27003 13272 27035
rect 13312 27003 13344 27035
rect 13384 27003 13416 27035
rect 13456 27003 13488 27035
rect 13528 27003 13560 27035
rect 13600 27003 13632 27035
rect 13672 27003 13704 27035
rect 13744 27003 13776 27035
rect 13816 27003 13848 27035
rect 13888 27003 13920 27035
rect 13960 27003 13992 27035
rect 14032 27003 14064 27035
rect 14104 27003 14136 27035
rect 14176 27003 14208 27035
rect 14248 27003 14280 27035
rect 14320 27003 14352 27035
rect 14392 27003 14424 27035
rect 14464 27003 14496 27035
rect 14536 27003 14568 27035
rect 14608 27003 14640 27035
rect 14680 27003 14712 27035
rect 14752 27003 14784 27035
rect 14824 27003 14856 27035
rect 14896 27003 14928 27035
rect 14968 27003 15000 27035
rect 15040 27003 15072 27035
rect 15112 27003 15144 27035
rect 15184 27003 15216 27035
rect 15256 27003 15288 27035
rect 15328 27003 15360 27035
rect 15400 27003 15432 27035
rect 15472 27003 15504 27035
rect 15544 27003 15576 27035
rect 15616 27003 15648 27035
rect 15688 27003 15720 27035
rect 15760 27003 15792 27035
rect 15832 27003 15864 27035
rect 15904 27003 15936 27035
rect 64 26931 96 26963
rect 136 26931 168 26963
rect 208 26931 240 26963
rect 280 26931 312 26963
rect 352 26931 384 26963
rect 424 26931 456 26963
rect 496 26931 528 26963
rect 568 26931 600 26963
rect 640 26931 672 26963
rect 712 26931 744 26963
rect 784 26931 816 26963
rect 856 26931 888 26963
rect 928 26931 960 26963
rect 1000 26931 1032 26963
rect 1072 26931 1104 26963
rect 1144 26931 1176 26963
rect 1216 26931 1248 26963
rect 1288 26931 1320 26963
rect 1360 26931 1392 26963
rect 1432 26931 1464 26963
rect 1504 26931 1536 26963
rect 1576 26931 1608 26963
rect 1648 26931 1680 26963
rect 1720 26931 1752 26963
rect 1792 26931 1824 26963
rect 1864 26931 1896 26963
rect 1936 26931 1968 26963
rect 2008 26931 2040 26963
rect 2080 26931 2112 26963
rect 2152 26931 2184 26963
rect 2224 26931 2256 26963
rect 2296 26931 2328 26963
rect 2368 26931 2400 26963
rect 2440 26931 2472 26963
rect 2512 26931 2544 26963
rect 2584 26931 2616 26963
rect 2656 26931 2688 26963
rect 2728 26931 2760 26963
rect 2800 26931 2832 26963
rect 2872 26931 2904 26963
rect 2944 26931 2976 26963
rect 3016 26931 3048 26963
rect 3088 26931 3120 26963
rect 3160 26931 3192 26963
rect 3232 26931 3264 26963
rect 3304 26931 3336 26963
rect 3376 26931 3408 26963
rect 3448 26931 3480 26963
rect 3520 26931 3552 26963
rect 3592 26931 3624 26963
rect 3664 26931 3696 26963
rect 3736 26931 3768 26963
rect 3808 26931 3840 26963
rect 3880 26931 3912 26963
rect 3952 26931 3984 26963
rect 4024 26931 4056 26963
rect 4096 26931 4128 26963
rect 4168 26931 4200 26963
rect 4240 26931 4272 26963
rect 4312 26931 4344 26963
rect 4384 26931 4416 26963
rect 4456 26931 4488 26963
rect 4528 26931 4560 26963
rect 4600 26931 4632 26963
rect 4672 26931 4704 26963
rect 4744 26931 4776 26963
rect 4816 26931 4848 26963
rect 4888 26931 4920 26963
rect 4960 26931 4992 26963
rect 5032 26931 5064 26963
rect 5104 26931 5136 26963
rect 5176 26931 5208 26963
rect 5248 26931 5280 26963
rect 5320 26931 5352 26963
rect 5392 26931 5424 26963
rect 5464 26931 5496 26963
rect 5536 26931 5568 26963
rect 5608 26931 5640 26963
rect 5680 26931 5712 26963
rect 5752 26931 5784 26963
rect 5824 26931 5856 26963
rect 5896 26931 5928 26963
rect 5968 26931 6000 26963
rect 6040 26931 6072 26963
rect 6112 26931 6144 26963
rect 6184 26931 6216 26963
rect 6256 26931 6288 26963
rect 6328 26931 6360 26963
rect 6400 26931 6432 26963
rect 6472 26931 6504 26963
rect 6544 26931 6576 26963
rect 6616 26931 6648 26963
rect 6688 26931 6720 26963
rect 6760 26931 6792 26963
rect 6832 26931 6864 26963
rect 6904 26931 6936 26963
rect 6976 26931 7008 26963
rect 7048 26931 7080 26963
rect 7120 26931 7152 26963
rect 7192 26931 7224 26963
rect 7264 26931 7296 26963
rect 7336 26931 7368 26963
rect 7408 26931 7440 26963
rect 7480 26931 7512 26963
rect 7552 26931 7584 26963
rect 7624 26931 7656 26963
rect 7696 26931 7728 26963
rect 7768 26931 7800 26963
rect 7840 26931 7872 26963
rect 7912 26931 7944 26963
rect 7984 26931 8016 26963
rect 8056 26931 8088 26963
rect 8128 26931 8160 26963
rect 8200 26931 8232 26963
rect 8272 26931 8304 26963
rect 8344 26931 8376 26963
rect 8416 26931 8448 26963
rect 8488 26931 8520 26963
rect 8560 26931 8592 26963
rect 8632 26931 8664 26963
rect 8704 26931 8736 26963
rect 8776 26931 8808 26963
rect 8848 26931 8880 26963
rect 8920 26931 8952 26963
rect 8992 26931 9024 26963
rect 9064 26931 9096 26963
rect 9136 26931 9168 26963
rect 9208 26931 9240 26963
rect 9280 26931 9312 26963
rect 9352 26931 9384 26963
rect 9424 26931 9456 26963
rect 9496 26931 9528 26963
rect 9568 26931 9600 26963
rect 9640 26931 9672 26963
rect 9712 26931 9744 26963
rect 9784 26931 9816 26963
rect 9856 26931 9888 26963
rect 9928 26931 9960 26963
rect 10000 26931 10032 26963
rect 10072 26931 10104 26963
rect 10144 26931 10176 26963
rect 10216 26931 10248 26963
rect 10288 26931 10320 26963
rect 10360 26931 10392 26963
rect 10432 26931 10464 26963
rect 10504 26931 10536 26963
rect 10576 26931 10608 26963
rect 10648 26931 10680 26963
rect 10720 26931 10752 26963
rect 10792 26931 10824 26963
rect 10864 26931 10896 26963
rect 10936 26931 10968 26963
rect 11008 26931 11040 26963
rect 11080 26931 11112 26963
rect 11152 26931 11184 26963
rect 11224 26931 11256 26963
rect 11296 26931 11328 26963
rect 11368 26931 11400 26963
rect 11440 26931 11472 26963
rect 11512 26931 11544 26963
rect 11584 26931 11616 26963
rect 11656 26931 11688 26963
rect 11728 26931 11760 26963
rect 11800 26931 11832 26963
rect 11872 26931 11904 26963
rect 11944 26931 11976 26963
rect 12016 26931 12048 26963
rect 12088 26931 12120 26963
rect 12160 26931 12192 26963
rect 12232 26931 12264 26963
rect 12304 26931 12336 26963
rect 12376 26931 12408 26963
rect 12448 26931 12480 26963
rect 12520 26931 12552 26963
rect 12592 26931 12624 26963
rect 12664 26931 12696 26963
rect 12736 26931 12768 26963
rect 12808 26931 12840 26963
rect 12880 26931 12912 26963
rect 12952 26931 12984 26963
rect 13024 26931 13056 26963
rect 13096 26931 13128 26963
rect 13168 26931 13200 26963
rect 13240 26931 13272 26963
rect 13312 26931 13344 26963
rect 13384 26931 13416 26963
rect 13456 26931 13488 26963
rect 13528 26931 13560 26963
rect 13600 26931 13632 26963
rect 13672 26931 13704 26963
rect 13744 26931 13776 26963
rect 13816 26931 13848 26963
rect 13888 26931 13920 26963
rect 13960 26931 13992 26963
rect 14032 26931 14064 26963
rect 14104 26931 14136 26963
rect 14176 26931 14208 26963
rect 14248 26931 14280 26963
rect 14320 26931 14352 26963
rect 14392 26931 14424 26963
rect 14464 26931 14496 26963
rect 14536 26931 14568 26963
rect 14608 26931 14640 26963
rect 14680 26931 14712 26963
rect 14752 26931 14784 26963
rect 14824 26931 14856 26963
rect 14896 26931 14928 26963
rect 14968 26931 15000 26963
rect 15040 26931 15072 26963
rect 15112 26931 15144 26963
rect 15184 26931 15216 26963
rect 15256 26931 15288 26963
rect 15328 26931 15360 26963
rect 15400 26931 15432 26963
rect 15472 26931 15504 26963
rect 15544 26931 15576 26963
rect 15616 26931 15648 26963
rect 15688 26931 15720 26963
rect 15760 26931 15792 26963
rect 15832 26931 15864 26963
rect 15904 26931 15936 26963
rect 64 26859 96 26891
rect 136 26859 168 26891
rect 208 26859 240 26891
rect 280 26859 312 26891
rect 352 26859 384 26891
rect 424 26859 456 26891
rect 496 26859 528 26891
rect 568 26859 600 26891
rect 640 26859 672 26891
rect 712 26859 744 26891
rect 784 26859 816 26891
rect 856 26859 888 26891
rect 928 26859 960 26891
rect 1000 26859 1032 26891
rect 1072 26859 1104 26891
rect 1144 26859 1176 26891
rect 1216 26859 1248 26891
rect 1288 26859 1320 26891
rect 1360 26859 1392 26891
rect 1432 26859 1464 26891
rect 1504 26859 1536 26891
rect 1576 26859 1608 26891
rect 1648 26859 1680 26891
rect 1720 26859 1752 26891
rect 1792 26859 1824 26891
rect 1864 26859 1896 26891
rect 1936 26859 1968 26891
rect 2008 26859 2040 26891
rect 2080 26859 2112 26891
rect 2152 26859 2184 26891
rect 2224 26859 2256 26891
rect 2296 26859 2328 26891
rect 2368 26859 2400 26891
rect 2440 26859 2472 26891
rect 2512 26859 2544 26891
rect 2584 26859 2616 26891
rect 2656 26859 2688 26891
rect 2728 26859 2760 26891
rect 2800 26859 2832 26891
rect 2872 26859 2904 26891
rect 2944 26859 2976 26891
rect 3016 26859 3048 26891
rect 3088 26859 3120 26891
rect 3160 26859 3192 26891
rect 3232 26859 3264 26891
rect 3304 26859 3336 26891
rect 3376 26859 3408 26891
rect 3448 26859 3480 26891
rect 3520 26859 3552 26891
rect 3592 26859 3624 26891
rect 3664 26859 3696 26891
rect 3736 26859 3768 26891
rect 3808 26859 3840 26891
rect 3880 26859 3912 26891
rect 3952 26859 3984 26891
rect 4024 26859 4056 26891
rect 4096 26859 4128 26891
rect 4168 26859 4200 26891
rect 4240 26859 4272 26891
rect 4312 26859 4344 26891
rect 4384 26859 4416 26891
rect 4456 26859 4488 26891
rect 4528 26859 4560 26891
rect 4600 26859 4632 26891
rect 4672 26859 4704 26891
rect 4744 26859 4776 26891
rect 4816 26859 4848 26891
rect 4888 26859 4920 26891
rect 4960 26859 4992 26891
rect 5032 26859 5064 26891
rect 5104 26859 5136 26891
rect 5176 26859 5208 26891
rect 5248 26859 5280 26891
rect 5320 26859 5352 26891
rect 5392 26859 5424 26891
rect 5464 26859 5496 26891
rect 5536 26859 5568 26891
rect 5608 26859 5640 26891
rect 5680 26859 5712 26891
rect 5752 26859 5784 26891
rect 5824 26859 5856 26891
rect 5896 26859 5928 26891
rect 5968 26859 6000 26891
rect 6040 26859 6072 26891
rect 6112 26859 6144 26891
rect 6184 26859 6216 26891
rect 6256 26859 6288 26891
rect 6328 26859 6360 26891
rect 6400 26859 6432 26891
rect 6472 26859 6504 26891
rect 6544 26859 6576 26891
rect 6616 26859 6648 26891
rect 6688 26859 6720 26891
rect 6760 26859 6792 26891
rect 6832 26859 6864 26891
rect 6904 26859 6936 26891
rect 6976 26859 7008 26891
rect 7048 26859 7080 26891
rect 7120 26859 7152 26891
rect 7192 26859 7224 26891
rect 7264 26859 7296 26891
rect 7336 26859 7368 26891
rect 7408 26859 7440 26891
rect 7480 26859 7512 26891
rect 7552 26859 7584 26891
rect 7624 26859 7656 26891
rect 7696 26859 7728 26891
rect 7768 26859 7800 26891
rect 7840 26859 7872 26891
rect 7912 26859 7944 26891
rect 7984 26859 8016 26891
rect 8056 26859 8088 26891
rect 8128 26859 8160 26891
rect 8200 26859 8232 26891
rect 8272 26859 8304 26891
rect 8344 26859 8376 26891
rect 8416 26859 8448 26891
rect 8488 26859 8520 26891
rect 8560 26859 8592 26891
rect 8632 26859 8664 26891
rect 8704 26859 8736 26891
rect 8776 26859 8808 26891
rect 8848 26859 8880 26891
rect 8920 26859 8952 26891
rect 8992 26859 9024 26891
rect 9064 26859 9096 26891
rect 9136 26859 9168 26891
rect 9208 26859 9240 26891
rect 9280 26859 9312 26891
rect 9352 26859 9384 26891
rect 9424 26859 9456 26891
rect 9496 26859 9528 26891
rect 9568 26859 9600 26891
rect 9640 26859 9672 26891
rect 9712 26859 9744 26891
rect 9784 26859 9816 26891
rect 9856 26859 9888 26891
rect 9928 26859 9960 26891
rect 10000 26859 10032 26891
rect 10072 26859 10104 26891
rect 10144 26859 10176 26891
rect 10216 26859 10248 26891
rect 10288 26859 10320 26891
rect 10360 26859 10392 26891
rect 10432 26859 10464 26891
rect 10504 26859 10536 26891
rect 10576 26859 10608 26891
rect 10648 26859 10680 26891
rect 10720 26859 10752 26891
rect 10792 26859 10824 26891
rect 10864 26859 10896 26891
rect 10936 26859 10968 26891
rect 11008 26859 11040 26891
rect 11080 26859 11112 26891
rect 11152 26859 11184 26891
rect 11224 26859 11256 26891
rect 11296 26859 11328 26891
rect 11368 26859 11400 26891
rect 11440 26859 11472 26891
rect 11512 26859 11544 26891
rect 11584 26859 11616 26891
rect 11656 26859 11688 26891
rect 11728 26859 11760 26891
rect 11800 26859 11832 26891
rect 11872 26859 11904 26891
rect 11944 26859 11976 26891
rect 12016 26859 12048 26891
rect 12088 26859 12120 26891
rect 12160 26859 12192 26891
rect 12232 26859 12264 26891
rect 12304 26859 12336 26891
rect 12376 26859 12408 26891
rect 12448 26859 12480 26891
rect 12520 26859 12552 26891
rect 12592 26859 12624 26891
rect 12664 26859 12696 26891
rect 12736 26859 12768 26891
rect 12808 26859 12840 26891
rect 12880 26859 12912 26891
rect 12952 26859 12984 26891
rect 13024 26859 13056 26891
rect 13096 26859 13128 26891
rect 13168 26859 13200 26891
rect 13240 26859 13272 26891
rect 13312 26859 13344 26891
rect 13384 26859 13416 26891
rect 13456 26859 13488 26891
rect 13528 26859 13560 26891
rect 13600 26859 13632 26891
rect 13672 26859 13704 26891
rect 13744 26859 13776 26891
rect 13816 26859 13848 26891
rect 13888 26859 13920 26891
rect 13960 26859 13992 26891
rect 14032 26859 14064 26891
rect 14104 26859 14136 26891
rect 14176 26859 14208 26891
rect 14248 26859 14280 26891
rect 14320 26859 14352 26891
rect 14392 26859 14424 26891
rect 14464 26859 14496 26891
rect 14536 26859 14568 26891
rect 14608 26859 14640 26891
rect 14680 26859 14712 26891
rect 14752 26859 14784 26891
rect 14824 26859 14856 26891
rect 14896 26859 14928 26891
rect 14968 26859 15000 26891
rect 15040 26859 15072 26891
rect 15112 26859 15144 26891
rect 15184 26859 15216 26891
rect 15256 26859 15288 26891
rect 15328 26859 15360 26891
rect 15400 26859 15432 26891
rect 15472 26859 15504 26891
rect 15544 26859 15576 26891
rect 15616 26859 15648 26891
rect 15688 26859 15720 26891
rect 15760 26859 15792 26891
rect 15832 26859 15864 26891
rect 15904 26859 15936 26891
rect 64 26787 96 26819
rect 136 26787 168 26819
rect 208 26787 240 26819
rect 280 26787 312 26819
rect 352 26787 384 26819
rect 424 26787 456 26819
rect 496 26787 528 26819
rect 568 26787 600 26819
rect 640 26787 672 26819
rect 712 26787 744 26819
rect 784 26787 816 26819
rect 856 26787 888 26819
rect 928 26787 960 26819
rect 1000 26787 1032 26819
rect 1072 26787 1104 26819
rect 1144 26787 1176 26819
rect 1216 26787 1248 26819
rect 1288 26787 1320 26819
rect 1360 26787 1392 26819
rect 1432 26787 1464 26819
rect 1504 26787 1536 26819
rect 1576 26787 1608 26819
rect 1648 26787 1680 26819
rect 1720 26787 1752 26819
rect 1792 26787 1824 26819
rect 1864 26787 1896 26819
rect 1936 26787 1968 26819
rect 2008 26787 2040 26819
rect 2080 26787 2112 26819
rect 2152 26787 2184 26819
rect 2224 26787 2256 26819
rect 2296 26787 2328 26819
rect 2368 26787 2400 26819
rect 2440 26787 2472 26819
rect 2512 26787 2544 26819
rect 2584 26787 2616 26819
rect 2656 26787 2688 26819
rect 2728 26787 2760 26819
rect 2800 26787 2832 26819
rect 2872 26787 2904 26819
rect 2944 26787 2976 26819
rect 3016 26787 3048 26819
rect 3088 26787 3120 26819
rect 3160 26787 3192 26819
rect 3232 26787 3264 26819
rect 3304 26787 3336 26819
rect 3376 26787 3408 26819
rect 3448 26787 3480 26819
rect 3520 26787 3552 26819
rect 3592 26787 3624 26819
rect 3664 26787 3696 26819
rect 3736 26787 3768 26819
rect 3808 26787 3840 26819
rect 3880 26787 3912 26819
rect 3952 26787 3984 26819
rect 4024 26787 4056 26819
rect 4096 26787 4128 26819
rect 4168 26787 4200 26819
rect 4240 26787 4272 26819
rect 4312 26787 4344 26819
rect 4384 26787 4416 26819
rect 4456 26787 4488 26819
rect 4528 26787 4560 26819
rect 4600 26787 4632 26819
rect 4672 26787 4704 26819
rect 4744 26787 4776 26819
rect 4816 26787 4848 26819
rect 4888 26787 4920 26819
rect 4960 26787 4992 26819
rect 5032 26787 5064 26819
rect 5104 26787 5136 26819
rect 5176 26787 5208 26819
rect 5248 26787 5280 26819
rect 5320 26787 5352 26819
rect 5392 26787 5424 26819
rect 5464 26787 5496 26819
rect 5536 26787 5568 26819
rect 5608 26787 5640 26819
rect 5680 26787 5712 26819
rect 5752 26787 5784 26819
rect 5824 26787 5856 26819
rect 5896 26787 5928 26819
rect 5968 26787 6000 26819
rect 6040 26787 6072 26819
rect 6112 26787 6144 26819
rect 6184 26787 6216 26819
rect 6256 26787 6288 26819
rect 6328 26787 6360 26819
rect 6400 26787 6432 26819
rect 6472 26787 6504 26819
rect 6544 26787 6576 26819
rect 6616 26787 6648 26819
rect 6688 26787 6720 26819
rect 6760 26787 6792 26819
rect 6832 26787 6864 26819
rect 6904 26787 6936 26819
rect 6976 26787 7008 26819
rect 7048 26787 7080 26819
rect 7120 26787 7152 26819
rect 7192 26787 7224 26819
rect 7264 26787 7296 26819
rect 7336 26787 7368 26819
rect 7408 26787 7440 26819
rect 7480 26787 7512 26819
rect 7552 26787 7584 26819
rect 7624 26787 7656 26819
rect 7696 26787 7728 26819
rect 7768 26787 7800 26819
rect 7840 26787 7872 26819
rect 7912 26787 7944 26819
rect 7984 26787 8016 26819
rect 8056 26787 8088 26819
rect 8128 26787 8160 26819
rect 8200 26787 8232 26819
rect 8272 26787 8304 26819
rect 8344 26787 8376 26819
rect 8416 26787 8448 26819
rect 8488 26787 8520 26819
rect 8560 26787 8592 26819
rect 8632 26787 8664 26819
rect 8704 26787 8736 26819
rect 8776 26787 8808 26819
rect 8848 26787 8880 26819
rect 8920 26787 8952 26819
rect 8992 26787 9024 26819
rect 9064 26787 9096 26819
rect 9136 26787 9168 26819
rect 9208 26787 9240 26819
rect 9280 26787 9312 26819
rect 9352 26787 9384 26819
rect 9424 26787 9456 26819
rect 9496 26787 9528 26819
rect 9568 26787 9600 26819
rect 9640 26787 9672 26819
rect 9712 26787 9744 26819
rect 9784 26787 9816 26819
rect 9856 26787 9888 26819
rect 9928 26787 9960 26819
rect 10000 26787 10032 26819
rect 10072 26787 10104 26819
rect 10144 26787 10176 26819
rect 10216 26787 10248 26819
rect 10288 26787 10320 26819
rect 10360 26787 10392 26819
rect 10432 26787 10464 26819
rect 10504 26787 10536 26819
rect 10576 26787 10608 26819
rect 10648 26787 10680 26819
rect 10720 26787 10752 26819
rect 10792 26787 10824 26819
rect 10864 26787 10896 26819
rect 10936 26787 10968 26819
rect 11008 26787 11040 26819
rect 11080 26787 11112 26819
rect 11152 26787 11184 26819
rect 11224 26787 11256 26819
rect 11296 26787 11328 26819
rect 11368 26787 11400 26819
rect 11440 26787 11472 26819
rect 11512 26787 11544 26819
rect 11584 26787 11616 26819
rect 11656 26787 11688 26819
rect 11728 26787 11760 26819
rect 11800 26787 11832 26819
rect 11872 26787 11904 26819
rect 11944 26787 11976 26819
rect 12016 26787 12048 26819
rect 12088 26787 12120 26819
rect 12160 26787 12192 26819
rect 12232 26787 12264 26819
rect 12304 26787 12336 26819
rect 12376 26787 12408 26819
rect 12448 26787 12480 26819
rect 12520 26787 12552 26819
rect 12592 26787 12624 26819
rect 12664 26787 12696 26819
rect 12736 26787 12768 26819
rect 12808 26787 12840 26819
rect 12880 26787 12912 26819
rect 12952 26787 12984 26819
rect 13024 26787 13056 26819
rect 13096 26787 13128 26819
rect 13168 26787 13200 26819
rect 13240 26787 13272 26819
rect 13312 26787 13344 26819
rect 13384 26787 13416 26819
rect 13456 26787 13488 26819
rect 13528 26787 13560 26819
rect 13600 26787 13632 26819
rect 13672 26787 13704 26819
rect 13744 26787 13776 26819
rect 13816 26787 13848 26819
rect 13888 26787 13920 26819
rect 13960 26787 13992 26819
rect 14032 26787 14064 26819
rect 14104 26787 14136 26819
rect 14176 26787 14208 26819
rect 14248 26787 14280 26819
rect 14320 26787 14352 26819
rect 14392 26787 14424 26819
rect 14464 26787 14496 26819
rect 14536 26787 14568 26819
rect 14608 26787 14640 26819
rect 14680 26787 14712 26819
rect 14752 26787 14784 26819
rect 14824 26787 14856 26819
rect 14896 26787 14928 26819
rect 14968 26787 15000 26819
rect 15040 26787 15072 26819
rect 15112 26787 15144 26819
rect 15184 26787 15216 26819
rect 15256 26787 15288 26819
rect 15328 26787 15360 26819
rect 15400 26787 15432 26819
rect 15472 26787 15504 26819
rect 15544 26787 15576 26819
rect 15616 26787 15648 26819
rect 15688 26787 15720 26819
rect 15760 26787 15792 26819
rect 15832 26787 15864 26819
rect 15904 26787 15936 26819
rect 64 26715 96 26747
rect 136 26715 168 26747
rect 208 26715 240 26747
rect 280 26715 312 26747
rect 352 26715 384 26747
rect 424 26715 456 26747
rect 496 26715 528 26747
rect 568 26715 600 26747
rect 640 26715 672 26747
rect 712 26715 744 26747
rect 784 26715 816 26747
rect 856 26715 888 26747
rect 928 26715 960 26747
rect 1000 26715 1032 26747
rect 1072 26715 1104 26747
rect 1144 26715 1176 26747
rect 1216 26715 1248 26747
rect 1288 26715 1320 26747
rect 1360 26715 1392 26747
rect 1432 26715 1464 26747
rect 1504 26715 1536 26747
rect 1576 26715 1608 26747
rect 1648 26715 1680 26747
rect 1720 26715 1752 26747
rect 1792 26715 1824 26747
rect 1864 26715 1896 26747
rect 1936 26715 1968 26747
rect 2008 26715 2040 26747
rect 2080 26715 2112 26747
rect 2152 26715 2184 26747
rect 2224 26715 2256 26747
rect 2296 26715 2328 26747
rect 2368 26715 2400 26747
rect 2440 26715 2472 26747
rect 2512 26715 2544 26747
rect 2584 26715 2616 26747
rect 2656 26715 2688 26747
rect 2728 26715 2760 26747
rect 2800 26715 2832 26747
rect 2872 26715 2904 26747
rect 2944 26715 2976 26747
rect 3016 26715 3048 26747
rect 3088 26715 3120 26747
rect 3160 26715 3192 26747
rect 3232 26715 3264 26747
rect 3304 26715 3336 26747
rect 3376 26715 3408 26747
rect 3448 26715 3480 26747
rect 3520 26715 3552 26747
rect 3592 26715 3624 26747
rect 3664 26715 3696 26747
rect 3736 26715 3768 26747
rect 3808 26715 3840 26747
rect 3880 26715 3912 26747
rect 3952 26715 3984 26747
rect 4024 26715 4056 26747
rect 4096 26715 4128 26747
rect 4168 26715 4200 26747
rect 4240 26715 4272 26747
rect 4312 26715 4344 26747
rect 4384 26715 4416 26747
rect 4456 26715 4488 26747
rect 4528 26715 4560 26747
rect 4600 26715 4632 26747
rect 4672 26715 4704 26747
rect 4744 26715 4776 26747
rect 4816 26715 4848 26747
rect 4888 26715 4920 26747
rect 4960 26715 4992 26747
rect 5032 26715 5064 26747
rect 5104 26715 5136 26747
rect 5176 26715 5208 26747
rect 5248 26715 5280 26747
rect 5320 26715 5352 26747
rect 5392 26715 5424 26747
rect 5464 26715 5496 26747
rect 5536 26715 5568 26747
rect 5608 26715 5640 26747
rect 5680 26715 5712 26747
rect 5752 26715 5784 26747
rect 5824 26715 5856 26747
rect 5896 26715 5928 26747
rect 5968 26715 6000 26747
rect 6040 26715 6072 26747
rect 6112 26715 6144 26747
rect 6184 26715 6216 26747
rect 6256 26715 6288 26747
rect 6328 26715 6360 26747
rect 6400 26715 6432 26747
rect 6472 26715 6504 26747
rect 6544 26715 6576 26747
rect 6616 26715 6648 26747
rect 6688 26715 6720 26747
rect 6760 26715 6792 26747
rect 6832 26715 6864 26747
rect 6904 26715 6936 26747
rect 6976 26715 7008 26747
rect 7048 26715 7080 26747
rect 7120 26715 7152 26747
rect 7192 26715 7224 26747
rect 7264 26715 7296 26747
rect 7336 26715 7368 26747
rect 7408 26715 7440 26747
rect 7480 26715 7512 26747
rect 7552 26715 7584 26747
rect 7624 26715 7656 26747
rect 7696 26715 7728 26747
rect 7768 26715 7800 26747
rect 7840 26715 7872 26747
rect 7912 26715 7944 26747
rect 7984 26715 8016 26747
rect 8056 26715 8088 26747
rect 8128 26715 8160 26747
rect 8200 26715 8232 26747
rect 8272 26715 8304 26747
rect 8344 26715 8376 26747
rect 8416 26715 8448 26747
rect 8488 26715 8520 26747
rect 8560 26715 8592 26747
rect 8632 26715 8664 26747
rect 8704 26715 8736 26747
rect 8776 26715 8808 26747
rect 8848 26715 8880 26747
rect 8920 26715 8952 26747
rect 8992 26715 9024 26747
rect 9064 26715 9096 26747
rect 9136 26715 9168 26747
rect 9208 26715 9240 26747
rect 9280 26715 9312 26747
rect 9352 26715 9384 26747
rect 9424 26715 9456 26747
rect 9496 26715 9528 26747
rect 9568 26715 9600 26747
rect 9640 26715 9672 26747
rect 9712 26715 9744 26747
rect 9784 26715 9816 26747
rect 9856 26715 9888 26747
rect 9928 26715 9960 26747
rect 10000 26715 10032 26747
rect 10072 26715 10104 26747
rect 10144 26715 10176 26747
rect 10216 26715 10248 26747
rect 10288 26715 10320 26747
rect 10360 26715 10392 26747
rect 10432 26715 10464 26747
rect 10504 26715 10536 26747
rect 10576 26715 10608 26747
rect 10648 26715 10680 26747
rect 10720 26715 10752 26747
rect 10792 26715 10824 26747
rect 10864 26715 10896 26747
rect 10936 26715 10968 26747
rect 11008 26715 11040 26747
rect 11080 26715 11112 26747
rect 11152 26715 11184 26747
rect 11224 26715 11256 26747
rect 11296 26715 11328 26747
rect 11368 26715 11400 26747
rect 11440 26715 11472 26747
rect 11512 26715 11544 26747
rect 11584 26715 11616 26747
rect 11656 26715 11688 26747
rect 11728 26715 11760 26747
rect 11800 26715 11832 26747
rect 11872 26715 11904 26747
rect 11944 26715 11976 26747
rect 12016 26715 12048 26747
rect 12088 26715 12120 26747
rect 12160 26715 12192 26747
rect 12232 26715 12264 26747
rect 12304 26715 12336 26747
rect 12376 26715 12408 26747
rect 12448 26715 12480 26747
rect 12520 26715 12552 26747
rect 12592 26715 12624 26747
rect 12664 26715 12696 26747
rect 12736 26715 12768 26747
rect 12808 26715 12840 26747
rect 12880 26715 12912 26747
rect 12952 26715 12984 26747
rect 13024 26715 13056 26747
rect 13096 26715 13128 26747
rect 13168 26715 13200 26747
rect 13240 26715 13272 26747
rect 13312 26715 13344 26747
rect 13384 26715 13416 26747
rect 13456 26715 13488 26747
rect 13528 26715 13560 26747
rect 13600 26715 13632 26747
rect 13672 26715 13704 26747
rect 13744 26715 13776 26747
rect 13816 26715 13848 26747
rect 13888 26715 13920 26747
rect 13960 26715 13992 26747
rect 14032 26715 14064 26747
rect 14104 26715 14136 26747
rect 14176 26715 14208 26747
rect 14248 26715 14280 26747
rect 14320 26715 14352 26747
rect 14392 26715 14424 26747
rect 14464 26715 14496 26747
rect 14536 26715 14568 26747
rect 14608 26715 14640 26747
rect 14680 26715 14712 26747
rect 14752 26715 14784 26747
rect 14824 26715 14856 26747
rect 14896 26715 14928 26747
rect 14968 26715 15000 26747
rect 15040 26715 15072 26747
rect 15112 26715 15144 26747
rect 15184 26715 15216 26747
rect 15256 26715 15288 26747
rect 15328 26715 15360 26747
rect 15400 26715 15432 26747
rect 15472 26715 15504 26747
rect 15544 26715 15576 26747
rect 15616 26715 15648 26747
rect 15688 26715 15720 26747
rect 15760 26715 15792 26747
rect 15832 26715 15864 26747
rect 15904 26715 15936 26747
rect 64 26643 96 26675
rect 136 26643 168 26675
rect 208 26643 240 26675
rect 280 26643 312 26675
rect 352 26643 384 26675
rect 424 26643 456 26675
rect 496 26643 528 26675
rect 568 26643 600 26675
rect 640 26643 672 26675
rect 712 26643 744 26675
rect 784 26643 816 26675
rect 856 26643 888 26675
rect 928 26643 960 26675
rect 1000 26643 1032 26675
rect 1072 26643 1104 26675
rect 1144 26643 1176 26675
rect 1216 26643 1248 26675
rect 1288 26643 1320 26675
rect 1360 26643 1392 26675
rect 1432 26643 1464 26675
rect 1504 26643 1536 26675
rect 1576 26643 1608 26675
rect 1648 26643 1680 26675
rect 1720 26643 1752 26675
rect 1792 26643 1824 26675
rect 1864 26643 1896 26675
rect 1936 26643 1968 26675
rect 2008 26643 2040 26675
rect 2080 26643 2112 26675
rect 2152 26643 2184 26675
rect 2224 26643 2256 26675
rect 2296 26643 2328 26675
rect 2368 26643 2400 26675
rect 2440 26643 2472 26675
rect 2512 26643 2544 26675
rect 2584 26643 2616 26675
rect 2656 26643 2688 26675
rect 2728 26643 2760 26675
rect 2800 26643 2832 26675
rect 2872 26643 2904 26675
rect 2944 26643 2976 26675
rect 3016 26643 3048 26675
rect 3088 26643 3120 26675
rect 3160 26643 3192 26675
rect 3232 26643 3264 26675
rect 3304 26643 3336 26675
rect 3376 26643 3408 26675
rect 3448 26643 3480 26675
rect 3520 26643 3552 26675
rect 3592 26643 3624 26675
rect 3664 26643 3696 26675
rect 3736 26643 3768 26675
rect 3808 26643 3840 26675
rect 3880 26643 3912 26675
rect 3952 26643 3984 26675
rect 4024 26643 4056 26675
rect 4096 26643 4128 26675
rect 4168 26643 4200 26675
rect 4240 26643 4272 26675
rect 4312 26643 4344 26675
rect 4384 26643 4416 26675
rect 4456 26643 4488 26675
rect 4528 26643 4560 26675
rect 4600 26643 4632 26675
rect 4672 26643 4704 26675
rect 4744 26643 4776 26675
rect 4816 26643 4848 26675
rect 4888 26643 4920 26675
rect 4960 26643 4992 26675
rect 5032 26643 5064 26675
rect 5104 26643 5136 26675
rect 5176 26643 5208 26675
rect 5248 26643 5280 26675
rect 5320 26643 5352 26675
rect 5392 26643 5424 26675
rect 5464 26643 5496 26675
rect 5536 26643 5568 26675
rect 5608 26643 5640 26675
rect 5680 26643 5712 26675
rect 5752 26643 5784 26675
rect 5824 26643 5856 26675
rect 5896 26643 5928 26675
rect 5968 26643 6000 26675
rect 6040 26643 6072 26675
rect 6112 26643 6144 26675
rect 6184 26643 6216 26675
rect 6256 26643 6288 26675
rect 6328 26643 6360 26675
rect 6400 26643 6432 26675
rect 6472 26643 6504 26675
rect 6544 26643 6576 26675
rect 6616 26643 6648 26675
rect 6688 26643 6720 26675
rect 6760 26643 6792 26675
rect 6832 26643 6864 26675
rect 6904 26643 6936 26675
rect 6976 26643 7008 26675
rect 7048 26643 7080 26675
rect 7120 26643 7152 26675
rect 7192 26643 7224 26675
rect 7264 26643 7296 26675
rect 7336 26643 7368 26675
rect 7408 26643 7440 26675
rect 7480 26643 7512 26675
rect 7552 26643 7584 26675
rect 7624 26643 7656 26675
rect 7696 26643 7728 26675
rect 7768 26643 7800 26675
rect 7840 26643 7872 26675
rect 7912 26643 7944 26675
rect 7984 26643 8016 26675
rect 8056 26643 8088 26675
rect 8128 26643 8160 26675
rect 8200 26643 8232 26675
rect 8272 26643 8304 26675
rect 8344 26643 8376 26675
rect 8416 26643 8448 26675
rect 8488 26643 8520 26675
rect 8560 26643 8592 26675
rect 8632 26643 8664 26675
rect 8704 26643 8736 26675
rect 8776 26643 8808 26675
rect 8848 26643 8880 26675
rect 8920 26643 8952 26675
rect 8992 26643 9024 26675
rect 9064 26643 9096 26675
rect 9136 26643 9168 26675
rect 9208 26643 9240 26675
rect 9280 26643 9312 26675
rect 9352 26643 9384 26675
rect 9424 26643 9456 26675
rect 9496 26643 9528 26675
rect 9568 26643 9600 26675
rect 9640 26643 9672 26675
rect 9712 26643 9744 26675
rect 9784 26643 9816 26675
rect 9856 26643 9888 26675
rect 9928 26643 9960 26675
rect 10000 26643 10032 26675
rect 10072 26643 10104 26675
rect 10144 26643 10176 26675
rect 10216 26643 10248 26675
rect 10288 26643 10320 26675
rect 10360 26643 10392 26675
rect 10432 26643 10464 26675
rect 10504 26643 10536 26675
rect 10576 26643 10608 26675
rect 10648 26643 10680 26675
rect 10720 26643 10752 26675
rect 10792 26643 10824 26675
rect 10864 26643 10896 26675
rect 10936 26643 10968 26675
rect 11008 26643 11040 26675
rect 11080 26643 11112 26675
rect 11152 26643 11184 26675
rect 11224 26643 11256 26675
rect 11296 26643 11328 26675
rect 11368 26643 11400 26675
rect 11440 26643 11472 26675
rect 11512 26643 11544 26675
rect 11584 26643 11616 26675
rect 11656 26643 11688 26675
rect 11728 26643 11760 26675
rect 11800 26643 11832 26675
rect 11872 26643 11904 26675
rect 11944 26643 11976 26675
rect 12016 26643 12048 26675
rect 12088 26643 12120 26675
rect 12160 26643 12192 26675
rect 12232 26643 12264 26675
rect 12304 26643 12336 26675
rect 12376 26643 12408 26675
rect 12448 26643 12480 26675
rect 12520 26643 12552 26675
rect 12592 26643 12624 26675
rect 12664 26643 12696 26675
rect 12736 26643 12768 26675
rect 12808 26643 12840 26675
rect 12880 26643 12912 26675
rect 12952 26643 12984 26675
rect 13024 26643 13056 26675
rect 13096 26643 13128 26675
rect 13168 26643 13200 26675
rect 13240 26643 13272 26675
rect 13312 26643 13344 26675
rect 13384 26643 13416 26675
rect 13456 26643 13488 26675
rect 13528 26643 13560 26675
rect 13600 26643 13632 26675
rect 13672 26643 13704 26675
rect 13744 26643 13776 26675
rect 13816 26643 13848 26675
rect 13888 26643 13920 26675
rect 13960 26643 13992 26675
rect 14032 26643 14064 26675
rect 14104 26643 14136 26675
rect 14176 26643 14208 26675
rect 14248 26643 14280 26675
rect 14320 26643 14352 26675
rect 14392 26643 14424 26675
rect 14464 26643 14496 26675
rect 14536 26643 14568 26675
rect 14608 26643 14640 26675
rect 14680 26643 14712 26675
rect 14752 26643 14784 26675
rect 14824 26643 14856 26675
rect 14896 26643 14928 26675
rect 14968 26643 15000 26675
rect 15040 26643 15072 26675
rect 15112 26643 15144 26675
rect 15184 26643 15216 26675
rect 15256 26643 15288 26675
rect 15328 26643 15360 26675
rect 15400 26643 15432 26675
rect 15472 26643 15504 26675
rect 15544 26643 15576 26675
rect 15616 26643 15648 26675
rect 15688 26643 15720 26675
rect 15760 26643 15792 26675
rect 15832 26643 15864 26675
rect 15904 26643 15936 26675
rect 64 26571 96 26603
rect 136 26571 168 26603
rect 208 26571 240 26603
rect 280 26571 312 26603
rect 352 26571 384 26603
rect 424 26571 456 26603
rect 496 26571 528 26603
rect 568 26571 600 26603
rect 640 26571 672 26603
rect 712 26571 744 26603
rect 784 26571 816 26603
rect 856 26571 888 26603
rect 928 26571 960 26603
rect 1000 26571 1032 26603
rect 1072 26571 1104 26603
rect 1144 26571 1176 26603
rect 1216 26571 1248 26603
rect 1288 26571 1320 26603
rect 1360 26571 1392 26603
rect 1432 26571 1464 26603
rect 1504 26571 1536 26603
rect 1576 26571 1608 26603
rect 1648 26571 1680 26603
rect 1720 26571 1752 26603
rect 1792 26571 1824 26603
rect 1864 26571 1896 26603
rect 1936 26571 1968 26603
rect 2008 26571 2040 26603
rect 2080 26571 2112 26603
rect 2152 26571 2184 26603
rect 2224 26571 2256 26603
rect 2296 26571 2328 26603
rect 2368 26571 2400 26603
rect 2440 26571 2472 26603
rect 2512 26571 2544 26603
rect 2584 26571 2616 26603
rect 2656 26571 2688 26603
rect 2728 26571 2760 26603
rect 2800 26571 2832 26603
rect 2872 26571 2904 26603
rect 2944 26571 2976 26603
rect 3016 26571 3048 26603
rect 3088 26571 3120 26603
rect 3160 26571 3192 26603
rect 3232 26571 3264 26603
rect 3304 26571 3336 26603
rect 3376 26571 3408 26603
rect 3448 26571 3480 26603
rect 3520 26571 3552 26603
rect 3592 26571 3624 26603
rect 3664 26571 3696 26603
rect 3736 26571 3768 26603
rect 3808 26571 3840 26603
rect 3880 26571 3912 26603
rect 3952 26571 3984 26603
rect 4024 26571 4056 26603
rect 4096 26571 4128 26603
rect 4168 26571 4200 26603
rect 4240 26571 4272 26603
rect 4312 26571 4344 26603
rect 4384 26571 4416 26603
rect 4456 26571 4488 26603
rect 4528 26571 4560 26603
rect 4600 26571 4632 26603
rect 4672 26571 4704 26603
rect 4744 26571 4776 26603
rect 4816 26571 4848 26603
rect 4888 26571 4920 26603
rect 4960 26571 4992 26603
rect 5032 26571 5064 26603
rect 5104 26571 5136 26603
rect 5176 26571 5208 26603
rect 5248 26571 5280 26603
rect 5320 26571 5352 26603
rect 5392 26571 5424 26603
rect 5464 26571 5496 26603
rect 5536 26571 5568 26603
rect 5608 26571 5640 26603
rect 5680 26571 5712 26603
rect 5752 26571 5784 26603
rect 5824 26571 5856 26603
rect 5896 26571 5928 26603
rect 5968 26571 6000 26603
rect 6040 26571 6072 26603
rect 6112 26571 6144 26603
rect 6184 26571 6216 26603
rect 6256 26571 6288 26603
rect 6328 26571 6360 26603
rect 6400 26571 6432 26603
rect 6472 26571 6504 26603
rect 6544 26571 6576 26603
rect 6616 26571 6648 26603
rect 6688 26571 6720 26603
rect 6760 26571 6792 26603
rect 6832 26571 6864 26603
rect 6904 26571 6936 26603
rect 6976 26571 7008 26603
rect 7048 26571 7080 26603
rect 7120 26571 7152 26603
rect 7192 26571 7224 26603
rect 7264 26571 7296 26603
rect 7336 26571 7368 26603
rect 7408 26571 7440 26603
rect 7480 26571 7512 26603
rect 7552 26571 7584 26603
rect 7624 26571 7656 26603
rect 7696 26571 7728 26603
rect 7768 26571 7800 26603
rect 7840 26571 7872 26603
rect 7912 26571 7944 26603
rect 7984 26571 8016 26603
rect 8056 26571 8088 26603
rect 8128 26571 8160 26603
rect 8200 26571 8232 26603
rect 8272 26571 8304 26603
rect 8344 26571 8376 26603
rect 8416 26571 8448 26603
rect 8488 26571 8520 26603
rect 8560 26571 8592 26603
rect 8632 26571 8664 26603
rect 8704 26571 8736 26603
rect 8776 26571 8808 26603
rect 8848 26571 8880 26603
rect 8920 26571 8952 26603
rect 8992 26571 9024 26603
rect 9064 26571 9096 26603
rect 9136 26571 9168 26603
rect 9208 26571 9240 26603
rect 9280 26571 9312 26603
rect 9352 26571 9384 26603
rect 9424 26571 9456 26603
rect 9496 26571 9528 26603
rect 9568 26571 9600 26603
rect 9640 26571 9672 26603
rect 9712 26571 9744 26603
rect 9784 26571 9816 26603
rect 9856 26571 9888 26603
rect 9928 26571 9960 26603
rect 10000 26571 10032 26603
rect 10072 26571 10104 26603
rect 10144 26571 10176 26603
rect 10216 26571 10248 26603
rect 10288 26571 10320 26603
rect 10360 26571 10392 26603
rect 10432 26571 10464 26603
rect 10504 26571 10536 26603
rect 10576 26571 10608 26603
rect 10648 26571 10680 26603
rect 10720 26571 10752 26603
rect 10792 26571 10824 26603
rect 10864 26571 10896 26603
rect 10936 26571 10968 26603
rect 11008 26571 11040 26603
rect 11080 26571 11112 26603
rect 11152 26571 11184 26603
rect 11224 26571 11256 26603
rect 11296 26571 11328 26603
rect 11368 26571 11400 26603
rect 11440 26571 11472 26603
rect 11512 26571 11544 26603
rect 11584 26571 11616 26603
rect 11656 26571 11688 26603
rect 11728 26571 11760 26603
rect 11800 26571 11832 26603
rect 11872 26571 11904 26603
rect 11944 26571 11976 26603
rect 12016 26571 12048 26603
rect 12088 26571 12120 26603
rect 12160 26571 12192 26603
rect 12232 26571 12264 26603
rect 12304 26571 12336 26603
rect 12376 26571 12408 26603
rect 12448 26571 12480 26603
rect 12520 26571 12552 26603
rect 12592 26571 12624 26603
rect 12664 26571 12696 26603
rect 12736 26571 12768 26603
rect 12808 26571 12840 26603
rect 12880 26571 12912 26603
rect 12952 26571 12984 26603
rect 13024 26571 13056 26603
rect 13096 26571 13128 26603
rect 13168 26571 13200 26603
rect 13240 26571 13272 26603
rect 13312 26571 13344 26603
rect 13384 26571 13416 26603
rect 13456 26571 13488 26603
rect 13528 26571 13560 26603
rect 13600 26571 13632 26603
rect 13672 26571 13704 26603
rect 13744 26571 13776 26603
rect 13816 26571 13848 26603
rect 13888 26571 13920 26603
rect 13960 26571 13992 26603
rect 14032 26571 14064 26603
rect 14104 26571 14136 26603
rect 14176 26571 14208 26603
rect 14248 26571 14280 26603
rect 14320 26571 14352 26603
rect 14392 26571 14424 26603
rect 14464 26571 14496 26603
rect 14536 26571 14568 26603
rect 14608 26571 14640 26603
rect 14680 26571 14712 26603
rect 14752 26571 14784 26603
rect 14824 26571 14856 26603
rect 14896 26571 14928 26603
rect 14968 26571 15000 26603
rect 15040 26571 15072 26603
rect 15112 26571 15144 26603
rect 15184 26571 15216 26603
rect 15256 26571 15288 26603
rect 15328 26571 15360 26603
rect 15400 26571 15432 26603
rect 15472 26571 15504 26603
rect 15544 26571 15576 26603
rect 15616 26571 15648 26603
rect 15688 26571 15720 26603
rect 15760 26571 15792 26603
rect 15832 26571 15864 26603
rect 15904 26571 15936 26603
rect 64 26499 96 26531
rect 136 26499 168 26531
rect 208 26499 240 26531
rect 280 26499 312 26531
rect 352 26499 384 26531
rect 424 26499 456 26531
rect 496 26499 528 26531
rect 568 26499 600 26531
rect 640 26499 672 26531
rect 712 26499 744 26531
rect 784 26499 816 26531
rect 856 26499 888 26531
rect 928 26499 960 26531
rect 1000 26499 1032 26531
rect 1072 26499 1104 26531
rect 1144 26499 1176 26531
rect 1216 26499 1248 26531
rect 1288 26499 1320 26531
rect 1360 26499 1392 26531
rect 1432 26499 1464 26531
rect 1504 26499 1536 26531
rect 1576 26499 1608 26531
rect 1648 26499 1680 26531
rect 1720 26499 1752 26531
rect 1792 26499 1824 26531
rect 1864 26499 1896 26531
rect 1936 26499 1968 26531
rect 2008 26499 2040 26531
rect 2080 26499 2112 26531
rect 2152 26499 2184 26531
rect 2224 26499 2256 26531
rect 2296 26499 2328 26531
rect 2368 26499 2400 26531
rect 2440 26499 2472 26531
rect 2512 26499 2544 26531
rect 2584 26499 2616 26531
rect 2656 26499 2688 26531
rect 2728 26499 2760 26531
rect 2800 26499 2832 26531
rect 2872 26499 2904 26531
rect 2944 26499 2976 26531
rect 3016 26499 3048 26531
rect 3088 26499 3120 26531
rect 3160 26499 3192 26531
rect 3232 26499 3264 26531
rect 3304 26499 3336 26531
rect 3376 26499 3408 26531
rect 3448 26499 3480 26531
rect 3520 26499 3552 26531
rect 3592 26499 3624 26531
rect 3664 26499 3696 26531
rect 3736 26499 3768 26531
rect 3808 26499 3840 26531
rect 3880 26499 3912 26531
rect 3952 26499 3984 26531
rect 4024 26499 4056 26531
rect 4096 26499 4128 26531
rect 4168 26499 4200 26531
rect 4240 26499 4272 26531
rect 4312 26499 4344 26531
rect 4384 26499 4416 26531
rect 4456 26499 4488 26531
rect 4528 26499 4560 26531
rect 4600 26499 4632 26531
rect 4672 26499 4704 26531
rect 4744 26499 4776 26531
rect 4816 26499 4848 26531
rect 4888 26499 4920 26531
rect 4960 26499 4992 26531
rect 5032 26499 5064 26531
rect 5104 26499 5136 26531
rect 5176 26499 5208 26531
rect 5248 26499 5280 26531
rect 5320 26499 5352 26531
rect 5392 26499 5424 26531
rect 5464 26499 5496 26531
rect 5536 26499 5568 26531
rect 5608 26499 5640 26531
rect 5680 26499 5712 26531
rect 5752 26499 5784 26531
rect 5824 26499 5856 26531
rect 5896 26499 5928 26531
rect 5968 26499 6000 26531
rect 6040 26499 6072 26531
rect 6112 26499 6144 26531
rect 6184 26499 6216 26531
rect 6256 26499 6288 26531
rect 6328 26499 6360 26531
rect 6400 26499 6432 26531
rect 6472 26499 6504 26531
rect 6544 26499 6576 26531
rect 6616 26499 6648 26531
rect 6688 26499 6720 26531
rect 6760 26499 6792 26531
rect 6832 26499 6864 26531
rect 6904 26499 6936 26531
rect 6976 26499 7008 26531
rect 7048 26499 7080 26531
rect 7120 26499 7152 26531
rect 7192 26499 7224 26531
rect 7264 26499 7296 26531
rect 7336 26499 7368 26531
rect 7408 26499 7440 26531
rect 7480 26499 7512 26531
rect 7552 26499 7584 26531
rect 7624 26499 7656 26531
rect 7696 26499 7728 26531
rect 7768 26499 7800 26531
rect 7840 26499 7872 26531
rect 7912 26499 7944 26531
rect 7984 26499 8016 26531
rect 8056 26499 8088 26531
rect 8128 26499 8160 26531
rect 8200 26499 8232 26531
rect 8272 26499 8304 26531
rect 8344 26499 8376 26531
rect 8416 26499 8448 26531
rect 8488 26499 8520 26531
rect 8560 26499 8592 26531
rect 8632 26499 8664 26531
rect 8704 26499 8736 26531
rect 8776 26499 8808 26531
rect 8848 26499 8880 26531
rect 8920 26499 8952 26531
rect 8992 26499 9024 26531
rect 9064 26499 9096 26531
rect 9136 26499 9168 26531
rect 9208 26499 9240 26531
rect 9280 26499 9312 26531
rect 9352 26499 9384 26531
rect 9424 26499 9456 26531
rect 9496 26499 9528 26531
rect 9568 26499 9600 26531
rect 9640 26499 9672 26531
rect 9712 26499 9744 26531
rect 9784 26499 9816 26531
rect 9856 26499 9888 26531
rect 9928 26499 9960 26531
rect 10000 26499 10032 26531
rect 10072 26499 10104 26531
rect 10144 26499 10176 26531
rect 10216 26499 10248 26531
rect 10288 26499 10320 26531
rect 10360 26499 10392 26531
rect 10432 26499 10464 26531
rect 10504 26499 10536 26531
rect 10576 26499 10608 26531
rect 10648 26499 10680 26531
rect 10720 26499 10752 26531
rect 10792 26499 10824 26531
rect 10864 26499 10896 26531
rect 10936 26499 10968 26531
rect 11008 26499 11040 26531
rect 11080 26499 11112 26531
rect 11152 26499 11184 26531
rect 11224 26499 11256 26531
rect 11296 26499 11328 26531
rect 11368 26499 11400 26531
rect 11440 26499 11472 26531
rect 11512 26499 11544 26531
rect 11584 26499 11616 26531
rect 11656 26499 11688 26531
rect 11728 26499 11760 26531
rect 11800 26499 11832 26531
rect 11872 26499 11904 26531
rect 11944 26499 11976 26531
rect 12016 26499 12048 26531
rect 12088 26499 12120 26531
rect 12160 26499 12192 26531
rect 12232 26499 12264 26531
rect 12304 26499 12336 26531
rect 12376 26499 12408 26531
rect 12448 26499 12480 26531
rect 12520 26499 12552 26531
rect 12592 26499 12624 26531
rect 12664 26499 12696 26531
rect 12736 26499 12768 26531
rect 12808 26499 12840 26531
rect 12880 26499 12912 26531
rect 12952 26499 12984 26531
rect 13024 26499 13056 26531
rect 13096 26499 13128 26531
rect 13168 26499 13200 26531
rect 13240 26499 13272 26531
rect 13312 26499 13344 26531
rect 13384 26499 13416 26531
rect 13456 26499 13488 26531
rect 13528 26499 13560 26531
rect 13600 26499 13632 26531
rect 13672 26499 13704 26531
rect 13744 26499 13776 26531
rect 13816 26499 13848 26531
rect 13888 26499 13920 26531
rect 13960 26499 13992 26531
rect 14032 26499 14064 26531
rect 14104 26499 14136 26531
rect 14176 26499 14208 26531
rect 14248 26499 14280 26531
rect 14320 26499 14352 26531
rect 14392 26499 14424 26531
rect 14464 26499 14496 26531
rect 14536 26499 14568 26531
rect 14608 26499 14640 26531
rect 14680 26499 14712 26531
rect 14752 26499 14784 26531
rect 14824 26499 14856 26531
rect 14896 26499 14928 26531
rect 14968 26499 15000 26531
rect 15040 26499 15072 26531
rect 15112 26499 15144 26531
rect 15184 26499 15216 26531
rect 15256 26499 15288 26531
rect 15328 26499 15360 26531
rect 15400 26499 15432 26531
rect 15472 26499 15504 26531
rect 15544 26499 15576 26531
rect 15616 26499 15648 26531
rect 15688 26499 15720 26531
rect 15760 26499 15792 26531
rect 15832 26499 15864 26531
rect 15904 26499 15936 26531
rect 64 26427 96 26459
rect 136 26427 168 26459
rect 208 26427 240 26459
rect 280 26427 312 26459
rect 352 26427 384 26459
rect 424 26427 456 26459
rect 496 26427 528 26459
rect 568 26427 600 26459
rect 640 26427 672 26459
rect 712 26427 744 26459
rect 784 26427 816 26459
rect 856 26427 888 26459
rect 928 26427 960 26459
rect 1000 26427 1032 26459
rect 1072 26427 1104 26459
rect 1144 26427 1176 26459
rect 1216 26427 1248 26459
rect 1288 26427 1320 26459
rect 1360 26427 1392 26459
rect 1432 26427 1464 26459
rect 1504 26427 1536 26459
rect 1576 26427 1608 26459
rect 1648 26427 1680 26459
rect 1720 26427 1752 26459
rect 1792 26427 1824 26459
rect 1864 26427 1896 26459
rect 1936 26427 1968 26459
rect 2008 26427 2040 26459
rect 2080 26427 2112 26459
rect 2152 26427 2184 26459
rect 2224 26427 2256 26459
rect 2296 26427 2328 26459
rect 2368 26427 2400 26459
rect 2440 26427 2472 26459
rect 2512 26427 2544 26459
rect 2584 26427 2616 26459
rect 2656 26427 2688 26459
rect 2728 26427 2760 26459
rect 2800 26427 2832 26459
rect 2872 26427 2904 26459
rect 2944 26427 2976 26459
rect 3016 26427 3048 26459
rect 3088 26427 3120 26459
rect 3160 26427 3192 26459
rect 3232 26427 3264 26459
rect 3304 26427 3336 26459
rect 3376 26427 3408 26459
rect 3448 26427 3480 26459
rect 3520 26427 3552 26459
rect 3592 26427 3624 26459
rect 3664 26427 3696 26459
rect 3736 26427 3768 26459
rect 3808 26427 3840 26459
rect 3880 26427 3912 26459
rect 3952 26427 3984 26459
rect 4024 26427 4056 26459
rect 4096 26427 4128 26459
rect 4168 26427 4200 26459
rect 4240 26427 4272 26459
rect 4312 26427 4344 26459
rect 4384 26427 4416 26459
rect 4456 26427 4488 26459
rect 4528 26427 4560 26459
rect 4600 26427 4632 26459
rect 4672 26427 4704 26459
rect 4744 26427 4776 26459
rect 4816 26427 4848 26459
rect 4888 26427 4920 26459
rect 4960 26427 4992 26459
rect 5032 26427 5064 26459
rect 5104 26427 5136 26459
rect 5176 26427 5208 26459
rect 5248 26427 5280 26459
rect 5320 26427 5352 26459
rect 5392 26427 5424 26459
rect 5464 26427 5496 26459
rect 5536 26427 5568 26459
rect 5608 26427 5640 26459
rect 5680 26427 5712 26459
rect 5752 26427 5784 26459
rect 5824 26427 5856 26459
rect 5896 26427 5928 26459
rect 5968 26427 6000 26459
rect 6040 26427 6072 26459
rect 6112 26427 6144 26459
rect 6184 26427 6216 26459
rect 6256 26427 6288 26459
rect 6328 26427 6360 26459
rect 6400 26427 6432 26459
rect 6472 26427 6504 26459
rect 6544 26427 6576 26459
rect 6616 26427 6648 26459
rect 6688 26427 6720 26459
rect 6760 26427 6792 26459
rect 6832 26427 6864 26459
rect 6904 26427 6936 26459
rect 6976 26427 7008 26459
rect 7048 26427 7080 26459
rect 7120 26427 7152 26459
rect 7192 26427 7224 26459
rect 7264 26427 7296 26459
rect 7336 26427 7368 26459
rect 7408 26427 7440 26459
rect 7480 26427 7512 26459
rect 7552 26427 7584 26459
rect 7624 26427 7656 26459
rect 7696 26427 7728 26459
rect 7768 26427 7800 26459
rect 7840 26427 7872 26459
rect 7912 26427 7944 26459
rect 7984 26427 8016 26459
rect 8056 26427 8088 26459
rect 8128 26427 8160 26459
rect 8200 26427 8232 26459
rect 8272 26427 8304 26459
rect 8344 26427 8376 26459
rect 8416 26427 8448 26459
rect 8488 26427 8520 26459
rect 8560 26427 8592 26459
rect 8632 26427 8664 26459
rect 8704 26427 8736 26459
rect 8776 26427 8808 26459
rect 8848 26427 8880 26459
rect 8920 26427 8952 26459
rect 8992 26427 9024 26459
rect 9064 26427 9096 26459
rect 9136 26427 9168 26459
rect 9208 26427 9240 26459
rect 9280 26427 9312 26459
rect 9352 26427 9384 26459
rect 9424 26427 9456 26459
rect 9496 26427 9528 26459
rect 9568 26427 9600 26459
rect 9640 26427 9672 26459
rect 9712 26427 9744 26459
rect 9784 26427 9816 26459
rect 9856 26427 9888 26459
rect 9928 26427 9960 26459
rect 10000 26427 10032 26459
rect 10072 26427 10104 26459
rect 10144 26427 10176 26459
rect 10216 26427 10248 26459
rect 10288 26427 10320 26459
rect 10360 26427 10392 26459
rect 10432 26427 10464 26459
rect 10504 26427 10536 26459
rect 10576 26427 10608 26459
rect 10648 26427 10680 26459
rect 10720 26427 10752 26459
rect 10792 26427 10824 26459
rect 10864 26427 10896 26459
rect 10936 26427 10968 26459
rect 11008 26427 11040 26459
rect 11080 26427 11112 26459
rect 11152 26427 11184 26459
rect 11224 26427 11256 26459
rect 11296 26427 11328 26459
rect 11368 26427 11400 26459
rect 11440 26427 11472 26459
rect 11512 26427 11544 26459
rect 11584 26427 11616 26459
rect 11656 26427 11688 26459
rect 11728 26427 11760 26459
rect 11800 26427 11832 26459
rect 11872 26427 11904 26459
rect 11944 26427 11976 26459
rect 12016 26427 12048 26459
rect 12088 26427 12120 26459
rect 12160 26427 12192 26459
rect 12232 26427 12264 26459
rect 12304 26427 12336 26459
rect 12376 26427 12408 26459
rect 12448 26427 12480 26459
rect 12520 26427 12552 26459
rect 12592 26427 12624 26459
rect 12664 26427 12696 26459
rect 12736 26427 12768 26459
rect 12808 26427 12840 26459
rect 12880 26427 12912 26459
rect 12952 26427 12984 26459
rect 13024 26427 13056 26459
rect 13096 26427 13128 26459
rect 13168 26427 13200 26459
rect 13240 26427 13272 26459
rect 13312 26427 13344 26459
rect 13384 26427 13416 26459
rect 13456 26427 13488 26459
rect 13528 26427 13560 26459
rect 13600 26427 13632 26459
rect 13672 26427 13704 26459
rect 13744 26427 13776 26459
rect 13816 26427 13848 26459
rect 13888 26427 13920 26459
rect 13960 26427 13992 26459
rect 14032 26427 14064 26459
rect 14104 26427 14136 26459
rect 14176 26427 14208 26459
rect 14248 26427 14280 26459
rect 14320 26427 14352 26459
rect 14392 26427 14424 26459
rect 14464 26427 14496 26459
rect 14536 26427 14568 26459
rect 14608 26427 14640 26459
rect 14680 26427 14712 26459
rect 14752 26427 14784 26459
rect 14824 26427 14856 26459
rect 14896 26427 14928 26459
rect 14968 26427 15000 26459
rect 15040 26427 15072 26459
rect 15112 26427 15144 26459
rect 15184 26427 15216 26459
rect 15256 26427 15288 26459
rect 15328 26427 15360 26459
rect 15400 26427 15432 26459
rect 15472 26427 15504 26459
rect 15544 26427 15576 26459
rect 15616 26427 15648 26459
rect 15688 26427 15720 26459
rect 15760 26427 15792 26459
rect 15832 26427 15864 26459
rect 15904 26427 15936 26459
rect 64 26355 96 26387
rect 136 26355 168 26387
rect 208 26355 240 26387
rect 280 26355 312 26387
rect 352 26355 384 26387
rect 424 26355 456 26387
rect 496 26355 528 26387
rect 568 26355 600 26387
rect 640 26355 672 26387
rect 712 26355 744 26387
rect 784 26355 816 26387
rect 856 26355 888 26387
rect 928 26355 960 26387
rect 1000 26355 1032 26387
rect 1072 26355 1104 26387
rect 1144 26355 1176 26387
rect 1216 26355 1248 26387
rect 1288 26355 1320 26387
rect 1360 26355 1392 26387
rect 1432 26355 1464 26387
rect 1504 26355 1536 26387
rect 1576 26355 1608 26387
rect 1648 26355 1680 26387
rect 1720 26355 1752 26387
rect 1792 26355 1824 26387
rect 1864 26355 1896 26387
rect 1936 26355 1968 26387
rect 2008 26355 2040 26387
rect 2080 26355 2112 26387
rect 2152 26355 2184 26387
rect 2224 26355 2256 26387
rect 2296 26355 2328 26387
rect 2368 26355 2400 26387
rect 2440 26355 2472 26387
rect 2512 26355 2544 26387
rect 2584 26355 2616 26387
rect 2656 26355 2688 26387
rect 2728 26355 2760 26387
rect 2800 26355 2832 26387
rect 2872 26355 2904 26387
rect 2944 26355 2976 26387
rect 3016 26355 3048 26387
rect 3088 26355 3120 26387
rect 3160 26355 3192 26387
rect 3232 26355 3264 26387
rect 3304 26355 3336 26387
rect 3376 26355 3408 26387
rect 3448 26355 3480 26387
rect 3520 26355 3552 26387
rect 3592 26355 3624 26387
rect 3664 26355 3696 26387
rect 3736 26355 3768 26387
rect 3808 26355 3840 26387
rect 3880 26355 3912 26387
rect 3952 26355 3984 26387
rect 4024 26355 4056 26387
rect 4096 26355 4128 26387
rect 4168 26355 4200 26387
rect 4240 26355 4272 26387
rect 4312 26355 4344 26387
rect 4384 26355 4416 26387
rect 4456 26355 4488 26387
rect 4528 26355 4560 26387
rect 4600 26355 4632 26387
rect 4672 26355 4704 26387
rect 4744 26355 4776 26387
rect 4816 26355 4848 26387
rect 4888 26355 4920 26387
rect 4960 26355 4992 26387
rect 5032 26355 5064 26387
rect 5104 26355 5136 26387
rect 5176 26355 5208 26387
rect 5248 26355 5280 26387
rect 5320 26355 5352 26387
rect 5392 26355 5424 26387
rect 5464 26355 5496 26387
rect 5536 26355 5568 26387
rect 5608 26355 5640 26387
rect 5680 26355 5712 26387
rect 5752 26355 5784 26387
rect 5824 26355 5856 26387
rect 5896 26355 5928 26387
rect 5968 26355 6000 26387
rect 6040 26355 6072 26387
rect 6112 26355 6144 26387
rect 6184 26355 6216 26387
rect 6256 26355 6288 26387
rect 6328 26355 6360 26387
rect 6400 26355 6432 26387
rect 6472 26355 6504 26387
rect 6544 26355 6576 26387
rect 6616 26355 6648 26387
rect 6688 26355 6720 26387
rect 6760 26355 6792 26387
rect 6832 26355 6864 26387
rect 6904 26355 6936 26387
rect 6976 26355 7008 26387
rect 7048 26355 7080 26387
rect 7120 26355 7152 26387
rect 7192 26355 7224 26387
rect 7264 26355 7296 26387
rect 7336 26355 7368 26387
rect 7408 26355 7440 26387
rect 7480 26355 7512 26387
rect 7552 26355 7584 26387
rect 7624 26355 7656 26387
rect 7696 26355 7728 26387
rect 7768 26355 7800 26387
rect 7840 26355 7872 26387
rect 7912 26355 7944 26387
rect 7984 26355 8016 26387
rect 8056 26355 8088 26387
rect 8128 26355 8160 26387
rect 8200 26355 8232 26387
rect 8272 26355 8304 26387
rect 8344 26355 8376 26387
rect 8416 26355 8448 26387
rect 8488 26355 8520 26387
rect 8560 26355 8592 26387
rect 8632 26355 8664 26387
rect 8704 26355 8736 26387
rect 8776 26355 8808 26387
rect 8848 26355 8880 26387
rect 8920 26355 8952 26387
rect 8992 26355 9024 26387
rect 9064 26355 9096 26387
rect 9136 26355 9168 26387
rect 9208 26355 9240 26387
rect 9280 26355 9312 26387
rect 9352 26355 9384 26387
rect 9424 26355 9456 26387
rect 9496 26355 9528 26387
rect 9568 26355 9600 26387
rect 9640 26355 9672 26387
rect 9712 26355 9744 26387
rect 9784 26355 9816 26387
rect 9856 26355 9888 26387
rect 9928 26355 9960 26387
rect 10000 26355 10032 26387
rect 10072 26355 10104 26387
rect 10144 26355 10176 26387
rect 10216 26355 10248 26387
rect 10288 26355 10320 26387
rect 10360 26355 10392 26387
rect 10432 26355 10464 26387
rect 10504 26355 10536 26387
rect 10576 26355 10608 26387
rect 10648 26355 10680 26387
rect 10720 26355 10752 26387
rect 10792 26355 10824 26387
rect 10864 26355 10896 26387
rect 10936 26355 10968 26387
rect 11008 26355 11040 26387
rect 11080 26355 11112 26387
rect 11152 26355 11184 26387
rect 11224 26355 11256 26387
rect 11296 26355 11328 26387
rect 11368 26355 11400 26387
rect 11440 26355 11472 26387
rect 11512 26355 11544 26387
rect 11584 26355 11616 26387
rect 11656 26355 11688 26387
rect 11728 26355 11760 26387
rect 11800 26355 11832 26387
rect 11872 26355 11904 26387
rect 11944 26355 11976 26387
rect 12016 26355 12048 26387
rect 12088 26355 12120 26387
rect 12160 26355 12192 26387
rect 12232 26355 12264 26387
rect 12304 26355 12336 26387
rect 12376 26355 12408 26387
rect 12448 26355 12480 26387
rect 12520 26355 12552 26387
rect 12592 26355 12624 26387
rect 12664 26355 12696 26387
rect 12736 26355 12768 26387
rect 12808 26355 12840 26387
rect 12880 26355 12912 26387
rect 12952 26355 12984 26387
rect 13024 26355 13056 26387
rect 13096 26355 13128 26387
rect 13168 26355 13200 26387
rect 13240 26355 13272 26387
rect 13312 26355 13344 26387
rect 13384 26355 13416 26387
rect 13456 26355 13488 26387
rect 13528 26355 13560 26387
rect 13600 26355 13632 26387
rect 13672 26355 13704 26387
rect 13744 26355 13776 26387
rect 13816 26355 13848 26387
rect 13888 26355 13920 26387
rect 13960 26355 13992 26387
rect 14032 26355 14064 26387
rect 14104 26355 14136 26387
rect 14176 26355 14208 26387
rect 14248 26355 14280 26387
rect 14320 26355 14352 26387
rect 14392 26355 14424 26387
rect 14464 26355 14496 26387
rect 14536 26355 14568 26387
rect 14608 26355 14640 26387
rect 14680 26355 14712 26387
rect 14752 26355 14784 26387
rect 14824 26355 14856 26387
rect 14896 26355 14928 26387
rect 14968 26355 15000 26387
rect 15040 26355 15072 26387
rect 15112 26355 15144 26387
rect 15184 26355 15216 26387
rect 15256 26355 15288 26387
rect 15328 26355 15360 26387
rect 15400 26355 15432 26387
rect 15472 26355 15504 26387
rect 15544 26355 15576 26387
rect 15616 26355 15648 26387
rect 15688 26355 15720 26387
rect 15760 26355 15792 26387
rect 15832 26355 15864 26387
rect 15904 26355 15936 26387
rect 64 26283 96 26315
rect 136 26283 168 26315
rect 208 26283 240 26315
rect 280 26283 312 26315
rect 352 26283 384 26315
rect 424 26283 456 26315
rect 496 26283 528 26315
rect 568 26283 600 26315
rect 640 26283 672 26315
rect 712 26283 744 26315
rect 784 26283 816 26315
rect 856 26283 888 26315
rect 928 26283 960 26315
rect 1000 26283 1032 26315
rect 1072 26283 1104 26315
rect 1144 26283 1176 26315
rect 1216 26283 1248 26315
rect 1288 26283 1320 26315
rect 1360 26283 1392 26315
rect 1432 26283 1464 26315
rect 1504 26283 1536 26315
rect 1576 26283 1608 26315
rect 1648 26283 1680 26315
rect 1720 26283 1752 26315
rect 1792 26283 1824 26315
rect 1864 26283 1896 26315
rect 1936 26283 1968 26315
rect 2008 26283 2040 26315
rect 2080 26283 2112 26315
rect 2152 26283 2184 26315
rect 2224 26283 2256 26315
rect 2296 26283 2328 26315
rect 2368 26283 2400 26315
rect 2440 26283 2472 26315
rect 2512 26283 2544 26315
rect 2584 26283 2616 26315
rect 2656 26283 2688 26315
rect 2728 26283 2760 26315
rect 2800 26283 2832 26315
rect 2872 26283 2904 26315
rect 2944 26283 2976 26315
rect 3016 26283 3048 26315
rect 3088 26283 3120 26315
rect 3160 26283 3192 26315
rect 3232 26283 3264 26315
rect 3304 26283 3336 26315
rect 3376 26283 3408 26315
rect 3448 26283 3480 26315
rect 3520 26283 3552 26315
rect 3592 26283 3624 26315
rect 3664 26283 3696 26315
rect 3736 26283 3768 26315
rect 3808 26283 3840 26315
rect 3880 26283 3912 26315
rect 3952 26283 3984 26315
rect 4024 26283 4056 26315
rect 4096 26283 4128 26315
rect 4168 26283 4200 26315
rect 4240 26283 4272 26315
rect 4312 26283 4344 26315
rect 4384 26283 4416 26315
rect 4456 26283 4488 26315
rect 4528 26283 4560 26315
rect 4600 26283 4632 26315
rect 4672 26283 4704 26315
rect 4744 26283 4776 26315
rect 4816 26283 4848 26315
rect 4888 26283 4920 26315
rect 4960 26283 4992 26315
rect 5032 26283 5064 26315
rect 5104 26283 5136 26315
rect 5176 26283 5208 26315
rect 5248 26283 5280 26315
rect 5320 26283 5352 26315
rect 5392 26283 5424 26315
rect 5464 26283 5496 26315
rect 5536 26283 5568 26315
rect 5608 26283 5640 26315
rect 5680 26283 5712 26315
rect 5752 26283 5784 26315
rect 5824 26283 5856 26315
rect 5896 26283 5928 26315
rect 5968 26283 6000 26315
rect 6040 26283 6072 26315
rect 6112 26283 6144 26315
rect 6184 26283 6216 26315
rect 6256 26283 6288 26315
rect 6328 26283 6360 26315
rect 6400 26283 6432 26315
rect 6472 26283 6504 26315
rect 6544 26283 6576 26315
rect 6616 26283 6648 26315
rect 6688 26283 6720 26315
rect 6760 26283 6792 26315
rect 6832 26283 6864 26315
rect 6904 26283 6936 26315
rect 6976 26283 7008 26315
rect 7048 26283 7080 26315
rect 7120 26283 7152 26315
rect 7192 26283 7224 26315
rect 7264 26283 7296 26315
rect 7336 26283 7368 26315
rect 7408 26283 7440 26315
rect 7480 26283 7512 26315
rect 7552 26283 7584 26315
rect 7624 26283 7656 26315
rect 7696 26283 7728 26315
rect 7768 26283 7800 26315
rect 7840 26283 7872 26315
rect 7912 26283 7944 26315
rect 7984 26283 8016 26315
rect 8056 26283 8088 26315
rect 8128 26283 8160 26315
rect 8200 26283 8232 26315
rect 8272 26283 8304 26315
rect 8344 26283 8376 26315
rect 8416 26283 8448 26315
rect 8488 26283 8520 26315
rect 8560 26283 8592 26315
rect 8632 26283 8664 26315
rect 8704 26283 8736 26315
rect 8776 26283 8808 26315
rect 8848 26283 8880 26315
rect 8920 26283 8952 26315
rect 8992 26283 9024 26315
rect 9064 26283 9096 26315
rect 9136 26283 9168 26315
rect 9208 26283 9240 26315
rect 9280 26283 9312 26315
rect 9352 26283 9384 26315
rect 9424 26283 9456 26315
rect 9496 26283 9528 26315
rect 9568 26283 9600 26315
rect 9640 26283 9672 26315
rect 9712 26283 9744 26315
rect 9784 26283 9816 26315
rect 9856 26283 9888 26315
rect 9928 26283 9960 26315
rect 10000 26283 10032 26315
rect 10072 26283 10104 26315
rect 10144 26283 10176 26315
rect 10216 26283 10248 26315
rect 10288 26283 10320 26315
rect 10360 26283 10392 26315
rect 10432 26283 10464 26315
rect 10504 26283 10536 26315
rect 10576 26283 10608 26315
rect 10648 26283 10680 26315
rect 10720 26283 10752 26315
rect 10792 26283 10824 26315
rect 10864 26283 10896 26315
rect 10936 26283 10968 26315
rect 11008 26283 11040 26315
rect 11080 26283 11112 26315
rect 11152 26283 11184 26315
rect 11224 26283 11256 26315
rect 11296 26283 11328 26315
rect 11368 26283 11400 26315
rect 11440 26283 11472 26315
rect 11512 26283 11544 26315
rect 11584 26283 11616 26315
rect 11656 26283 11688 26315
rect 11728 26283 11760 26315
rect 11800 26283 11832 26315
rect 11872 26283 11904 26315
rect 11944 26283 11976 26315
rect 12016 26283 12048 26315
rect 12088 26283 12120 26315
rect 12160 26283 12192 26315
rect 12232 26283 12264 26315
rect 12304 26283 12336 26315
rect 12376 26283 12408 26315
rect 12448 26283 12480 26315
rect 12520 26283 12552 26315
rect 12592 26283 12624 26315
rect 12664 26283 12696 26315
rect 12736 26283 12768 26315
rect 12808 26283 12840 26315
rect 12880 26283 12912 26315
rect 12952 26283 12984 26315
rect 13024 26283 13056 26315
rect 13096 26283 13128 26315
rect 13168 26283 13200 26315
rect 13240 26283 13272 26315
rect 13312 26283 13344 26315
rect 13384 26283 13416 26315
rect 13456 26283 13488 26315
rect 13528 26283 13560 26315
rect 13600 26283 13632 26315
rect 13672 26283 13704 26315
rect 13744 26283 13776 26315
rect 13816 26283 13848 26315
rect 13888 26283 13920 26315
rect 13960 26283 13992 26315
rect 14032 26283 14064 26315
rect 14104 26283 14136 26315
rect 14176 26283 14208 26315
rect 14248 26283 14280 26315
rect 14320 26283 14352 26315
rect 14392 26283 14424 26315
rect 14464 26283 14496 26315
rect 14536 26283 14568 26315
rect 14608 26283 14640 26315
rect 14680 26283 14712 26315
rect 14752 26283 14784 26315
rect 14824 26283 14856 26315
rect 14896 26283 14928 26315
rect 14968 26283 15000 26315
rect 15040 26283 15072 26315
rect 15112 26283 15144 26315
rect 15184 26283 15216 26315
rect 15256 26283 15288 26315
rect 15328 26283 15360 26315
rect 15400 26283 15432 26315
rect 15472 26283 15504 26315
rect 15544 26283 15576 26315
rect 15616 26283 15648 26315
rect 15688 26283 15720 26315
rect 15760 26283 15792 26315
rect 15832 26283 15864 26315
rect 15904 26283 15936 26315
rect 64 26211 96 26243
rect 136 26211 168 26243
rect 208 26211 240 26243
rect 280 26211 312 26243
rect 352 26211 384 26243
rect 424 26211 456 26243
rect 496 26211 528 26243
rect 568 26211 600 26243
rect 640 26211 672 26243
rect 712 26211 744 26243
rect 784 26211 816 26243
rect 856 26211 888 26243
rect 928 26211 960 26243
rect 1000 26211 1032 26243
rect 1072 26211 1104 26243
rect 1144 26211 1176 26243
rect 1216 26211 1248 26243
rect 1288 26211 1320 26243
rect 1360 26211 1392 26243
rect 1432 26211 1464 26243
rect 1504 26211 1536 26243
rect 1576 26211 1608 26243
rect 1648 26211 1680 26243
rect 1720 26211 1752 26243
rect 1792 26211 1824 26243
rect 1864 26211 1896 26243
rect 1936 26211 1968 26243
rect 2008 26211 2040 26243
rect 2080 26211 2112 26243
rect 2152 26211 2184 26243
rect 2224 26211 2256 26243
rect 2296 26211 2328 26243
rect 2368 26211 2400 26243
rect 2440 26211 2472 26243
rect 2512 26211 2544 26243
rect 2584 26211 2616 26243
rect 2656 26211 2688 26243
rect 2728 26211 2760 26243
rect 2800 26211 2832 26243
rect 2872 26211 2904 26243
rect 2944 26211 2976 26243
rect 3016 26211 3048 26243
rect 3088 26211 3120 26243
rect 3160 26211 3192 26243
rect 3232 26211 3264 26243
rect 3304 26211 3336 26243
rect 3376 26211 3408 26243
rect 3448 26211 3480 26243
rect 3520 26211 3552 26243
rect 3592 26211 3624 26243
rect 3664 26211 3696 26243
rect 3736 26211 3768 26243
rect 3808 26211 3840 26243
rect 3880 26211 3912 26243
rect 3952 26211 3984 26243
rect 4024 26211 4056 26243
rect 4096 26211 4128 26243
rect 4168 26211 4200 26243
rect 4240 26211 4272 26243
rect 4312 26211 4344 26243
rect 4384 26211 4416 26243
rect 4456 26211 4488 26243
rect 4528 26211 4560 26243
rect 4600 26211 4632 26243
rect 4672 26211 4704 26243
rect 4744 26211 4776 26243
rect 4816 26211 4848 26243
rect 4888 26211 4920 26243
rect 4960 26211 4992 26243
rect 5032 26211 5064 26243
rect 5104 26211 5136 26243
rect 5176 26211 5208 26243
rect 5248 26211 5280 26243
rect 5320 26211 5352 26243
rect 5392 26211 5424 26243
rect 5464 26211 5496 26243
rect 5536 26211 5568 26243
rect 5608 26211 5640 26243
rect 5680 26211 5712 26243
rect 5752 26211 5784 26243
rect 5824 26211 5856 26243
rect 5896 26211 5928 26243
rect 5968 26211 6000 26243
rect 6040 26211 6072 26243
rect 6112 26211 6144 26243
rect 6184 26211 6216 26243
rect 6256 26211 6288 26243
rect 6328 26211 6360 26243
rect 6400 26211 6432 26243
rect 6472 26211 6504 26243
rect 6544 26211 6576 26243
rect 6616 26211 6648 26243
rect 6688 26211 6720 26243
rect 6760 26211 6792 26243
rect 6832 26211 6864 26243
rect 6904 26211 6936 26243
rect 6976 26211 7008 26243
rect 7048 26211 7080 26243
rect 7120 26211 7152 26243
rect 7192 26211 7224 26243
rect 7264 26211 7296 26243
rect 7336 26211 7368 26243
rect 7408 26211 7440 26243
rect 7480 26211 7512 26243
rect 7552 26211 7584 26243
rect 7624 26211 7656 26243
rect 7696 26211 7728 26243
rect 7768 26211 7800 26243
rect 7840 26211 7872 26243
rect 7912 26211 7944 26243
rect 7984 26211 8016 26243
rect 8056 26211 8088 26243
rect 8128 26211 8160 26243
rect 8200 26211 8232 26243
rect 8272 26211 8304 26243
rect 8344 26211 8376 26243
rect 8416 26211 8448 26243
rect 8488 26211 8520 26243
rect 8560 26211 8592 26243
rect 8632 26211 8664 26243
rect 8704 26211 8736 26243
rect 8776 26211 8808 26243
rect 8848 26211 8880 26243
rect 8920 26211 8952 26243
rect 8992 26211 9024 26243
rect 9064 26211 9096 26243
rect 9136 26211 9168 26243
rect 9208 26211 9240 26243
rect 9280 26211 9312 26243
rect 9352 26211 9384 26243
rect 9424 26211 9456 26243
rect 9496 26211 9528 26243
rect 9568 26211 9600 26243
rect 9640 26211 9672 26243
rect 9712 26211 9744 26243
rect 9784 26211 9816 26243
rect 9856 26211 9888 26243
rect 9928 26211 9960 26243
rect 10000 26211 10032 26243
rect 10072 26211 10104 26243
rect 10144 26211 10176 26243
rect 10216 26211 10248 26243
rect 10288 26211 10320 26243
rect 10360 26211 10392 26243
rect 10432 26211 10464 26243
rect 10504 26211 10536 26243
rect 10576 26211 10608 26243
rect 10648 26211 10680 26243
rect 10720 26211 10752 26243
rect 10792 26211 10824 26243
rect 10864 26211 10896 26243
rect 10936 26211 10968 26243
rect 11008 26211 11040 26243
rect 11080 26211 11112 26243
rect 11152 26211 11184 26243
rect 11224 26211 11256 26243
rect 11296 26211 11328 26243
rect 11368 26211 11400 26243
rect 11440 26211 11472 26243
rect 11512 26211 11544 26243
rect 11584 26211 11616 26243
rect 11656 26211 11688 26243
rect 11728 26211 11760 26243
rect 11800 26211 11832 26243
rect 11872 26211 11904 26243
rect 11944 26211 11976 26243
rect 12016 26211 12048 26243
rect 12088 26211 12120 26243
rect 12160 26211 12192 26243
rect 12232 26211 12264 26243
rect 12304 26211 12336 26243
rect 12376 26211 12408 26243
rect 12448 26211 12480 26243
rect 12520 26211 12552 26243
rect 12592 26211 12624 26243
rect 12664 26211 12696 26243
rect 12736 26211 12768 26243
rect 12808 26211 12840 26243
rect 12880 26211 12912 26243
rect 12952 26211 12984 26243
rect 13024 26211 13056 26243
rect 13096 26211 13128 26243
rect 13168 26211 13200 26243
rect 13240 26211 13272 26243
rect 13312 26211 13344 26243
rect 13384 26211 13416 26243
rect 13456 26211 13488 26243
rect 13528 26211 13560 26243
rect 13600 26211 13632 26243
rect 13672 26211 13704 26243
rect 13744 26211 13776 26243
rect 13816 26211 13848 26243
rect 13888 26211 13920 26243
rect 13960 26211 13992 26243
rect 14032 26211 14064 26243
rect 14104 26211 14136 26243
rect 14176 26211 14208 26243
rect 14248 26211 14280 26243
rect 14320 26211 14352 26243
rect 14392 26211 14424 26243
rect 14464 26211 14496 26243
rect 14536 26211 14568 26243
rect 14608 26211 14640 26243
rect 14680 26211 14712 26243
rect 14752 26211 14784 26243
rect 14824 26211 14856 26243
rect 14896 26211 14928 26243
rect 14968 26211 15000 26243
rect 15040 26211 15072 26243
rect 15112 26211 15144 26243
rect 15184 26211 15216 26243
rect 15256 26211 15288 26243
rect 15328 26211 15360 26243
rect 15400 26211 15432 26243
rect 15472 26211 15504 26243
rect 15544 26211 15576 26243
rect 15616 26211 15648 26243
rect 15688 26211 15720 26243
rect 15760 26211 15792 26243
rect 15832 26211 15864 26243
rect 15904 26211 15936 26243
rect 64 26139 96 26171
rect 136 26139 168 26171
rect 208 26139 240 26171
rect 280 26139 312 26171
rect 352 26139 384 26171
rect 424 26139 456 26171
rect 496 26139 528 26171
rect 568 26139 600 26171
rect 640 26139 672 26171
rect 712 26139 744 26171
rect 784 26139 816 26171
rect 856 26139 888 26171
rect 928 26139 960 26171
rect 1000 26139 1032 26171
rect 1072 26139 1104 26171
rect 1144 26139 1176 26171
rect 1216 26139 1248 26171
rect 1288 26139 1320 26171
rect 1360 26139 1392 26171
rect 1432 26139 1464 26171
rect 1504 26139 1536 26171
rect 1576 26139 1608 26171
rect 1648 26139 1680 26171
rect 1720 26139 1752 26171
rect 1792 26139 1824 26171
rect 1864 26139 1896 26171
rect 1936 26139 1968 26171
rect 2008 26139 2040 26171
rect 2080 26139 2112 26171
rect 2152 26139 2184 26171
rect 2224 26139 2256 26171
rect 2296 26139 2328 26171
rect 2368 26139 2400 26171
rect 2440 26139 2472 26171
rect 2512 26139 2544 26171
rect 2584 26139 2616 26171
rect 2656 26139 2688 26171
rect 2728 26139 2760 26171
rect 2800 26139 2832 26171
rect 2872 26139 2904 26171
rect 2944 26139 2976 26171
rect 3016 26139 3048 26171
rect 3088 26139 3120 26171
rect 3160 26139 3192 26171
rect 3232 26139 3264 26171
rect 3304 26139 3336 26171
rect 3376 26139 3408 26171
rect 3448 26139 3480 26171
rect 3520 26139 3552 26171
rect 3592 26139 3624 26171
rect 3664 26139 3696 26171
rect 3736 26139 3768 26171
rect 3808 26139 3840 26171
rect 3880 26139 3912 26171
rect 3952 26139 3984 26171
rect 4024 26139 4056 26171
rect 4096 26139 4128 26171
rect 4168 26139 4200 26171
rect 4240 26139 4272 26171
rect 4312 26139 4344 26171
rect 4384 26139 4416 26171
rect 4456 26139 4488 26171
rect 4528 26139 4560 26171
rect 4600 26139 4632 26171
rect 4672 26139 4704 26171
rect 4744 26139 4776 26171
rect 4816 26139 4848 26171
rect 4888 26139 4920 26171
rect 4960 26139 4992 26171
rect 5032 26139 5064 26171
rect 5104 26139 5136 26171
rect 5176 26139 5208 26171
rect 5248 26139 5280 26171
rect 5320 26139 5352 26171
rect 5392 26139 5424 26171
rect 5464 26139 5496 26171
rect 5536 26139 5568 26171
rect 5608 26139 5640 26171
rect 5680 26139 5712 26171
rect 5752 26139 5784 26171
rect 5824 26139 5856 26171
rect 5896 26139 5928 26171
rect 5968 26139 6000 26171
rect 6040 26139 6072 26171
rect 6112 26139 6144 26171
rect 6184 26139 6216 26171
rect 6256 26139 6288 26171
rect 6328 26139 6360 26171
rect 6400 26139 6432 26171
rect 6472 26139 6504 26171
rect 6544 26139 6576 26171
rect 6616 26139 6648 26171
rect 6688 26139 6720 26171
rect 6760 26139 6792 26171
rect 6832 26139 6864 26171
rect 6904 26139 6936 26171
rect 6976 26139 7008 26171
rect 7048 26139 7080 26171
rect 7120 26139 7152 26171
rect 7192 26139 7224 26171
rect 7264 26139 7296 26171
rect 7336 26139 7368 26171
rect 7408 26139 7440 26171
rect 7480 26139 7512 26171
rect 7552 26139 7584 26171
rect 7624 26139 7656 26171
rect 7696 26139 7728 26171
rect 7768 26139 7800 26171
rect 7840 26139 7872 26171
rect 7912 26139 7944 26171
rect 7984 26139 8016 26171
rect 8056 26139 8088 26171
rect 8128 26139 8160 26171
rect 8200 26139 8232 26171
rect 8272 26139 8304 26171
rect 8344 26139 8376 26171
rect 8416 26139 8448 26171
rect 8488 26139 8520 26171
rect 8560 26139 8592 26171
rect 8632 26139 8664 26171
rect 8704 26139 8736 26171
rect 8776 26139 8808 26171
rect 8848 26139 8880 26171
rect 8920 26139 8952 26171
rect 8992 26139 9024 26171
rect 9064 26139 9096 26171
rect 9136 26139 9168 26171
rect 9208 26139 9240 26171
rect 9280 26139 9312 26171
rect 9352 26139 9384 26171
rect 9424 26139 9456 26171
rect 9496 26139 9528 26171
rect 9568 26139 9600 26171
rect 9640 26139 9672 26171
rect 9712 26139 9744 26171
rect 9784 26139 9816 26171
rect 9856 26139 9888 26171
rect 9928 26139 9960 26171
rect 10000 26139 10032 26171
rect 10072 26139 10104 26171
rect 10144 26139 10176 26171
rect 10216 26139 10248 26171
rect 10288 26139 10320 26171
rect 10360 26139 10392 26171
rect 10432 26139 10464 26171
rect 10504 26139 10536 26171
rect 10576 26139 10608 26171
rect 10648 26139 10680 26171
rect 10720 26139 10752 26171
rect 10792 26139 10824 26171
rect 10864 26139 10896 26171
rect 10936 26139 10968 26171
rect 11008 26139 11040 26171
rect 11080 26139 11112 26171
rect 11152 26139 11184 26171
rect 11224 26139 11256 26171
rect 11296 26139 11328 26171
rect 11368 26139 11400 26171
rect 11440 26139 11472 26171
rect 11512 26139 11544 26171
rect 11584 26139 11616 26171
rect 11656 26139 11688 26171
rect 11728 26139 11760 26171
rect 11800 26139 11832 26171
rect 11872 26139 11904 26171
rect 11944 26139 11976 26171
rect 12016 26139 12048 26171
rect 12088 26139 12120 26171
rect 12160 26139 12192 26171
rect 12232 26139 12264 26171
rect 12304 26139 12336 26171
rect 12376 26139 12408 26171
rect 12448 26139 12480 26171
rect 12520 26139 12552 26171
rect 12592 26139 12624 26171
rect 12664 26139 12696 26171
rect 12736 26139 12768 26171
rect 12808 26139 12840 26171
rect 12880 26139 12912 26171
rect 12952 26139 12984 26171
rect 13024 26139 13056 26171
rect 13096 26139 13128 26171
rect 13168 26139 13200 26171
rect 13240 26139 13272 26171
rect 13312 26139 13344 26171
rect 13384 26139 13416 26171
rect 13456 26139 13488 26171
rect 13528 26139 13560 26171
rect 13600 26139 13632 26171
rect 13672 26139 13704 26171
rect 13744 26139 13776 26171
rect 13816 26139 13848 26171
rect 13888 26139 13920 26171
rect 13960 26139 13992 26171
rect 14032 26139 14064 26171
rect 14104 26139 14136 26171
rect 14176 26139 14208 26171
rect 14248 26139 14280 26171
rect 14320 26139 14352 26171
rect 14392 26139 14424 26171
rect 14464 26139 14496 26171
rect 14536 26139 14568 26171
rect 14608 26139 14640 26171
rect 14680 26139 14712 26171
rect 14752 26139 14784 26171
rect 14824 26139 14856 26171
rect 14896 26139 14928 26171
rect 14968 26139 15000 26171
rect 15040 26139 15072 26171
rect 15112 26139 15144 26171
rect 15184 26139 15216 26171
rect 15256 26139 15288 26171
rect 15328 26139 15360 26171
rect 15400 26139 15432 26171
rect 15472 26139 15504 26171
rect 15544 26139 15576 26171
rect 15616 26139 15648 26171
rect 15688 26139 15720 26171
rect 15760 26139 15792 26171
rect 15832 26139 15864 26171
rect 15904 26139 15936 26171
rect 64 26067 96 26099
rect 136 26067 168 26099
rect 208 26067 240 26099
rect 280 26067 312 26099
rect 352 26067 384 26099
rect 424 26067 456 26099
rect 496 26067 528 26099
rect 568 26067 600 26099
rect 640 26067 672 26099
rect 712 26067 744 26099
rect 784 26067 816 26099
rect 856 26067 888 26099
rect 928 26067 960 26099
rect 1000 26067 1032 26099
rect 1072 26067 1104 26099
rect 1144 26067 1176 26099
rect 1216 26067 1248 26099
rect 1288 26067 1320 26099
rect 1360 26067 1392 26099
rect 1432 26067 1464 26099
rect 1504 26067 1536 26099
rect 1576 26067 1608 26099
rect 1648 26067 1680 26099
rect 1720 26067 1752 26099
rect 1792 26067 1824 26099
rect 1864 26067 1896 26099
rect 1936 26067 1968 26099
rect 2008 26067 2040 26099
rect 2080 26067 2112 26099
rect 2152 26067 2184 26099
rect 2224 26067 2256 26099
rect 2296 26067 2328 26099
rect 2368 26067 2400 26099
rect 2440 26067 2472 26099
rect 2512 26067 2544 26099
rect 2584 26067 2616 26099
rect 2656 26067 2688 26099
rect 2728 26067 2760 26099
rect 2800 26067 2832 26099
rect 2872 26067 2904 26099
rect 2944 26067 2976 26099
rect 3016 26067 3048 26099
rect 3088 26067 3120 26099
rect 3160 26067 3192 26099
rect 3232 26067 3264 26099
rect 3304 26067 3336 26099
rect 3376 26067 3408 26099
rect 3448 26067 3480 26099
rect 3520 26067 3552 26099
rect 3592 26067 3624 26099
rect 3664 26067 3696 26099
rect 3736 26067 3768 26099
rect 3808 26067 3840 26099
rect 3880 26067 3912 26099
rect 3952 26067 3984 26099
rect 4024 26067 4056 26099
rect 4096 26067 4128 26099
rect 4168 26067 4200 26099
rect 4240 26067 4272 26099
rect 4312 26067 4344 26099
rect 4384 26067 4416 26099
rect 4456 26067 4488 26099
rect 4528 26067 4560 26099
rect 4600 26067 4632 26099
rect 4672 26067 4704 26099
rect 4744 26067 4776 26099
rect 4816 26067 4848 26099
rect 4888 26067 4920 26099
rect 4960 26067 4992 26099
rect 5032 26067 5064 26099
rect 5104 26067 5136 26099
rect 5176 26067 5208 26099
rect 5248 26067 5280 26099
rect 5320 26067 5352 26099
rect 5392 26067 5424 26099
rect 5464 26067 5496 26099
rect 5536 26067 5568 26099
rect 5608 26067 5640 26099
rect 5680 26067 5712 26099
rect 5752 26067 5784 26099
rect 5824 26067 5856 26099
rect 5896 26067 5928 26099
rect 5968 26067 6000 26099
rect 6040 26067 6072 26099
rect 6112 26067 6144 26099
rect 6184 26067 6216 26099
rect 6256 26067 6288 26099
rect 6328 26067 6360 26099
rect 6400 26067 6432 26099
rect 6472 26067 6504 26099
rect 6544 26067 6576 26099
rect 6616 26067 6648 26099
rect 6688 26067 6720 26099
rect 6760 26067 6792 26099
rect 6832 26067 6864 26099
rect 6904 26067 6936 26099
rect 6976 26067 7008 26099
rect 7048 26067 7080 26099
rect 7120 26067 7152 26099
rect 7192 26067 7224 26099
rect 7264 26067 7296 26099
rect 7336 26067 7368 26099
rect 7408 26067 7440 26099
rect 7480 26067 7512 26099
rect 7552 26067 7584 26099
rect 7624 26067 7656 26099
rect 7696 26067 7728 26099
rect 7768 26067 7800 26099
rect 7840 26067 7872 26099
rect 7912 26067 7944 26099
rect 7984 26067 8016 26099
rect 8056 26067 8088 26099
rect 8128 26067 8160 26099
rect 8200 26067 8232 26099
rect 8272 26067 8304 26099
rect 8344 26067 8376 26099
rect 8416 26067 8448 26099
rect 8488 26067 8520 26099
rect 8560 26067 8592 26099
rect 8632 26067 8664 26099
rect 8704 26067 8736 26099
rect 8776 26067 8808 26099
rect 8848 26067 8880 26099
rect 8920 26067 8952 26099
rect 8992 26067 9024 26099
rect 9064 26067 9096 26099
rect 9136 26067 9168 26099
rect 9208 26067 9240 26099
rect 9280 26067 9312 26099
rect 9352 26067 9384 26099
rect 9424 26067 9456 26099
rect 9496 26067 9528 26099
rect 9568 26067 9600 26099
rect 9640 26067 9672 26099
rect 9712 26067 9744 26099
rect 9784 26067 9816 26099
rect 9856 26067 9888 26099
rect 9928 26067 9960 26099
rect 10000 26067 10032 26099
rect 10072 26067 10104 26099
rect 10144 26067 10176 26099
rect 10216 26067 10248 26099
rect 10288 26067 10320 26099
rect 10360 26067 10392 26099
rect 10432 26067 10464 26099
rect 10504 26067 10536 26099
rect 10576 26067 10608 26099
rect 10648 26067 10680 26099
rect 10720 26067 10752 26099
rect 10792 26067 10824 26099
rect 10864 26067 10896 26099
rect 10936 26067 10968 26099
rect 11008 26067 11040 26099
rect 11080 26067 11112 26099
rect 11152 26067 11184 26099
rect 11224 26067 11256 26099
rect 11296 26067 11328 26099
rect 11368 26067 11400 26099
rect 11440 26067 11472 26099
rect 11512 26067 11544 26099
rect 11584 26067 11616 26099
rect 11656 26067 11688 26099
rect 11728 26067 11760 26099
rect 11800 26067 11832 26099
rect 11872 26067 11904 26099
rect 11944 26067 11976 26099
rect 12016 26067 12048 26099
rect 12088 26067 12120 26099
rect 12160 26067 12192 26099
rect 12232 26067 12264 26099
rect 12304 26067 12336 26099
rect 12376 26067 12408 26099
rect 12448 26067 12480 26099
rect 12520 26067 12552 26099
rect 12592 26067 12624 26099
rect 12664 26067 12696 26099
rect 12736 26067 12768 26099
rect 12808 26067 12840 26099
rect 12880 26067 12912 26099
rect 12952 26067 12984 26099
rect 13024 26067 13056 26099
rect 13096 26067 13128 26099
rect 13168 26067 13200 26099
rect 13240 26067 13272 26099
rect 13312 26067 13344 26099
rect 13384 26067 13416 26099
rect 13456 26067 13488 26099
rect 13528 26067 13560 26099
rect 13600 26067 13632 26099
rect 13672 26067 13704 26099
rect 13744 26067 13776 26099
rect 13816 26067 13848 26099
rect 13888 26067 13920 26099
rect 13960 26067 13992 26099
rect 14032 26067 14064 26099
rect 14104 26067 14136 26099
rect 14176 26067 14208 26099
rect 14248 26067 14280 26099
rect 14320 26067 14352 26099
rect 14392 26067 14424 26099
rect 14464 26067 14496 26099
rect 14536 26067 14568 26099
rect 14608 26067 14640 26099
rect 14680 26067 14712 26099
rect 14752 26067 14784 26099
rect 14824 26067 14856 26099
rect 14896 26067 14928 26099
rect 14968 26067 15000 26099
rect 15040 26067 15072 26099
rect 15112 26067 15144 26099
rect 15184 26067 15216 26099
rect 15256 26067 15288 26099
rect 15328 26067 15360 26099
rect 15400 26067 15432 26099
rect 15472 26067 15504 26099
rect 15544 26067 15576 26099
rect 15616 26067 15648 26099
rect 15688 26067 15720 26099
rect 15760 26067 15792 26099
rect 15832 26067 15864 26099
rect 15904 26067 15936 26099
rect 64 25995 96 26027
rect 136 25995 168 26027
rect 208 25995 240 26027
rect 280 25995 312 26027
rect 352 25995 384 26027
rect 424 25995 456 26027
rect 496 25995 528 26027
rect 568 25995 600 26027
rect 640 25995 672 26027
rect 712 25995 744 26027
rect 784 25995 816 26027
rect 856 25995 888 26027
rect 928 25995 960 26027
rect 1000 25995 1032 26027
rect 1072 25995 1104 26027
rect 1144 25995 1176 26027
rect 1216 25995 1248 26027
rect 1288 25995 1320 26027
rect 1360 25995 1392 26027
rect 1432 25995 1464 26027
rect 1504 25995 1536 26027
rect 1576 25995 1608 26027
rect 1648 25995 1680 26027
rect 1720 25995 1752 26027
rect 1792 25995 1824 26027
rect 1864 25995 1896 26027
rect 1936 25995 1968 26027
rect 2008 25995 2040 26027
rect 2080 25995 2112 26027
rect 2152 25995 2184 26027
rect 2224 25995 2256 26027
rect 2296 25995 2328 26027
rect 2368 25995 2400 26027
rect 2440 25995 2472 26027
rect 2512 25995 2544 26027
rect 2584 25995 2616 26027
rect 2656 25995 2688 26027
rect 2728 25995 2760 26027
rect 2800 25995 2832 26027
rect 2872 25995 2904 26027
rect 2944 25995 2976 26027
rect 3016 25995 3048 26027
rect 3088 25995 3120 26027
rect 3160 25995 3192 26027
rect 3232 25995 3264 26027
rect 3304 25995 3336 26027
rect 3376 25995 3408 26027
rect 3448 25995 3480 26027
rect 3520 25995 3552 26027
rect 3592 25995 3624 26027
rect 3664 25995 3696 26027
rect 3736 25995 3768 26027
rect 3808 25995 3840 26027
rect 3880 25995 3912 26027
rect 3952 25995 3984 26027
rect 4024 25995 4056 26027
rect 4096 25995 4128 26027
rect 4168 25995 4200 26027
rect 4240 25995 4272 26027
rect 4312 25995 4344 26027
rect 4384 25995 4416 26027
rect 4456 25995 4488 26027
rect 4528 25995 4560 26027
rect 4600 25995 4632 26027
rect 4672 25995 4704 26027
rect 4744 25995 4776 26027
rect 4816 25995 4848 26027
rect 4888 25995 4920 26027
rect 4960 25995 4992 26027
rect 5032 25995 5064 26027
rect 5104 25995 5136 26027
rect 5176 25995 5208 26027
rect 5248 25995 5280 26027
rect 5320 25995 5352 26027
rect 5392 25995 5424 26027
rect 5464 25995 5496 26027
rect 5536 25995 5568 26027
rect 5608 25995 5640 26027
rect 5680 25995 5712 26027
rect 5752 25995 5784 26027
rect 5824 25995 5856 26027
rect 5896 25995 5928 26027
rect 5968 25995 6000 26027
rect 6040 25995 6072 26027
rect 6112 25995 6144 26027
rect 6184 25995 6216 26027
rect 6256 25995 6288 26027
rect 6328 25995 6360 26027
rect 6400 25995 6432 26027
rect 6472 25995 6504 26027
rect 6544 25995 6576 26027
rect 6616 25995 6648 26027
rect 6688 25995 6720 26027
rect 6760 25995 6792 26027
rect 6832 25995 6864 26027
rect 6904 25995 6936 26027
rect 6976 25995 7008 26027
rect 7048 25995 7080 26027
rect 7120 25995 7152 26027
rect 7192 25995 7224 26027
rect 7264 25995 7296 26027
rect 7336 25995 7368 26027
rect 7408 25995 7440 26027
rect 7480 25995 7512 26027
rect 7552 25995 7584 26027
rect 7624 25995 7656 26027
rect 7696 25995 7728 26027
rect 7768 25995 7800 26027
rect 7840 25995 7872 26027
rect 7912 25995 7944 26027
rect 7984 25995 8016 26027
rect 8056 25995 8088 26027
rect 8128 25995 8160 26027
rect 8200 25995 8232 26027
rect 8272 25995 8304 26027
rect 8344 25995 8376 26027
rect 8416 25995 8448 26027
rect 8488 25995 8520 26027
rect 8560 25995 8592 26027
rect 8632 25995 8664 26027
rect 8704 25995 8736 26027
rect 8776 25995 8808 26027
rect 8848 25995 8880 26027
rect 8920 25995 8952 26027
rect 8992 25995 9024 26027
rect 9064 25995 9096 26027
rect 9136 25995 9168 26027
rect 9208 25995 9240 26027
rect 9280 25995 9312 26027
rect 9352 25995 9384 26027
rect 9424 25995 9456 26027
rect 9496 25995 9528 26027
rect 9568 25995 9600 26027
rect 9640 25995 9672 26027
rect 9712 25995 9744 26027
rect 9784 25995 9816 26027
rect 9856 25995 9888 26027
rect 9928 25995 9960 26027
rect 10000 25995 10032 26027
rect 10072 25995 10104 26027
rect 10144 25995 10176 26027
rect 10216 25995 10248 26027
rect 10288 25995 10320 26027
rect 10360 25995 10392 26027
rect 10432 25995 10464 26027
rect 10504 25995 10536 26027
rect 10576 25995 10608 26027
rect 10648 25995 10680 26027
rect 10720 25995 10752 26027
rect 10792 25995 10824 26027
rect 10864 25995 10896 26027
rect 10936 25995 10968 26027
rect 11008 25995 11040 26027
rect 11080 25995 11112 26027
rect 11152 25995 11184 26027
rect 11224 25995 11256 26027
rect 11296 25995 11328 26027
rect 11368 25995 11400 26027
rect 11440 25995 11472 26027
rect 11512 25995 11544 26027
rect 11584 25995 11616 26027
rect 11656 25995 11688 26027
rect 11728 25995 11760 26027
rect 11800 25995 11832 26027
rect 11872 25995 11904 26027
rect 11944 25995 11976 26027
rect 12016 25995 12048 26027
rect 12088 25995 12120 26027
rect 12160 25995 12192 26027
rect 12232 25995 12264 26027
rect 12304 25995 12336 26027
rect 12376 25995 12408 26027
rect 12448 25995 12480 26027
rect 12520 25995 12552 26027
rect 12592 25995 12624 26027
rect 12664 25995 12696 26027
rect 12736 25995 12768 26027
rect 12808 25995 12840 26027
rect 12880 25995 12912 26027
rect 12952 25995 12984 26027
rect 13024 25995 13056 26027
rect 13096 25995 13128 26027
rect 13168 25995 13200 26027
rect 13240 25995 13272 26027
rect 13312 25995 13344 26027
rect 13384 25995 13416 26027
rect 13456 25995 13488 26027
rect 13528 25995 13560 26027
rect 13600 25995 13632 26027
rect 13672 25995 13704 26027
rect 13744 25995 13776 26027
rect 13816 25995 13848 26027
rect 13888 25995 13920 26027
rect 13960 25995 13992 26027
rect 14032 25995 14064 26027
rect 14104 25995 14136 26027
rect 14176 25995 14208 26027
rect 14248 25995 14280 26027
rect 14320 25995 14352 26027
rect 14392 25995 14424 26027
rect 14464 25995 14496 26027
rect 14536 25995 14568 26027
rect 14608 25995 14640 26027
rect 14680 25995 14712 26027
rect 14752 25995 14784 26027
rect 14824 25995 14856 26027
rect 14896 25995 14928 26027
rect 14968 25995 15000 26027
rect 15040 25995 15072 26027
rect 15112 25995 15144 26027
rect 15184 25995 15216 26027
rect 15256 25995 15288 26027
rect 15328 25995 15360 26027
rect 15400 25995 15432 26027
rect 15472 25995 15504 26027
rect 15544 25995 15576 26027
rect 15616 25995 15648 26027
rect 15688 25995 15720 26027
rect 15760 25995 15792 26027
rect 15832 25995 15864 26027
rect 15904 25995 15936 26027
rect 64 25923 96 25955
rect 136 25923 168 25955
rect 208 25923 240 25955
rect 280 25923 312 25955
rect 352 25923 384 25955
rect 424 25923 456 25955
rect 496 25923 528 25955
rect 568 25923 600 25955
rect 640 25923 672 25955
rect 712 25923 744 25955
rect 784 25923 816 25955
rect 856 25923 888 25955
rect 928 25923 960 25955
rect 1000 25923 1032 25955
rect 1072 25923 1104 25955
rect 1144 25923 1176 25955
rect 1216 25923 1248 25955
rect 1288 25923 1320 25955
rect 1360 25923 1392 25955
rect 1432 25923 1464 25955
rect 1504 25923 1536 25955
rect 1576 25923 1608 25955
rect 1648 25923 1680 25955
rect 1720 25923 1752 25955
rect 1792 25923 1824 25955
rect 1864 25923 1896 25955
rect 1936 25923 1968 25955
rect 2008 25923 2040 25955
rect 2080 25923 2112 25955
rect 2152 25923 2184 25955
rect 2224 25923 2256 25955
rect 2296 25923 2328 25955
rect 2368 25923 2400 25955
rect 2440 25923 2472 25955
rect 2512 25923 2544 25955
rect 2584 25923 2616 25955
rect 2656 25923 2688 25955
rect 2728 25923 2760 25955
rect 2800 25923 2832 25955
rect 2872 25923 2904 25955
rect 2944 25923 2976 25955
rect 3016 25923 3048 25955
rect 3088 25923 3120 25955
rect 3160 25923 3192 25955
rect 3232 25923 3264 25955
rect 3304 25923 3336 25955
rect 3376 25923 3408 25955
rect 3448 25923 3480 25955
rect 3520 25923 3552 25955
rect 3592 25923 3624 25955
rect 3664 25923 3696 25955
rect 3736 25923 3768 25955
rect 3808 25923 3840 25955
rect 3880 25923 3912 25955
rect 3952 25923 3984 25955
rect 4024 25923 4056 25955
rect 4096 25923 4128 25955
rect 4168 25923 4200 25955
rect 4240 25923 4272 25955
rect 4312 25923 4344 25955
rect 4384 25923 4416 25955
rect 4456 25923 4488 25955
rect 4528 25923 4560 25955
rect 4600 25923 4632 25955
rect 4672 25923 4704 25955
rect 4744 25923 4776 25955
rect 4816 25923 4848 25955
rect 4888 25923 4920 25955
rect 4960 25923 4992 25955
rect 5032 25923 5064 25955
rect 5104 25923 5136 25955
rect 5176 25923 5208 25955
rect 5248 25923 5280 25955
rect 5320 25923 5352 25955
rect 5392 25923 5424 25955
rect 5464 25923 5496 25955
rect 5536 25923 5568 25955
rect 5608 25923 5640 25955
rect 5680 25923 5712 25955
rect 5752 25923 5784 25955
rect 5824 25923 5856 25955
rect 5896 25923 5928 25955
rect 5968 25923 6000 25955
rect 6040 25923 6072 25955
rect 6112 25923 6144 25955
rect 6184 25923 6216 25955
rect 6256 25923 6288 25955
rect 6328 25923 6360 25955
rect 6400 25923 6432 25955
rect 6472 25923 6504 25955
rect 6544 25923 6576 25955
rect 6616 25923 6648 25955
rect 6688 25923 6720 25955
rect 6760 25923 6792 25955
rect 6832 25923 6864 25955
rect 6904 25923 6936 25955
rect 6976 25923 7008 25955
rect 7048 25923 7080 25955
rect 7120 25923 7152 25955
rect 7192 25923 7224 25955
rect 7264 25923 7296 25955
rect 7336 25923 7368 25955
rect 7408 25923 7440 25955
rect 7480 25923 7512 25955
rect 7552 25923 7584 25955
rect 7624 25923 7656 25955
rect 7696 25923 7728 25955
rect 7768 25923 7800 25955
rect 7840 25923 7872 25955
rect 7912 25923 7944 25955
rect 7984 25923 8016 25955
rect 8056 25923 8088 25955
rect 8128 25923 8160 25955
rect 8200 25923 8232 25955
rect 8272 25923 8304 25955
rect 8344 25923 8376 25955
rect 8416 25923 8448 25955
rect 8488 25923 8520 25955
rect 8560 25923 8592 25955
rect 8632 25923 8664 25955
rect 8704 25923 8736 25955
rect 8776 25923 8808 25955
rect 8848 25923 8880 25955
rect 8920 25923 8952 25955
rect 8992 25923 9024 25955
rect 9064 25923 9096 25955
rect 9136 25923 9168 25955
rect 9208 25923 9240 25955
rect 9280 25923 9312 25955
rect 9352 25923 9384 25955
rect 9424 25923 9456 25955
rect 9496 25923 9528 25955
rect 9568 25923 9600 25955
rect 9640 25923 9672 25955
rect 9712 25923 9744 25955
rect 9784 25923 9816 25955
rect 9856 25923 9888 25955
rect 9928 25923 9960 25955
rect 10000 25923 10032 25955
rect 10072 25923 10104 25955
rect 10144 25923 10176 25955
rect 10216 25923 10248 25955
rect 10288 25923 10320 25955
rect 10360 25923 10392 25955
rect 10432 25923 10464 25955
rect 10504 25923 10536 25955
rect 10576 25923 10608 25955
rect 10648 25923 10680 25955
rect 10720 25923 10752 25955
rect 10792 25923 10824 25955
rect 10864 25923 10896 25955
rect 10936 25923 10968 25955
rect 11008 25923 11040 25955
rect 11080 25923 11112 25955
rect 11152 25923 11184 25955
rect 11224 25923 11256 25955
rect 11296 25923 11328 25955
rect 11368 25923 11400 25955
rect 11440 25923 11472 25955
rect 11512 25923 11544 25955
rect 11584 25923 11616 25955
rect 11656 25923 11688 25955
rect 11728 25923 11760 25955
rect 11800 25923 11832 25955
rect 11872 25923 11904 25955
rect 11944 25923 11976 25955
rect 12016 25923 12048 25955
rect 12088 25923 12120 25955
rect 12160 25923 12192 25955
rect 12232 25923 12264 25955
rect 12304 25923 12336 25955
rect 12376 25923 12408 25955
rect 12448 25923 12480 25955
rect 12520 25923 12552 25955
rect 12592 25923 12624 25955
rect 12664 25923 12696 25955
rect 12736 25923 12768 25955
rect 12808 25923 12840 25955
rect 12880 25923 12912 25955
rect 12952 25923 12984 25955
rect 13024 25923 13056 25955
rect 13096 25923 13128 25955
rect 13168 25923 13200 25955
rect 13240 25923 13272 25955
rect 13312 25923 13344 25955
rect 13384 25923 13416 25955
rect 13456 25923 13488 25955
rect 13528 25923 13560 25955
rect 13600 25923 13632 25955
rect 13672 25923 13704 25955
rect 13744 25923 13776 25955
rect 13816 25923 13848 25955
rect 13888 25923 13920 25955
rect 13960 25923 13992 25955
rect 14032 25923 14064 25955
rect 14104 25923 14136 25955
rect 14176 25923 14208 25955
rect 14248 25923 14280 25955
rect 14320 25923 14352 25955
rect 14392 25923 14424 25955
rect 14464 25923 14496 25955
rect 14536 25923 14568 25955
rect 14608 25923 14640 25955
rect 14680 25923 14712 25955
rect 14752 25923 14784 25955
rect 14824 25923 14856 25955
rect 14896 25923 14928 25955
rect 14968 25923 15000 25955
rect 15040 25923 15072 25955
rect 15112 25923 15144 25955
rect 15184 25923 15216 25955
rect 15256 25923 15288 25955
rect 15328 25923 15360 25955
rect 15400 25923 15432 25955
rect 15472 25923 15504 25955
rect 15544 25923 15576 25955
rect 15616 25923 15648 25955
rect 15688 25923 15720 25955
rect 15760 25923 15792 25955
rect 15832 25923 15864 25955
rect 15904 25923 15936 25955
rect 64 25851 96 25883
rect 136 25851 168 25883
rect 208 25851 240 25883
rect 280 25851 312 25883
rect 352 25851 384 25883
rect 424 25851 456 25883
rect 496 25851 528 25883
rect 568 25851 600 25883
rect 640 25851 672 25883
rect 712 25851 744 25883
rect 784 25851 816 25883
rect 856 25851 888 25883
rect 928 25851 960 25883
rect 1000 25851 1032 25883
rect 1072 25851 1104 25883
rect 1144 25851 1176 25883
rect 1216 25851 1248 25883
rect 1288 25851 1320 25883
rect 1360 25851 1392 25883
rect 1432 25851 1464 25883
rect 1504 25851 1536 25883
rect 1576 25851 1608 25883
rect 1648 25851 1680 25883
rect 1720 25851 1752 25883
rect 1792 25851 1824 25883
rect 1864 25851 1896 25883
rect 1936 25851 1968 25883
rect 2008 25851 2040 25883
rect 2080 25851 2112 25883
rect 2152 25851 2184 25883
rect 2224 25851 2256 25883
rect 2296 25851 2328 25883
rect 2368 25851 2400 25883
rect 2440 25851 2472 25883
rect 2512 25851 2544 25883
rect 2584 25851 2616 25883
rect 2656 25851 2688 25883
rect 2728 25851 2760 25883
rect 2800 25851 2832 25883
rect 2872 25851 2904 25883
rect 2944 25851 2976 25883
rect 3016 25851 3048 25883
rect 3088 25851 3120 25883
rect 3160 25851 3192 25883
rect 3232 25851 3264 25883
rect 3304 25851 3336 25883
rect 3376 25851 3408 25883
rect 3448 25851 3480 25883
rect 3520 25851 3552 25883
rect 3592 25851 3624 25883
rect 3664 25851 3696 25883
rect 3736 25851 3768 25883
rect 3808 25851 3840 25883
rect 3880 25851 3912 25883
rect 3952 25851 3984 25883
rect 4024 25851 4056 25883
rect 4096 25851 4128 25883
rect 4168 25851 4200 25883
rect 4240 25851 4272 25883
rect 4312 25851 4344 25883
rect 4384 25851 4416 25883
rect 4456 25851 4488 25883
rect 4528 25851 4560 25883
rect 4600 25851 4632 25883
rect 4672 25851 4704 25883
rect 4744 25851 4776 25883
rect 4816 25851 4848 25883
rect 4888 25851 4920 25883
rect 4960 25851 4992 25883
rect 5032 25851 5064 25883
rect 5104 25851 5136 25883
rect 5176 25851 5208 25883
rect 5248 25851 5280 25883
rect 5320 25851 5352 25883
rect 5392 25851 5424 25883
rect 5464 25851 5496 25883
rect 5536 25851 5568 25883
rect 5608 25851 5640 25883
rect 5680 25851 5712 25883
rect 5752 25851 5784 25883
rect 5824 25851 5856 25883
rect 5896 25851 5928 25883
rect 5968 25851 6000 25883
rect 6040 25851 6072 25883
rect 6112 25851 6144 25883
rect 6184 25851 6216 25883
rect 6256 25851 6288 25883
rect 6328 25851 6360 25883
rect 6400 25851 6432 25883
rect 6472 25851 6504 25883
rect 6544 25851 6576 25883
rect 6616 25851 6648 25883
rect 6688 25851 6720 25883
rect 6760 25851 6792 25883
rect 6832 25851 6864 25883
rect 6904 25851 6936 25883
rect 6976 25851 7008 25883
rect 7048 25851 7080 25883
rect 7120 25851 7152 25883
rect 7192 25851 7224 25883
rect 7264 25851 7296 25883
rect 7336 25851 7368 25883
rect 7408 25851 7440 25883
rect 7480 25851 7512 25883
rect 7552 25851 7584 25883
rect 7624 25851 7656 25883
rect 7696 25851 7728 25883
rect 7768 25851 7800 25883
rect 7840 25851 7872 25883
rect 7912 25851 7944 25883
rect 7984 25851 8016 25883
rect 8056 25851 8088 25883
rect 8128 25851 8160 25883
rect 8200 25851 8232 25883
rect 8272 25851 8304 25883
rect 8344 25851 8376 25883
rect 8416 25851 8448 25883
rect 8488 25851 8520 25883
rect 8560 25851 8592 25883
rect 8632 25851 8664 25883
rect 8704 25851 8736 25883
rect 8776 25851 8808 25883
rect 8848 25851 8880 25883
rect 8920 25851 8952 25883
rect 8992 25851 9024 25883
rect 9064 25851 9096 25883
rect 9136 25851 9168 25883
rect 9208 25851 9240 25883
rect 9280 25851 9312 25883
rect 9352 25851 9384 25883
rect 9424 25851 9456 25883
rect 9496 25851 9528 25883
rect 9568 25851 9600 25883
rect 9640 25851 9672 25883
rect 9712 25851 9744 25883
rect 9784 25851 9816 25883
rect 9856 25851 9888 25883
rect 9928 25851 9960 25883
rect 10000 25851 10032 25883
rect 10072 25851 10104 25883
rect 10144 25851 10176 25883
rect 10216 25851 10248 25883
rect 10288 25851 10320 25883
rect 10360 25851 10392 25883
rect 10432 25851 10464 25883
rect 10504 25851 10536 25883
rect 10576 25851 10608 25883
rect 10648 25851 10680 25883
rect 10720 25851 10752 25883
rect 10792 25851 10824 25883
rect 10864 25851 10896 25883
rect 10936 25851 10968 25883
rect 11008 25851 11040 25883
rect 11080 25851 11112 25883
rect 11152 25851 11184 25883
rect 11224 25851 11256 25883
rect 11296 25851 11328 25883
rect 11368 25851 11400 25883
rect 11440 25851 11472 25883
rect 11512 25851 11544 25883
rect 11584 25851 11616 25883
rect 11656 25851 11688 25883
rect 11728 25851 11760 25883
rect 11800 25851 11832 25883
rect 11872 25851 11904 25883
rect 11944 25851 11976 25883
rect 12016 25851 12048 25883
rect 12088 25851 12120 25883
rect 12160 25851 12192 25883
rect 12232 25851 12264 25883
rect 12304 25851 12336 25883
rect 12376 25851 12408 25883
rect 12448 25851 12480 25883
rect 12520 25851 12552 25883
rect 12592 25851 12624 25883
rect 12664 25851 12696 25883
rect 12736 25851 12768 25883
rect 12808 25851 12840 25883
rect 12880 25851 12912 25883
rect 12952 25851 12984 25883
rect 13024 25851 13056 25883
rect 13096 25851 13128 25883
rect 13168 25851 13200 25883
rect 13240 25851 13272 25883
rect 13312 25851 13344 25883
rect 13384 25851 13416 25883
rect 13456 25851 13488 25883
rect 13528 25851 13560 25883
rect 13600 25851 13632 25883
rect 13672 25851 13704 25883
rect 13744 25851 13776 25883
rect 13816 25851 13848 25883
rect 13888 25851 13920 25883
rect 13960 25851 13992 25883
rect 14032 25851 14064 25883
rect 14104 25851 14136 25883
rect 14176 25851 14208 25883
rect 14248 25851 14280 25883
rect 14320 25851 14352 25883
rect 14392 25851 14424 25883
rect 14464 25851 14496 25883
rect 14536 25851 14568 25883
rect 14608 25851 14640 25883
rect 14680 25851 14712 25883
rect 14752 25851 14784 25883
rect 14824 25851 14856 25883
rect 14896 25851 14928 25883
rect 14968 25851 15000 25883
rect 15040 25851 15072 25883
rect 15112 25851 15144 25883
rect 15184 25851 15216 25883
rect 15256 25851 15288 25883
rect 15328 25851 15360 25883
rect 15400 25851 15432 25883
rect 15472 25851 15504 25883
rect 15544 25851 15576 25883
rect 15616 25851 15648 25883
rect 15688 25851 15720 25883
rect 15760 25851 15792 25883
rect 15832 25851 15864 25883
rect 15904 25851 15936 25883
rect 64 25779 96 25811
rect 136 25779 168 25811
rect 208 25779 240 25811
rect 280 25779 312 25811
rect 352 25779 384 25811
rect 424 25779 456 25811
rect 496 25779 528 25811
rect 568 25779 600 25811
rect 640 25779 672 25811
rect 712 25779 744 25811
rect 784 25779 816 25811
rect 856 25779 888 25811
rect 928 25779 960 25811
rect 1000 25779 1032 25811
rect 1072 25779 1104 25811
rect 1144 25779 1176 25811
rect 1216 25779 1248 25811
rect 1288 25779 1320 25811
rect 1360 25779 1392 25811
rect 1432 25779 1464 25811
rect 1504 25779 1536 25811
rect 1576 25779 1608 25811
rect 1648 25779 1680 25811
rect 1720 25779 1752 25811
rect 1792 25779 1824 25811
rect 1864 25779 1896 25811
rect 1936 25779 1968 25811
rect 2008 25779 2040 25811
rect 2080 25779 2112 25811
rect 2152 25779 2184 25811
rect 2224 25779 2256 25811
rect 2296 25779 2328 25811
rect 2368 25779 2400 25811
rect 2440 25779 2472 25811
rect 2512 25779 2544 25811
rect 2584 25779 2616 25811
rect 2656 25779 2688 25811
rect 2728 25779 2760 25811
rect 2800 25779 2832 25811
rect 2872 25779 2904 25811
rect 2944 25779 2976 25811
rect 3016 25779 3048 25811
rect 3088 25779 3120 25811
rect 3160 25779 3192 25811
rect 3232 25779 3264 25811
rect 3304 25779 3336 25811
rect 3376 25779 3408 25811
rect 3448 25779 3480 25811
rect 3520 25779 3552 25811
rect 3592 25779 3624 25811
rect 3664 25779 3696 25811
rect 3736 25779 3768 25811
rect 3808 25779 3840 25811
rect 3880 25779 3912 25811
rect 3952 25779 3984 25811
rect 4024 25779 4056 25811
rect 4096 25779 4128 25811
rect 4168 25779 4200 25811
rect 4240 25779 4272 25811
rect 4312 25779 4344 25811
rect 4384 25779 4416 25811
rect 4456 25779 4488 25811
rect 4528 25779 4560 25811
rect 4600 25779 4632 25811
rect 4672 25779 4704 25811
rect 4744 25779 4776 25811
rect 4816 25779 4848 25811
rect 4888 25779 4920 25811
rect 4960 25779 4992 25811
rect 5032 25779 5064 25811
rect 5104 25779 5136 25811
rect 5176 25779 5208 25811
rect 5248 25779 5280 25811
rect 5320 25779 5352 25811
rect 5392 25779 5424 25811
rect 5464 25779 5496 25811
rect 5536 25779 5568 25811
rect 5608 25779 5640 25811
rect 5680 25779 5712 25811
rect 5752 25779 5784 25811
rect 5824 25779 5856 25811
rect 5896 25779 5928 25811
rect 5968 25779 6000 25811
rect 6040 25779 6072 25811
rect 6112 25779 6144 25811
rect 6184 25779 6216 25811
rect 6256 25779 6288 25811
rect 6328 25779 6360 25811
rect 6400 25779 6432 25811
rect 6472 25779 6504 25811
rect 6544 25779 6576 25811
rect 6616 25779 6648 25811
rect 6688 25779 6720 25811
rect 6760 25779 6792 25811
rect 6832 25779 6864 25811
rect 6904 25779 6936 25811
rect 6976 25779 7008 25811
rect 7048 25779 7080 25811
rect 7120 25779 7152 25811
rect 7192 25779 7224 25811
rect 7264 25779 7296 25811
rect 7336 25779 7368 25811
rect 7408 25779 7440 25811
rect 7480 25779 7512 25811
rect 7552 25779 7584 25811
rect 7624 25779 7656 25811
rect 7696 25779 7728 25811
rect 7768 25779 7800 25811
rect 7840 25779 7872 25811
rect 7912 25779 7944 25811
rect 7984 25779 8016 25811
rect 8056 25779 8088 25811
rect 8128 25779 8160 25811
rect 8200 25779 8232 25811
rect 8272 25779 8304 25811
rect 8344 25779 8376 25811
rect 8416 25779 8448 25811
rect 8488 25779 8520 25811
rect 8560 25779 8592 25811
rect 8632 25779 8664 25811
rect 8704 25779 8736 25811
rect 8776 25779 8808 25811
rect 8848 25779 8880 25811
rect 8920 25779 8952 25811
rect 8992 25779 9024 25811
rect 9064 25779 9096 25811
rect 9136 25779 9168 25811
rect 9208 25779 9240 25811
rect 9280 25779 9312 25811
rect 9352 25779 9384 25811
rect 9424 25779 9456 25811
rect 9496 25779 9528 25811
rect 9568 25779 9600 25811
rect 9640 25779 9672 25811
rect 9712 25779 9744 25811
rect 9784 25779 9816 25811
rect 9856 25779 9888 25811
rect 9928 25779 9960 25811
rect 10000 25779 10032 25811
rect 10072 25779 10104 25811
rect 10144 25779 10176 25811
rect 10216 25779 10248 25811
rect 10288 25779 10320 25811
rect 10360 25779 10392 25811
rect 10432 25779 10464 25811
rect 10504 25779 10536 25811
rect 10576 25779 10608 25811
rect 10648 25779 10680 25811
rect 10720 25779 10752 25811
rect 10792 25779 10824 25811
rect 10864 25779 10896 25811
rect 10936 25779 10968 25811
rect 11008 25779 11040 25811
rect 11080 25779 11112 25811
rect 11152 25779 11184 25811
rect 11224 25779 11256 25811
rect 11296 25779 11328 25811
rect 11368 25779 11400 25811
rect 11440 25779 11472 25811
rect 11512 25779 11544 25811
rect 11584 25779 11616 25811
rect 11656 25779 11688 25811
rect 11728 25779 11760 25811
rect 11800 25779 11832 25811
rect 11872 25779 11904 25811
rect 11944 25779 11976 25811
rect 12016 25779 12048 25811
rect 12088 25779 12120 25811
rect 12160 25779 12192 25811
rect 12232 25779 12264 25811
rect 12304 25779 12336 25811
rect 12376 25779 12408 25811
rect 12448 25779 12480 25811
rect 12520 25779 12552 25811
rect 12592 25779 12624 25811
rect 12664 25779 12696 25811
rect 12736 25779 12768 25811
rect 12808 25779 12840 25811
rect 12880 25779 12912 25811
rect 12952 25779 12984 25811
rect 13024 25779 13056 25811
rect 13096 25779 13128 25811
rect 13168 25779 13200 25811
rect 13240 25779 13272 25811
rect 13312 25779 13344 25811
rect 13384 25779 13416 25811
rect 13456 25779 13488 25811
rect 13528 25779 13560 25811
rect 13600 25779 13632 25811
rect 13672 25779 13704 25811
rect 13744 25779 13776 25811
rect 13816 25779 13848 25811
rect 13888 25779 13920 25811
rect 13960 25779 13992 25811
rect 14032 25779 14064 25811
rect 14104 25779 14136 25811
rect 14176 25779 14208 25811
rect 14248 25779 14280 25811
rect 14320 25779 14352 25811
rect 14392 25779 14424 25811
rect 14464 25779 14496 25811
rect 14536 25779 14568 25811
rect 14608 25779 14640 25811
rect 14680 25779 14712 25811
rect 14752 25779 14784 25811
rect 14824 25779 14856 25811
rect 14896 25779 14928 25811
rect 14968 25779 15000 25811
rect 15040 25779 15072 25811
rect 15112 25779 15144 25811
rect 15184 25779 15216 25811
rect 15256 25779 15288 25811
rect 15328 25779 15360 25811
rect 15400 25779 15432 25811
rect 15472 25779 15504 25811
rect 15544 25779 15576 25811
rect 15616 25779 15648 25811
rect 15688 25779 15720 25811
rect 15760 25779 15792 25811
rect 15832 25779 15864 25811
rect 15904 25779 15936 25811
rect 64 25707 96 25739
rect 136 25707 168 25739
rect 208 25707 240 25739
rect 280 25707 312 25739
rect 352 25707 384 25739
rect 424 25707 456 25739
rect 496 25707 528 25739
rect 568 25707 600 25739
rect 640 25707 672 25739
rect 712 25707 744 25739
rect 784 25707 816 25739
rect 856 25707 888 25739
rect 928 25707 960 25739
rect 1000 25707 1032 25739
rect 1072 25707 1104 25739
rect 1144 25707 1176 25739
rect 1216 25707 1248 25739
rect 1288 25707 1320 25739
rect 1360 25707 1392 25739
rect 1432 25707 1464 25739
rect 1504 25707 1536 25739
rect 1576 25707 1608 25739
rect 1648 25707 1680 25739
rect 1720 25707 1752 25739
rect 1792 25707 1824 25739
rect 1864 25707 1896 25739
rect 1936 25707 1968 25739
rect 2008 25707 2040 25739
rect 2080 25707 2112 25739
rect 2152 25707 2184 25739
rect 2224 25707 2256 25739
rect 2296 25707 2328 25739
rect 2368 25707 2400 25739
rect 2440 25707 2472 25739
rect 2512 25707 2544 25739
rect 2584 25707 2616 25739
rect 2656 25707 2688 25739
rect 2728 25707 2760 25739
rect 2800 25707 2832 25739
rect 2872 25707 2904 25739
rect 2944 25707 2976 25739
rect 3016 25707 3048 25739
rect 3088 25707 3120 25739
rect 3160 25707 3192 25739
rect 3232 25707 3264 25739
rect 3304 25707 3336 25739
rect 3376 25707 3408 25739
rect 3448 25707 3480 25739
rect 3520 25707 3552 25739
rect 3592 25707 3624 25739
rect 3664 25707 3696 25739
rect 3736 25707 3768 25739
rect 3808 25707 3840 25739
rect 3880 25707 3912 25739
rect 3952 25707 3984 25739
rect 4024 25707 4056 25739
rect 4096 25707 4128 25739
rect 4168 25707 4200 25739
rect 4240 25707 4272 25739
rect 4312 25707 4344 25739
rect 4384 25707 4416 25739
rect 4456 25707 4488 25739
rect 4528 25707 4560 25739
rect 4600 25707 4632 25739
rect 4672 25707 4704 25739
rect 4744 25707 4776 25739
rect 4816 25707 4848 25739
rect 4888 25707 4920 25739
rect 4960 25707 4992 25739
rect 5032 25707 5064 25739
rect 5104 25707 5136 25739
rect 5176 25707 5208 25739
rect 5248 25707 5280 25739
rect 5320 25707 5352 25739
rect 5392 25707 5424 25739
rect 5464 25707 5496 25739
rect 5536 25707 5568 25739
rect 5608 25707 5640 25739
rect 5680 25707 5712 25739
rect 5752 25707 5784 25739
rect 5824 25707 5856 25739
rect 5896 25707 5928 25739
rect 5968 25707 6000 25739
rect 6040 25707 6072 25739
rect 6112 25707 6144 25739
rect 6184 25707 6216 25739
rect 6256 25707 6288 25739
rect 6328 25707 6360 25739
rect 6400 25707 6432 25739
rect 6472 25707 6504 25739
rect 6544 25707 6576 25739
rect 6616 25707 6648 25739
rect 6688 25707 6720 25739
rect 6760 25707 6792 25739
rect 6832 25707 6864 25739
rect 6904 25707 6936 25739
rect 6976 25707 7008 25739
rect 7048 25707 7080 25739
rect 7120 25707 7152 25739
rect 7192 25707 7224 25739
rect 7264 25707 7296 25739
rect 7336 25707 7368 25739
rect 7408 25707 7440 25739
rect 7480 25707 7512 25739
rect 7552 25707 7584 25739
rect 7624 25707 7656 25739
rect 7696 25707 7728 25739
rect 7768 25707 7800 25739
rect 7840 25707 7872 25739
rect 7912 25707 7944 25739
rect 7984 25707 8016 25739
rect 8056 25707 8088 25739
rect 8128 25707 8160 25739
rect 8200 25707 8232 25739
rect 8272 25707 8304 25739
rect 8344 25707 8376 25739
rect 8416 25707 8448 25739
rect 8488 25707 8520 25739
rect 8560 25707 8592 25739
rect 8632 25707 8664 25739
rect 8704 25707 8736 25739
rect 8776 25707 8808 25739
rect 8848 25707 8880 25739
rect 8920 25707 8952 25739
rect 8992 25707 9024 25739
rect 9064 25707 9096 25739
rect 9136 25707 9168 25739
rect 9208 25707 9240 25739
rect 9280 25707 9312 25739
rect 9352 25707 9384 25739
rect 9424 25707 9456 25739
rect 9496 25707 9528 25739
rect 9568 25707 9600 25739
rect 9640 25707 9672 25739
rect 9712 25707 9744 25739
rect 9784 25707 9816 25739
rect 9856 25707 9888 25739
rect 9928 25707 9960 25739
rect 10000 25707 10032 25739
rect 10072 25707 10104 25739
rect 10144 25707 10176 25739
rect 10216 25707 10248 25739
rect 10288 25707 10320 25739
rect 10360 25707 10392 25739
rect 10432 25707 10464 25739
rect 10504 25707 10536 25739
rect 10576 25707 10608 25739
rect 10648 25707 10680 25739
rect 10720 25707 10752 25739
rect 10792 25707 10824 25739
rect 10864 25707 10896 25739
rect 10936 25707 10968 25739
rect 11008 25707 11040 25739
rect 11080 25707 11112 25739
rect 11152 25707 11184 25739
rect 11224 25707 11256 25739
rect 11296 25707 11328 25739
rect 11368 25707 11400 25739
rect 11440 25707 11472 25739
rect 11512 25707 11544 25739
rect 11584 25707 11616 25739
rect 11656 25707 11688 25739
rect 11728 25707 11760 25739
rect 11800 25707 11832 25739
rect 11872 25707 11904 25739
rect 11944 25707 11976 25739
rect 12016 25707 12048 25739
rect 12088 25707 12120 25739
rect 12160 25707 12192 25739
rect 12232 25707 12264 25739
rect 12304 25707 12336 25739
rect 12376 25707 12408 25739
rect 12448 25707 12480 25739
rect 12520 25707 12552 25739
rect 12592 25707 12624 25739
rect 12664 25707 12696 25739
rect 12736 25707 12768 25739
rect 12808 25707 12840 25739
rect 12880 25707 12912 25739
rect 12952 25707 12984 25739
rect 13024 25707 13056 25739
rect 13096 25707 13128 25739
rect 13168 25707 13200 25739
rect 13240 25707 13272 25739
rect 13312 25707 13344 25739
rect 13384 25707 13416 25739
rect 13456 25707 13488 25739
rect 13528 25707 13560 25739
rect 13600 25707 13632 25739
rect 13672 25707 13704 25739
rect 13744 25707 13776 25739
rect 13816 25707 13848 25739
rect 13888 25707 13920 25739
rect 13960 25707 13992 25739
rect 14032 25707 14064 25739
rect 14104 25707 14136 25739
rect 14176 25707 14208 25739
rect 14248 25707 14280 25739
rect 14320 25707 14352 25739
rect 14392 25707 14424 25739
rect 14464 25707 14496 25739
rect 14536 25707 14568 25739
rect 14608 25707 14640 25739
rect 14680 25707 14712 25739
rect 14752 25707 14784 25739
rect 14824 25707 14856 25739
rect 14896 25707 14928 25739
rect 14968 25707 15000 25739
rect 15040 25707 15072 25739
rect 15112 25707 15144 25739
rect 15184 25707 15216 25739
rect 15256 25707 15288 25739
rect 15328 25707 15360 25739
rect 15400 25707 15432 25739
rect 15472 25707 15504 25739
rect 15544 25707 15576 25739
rect 15616 25707 15648 25739
rect 15688 25707 15720 25739
rect 15760 25707 15792 25739
rect 15832 25707 15864 25739
rect 15904 25707 15936 25739
rect 64 25635 96 25667
rect 136 25635 168 25667
rect 208 25635 240 25667
rect 280 25635 312 25667
rect 352 25635 384 25667
rect 424 25635 456 25667
rect 496 25635 528 25667
rect 568 25635 600 25667
rect 640 25635 672 25667
rect 712 25635 744 25667
rect 784 25635 816 25667
rect 856 25635 888 25667
rect 928 25635 960 25667
rect 1000 25635 1032 25667
rect 1072 25635 1104 25667
rect 1144 25635 1176 25667
rect 1216 25635 1248 25667
rect 1288 25635 1320 25667
rect 1360 25635 1392 25667
rect 1432 25635 1464 25667
rect 1504 25635 1536 25667
rect 1576 25635 1608 25667
rect 1648 25635 1680 25667
rect 1720 25635 1752 25667
rect 1792 25635 1824 25667
rect 1864 25635 1896 25667
rect 1936 25635 1968 25667
rect 2008 25635 2040 25667
rect 2080 25635 2112 25667
rect 2152 25635 2184 25667
rect 2224 25635 2256 25667
rect 2296 25635 2328 25667
rect 2368 25635 2400 25667
rect 2440 25635 2472 25667
rect 2512 25635 2544 25667
rect 2584 25635 2616 25667
rect 2656 25635 2688 25667
rect 2728 25635 2760 25667
rect 2800 25635 2832 25667
rect 2872 25635 2904 25667
rect 2944 25635 2976 25667
rect 3016 25635 3048 25667
rect 3088 25635 3120 25667
rect 3160 25635 3192 25667
rect 3232 25635 3264 25667
rect 3304 25635 3336 25667
rect 3376 25635 3408 25667
rect 3448 25635 3480 25667
rect 3520 25635 3552 25667
rect 3592 25635 3624 25667
rect 3664 25635 3696 25667
rect 3736 25635 3768 25667
rect 3808 25635 3840 25667
rect 3880 25635 3912 25667
rect 3952 25635 3984 25667
rect 4024 25635 4056 25667
rect 4096 25635 4128 25667
rect 4168 25635 4200 25667
rect 4240 25635 4272 25667
rect 4312 25635 4344 25667
rect 4384 25635 4416 25667
rect 4456 25635 4488 25667
rect 4528 25635 4560 25667
rect 4600 25635 4632 25667
rect 4672 25635 4704 25667
rect 4744 25635 4776 25667
rect 4816 25635 4848 25667
rect 4888 25635 4920 25667
rect 4960 25635 4992 25667
rect 5032 25635 5064 25667
rect 5104 25635 5136 25667
rect 5176 25635 5208 25667
rect 5248 25635 5280 25667
rect 5320 25635 5352 25667
rect 5392 25635 5424 25667
rect 5464 25635 5496 25667
rect 5536 25635 5568 25667
rect 5608 25635 5640 25667
rect 5680 25635 5712 25667
rect 5752 25635 5784 25667
rect 5824 25635 5856 25667
rect 5896 25635 5928 25667
rect 5968 25635 6000 25667
rect 6040 25635 6072 25667
rect 6112 25635 6144 25667
rect 6184 25635 6216 25667
rect 6256 25635 6288 25667
rect 6328 25635 6360 25667
rect 6400 25635 6432 25667
rect 6472 25635 6504 25667
rect 6544 25635 6576 25667
rect 6616 25635 6648 25667
rect 6688 25635 6720 25667
rect 6760 25635 6792 25667
rect 6832 25635 6864 25667
rect 6904 25635 6936 25667
rect 6976 25635 7008 25667
rect 7048 25635 7080 25667
rect 7120 25635 7152 25667
rect 7192 25635 7224 25667
rect 7264 25635 7296 25667
rect 7336 25635 7368 25667
rect 7408 25635 7440 25667
rect 7480 25635 7512 25667
rect 7552 25635 7584 25667
rect 7624 25635 7656 25667
rect 7696 25635 7728 25667
rect 7768 25635 7800 25667
rect 7840 25635 7872 25667
rect 7912 25635 7944 25667
rect 7984 25635 8016 25667
rect 8056 25635 8088 25667
rect 8128 25635 8160 25667
rect 8200 25635 8232 25667
rect 8272 25635 8304 25667
rect 8344 25635 8376 25667
rect 8416 25635 8448 25667
rect 8488 25635 8520 25667
rect 8560 25635 8592 25667
rect 8632 25635 8664 25667
rect 8704 25635 8736 25667
rect 8776 25635 8808 25667
rect 8848 25635 8880 25667
rect 8920 25635 8952 25667
rect 8992 25635 9024 25667
rect 9064 25635 9096 25667
rect 9136 25635 9168 25667
rect 9208 25635 9240 25667
rect 9280 25635 9312 25667
rect 9352 25635 9384 25667
rect 9424 25635 9456 25667
rect 9496 25635 9528 25667
rect 9568 25635 9600 25667
rect 9640 25635 9672 25667
rect 9712 25635 9744 25667
rect 9784 25635 9816 25667
rect 9856 25635 9888 25667
rect 9928 25635 9960 25667
rect 10000 25635 10032 25667
rect 10072 25635 10104 25667
rect 10144 25635 10176 25667
rect 10216 25635 10248 25667
rect 10288 25635 10320 25667
rect 10360 25635 10392 25667
rect 10432 25635 10464 25667
rect 10504 25635 10536 25667
rect 10576 25635 10608 25667
rect 10648 25635 10680 25667
rect 10720 25635 10752 25667
rect 10792 25635 10824 25667
rect 10864 25635 10896 25667
rect 10936 25635 10968 25667
rect 11008 25635 11040 25667
rect 11080 25635 11112 25667
rect 11152 25635 11184 25667
rect 11224 25635 11256 25667
rect 11296 25635 11328 25667
rect 11368 25635 11400 25667
rect 11440 25635 11472 25667
rect 11512 25635 11544 25667
rect 11584 25635 11616 25667
rect 11656 25635 11688 25667
rect 11728 25635 11760 25667
rect 11800 25635 11832 25667
rect 11872 25635 11904 25667
rect 11944 25635 11976 25667
rect 12016 25635 12048 25667
rect 12088 25635 12120 25667
rect 12160 25635 12192 25667
rect 12232 25635 12264 25667
rect 12304 25635 12336 25667
rect 12376 25635 12408 25667
rect 12448 25635 12480 25667
rect 12520 25635 12552 25667
rect 12592 25635 12624 25667
rect 12664 25635 12696 25667
rect 12736 25635 12768 25667
rect 12808 25635 12840 25667
rect 12880 25635 12912 25667
rect 12952 25635 12984 25667
rect 13024 25635 13056 25667
rect 13096 25635 13128 25667
rect 13168 25635 13200 25667
rect 13240 25635 13272 25667
rect 13312 25635 13344 25667
rect 13384 25635 13416 25667
rect 13456 25635 13488 25667
rect 13528 25635 13560 25667
rect 13600 25635 13632 25667
rect 13672 25635 13704 25667
rect 13744 25635 13776 25667
rect 13816 25635 13848 25667
rect 13888 25635 13920 25667
rect 13960 25635 13992 25667
rect 14032 25635 14064 25667
rect 14104 25635 14136 25667
rect 14176 25635 14208 25667
rect 14248 25635 14280 25667
rect 14320 25635 14352 25667
rect 14392 25635 14424 25667
rect 14464 25635 14496 25667
rect 14536 25635 14568 25667
rect 14608 25635 14640 25667
rect 14680 25635 14712 25667
rect 14752 25635 14784 25667
rect 14824 25635 14856 25667
rect 14896 25635 14928 25667
rect 14968 25635 15000 25667
rect 15040 25635 15072 25667
rect 15112 25635 15144 25667
rect 15184 25635 15216 25667
rect 15256 25635 15288 25667
rect 15328 25635 15360 25667
rect 15400 25635 15432 25667
rect 15472 25635 15504 25667
rect 15544 25635 15576 25667
rect 15616 25635 15648 25667
rect 15688 25635 15720 25667
rect 15760 25635 15792 25667
rect 15832 25635 15864 25667
rect 15904 25635 15936 25667
rect 64 25563 96 25595
rect 136 25563 168 25595
rect 208 25563 240 25595
rect 280 25563 312 25595
rect 352 25563 384 25595
rect 424 25563 456 25595
rect 496 25563 528 25595
rect 568 25563 600 25595
rect 640 25563 672 25595
rect 712 25563 744 25595
rect 784 25563 816 25595
rect 856 25563 888 25595
rect 928 25563 960 25595
rect 1000 25563 1032 25595
rect 1072 25563 1104 25595
rect 1144 25563 1176 25595
rect 1216 25563 1248 25595
rect 1288 25563 1320 25595
rect 1360 25563 1392 25595
rect 1432 25563 1464 25595
rect 1504 25563 1536 25595
rect 1576 25563 1608 25595
rect 1648 25563 1680 25595
rect 1720 25563 1752 25595
rect 1792 25563 1824 25595
rect 1864 25563 1896 25595
rect 1936 25563 1968 25595
rect 2008 25563 2040 25595
rect 2080 25563 2112 25595
rect 2152 25563 2184 25595
rect 2224 25563 2256 25595
rect 2296 25563 2328 25595
rect 2368 25563 2400 25595
rect 2440 25563 2472 25595
rect 2512 25563 2544 25595
rect 2584 25563 2616 25595
rect 2656 25563 2688 25595
rect 2728 25563 2760 25595
rect 2800 25563 2832 25595
rect 2872 25563 2904 25595
rect 2944 25563 2976 25595
rect 3016 25563 3048 25595
rect 3088 25563 3120 25595
rect 3160 25563 3192 25595
rect 3232 25563 3264 25595
rect 3304 25563 3336 25595
rect 3376 25563 3408 25595
rect 3448 25563 3480 25595
rect 3520 25563 3552 25595
rect 3592 25563 3624 25595
rect 3664 25563 3696 25595
rect 3736 25563 3768 25595
rect 3808 25563 3840 25595
rect 3880 25563 3912 25595
rect 3952 25563 3984 25595
rect 4024 25563 4056 25595
rect 4096 25563 4128 25595
rect 4168 25563 4200 25595
rect 4240 25563 4272 25595
rect 4312 25563 4344 25595
rect 4384 25563 4416 25595
rect 4456 25563 4488 25595
rect 4528 25563 4560 25595
rect 4600 25563 4632 25595
rect 4672 25563 4704 25595
rect 4744 25563 4776 25595
rect 4816 25563 4848 25595
rect 4888 25563 4920 25595
rect 4960 25563 4992 25595
rect 5032 25563 5064 25595
rect 5104 25563 5136 25595
rect 5176 25563 5208 25595
rect 5248 25563 5280 25595
rect 5320 25563 5352 25595
rect 5392 25563 5424 25595
rect 5464 25563 5496 25595
rect 5536 25563 5568 25595
rect 5608 25563 5640 25595
rect 5680 25563 5712 25595
rect 5752 25563 5784 25595
rect 5824 25563 5856 25595
rect 5896 25563 5928 25595
rect 5968 25563 6000 25595
rect 6040 25563 6072 25595
rect 6112 25563 6144 25595
rect 6184 25563 6216 25595
rect 6256 25563 6288 25595
rect 6328 25563 6360 25595
rect 6400 25563 6432 25595
rect 6472 25563 6504 25595
rect 6544 25563 6576 25595
rect 6616 25563 6648 25595
rect 6688 25563 6720 25595
rect 6760 25563 6792 25595
rect 6832 25563 6864 25595
rect 6904 25563 6936 25595
rect 6976 25563 7008 25595
rect 7048 25563 7080 25595
rect 7120 25563 7152 25595
rect 7192 25563 7224 25595
rect 7264 25563 7296 25595
rect 7336 25563 7368 25595
rect 7408 25563 7440 25595
rect 7480 25563 7512 25595
rect 7552 25563 7584 25595
rect 7624 25563 7656 25595
rect 7696 25563 7728 25595
rect 7768 25563 7800 25595
rect 7840 25563 7872 25595
rect 7912 25563 7944 25595
rect 7984 25563 8016 25595
rect 8056 25563 8088 25595
rect 8128 25563 8160 25595
rect 8200 25563 8232 25595
rect 8272 25563 8304 25595
rect 8344 25563 8376 25595
rect 8416 25563 8448 25595
rect 8488 25563 8520 25595
rect 8560 25563 8592 25595
rect 8632 25563 8664 25595
rect 8704 25563 8736 25595
rect 8776 25563 8808 25595
rect 8848 25563 8880 25595
rect 8920 25563 8952 25595
rect 8992 25563 9024 25595
rect 9064 25563 9096 25595
rect 9136 25563 9168 25595
rect 9208 25563 9240 25595
rect 9280 25563 9312 25595
rect 9352 25563 9384 25595
rect 9424 25563 9456 25595
rect 9496 25563 9528 25595
rect 9568 25563 9600 25595
rect 9640 25563 9672 25595
rect 9712 25563 9744 25595
rect 9784 25563 9816 25595
rect 9856 25563 9888 25595
rect 9928 25563 9960 25595
rect 10000 25563 10032 25595
rect 10072 25563 10104 25595
rect 10144 25563 10176 25595
rect 10216 25563 10248 25595
rect 10288 25563 10320 25595
rect 10360 25563 10392 25595
rect 10432 25563 10464 25595
rect 10504 25563 10536 25595
rect 10576 25563 10608 25595
rect 10648 25563 10680 25595
rect 10720 25563 10752 25595
rect 10792 25563 10824 25595
rect 10864 25563 10896 25595
rect 10936 25563 10968 25595
rect 11008 25563 11040 25595
rect 11080 25563 11112 25595
rect 11152 25563 11184 25595
rect 11224 25563 11256 25595
rect 11296 25563 11328 25595
rect 11368 25563 11400 25595
rect 11440 25563 11472 25595
rect 11512 25563 11544 25595
rect 11584 25563 11616 25595
rect 11656 25563 11688 25595
rect 11728 25563 11760 25595
rect 11800 25563 11832 25595
rect 11872 25563 11904 25595
rect 11944 25563 11976 25595
rect 12016 25563 12048 25595
rect 12088 25563 12120 25595
rect 12160 25563 12192 25595
rect 12232 25563 12264 25595
rect 12304 25563 12336 25595
rect 12376 25563 12408 25595
rect 12448 25563 12480 25595
rect 12520 25563 12552 25595
rect 12592 25563 12624 25595
rect 12664 25563 12696 25595
rect 12736 25563 12768 25595
rect 12808 25563 12840 25595
rect 12880 25563 12912 25595
rect 12952 25563 12984 25595
rect 13024 25563 13056 25595
rect 13096 25563 13128 25595
rect 13168 25563 13200 25595
rect 13240 25563 13272 25595
rect 13312 25563 13344 25595
rect 13384 25563 13416 25595
rect 13456 25563 13488 25595
rect 13528 25563 13560 25595
rect 13600 25563 13632 25595
rect 13672 25563 13704 25595
rect 13744 25563 13776 25595
rect 13816 25563 13848 25595
rect 13888 25563 13920 25595
rect 13960 25563 13992 25595
rect 14032 25563 14064 25595
rect 14104 25563 14136 25595
rect 14176 25563 14208 25595
rect 14248 25563 14280 25595
rect 14320 25563 14352 25595
rect 14392 25563 14424 25595
rect 14464 25563 14496 25595
rect 14536 25563 14568 25595
rect 14608 25563 14640 25595
rect 14680 25563 14712 25595
rect 14752 25563 14784 25595
rect 14824 25563 14856 25595
rect 14896 25563 14928 25595
rect 14968 25563 15000 25595
rect 15040 25563 15072 25595
rect 15112 25563 15144 25595
rect 15184 25563 15216 25595
rect 15256 25563 15288 25595
rect 15328 25563 15360 25595
rect 15400 25563 15432 25595
rect 15472 25563 15504 25595
rect 15544 25563 15576 25595
rect 15616 25563 15648 25595
rect 15688 25563 15720 25595
rect 15760 25563 15792 25595
rect 15832 25563 15864 25595
rect 15904 25563 15936 25595
rect 64 25491 96 25523
rect 136 25491 168 25523
rect 208 25491 240 25523
rect 280 25491 312 25523
rect 352 25491 384 25523
rect 424 25491 456 25523
rect 496 25491 528 25523
rect 568 25491 600 25523
rect 640 25491 672 25523
rect 712 25491 744 25523
rect 784 25491 816 25523
rect 856 25491 888 25523
rect 928 25491 960 25523
rect 1000 25491 1032 25523
rect 1072 25491 1104 25523
rect 1144 25491 1176 25523
rect 1216 25491 1248 25523
rect 1288 25491 1320 25523
rect 1360 25491 1392 25523
rect 1432 25491 1464 25523
rect 1504 25491 1536 25523
rect 1576 25491 1608 25523
rect 1648 25491 1680 25523
rect 1720 25491 1752 25523
rect 1792 25491 1824 25523
rect 1864 25491 1896 25523
rect 1936 25491 1968 25523
rect 2008 25491 2040 25523
rect 2080 25491 2112 25523
rect 2152 25491 2184 25523
rect 2224 25491 2256 25523
rect 2296 25491 2328 25523
rect 2368 25491 2400 25523
rect 2440 25491 2472 25523
rect 2512 25491 2544 25523
rect 2584 25491 2616 25523
rect 2656 25491 2688 25523
rect 2728 25491 2760 25523
rect 2800 25491 2832 25523
rect 2872 25491 2904 25523
rect 2944 25491 2976 25523
rect 3016 25491 3048 25523
rect 3088 25491 3120 25523
rect 3160 25491 3192 25523
rect 3232 25491 3264 25523
rect 3304 25491 3336 25523
rect 3376 25491 3408 25523
rect 3448 25491 3480 25523
rect 3520 25491 3552 25523
rect 3592 25491 3624 25523
rect 3664 25491 3696 25523
rect 3736 25491 3768 25523
rect 3808 25491 3840 25523
rect 3880 25491 3912 25523
rect 3952 25491 3984 25523
rect 4024 25491 4056 25523
rect 4096 25491 4128 25523
rect 4168 25491 4200 25523
rect 4240 25491 4272 25523
rect 4312 25491 4344 25523
rect 4384 25491 4416 25523
rect 4456 25491 4488 25523
rect 4528 25491 4560 25523
rect 4600 25491 4632 25523
rect 4672 25491 4704 25523
rect 4744 25491 4776 25523
rect 4816 25491 4848 25523
rect 4888 25491 4920 25523
rect 4960 25491 4992 25523
rect 5032 25491 5064 25523
rect 5104 25491 5136 25523
rect 5176 25491 5208 25523
rect 5248 25491 5280 25523
rect 5320 25491 5352 25523
rect 5392 25491 5424 25523
rect 5464 25491 5496 25523
rect 5536 25491 5568 25523
rect 5608 25491 5640 25523
rect 5680 25491 5712 25523
rect 5752 25491 5784 25523
rect 5824 25491 5856 25523
rect 5896 25491 5928 25523
rect 5968 25491 6000 25523
rect 6040 25491 6072 25523
rect 6112 25491 6144 25523
rect 6184 25491 6216 25523
rect 6256 25491 6288 25523
rect 6328 25491 6360 25523
rect 6400 25491 6432 25523
rect 6472 25491 6504 25523
rect 6544 25491 6576 25523
rect 6616 25491 6648 25523
rect 6688 25491 6720 25523
rect 6760 25491 6792 25523
rect 6832 25491 6864 25523
rect 6904 25491 6936 25523
rect 6976 25491 7008 25523
rect 7048 25491 7080 25523
rect 7120 25491 7152 25523
rect 7192 25491 7224 25523
rect 7264 25491 7296 25523
rect 7336 25491 7368 25523
rect 7408 25491 7440 25523
rect 7480 25491 7512 25523
rect 7552 25491 7584 25523
rect 7624 25491 7656 25523
rect 7696 25491 7728 25523
rect 7768 25491 7800 25523
rect 7840 25491 7872 25523
rect 7912 25491 7944 25523
rect 7984 25491 8016 25523
rect 8056 25491 8088 25523
rect 8128 25491 8160 25523
rect 8200 25491 8232 25523
rect 8272 25491 8304 25523
rect 8344 25491 8376 25523
rect 8416 25491 8448 25523
rect 8488 25491 8520 25523
rect 8560 25491 8592 25523
rect 8632 25491 8664 25523
rect 8704 25491 8736 25523
rect 8776 25491 8808 25523
rect 8848 25491 8880 25523
rect 8920 25491 8952 25523
rect 8992 25491 9024 25523
rect 9064 25491 9096 25523
rect 9136 25491 9168 25523
rect 9208 25491 9240 25523
rect 9280 25491 9312 25523
rect 9352 25491 9384 25523
rect 9424 25491 9456 25523
rect 9496 25491 9528 25523
rect 9568 25491 9600 25523
rect 9640 25491 9672 25523
rect 9712 25491 9744 25523
rect 9784 25491 9816 25523
rect 9856 25491 9888 25523
rect 9928 25491 9960 25523
rect 10000 25491 10032 25523
rect 10072 25491 10104 25523
rect 10144 25491 10176 25523
rect 10216 25491 10248 25523
rect 10288 25491 10320 25523
rect 10360 25491 10392 25523
rect 10432 25491 10464 25523
rect 10504 25491 10536 25523
rect 10576 25491 10608 25523
rect 10648 25491 10680 25523
rect 10720 25491 10752 25523
rect 10792 25491 10824 25523
rect 10864 25491 10896 25523
rect 10936 25491 10968 25523
rect 11008 25491 11040 25523
rect 11080 25491 11112 25523
rect 11152 25491 11184 25523
rect 11224 25491 11256 25523
rect 11296 25491 11328 25523
rect 11368 25491 11400 25523
rect 11440 25491 11472 25523
rect 11512 25491 11544 25523
rect 11584 25491 11616 25523
rect 11656 25491 11688 25523
rect 11728 25491 11760 25523
rect 11800 25491 11832 25523
rect 11872 25491 11904 25523
rect 11944 25491 11976 25523
rect 12016 25491 12048 25523
rect 12088 25491 12120 25523
rect 12160 25491 12192 25523
rect 12232 25491 12264 25523
rect 12304 25491 12336 25523
rect 12376 25491 12408 25523
rect 12448 25491 12480 25523
rect 12520 25491 12552 25523
rect 12592 25491 12624 25523
rect 12664 25491 12696 25523
rect 12736 25491 12768 25523
rect 12808 25491 12840 25523
rect 12880 25491 12912 25523
rect 12952 25491 12984 25523
rect 13024 25491 13056 25523
rect 13096 25491 13128 25523
rect 13168 25491 13200 25523
rect 13240 25491 13272 25523
rect 13312 25491 13344 25523
rect 13384 25491 13416 25523
rect 13456 25491 13488 25523
rect 13528 25491 13560 25523
rect 13600 25491 13632 25523
rect 13672 25491 13704 25523
rect 13744 25491 13776 25523
rect 13816 25491 13848 25523
rect 13888 25491 13920 25523
rect 13960 25491 13992 25523
rect 14032 25491 14064 25523
rect 14104 25491 14136 25523
rect 14176 25491 14208 25523
rect 14248 25491 14280 25523
rect 14320 25491 14352 25523
rect 14392 25491 14424 25523
rect 14464 25491 14496 25523
rect 14536 25491 14568 25523
rect 14608 25491 14640 25523
rect 14680 25491 14712 25523
rect 14752 25491 14784 25523
rect 14824 25491 14856 25523
rect 14896 25491 14928 25523
rect 14968 25491 15000 25523
rect 15040 25491 15072 25523
rect 15112 25491 15144 25523
rect 15184 25491 15216 25523
rect 15256 25491 15288 25523
rect 15328 25491 15360 25523
rect 15400 25491 15432 25523
rect 15472 25491 15504 25523
rect 15544 25491 15576 25523
rect 15616 25491 15648 25523
rect 15688 25491 15720 25523
rect 15760 25491 15792 25523
rect 15832 25491 15864 25523
rect 15904 25491 15936 25523
rect 64 25419 96 25451
rect 136 25419 168 25451
rect 208 25419 240 25451
rect 280 25419 312 25451
rect 352 25419 384 25451
rect 424 25419 456 25451
rect 496 25419 528 25451
rect 568 25419 600 25451
rect 640 25419 672 25451
rect 712 25419 744 25451
rect 784 25419 816 25451
rect 856 25419 888 25451
rect 928 25419 960 25451
rect 1000 25419 1032 25451
rect 1072 25419 1104 25451
rect 1144 25419 1176 25451
rect 1216 25419 1248 25451
rect 1288 25419 1320 25451
rect 1360 25419 1392 25451
rect 1432 25419 1464 25451
rect 1504 25419 1536 25451
rect 1576 25419 1608 25451
rect 1648 25419 1680 25451
rect 1720 25419 1752 25451
rect 1792 25419 1824 25451
rect 1864 25419 1896 25451
rect 1936 25419 1968 25451
rect 2008 25419 2040 25451
rect 2080 25419 2112 25451
rect 2152 25419 2184 25451
rect 2224 25419 2256 25451
rect 2296 25419 2328 25451
rect 2368 25419 2400 25451
rect 2440 25419 2472 25451
rect 2512 25419 2544 25451
rect 2584 25419 2616 25451
rect 2656 25419 2688 25451
rect 2728 25419 2760 25451
rect 2800 25419 2832 25451
rect 2872 25419 2904 25451
rect 2944 25419 2976 25451
rect 3016 25419 3048 25451
rect 3088 25419 3120 25451
rect 3160 25419 3192 25451
rect 3232 25419 3264 25451
rect 3304 25419 3336 25451
rect 3376 25419 3408 25451
rect 3448 25419 3480 25451
rect 3520 25419 3552 25451
rect 3592 25419 3624 25451
rect 3664 25419 3696 25451
rect 3736 25419 3768 25451
rect 3808 25419 3840 25451
rect 3880 25419 3912 25451
rect 3952 25419 3984 25451
rect 4024 25419 4056 25451
rect 4096 25419 4128 25451
rect 4168 25419 4200 25451
rect 4240 25419 4272 25451
rect 4312 25419 4344 25451
rect 4384 25419 4416 25451
rect 4456 25419 4488 25451
rect 4528 25419 4560 25451
rect 4600 25419 4632 25451
rect 4672 25419 4704 25451
rect 4744 25419 4776 25451
rect 4816 25419 4848 25451
rect 4888 25419 4920 25451
rect 4960 25419 4992 25451
rect 5032 25419 5064 25451
rect 5104 25419 5136 25451
rect 5176 25419 5208 25451
rect 5248 25419 5280 25451
rect 5320 25419 5352 25451
rect 5392 25419 5424 25451
rect 5464 25419 5496 25451
rect 5536 25419 5568 25451
rect 5608 25419 5640 25451
rect 5680 25419 5712 25451
rect 5752 25419 5784 25451
rect 5824 25419 5856 25451
rect 5896 25419 5928 25451
rect 5968 25419 6000 25451
rect 6040 25419 6072 25451
rect 6112 25419 6144 25451
rect 6184 25419 6216 25451
rect 6256 25419 6288 25451
rect 6328 25419 6360 25451
rect 6400 25419 6432 25451
rect 6472 25419 6504 25451
rect 6544 25419 6576 25451
rect 6616 25419 6648 25451
rect 6688 25419 6720 25451
rect 6760 25419 6792 25451
rect 6832 25419 6864 25451
rect 6904 25419 6936 25451
rect 6976 25419 7008 25451
rect 7048 25419 7080 25451
rect 7120 25419 7152 25451
rect 7192 25419 7224 25451
rect 7264 25419 7296 25451
rect 7336 25419 7368 25451
rect 7408 25419 7440 25451
rect 7480 25419 7512 25451
rect 7552 25419 7584 25451
rect 7624 25419 7656 25451
rect 7696 25419 7728 25451
rect 7768 25419 7800 25451
rect 7840 25419 7872 25451
rect 7912 25419 7944 25451
rect 7984 25419 8016 25451
rect 8056 25419 8088 25451
rect 8128 25419 8160 25451
rect 8200 25419 8232 25451
rect 8272 25419 8304 25451
rect 8344 25419 8376 25451
rect 8416 25419 8448 25451
rect 8488 25419 8520 25451
rect 8560 25419 8592 25451
rect 8632 25419 8664 25451
rect 8704 25419 8736 25451
rect 8776 25419 8808 25451
rect 8848 25419 8880 25451
rect 8920 25419 8952 25451
rect 8992 25419 9024 25451
rect 9064 25419 9096 25451
rect 9136 25419 9168 25451
rect 9208 25419 9240 25451
rect 9280 25419 9312 25451
rect 9352 25419 9384 25451
rect 9424 25419 9456 25451
rect 9496 25419 9528 25451
rect 9568 25419 9600 25451
rect 9640 25419 9672 25451
rect 9712 25419 9744 25451
rect 9784 25419 9816 25451
rect 9856 25419 9888 25451
rect 9928 25419 9960 25451
rect 10000 25419 10032 25451
rect 10072 25419 10104 25451
rect 10144 25419 10176 25451
rect 10216 25419 10248 25451
rect 10288 25419 10320 25451
rect 10360 25419 10392 25451
rect 10432 25419 10464 25451
rect 10504 25419 10536 25451
rect 10576 25419 10608 25451
rect 10648 25419 10680 25451
rect 10720 25419 10752 25451
rect 10792 25419 10824 25451
rect 10864 25419 10896 25451
rect 10936 25419 10968 25451
rect 11008 25419 11040 25451
rect 11080 25419 11112 25451
rect 11152 25419 11184 25451
rect 11224 25419 11256 25451
rect 11296 25419 11328 25451
rect 11368 25419 11400 25451
rect 11440 25419 11472 25451
rect 11512 25419 11544 25451
rect 11584 25419 11616 25451
rect 11656 25419 11688 25451
rect 11728 25419 11760 25451
rect 11800 25419 11832 25451
rect 11872 25419 11904 25451
rect 11944 25419 11976 25451
rect 12016 25419 12048 25451
rect 12088 25419 12120 25451
rect 12160 25419 12192 25451
rect 12232 25419 12264 25451
rect 12304 25419 12336 25451
rect 12376 25419 12408 25451
rect 12448 25419 12480 25451
rect 12520 25419 12552 25451
rect 12592 25419 12624 25451
rect 12664 25419 12696 25451
rect 12736 25419 12768 25451
rect 12808 25419 12840 25451
rect 12880 25419 12912 25451
rect 12952 25419 12984 25451
rect 13024 25419 13056 25451
rect 13096 25419 13128 25451
rect 13168 25419 13200 25451
rect 13240 25419 13272 25451
rect 13312 25419 13344 25451
rect 13384 25419 13416 25451
rect 13456 25419 13488 25451
rect 13528 25419 13560 25451
rect 13600 25419 13632 25451
rect 13672 25419 13704 25451
rect 13744 25419 13776 25451
rect 13816 25419 13848 25451
rect 13888 25419 13920 25451
rect 13960 25419 13992 25451
rect 14032 25419 14064 25451
rect 14104 25419 14136 25451
rect 14176 25419 14208 25451
rect 14248 25419 14280 25451
rect 14320 25419 14352 25451
rect 14392 25419 14424 25451
rect 14464 25419 14496 25451
rect 14536 25419 14568 25451
rect 14608 25419 14640 25451
rect 14680 25419 14712 25451
rect 14752 25419 14784 25451
rect 14824 25419 14856 25451
rect 14896 25419 14928 25451
rect 14968 25419 15000 25451
rect 15040 25419 15072 25451
rect 15112 25419 15144 25451
rect 15184 25419 15216 25451
rect 15256 25419 15288 25451
rect 15328 25419 15360 25451
rect 15400 25419 15432 25451
rect 15472 25419 15504 25451
rect 15544 25419 15576 25451
rect 15616 25419 15648 25451
rect 15688 25419 15720 25451
rect 15760 25419 15792 25451
rect 15832 25419 15864 25451
rect 15904 25419 15936 25451
rect 64 25347 96 25379
rect 136 25347 168 25379
rect 208 25347 240 25379
rect 280 25347 312 25379
rect 352 25347 384 25379
rect 424 25347 456 25379
rect 496 25347 528 25379
rect 568 25347 600 25379
rect 640 25347 672 25379
rect 712 25347 744 25379
rect 784 25347 816 25379
rect 856 25347 888 25379
rect 928 25347 960 25379
rect 1000 25347 1032 25379
rect 1072 25347 1104 25379
rect 1144 25347 1176 25379
rect 1216 25347 1248 25379
rect 1288 25347 1320 25379
rect 1360 25347 1392 25379
rect 1432 25347 1464 25379
rect 1504 25347 1536 25379
rect 1576 25347 1608 25379
rect 1648 25347 1680 25379
rect 1720 25347 1752 25379
rect 1792 25347 1824 25379
rect 1864 25347 1896 25379
rect 1936 25347 1968 25379
rect 2008 25347 2040 25379
rect 2080 25347 2112 25379
rect 2152 25347 2184 25379
rect 2224 25347 2256 25379
rect 2296 25347 2328 25379
rect 2368 25347 2400 25379
rect 2440 25347 2472 25379
rect 2512 25347 2544 25379
rect 2584 25347 2616 25379
rect 2656 25347 2688 25379
rect 2728 25347 2760 25379
rect 2800 25347 2832 25379
rect 2872 25347 2904 25379
rect 2944 25347 2976 25379
rect 3016 25347 3048 25379
rect 3088 25347 3120 25379
rect 3160 25347 3192 25379
rect 3232 25347 3264 25379
rect 3304 25347 3336 25379
rect 3376 25347 3408 25379
rect 3448 25347 3480 25379
rect 3520 25347 3552 25379
rect 3592 25347 3624 25379
rect 3664 25347 3696 25379
rect 3736 25347 3768 25379
rect 3808 25347 3840 25379
rect 3880 25347 3912 25379
rect 3952 25347 3984 25379
rect 4024 25347 4056 25379
rect 4096 25347 4128 25379
rect 4168 25347 4200 25379
rect 4240 25347 4272 25379
rect 4312 25347 4344 25379
rect 4384 25347 4416 25379
rect 4456 25347 4488 25379
rect 4528 25347 4560 25379
rect 4600 25347 4632 25379
rect 4672 25347 4704 25379
rect 4744 25347 4776 25379
rect 4816 25347 4848 25379
rect 4888 25347 4920 25379
rect 4960 25347 4992 25379
rect 5032 25347 5064 25379
rect 5104 25347 5136 25379
rect 5176 25347 5208 25379
rect 5248 25347 5280 25379
rect 5320 25347 5352 25379
rect 5392 25347 5424 25379
rect 5464 25347 5496 25379
rect 5536 25347 5568 25379
rect 5608 25347 5640 25379
rect 5680 25347 5712 25379
rect 5752 25347 5784 25379
rect 5824 25347 5856 25379
rect 5896 25347 5928 25379
rect 5968 25347 6000 25379
rect 6040 25347 6072 25379
rect 6112 25347 6144 25379
rect 6184 25347 6216 25379
rect 6256 25347 6288 25379
rect 6328 25347 6360 25379
rect 6400 25347 6432 25379
rect 6472 25347 6504 25379
rect 6544 25347 6576 25379
rect 6616 25347 6648 25379
rect 6688 25347 6720 25379
rect 6760 25347 6792 25379
rect 6832 25347 6864 25379
rect 6904 25347 6936 25379
rect 6976 25347 7008 25379
rect 7048 25347 7080 25379
rect 7120 25347 7152 25379
rect 7192 25347 7224 25379
rect 7264 25347 7296 25379
rect 7336 25347 7368 25379
rect 7408 25347 7440 25379
rect 7480 25347 7512 25379
rect 7552 25347 7584 25379
rect 7624 25347 7656 25379
rect 7696 25347 7728 25379
rect 7768 25347 7800 25379
rect 7840 25347 7872 25379
rect 7912 25347 7944 25379
rect 7984 25347 8016 25379
rect 8056 25347 8088 25379
rect 8128 25347 8160 25379
rect 8200 25347 8232 25379
rect 8272 25347 8304 25379
rect 8344 25347 8376 25379
rect 8416 25347 8448 25379
rect 8488 25347 8520 25379
rect 8560 25347 8592 25379
rect 8632 25347 8664 25379
rect 8704 25347 8736 25379
rect 8776 25347 8808 25379
rect 8848 25347 8880 25379
rect 8920 25347 8952 25379
rect 8992 25347 9024 25379
rect 9064 25347 9096 25379
rect 9136 25347 9168 25379
rect 9208 25347 9240 25379
rect 9280 25347 9312 25379
rect 9352 25347 9384 25379
rect 9424 25347 9456 25379
rect 9496 25347 9528 25379
rect 9568 25347 9600 25379
rect 9640 25347 9672 25379
rect 9712 25347 9744 25379
rect 9784 25347 9816 25379
rect 9856 25347 9888 25379
rect 9928 25347 9960 25379
rect 10000 25347 10032 25379
rect 10072 25347 10104 25379
rect 10144 25347 10176 25379
rect 10216 25347 10248 25379
rect 10288 25347 10320 25379
rect 10360 25347 10392 25379
rect 10432 25347 10464 25379
rect 10504 25347 10536 25379
rect 10576 25347 10608 25379
rect 10648 25347 10680 25379
rect 10720 25347 10752 25379
rect 10792 25347 10824 25379
rect 10864 25347 10896 25379
rect 10936 25347 10968 25379
rect 11008 25347 11040 25379
rect 11080 25347 11112 25379
rect 11152 25347 11184 25379
rect 11224 25347 11256 25379
rect 11296 25347 11328 25379
rect 11368 25347 11400 25379
rect 11440 25347 11472 25379
rect 11512 25347 11544 25379
rect 11584 25347 11616 25379
rect 11656 25347 11688 25379
rect 11728 25347 11760 25379
rect 11800 25347 11832 25379
rect 11872 25347 11904 25379
rect 11944 25347 11976 25379
rect 12016 25347 12048 25379
rect 12088 25347 12120 25379
rect 12160 25347 12192 25379
rect 12232 25347 12264 25379
rect 12304 25347 12336 25379
rect 12376 25347 12408 25379
rect 12448 25347 12480 25379
rect 12520 25347 12552 25379
rect 12592 25347 12624 25379
rect 12664 25347 12696 25379
rect 12736 25347 12768 25379
rect 12808 25347 12840 25379
rect 12880 25347 12912 25379
rect 12952 25347 12984 25379
rect 13024 25347 13056 25379
rect 13096 25347 13128 25379
rect 13168 25347 13200 25379
rect 13240 25347 13272 25379
rect 13312 25347 13344 25379
rect 13384 25347 13416 25379
rect 13456 25347 13488 25379
rect 13528 25347 13560 25379
rect 13600 25347 13632 25379
rect 13672 25347 13704 25379
rect 13744 25347 13776 25379
rect 13816 25347 13848 25379
rect 13888 25347 13920 25379
rect 13960 25347 13992 25379
rect 14032 25347 14064 25379
rect 14104 25347 14136 25379
rect 14176 25347 14208 25379
rect 14248 25347 14280 25379
rect 14320 25347 14352 25379
rect 14392 25347 14424 25379
rect 14464 25347 14496 25379
rect 14536 25347 14568 25379
rect 14608 25347 14640 25379
rect 14680 25347 14712 25379
rect 14752 25347 14784 25379
rect 14824 25347 14856 25379
rect 14896 25347 14928 25379
rect 14968 25347 15000 25379
rect 15040 25347 15072 25379
rect 15112 25347 15144 25379
rect 15184 25347 15216 25379
rect 15256 25347 15288 25379
rect 15328 25347 15360 25379
rect 15400 25347 15432 25379
rect 15472 25347 15504 25379
rect 15544 25347 15576 25379
rect 15616 25347 15648 25379
rect 15688 25347 15720 25379
rect 15760 25347 15792 25379
rect 15832 25347 15864 25379
rect 15904 25347 15936 25379
rect 64 25275 96 25307
rect 136 25275 168 25307
rect 208 25275 240 25307
rect 280 25275 312 25307
rect 352 25275 384 25307
rect 424 25275 456 25307
rect 496 25275 528 25307
rect 568 25275 600 25307
rect 640 25275 672 25307
rect 712 25275 744 25307
rect 784 25275 816 25307
rect 856 25275 888 25307
rect 928 25275 960 25307
rect 1000 25275 1032 25307
rect 1072 25275 1104 25307
rect 1144 25275 1176 25307
rect 1216 25275 1248 25307
rect 1288 25275 1320 25307
rect 1360 25275 1392 25307
rect 1432 25275 1464 25307
rect 1504 25275 1536 25307
rect 1576 25275 1608 25307
rect 1648 25275 1680 25307
rect 1720 25275 1752 25307
rect 1792 25275 1824 25307
rect 1864 25275 1896 25307
rect 1936 25275 1968 25307
rect 2008 25275 2040 25307
rect 2080 25275 2112 25307
rect 2152 25275 2184 25307
rect 2224 25275 2256 25307
rect 2296 25275 2328 25307
rect 2368 25275 2400 25307
rect 2440 25275 2472 25307
rect 2512 25275 2544 25307
rect 2584 25275 2616 25307
rect 2656 25275 2688 25307
rect 2728 25275 2760 25307
rect 2800 25275 2832 25307
rect 2872 25275 2904 25307
rect 2944 25275 2976 25307
rect 3016 25275 3048 25307
rect 3088 25275 3120 25307
rect 3160 25275 3192 25307
rect 3232 25275 3264 25307
rect 3304 25275 3336 25307
rect 3376 25275 3408 25307
rect 3448 25275 3480 25307
rect 3520 25275 3552 25307
rect 3592 25275 3624 25307
rect 3664 25275 3696 25307
rect 3736 25275 3768 25307
rect 3808 25275 3840 25307
rect 3880 25275 3912 25307
rect 3952 25275 3984 25307
rect 4024 25275 4056 25307
rect 4096 25275 4128 25307
rect 4168 25275 4200 25307
rect 4240 25275 4272 25307
rect 4312 25275 4344 25307
rect 4384 25275 4416 25307
rect 4456 25275 4488 25307
rect 4528 25275 4560 25307
rect 4600 25275 4632 25307
rect 4672 25275 4704 25307
rect 4744 25275 4776 25307
rect 4816 25275 4848 25307
rect 4888 25275 4920 25307
rect 4960 25275 4992 25307
rect 5032 25275 5064 25307
rect 5104 25275 5136 25307
rect 5176 25275 5208 25307
rect 5248 25275 5280 25307
rect 5320 25275 5352 25307
rect 5392 25275 5424 25307
rect 5464 25275 5496 25307
rect 5536 25275 5568 25307
rect 5608 25275 5640 25307
rect 5680 25275 5712 25307
rect 5752 25275 5784 25307
rect 5824 25275 5856 25307
rect 5896 25275 5928 25307
rect 5968 25275 6000 25307
rect 6040 25275 6072 25307
rect 6112 25275 6144 25307
rect 6184 25275 6216 25307
rect 6256 25275 6288 25307
rect 6328 25275 6360 25307
rect 6400 25275 6432 25307
rect 6472 25275 6504 25307
rect 6544 25275 6576 25307
rect 6616 25275 6648 25307
rect 6688 25275 6720 25307
rect 6760 25275 6792 25307
rect 6832 25275 6864 25307
rect 6904 25275 6936 25307
rect 6976 25275 7008 25307
rect 7048 25275 7080 25307
rect 7120 25275 7152 25307
rect 7192 25275 7224 25307
rect 7264 25275 7296 25307
rect 7336 25275 7368 25307
rect 7408 25275 7440 25307
rect 7480 25275 7512 25307
rect 7552 25275 7584 25307
rect 7624 25275 7656 25307
rect 7696 25275 7728 25307
rect 7768 25275 7800 25307
rect 7840 25275 7872 25307
rect 7912 25275 7944 25307
rect 7984 25275 8016 25307
rect 8056 25275 8088 25307
rect 8128 25275 8160 25307
rect 8200 25275 8232 25307
rect 8272 25275 8304 25307
rect 8344 25275 8376 25307
rect 8416 25275 8448 25307
rect 8488 25275 8520 25307
rect 8560 25275 8592 25307
rect 8632 25275 8664 25307
rect 8704 25275 8736 25307
rect 8776 25275 8808 25307
rect 8848 25275 8880 25307
rect 8920 25275 8952 25307
rect 8992 25275 9024 25307
rect 9064 25275 9096 25307
rect 9136 25275 9168 25307
rect 9208 25275 9240 25307
rect 9280 25275 9312 25307
rect 9352 25275 9384 25307
rect 9424 25275 9456 25307
rect 9496 25275 9528 25307
rect 9568 25275 9600 25307
rect 9640 25275 9672 25307
rect 9712 25275 9744 25307
rect 9784 25275 9816 25307
rect 9856 25275 9888 25307
rect 9928 25275 9960 25307
rect 10000 25275 10032 25307
rect 10072 25275 10104 25307
rect 10144 25275 10176 25307
rect 10216 25275 10248 25307
rect 10288 25275 10320 25307
rect 10360 25275 10392 25307
rect 10432 25275 10464 25307
rect 10504 25275 10536 25307
rect 10576 25275 10608 25307
rect 10648 25275 10680 25307
rect 10720 25275 10752 25307
rect 10792 25275 10824 25307
rect 10864 25275 10896 25307
rect 10936 25275 10968 25307
rect 11008 25275 11040 25307
rect 11080 25275 11112 25307
rect 11152 25275 11184 25307
rect 11224 25275 11256 25307
rect 11296 25275 11328 25307
rect 11368 25275 11400 25307
rect 11440 25275 11472 25307
rect 11512 25275 11544 25307
rect 11584 25275 11616 25307
rect 11656 25275 11688 25307
rect 11728 25275 11760 25307
rect 11800 25275 11832 25307
rect 11872 25275 11904 25307
rect 11944 25275 11976 25307
rect 12016 25275 12048 25307
rect 12088 25275 12120 25307
rect 12160 25275 12192 25307
rect 12232 25275 12264 25307
rect 12304 25275 12336 25307
rect 12376 25275 12408 25307
rect 12448 25275 12480 25307
rect 12520 25275 12552 25307
rect 12592 25275 12624 25307
rect 12664 25275 12696 25307
rect 12736 25275 12768 25307
rect 12808 25275 12840 25307
rect 12880 25275 12912 25307
rect 12952 25275 12984 25307
rect 13024 25275 13056 25307
rect 13096 25275 13128 25307
rect 13168 25275 13200 25307
rect 13240 25275 13272 25307
rect 13312 25275 13344 25307
rect 13384 25275 13416 25307
rect 13456 25275 13488 25307
rect 13528 25275 13560 25307
rect 13600 25275 13632 25307
rect 13672 25275 13704 25307
rect 13744 25275 13776 25307
rect 13816 25275 13848 25307
rect 13888 25275 13920 25307
rect 13960 25275 13992 25307
rect 14032 25275 14064 25307
rect 14104 25275 14136 25307
rect 14176 25275 14208 25307
rect 14248 25275 14280 25307
rect 14320 25275 14352 25307
rect 14392 25275 14424 25307
rect 14464 25275 14496 25307
rect 14536 25275 14568 25307
rect 14608 25275 14640 25307
rect 14680 25275 14712 25307
rect 14752 25275 14784 25307
rect 14824 25275 14856 25307
rect 14896 25275 14928 25307
rect 14968 25275 15000 25307
rect 15040 25275 15072 25307
rect 15112 25275 15144 25307
rect 15184 25275 15216 25307
rect 15256 25275 15288 25307
rect 15328 25275 15360 25307
rect 15400 25275 15432 25307
rect 15472 25275 15504 25307
rect 15544 25275 15576 25307
rect 15616 25275 15648 25307
rect 15688 25275 15720 25307
rect 15760 25275 15792 25307
rect 15832 25275 15864 25307
rect 15904 25275 15936 25307
rect 64 25203 96 25235
rect 136 25203 168 25235
rect 208 25203 240 25235
rect 280 25203 312 25235
rect 352 25203 384 25235
rect 424 25203 456 25235
rect 496 25203 528 25235
rect 568 25203 600 25235
rect 640 25203 672 25235
rect 712 25203 744 25235
rect 784 25203 816 25235
rect 856 25203 888 25235
rect 928 25203 960 25235
rect 1000 25203 1032 25235
rect 1072 25203 1104 25235
rect 1144 25203 1176 25235
rect 1216 25203 1248 25235
rect 1288 25203 1320 25235
rect 1360 25203 1392 25235
rect 1432 25203 1464 25235
rect 1504 25203 1536 25235
rect 1576 25203 1608 25235
rect 1648 25203 1680 25235
rect 1720 25203 1752 25235
rect 1792 25203 1824 25235
rect 1864 25203 1896 25235
rect 1936 25203 1968 25235
rect 2008 25203 2040 25235
rect 2080 25203 2112 25235
rect 2152 25203 2184 25235
rect 2224 25203 2256 25235
rect 2296 25203 2328 25235
rect 2368 25203 2400 25235
rect 2440 25203 2472 25235
rect 2512 25203 2544 25235
rect 2584 25203 2616 25235
rect 2656 25203 2688 25235
rect 2728 25203 2760 25235
rect 2800 25203 2832 25235
rect 2872 25203 2904 25235
rect 2944 25203 2976 25235
rect 3016 25203 3048 25235
rect 3088 25203 3120 25235
rect 3160 25203 3192 25235
rect 3232 25203 3264 25235
rect 3304 25203 3336 25235
rect 3376 25203 3408 25235
rect 3448 25203 3480 25235
rect 3520 25203 3552 25235
rect 3592 25203 3624 25235
rect 3664 25203 3696 25235
rect 3736 25203 3768 25235
rect 3808 25203 3840 25235
rect 3880 25203 3912 25235
rect 3952 25203 3984 25235
rect 4024 25203 4056 25235
rect 4096 25203 4128 25235
rect 4168 25203 4200 25235
rect 4240 25203 4272 25235
rect 4312 25203 4344 25235
rect 4384 25203 4416 25235
rect 4456 25203 4488 25235
rect 4528 25203 4560 25235
rect 4600 25203 4632 25235
rect 4672 25203 4704 25235
rect 4744 25203 4776 25235
rect 4816 25203 4848 25235
rect 4888 25203 4920 25235
rect 4960 25203 4992 25235
rect 5032 25203 5064 25235
rect 5104 25203 5136 25235
rect 5176 25203 5208 25235
rect 5248 25203 5280 25235
rect 5320 25203 5352 25235
rect 5392 25203 5424 25235
rect 5464 25203 5496 25235
rect 5536 25203 5568 25235
rect 5608 25203 5640 25235
rect 5680 25203 5712 25235
rect 5752 25203 5784 25235
rect 5824 25203 5856 25235
rect 5896 25203 5928 25235
rect 5968 25203 6000 25235
rect 6040 25203 6072 25235
rect 6112 25203 6144 25235
rect 6184 25203 6216 25235
rect 6256 25203 6288 25235
rect 6328 25203 6360 25235
rect 6400 25203 6432 25235
rect 6472 25203 6504 25235
rect 6544 25203 6576 25235
rect 6616 25203 6648 25235
rect 6688 25203 6720 25235
rect 6760 25203 6792 25235
rect 6832 25203 6864 25235
rect 6904 25203 6936 25235
rect 6976 25203 7008 25235
rect 7048 25203 7080 25235
rect 7120 25203 7152 25235
rect 7192 25203 7224 25235
rect 7264 25203 7296 25235
rect 7336 25203 7368 25235
rect 7408 25203 7440 25235
rect 7480 25203 7512 25235
rect 7552 25203 7584 25235
rect 7624 25203 7656 25235
rect 7696 25203 7728 25235
rect 7768 25203 7800 25235
rect 7840 25203 7872 25235
rect 7912 25203 7944 25235
rect 7984 25203 8016 25235
rect 8056 25203 8088 25235
rect 8128 25203 8160 25235
rect 8200 25203 8232 25235
rect 8272 25203 8304 25235
rect 8344 25203 8376 25235
rect 8416 25203 8448 25235
rect 8488 25203 8520 25235
rect 8560 25203 8592 25235
rect 8632 25203 8664 25235
rect 8704 25203 8736 25235
rect 8776 25203 8808 25235
rect 8848 25203 8880 25235
rect 8920 25203 8952 25235
rect 8992 25203 9024 25235
rect 9064 25203 9096 25235
rect 9136 25203 9168 25235
rect 9208 25203 9240 25235
rect 9280 25203 9312 25235
rect 9352 25203 9384 25235
rect 9424 25203 9456 25235
rect 9496 25203 9528 25235
rect 9568 25203 9600 25235
rect 9640 25203 9672 25235
rect 9712 25203 9744 25235
rect 9784 25203 9816 25235
rect 9856 25203 9888 25235
rect 9928 25203 9960 25235
rect 10000 25203 10032 25235
rect 10072 25203 10104 25235
rect 10144 25203 10176 25235
rect 10216 25203 10248 25235
rect 10288 25203 10320 25235
rect 10360 25203 10392 25235
rect 10432 25203 10464 25235
rect 10504 25203 10536 25235
rect 10576 25203 10608 25235
rect 10648 25203 10680 25235
rect 10720 25203 10752 25235
rect 10792 25203 10824 25235
rect 10864 25203 10896 25235
rect 10936 25203 10968 25235
rect 11008 25203 11040 25235
rect 11080 25203 11112 25235
rect 11152 25203 11184 25235
rect 11224 25203 11256 25235
rect 11296 25203 11328 25235
rect 11368 25203 11400 25235
rect 11440 25203 11472 25235
rect 11512 25203 11544 25235
rect 11584 25203 11616 25235
rect 11656 25203 11688 25235
rect 11728 25203 11760 25235
rect 11800 25203 11832 25235
rect 11872 25203 11904 25235
rect 11944 25203 11976 25235
rect 12016 25203 12048 25235
rect 12088 25203 12120 25235
rect 12160 25203 12192 25235
rect 12232 25203 12264 25235
rect 12304 25203 12336 25235
rect 12376 25203 12408 25235
rect 12448 25203 12480 25235
rect 12520 25203 12552 25235
rect 12592 25203 12624 25235
rect 12664 25203 12696 25235
rect 12736 25203 12768 25235
rect 12808 25203 12840 25235
rect 12880 25203 12912 25235
rect 12952 25203 12984 25235
rect 13024 25203 13056 25235
rect 13096 25203 13128 25235
rect 13168 25203 13200 25235
rect 13240 25203 13272 25235
rect 13312 25203 13344 25235
rect 13384 25203 13416 25235
rect 13456 25203 13488 25235
rect 13528 25203 13560 25235
rect 13600 25203 13632 25235
rect 13672 25203 13704 25235
rect 13744 25203 13776 25235
rect 13816 25203 13848 25235
rect 13888 25203 13920 25235
rect 13960 25203 13992 25235
rect 14032 25203 14064 25235
rect 14104 25203 14136 25235
rect 14176 25203 14208 25235
rect 14248 25203 14280 25235
rect 14320 25203 14352 25235
rect 14392 25203 14424 25235
rect 14464 25203 14496 25235
rect 14536 25203 14568 25235
rect 14608 25203 14640 25235
rect 14680 25203 14712 25235
rect 14752 25203 14784 25235
rect 14824 25203 14856 25235
rect 14896 25203 14928 25235
rect 14968 25203 15000 25235
rect 15040 25203 15072 25235
rect 15112 25203 15144 25235
rect 15184 25203 15216 25235
rect 15256 25203 15288 25235
rect 15328 25203 15360 25235
rect 15400 25203 15432 25235
rect 15472 25203 15504 25235
rect 15544 25203 15576 25235
rect 15616 25203 15648 25235
rect 15688 25203 15720 25235
rect 15760 25203 15792 25235
rect 15832 25203 15864 25235
rect 15904 25203 15936 25235
rect 64 25131 96 25163
rect 136 25131 168 25163
rect 208 25131 240 25163
rect 280 25131 312 25163
rect 352 25131 384 25163
rect 424 25131 456 25163
rect 496 25131 528 25163
rect 568 25131 600 25163
rect 640 25131 672 25163
rect 712 25131 744 25163
rect 784 25131 816 25163
rect 856 25131 888 25163
rect 928 25131 960 25163
rect 1000 25131 1032 25163
rect 1072 25131 1104 25163
rect 1144 25131 1176 25163
rect 1216 25131 1248 25163
rect 1288 25131 1320 25163
rect 1360 25131 1392 25163
rect 1432 25131 1464 25163
rect 1504 25131 1536 25163
rect 1576 25131 1608 25163
rect 1648 25131 1680 25163
rect 1720 25131 1752 25163
rect 1792 25131 1824 25163
rect 1864 25131 1896 25163
rect 1936 25131 1968 25163
rect 2008 25131 2040 25163
rect 2080 25131 2112 25163
rect 2152 25131 2184 25163
rect 2224 25131 2256 25163
rect 2296 25131 2328 25163
rect 2368 25131 2400 25163
rect 2440 25131 2472 25163
rect 2512 25131 2544 25163
rect 2584 25131 2616 25163
rect 2656 25131 2688 25163
rect 2728 25131 2760 25163
rect 2800 25131 2832 25163
rect 2872 25131 2904 25163
rect 2944 25131 2976 25163
rect 3016 25131 3048 25163
rect 3088 25131 3120 25163
rect 3160 25131 3192 25163
rect 3232 25131 3264 25163
rect 3304 25131 3336 25163
rect 3376 25131 3408 25163
rect 3448 25131 3480 25163
rect 3520 25131 3552 25163
rect 3592 25131 3624 25163
rect 3664 25131 3696 25163
rect 3736 25131 3768 25163
rect 3808 25131 3840 25163
rect 3880 25131 3912 25163
rect 3952 25131 3984 25163
rect 4024 25131 4056 25163
rect 4096 25131 4128 25163
rect 4168 25131 4200 25163
rect 4240 25131 4272 25163
rect 4312 25131 4344 25163
rect 4384 25131 4416 25163
rect 4456 25131 4488 25163
rect 4528 25131 4560 25163
rect 4600 25131 4632 25163
rect 4672 25131 4704 25163
rect 4744 25131 4776 25163
rect 4816 25131 4848 25163
rect 4888 25131 4920 25163
rect 4960 25131 4992 25163
rect 5032 25131 5064 25163
rect 5104 25131 5136 25163
rect 5176 25131 5208 25163
rect 5248 25131 5280 25163
rect 5320 25131 5352 25163
rect 5392 25131 5424 25163
rect 5464 25131 5496 25163
rect 5536 25131 5568 25163
rect 5608 25131 5640 25163
rect 5680 25131 5712 25163
rect 5752 25131 5784 25163
rect 5824 25131 5856 25163
rect 5896 25131 5928 25163
rect 5968 25131 6000 25163
rect 6040 25131 6072 25163
rect 6112 25131 6144 25163
rect 6184 25131 6216 25163
rect 6256 25131 6288 25163
rect 6328 25131 6360 25163
rect 6400 25131 6432 25163
rect 6472 25131 6504 25163
rect 6544 25131 6576 25163
rect 6616 25131 6648 25163
rect 6688 25131 6720 25163
rect 6760 25131 6792 25163
rect 6832 25131 6864 25163
rect 6904 25131 6936 25163
rect 6976 25131 7008 25163
rect 7048 25131 7080 25163
rect 7120 25131 7152 25163
rect 7192 25131 7224 25163
rect 7264 25131 7296 25163
rect 7336 25131 7368 25163
rect 7408 25131 7440 25163
rect 7480 25131 7512 25163
rect 7552 25131 7584 25163
rect 7624 25131 7656 25163
rect 7696 25131 7728 25163
rect 7768 25131 7800 25163
rect 7840 25131 7872 25163
rect 7912 25131 7944 25163
rect 7984 25131 8016 25163
rect 8056 25131 8088 25163
rect 8128 25131 8160 25163
rect 8200 25131 8232 25163
rect 8272 25131 8304 25163
rect 8344 25131 8376 25163
rect 8416 25131 8448 25163
rect 8488 25131 8520 25163
rect 8560 25131 8592 25163
rect 8632 25131 8664 25163
rect 8704 25131 8736 25163
rect 8776 25131 8808 25163
rect 8848 25131 8880 25163
rect 8920 25131 8952 25163
rect 8992 25131 9024 25163
rect 9064 25131 9096 25163
rect 9136 25131 9168 25163
rect 9208 25131 9240 25163
rect 9280 25131 9312 25163
rect 9352 25131 9384 25163
rect 9424 25131 9456 25163
rect 9496 25131 9528 25163
rect 9568 25131 9600 25163
rect 9640 25131 9672 25163
rect 9712 25131 9744 25163
rect 9784 25131 9816 25163
rect 9856 25131 9888 25163
rect 9928 25131 9960 25163
rect 10000 25131 10032 25163
rect 10072 25131 10104 25163
rect 10144 25131 10176 25163
rect 10216 25131 10248 25163
rect 10288 25131 10320 25163
rect 10360 25131 10392 25163
rect 10432 25131 10464 25163
rect 10504 25131 10536 25163
rect 10576 25131 10608 25163
rect 10648 25131 10680 25163
rect 10720 25131 10752 25163
rect 10792 25131 10824 25163
rect 10864 25131 10896 25163
rect 10936 25131 10968 25163
rect 11008 25131 11040 25163
rect 11080 25131 11112 25163
rect 11152 25131 11184 25163
rect 11224 25131 11256 25163
rect 11296 25131 11328 25163
rect 11368 25131 11400 25163
rect 11440 25131 11472 25163
rect 11512 25131 11544 25163
rect 11584 25131 11616 25163
rect 11656 25131 11688 25163
rect 11728 25131 11760 25163
rect 11800 25131 11832 25163
rect 11872 25131 11904 25163
rect 11944 25131 11976 25163
rect 12016 25131 12048 25163
rect 12088 25131 12120 25163
rect 12160 25131 12192 25163
rect 12232 25131 12264 25163
rect 12304 25131 12336 25163
rect 12376 25131 12408 25163
rect 12448 25131 12480 25163
rect 12520 25131 12552 25163
rect 12592 25131 12624 25163
rect 12664 25131 12696 25163
rect 12736 25131 12768 25163
rect 12808 25131 12840 25163
rect 12880 25131 12912 25163
rect 12952 25131 12984 25163
rect 13024 25131 13056 25163
rect 13096 25131 13128 25163
rect 13168 25131 13200 25163
rect 13240 25131 13272 25163
rect 13312 25131 13344 25163
rect 13384 25131 13416 25163
rect 13456 25131 13488 25163
rect 13528 25131 13560 25163
rect 13600 25131 13632 25163
rect 13672 25131 13704 25163
rect 13744 25131 13776 25163
rect 13816 25131 13848 25163
rect 13888 25131 13920 25163
rect 13960 25131 13992 25163
rect 14032 25131 14064 25163
rect 14104 25131 14136 25163
rect 14176 25131 14208 25163
rect 14248 25131 14280 25163
rect 14320 25131 14352 25163
rect 14392 25131 14424 25163
rect 14464 25131 14496 25163
rect 14536 25131 14568 25163
rect 14608 25131 14640 25163
rect 14680 25131 14712 25163
rect 14752 25131 14784 25163
rect 14824 25131 14856 25163
rect 14896 25131 14928 25163
rect 14968 25131 15000 25163
rect 15040 25131 15072 25163
rect 15112 25131 15144 25163
rect 15184 25131 15216 25163
rect 15256 25131 15288 25163
rect 15328 25131 15360 25163
rect 15400 25131 15432 25163
rect 15472 25131 15504 25163
rect 15544 25131 15576 25163
rect 15616 25131 15648 25163
rect 15688 25131 15720 25163
rect 15760 25131 15792 25163
rect 15832 25131 15864 25163
rect 15904 25131 15936 25163
rect 64 25059 96 25091
rect 136 25059 168 25091
rect 208 25059 240 25091
rect 280 25059 312 25091
rect 352 25059 384 25091
rect 424 25059 456 25091
rect 496 25059 528 25091
rect 568 25059 600 25091
rect 640 25059 672 25091
rect 712 25059 744 25091
rect 784 25059 816 25091
rect 856 25059 888 25091
rect 928 25059 960 25091
rect 1000 25059 1032 25091
rect 1072 25059 1104 25091
rect 1144 25059 1176 25091
rect 1216 25059 1248 25091
rect 1288 25059 1320 25091
rect 1360 25059 1392 25091
rect 1432 25059 1464 25091
rect 1504 25059 1536 25091
rect 1576 25059 1608 25091
rect 1648 25059 1680 25091
rect 1720 25059 1752 25091
rect 1792 25059 1824 25091
rect 1864 25059 1896 25091
rect 1936 25059 1968 25091
rect 2008 25059 2040 25091
rect 2080 25059 2112 25091
rect 2152 25059 2184 25091
rect 2224 25059 2256 25091
rect 2296 25059 2328 25091
rect 2368 25059 2400 25091
rect 2440 25059 2472 25091
rect 2512 25059 2544 25091
rect 2584 25059 2616 25091
rect 2656 25059 2688 25091
rect 2728 25059 2760 25091
rect 2800 25059 2832 25091
rect 2872 25059 2904 25091
rect 2944 25059 2976 25091
rect 3016 25059 3048 25091
rect 3088 25059 3120 25091
rect 3160 25059 3192 25091
rect 3232 25059 3264 25091
rect 3304 25059 3336 25091
rect 3376 25059 3408 25091
rect 3448 25059 3480 25091
rect 3520 25059 3552 25091
rect 3592 25059 3624 25091
rect 3664 25059 3696 25091
rect 3736 25059 3768 25091
rect 3808 25059 3840 25091
rect 3880 25059 3912 25091
rect 3952 25059 3984 25091
rect 4024 25059 4056 25091
rect 4096 25059 4128 25091
rect 4168 25059 4200 25091
rect 4240 25059 4272 25091
rect 4312 25059 4344 25091
rect 4384 25059 4416 25091
rect 4456 25059 4488 25091
rect 4528 25059 4560 25091
rect 4600 25059 4632 25091
rect 4672 25059 4704 25091
rect 4744 25059 4776 25091
rect 4816 25059 4848 25091
rect 4888 25059 4920 25091
rect 4960 25059 4992 25091
rect 5032 25059 5064 25091
rect 5104 25059 5136 25091
rect 5176 25059 5208 25091
rect 5248 25059 5280 25091
rect 5320 25059 5352 25091
rect 5392 25059 5424 25091
rect 5464 25059 5496 25091
rect 5536 25059 5568 25091
rect 5608 25059 5640 25091
rect 5680 25059 5712 25091
rect 5752 25059 5784 25091
rect 5824 25059 5856 25091
rect 5896 25059 5928 25091
rect 5968 25059 6000 25091
rect 6040 25059 6072 25091
rect 6112 25059 6144 25091
rect 6184 25059 6216 25091
rect 6256 25059 6288 25091
rect 6328 25059 6360 25091
rect 6400 25059 6432 25091
rect 6472 25059 6504 25091
rect 6544 25059 6576 25091
rect 6616 25059 6648 25091
rect 6688 25059 6720 25091
rect 6760 25059 6792 25091
rect 6832 25059 6864 25091
rect 6904 25059 6936 25091
rect 6976 25059 7008 25091
rect 7048 25059 7080 25091
rect 7120 25059 7152 25091
rect 7192 25059 7224 25091
rect 7264 25059 7296 25091
rect 7336 25059 7368 25091
rect 7408 25059 7440 25091
rect 7480 25059 7512 25091
rect 7552 25059 7584 25091
rect 7624 25059 7656 25091
rect 7696 25059 7728 25091
rect 7768 25059 7800 25091
rect 7840 25059 7872 25091
rect 7912 25059 7944 25091
rect 7984 25059 8016 25091
rect 8056 25059 8088 25091
rect 8128 25059 8160 25091
rect 8200 25059 8232 25091
rect 8272 25059 8304 25091
rect 8344 25059 8376 25091
rect 8416 25059 8448 25091
rect 8488 25059 8520 25091
rect 8560 25059 8592 25091
rect 8632 25059 8664 25091
rect 8704 25059 8736 25091
rect 8776 25059 8808 25091
rect 8848 25059 8880 25091
rect 8920 25059 8952 25091
rect 8992 25059 9024 25091
rect 9064 25059 9096 25091
rect 9136 25059 9168 25091
rect 9208 25059 9240 25091
rect 9280 25059 9312 25091
rect 9352 25059 9384 25091
rect 9424 25059 9456 25091
rect 9496 25059 9528 25091
rect 9568 25059 9600 25091
rect 9640 25059 9672 25091
rect 9712 25059 9744 25091
rect 9784 25059 9816 25091
rect 9856 25059 9888 25091
rect 9928 25059 9960 25091
rect 10000 25059 10032 25091
rect 10072 25059 10104 25091
rect 10144 25059 10176 25091
rect 10216 25059 10248 25091
rect 10288 25059 10320 25091
rect 10360 25059 10392 25091
rect 10432 25059 10464 25091
rect 10504 25059 10536 25091
rect 10576 25059 10608 25091
rect 10648 25059 10680 25091
rect 10720 25059 10752 25091
rect 10792 25059 10824 25091
rect 10864 25059 10896 25091
rect 10936 25059 10968 25091
rect 11008 25059 11040 25091
rect 11080 25059 11112 25091
rect 11152 25059 11184 25091
rect 11224 25059 11256 25091
rect 11296 25059 11328 25091
rect 11368 25059 11400 25091
rect 11440 25059 11472 25091
rect 11512 25059 11544 25091
rect 11584 25059 11616 25091
rect 11656 25059 11688 25091
rect 11728 25059 11760 25091
rect 11800 25059 11832 25091
rect 11872 25059 11904 25091
rect 11944 25059 11976 25091
rect 12016 25059 12048 25091
rect 12088 25059 12120 25091
rect 12160 25059 12192 25091
rect 12232 25059 12264 25091
rect 12304 25059 12336 25091
rect 12376 25059 12408 25091
rect 12448 25059 12480 25091
rect 12520 25059 12552 25091
rect 12592 25059 12624 25091
rect 12664 25059 12696 25091
rect 12736 25059 12768 25091
rect 12808 25059 12840 25091
rect 12880 25059 12912 25091
rect 12952 25059 12984 25091
rect 13024 25059 13056 25091
rect 13096 25059 13128 25091
rect 13168 25059 13200 25091
rect 13240 25059 13272 25091
rect 13312 25059 13344 25091
rect 13384 25059 13416 25091
rect 13456 25059 13488 25091
rect 13528 25059 13560 25091
rect 13600 25059 13632 25091
rect 13672 25059 13704 25091
rect 13744 25059 13776 25091
rect 13816 25059 13848 25091
rect 13888 25059 13920 25091
rect 13960 25059 13992 25091
rect 14032 25059 14064 25091
rect 14104 25059 14136 25091
rect 14176 25059 14208 25091
rect 14248 25059 14280 25091
rect 14320 25059 14352 25091
rect 14392 25059 14424 25091
rect 14464 25059 14496 25091
rect 14536 25059 14568 25091
rect 14608 25059 14640 25091
rect 14680 25059 14712 25091
rect 14752 25059 14784 25091
rect 14824 25059 14856 25091
rect 14896 25059 14928 25091
rect 14968 25059 15000 25091
rect 15040 25059 15072 25091
rect 15112 25059 15144 25091
rect 15184 25059 15216 25091
rect 15256 25059 15288 25091
rect 15328 25059 15360 25091
rect 15400 25059 15432 25091
rect 15472 25059 15504 25091
rect 15544 25059 15576 25091
rect 15616 25059 15648 25091
rect 15688 25059 15720 25091
rect 15760 25059 15792 25091
rect 15832 25059 15864 25091
rect 15904 25059 15936 25091
rect 64 24987 96 25019
rect 136 24987 168 25019
rect 208 24987 240 25019
rect 280 24987 312 25019
rect 352 24987 384 25019
rect 424 24987 456 25019
rect 496 24987 528 25019
rect 568 24987 600 25019
rect 640 24987 672 25019
rect 712 24987 744 25019
rect 784 24987 816 25019
rect 856 24987 888 25019
rect 928 24987 960 25019
rect 1000 24987 1032 25019
rect 1072 24987 1104 25019
rect 1144 24987 1176 25019
rect 1216 24987 1248 25019
rect 1288 24987 1320 25019
rect 1360 24987 1392 25019
rect 1432 24987 1464 25019
rect 1504 24987 1536 25019
rect 1576 24987 1608 25019
rect 1648 24987 1680 25019
rect 1720 24987 1752 25019
rect 1792 24987 1824 25019
rect 1864 24987 1896 25019
rect 1936 24987 1968 25019
rect 2008 24987 2040 25019
rect 2080 24987 2112 25019
rect 2152 24987 2184 25019
rect 2224 24987 2256 25019
rect 2296 24987 2328 25019
rect 2368 24987 2400 25019
rect 2440 24987 2472 25019
rect 2512 24987 2544 25019
rect 2584 24987 2616 25019
rect 2656 24987 2688 25019
rect 2728 24987 2760 25019
rect 2800 24987 2832 25019
rect 2872 24987 2904 25019
rect 2944 24987 2976 25019
rect 3016 24987 3048 25019
rect 3088 24987 3120 25019
rect 3160 24987 3192 25019
rect 3232 24987 3264 25019
rect 3304 24987 3336 25019
rect 3376 24987 3408 25019
rect 3448 24987 3480 25019
rect 3520 24987 3552 25019
rect 3592 24987 3624 25019
rect 3664 24987 3696 25019
rect 3736 24987 3768 25019
rect 3808 24987 3840 25019
rect 3880 24987 3912 25019
rect 3952 24987 3984 25019
rect 4024 24987 4056 25019
rect 4096 24987 4128 25019
rect 4168 24987 4200 25019
rect 4240 24987 4272 25019
rect 4312 24987 4344 25019
rect 4384 24987 4416 25019
rect 4456 24987 4488 25019
rect 4528 24987 4560 25019
rect 4600 24987 4632 25019
rect 4672 24987 4704 25019
rect 4744 24987 4776 25019
rect 4816 24987 4848 25019
rect 4888 24987 4920 25019
rect 4960 24987 4992 25019
rect 5032 24987 5064 25019
rect 5104 24987 5136 25019
rect 5176 24987 5208 25019
rect 5248 24987 5280 25019
rect 5320 24987 5352 25019
rect 5392 24987 5424 25019
rect 5464 24987 5496 25019
rect 5536 24987 5568 25019
rect 5608 24987 5640 25019
rect 5680 24987 5712 25019
rect 5752 24987 5784 25019
rect 5824 24987 5856 25019
rect 5896 24987 5928 25019
rect 5968 24987 6000 25019
rect 6040 24987 6072 25019
rect 6112 24987 6144 25019
rect 6184 24987 6216 25019
rect 6256 24987 6288 25019
rect 6328 24987 6360 25019
rect 6400 24987 6432 25019
rect 6472 24987 6504 25019
rect 6544 24987 6576 25019
rect 6616 24987 6648 25019
rect 6688 24987 6720 25019
rect 6760 24987 6792 25019
rect 6832 24987 6864 25019
rect 6904 24987 6936 25019
rect 6976 24987 7008 25019
rect 7048 24987 7080 25019
rect 7120 24987 7152 25019
rect 7192 24987 7224 25019
rect 7264 24987 7296 25019
rect 7336 24987 7368 25019
rect 7408 24987 7440 25019
rect 7480 24987 7512 25019
rect 7552 24987 7584 25019
rect 7624 24987 7656 25019
rect 7696 24987 7728 25019
rect 7768 24987 7800 25019
rect 7840 24987 7872 25019
rect 7912 24987 7944 25019
rect 7984 24987 8016 25019
rect 8056 24987 8088 25019
rect 8128 24987 8160 25019
rect 8200 24987 8232 25019
rect 8272 24987 8304 25019
rect 8344 24987 8376 25019
rect 8416 24987 8448 25019
rect 8488 24987 8520 25019
rect 8560 24987 8592 25019
rect 8632 24987 8664 25019
rect 8704 24987 8736 25019
rect 8776 24987 8808 25019
rect 8848 24987 8880 25019
rect 8920 24987 8952 25019
rect 8992 24987 9024 25019
rect 9064 24987 9096 25019
rect 9136 24987 9168 25019
rect 9208 24987 9240 25019
rect 9280 24987 9312 25019
rect 9352 24987 9384 25019
rect 9424 24987 9456 25019
rect 9496 24987 9528 25019
rect 9568 24987 9600 25019
rect 9640 24987 9672 25019
rect 9712 24987 9744 25019
rect 9784 24987 9816 25019
rect 9856 24987 9888 25019
rect 9928 24987 9960 25019
rect 10000 24987 10032 25019
rect 10072 24987 10104 25019
rect 10144 24987 10176 25019
rect 10216 24987 10248 25019
rect 10288 24987 10320 25019
rect 10360 24987 10392 25019
rect 10432 24987 10464 25019
rect 10504 24987 10536 25019
rect 10576 24987 10608 25019
rect 10648 24987 10680 25019
rect 10720 24987 10752 25019
rect 10792 24987 10824 25019
rect 10864 24987 10896 25019
rect 10936 24987 10968 25019
rect 11008 24987 11040 25019
rect 11080 24987 11112 25019
rect 11152 24987 11184 25019
rect 11224 24987 11256 25019
rect 11296 24987 11328 25019
rect 11368 24987 11400 25019
rect 11440 24987 11472 25019
rect 11512 24987 11544 25019
rect 11584 24987 11616 25019
rect 11656 24987 11688 25019
rect 11728 24987 11760 25019
rect 11800 24987 11832 25019
rect 11872 24987 11904 25019
rect 11944 24987 11976 25019
rect 12016 24987 12048 25019
rect 12088 24987 12120 25019
rect 12160 24987 12192 25019
rect 12232 24987 12264 25019
rect 12304 24987 12336 25019
rect 12376 24987 12408 25019
rect 12448 24987 12480 25019
rect 12520 24987 12552 25019
rect 12592 24987 12624 25019
rect 12664 24987 12696 25019
rect 12736 24987 12768 25019
rect 12808 24987 12840 25019
rect 12880 24987 12912 25019
rect 12952 24987 12984 25019
rect 13024 24987 13056 25019
rect 13096 24987 13128 25019
rect 13168 24987 13200 25019
rect 13240 24987 13272 25019
rect 13312 24987 13344 25019
rect 13384 24987 13416 25019
rect 13456 24987 13488 25019
rect 13528 24987 13560 25019
rect 13600 24987 13632 25019
rect 13672 24987 13704 25019
rect 13744 24987 13776 25019
rect 13816 24987 13848 25019
rect 13888 24987 13920 25019
rect 13960 24987 13992 25019
rect 14032 24987 14064 25019
rect 14104 24987 14136 25019
rect 14176 24987 14208 25019
rect 14248 24987 14280 25019
rect 14320 24987 14352 25019
rect 14392 24987 14424 25019
rect 14464 24987 14496 25019
rect 14536 24987 14568 25019
rect 14608 24987 14640 25019
rect 14680 24987 14712 25019
rect 14752 24987 14784 25019
rect 14824 24987 14856 25019
rect 14896 24987 14928 25019
rect 14968 24987 15000 25019
rect 15040 24987 15072 25019
rect 15112 24987 15144 25019
rect 15184 24987 15216 25019
rect 15256 24987 15288 25019
rect 15328 24987 15360 25019
rect 15400 24987 15432 25019
rect 15472 24987 15504 25019
rect 15544 24987 15576 25019
rect 15616 24987 15648 25019
rect 15688 24987 15720 25019
rect 15760 24987 15792 25019
rect 15832 24987 15864 25019
rect 15904 24987 15936 25019
rect 64 24915 96 24947
rect 136 24915 168 24947
rect 208 24915 240 24947
rect 280 24915 312 24947
rect 352 24915 384 24947
rect 424 24915 456 24947
rect 496 24915 528 24947
rect 568 24915 600 24947
rect 640 24915 672 24947
rect 712 24915 744 24947
rect 784 24915 816 24947
rect 856 24915 888 24947
rect 928 24915 960 24947
rect 1000 24915 1032 24947
rect 1072 24915 1104 24947
rect 1144 24915 1176 24947
rect 1216 24915 1248 24947
rect 1288 24915 1320 24947
rect 1360 24915 1392 24947
rect 1432 24915 1464 24947
rect 1504 24915 1536 24947
rect 1576 24915 1608 24947
rect 1648 24915 1680 24947
rect 1720 24915 1752 24947
rect 1792 24915 1824 24947
rect 1864 24915 1896 24947
rect 1936 24915 1968 24947
rect 2008 24915 2040 24947
rect 2080 24915 2112 24947
rect 2152 24915 2184 24947
rect 2224 24915 2256 24947
rect 2296 24915 2328 24947
rect 2368 24915 2400 24947
rect 2440 24915 2472 24947
rect 2512 24915 2544 24947
rect 2584 24915 2616 24947
rect 2656 24915 2688 24947
rect 2728 24915 2760 24947
rect 2800 24915 2832 24947
rect 2872 24915 2904 24947
rect 2944 24915 2976 24947
rect 3016 24915 3048 24947
rect 3088 24915 3120 24947
rect 3160 24915 3192 24947
rect 3232 24915 3264 24947
rect 3304 24915 3336 24947
rect 3376 24915 3408 24947
rect 3448 24915 3480 24947
rect 3520 24915 3552 24947
rect 3592 24915 3624 24947
rect 3664 24915 3696 24947
rect 3736 24915 3768 24947
rect 3808 24915 3840 24947
rect 3880 24915 3912 24947
rect 3952 24915 3984 24947
rect 4024 24915 4056 24947
rect 4096 24915 4128 24947
rect 4168 24915 4200 24947
rect 4240 24915 4272 24947
rect 4312 24915 4344 24947
rect 4384 24915 4416 24947
rect 4456 24915 4488 24947
rect 4528 24915 4560 24947
rect 4600 24915 4632 24947
rect 4672 24915 4704 24947
rect 4744 24915 4776 24947
rect 4816 24915 4848 24947
rect 4888 24915 4920 24947
rect 4960 24915 4992 24947
rect 5032 24915 5064 24947
rect 5104 24915 5136 24947
rect 5176 24915 5208 24947
rect 5248 24915 5280 24947
rect 5320 24915 5352 24947
rect 5392 24915 5424 24947
rect 5464 24915 5496 24947
rect 5536 24915 5568 24947
rect 5608 24915 5640 24947
rect 5680 24915 5712 24947
rect 5752 24915 5784 24947
rect 5824 24915 5856 24947
rect 5896 24915 5928 24947
rect 5968 24915 6000 24947
rect 6040 24915 6072 24947
rect 6112 24915 6144 24947
rect 6184 24915 6216 24947
rect 6256 24915 6288 24947
rect 6328 24915 6360 24947
rect 6400 24915 6432 24947
rect 6472 24915 6504 24947
rect 6544 24915 6576 24947
rect 6616 24915 6648 24947
rect 6688 24915 6720 24947
rect 6760 24915 6792 24947
rect 6832 24915 6864 24947
rect 6904 24915 6936 24947
rect 6976 24915 7008 24947
rect 7048 24915 7080 24947
rect 7120 24915 7152 24947
rect 7192 24915 7224 24947
rect 7264 24915 7296 24947
rect 7336 24915 7368 24947
rect 7408 24915 7440 24947
rect 7480 24915 7512 24947
rect 7552 24915 7584 24947
rect 7624 24915 7656 24947
rect 7696 24915 7728 24947
rect 7768 24915 7800 24947
rect 7840 24915 7872 24947
rect 7912 24915 7944 24947
rect 7984 24915 8016 24947
rect 8056 24915 8088 24947
rect 8128 24915 8160 24947
rect 8200 24915 8232 24947
rect 8272 24915 8304 24947
rect 8344 24915 8376 24947
rect 8416 24915 8448 24947
rect 8488 24915 8520 24947
rect 8560 24915 8592 24947
rect 8632 24915 8664 24947
rect 8704 24915 8736 24947
rect 8776 24915 8808 24947
rect 8848 24915 8880 24947
rect 8920 24915 8952 24947
rect 8992 24915 9024 24947
rect 9064 24915 9096 24947
rect 9136 24915 9168 24947
rect 9208 24915 9240 24947
rect 9280 24915 9312 24947
rect 9352 24915 9384 24947
rect 9424 24915 9456 24947
rect 9496 24915 9528 24947
rect 9568 24915 9600 24947
rect 9640 24915 9672 24947
rect 9712 24915 9744 24947
rect 9784 24915 9816 24947
rect 9856 24915 9888 24947
rect 9928 24915 9960 24947
rect 10000 24915 10032 24947
rect 10072 24915 10104 24947
rect 10144 24915 10176 24947
rect 10216 24915 10248 24947
rect 10288 24915 10320 24947
rect 10360 24915 10392 24947
rect 10432 24915 10464 24947
rect 10504 24915 10536 24947
rect 10576 24915 10608 24947
rect 10648 24915 10680 24947
rect 10720 24915 10752 24947
rect 10792 24915 10824 24947
rect 10864 24915 10896 24947
rect 10936 24915 10968 24947
rect 11008 24915 11040 24947
rect 11080 24915 11112 24947
rect 11152 24915 11184 24947
rect 11224 24915 11256 24947
rect 11296 24915 11328 24947
rect 11368 24915 11400 24947
rect 11440 24915 11472 24947
rect 11512 24915 11544 24947
rect 11584 24915 11616 24947
rect 11656 24915 11688 24947
rect 11728 24915 11760 24947
rect 11800 24915 11832 24947
rect 11872 24915 11904 24947
rect 11944 24915 11976 24947
rect 12016 24915 12048 24947
rect 12088 24915 12120 24947
rect 12160 24915 12192 24947
rect 12232 24915 12264 24947
rect 12304 24915 12336 24947
rect 12376 24915 12408 24947
rect 12448 24915 12480 24947
rect 12520 24915 12552 24947
rect 12592 24915 12624 24947
rect 12664 24915 12696 24947
rect 12736 24915 12768 24947
rect 12808 24915 12840 24947
rect 12880 24915 12912 24947
rect 12952 24915 12984 24947
rect 13024 24915 13056 24947
rect 13096 24915 13128 24947
rect 13168 24915 13200 24947
rect 13240 24915 13272 24947
rect 13312 24915 13344 24947
rect 13384 24915 13416 24947
rect 13456 24915 13488 24947
rect 13528 24915 13560 24947
rect 13600 24915 13632 24947
rect 13672 24915 13704 24947
rect 13744 24915 13776 24947
rect 13816 24915 13848 24947
rect 13888 24915 13920 24947
rect 13960 24915 13992 24947
rect 14032 24915 14064 24947
rect 14104 24915 14136 24947
rect 14176 24915 14208 24947
rect 14248 24915 14280 24947
rect 14320 24915 14352 24947
rect 14392 24915 14424 24947
rect 14464 24915 14496 24947
rect 14536 24915 14568 24947
rect 14608 24915 14640 24947
rect 14680 24915 14712 24947
rect 14752 24915 14784 24947
rect 14824 24915 14856 24947
rect 14896 24915 14928 24947
rect 14968 24915 15000 24947
rect 15040 24915 15072 24947
rect 15112 24915 15144 24947
rect 15184 24915 15216 24947
rect 15256 24915 15288 24947
rect 15328 24915 15360 24947
rect 15400 24915 15432 24947
rect 15472 24915 15504 24947
rect 15544 24915 15576 24947
rect 15616 24915 15648 24947
rect 15688 24915 15720 24947
rect 15760 24915 15792 24947
rect 15832 24915 15864 24947
rect 15904 24915 15936 24947
rect 64 24843 96 24875
rect 136 24843 168 24875
rect 208 24843 240 24875
rect 280 24843 312 24875
rect 352 24843 384 24875
rect 424 24843 456 24875
rect 496 24843 528 24875
rect 568 24843 600 24875
rect 640 24843 672 24875
rect 712 24843 744 24875
rect 784 24843 816 24875
rect 856 24843 888 24875
rect 928 24843 960 24875
rect 1000 24843 1032 24875
rect 1072 24843 1104 24875
rect 1144 24843 1176 24875
rect 1216 24843 1248 24875
rect 1288 24843 1320 24875
rect 1360 24843 1392 24875
rect 1432 24843 1464 24875
rect 1504 24843 1536 24875
rect 1576 24843 1608 24875
rect 1648 24843 1680 24875
rect 1720 24843 1752 24875
rect 1792 24843 1824 24875
rect 1864 24843 1896 24875
rect 1936 24843 1968 24875
rect 2008 24843 2040 24875
rect 2080 24843 2112 24875
rect 2152 24843 2184 24875
rect 2224 24843 2256 24875
rect 2296 24843 2328 24875
rect 2368 24843 2400 24875
rect 2440 24843 2472 24875
rect 2512 24843 2544 24875
rect 2584 24843 2616 24875
rect 2656 24843 2688 24875
rect 2728 24843 2760 24875
rect 2800 24843 2832 24875
rect 2872 24843 2904 24875
rect 2944 24843 2976 24875
rect 3016 24843 3048 24875
rect 3088 24843 3120 24875
rect 3160 24843 3192 24875
rect 3232 24843 3264 24875
rect 3304 24843 3336 24875
rect 3376 24843 3408 24875
rect 3448 24843 3480 24875
rect 3520 24843 3552 24875
rect 3592 24843 3624 24875
rect 3664 24843 3696 24875
rect 3736 24843 3768 24875
rect 3808 24843 3840 24875
rect 3880 24843 3912 24875
rect 3952 24843 3984 24875
rect 4024 24843 4056 24875
rect 4096 24843 4128 24875
rect 4168 24843 4200 24875
rect 4240 24843 4272 24875
rect 4312 24843 4344 24875
rect 4384 24843 4416 24875
rect 4456 24843 4488 24875
rect 4528 24843 4560 24875
rect 4600 24843 4632 24875
rect 4672 24843 4704 24875
rect 4744 24843 4776 24875
rect 4816 24843 4848 24875
rect 4888 24843 4920 24875
rect 4960 24843 4992 24875
rect 5032 24843 5064 24875
rect 5104 24843 5136 24875
rect 5176 24843 5208 24875
rect 5248 24843 5280 24875
rect 5320 24843 5352 24875
rect 5392 24843 5424 24875
rect 5464 24843 5496 24875
rect 5536 24843 5568 24875
rect 5608 24843 5640 24875
rect 5680 24843 5712 24875
rect 5752 24843 5784 24875
rect 5824 24843 5856 24875
rect 5896 24843 5928 24875
rect 5968 24843 6000 24875
rect 6040 24843 6072 24875
rect 6112 24843 6144 24875
rect 6184 24843 6216 24875
rect 6256 24843 6288 24875
rect 6328 24843 6360 24875
rect 6400 24843 6432 24875
rect 6472 24843 6504 24875
rect 6544 24843 6576 24875
rect 6616 24843 6648 24875
rect 6688 24843 6720 24875
rect 6760 24843 6792 24875
rect 6832 24843 6864 24875
rect 6904 24843 6936 24875
rect 6976 24843 7008 24875
rect 7048 24843 7080 24875
rect 7120 24843 7152 24875
rect 7192 24843 7224 24875
rect 7264 24843 7296 24875
rect 7336 24843 7368 24875
rect 7408 24843 7440 24875
rect 7480 24843 7512 24875
rect 7552 24843 7584 24875
rect 7624 24843 7656 24875
rect 7696 24843 7728 24875
rect 7768 24843 7800 24875
rect 7840 24843 7872 24875
rect 7912 24843 7944 24875
rect 7984 24843 8016 24875
rect 8056 24843 8088 24875
rect 8128 24843 8160 24875
rect 8200 24843 8232 24875
rect 8272 24843 8304 24875
rect 8344 24843 8376 24875
rect 8416 24843 8448 24875
rect 8488 24843 8520 24875
rect 8560 24843 8592 24875
rect 8632 24843 8664 24875
rect 8704 24843 8736 24875
rect 8776 24843 8808 24875
rect 8848 24843 8880 24875
rect 8920 24843 8952 24875
rect 8992 24843 9024 24875
rect 9064 24843 9096 24875
rect 9136 24843 9168 24875
rect 9208 24843 9240 24875
rect 9280 24843 9312 24875
rect 9352 24843 9384 24875
rect 9424 24843 9456 24875
rect 9496 24843 9528 24875
rect 9568 24843 9600 24875
rect 9640 24843 9672 24875
rect 9712 24843 9744 24875
rect 9784 24843 9816 24875
rect 9856 24843 9888 24875
rect 9928 24843 9960 24875
rect 10000 24843 10032 24875
rect 10072 24843 10104 24875
rect 10144 24843 10176 24875
rect 10216 24843 10248 24875
rect 10288 24843 10320 24875
rect 10360 24843 10392 24875
rect 10432 24843 10464 24875
rect 10504 24843 10536 24875
rect 10576 24843 10608 24875
rect 10648 24843 10680 24875
rect 10720 24843 10752 24875
rect 10792 24843 10824 24875
rect 10864 24843 10896 24875
rect 10936 24843 10968 24875
rect 11008 24843 11040 24875
rect 11080 24843 11112 24875
rect 11152 24843 11184 24875
rect 11224 24843 11256 24875
rect 11296 24843 11328 24875
rect 11368 24843 11400 24875
rect 11440 24843 11472 24875
rect 11512 24843 11544 24875
rect 11584 24843 11616 24875
rect 11656 24843 11688 24875
rect 11728 24843 11760 24875
rect 11800 24843 11832 24875
rect 11872 24843 11904 24875
rect 11944 24843 11976 24875
rect 12016 24843 12048 24875
rect 12088 24843 12120 24875
rect 12160 24843 12192 24875
rect 12232 24843 12264 24875
rect 12304 24843 12336 24875
rect 12376 24843 12408 24875
rect 12448 24843 12480 24875
rect 12520 24843 12552 24875
rect 12592 24843 12624 24875
rect 12664 24843 12696 24875
rect 12736 24843 12768 24875
rect 12808 24843 12840 24875
rect 12880 24843 12912 24875
rect 12952 24843 12984 24875
rect 13024 24843 13056 24875
rect 13096 24843 13128 24875
rect 13168 24843 13200 24875
rect 13240 24843 13272 24875
rect 13312 24843 13344 24875
rect 13384 24843 13416 24875
rect 13456 24843 13488 24875
rect 13528 24843 13560 24875
rect 13600 24843 13632 24875
rect 13672 24843 13704 24875
rect 13744 24843 13776 24875
rect 13816 24843 13848 24875
rect 13888 24843 13920 24875
rect 13960 24843 13992 24875
rect 14032 24843 14064 24875
rect 14104 24843 14136 24875
rect 14176 24843 14208 24875
rect 14248 24843 14280 24875
rect 14320 24843 14352 24875
rect 14392 24843 14424 24875
rect 14464 24843 14496 24875
rect 14536 24843 14568 24875
rect 14608 24843 14640 24875
rect 14680 24843 14712 24875
rect 14752 24843 14784 24875
rect 14824 24843 14856 24875
rect 14896 24843 14928 24875
rect 14968 24843 15000 24875
rect 15040 24843 15072 24875
rect 15112 24843 15144 24875
rect 15184 24843 15216 24875
rect 15256 24843 15288 24875
rect 15328 24843 15360 24875
rect 15400 24843 15432 24875
rect 15472 24843 15504 24875
rect 15544 24843 15576 24875
rect 15616 24843 15648 24875
rect 15688 24843 15720 24875
rect 15760 24843 15792 24875
rect 15832 24843 15864 24875
rect 15904 24843 15936 24875
rect 64 24771 96 24803
rect 136 24771 168 24803
rect 208 24771 240 24803
rect 280 24771 312 24803
rect 352 24771 384 24803
rect 424 24771 456 24803
rect 496 24771 528 24803
rect 568 24771 600 24803
rect 640 24771 672 24803
rect 712 24771 744 24803
rect 784 24771 816 24803
rect 856 24771 888 24803
rect 928 24771 960 24803
rect 1000 24771 1032 24803
rect 1072 24771 1104 24803
rect 1144 24771 1176 24803
rect 1216 24771 1248 24803
rect 1288 24771 1320 24803
rect 1360 24771 1392 24803
rect 1432 24771 1464 24803
rect 1504 24771 1536 24803
rect 1576 24771 1608 24803
rect 1648 24771 1680 24803
rect 1720 24771 1752 24803
rect 1792 24771 1824 24803
rect 1864 24771 1896 24803
rect 1936 24771 1968 24803
rect 2008 24771 2040 24803
rect 2080 24771 2112 24803
rect 2152 24771 2184 24803
rect 2224 24771 2256 24803
rect 2296 24771 2328 24803
rect 2368 24771 2400 24803
rect 2440 24771 2472 24803
rect 2512 24771 2544 24803
rect 2584 24771 2616 24803
rect 2656 24771 2688 24803
rect 2728 24771 2760 24803
rect 2800 24771 2832 24803
rect 2872 24771 2904 24803
rect 2944 24771 2976 24803
rect 3016 24771 3048 24803
rect 3088 24771 3120 24803
rect 3160 24771 3192 24803
rect 3232 24771 3264 24803
rect 3304 24771 3336 24803
rect 3376 24771 3408 24803
rect 3448 24771 3480 24803
rect 3520 24771 3552 24803
rect 3592 24771 3624 24803
rect 3664 24771 3696 24803
rect 3736 24771 3768 24803
rect 3808 24771 3840 24803
rect 3880 24771 3912 24803
rect 3952 24771 3984 24803
rect 4024 24771 4056 24803
rect 4096 24771 4128 24803
rect 4168 24771 4200 24803
rect 4240 24771 4272 24803
rect 4312 24771 4344 24803
rect 4384 24771 4416 24803
rect 4456 24771 4488 24803
rect 4528 24771 4560 24803
rect 4600 24771 4632 24803
rect 4672 24771 4704 24803
rect 4744 24771 4776 24803
rect 4816 24771 4848 24803
rect 4888 24771 4920 24803
rect 4960 24771 4992 24803
rect 5032 24771 5064 24803
rect 5104 24771 5136 24803
rect 5176 24771 5208 24803
rect 5248 24771 5280 24803
rect 5320 24771 5352 24803
rect 5392 24771 5424 24803
rect 5464 24771 5496 24803
rect 5536 24771 5568 24803
rect 5608 24771 5640 24803
rect 5680 24771 5712 24803
rect 5752 24771 5784 24803
rect 5824 24771 5856 24803
rect 5896 24771 5928 24803
rect 5968 24771 6000 24803
rect 6040 24771 6072 24803
rect 6112 24771 6144 24803
rect 6184 24771 6216 24803
rect 6256 24771 6288 24803
rect 6328 24771 6360 24803
rect 6400 24771 6432 24803
rect 6472 24771 6504 24803
rect 6544 24771 6576 24803
rect 6616 24771 6648 24803
rect 6688 24771 6720 24803
rect 6760 24771 6792 24803
rect 6832 24771 6864 24803
rect 6904 24771 6936 24803
rect 6976 24771 7008 24803
rect 7048 24771 7080 24803
rect 7120 24771 7152 24803
rect 7192 24771 7224 24803
rect 7264 24771 7296 24803
rect 7336 24771 7368 24803
rect 7408 24771 7440 24803
rect 7480 24771 7512 24803
rect 7552 24771 7584 24803
rect 7624 24771 7656 24803
rect 7696 24771 7728 24803
rect 7768 24771 7800 24803
rect 7840 24771 7872 24803
rect 7912 24771 7944 24803
rect 7984 24771 8016 24803
rect 8056 24771 8088 24803
rect 8128 24771 8160 24803
rect 8200 24771 8232 24803
rect 8272 24771 8304 24803
rect 8344 24771 8376 24803
rect 8416 24771 8448 24803
rect 8488 24771 8520 24803
rect 8560 24771 8592 24803
rect 8632 24771 8664 24803
rect 8704 24771 8736 24803
rect 8776 24771 8808 24803
rect 8848 24771 8880 24803
rect 8920 24771 8952 24803
rect 8992 24771 9024 24803
rect 9064 24771 9096 24803
rect 9136 24771 9168 24803
rect 9208 24771 9240 24803
rect 9280 24771 9312 24803
rect 9352 24771 9384 24803
rect 9424 24771 9456 24803
rect 9496 24771 9528 24803
rect 9568 24771 9600 24803
rect 9640 24771 9672 24803
rect 9712 24771 9744 24803
rect 9784 24771 9816 24803
rect 9856 24771 9888 24803
rect 9928 24771 9960 24803
rect 10000 24771 10032 24803
rect 10072 24771 10104 24803
rect 10144 24771 10176 24803
rect 10216 24771 10248 24803
rect 10288 24771 10320 24803
rect 10360 24771 10392 24803
rect 10432 24771 10464 24803
rect 10504 24771 10536 24803
rect 10576 24771 10608 24803
rect 10648 24771 10680 24803
rect 10720 24771 10752 24803
rect 10792 24771 10824 24803
rect 10864 24771 10896 24803
rect 10936 24771 10968 24803
rect 11008 24771 11040 24803
rect 11080 24771 11112 24803
rect 11152 24771 11184 24803
rect 11224 24771 11256 24803
rect 11296 24771 11328 24803
rect 11368 24771 11400 24803
rect 11440 24771 11472 24803
rect 11512 24771 11544 24803
rect 11584 24771 11616 24803
rect 11656 24771 11688 24803
rect 11728 24771 11760 24803
rect 11800 24771 11832 24803
rect 11872 24771 11904 24803
rect 11944 24771 11976 24803
rect 12016 24771 12048 24803
rect 12088 24771 12120 24803
rect 12160 24771 12192 24803
rect 12232 24771 12264 24803
rect 12304 24771 12336 24803
rect 12376 24771 12408 24803
rect 12448 24771 12480 24803
rect 12520 24771 12552 24803
rect 12592 24771 12624 24803
rect 12664 24771 12696 24803
rect 12736 24771 12768 24803
rect 12808 24771 12840 24803
rect 12880 24771 12912 24803
rect 12952 24771 12984 24803
rect 13024 24771 13056 24803
rect 13096 24771 13128 24803
rect 13168 24771 13200 24803
rect 13240 24771 13272 24803
rect 13312 24771 13344 24803
rect 13384 24771 13416 24803
rect 13456 24771 13488 24803
rect 13528 24771 13560 24803
rect 13600 24771 13632 24803
rect 13672 24771 13704 24803
rect 13744 24771 13776 24803
rect 13816 24771 13848 24803
rect 13888 24771 13920 24803
rect 13960 24771 13992 24803
rect 14032 24771 14064 24803
rect 14104 24771 14136 24803
rect 14176 24771 14208 24803
rect 14248 24771 14280 24803
rect 14320 24771 14352 24803
rect 14392 24771 14424 24803
rect 14464 24771 14496 24803
rect 14536 24771 14568 24803
rect 14608 24771 14640 24803
rect 14680 24771 14712 24803
rect 14752 24771 14784 24803
rect 14824 24771 14856 24803
rect 14896 24771 14928 24803
rect 14968 24771 15000 24803
rect 15040 24771 15072 24803
rect 15112 24771 15144 24803
rect 15184 24771 15216 24803
rect 15256 24771 15288 24803
rect 15328 24771 15360 24803
rect 15400 24771 15432 24803
rect 15472 24771 15504 24803
rect 15544 24771 15576 24803
rect 15616 24771 15648 24803
rect 15688 24771 15720 24803
rect 15760 24771 15792 24803
rect 15832 24771 15864 24803
rect 15904 24771 15936 24803
rect 64 24699 96 24731
rect 136 24699 168 24731
rect 208 24699 240 24731
rect 280 24699 312 24731
rect 352 24699 384 24731
rect 424 24699 456 24731
rect 496 24699 528 24731
rect 568 24699 600 24731
rect 640 24699 672 24731
rect 712 24699 744 24731
rect 784 24699 816 24731
rect 856 24699 888 24731
rect 928 24699 960 24731
rect 1000 24699 1032 24731
rect 1072 24699 1104 24731
rect 1144 24699 1176 24731
rect 1216 24699 1248 24731
rect 1288 24699 1320 24731
rect 1360 24699 1392 24731
rect 1432 24699 1464 24731
rect 1504 24699 1536 24731
rect 1576 24699 1608 24731
rect 1648 24699 1680 24731
rect 1720 24699 1752 24731
rect 1792 24699 1824 24731
rect 1864 24699 1896 24731
rect 1936 24699 1968 24731
rect 2008 24699 2040 24731
rect 2080 24699 2112 24731
rect 2152 24699 2184 24731
rect 2224 24699 2256 24731
rect 2296 24699 2328 24731
rect 2368 24699 2400 24731
rect 2440 24699 2472 24731
rect 2512 24699 2544 24731
rect 2584 24699 2616 24731
rect 2656 24699 2688 24731
rect 2728 24699 2760 24731
rect 2800 24699 2832 24731
rect 2872 24699 2904 24731
rect 2944 24699 2976 24731
rect 3016 24699 3048 24731
rect 3088 24699 3120 24731
rect 3160 24699 3192 24731
rect 3232 24699 3264 24731
rect 3304 24699 3336 24731
rect 3376 24699 3408 24731
rect 3448 24699 3480 24731
rect 3520 24699 3552 24731
rect 3592 24699 3624 24731
rect 3664 24699 3696 24731
rect 3736 24699 3768 24731
rect 3808 24699 3840 24731
rect 3880 24699 3912 24731
rect 3952 24699 3984 24731
rect 4024 24699 4056 24731
rect 4096 24699 4128 24731
rect 4168 24699 4200 24731
rect 4240 24699 4272 24731
rect 4312 24699 4344 24731
rect 4384 24699 4416 24731
rect 4456 24699 4488 24731
rect 4528 24699 4560 24731
rect 4600 24699 4632 24731
rect 4672 24699 4704 24731
rect 4744 24699 4776 24731
rect 4816 24699 4848 24731
rect 4888 24699 4920 24731
rect 4960 24699 4992 24731
rect 5032 24699 5064 24731
rect 5104 24699 5136 24731
rect 5176 24699 5208 24731
rect 5248 24699 5280 24731
rect 5320 24699 5352 24731
rect 5392 24699 5424 24731
rect 5464 24699 5496 24731
rect 5536 24699 5568 24731
rect 5608 24699 5640 24731
rect 5680 24699 5712 24731
rect 5752 24699 5784 24731
rect 5824 24699 5856 24731
rect 5896 24699 5928 24731
rect 5968 24699 6000 24731
rect 6040 24699 6072 24731
rect 6112 24699 6144 24731
rect 6184 24699 6216 24731
rect 6256 24699 6288 24731
rect 6328 24699 6360 24731
rect 6400 24699 6432 24731
rect 6472 24699 6504 24731
rect 6544 24699 6576 24731
rect 6616 24699 6648 24731
rect 6688 24699 6720 24731
rect 6760 24699 6792 24731
rect 6832 24699 6864 24731
rect 6904 24699 6936 24731
rect 6976 24699 7008 24731
rect 7048 24699 7080 24731
rect 7120 24699 7152 24731
rect 7192 24699 7224 24731
rect 7264 24699 7296 24731
rect 7336 24699 7368 24731
rect 7408 24699 7440 24731
rect 7480 24699 7512 24731
rect 7552 24699 7584 24731
rect 7624 24699 7656 24731
rect 7696 24699 7728 24731
rect 7768 24699 7800 24731
rect 7840 24699 7872 24731
rect 7912 24699 7944 24731
rect 7984 24699 8016 24731
rect 8056 24699 8088 24731
rect 8128 24699 8160 24731
rect 8200 24699 8232 24731
rect 8272 24699 8304 24731
rect 8344 24699 8376 24731
rect 8416 24699 8448 24731
rect 8488 24699 8520 24731
rect 8560 24699 8592 24731
rect 8632 24699 8664 24731
rect 8704 24699 8736 24731
rect 8776 24699 8808 24731
rect 8848 24699 8880 24731
rect 8920 24699 8952 24731
rect 8992 24699 9024 24731
rect 9064 24699 9096 24731
rect 9136 24699 9168 24731
rect 9208 24699 9240 24731
rect 9280 24699 9312 24731
rect 9352 24699 9384 24731
rect 9424 24699 9456 24731
rect 9496 24699 9528 24731
rect 9568 24699 9600 24731
rect 9640 24699 9672 24731
rect 9712 24699 9744 24731
rect 9784 24699 9816 24731
rect 9856 24699 9888 24731
rect 9928 24699 9960 24731
rect 10000 24699 10032 24731
rect 10072 24699 10104 24731
rect 10144 24699 10176 24731
rect 10216 24699 10248 24731
rect 10288 24699 10320 24731
rect 10360 24699 10392 24731
rect 10432 24699 10464 24731
rect 10504 24699 10536 24731
rect 10576 24699 10608 24731
rect 10648 24699 10680 24731
rect 10720 24699 10752 24731
rect 10792 24699 10824 24731
rect 10864 24699 10896 24731
rect 10936 24699 10968 24731
rect 11008 24699 11040 24731
rect 11080 24699 11112 24731
rect 11152 24699 11184 24731
rect 11224 24699 11256 24731
rect 11296 24699 11328 24731
rect 11368 24699 11400 24731
rect 11440 24699 11472 24731
rect 11512 24699 11544 24731
rect 11584 24699 11616 24731
rect 11656 24699 11688 24731
rect 11728 24699 11760 24731
rect 11800 24699 11832 24731
rect 11872 24699 11904 24731
rect 11944 24699 11976 24731
rect 12016 24699 12048 24731
rect 12088 24699 12120 24731
rect 12160 24699 12192 24731
rect 12232 24699 12264 24731
rect 12304 24699 12336 24731
rect 12376 24699 12408 24731
rect 12448 24699 12480 24731
rect 12520 24699 12552 24731
rect 12592 24699 12624 24731
rect 12664 24699 12696 24731
rect 12736 24699 12768 24731
rect 12808 24699 12840 24731
rect 12880 24699 12912 24731
rect 12952 24699 12984 24731
rect 13024 24699 13056 24731
rect 13096 24699 13128 24731
rect 13168 24699 13200 24731
rect 13240 24699 13272 24731
rect 13312 24699 13344 24731
rect 13384 24699 13416 24731
rect 13456 24699 13488 24731
rect 13528 24699 13560 24731
rect 13600 24699 13632 24731
rect 13672 24699 13704 24731
rect 13744 24699 13776 24731
rect 13816 24699 13848 24731
rect 13888 24699 13920 24731
rect 13960 24699 13992 24731
rect 14032 24699 14064 24731
rect 14104 24699 14136 24731
rect 14176 24699 14208 24731
rect 14248 24699 14280 24731
rect 14320 24699 14352 24731
rect 14392 24699 14424 24731
rect 14464 24699 14496 24731
rect 14536 24699 14568 24731
rect 14608 24699 14640 24731
rect 14680 24699 14712 24731
rect 14752 24699 14784 24731
rect 14824 24699 14856 24731
rect 14896 24699 14928 24731
rect 14968 24699 15000 24731
rect 15040 24699 15072 24731
rect 15112 24699 15144 24731
rect 15184 24699 15216 24731
rect 15256 24699 15288 24731
rect 15328 24699 15360 24731
rect 15400 24699 15432 24731
rect 15472 24699 15504 24731
rect 15544 24699 15576 24731
rect 15616 24699 15648 24731
rect 15688 24699 15720 24731
rect 15760 24699 15792 24731
rect 15832 24699 15864 24731
rect 15904 24699 15936 24731
rect 64 24627 96 24659
rect 136 24627 168 24659
rect 208 24627 240 24659
rect 280 24627 312 24659
rect 352 24627 384 24659
rect 424 24627 456 24659
rect 496 24627 528 24659
rect 568 24627 600 24659
rect 640 24627 672 24659
rect 712 24627 744 24659
rect 784 24627 816 24659
rect 856 24627 888 24659
rect 928 24627 960 24659
rect 1000 24627 1032 24659
rect 1072 24627 1104 24659
rect 1144 24627 1176 24659
rect 1216 24627 1248 24659
rect 1288 24627 1320 24659
rect 1360 24627 1392 24659
rect 1432 24627 1464 24659
rect 1504 24627 1536 24659
rect 1576 24627 1608 24659
rect 1648 24627 1680 24659
rect 1720 24627 1752 24659
rect 1792 24627 1824 24659
rect 1864 24627 1896 24659
rect 1936 24627 1968 24659
rect 2008 24627 2040 24659
rect 2080 24627 2112 24659
rect 2152 24627 2184 24659
rect 2224 24627 2256 24659
rect 2296 24627 2328 24659
rect 2368 24627 2400 24659
rect 2440 24627 2472 24659
rect 2512 24627 2544 24659
rect 2584 24627 2616 24659
rect 2656 24627 2688 24659
rect 2728 24627 2760 24659
rect 2800 24627 2832 24659
rect 2872 24627 2904 24659
rect 2944 24627 2976 24659
rect 3016 24627 3048 24659
rect 3088 24627 3120 24659
rect 3160 24627 3192 24659
rect 3232 24627 3264 24659
rect 3304 24627 3336 24659
rect 3376 24627 3408 24659
rect 3448 24627 3480 24659
rect 3520 24627 3552 24659
rect 3592 24627 3624 24659
rect 3664 24627 3696 24659
rect 3736 24627 3768 24659
rect 3808 24627 3840 24659
rect 3880 24627 3912 24659
rect 3952 24627 3984 24659
rect 4024 24627 4056 24659
rect 4096 24627 4128 24659
rect 4168 24627 4200 24659
rect 4240 24627 4272 24659
rect 4312 24627 4344 24659
rect 4384 24627 4416 24659
rect 4456 24627 4488 24659
rect 4528 24627 4560 24659
rect 4600 24627 4632 24659
rect 4672 24627 4704 24659
rect 4744 24627 4776 24659
rect 4816 24627 4848 24659
rect 4888 24627 4920 24659
rect 4960 24627 4992 24659
rect 5032 24627 5064 24659
rect 5104 24627 5136 24659
rect 5176 24627 5208 24659
rect 5248 24627 5280 24659
rect 5320 24627 5352 24659
rect 5392 24627 5424 24659
rect 5464 24627 5496 24659
rect 5536 24627 5568 24659
rect 5608 24627 5640 24659
rect 5680 24627 5712 24659
rect 5752 24627 5784 24659
rect 5824 24627 5856 24659
rect 5896 24627 5928 24659
rect 5968 24627 6000 24659
rect 6040 24627 6072 24659
rect 6112 24627 6144 24659
rect 6184 24627 6216 24659
rect 6256 24627 6288 24659
rect 6328 24627 6360 24659
rect 6400 24627 6432 24659
rect 6472 24627 6504 24659
rect 6544 24627 6576 24659
rect 6616 24627 6648 24659
rect 6688 24627 6720 24659
rect 6760 24627 6792 24659
rect 6832 24627 6864 24659
rect 6904 24627 6936 24659
rect 6976 24627 7008 24659
rect 7048 24627 7080 24659
rect 7120 24627 7152 24659
rect 7192 24627 7224 24659
rect 7264 24627 7296 24659
rect 7336 24627 7368 24659
rect 7408 24627 7440 24659
rect 7480 24627 7512 24659
rect 7552 24627 7584 24659
rect 7624 24627 7656 24659
rect 7696 24627 7728 24659
rect 7768 24627 7800 24659
rect 7840 24627 7872 24659
rect 7912 24627 7944 24659
rect 7984 24627 8016 24659
rect 8056 24627 8088 24659
rect 8128 24627 8160 24659
rect 8200 24627 8232 24659
rect 8272 24627 8304 24659
rect 8344 24627 8376 24659
rect 8416 24627 8448 24659
rect 8488 24627 8520 24659
rect 8560 24627 8592 24659
rect 8632 24627 8664 24659
rect 8704 24627 8736 24659
rect 8776 24627 8808 24659
rect 8848 24627 8880 24659
rect 8920 24627 8952 24659
rect 8992 24627 9024 24659
rect 9064 24627 9096 24659
rect 9136 24627 9168 24659
rect 9208 24627 9240 24659
rect 9280 24627 9312 24659
rect 9352 24627 9384 24659
rect 9424 24627 9456 24659
rect 9496 24627 9528 24659
rect 9568 24627 9600 24659
rect 9640 24627 9672 24659
rect 9712 24627 9744 24659
rect 9784 24627 9816 24659
rect 9856 24627 9888 24659
rect 9928 24627 9960 24659
rect 10000 24627 10032 24659
rect 10072 24627 10104 24659
rect 10144 24627 10176 24659
rect 10216 24627 10248 24659
rect 10288 24627 10320 24659
rect 10360 24627 10392 24659
rect 10432 24627 10464 24659
rect 10504 24627 10536 24659
rect 10576 24627 10608 24659
rect 10648 24627 10680 24659
rect 10720 24627 10752 24659
rect 10792 24627 10824 24659
rect 10864 24627 10896 24659
rect 10936 24627 10968 24659
rect 11008 24627 11040 24659
rect 11080 24627 11112 24659
rect 11152 24627 11184 24659
rect 11224 24627 11256 24659
rect 11296 24627 11328 24659
rect 11368 24627 11400 24659
rect 11440 24627 11472 24659
rect 11512 24627 11544 24659
rect 11584 24627 11616 24659
rect 11656 24627 11688 24659
rect 11728 24627 11760 24659
rect 11800 24627 11832 24659
rect 11872 24627 11904 24659
rect 11944 24627 11976 24659
rect 12016 24627 12048 24659
rect 12088 24627 12120 24659
rect 12160 24627 12192 24659
rect 12232 24627 12264 24659
rect 12304 24627 12336 24659
rect 12376 24627 12408 24659
rect 12448 24627 12480 24659
rect 12520 24627 12552 24659
rect 12592 24627 12624 24659
rect 12664 24627 12696 24659
rect 12736 24627 12768 24659
rect 12808 24627 12840 24659
rect 12880 24627 12912 24659
rect 12952 24627 12984 24659
rect 13024 24627 13056 24659
rect 13096 24627 13128 24659
rect 13168 24627 13200 24659
rect 13240 24627 13272 24659
rect 13312 24627 13344 24659
rect 13384 24627 13416 24659
rect 13456 24627 13488 24659
rect 13528 24627 13560 24659
rect 13600 24627 13632 24659
rect 13672 24627 13704 24659
rect 13744 24627 13776 24659
rect 13816 24627 13848 24659
rect 13888 24627 13920 24659
rect 13960 24627 13992 24659
rect 14032 24627 14064 24659
rect 14104 24627 14136 24659
rect 14176 24627 14208 24659
rect 14248 24627 14280 24659
rect 14320 24627 14352 24659
rect 14392 24627 14424 24659
rect 14464 24627 14496 24659
rect 14536 24627 14568 24659
rect 14608 24627 14640 24659
rect 14680 24627 14712 24659
rect 14752 24627 14784 24659
rect 14824 24627 14856 24659
rect 14896 24627 14928 24659
rect 14968 24627 15000 24659
rect 15040 24627 15072 24659
rect 15112 24627 15144 24659
rect 15184 24627 15216 24659
rect 15256 24627 15288 24659
rect 15328 24627 15360 24659
rect 15400 24627 15432 24659
rect 15472 24627 15504 24659
rect 15544 24627 15576 24659
rect 15616 24627 15648 24659
rect 15688 24627 15720 24659
rect 15760 24627 15792 24659
rect 15832 24627 15864 24659
rect 15904 24627 15936 24659
rect 64 24555 96 24587
rect 136 24555 168 24587
rect 208 24555 240 24587
rect 280 24555 312 24587
rect 352 24555 384 24587
rect 424 24555 456 24587
rect 496 24555 528 24587
rect 568 24555 600 24587
rect 640 24555 672 24587
rect 712 24555 744 24587
rect 784 24555 816 24587
rect 856 24555 888 24587
rect 928 24555 960 24587
rect 1000 24555 1032 24587
rect 1072 24555 1104 24587
rect 1144 24555 1176 24587
rect 1216 24555 1248 24587
rect 1288 24555 1320 24587
rect 1360 24555 1392 24587
rect 1432 24555 1464 24587
rect 1504 24555 1536 24587
rect 1576 24555 1608 24587
rect 1648 24555 1680 24587
rect 1720 24555 1752 24587
rect 1792 24555 1824 24587
rect 1864 24555 1896 24587
rect 1936 24555 1968 24587
rect 2008 24555 2040 24587
rect 2080 24555 2112 24587
rect 2152 24555 2184 24587
rect 2224 24555 2256 24587
rect 2296 24555 2328 24587
rect 2368 24555 2400 24587
rect 2440 24555 2472 24587
rect 2512 24555 2544 24587
rect 2584 24555 2616 24587
rect 2656 24555 2688 24587
rect 2728 24555 2760 24587
rect 2800 24555 2832 24587
rect 2872 24555 2904 24587
rect 2944 24555 2976 24587
rect 3016 24555 3048 24587
rect 3088 24555 3120 24587
rect 3160 24555 3192 24587
rect 3232 24555 3264 24587
rect 3304 24555 3336 24587
rect 3376 24555 3408 24587
rect 3448 24555 3480 24587
rect 3520 24555 3552 24587
rect 3592 24555 3624 24587
rect 3664 24555 3696 24587
rect 3736 24555 3768 24587
rect 3808 24555 3840 24587
rect 3880 24555 3912 24587
rect 3952 24555 3984 24587
rect 4024 24555 4056 24587
rect 4096 24555 4128 24587
rect 4168 24555 4200 24587
rect 4240 24555 4272 24587
rect 4312 24555 4344 24587
rect 4384 24555 4416 24587
rect 4456 24555 4488 24587
rect 4528 24555 4560 24587
rect 4600 24555 4632 24587
rect 4672 24555 4704 24587
rect 4744 24555 4776 24587
rect 4816 24555 4848 24587
rect 4888 24555 4920 24587
rect 4960 24555 4992 24587
rect 5032 24555 5064 24587
rect 5104 24555 5136 24587
rect 5176 24555 5208 24587
rect 5248 24555 5280 24587
rect 5320 24555 5352 24587
rect 5392 24555 5424 24587
rect 5464 24555 5496 24587
rect 5536 24555 5568 24587
rect 5608 24555 5640 24587
rect 5680 24555 5712 24587
rect 5752 24555 5784 24587
rect 5824 24555 5856 24587
rect 5896 24555 5928 24587
rect 5968 24555 6000 24587
rect 6040 24555 6072 24587
rect 6112 24555 6144 24587
rect 6184 24555 6216 24587
rect 6256 24555 6288 24587
rect 6328 24555 6360 24587
rect 6400 24555 6432 24587
rect 6472 24555 6504 24587
rect 6544 24555 6576 24587
rect 6616 24555 6648 24587
rect 6688 24555 6720 24587
rect 6760 24555 6792 24587
rect 6832 24555 6864 24587
rect 6904 24555 6936 24587
rect 6976 24555 7008 24587
rect 7048 24555 7080 24587
rect 7120 24555 7152 24587
rect 7192 24555 7224 24587
rect 7264 24555 7296 24587
rect 7336 24555 7368 24587
rect 7408 24555 7440 24587
rect 7480 24555 7512 24587
rect 7552 24555 7584 24587
rect 7624 24555 7656 24587
rect 7696 24555 7728 24587
rect 7768 24555 7800 24587
rect 7840 24555 7872 24587
rect 7912 24555 7944 24587
rect 7984 24555 8016 24587
rect 8056 24555 8088 24587
rect 8128 24555 8160 24587
rect 8200 24555 8232 24587
rect 8272 24555 8304 24587
rect 8344 24555 8376 24587
rect 8416 24555 8448 24587
rect 8488 24555 8520 24587
rect 8560 24555 8592 24587
rect 8632 24555 8664 24587
rect 8704 24555 8736 24587
rect 8776 24555 8808 24587
rect 8848 24555 8880 24587
rect 8920 24555 8952 24587
rect 8992 24555 9024 24587
rect 9064 24555 9096 24587
rect 9136 24555 9168 24587
rect 9208 24555 9240 24587
rect 9280 24555 9312 24587
rect 9352 24555 9384 24587
rect 9424 24555 9456 24587
rect 9496 24555 9528 24587
rect 9568 24555 9600 24587
rect 9640 24555 9672 24587
rect 9712 24555 9744 24587
rect 9784 24555 9816 24587
rect 9856 24555 9888 24587
rect 9928 24555 9960 24587
rect 10000 24555 10032 24587
rect 10072 24555 10104 24587
rect 10144 24555 10176 24587
rect 10216 24555 10248 24587
rect 10288 24555 10320 24587
rect 10360 24555 10392 24587
rect 10432 24555 10464 24587
rect 10504 24555 10536 24587
rect 10576 24555 10608 24587
rect 10648 24555 10680 24587
rect 10720 24555 10752 24587
rect 10792 24555 10824 24587
rect 10864 24555 10896 24587
rect 10936 24555 10968 24587
rect 11008 24555 11040 24587
rect 11080 24555 11112 24587
rect 11152 24555 11184 24587
rect 11224 24555 11256 24587
rect 11296 24555 11328 24587
rect 11368 24555 11400 24587
rect 11440 24555 11472 24587
rect 11512 24555 11544 24587
rect 11584 24555 11616 24587
rect 11656 24555 11688 24587
rect 11728 24555 11760 24587
rect 11800 24555 11832 24587
rect 11872 24555 11904 24587
rect 11944 24555 11976 24587
rect 12016 24555 12048 24587
rect 12088 24555 12120 24587
rect 12160 24555 12192 24587
rect 12232 24555 12264 24587
rect 12304 24555 12336 24587
rect 12376 24555 12408 24587
rect 12448 24555 12480 24587
rect 12520 24555 12552 24587
rect 12592 24555 12624 24587
rect 12664 24555 12696 24587
rect 12736 24555 12768 24587
rect 12808 24555 12840 24587
rect 12880 24555 12912 24587
rect 12952 24555 12984 24587
rect 13024 24555 13056 24587
rect 13096 24555 13128 24587
rect 13168 24555 13200 24587
rect 13240 24555 13272 24587
rect 13312 24555 13344 24587
rect 13384 24555 13416 24587
rect 13456 24555 13488 24587
rect 13528 24555 13560 24587
rect 13600 24555 13632 24587
rect 13672 24555 13704 24587
rect 13744 24555 13776 24587
rect 13816 24555 13848 24587
rect 13888 24555 13920 24587
rect 13960 24555 13992 24587
rect 14032 24555 14064 24587
rect 14104 24555 14136 24587
rect 14176 24555 14208 24587
rect 14248 24555 14280 24587
rect 14320 24555 14352 24587
rect 14392 24555 14424 24587
rect 14464 24555 14496 24587
rect 14536 24555 14568 24587
rect 14608 24555 14640 24587
rect 14680 24555 14712 24587
rect 14752 24555 14784 24587
rect 14824 24555 14856 24587
rect 14896 24555 14928 24587
rect 14968 24555 15000 24587
rect 15040 24555 15072 24587
rect 15112 24555 15144 24587
rect 15184 24555 15216 24587
rect 15256 24555 15288 24587
rect 15328 24555 15360 24587
rect 15400 24555 15432 24587
rect 15472 24555 15504 24587
rect 15544 24555 15576 24587
rect 15616 24555 15648 24587
rect 15688 24555 15720 24587
rect 15760 24555 15792 24587
rect 15832 24555 15864 24587
rect 15904 24555 15936 24587
rect 64 24483 96 24515
rect 136 24483 168 24515
rect 208 24483 240 24515
rect 280 24483 312 24515
rect 352 24483 384 24515
rect 424 24483 456 24515
rect 496 24483 528 24515
rect 568 24483 600 24515
rect 640 24483 672 24515
rect 712 24483 744 24515
rect 784 24483 816 24515
rect 856 24483 888 24515
rect 928 24483 960 24515
rect 1000 24483 1032 24515
rect 1072 24483 1104 24515
rect 1144 24483 1176 24515
rect 1216 24483 1248 24515
rect 1288 24483 1320 24515
rect 1360 24483 1392 24515
rect 1432 24483 1464 24515
rect 1504 24483 1536 24515
rect 1576 24483 1608 24515
rect 1648 24483 1680 24515
rect 1720 24483 1752 24515
rect 1792 24483 1824 24515
rect 1864 24483 1896 24515
rect 1936 24483 1968 24515
rect 2008 24483 2040 24515
rect 2080 24483 2112 24515
rect 2152 24483 2184 24515
rect 2224 24483 2256 24515
rect 2296 24483 2328 24515
rect 2368 24483 2400 24515
rect 2440 24483 2472 24515
rect 2512 24483 2544 24515
rect 2584 24483 2616 24515
rect 2656 24483 2688 24515
rect 2728 24483 2760 24515
rect 2800 24483 2832 24515
rect 2872 24483 2904 24515
rect 2944 24483 2976 24515
rect 3016 24483 3048 24515
rect 3088 24483 3120 24515
rect 3160 24483 3192 24515
rect 3232 24483 3264 24515
rect 3304 24483 3336 24515
rect 3376 24483 3408 24515
rect 3448 24483 3480 24515
rect 3520 24483 3552 24515
rect 3592 24483 3624 24515
rect 3664 24483 3696 24515
rect 3736 24483 3768 24515
rect 3808 24483 3840 24515
rect 3880 24483 3912 24515
rect 3952 24483 3984 24515
rect 4024 24483 4056 24515
rect 4096 24483 4128 24515
rect 4168 24483 4200 24515
rect 4240 24483 4272 24515
rect 4312 24483 4344 24515
rect 4384 24483 4416 24515
rect 4456 24483 4488 24515
rect 4528 24483 4560 24515
rect 4600 24483 4632 24515
rect 4672 24483 4704 24515
rect 4744 24483 4776 24515
rect 4816 24483 4848 24515
rect 4888 24483 4920 24515
rect 4960 24483 4992 24515
rect 5032 24483 5064 24515
rect 5104 24483 5136 24515
rect 5176 24483 5208 24515
rect 5248 24483 5280 24515
rect 5320 24483 5352 24515
rect 5392 24483 5424 24515
rect 5464 24483 5496 24515
rect 5536 24483 5568 24515
rect 5608 24483 5640 24515
rect 5680 24483 5712 24515
rect 5752 24483 5784 24515
rect 5824 24483 5856 24515
rect 5896 24483 5928 24515
rect 5968 24483 6000 24515
rect 6040 24483 6072 24515
rect 6112 24483 6144 24515
rect 6184 24483 6216 24515
rect 6256 24483 6288 24515
rect 6328 24483 6360 24515
rect 6400 24483 6432 24515
rect 6472 24483 6504 24515
rect 6544 24483 6576 24515
rect 6616 24483 6648 24515
rect 6688 24483 6720 24515
rect 6760 24483 6792 24515
rect 6832 24483 6864 24515
rect 6904 24483 6936 24515
rect 6976 24483 7008 24515
rect 7048 24483 7080 24515
rect 7120 24483 7152 24515
rect 7192 24483 7224 24515
rect 7264 24483 7296 24515
rect 7336 24483 7368 24515
rect 7408 24483 7440 24515
rect 7480 24483 7512 24515
rect 7552 24483 7584 24515
rect 7624 24483 7656 24515
rect 7696 24483 7728 24515
rect 7768 24483 7800 24515
rect 7840 24483 7872 24515
rect 7912 24483 7944 24515
rect 7984 24483 8016 24515
rect 8056 24483 8088 24515
rect 8128 24483 8160 24515
rect 8200 24483 8232 24515
rect 8272 24483 8304 24515
rect 8344 24483 8376 24515
rect 8416 24483 8448 24515
rect 8488 24483 8520 24515
rect 8560 24483 8592 24515
rect 8632 24483 8664 24515
rect 8704 24483 8736 24515
rect 8776 24483 8808 24515
rect 8848 24483 8880 24515
rect 8920 24483 8952 24515
rect 8992 24483 9024 24515
rect 9064 24483 9096 24515
rect 9136 24483 9168 24515
rect 9208 24483 9240 24515
rect 9280 24483 9312 24515
rect 9352 24483 9384 24515
rect 9424 24483 9456 24515
rect 9496 24483 9528 24515
rect 9568 24483 9600 24515
rect 9640 24483 9672 24515
rect 9712 24483 9744 24515
rect 9784 24483 9816 24515
rect 9856 24483 9888 24515
rect 9928 24483 9960 24515
rect 10000 24483 10032 24515
rect 10072 24483 10104 24515
rect 10144 24483 10176 24515
rect 10216 24483 10248 24515
rect 10288 24483 10320 24515
rect 10360 24483 10392 24515
rect 10432 24483 10464 24515
rect 10504 24483 10536 24515
rect 10576 24483 10608 24515
rect 10648 24483 10680 24515
rect 10720 24483 10752 24515
rect 10792 24483 10824 24515
rect 10864 24483 10896 24515
rect 10936 24483 10968 24515
rect 11008 24483 11040 24515
rect 11080 24483 11112 24515
rect 11152 24483 11184 24515
rect 11224 24483 11256 24515
rect 11296 24483 11328 24515
rect 11368 24483 11400 24515
rect 11440 24483 11472 24515
rect 11512 24483 11544 24515
rect 11584 24483 11616 24515
rect 11656 24483 11688 24515
rect 11728 24483 11760 24515
rect 11800 24483 11832 24515
rect 11872 24483 11904 24515
rect 11944 24483 11976 24515
rect 12016 24483 12048 24515
rect 12088 24483 12120 24515
rect 12160 24483 12192 24515
rect 12232 24483 12264 24515
rect 12304 24483 12336 24515
rect 12376 24483 12408 24515
rect 12448 24483 12480 24515
rect 12520 24483 12552 24515
rect 12592 24483 12624 24515
rect 12664 24483 12696 24515
rect 12736 24483 12768 24515
rect 12808 24483 12840 24515
rect 12880 24483 12912 24515
rect 12952 24483 12984 24515
rect 13024 24483 13056 24515
rect 13096 24483 13128 24515
rect 13168 24483 13200 24515
rect 13240 24483 13272 24515
rect 13312 24483 13344 24515
rect 13384 24483 13416 24515
rect 13456 24483 13488 24515
rect 13528 24483 13560 24515
rect 13600 24483 13632 24515
rect 13672 24483 13704 24515
rect 13744 24483 13776 24515
rect 13816 24483 13848 24515
rect 13888 24483 13920 24515
rect 13960 24483 13992 24515
rect 14032 24483 14064 24515
rect 14104 24483 14136 24515
rect 14176 24483 14208 24515
rect 14248 24483 14280 24515
rect 14320 24483 14352 24515
rect 14392 24483 14424 24515
rect 14464 24483 14496 24515
rect 14536 24483 14568 24515
rect 14608 24483 14640 24515
rect 14680 24483 14712 24515
rect 14752 24483 14784 24515
rect 14824 24483 14856 24515
rect 14896 24483 14928 24515
rect 14968 24483 15000 24515
rect 15040 24483 15072 24515
rect 15112 24483 15144 24515
rect 15184 24483 15216 24515
rect 15256 24483 15288 24515
rect 15328 24483 15360 24515
rect 15400 24483 15432 24515
rect 15472 24483 15504 24515
rect 15544 24483 15576 24515
rect 15616 24483 15648 24515
rect 15688 24483 15720 24515
rect 15760 24483 15792 24515
rect 15832 24483 15864 24515
rect 15904 24483 15936 24515
rect 64 24411 96 24443
rect 136 24411 168 24443
rect 208 24411 240 24443
rect 280 24411 312 24443
rect 352 24411 384 24443
rect 424 24411 456 24443
rect 496 24411 528 24443
rect 568 24411 600 24443
rect 640 24411 672 24443
rect 712 24411 744 24443
rect 784 24411 816 24443
rect 856 24411 888 24443
rect 928 24411 960 24443
rect 1000 24411 1032 24443
rect 1072 24411 1104 24443
rect 1144 24411 1176 24443
rect 1216 24411 1248 24443
rect 1288 24411 1320 24443
rect 1360 24411 1392 24443
rect 1432 24411 1464 24443
rect 1504 24411 1536 24443
rect 1576 24411 1608 24443
rect 1648 24411 1680 24443
rect 1720 24411 1752 24443
rect 1792 24411 1824 24443
rect 1864 24411 1896 24443
rect 1936 24411 1968 24443
rect 2008 24411 2040 24443
rect 2080 24411 2112 24443
rect 2152 24411 2184 24443
rect 2224 24411 2256 24443
rect 2296 24411 2328 24443
rect 2368 24411 2400 24443
rect 2440 24411 2472 24443
rect 2512 24411 2544 24443
rect 2584 24411 2616 24443
rect 2656 24411 2688 24443
rect 2728 24411 2760 24443
rect 2800 24411 2832 24443
rect 2872 24411 2904 24443
rect 2944 24411 2976 24443
rect 3016 24411 3048 24443
rect 3088 24411 3120 24443
rect 3160 24411 3192 24443
rect 3232 24411 3264 24443
rect 3304 24411 3336 24443
rect 3376 24411 3408 24443
rect 3448 24411 3480 24443
rect 3520 24411 3552 24443
rect 3592 24411 3624 24443
rect 3664 24411 3696 24443
rect 3736 24411 3768 24443
rect 3808 24411 3840 24443
rect 3880 24411 3912 24443
rect 3952 24411 3984 24443
rect 4024 24411 4056 24443
rect 4096 24411 4128 24443
rect 4168 24411 4200 24443
rect 4240 24411 4272 24443
rect 4312 24411 4344 24443
rect 4384 24411 4416 24443
rect 4456 24411 4488 24443
rect 4528 24411 4560 24443
rect 4600 24411 4632 24443
rect 4672 24411 4704 24443
rect 4744 24411 4776 24443
rect 4816 24411 4848 24443
rect 4888 24411 4920 24443
rect 4960 24411 4992 24443
rect 5032 24411 5064 24443
rect 5104 24411 5136 24443
rect 5176 24411 5208 24443
rect 5248 24411 5280 24443
rect 5320 24411 5352 24443
rect 5392 24411 5424 24443
rect 5464 24411 5496 24443
rect 5536 24411 5568 24443
rect 5608 24411 5640 24443
rect 5680 24411 5712 24443
rect 5752 24411 5784 24443
rect 5824 24411 5856 24443
rect 5896 24411 5928 24443
rect 5968 24411 6000 24443
rect 6040 24411 6072 24443
rect 6112 24411 6144 24443
rect 6184 24411 6216 24443
rect 6256 24411 6288 24443
rect 6328 24411 6360 24443
rect 6400 24411 6432 24443
rect 6472 24411 6504 24443
rect 6544 24411 6576 24443
rect 6616 24411 6648 24443
rect 6688 24411 6720 24443
rect 6760 24411 6792 24443
rect 6832 24411 6864 24443
rect 6904 24411 6936 24443
rect 6976 24411 7008 24443
rect 7048 24411 7080 24443
rect 7120 24411 7152 24443
rect 7192 24411 7224 24443
rect 7264 24411 7296 24443
rect 7336 24411 7368 24443
rect 7408 24411 7440 24443
rect 7480 24411 7512 24443
rect 7552 24411 7584 24443
rect 7624 24411 7656 24443
rect 7696 24411 7728 24443
rect 7768 24411 7800 24443
rect 7840 24411 7872 24443
rect 7912 24411 7944 24443
rect 7984 24411 8016 24443
rect 8056 24411 8088 24443
rect 8128 24411 8160 24443
rect 8200 24411 8232 24443
rect 8272 24411 8304 24443
rect 8344 24411 8376 24443
rect 8416 24411 8448 24443
rect 8488 24411 8520 24443
rect 8560 24411 8592 24443
rect 8632 24411 8664 24443
rect 8704 24411 8736 24443
rect 8776 24411 8808 24443
rect 8848 24411 8880 24443
rect 8920 24411 8952 24443
rect 8992 24411 9024 24443
rect 9064 24411 9096 24443
rect 9136 24411 9168 24443
rect 9208 24411 9240 24443
rect 9280 24411 9312 24443
rect 9352 24411 9384 24443
rect 9424 24411 9456 24443
rect 9496 24411 9528 24443
rect 9568 24411 9600 24443
rect 9640 24411 9672 24443
rect 9712 24411 9744 24443
rect 9784 24411 9816 24443
rect 9856 24411 9888 24443
rect 9928 24411 9960 24443
rect 10000 24411 10032 24443
rect 10072 24411 10104 24443
rect 10144 24411 10176 24443
rect 10216 24411 10248 24443
rect 10288 24411 10320 24443
rect 10360 24411 10392 24443
rect 10432 24411 10464 24443
rect 10504 24411 10536 24443
rect 10576 24411 10608 24443
rect 10648 24411 10680 24443
rect 10720 24411 10752 24443
rect 10792 24411 10824 24443
rect 10864 24411 10896 24443
rect 10936 24411 10968 24443
rect 11008 24411 11040 24443
rect 11080 24411 11112 24443
rect 11152 24411 11184 24443
rect 11224 24411 11256 24443
rect 11296 24411 11328 24443
rect 11368 24411 11400 24443
rect 11440 24411 11472 24443
rect 11512 24411 11544 24443
rect 11584 24411 11616 24443
rect 11656 24411 11688 24443
rect 11728 24411 11760 24443
rect 11800 24411 11832 24443
rect 11872 24411 11904 24443
rect 11944 24411 11976 24443
rect 12016 24411 12048 24443
rect 12088 24411 12120 24443
rect 12160 24411 12192 24443
rect 12232 24411 12264 24443
rect 12304 24411 12336 24443
rect 12376 24411 12408 24443
rect 12448 24411 12480 24443
rect 12520 24411 12552 24443
rect 12592 24411 12624 24443
rect 12664 24411 12696 24443
rect 12736 24411 12768 24443
rect 12808 24411 12840 24443
rect 12880 24411 12912 24443
rect 12952 24411 12984 24443
rect 13024 24411 13056 24443
rect 13096 24411 13128 24443
rect 13168 24411 13200 24443
rect 13240 24411 13272 24443
rect 13312 24411 13344 24443
rect 13384 24411 13416 24443
rect 13456 24411 13488 24443
rect 13528 24411 13560 24443
rect 13600 24411 13632 24443
rect 13672 24411 13704 24443
rect 13744 24411 13776 24443
rect 13816 24411 13848 24443
rect 13888 24411 13920 24443
rect 13960 24411 13992 24443
rect 14032 24411 14064 24443
rect 14104 24411 14136 24443
rect 14176 24411 14208 24443
rect 14248 24411 14280 24443
rect 14320 24411 14352 24443
rect 14392 24411 14424 24443
rect 14464 24411 14496 24443
rect 14536 24411 14568 24443
rect 14608 24411 14640 24443
rect 14680 24411 14712 24443
rect 14752 24411 14784 24443
rect 14824 24411 14856 24443
rect 14896 24411 14928 24443
rect 14968 24411 15000 24443
rect 15040 24411 15072 24443
rect 15112 24411 15144 24443
rect 15184 24411 15216 24443
rect 15256 24411 15288 24443
rect 15328 24411 15360 24443
rect 15400 24411 15432 24443
rect 15472 24411 15504 24443
rect 15544 24411 15576 24443
rect 15616 24411 15648 24443
rect 15688 24411 15720 24443
rect 15760 24411 15792 24443
rect 15832 24411 15864 24443
rect 15904 24411 15936 24443
rect 64 24339 96 24371
rect 136 24339 168 24371
rect 208 24339 240 24371
rect 280 24339 312 24371
rect 352 24339 384 24371
rect 424 24339 456 24371
rect 496 24339 528 24371
rect 568 24339 600 24371
rect 640 24339 672 24371
rect 712 24339 744 24371
rect 784 24339 816 24371
rect 856 24339 888 24371
rect 928 24339 960 24371
rect 1000 24339 1032 24371
rect 1072 24339 1104 24371
rect 1144 24339 1176 24371
rect 1216 24339 1248 24371
rect 1288 24339 1320 24371
rect 1360 24339 1392 24371
rect 1432 24339 1464 24371
rect 1504 24339 1536 24371
rect 1576 24339 1608 24371
rect 1648 24339 1680 24371
rect 1720 24339 1752 24371
rect 1792 24339 1824 24371
rect 1864 24339 1896 24371
rect 1936 24339 1968 24371
rect 2008 24339 2040 24371
rect 2080 24339 2112 24371
rect 2152 24339 2184 24371
rect 2224 24339 2256 24371
rect 2296 24339 2328 24371
rect 2368 24339 2400 24371
rect 2440 24339 2472 24371
rect 2512 24339 2544 24371
rect 2584 24339 2616 24371
rect 2656 24339 2688 24371
rect 2728 24339 2760 24371
rect 2800 24339 2832 24371
rect 2872 24339 2904 24371
rect 2944 24339 2976 24371
rect 3016 24339 3048 24371
rect 3088 24339 3120 24371
rect 3160 24339 3192 24371
rect 3232 24339 3264 24371
rect 3304 24339 3336 24371
rect 3376 24339 3408 24371
rect 3448 24339 3480 24371
rect 3520 24339 3552 24371
rect 3592 24339 3624 24371
rect 3664 24339 3696 24371
rect 3736 24339 3768 24371
rect 3808 24339 3840 24371
rect 3880 24339 3912 24371
rect 3952 24339 3984 24371
rect 4024 24339 4056 24371
rect 4096 24339 4128 24371
rect 4168 24339 4200 24371
rect 4240 24339 4272 24371
rect 4312 24339 4344 24371
rect 4384 24339 4416 24371
rect 4456 24339 4488 24371
rect 4528 24339 4560 24371
rect 4600 24339 4632 24371
rect 4672 24339 4704 24371
rect 4744 24339 4776 24371
rect 4816 24339 4848 24371
rect 4888 24339 4920 24371
rect 4960 24339 4992 24371
rect 5032 24339 5064 24371
rect 5104 24339 5136 24371
rect 5176 24339 5208 24371
rect 5248 24339 5280 24371
rect 5320 24339 5352 24371
rect 5392 24339 5424 24371
rect 5464 24339 5496 24371
rect 5536 24339 5568 24371
rect 5608 24339 5640 24371
rect 5680 24339 5712 24371
rect 5752 24339 5784 24371
rect 5824 24339 5856 24371
rect 5896 24339 5928 24371
rect 5968 24339 6000 24371
rect 6040 24339 6072 24371
rect 6112 24339 6144 24371
rect 6184 24339 6216 24371
rect 6256 24339 6288 24371
rect 6328 24339 6360 24371
rect 6400 24339 6432 24371
rect 6472 24339 6504 24371
rect 6544 24339 6576 24371
rect 6616 24339 6648 24371
rect 6688 24339 6720 24371
rect 6760 24339 6792 24371
rect 6832 24339 6864 24371
rect 6904 24339 6936 24371
rect 6976 24339 7008 24371
rect 7048 24339 7080 24371
rect 7120 24339 7152 24371
rect 7192 24339 7224 24371
rect 7264 24339 7296 24371
rect 7336 24339 7368 24371
rect 7408 24339 7440 24371
rect 7480 24339 7512 24371
rect 7552 24339 7584 24371
rect 7624 24339 7656 24371
rect 7696 24339 7728 24371
rect 7768 24339 7800 24371
rect 7840 24339 7872 24371
rect 7912 24339 7944 24371
rect 7984 24339 8016 24371
rect 8056 24339 8088 24371
rect 8128 24339 8160 24371
rect 8200 24339 8232 24371
rect 8272 24339 8304 24371
rect 8344 24339 8376 24371
rect 8416 24339 8448 24371
rect 8488 24339 8520 24371
rect 8560 24339 8592 24371
rect 8632 24339 8664 24371
rect 8704 24339 8736 24371
rect 8776 24339 8808 24371
rect 8848 24339 8880 24371
rect 8920 24339 8952 24371
rect 8992 24339 9024 24371
rect 9064 24339 9096 24371
rect 9136 24339 9168 24371
rect 9208 24339 9240 24371
rect 9280 24339 9312 24371
rect 9352 24339 9384 24371
rect 9424 24339 9456 24371
rect 9496 24339 9528 24371
rect 9568 24339 9600 24371
rect 9640 24339 9672 24371
rect 9712 24339 9744 24371
rect 9784 24339 9816 24371
rect 9856 24339 9888 24371
rect 9928 24339 9960 24371
rect 10000 24339 10032 24371
rect 10072 24339 10104 24371
rect 10144 24339 10176 24371
rect 10216 24339 10248 24371
rect 10288 24339 10320 24371
rect 10360 24339 10392 24371
rect 10432 24339 10464 24371
rect 10504 24339 10536 24371
rect 10576 24339 10608 24371
rect 10648 24339 10680 24371
rect 10720 24339 10752 24371
rect 10792 24339 10824 24371
rect 10864 24339 10896 24371
rect 10936 24339 10968 24371
rect 11008 24339 11040 24371
rect 11080 24339 11112 24371
rect 11152 24339 11184 24371
rect 11224 24339 11256 24371
rect 11296 24339 11328 24371
rect 11368 24339 11400 24371
rect 11440 24339 11472 24371
rect 11512 24339 11544 24371
rect 11584 24339 11616 24371
rect 11656 24339 11688 24371
rect 11728 24339 11760 24371
rect 11800 24339 11832 24371
rect 11872 24339 11904 24371
rect 11944 24339 11976 24371
rect 12016 24339 12048 24371
rect 12088 24339 12120 24371
rect 12160 24339 12192 24371
rect 12232 24339 12264 24371
rect 12304 24339 12336 24371
rect 12376 24339 12408 24371
rect 12448 24339 12480 24371
rect 12520 24339 12552 24371
rect 12592 24339 12624 24371
rect 12664 24339 12696 24371
rect 12736 24339 12768 24371
rect 12808 24339 12840 24371
rect 12880 24339 12912 24371
rect 12952 24339 12984 24371
rect 13024 24339 13056 24371
rect 13096 24339 13128 24371
rect 13168 24339 13200 24371
rect 13240 24339 13272 24371
rect 13312 24339 13344 24371
rect 13384 24339 13416 24371
rect 13456 24339 13488 24371
rect 13528 24339 13560 24371
rect 13600 24339 13632 24371
rect 13672 24339 13704 24371
rect 13744 24339 13776 24371
rect 13816 24339 13848 24371
rect 13888 24339 13920 24371
rect 13960 24339 13992 24371
rect 14032 24339 14064 24371
rect 14104 24339 14136 24371
rect 14176 24339 14208 24371
rect 14248 24339 14280 24371
rect 14320 24339 14352 24371
rect 14392 24339 14424 24371
rect 14464 24339 14496 24371
rect 14536 24339 14568 24371
rect 14608 24339 14640 24371
rect 14680 24339 14712 24371
rect 14752 24339 14784 24371
rect 14824 24339 14856 24371
rect 14896 24339 14928 24371
rect 14968 24339 15000 24371
rect 15040 24339 15072 24371
rect 15112 24339 15144 24371
rect 15184 24339 15216 24371
rect 15256 24339 15288 24371
rect 15328 24339 15360 24371
rect 15400 24339 15432 24371
rect 15472 24339 15504 24371
rect 15544 24339 15576 24371
rect 15616 24339 15648 24371
rect 15688 24339 15720 24371
rect 15760 24339 15792 24371
rect 15832 24339 15864 24371
rect 15904 24339 15936 24371
rect 64 24267 96 24299
rect 136 24267 168 24299
rect 208 24267 240 24299
rect 280 24267 312 24299
rect 352 24267 384 24299
rect 424 24267 456 24299
rect 496 24267 528 24299
rect 568 24267 600 24299
rect 640 24267 672 24299
rect 712 24267 744 24299
rect 784 24267 816 24299
rect 856 24267 888 24299
rect 928 24267 960 24299
rect 1000 24267 1032 24299
rect 1072 24267 1104 24299
rect 1144 24267 1176 24299
rect 1216 24267 1248 24299
rect 1288 24267 1320 24299
rect 1360 24267 1392 24299
rect 1432 24267 1464 24299
rect 1504 24267 1536 24299
rect 1576 24267 1608 24299
rect 1648 24267 1680 24299
rect 1720 24267 1752 24299
rect 1792 24267 1824 24299
rect 1864 24267 1896 24299
rect 1936 24267 1968 24299
rect 2008 24267 2040 24299
rect 2080 24267 2112 24299
rect 2152 24267 2184 24299
rect 2224 24267 2256 24299
rect 2296 24267 2328 24299
rect 2368 24267 2400 24299
rect 2440 24267 2472 24299
rect 2512 24267 2544 24299
rect 2584 24267 2616 24299
rect 2656 24267 2688 24299
rect 2728 24267 2760 24299
rect 2800 24267 2832 24299
rect 2872 24267 2904 24299
rect 2944 24267 2976 24299
rect 3016 24267 3048 24299
rect 3088 24267 3120 24299
rect 3160 24267 3192 24299
rect 3232 24267 3264 24299
rect 3304 24267 3336 24299
rect 3376 24267 3408 24299
rect 3448 24267 3480 24299
rect 3520 24267 3552 24299
rect 3592 24267 3624 24299
rect 3664 24267 3696 24299
rect 3736 24267 3768 24299
rect 3808 24267 3840 24299
rect 3880 24267 3912 24299
rect 3952 24267 3984 24299
rect 4024 24267 4056 24299
rect 4096 24267 4128 24299
rect 4168 24267 4200 24299
rect 4240 24267 4272 24299
rect 4312 24267 4344 24299
rect 4384 24267 4416 24299
rect 4456 24267 4488 24299
rect 4528 24267 4560 24299
rect 4600 24267 4632 24299
rect 4672 24267 4704 24299
rect 4744 24267 4776 24299
rect 4816 24267 4848 24299
rect 4888 24267 4920 24299
rect 4960 24267 4992 24299
rect 5032 24267 5064 24299
rect 5104 24267 5136 24299
rect 5176 24267 5208 24299
rect 5248 24267 5280 24299
rect 5320 24267 5352 24299
rect 5392 24267 5424 24299
rect 5464 24267 5496 24299
rect 5536 24267 5568 24299
rect 5608 24267 5640 24299
rect 5680 24267 5712 24299
rect 5752 24267 5784 24299
rect 5824 24267 5856 24299
rect 5896 24267 5928 24299
rect 5968 24267 6000 24299
rect 6040 24267 6072 24299
rect 6112 24267 6144 24299
rect 6184 24267 6216 24299
rect 6256 24267 6288 24299
rect 6328 24267 6360 24299
rect 6400 24267 6432 24299
rect 6472 24267 6504 24299
rect 6544 24267 6576 24299
rect 6616 24267 6648 24299
rect 6688 24267 6720 24299
rect 6760 24267 6792 24299
rect 6832 24267 6864 24299
rect 6904 24267 6936 24299
rect 6976 24267 7008 24299
rect 7048 24267 7080 24299
rect 7120 24267 7152 24299
rect 7192 24267 7224 24299
rect 7264 24267 7296 24299
rect 7336 24267 7368 24299
rect 7408 24267 7440 24299
rect 7480 24267 7512 24299
rect 7552 24267 7584 24299
rect 7624 24267 7656 24299
rect 7696 24267 7728 24299
rect 7768 24267 7800 24299
rect 7840 24267 7872 24299
rect 7912 24267 7944 24299
rect 7984 24267 8016 24299
rect 8056 24267 8088 24299
rect 8128 24267 8160 24299
rect 8200 24267 8232 24299
rect 8272 24267 8304 24299
rect 8344 24267 8376 24299
rect 8416 24267 8448 24299
rect 8488 24267 8520 24299
rect 8560 24267 8592 24299
rect 8632 24267 8664 24299
rect 8704 24267 8736 24299
rect 8776 24267 8808 24299
rect 8848 24267 8880 24299
rect 8920 24267 8952 24299
rect 8992 24267 9024 24299
rect 9064 24267 9096 24299
rect 9136 24267 9168 24299
rect 9208 24267 9240 24299
rect 9280 24267 9312 24299
rect 9352 24267 9384 24299
rect 9424 24267 9456 24299
rect 9496 24267 9528 24299
rect 9568 24267 9600 24299
rect 9640 24267 9672 24299
rect 9712 24267 9744 24299
rect 9784 24267 9816 24299
rect 9856 24267 9888 24299
rect 9928 24267 9960 24299
rect 10000 24267 10032 24299
rect 10072 24267 10104 24299
rect 10144 24267 10176 24299
rect 10216 24267 10248 24299
rect 10288 24267 10320 24299
rect 10360 24267 10392 24299
rect 10432 24267 10464 24299
rect 10504 24267 10536 24299
rect 10576 24267 10608 24299
rect 10648 24267 10680 24299
rect 10720 24267 10752 24299
rect 10792 24267 10824 24299
rect 10864 24267 10896 24299
rect 10936 24267 10968 24299
rect 11008 24267 11040 24299
rect 11080 24267 11112 24299
rect 11152 24267 11184 24299
rect 11224 24267 11256 24299
rect 11296 24267 11328 24299
rect 11368 24267 11400 24299
rect 11440 24267 11472 24299
rect 11512 24267 11544 24299
rect 11584 24267 11616 24299
rect 11656 24267 11688 24299
rect 11728 24267 11760 24299
rect 11800 24267 11832 24299
rect 11872 24267 11904 24299
rect 11944 24267 11976 24299
rect 12016 24267 12048 24299
rect 12088 24267 12120 24299
rect 12160 24267 12192 24299
rect 12232 24267 12264 24299
rect 12304 24267 12336 24299
rect 12376 24267 12408 24299
rect 12448 24267 12480 24299
rect 12520 24267 12552 24299
rect 12592 24267 12624 24299
rect 12664 24267 12696 24299
rect 12736 24267 12768 24299
rect 12808 24267 12840 24299
rect 12880 24267 12912 24299
rect 12952 24267 12984 24299
rect 13024 24267 13056 24299
rect 13096 24267 13128 24299
rect 13168 24267 13200 24299
rect 13240 24267 13272 24299
rect 13312 24267 13344 24299
rect 13384 24267 13416 24299
rect 13456 24267 13488 24299
rect 13528 24267 13560 24299
rect 13600 24267 13632 24299
rect 13672 24267 13704 24299
rect 13744 24267 13776 24299
rect 13816 24267 13848 24299
rect 13888 24267 13920 24299
rect 13960 24267 13992 24299
rect 14032 24267 14064 24299
rect 14104 24267 14136 24299
rect 14176 24267 14208 24299
rect 14248 24267 14280 24299
rect 14320 24267 14352 24299
rect 14392 24267 14424 24299
rect 14464 24267 14496 24299
rect 14536 24267 14568 24299
rect 14608 24267 14640 24299
rect 14680 24267 14712 24299
rect 14752 24267 14784 24299
rect 14824 24267 14856 24299
rect 14896 24267 14928 24299
rect 14968 24267 15000 24299
rect 15040 24267 15072 24299
rect 15112 24267 15144 24299
rect 15184 24267 15216 24299
rect 15256 24267 15288 24299
rect 15328 24267 15360 24299
rect 15400 24267 15432 24299
rect 15472 24267 15504 24299
rect 15544 24267 15576 24299
rect 15616 24267 15648 24299
rect 15688 24267 15720 24299
rect 15760 24267 15792 24299
rect 15832 24267 15864 24299
rect 15904 24267 15936 24299
rect 64 24195 96 24227
rect 136 24195 168 24227
rect 208 24195 240 24227
rect 280 24195 312 24227
rect 352 24195 384 24227
rect 424 24195 456 24227
rect 496 24195 528 24227
rect 568 24195 600 24227
rect 640 24195 672 24227
rect 712 24195 744 24227
rect 784 24195 816 24227
rect 856 24195 888 24227
rect 928 24195 960 24227
rect 1000 24195 1032 24227
rect 1072 24195 1104 24227
rect 1144 24195 1176 24227
rect 1216 24195 1248 24227
rect 1288 24195 1320 24227
rect 1360 24195 1392 24227
rect 1432 24195 1464 24227
rect 1504 24195 1536 24227
rect 1576 24195 1608 24227
rect 1648 24195 1680 24227
rect 1720 24195 1752 24227
rect 1792 24195 1824 24227
rect 1864 24195 1896 24227
rect 1936 24195 1968 24227
rect 2008 24195 2040 24227
rect 2080 24195 2112 24227
rect 2152 24195 2184 24227
rect 2224 24195 2256 24227
rect 2296 24195 2328 24227
rect 2368 24195 2400 24227
rect 2440 24195 2472 24227
rect 2512 24195 2544 24227
rect 2584 24195 2616 24227
rect 2656 24195 2688 24227
rect 2728 24195 2760 24227
rect 2800 24195 2832 24227
rect 2872 24195 2904 24227
rect 2944 24195 2976 24227
rect 3016 24195 3048 24227
rect 3088 24195 3120 24227
rect 3160 24195 3192 24227
rect 3232 24195 3264 24227
rect 3304 24195 3336 24227
rect 3376 24195 3408 24227
rect 3448 24195 3480 24227
rect 3520 24195 3552 24227
rect 3592 24195 3624 24227
rect 3664 24195 3696 24227
rect 3736 24195 3768 24227
rect 3808 24195 3840 24227
rect 3880 24195 3912 24227
rect 3952 24195 3984 24227
rect 4024 24195 4056 24227
rect 4096 24195 4128 24227
rect 4168 24195 4200 24227
rect 4240 24195 4272 24227
rect 4312 24195 4344 24227
rect 4384 24195 4416 24227
rect 4456 24195 4488 24227
rect 4528 24195 4560 24227
rect 4600 24195 4632 24227
rect 4672 24195 4704 24227
rect 4744 24195 4776 24227
rect 4816 24195 4848 24227
rect 4888 24195 4920 24227
rect 4960 24195 4992 24227
rect 5032 24195 5064 24227
rect 5104 24195 5136 24227
rect 5176 24195 5208 24227
rect 5248 24195 5280 24227
rect 5320 24195 5352 24227
rect 5392 24195 5424 24227
rect 5464 24195 5496 24227
rect 5536 24195 5568 24227
rect 5608 24195 5640 24227
rect 5680 24195 5712 24227
rect 5752 24195 5784 24227
rect 5824 24195 5856 24227
rect 5896 24195 5928 24227
rect 5968 24195 6000 24227
rect 6040 24195 6072 24227
rect 6112 24195 6144 24227
rect 6184 24195 6216 24227
rect 6256 24195 6288 24227
rect 6328 24195 6360 24227
rect 6400 24195 6432 24227
rect 6472 24195 6504 24227
rect 6544 24195 6576 24227
rect 6616 24195 6648 24227
rect 6688 24195 6720 24227
rect 6760 24195 6792 24227
rect 6832 24195 6864 24227
rect 6904 24195 6936 24227
rect 6976 24195 7008 24227
rect 7048 24195 7080 24227
rect 7120 24195 7152 24227
rect 7192 24195 7224 24227
rect 7264 24195 7296 24227
rect 7336 24195 7368 24227
rect 7408 24195 7440 24227
rect 7480 24195 7512 24227
rect 7552 24195 7584 24227
rect 7624 24195 7656 24227
rect 7696 24195 7728 24227
rect 7768 24195 7800 24227
rect 7840 24195 7872 24227
rect 7912 24195 7944 24227
rect 7984 24195 8016 24227
rect 8056 24195 8088 24227
rect 8128 24195 8160 24227
rect 8200 24195 8232 24227
rect 8272 24195 8304 24227
rect 8344 24195 8376 24227
rect 8416 24195 8448 24227
rect 8488 24195 8520 24227
rect 8560 24195 8592 24227
rect 8632 24195 8664 24227
rect 8704 24195 8736 24227
rect 8776 24195 8808 24227
rect 8848 24195 8880 24227
rect 8920 24195 8952 24227
rect 8992 24195 9024 24227
rect 9064 24195 9096 24227
rect 9136 24195 9168 24227
rect 9208 24195 9240 24227
rect 9280 24195 9312 24227
rect 9352 24195 9384 24227
rect 9424 24195 9456 24227
rect 9496 24195 9528 24227
rect 9568 24195 9600 24227
rect 9640 24195 9672 24227
rect 9712 24195 9744 24227
rect 9784 24195 9816 24227
rect 9856 24195 9888 24227
rect 9928 24195 9960 24227
rect 10000 24195 10032 24227
rect 10072 24195 10104 24227
rect 10144 24195 10176 24227
rect 10216 24195 10248 24227
rect 10288 24195 10320 24227
rect 10360 24195 10392 24227
rect 10432 24195 10464 24227
rect 10504 24195 10536 24227
rect 10576 24195 10608 24227
rect 10648 24195 10680 24227
rect 10720 24195 10752 24227
rect 10792 24195 10824 24227
rect 10864 24195 10896 24227
rect 10936 24195 10968 24227
rect 11008 24195 11040 24227
rect 11080 24195 11112 24227
rect 11152 24195 11184 24227
rect 11224 24195 11256 24227
rect 11296 24195 11328 24227
rect 11368 24195 11400 24227
rect 11440 24195 11472 24227
rect 11512 24195 11544 24227
rect 11584 24195 11616 24227
rect 11656 24195 11688 24227
rect 11728 24195 11760 24227
rect 11800 24195 11832 24227
rect 11872 24195 11904 24227
rect 11944 24195 11976 24227
rect 12016 24195 12048 24227
rect 12088 24195 12120 24227
rect 12160 24195 12192 24227
rect 12232 24195 12264 24227
rect 12304 24195 12336 24227
rect 12376 24195 12408 24227
rect 12448 24195 12480 24227
rect 12520 24195 12552 24227
rect 12592 24195 12624 24227
rect 12664 24195 12696 24227
rect 12736 24195 12768 24227
rect 12808 24195 12840 24227
rect 12880 24195 12912 24227
rect 12952 24195 12984 24227
rect 13024 24195 13056 24227
rect 13096 24195 13128 24227
rect 13168 24195 13200 24227
rect 13240 24195 13272 24227
rect 13312 24195 13344 24227
rect 13384 24195 13416 24227
rect 13456 24195 13488 24227
rect 13528 24195 13560 24227
rect 13600 24195 13632 24227
rect 13672 24195 13704 24227
rect 13744 24195 13776 24227
rect 13816 24195 13848 24227
rect 13888 24195 13920 24227
rect 13960 24195 13992 24227
rect 14032 24195 14064 24227
rect 14104 24195 14136 24227
rect 14176 24195 14208 24227
rect 14248 24195 14280 24227
rect 14320 24195 14352 24227
rect 14392 24195 14424 24227
rect 14464 24195 14496 24227
rect 14536 24195 14568 24227
rect 14608 24195 14640 24227
rect 14680 24195 14712 24227
rect 14752 24195 14784 24227
rect 14824 24195 14856 24227
rect 14896 24195 14928 24227
rect 14968 24195 15000 24227
rect 15040 24195 15072 24227
rect 15112 24195 15144 24227
rect 15184 24195 15216 24227
rect 15256 24195 15288 24227
rect 15328 24195 15360 24227
rect 15400 24195 15432 24227
rect 15472 24195 15504 24227
rect 15544 24195 15576 24227
rect 15616 24195 15648 24227
rect 15688 24195 15720 24227
rect 15760 24195 15792 24227
rect 15832 24195 15864 24227
rect 15904 24195 15936 24227
rect 64 24123 96 24155
rect 136 24123 168 24155
rect 208 24123 240 24155
rect 280 24123 312 24155
rect 352 24123 384 24155
rect 424 24123 456 24155
rect 496 24123 528 24155
rect 568 24123 600 24155
rect 640 24123 672 24155
rect 712 24123 744 24155
rect 784 24123 816 24155
rect 856 24123 888 24155
rect 928 24123 960 24155
rect 1000 24123 1032 24155
rect 1072 24123 1104 24155
rect 1144 24123 1176 24155
rect 1216 24123 1248 24155
rect 1288 24123 1320 24155
rect 1360 24123 1392 24155
rect 1432 24123 1464 24155
rect 1504 24123 1536 24155
rect 1576 24123 1608 24155
rect 1648 24123 1680 24155
rect 1720 24123 1752 24155
rect 1792 24123 1824 24155
rect 1864 24123 1896 24155
rect 1936 24123 1968 24155
rect 2008 24123 2040 24155
rect 2080 24123 2112 24155
rect 2152 24123 2184 24155
rect 2224 24123 2256 24155
rect 2296 24123 2328 24155
rect 2368 24123 2400 24155
rect 2440 24123 2472 24155
rect 2512 24123 2544 24155
rect 2584 24123 2616 24155
rect 2656 24123 2688 24155
rect 2728 24123 2760 24155
rect 2800 24123 2832 24155
rect 2872 24123 2904 24155
rect 2944 24123 2976 24155
rect 3016 24123 3048 24155
rect 3088 24123 3120 24155
rect 3160 24123 3192 24155
rect 3232 24123 3264 24155
rect 3304 24123 3336 24155
rect 3376 24123 3408 24155
rect 3448 24123 3480 24155
rect 3520 24123 3552 24155
rect 3592 24123 3624 24155
rect 3664 24123 3696 24155
rect 3736 24123 3768 24155
rect 3808 24123 3840 24155
rect 3880 24123 3912 24155
rect 3952 24123 3984 24155
rect 4024 24123 4056 24155
rect 4096 24123 4128 24155
rect 4168 24123 4200 24155
rect 4240 24123 4272 24155
rect 4312 24123 4344 24155
rect 4384 24123 4416 24155
rect 4456 24123 4488 24155
rect 4528 24123 4560 24155
rect 4600 24123 4632 24155
rect 4672 24123 4704 24155
rect 4744 24123 4776 24155
rect 4816 24123 4848 24155
rect 4888 24123 4920 24155
rect 4960 24123 4992 24155
rect 5032 24123 5064 24155
rect 5104 24123 5136 24155
rect 5176 24123 5208 24155
rect 5248 24123 5280 24155
rect 5320 24123 5352 24155
rect 5392 24123 5424 24155
rect 5464 24123 5496 24155
rect 5536 24123 5568 24155
rect 5608 24123 5640 24155
rect 5680 24123 5712 24155
rect 5752 24123 5784 24155
rect 5824 24123 5856 24155
rect 5896 24123 5928 24155
rect 5968 24123 6000 24155
rect 6040 24123 6072 24155
rect 6112 24123 6144 24155
rect 6184 24123 6216 24155
rect 6256 24123 6288 24155
rect 6328 24123 6360 24155
rect 6400 24123 6432 24155
rect 6472 24123 6504 24155
rect 6544 24123 6576 24155
rect 6616 24123 6648 24155
rect 6688 24123 6720 24155
rect 6760 24123 6792 24155
rect 6832 24123 6864 24155
rect 6904 24123 6936 24155
rect 6976 24123 7008 24155
rect 7048 24123 7080 24155
rect 7120 24123 7152 24155
rect 7192 24123 7224 24155
rect 7264 24123 7296 24155
rect 7336 24123 7368 24155
rect 7408 24123 7440 24155
rect 7480 24123 7512 24155
rect 7552 24123 7584 24155
rect 7624 24123 7656 24155
rect 7696 24123 7728 24155
rect 7768 24123 7800 24155
rect 7840 24123 7872 24155
rect 7912 24123 7944 24155
rect 7984 24123 8016 24155
rect 8056 24123 8088 24155
rect 8128 24123 8160 24155
rect 8200 24123 8232 24155
rect 8272 24123 8304 24155
rect 8344 24123 8376 24155
rect 8416 24123 8448 24155
rect 8488 24123 8520 24155
rect 8560 24123 8592 24155
rect 8632 24123 8664 24155
rect 8704 24123 8736 24155
rect 8776 24123 8808 24155
rect 8848 24123 8880 24155
rect 8920 24123 8952 24155
rect 8992 24123 9024 24155
rect 9064 24123 9096 24155
rect 9136 24123 9168 24155
rect 9208 24123 9240 24155
rect 9280 24123 9312 24155
rect 9352 24123 9384 24155
rect 9424 24123 9456 24155
rect 9496 24123 9528 24155
rect 9568 24123 9600 24155
rect 9640 24123 9672 24155
rect 9712 24123 9744 24155
rect 9784 24123 9816 24155
rect 9856 24123 9888 24155
rect 9928 24123 9960 24155
rect 10000 24123 10032 24155
rect 10072 24123 10104 24155
rect 10144 24123 10176 24155
rect 10216 24123 10248 24155
rect 10288 24123 10320 24155
rect 10360 24123 10392 24155
rect 10432 24123 10464 24155
rect 10504 24123 10536 24155
rect 10576 24123 10608 24155
rect 10648 24123 10680 24155
rect 10720 24123 10752 24155
rect 10792 24123 10824 24155
rect 10864 24123 10896 24155
rect 10936 24123 10968 24155
rect 11008 24123 11040 24155
rect 11080 24123 11112 24155
rect 11152 24123 11184 24155
rect 11224 24123 11256 24155
rect 11296 24123 11328 24155
rect 11368 24123 11400 24155
rect 11440 24123 11472 24155
rect 11512 24123 11544 24155
rect 11584 24123 11616 24155
rect 11656 24123 11688 24155
rect 11728 24123 11760 24155
rect 11800 24123 11832 24155
rect 11872 24123 11904 24155
rect 11944 24123 11976 24155
rect 12016 24123 12048 24155
rect 12088 24123 12120 24155
rect 12160 24123 12192 24155
rect 12232 24123 12264 24155
rect 12304 24123 12336 24155
rect 12376 24123 12408 24155
rect 12448 24123 12480 24155
rect 12520 24123 12552 24155
rect 12592 24123 12624 24155
rect 12664 24123 12696 24155
rect 12736 24123 12768 24155
rect 12808 24123 12840 24155
rect 12880 24123 12912 24155
rect 12952 24123 12984 24155
rect 13024 24123 13056 24155
rect 13096 24123 13128 24155
rect 13168 24123 13200 24155
rect 13240 24123 13272 24155
rect 13312 24123 13344 24155
rect 13384 24123 13416 24155
rect 13456 24123 13488 24155
rect 13528 24123 13560 24155
rect 13600 24123 13632 24155
rect 13672 24123 13704 24155
rect 13744 24123 13776 24155
rect 13816 24123 13848 24155
rect 13888 24123 13920 24155
rect 13960 24123 13992 24155
rect 14032 24123 14064 24155
rect 14104 24123 14136 24155
rect 14176 24123 14208 24155
rect 14248 24123 14280 24155
rect 14320 24123 14352 24155
rect 14392 24123 14424 24155
rect 14464 24123 14496 24155
rect 14536 24123 14568 24155
rect 14608 24123 14640 24155
rect 14680 24123 14712 24155
rect 14752 24123 14784 24155
rect 14824 24123 14856 24155
rect 14896 24123 14928 24155
rect 14968 24123 15000 24155
rect 15040 24123 15072 24155
rect 15112 24123 15144 24155
rect 15184 24123 15216 24155
rect 15256 24123 15288 24155
rect 15328 24123 15360 24155
rect 15400 24123 15432 24155
rect 15472 24123 15504 24155
rect 15544 24123 15576 24155
rect 15616 24123 15648 24155
rect 15688 24123 15720 24155
rect 15760 24123 15792 24155
rect 15832 24123 15864 24155
rect 15904 24123 15936 24155
rect 64 24051 96 24083
rect 136 24051 168 24083
rect 208 24051 240 24083
rect 280 24051 312 24083
rect 352 24051 384 24083
rect 424 24051 456 24083
rect 496 24051 528 24083
rect 568 24051 600 24083
rect 640 24051 672 24083
rect 712 24051 744 24083
rect 784 24051 816 24083
rect 856 24051 888 24083
rect 928 24051 960 24083
rect 1000 24051 1032 24083
rect 1072 24051 1104 24083
rect 1144 24051 1176 24083
rect 1216 24051 1248 24083
rect 1288 24051 1320 24083
rect 1360 24051 1392 24083
rect 1432 24051 1464 24083
rect 1504 24051 1536 24083
rect 1576 24051 1608 24083
rect 1648 24051 1680 24083
rect 1720 24051 1752 24083
rect 1792 24051 1824 24083
rect 1864 24051 1896 24083
rect 1936 24051 1968 24083
rect 2008 24051 2040 24083
rect 2080 24051 2112 24083
rect 2152 24051 2184 24083
rect 2224 24051 2256 24083
rect 2296 24051 2328 24083
rect 2368 24051 2400 24083
rect 2440 24051 2472 24083
rect 2512 24051 2544 24083
rect 2584 24051 2616 24083
rect 2656 24051 2688 24083
rect 2728 24051 2760 24083
rect 2800 24051 2832 24083
rect 2872 24051 2904 24083
rect 2944 24051 2976 24083
rect 3016 24051 3048 24083
rect 3088 24051 3120 24083
rect 3160 24051 3192 24083
rect 3232 24051 3264 24083
rect 3304 24051 3336 24083
rect 3376 24051 3408 24083
rect 3448 24051 3480 24083
rect 3520 24051 3552 24083
rect 3592 24051 3624 24083
rect 3664 24051 3696 24083
rect 3736 24051 3768 24083
rect 3808 24051 3840 24083
rect 3880 24051 3912 24083
rect 3952 24051 3984 24083
rect 4024 24051 4056 24083
rect 4096 24051 4128 24083
rect 4168 24051 4200 24083
rect 4240 24051 4272 24083
rect 4312 24051 4344 24083
rect 4384 24051 4416 24083
rect 4456 24051 4488 24083
rect 4528 24051 4560 24083
rect 4600 24051 4632 24083
rect 4672 24051 4704 24083
rect 4744 24051 4776 24083
rect 4816 24051 4848 24083
rect 4888 24051 4920 24083
rect 4960 24051 4992 24083
rect 5032 24051 5064 24083
rect 5104 24051 5136 24083
rect 5176 24051 5208 24083
rect 5248 24051 5280 24083
rect 5320 24051 5352 24083
rect 5392 24051 5424 24083
rect 5464 24051 5496 24083
rect 5536 24051 5568 24083
rect 5608 24051 5640 24083
rect 5680 24051 5712 24083
rect 5752 24051 5784 24083
rect 5824 24051 5856 24083
rect 5896 24051 5928 24083
rect 5968 24051 6000 24083
rect 6040 24051 6072 24083
rect 6112 24051 6144 24083
rect 6184 24051 6216 24083
rect 6256 24051 6288 24083
rect 6328 24051 6360 24083
rect 6400 24051 6432 24083
rect 6472 24051 6504 24083
rect 6544 24051 6576 24083
rect 6616 24051 6648 24083
rect 6688 24051 6720 24083
rect 6760 24051 6792 24083
rect 6832 24051 6864 24083
rect 6904 24051 6936 24083
rect 6976 24051 7008 24083
rect 7048 24051 7080 24083
rect 7120 24051 7152 24083
rect 7192 24051 7224 24083
rect 7264 24051 7296 24083
rect 7336 24051 7368 24083
rect 7408 24051 7440 24083
rect 7480 24051 7512 24083
rect 7552 24051 7584 24083
rect 7624 24051 7656 24083
rect 7696 24051 7728 24083
rect 7768 24051 7800 24083
rect 7840 24051 7872 24083
rect 7912 24051 7944 24083
rect 7984 24051 8016 24083
rect 8056 24051 8088 24083
rect 8128 24051 8160 24083
rect 8200 24051 8232 24083
rect 8272 24051 8304 24083
rect 8344 24051 8376 24083
rect 8416 24051 8448 24083
rect 8488 24051 8520 24083
rect 8560 24051 8592 24083
rect 8632 24051 8664 24083
rect 8704 24051 8736 24083
rect 8776 24051 8808 24083
rect 8848 24051 8880 24083
rect 8920 24051 8952 24083
rect 8992 24051 9024 24083
rect 9064 24051 9096 24083
rect 9136 24051 9168 24083
rect 9208 24051 9240 24083
rect 9280 24051 9312 24083
rect 9352 24051 9384 24083
rect 9424 24051 9456 24083
rect 9496 24051 9528 24083
rect 9568 24051 9600 24083
rect 9640 24051 9672 24083
rect 9712 24051 9744 24083
rect 9784 24051 9816 24083
rect 9856 24051 9888 24083
rect 9928 24051 9960 24083
rect 10000 24051 10032 24083
rect 10072 24051 10104 24083
rect 10144 24051 10176 24083
rect 10216 24051 10248 24083
rect 10288 24051 10320 24083
rect 10360 24051 10392 24083
rect 10432 24051 10464 24083
rect 10504 24051 10536 24083
rect 10576 24051 10608 24083
rect 10648 24051 10680 24083
rect 10720 24051 10752 24083
rect 10792 24051 10824 24083
rect 10864 24051 10896 24083
rect 10936 24051 10968 24083
rect 11008 24051 11040 24083
rect 11080 24051 11112 24083
rect 11152 24051 11184 24083
rect 11224 24051 11256 24083
rect 11296 24051 11328 24083
rect 11368 24051 11400 24083
rect 11440 24051 11472 24083
rect 11512 24051 11544 24083
rect 11584 24051 11616 24083
rect 11656 24051 11688 24083
rect 11728 24051 11760 24083
rect 11800 24051 11832 24083
rect 11872 24051 11904 24083
rect 11944 24051 11976 24083
rect 12016 24051 12048 24083
rect 12088 24051 12120 24083
rect 12160 24051 12192 24083
rect 12232 24051 12264 24083
rect 12304 24051 12336 24083
rect 12376 24051 12408 24083
rect 12448 24051 12480 24083
rect 12520 24051 12552 24083
rect 12592 24051 12624 24083
rect 12664 24051 12696 24083
rect 12736 24051 12768 24083
rect 12808 24051 12840 24083
rect 12880 24051 12912 24083
rect 12952 24051 12984 24083
rect 13024 24051 13056 24083
rect 13096 24051 13128 24083
rect 13168 24051 13200 24083
rect 13240 24051 13272 24083
rect 13312 24051 13344 24083
rect 13384 24051 13416 24083
rect 13456 24051 13488 24083
rect 13528 24051 13560 24083
rect 13600 24051 13632 24083
rect 13672 24051 13704 24083
rect 13744 24051 13776 24083
rect 13816 24051 13848 24083
rect 13888 24051 13920 24083
rect 13960 24051 13992 24083
rect 14032 24051 14064 24083
rect 14104 24051 14136 24083
rect 14176 24051 14208 24083
rect 14248 24051 14280 24083
rect 14320 24051 14352 24083
rect 14392 24051 14424 24083
rect 14464 24051 14496 24083
rect 14536 24051 14568 24083
rect 14608 24051 14640 24083
rect 14680 24051 14712 24083
rect 14752 24051 14784 24083
rect 14824 24051 14856 24083
rect 14896 24051 14928 24083
rect 14968 24051 15000 24083
rect 15040 24051 15072 24083
rect 15112 24051 15144 24083
rect 15184 24051 15216 24083
rect 15256 24051 15288 24083
rect 15328 24051 15360 24083
rect 15400 24051 15432 24083
rect 15472 24051 15504 24083
rect 15544 24051 15576 24083
rect 15616 24051 15648 24083
rect 15688 24051 15720 24083
rect 15760 24051 15792 24083
rect 15832 24051 15864 24083
rect 15904 24051 15936 24083
rect 64 23979 96 24011
rect 136 23979 168 24011
rect 208 23979 240 24011
rect 280 23979 312 24011
rect 352 23979 384 24011
rect 424 23979 456 24011
rect 496 23979 528 24011
rect 568 23979 600 24011
rect 640 23979 672 24011
rect 712 23979 744 24011
rect 784 23979 816 24011
rect 856 23979 888 24011
rect 928 23979 960 24011
rect 1000 23979 1032 24011
rect 1072 23979 1104 24011
rect 1144 23979 1176 24011
rect 1216 23979 1248 24011
rect 1288 23979 1320 24011
rect 1360 23979 1392 24011
rect 1432 23979 1464 24011
rect 1504 23979 1536 24011
rect 1576 23979 1608 24011
rect 1648 23979 1680 24011
rect 1720 23979 1752 24011
rect 1792 23979 1824 24011
rect 1864 23979 1896 24011
rect 1936 23979 1968 24011
rect 2008 23979 2040 24011
rect 2080 23979 2112 24011
rect 2152 23979 2184 24011
rect 2224 23979 2256 24011
rect 2296 23979 2328 24011
rect 2368 23979 2400 24011
rect 2440 23979 2472 24011
rect 2512 23979 2544 24011
rect 2584 23979 2616 24011
rect 2656 23979 2688 24011
rect 2728 23979 2760 24011
rect 2800 23979 2832 24011
rect 2872 23979 2904 24011
rect 2944 23979 2976 24011
rect 3016 23979 3048 24011
rect 3088 23979 3120 24011
rect 3160 23979 3192 24011
rect 3232 23979 3264 24011
rect 3304 23979 3336 24011
rect 3376 23979 3408 24011
rect 3448 23979 3480 24011
rect 3520 23979 3552 24011
rect 3592 23979 3624 24011
rect 3664 23979 3696 24011
rect 3736 23979 3768 24011
rect 3808 23979 3840 24011
rect 3880 23979 3912 24011
rect 3952 23979 3984 24011
rect 4024 23979 4056 24011
rect 4096 23979 4128 24011
rect 4168 23979 4200 24011
rect 4240 23979 4272 24011
rect 4312 23979 4344 24011
rect 4384 23979 4416 24011
rect 4456 23979 4488 24011
rect 4528 23979 4560 24011
rect 4600 23979 4632 24011
rect 4672 23979 4704 24011
rect 4744 23979 4776 24011
rect 4816 23979 4848 24011
rect 4888 23979 4920 24011
rect 4960 23979 4992 24011
rect 5032 23979 5064 24011
rect 5104 23979 5136 24011
rect 5176 23979 5208 24011
rect 5248 23979 5280 24011
rect 5320 23979 5352 24011
rect 5392 23979 5424 24011
rect 5464 23979 5496 24011
rect 5536 23979 5568 24011
rect 5608 23979 5640 24011
rect 5680 23979 5712 24011
rect 5752 23979 5784 24011
rect 5824 23979 5856 24011
rect 5896 23979 5928 24011
rect 5968 23979 6000 24011
rect 6040 23979 6072 24011
rect 6112 23979 6144 24011
rect 6184 23979 6216 24011
rect 6256 23979 6288 24011
rect 6328 23979 6360 24011
rect 6400 23979 6432 24011
rect 6472 23979 6504 24011
rect 6544 23979 6576 24011
rect 6616 23979 6648 24011
rect 6688 23979 6720 24011
rect 6760 23979 6792 24011
rect 6832 23979 6864 24011
rect 6904 23979 6936 24011
rect 6976 23979 7008 24011
rect 7048 23979 7080 24011
rect 7120 23979 7152 24011
rect 7192 23979 7224 24011
rect 7264 23979 7296 24011
rect 7336 23979 7368 24011
rect 7408 23979 7440 24011
rect 7480 23979 7512 24011
rect 7552 23979 7584 24011
rect 7624 23979 7656 24011
rect 7696 23979 7728 24011
rect 7768 23979 7800 24011
rect 7840 23979 7872 24011
rect 7912 23979 7944 24011
rect 7984 23979 8016 24011
rect 8056 23979 8088 24011
rect 8128 23979 8160 24011
rect 8200 23979 8232 24011
rect 8272 23979 8304 24011
rect 8344 23979 8376 24011
rect 8416 23979 8448 24011
rect 8488 23979 8520 24011
rect 8560 23979 8592 24011
rect 8632 23979 8664 24011
rect 8704 23979 8736 24011
rect 8776 23979 8808 24011
rect 8848 23979 8880 24011
rect 8920 23979 8952 24011
rect 8992 23979 9024 24011
rect 9064 23979 9096 24011
rect 9136 23979 9168 24011
rect 9208 23979 9240 24011
rect 9280 23979 9312 24011
rect 9352 23979 9384 24011
rect 9424 23979 9456 24011
rect 9496 23979 9528 24011
rect 9568 23979 9600 24011
rect 9640 23979 9672 24011
rect 9712 23979 9744 24011
rect 9784 23979 9816 24011
rect 9856 23979 9888 24011
rect 9928 23979 9960 24011
rect 10000 23979 10032 24011
rect 10072 23979 10104 24011
rect 10144 23979 10176 24011
rect 10216 23979 10248 24011
rect 10288 23979 10320 24011
rect 10360 23979 10392 24011
rect 10432 23979 10464 24011
rect 10504 23979 10536 24011
rect 10576 23979 10608 24011
rect 10648 23979 10680 24011
rect 10720 23979 10752 24011
rect 10792 23979 10824 24011
rect 10864 23979 10896 24011
rect 10936 23979 10968 24011
rect 11008 23979 11040 24011
rect 11080 23979 11112 24011
rect 11152 23979 11184 24011
rect 11224 23979 11256 24011
rect 11296 23979 11328 24011
rect 11368 23979 11400 24011
rect 11440 23979 11472 24011
rect 11512 23979 11544 24011
rect 11584 23979 11616 24011
rect 11656 23979 11688 24011
rect 11728 23979 11760 24011
rect 11800 23979 11832 24011
rect 11872 23979 11904 24011
rect 11944 23979 11976 24011
rect 12016 23979 12048 24011
rect 12088 23979 12120 24011
rect 12160 23979 12192 24011
rect 12232 23979 12264 24011
rect 12304 23979 12336 24011
rect 12376 23979 12408 24011
rect 12448 23979 12480 24011
rect 12520 23979 12552 24011
rect 12592 23979 12624 24011
rect 12664 23979 12696 24011
rect 12736 23979 12768 24011
rect 12808 23979 12840 24011
rect 12880 23979 12912 24011
rect 12952 23979 12984 24011
rect 13024 23979 13056 24011
rect 13096 23979 13128 24011
rect 13168 23979 13200 24011
rect 13240 23979 13272 24011
rect 13312 23979 13344 24011
rect 13384 23979 13416 24011
rect 13456 23979 13488 24011
rect 13528 23979 13560 24011
rect 13600 23979 13632 24011
rect 13672 23979 13704 24011
rect 13744 23979 13776 24011
rect 13816 23979 13848 24011
rect 13888 23979 13920 24011
rect 13960 23979 13992 24011
rect 14032 23979 14064 24011
rect 14104 23979 14136 24011
rect 14176 23979 14208 24011
rect 14248 23979 14280 24011
rect 14320 23979 14352 24011
rect 14392 23979 14424 24011
rect 14464 23979 14496 24011
rect 14536 23979 14568 24011
rect 14608 23979 14640 24011
rect 14680 23979 14712 24011
rect 14752 23979 14784 24011
rect 14824 23979 14856 24011
rect 14896 23979 14928 24011
rect 14968 23979 15000 24011
rect 15040 23979 15072 24011
rect 15112 23979 15144 24011
rect 15184 23979 15216 24011
rect 15256 23979 15288 24011
rect 15328 23979 15360 24011
rect 15400 23979 15432 24011
rect 15472 23979 15504 24011
rect 15544 23979 15576 24011
rect 15616 23979 15648 24011
rect 15688 23979 15720 24011
rect 15760 23979 15792 24011
rect 15832 23979 15864 24011
rect 15904 23979 15936 24011
rect 64 23907 96 23939
rect 136 23907 168 23939
rect 208 23907 240 23939
rect 280 23907 312 23939
rect 352 23907 384 23939
rect 424 23907 456 23939
rect 496 23907 528 23939
rect 568 23907 600 23939
rect 640 23907 672 23939
rect 712 23907 744 23939
rect 784 23907 816 23939
rect 856 23907 888 23939
rect 928 23907 960 23939
rect 1000 23907 1032 23939
rect 1072 23907 1104 23939
rect 1144 23907 1176 23939
rect 1216 23907 1248 23939
rect 1288 23907 1320 23939
rect 1360 23907 1392 23939
rect 1432 23907 1464 23939
rect 1504 23907 1536 23939
rect 1576 23907 1608 23939
rect 1648 23907 1680 23939
rect 1720 23907 1752 23939
rect 1792 23907 1824 23939
rect 1864 23907 1896 23939
rect 1936 23907 1968 23939
rect 2008 23907 2040 23939
rect 2080 23907 2112 23939
rect 2152 23907 2184 23939
rect 2224 23907 2256 23939
rect 2296 23907 2328 23939
rect 2368 23907 2400 23939
rect 2440 23907 2472 23939
rect 2512 23907 2544 23939
rect 2584 23907 2616 23939
rect 2656 23907 2688 23939
rect 2728 23907 2760 23939
rect 2800 23907 2832 23939
rect 2872 23907 2904 23939
rect 2944 23907 2976 23939
rect 3016 23907 3048 23939
rect 3088 23907 3120 23939
rect 3160 23907 3192 23939
rect 3232 23907 3264 23939
rect 3304 23907 3336 23939
rect 3376 23907 3408 23939
rect 3448 23907 3480 23939
rect 3520 23907 3552 23939
rect 3592 23907 3624 23939
rect 3664 23907 3696 23939
rect 3736 23907 3768 23939
rect 3808 23907 3840 23939
rect 3880 23907 3912 23939
rect 3952 23907 3984 23939
rect 4024 23907 4056 23939
rect 4096 23907 4128 23939
rect 4168 23907 4200 23939
rect 4240 23907 4272 23939
rect 4312 23907 4344 23939
rect 4384 23907 4416 23939
rect 4456 23907 4488 23939
rect 4528 23907 4560 23939
rect 4600 23907 4632 23939
rect 4672 23907 4704 23939
rect 4744 23907 4776 23939
rect 4816 23907 4848 23939
rect 4888 23907 4920 23939
rect 4960 23907 4992 23939
rect 5032 23907 5064 23939
rect 5104 23907 5136 23939
rect 5176 23907 5208 23939
rect 5248 23907 5280 23939
rect 5320 23907 5352 23939
rect 5392 23907 5424 23939
rect 5464 23907 5496 23939
rect 5536 23907 5568 23939
rect 5608 23907 5640 23939
rect 5680 23907 5712 23939
rect 5752 23907 5784 23939
rect 5824 23907 5856 23939
rect 5896 23907 5928 23939
rect 5968 23907 6000 23939
rect 6040 23907 6072 23939
rect 6112 23907 6144 23939
rect 6184 23907 6216 23939
rect 6256 23907 6288 23939
rect 6328 23907 6360 23939
rect 6400 23907 6432 23939
rect 6472 23907 6504 23939
rect 6544 23907 6576 23939
rect 6616 23907 6648 23939
rect 6688 23907 6720 23939
rect 6760 23907 6792 23939
rect 6832 23907 6864 23939
rect 6904 23907 6936 23939
rect 6976 23907 7008 23939
rect 7048 23907 7080 23939
rect 7120 23907 7152 23939
rect 7192 23907 7224 23939
rect 7264 23907 7296 23939
rect 7336 23907 7368 23939
rect 7408 23907 7440 23939
rect 7480 23907 7512 23939
rect 7552 23907 7584 23939
rect 7624 23907 7656 23939
rect 7696 23907 7728 23939
rect 7768 23907 7800 23939
rect 7840 23907 7872 23939
rect 7912 23907 7944 23939
rect 7984 23907 8016 23939
rect 8056 23907 8088 23939
rect 8128 23907 8160 23939
rect 8200 23907 8232 23939
rect 8272 23907 8304 23939
rect 8344 23907 8376 23939
rect 8416 23907 8448 23939
rect 8488 23907 8520 23939
rect 8560 23907 8592 23939
rect 8632 23907 8664 23939
rect 8704 23907 8736 23939
rect 8776 23907 8808 23939
rect 8848 23907 8880 23939
rect 8920 23907 8952 23939
rect 8992 23907 9024 23939
rect 9064 23907 9096 23939
rect 9136 23907 9168 23939
rect 9208 23907 9240 23939
rect 9280 23907 9312 23939
rect 9352 23907 9384 23939
rect 9424 23907 9456 23939
rect 9496 23907 9528 23939
rect 9568 23907 9600 23939
rect 9640 23907 9672 23939
rect 9712 23907 9744 23939
rect 9784 23907 9816 23939
rect 9856 23907 9888 23939
rect 9928 23907 9960 23939
rect 10000 23907 10032 23939
rect 10072 23907 10104 23939
rect 10144 23907 10176 23939
rect 10216 23907 10248 23939
rect 10288 23907 10320 23939
rect 10360 23907 10392 23939
rect 10432 23907 10464 23939
rect 10504 23907 10536 23939
rect 10576 23907 10608 23939
rect 10648 23907 10680 23939
rect 10720 23907 10752 23939
rect 10792 23907 10824 23939
rect 10864 23907 10896 23939
rect 10936 23907 10968 23939
rect 11008 23907 11040 23939
rect 11080 23907 11112 23939
rect 11152 23907 11184 23939
rect 11224 23907 11256 23939
rect 11296 23907 11328 23939
rect 11368 23907 11400 23939
rect 11440 23907 11472 23939
rect 11512 23907 11544 23939
rect 11584 23907 11616 23939
rect 11656 23907 11688 23939
rect 11728 23907 11760 23939
rect 11800 23907 11832 23939
rect 11872 23907 11904 23939
rect 11944 23907 11976 23939
rect 12016 23907 12048 23939
rect 12088 23907 12120 23939
rect 12160 23907 12192 23939
rect 12232 23907 12264 23939
rect 12304 23907 12336 23939
rect 12376 23907 12408 23939
rect 12448 23907 12480 23939
rect 12520 23907 12552 23939
rect 12592 23907 12624 23939
rect 12664 23907 12696 23939
rect 12736 23907 12768 23939
rect 12808 23907 12840 23939
rect 12880 23907 12912 23939
rect 12952 23907 12984 23939
rect 13024 23907 13056 23939
rect 13096 23907 13128 23939
rect 13168 23907 13200 23939
rect 13240 23907 13272 23939
rect 13312 23907 13344 23939
rect 13384 23907 13416 23939
rect 13456 23907 13488 23939
rect 13528 23907 13560 23939
rect 13600 23907 13632 23939
rect 13672 23907 13704 23939
rect 13744 23907 13776 23939
rect 13816 23907 13848 23939
rect 13888 23907 13920 23939
rect 13960 23907 13992 23939
rect 14032 23907 14064 23939
rect 14104 23907 14136 23939
rect 14176 23907 14208 23939
rect 14248 23907 14280 23939
rect 14320 23907 14352 23939
rect 14392 23907 14424 23939
rect 14464 23907 14496 23939
rect 14536 23907 14568 23939
rect 14608 23907 14640 23939
rect 14680 23907 14712 23939
rect 14752 23907 14784 23939
rect 14824 23907 14856 23939
rect 14896 23907 14928 23939
rect 14968 23907 15000 23939
rect 15040 23907 15072 23939
rect 15112 23907 15144 23939
rect 15184 23907 15216 23939
rect 15256 23907 15288 23939
rect 15328 23907 15360 23939
rect 15400 23907 15432 23939
rect 15472 23907 15504 23939
rect 15544 23907 15576 23939
rect 15616 23907 15648 23939
rect 15688 23907 15720 23939
rect 15760 23907 15792 23939
rect 15832 23907 15864 23939
rect 15904 23907 15936 23939
rect 64 23835 96 23867
rect 136 23835 168 23867
rect 208 23835 240 23867
rect 280 23835 312 23867
rect 352 23835 384 23867
rect 424 23835 456 23867
rect 496 23835 528 23867
rect 568 23835 600 23867
rect 640 23835 672 23867
rect 712 23835 744 23867
rect 784 23835 816 23867
rect 856 23835 888 23867
rect 928 23835 960 23867
rect 1000 23835 1032 23867
rect 1072 23835 1104 23867
rect 1144 23835 1176 23867
rect 1216 23835 1248 23867
rect 1288 23835 1320 23867
rect 1360 23835 1392 23867
rect 1432 23835 1464 23867
rect 1504 23835 1536 23867
rect 1576 23835 1608 23867
rect 1648 23835 1680 23867
rect 1720 23835 1752 23867
rect 1792 23835 1824 23867
rect 1864 23835 1896 23867
rect 1936 23835 1968 23867
rect 2008 23835 2040 23867
rect 2080 23835 2112 23867
rect 2152 23835 2184 23867
rect 2224 23835 2256 23867
rect 2296 23835 2328 23867
rect 2368 23835 2400 23867
rect 2440 23835 2472 23867
rect 2512 23835 2544 23867
rect 2584 23835 2616 23867
rect 2656 23835 2688 23867
rect 2728 23835 2760 23867
rect 2800 23835 2832 23867
rect 2872 23835 2904 23867
rect 2944 23835 2976 23867
rect 3016 23835 3048 23867
rect 3088 23835 3120 23867
rect 3160 23835 3192 23867
rect 3232 23835 3264 23867
rect 3304 23835 3336 23867
rect 3376 23835 3408 23867
rect 3448 23835 3480 23867
rect 3520 23835 3552 23867
rect 3592 23835 3624 23867
rect 3664 23835 3696 23867
rect 3736 23835 3768 23867
rect 3808 23835 3840 23867
rect 3880 23835 3912 23867
rect 3952 23835 3984 23867
rect 4024 23835 4056 23867
rect 4096 23835 4128 23867
rect 4168 23835 4200 23867
rect 4240 23835 4272 23867
rect 4312 23835 4344 23867
rect 4384 23835 4416 23867
rect 4456 23835 4488 23867
rect 4528 23835 4560 23867
rect 4600 23835 4632 23867
rect 4672 23835 4704 23867
rect 4744 23835 4776 23867
rect 4816 23835 4848 23867
rect 4888 23835 4920 23867
rect 4960 23835 4992 23867
rect 5032 23835 5064 23867
rect 5104 23835 5136 23867
rect 5176 23835 5208 23867
rect 5248 23835 5280 23867
rect 5320 23835 5352 23867
rect 5392 23835 5424 23867
rect 5464 23835 5496 23867
rect 5536 23835 5568 23867
rect 5608 23835 5640 23867
rect 5680 23835 5712 23867
rect 5752 23835 5784 23867
rect 5824 23835 5856 23867
rect 5896 23835 5928 23867
rect 5968 23835 6000 23867
rect 6040 23835 6072 23867
rect 6112 23835 6144 23867
rect 6184 23835 6216 23867
rect 6256 23835 6288 23867
rect 6328 23835 6360 23867
rect 6400 23835 6432 23867
rect 6472 23835 6504 23867
rect 6544 23835 6576 23867
rect 6616 23835 6648 23867
rect 6688 23835 6720 23867
rect 6760 23835 6792 23867
rect 6832 23835 6864 23867
rect 6904 23835 6936 23867
rect 6976 23835 7008 23867
rect 7048 23835 7080 23867
rect 7120 23835 7152 23867
rect 7192 23835 7224 23867
rect 7264 23835 7296 23867
rect 7336 23835 7368 23867
rect 7408 23835 7440 23867
rect 7480 23835 7512 23867
rect 7552 23835 7584 23867
rect 7624 23835 7656 23867
rect 7696 23835 7728 23867
rect 7768 23835 7800 23867
rect 7840 23835 7872 23867
rect 7912 23835 7944 23867
rect 7984 23835 8016 23867
rect 8056 23835 8088 23867
rect 8128 23835 8160 23867
rect 8200 23835 8232 23867
rect 8272 23835 8304 23867
rect 8344 23835 8376 23867
rect 8416 23835 8448 23867
rect 8488 23835 8520 23867
rect 8560 23835 8592 23867
rect 8632 23835 8664 23867
rect 8704 23835 8736 23867
rect 8776 23835 8808 23867
rect 8848 23835 8880 23867
rect 8920 23835 8952 23867
rect 8992 23835 9024 23867
rect 9064 23835 9096 23867
rect 9136 23835 9168 23867
rect 9208 23835 9240 23867
rect 9280 23835 9312 23867
rect 9352 23835 9384 23867
rect 9424 23835 9456 23867
rect 9496 23835 9528 23867
rect 9568 23835 9600 23867
rect 9640 23835 9672 23867
rect 9712 23835 9744 23867
rect 9784 23835 9816 23867
rect 9856 23835 9888 23867
rect 9928 23835 9960 23867
rect 10000 23835 10032 23867
rect 10072 23835 10104 23867
rect 10144 23835 10176 23867
rect 10216 23835 10248 23867
rect 10288 23835 10320 23867
rect 10360 23835 10392 23867
rect 10432 23835 10464 23867
rect 10504 23835 10536 23867
rect 10576 23835 10608 23867
rect 10648 23835 10680 23867
rect 10720 23835 10752 23867
rect 10792 23835 10824 23867
rect 10864 23835 10896 23867
rect 10936 23835 10968 23867
rect 11008 23835 11040 23867
rect 11080 23835 11112 23867
rect 11152 23835 11184 23867
rect 11224 23835 11256 23867
rect 11296 23835 11328 23867
rect 11368 23835 11400 23867
rect 11440 23835 11472 23867
rect 11512 23835 11544 23867
rect 11584 23835 11616 23867
rect 11656 23835 11688 23867
rect 11728 23835 11760 23867
rect 11800 23835 11832 23867
rect 11872 23835 11904 23867
rect 11944 23835 11976 23867
rect 12016 23835 12048 23867
rect 12088 23835 12120 23867
rect 12160 23835 12192 23867
rect 12232 23835 12264 23867
rect 12304 23835 12336 23867
rect 12376 23835 12408 23867
rect 12448 23835 12480 23867
rect 12520 23835 12552 23867
rect 12592 23835 12624 23867
rect 12664 23835 12696 23867
rect 12736 23835 12768 23867
rect 12808 23835 12840 23867
rect 12880 23835 12912 23867
rect 12952 23835 12984 23867
rect 13024 23835 13056 23867
rect 13096 23835 13128 23867
rect 13168 23835 13200 23867
rect 13240 23835 13272 23867
rect 13312 23835 13344 23867
rect 13384 23835 13416 23867
rect 13456 23835 13488 23867
rect 13528 23835 13560 23867
rect 13600 23835 13632 23867
rect 13672 23835 13704 23867
rect 13744 23835 13776 23867
rect 13816 23835 13848 23867
rect 13888 23835 13920 23867
rect 13960 23835 13992 23867
rect 14032 23835 14064 23867
rect 14104 23835 14136 23867
rect 14176 23835 14208 23867
rect 14248 23835 14280 23867
rect 14320 23835 14352 23867
rect 14392 23835 14424 23867
rect 14464 23835 14496 23867
rect 14536 23835 14568 23867
rect 14608 23835 14640 23867
rect 14680 23835 14712 23867
rect 14752 23835 14784 23867
rect 14824 23835 14856 23867
rect 14896 23835 14928 23867
rect 14968 23835 15000 23867
rect 15040 23835 15072 23867
rect 15112 23835 15144 23867
rect 15184 23835 15216 23867
rect 15256 23835 15288 23867
rect 15328 23835 15360 23867
rect 15400 23835 15432 23867
rect 15472 23835 15504 23867
rect 15544 23835 15576 23867
rect 15616 23835 15648 23867
rect 15688 23835 15720 23867
rect 15760 23835 15792 23867
rect 15832 23835 15864 23867
rect 15904 23835 15936 23867
rect 64 23763 96 23795
rect 136 23763 168 23795
rect 208 23763 240 23795
rect 280 23763 312 23795
rect 352 23763 384 23795
rect 424 23763 456 23795
rect 496 23763 528 23795
rect 568 23763 600 23795
rect 640 23763 672 23795
rect 712 23763 744 23795
rect 784 23763 816 23795
rect 856 23763 888 23795
rect 928 23763 960 23795
rect 1000 23763 1032 23795
rect 1072 23763 1104 23795
rect 1144 23763 1176 23795
rect 1216 23763 1248 23795
rect 1288 23763 1320 23795
rect 1360 23763 1392 23795
rect 1432 23763 1464 23795
rect 1504 23763 1536 23795
rect 1576 23763 1608 23795
rect 1648 23763 1680 23795
rect 1720 23763 1752 23795
rect 1792 23763 1824 23795
rect 1864 23763 1896 23795
rect 1936 23763 1968 23795
rect 2008 23763 2040 23795
rect 2080 23763 2112 23795
rect 2152 23763 2184 23795
rect 2224 23763 2256 23795
rect 2296 23763 2328 23795
rect 2368 23763 2400 23795
rect 2440 23763 2472 23795
rect 2512 23763 2544 23795
rect 2584 23763 2616 23795
rect 2656 23763 2688 23795
rect 2728 23763 2760 23795
rect 2800 23763 2832 23795
rect 2872 23763 2904 23795
rect 2944 23763 2976 23795
rect 3016 23763 3048 23795
rect 3088 23763 3120 23795
rect 3160 23763 3192 23795
rect 3232 23763 3264 23795
rect 3304 23763 3336 23795
rect 3376 23763 3408 23795
rect 3448 23763 3480 23795
rect 3520 23763 3552 23795
rect 3592 23763 3624 23795
rect 3664 23763 3696 23795
rect 3736 23763 3768 23795
rect 3808 23763 3840 23795
rect 3880 23763 3912 23795
rect 3952 23763 3984 23795
rect 4024 23763 4056 23795
rect 4096 23763 4128 23795
rect 4168 23763 4200 23795
rect 4240 23763 4272 23795
rect 4312 23763 4344 23795
rect 4384 23763 4416 23795
rect 4456 23763 4488 23795
rect 4528 23763 4560 23795
rect 4600 23763 4632 23795
rect 4672 23763 4704 23795
rect 4744 23763 4776 23795
rect 4816 23763 4848 23795
rect 4888 23763 4920 23795
rect 4960 23763 4992 23795
rect 5032 23763 5064 23795
rect 5104 23763 5136 23795
rect 5176 23763 5208 23795
rect 5248 23763 5280 23795
rect 5320 23763 5352 23795
rect 5392 23763 5424 23795
rect 5464 23763 5496 23795
rect 5536 23763 5568 23795
rect 5608 23763 5640 23795
rect 5680 23763 5712 23795
rect 5752 23763 5784 23795
rect 5824 23763 5856 23795
rect 5896 23763 5928 23795
rect 5968 23763 6000 23795
rect 6040 23763 6072 23795
rect 6112 23763 6144 23795
rect 6184 23763 6216 23795
rect 6256 23763 6288 23795
rect 6328 23763 6360 23795
rect 6400 23763 6432 23795
rect 6472 23763 6504 23795
rect 6544 23763 6576 23795
rect 6616 23763 6648 23795
rect 6688 23763 6720 23795
rect 6760 23763 6792 23795
rect 6832 23763 6864 23795
rect 6904 23763 6936 23795
rect 6976 23763 7008 23795
rect 7048 23763 7080 23795
rect 7120 23763 7152 23795
rect 7192 23763 7224 23795
rect 7264 23763 7296 23795
rect 7336 23763 7368 23795
rect 7408 23763 7440 23795
rect 7480 23763 7512 23795
rect 7552 23763 7584 23795
rect 7624 23763 7656 23795
rect 7696 23763 7728 23795
rect 7768 23763 7800 23795
rect 7840 23763 7872 23795
rect 7912 23763 7944 23795
rect 7984 23763 8016 23795
rect 8056 23763 8088 23795
rect 8128 23763 8160 23795
rect 8200 23763 8232 23795
rect 8272 23763 8304 23795
rect 8344 23763 8376 23795
rect 8416 23763 8448 23795
rect 8488 23763 8520 23795
rect 8560 23763 8592 23795
rect 8632 23763 8664 23795
rect 8704 23763 8736 23795
rect 8776 23763 8808 23795
rect 8848 23763 8880 23795
rect 8920 23763 8952 23795
rect 8992 23763 9024 23795
rect 9064 23763 9096 23795
rect 9136 23763 9168 23795
rect 9208 23763 9240 23795
rect 9280 23763 9312 23795
rect 9352 23763 9384 23795
rect 9424 23763 9456 23795
rect 9496 23763 9528 23795
rect 9568 23763 9600 23795
rect 9640 23763 9672 23795
rect 9712 23763 9744 23795
rect 9784 23763 9816 23795
rect 9856 23763 9888 23795
rect 9928 23763 9960 23795
rect 10000 23763 10032 23795
rect 10072 23763 10104 23795
rect 10144 23763 10176 23795
rect 10216 23763 10248 23795
rect 10288 23763 10320 23795
rect 10360 23763 10392 23795
rect 10432 23763 10464 23795
rect 10504 23763 10536 23795
rect 10576 23763 10608 23795
rect 10648 23763 10680 23795
rect 10720 23763 10752 23795
rect 10792 23763 10824 23795
rect 10864 23763 10896 23795
rect 10936 23763 10968 23795
rect 11008 23763 11040 23795
rect 11080 23763 11112 23795
rect 11152 23763 11184 23795
rect 11224 23763 11256 23795
rect 11296 23763 11328 23795
rect 11368 23763 11400 23795
rect 11440 23763 11472 23795
rect 11512 23763 11544 23795
rect 11584 23763 11616 23795
rect 11656 23763 11688 23795
rect 11728 23763 11760 23795
rect 11800 23763 11832 23795
rect 11872 23763 11904 23795
rect 11944 23763 11976 23795
rect 12016 23763 12048 23795
rect 12088 23763 12120 23795
rect 12160 23763 12192 23795
rect 12232 23763 12264 23795
rect 12304 23763 12336 23795
rect 12376 23763 12408 23795
rect 12448 23763 12480 23795
rect 12520 23763 12552 23795
rect 12592 23763 12624 23795
rect 12664 23763 12696 23795
rect 12736 23763 12768 23795
rect 12808 23763 12840 23795
rect 12880 23763 12912 23795
rect 12952 23763 12984 23795
rect 13024 23763 13056 23795
rect 13096 23763 13128 23795
rect 13168 23763 13200 23795
rect 13240 23763 13272 23795
rect 13312 23763 13344 23795
rect 13384 23763 13416 23795
rect 13456 23763 13488 23795
rect 13528 23763 13560 23795
rect 13600 23763 13632 23795
rect 13672 23763 13704 23795
rect 13744 23763 13776 23795
rect 13816 23763 13848 23795
rect 13888 23763 13920 23795
rect 13960 23763 13992 23795
rect 14032 23763 14064 23795
rect 14104 23763 14136 23795
rect 14176 23763 14208 23795
rect 14248 23763 14280 23795
rect 14320 23763 14352 23795
rect 14392 23763 14424 23795
rect 14464 23763 14496 23795
rect 14536 23763 14568 23795
rect 14608 23763 14640 23795
rect 14680 23763 14712 23795
rect 14752 23763 14784 23795
rect 14824 23763 14856 23795
rect 14896 23763 14928 23795
rect 14968 23763 15000 23795
rect 15040 23763 15072 23795
rect 15112 23763 15144 23795
rect 15184 23763 15216 23795
rect 15256 23763 15288 23795
rect 15328 23763 15360 23795
rect 15400 23763 15432 23795
rect 15472 23763 15504 23795
rect 15544 23763 15576 23795
rect 15616 23763 15648 23795
rect 15688 23763 15720 23795
rect 15760 23763 15792 23795
rect 15832 23763 15864 23795
rect 15904 23763 15936 23795
rect 64 23691 96 23723
rect 136 23691 168 23723
rect 208 23691 240 23723
rect 280 23691 312 23723
rect 352 23691 384 23723
rect 424 23691 456 23723
rect 496 23691 528 23723
rect 568 23691 600 23723
rect 640 23691 672 23723
rect 712 23691 744 23723
rect 784 23691 816 23723
rect 856 23691 888 23723
rect 928 23691 960 23723
rect 1000 23691 1032 23723
rect 1072 23691 1104 23723
rect 1144 23691 1176 23723
rect 1216 23691 1248 23723
rect 1288 23691 1320 23723
rect 1360 23691 1392 23723
rect 1432 23691 1464 23723
rect 1504 23691 1536 23723
rect 1576 23691 1608 23723
rect 1648 23691 1680 23723
rect 1720 23691 1752 23723
rect 1792 23691 1824 23723
rect 1864 23691 1896 23723
rect 1936 23691 1968 23723
rect 2008 23691 2040 23723
rect 2080 23691 2112 23723
rect 2152 23691 2184 23723
rect 2224 23691 2256 23723
rect 2296 23691 2328 23723
rect 2368 23691 2400 23723
rect 2440 23691 2472 23723
rect 2512 23691 2544 23723
rect 2584 23691 2616 23723
rect 2656 23691 2688 23723
rect 2728 23691 2760 23723
rect 2800 23691 2832 23723
rect 2872 23691 2904 23723
rect 2944 23691 2976 23723
rect 3016 23691 3048 23723
rect 3088 23691 3120 23723
rect 3160 23691 3192 23723
rect 3232 23691 3264 23723
rect 3304 23691 3336 23723
rect 3376 23691 3408 23723
rect 3448 23691 3480 23723
rect 3520 23691 3552 23723
rect 3592 23691 3624 23723
rect 3664 23691 3696 23723
rect 3736 23691 3768 23723
rect 3808 23691 3840 23723
rect 3880 23691 3912 23723
rect 3952 23691 3984 23723
rect 4024 23691 4056 23723
rect 4096 23691 4128 23723
rect 4168 23691 4200 23723
rect 4240 23691 4272 23723
rect 4312 23691 4344 23723
rect 4384 23691 4416 23723
rect 4456 23691 4488 23723
rect 4528 23691 4560 23723
rect 4600 23691 4632 23723
rect 4672 23691 4704 23723
rect 4744 23691 4776 23723
rect 4816 23691 4848 23723
rect 4888 23691 4920 23723
rect 4960 23691 4992 23723
rect 5032 23691 5064 23723
rect 5104 23691 5136 23723
rect 5176 23691 5208 23723
rect 5248 23691 5280 23723
rect 5320 23691 5352 23723
rect 5392 23691 5424 23723
rect 5464 23691 5496 23723
rect 5536 23691 5568 23723
rect 5608 23691 5640 23723
rect 5680 23691 5712 23723
rect 5752 23691 5784 23723
rect 5824 23691 5856 23723
rect 5896 23691 5928 23723
rect 5968 23691 6000 23723
rect 6040 23691 6072 23723
rect 6112 23691 6144 23723
rect 6184 23691 6216 23723
rect 6256 23691 6288 23723
rect 6328 23691 6360 23723
rect 6400 23691 6432 23723
rect 6472 23691 6504 23723
rect 6544 23691 6576 23723
rect 6616 23691 6648 23723
rect 6688 23691 6720 23723
rect 6760 23691 6792 23723
rect 6832 23691 6864 23723
rect 6904 23691 6936 23723
rect 6976 23691 7008 23723
rect 7048 23691 7080 23723
rect 7120 23691 7152 23723
rect 7192 23691 7224 23723
rect 7264 23691 7296 23723
rect 7336 23691 7368 23723
rect 7408 23691 7440 23723
rect 7480 23691 7512 23723
rect 7552 23691 7584 23723
rect 7624 23691 7656 23723
rect 7696 23691 7728 23723
rect 7768 23691 7800 23723
rect 7840 23691 7872 23723
rect 7912 23691 7944 23723
rect 7984 23691 8016 23723
rect 8056 23691 8088 23723
rect 8128 23691 8160 23723
rect 8200 23691 8232 23723
rect 8272 23691 8304 23723
rect 8344 23691 8376 23723
rect 8416 23691 8448 23723
rect 8488 23691 8520 23723
rect 8560 23691 8592 23723
rect 8632 23691 8664 23723
rect 8704 23691 8736 23723
rect 8776 23691 8808 23723
rect 8848 23691 8880 23723
rect 8920 23691 8952 23723
rect 8992 23691 9024 23723
rect 9064 23691 9096 23723
rect 9136 23691 9168 23723
rect 9208 23691 9240 23723
rect 9280 23691 9312 23723
rect 9352 23691 9384 23723
rect 9424 23691 9456 23723
rect 9496 23691 9528 23723
rect 9568 23691 9600 23723
rect 9640 23691 9672 23723
rect 9712 23691 9744 23723
rect 9784 23691 9816 23723
rect 9856 23691 9888 23723
rect 9928 23691 9960 23723
rect 10000 23691 10032 23723
rect 10072 23691 10104 23723
rect 10144 23691 10176 23723
rect 10216 23691 10248 23723
rect 10288 23691 10320 23723
rect 10360 23691 10392 23723
rect 10432 23691 10464 23723
rect 10504 23691 10536 23723
rect 10576 23691 10608 23723
rect 10648 23691 10680 23723
rect 10720 23691 10752 23723
rect 10792 23691 10824 23723
rect 10864 23691 10896 23723
rect 10936 23691 10968 23723
rect 11008 23691 11040 23723
rect 11080 23691 11112 23723
rect 11152 23691 11184 23723
rect 11224 23691 11256 23723
rect 11296 23691 11328 23723
rect 11368 23691 11400 23723
rect 11440 23691 11472 23723
rect 11512 23691 11544 23723
rect 11584 23691 11616 23723
rect 11656 23691 11688 23723
rect 11728 23691 11760 23723
rect 11800 23691 11832 23723
rect 11872 23691 11904 23723
rect 11944 23691 11976 23723
rect 12016 23691 12048 23723
rect 12088 23691 12120 23723
rect 12160 23691 12192 23723
rect 12232 23691 12264 23723
rect 12304 23691 12336 23723
rect 12376 23691 12408 23723
rect 12448 23691 12480 23723
rect 12520 23691 12552 23723
rect 12592 23691 12624 23723
rect 12664 23691 12696 23723
rect 12736 23691 12768 23723
rect 12808 23691 12840 23723
rect 12880 23691 12912 23723
rect 12952 23691 12984 23723
rect 13024 23691 13056 23723
rect 13096 23691 13128 23723
rect 13168 23691 13200 23723
rect 13240 23691 13272 23723
rect 13312 23691 13344 23723
rect 13384 23691 13416 23723
rect 13456 23691 13488 23723
rect 13528 23691 13560 23723
rect 13600 23691 13632 23723
rect 13672 23691 13704 23723
rect 13744 23691 13776 23723
rect 13816 23691 13848 23723
rect 13888 23691 13920 23723
rect 13960 23691 13992 23723
rect 14032 23691 14064 23723
rect 14104 23691 14136 23723
rect 14176 23691 14208 23723
rect 14248 23691 14280 23723
rect 14320 23691 14352 23723
rect 14392 23691 14424 23723
rect 14464 23691 14496 23723
rect 14536 23691 14568 23723
rect 14608 23691 14640 23723
rect 14680 23691 14712 23723
rect 14752 23691 14784 23723
rect 14824 23691 14856 23723
rect 14896 23691 14928 23723
rect 14968 23691 15000 23723
rect 15040 23691 15072 23723
rect 15112 23691 15144 23723
rect 15184 23691 15216 23723
rect 15256 23691 15288 23723
rect 15328 23691 15360 23723
rect 15400 23691 15432 23723
rect 15472 23691 15504 23723
rect 15544 23691 15576 23723
rect 15616 23691 15648 23723
rect 15688 23691 15720 23723
rect 15760 23691 15792 23723
rect 15832 23691 15864 23723
rect 15904 23691 15936 23723
rect 64 23619 96 23651
rect 136 23619 168 23651
rect 208 23619 240 23651
rect 280 23619 312 23651
rect 352 23619 384 23651
rect 424 23619 456 23651
rect 496 23619 528 23651
rect 568 23619 600 23651
rect 640 23619 672 23651
rect 712 23619 744 23651
rect 784 23619 816 23651
rect 856 23619 888 23651
rect 928 23619 960 23651
rect 1000 23619 1032 23651
rect 1072 23619 1104 23651
rect 1144 23619 1176 23651
rect 1216 23619 1248 23651
rect 1288 23619 1320 23651
rect 1360 23619 1392 23651
rect 1432 23619 1464 23651
rect 1504 23619 1536 23651
rect 1576 23619 1608 23651
rect 1648 23619 1680 23651
rect 1720 23619 1752 23651
rect 1792 23619 1824 23651
rect 1864 23619 1896 23651
rect 1936 23619 1968 23651
rect 2008 23619 2040 23651
rect 2080 23619 2112 23651
rect 2152 23619 2184 23651
rect 2224 23619 2256 23651
rect 2296 23619 2328 23651
rect 2368 23619 2400 23651
rect 2440 23619 2472 23651
rect 2512 23619 2544 23651
rect 2584 23619 2616 23651
rect 2656 23619 2688 23651
rect 2728 23619 2760 23651
rect 2800 23619 2832 23651
rect 2872 23619 2904 23651
rect 2944 23619 2976 23651
rect 3016 23619 3048 23651
rect 3088 23619 3120 23651
rect 3160 23619 3192 23651
rect 3232 23619 3264 23651
rect 3304 23619 3336 23651
rect 3376 23619 3408 23651
rect 3448 23619 3480 23651
rect 3520 23619 3552 23651
rect 3592 23619 3624 23651
rect 3664 23619 3696 23651
rect 3736 23619 3768 23651
rect 3808 23619 3840 23651
rect 3880 23619 3912 23651
rect 3952 23619 3984 23651
rect 4024 23619 4056 23651
rect 4096 23619 4128 23651
rect 4168 23619 4200 23651
rect 4240 23619 4272 23651
rect 4312 23619 4344 23651
rect 4384 23619 4416 23651
rect 4456 23619 4488 23651
rect 4528 23619 4560 23651
rect 4600 23619 4632 23651
rect 4672 23619 4704 23651
rect 4744 23619 4776 23651
rect 4816 23619 4848 23651
rect 4888 23619 4920 23651
rect 4960 23619 4992 23651
rect 5032 23619 5064 23651
rect 5104 23619 5136 23651
rect 5176 23619 5208 23651
rect 5248 23619 5280 23651
rect 5320 23619 5352 23651
rect 5392 23619 5424 23651
rect 5464 23619 5496 23651
rect 5536 23619 5568 23651
rect 5608 23619 5640 23651
rect 5680 23619 5712 23651
rect 5752 23619 5784 23651
rect 5824 23619 5856 23651
rect 5896 23619 5928 23651
rect 5968 23619 6000 23651
rect 6040 23619 6072 23651
rect 6112 23619 6144 23651
rect 6184 23619 6216 23651
rect 6256 23619 6288 23651
rect 6328 23619 6360 23651
rect 6400 23619 6432 23651
rect 6472 23619 6504 23651
rect 6544 23619 6576 23651
rect 6616 23619 6648 23651
rect 6688 23619 6720 23651
rect 6760 23619 6792 23651
rect 6832 23619 6864 23651
rect 6904 23619 6936 23651
rect 6976 23619 7008 23651
rect 7048 23619 7080 23651
rect 7120 23619 7152 23651
rect 7192 23619 7224 23651
rect 7264 23619 7296 23651
rect 7336 23619 7368 23651
rect 7408 23619 7440 23651
rect 7480 23619 7512 23651
rect 7552 23619 7584 23651
rect 7624 23619 7656 23651
rect 7696 23619 7728 23651
rect 7768 23619 7800 23651
rect 7840 23619 7872 23651
rect 7912 23619 7944 23651
rect 7984 23619 8016 23651
rect 8056 23619 8088 23651
rect 8128 23619 8160 23651
rect 8200 23619 8232 23651
rect 8272 23619 8304 23651
rect 8344 23619 8376 23651
rect 8416 23619 8448 23651
rect 8488 23619 8520 23651
rect 8560 23619 8592 23651
rect 8632 23619 8664 23651
rect 8704 23619 8736 23651
rect 8776 23619 8808 23651
rect 8848 23619 8880 23651
rect 8920 23619 8952 23651
rect 8992 23619 9024 23651
rect 9064 23619 9096 23651
rect 9136 23619 9168 23651
rect 9208 23619 9240 23651
rect 9280 23619 9312 23651
rect 9352 23619 9384 23651
rect 9424 23619 9456 23651
rect 9496 23619 9528 23651
rect 9568 23619 9600 23651
rect 9640 23619 9672 23651
rect 9712 23619 9744 23651
rect 9784 23619 9816 23651
rect 9856 23619 9888 23651
rect 9928 23619 9960 23651
rect 10000 23619 10032 23651
rect 10072 23619 10104 23651
rect 10144 23619 10176 23651
rect 10216 23619 10248 23651
rect 10288 23619 10320 23651
rect 10360 23619 10392 23651
rect 10432 23619 10464 23651
rect 10504 23619 10536 23651
rect 10576 23619 10608 23651
rect 10648 23619 10680 23651
rect 10720 23619 10752 23651
rect 10792 23619 10824 23651
rect 10864 23619 10896 23651
rect 10936 23619 10968 23651
rect 11008 23619 11040 23651
rect 11080 23619 11112 23651
rect 11152 23619 11184 23651
rect 11224 23619 11256 23651
rect 11296 23619 11328 23651
rect 11368 23619 11400 23651
rect 11440 23619 11472 23651
rect 11512 23619 11544 23651
rect 11584 23619 11616 23651
rect 11656 23619 11688 23651
rect 11728 23619 11760 23651
rect 11800 23619 11832 23651
rect 11872 23619 11904 23651
rect 11944 23619 11976 23651
rect 12016 23619 12048 23651
rect 12088 23619 12120 23651
rect 12160 23619 12192 23651
rect 12232 23619 12264 23651
rect 12304 23619 12336 23651
rect 12376 23619 12408 23651
rect 12448 23619 12480 23651
rect 12520 23619 12552 23651
rect 12592 23619 12624 23651
rect 12664 23619 12696 23651
rect 12736 23619 12768 23651
rect 12808 23619 12840 23651
rect 12880 23619 12912 23651
rect 12952 23619 12984 23651
rect 13024 23619 13056 23651
rect 13096 23619 13128 23651
rect 13168 23619 13200 23651
rect 13240 23619 13272 23651
rect 13312 23619 13344 23651
rect 13384 23619 13416 23651
rect 13456 23619 13488 23651
rect 13528 23619 13560 23651
rect 13600 23619 13632 23651
rect 13672 23619 13704 23651
rect 13744 23619 13776 23651
rect 13816 23619 13848 23651
rect 13888 23619 13920 23651
rect 13960 23619 13992 23651
rect 14032 23619 14064 23651
rect 14104 23619 14136 23651
rect 14176 23619 14208 23651
rect 14248 23619 14280 23651
rect 14320 23619 14352 23651
rect 14392 23619 14424 23651
rect 14464 23619 14496 23651
rect 14536 23619 14568 23651
rect 14608 23619 14640 23651
rect 14680 23619 14712 23651
rect 14752 23619 14784 23651
rect 14824 23619 14856 23651
rect 14896 23619 14928 23651
rect 14968 23619 15000 23651
rect 15040 23619 15072 23651
rect 15112 23619 15144 23651
rect 15184 23619 15216 23651
rect 15256 23619 15288 23651
rect 15328 23619 15360 23651
rect 15400 23619 15432 23651
rect 15472 23619 15504 23651
rect 15544 23619 15576 23651
rect 15616 23619 15648 23651
rect 15688 23619 15720 23651
rect 15760 23619 15792 23651
rect 15832 23619 15864 23651
rect 15904 23619 15936 23651
rect 64 23547 96 23579
rect 136 23547 168 23579
rect 208 23547 240 23579
rect 280 23547 312 23579
rect 352 23547 384 23579
rect 424 23547 456 23579
rect 496 23547 528 23579
rect 568 23547 600 23579
rect 640 23547 672 23579
rect 712 23547 744 23579
rect 784 23547 816 23579
rect 856 23547 888 23579
rect 928 23547 960 23579
rect 1000 23547 1032 23579
rect 1072 23547 1104 23579
rect 1144 23547 1176 23579
rect 1216 23547 1248 23579
rect 1288 23547 1320 23579
rect 1360 23547 1392 23579
rect 1432 23547 1464 23579
rect 1504 23547 1536 23579
rect 1576 23547 1608 23579
rect 1648 23547 1680 23579
rect 1720 23547 1752 23579
rect 1792 23547 1824 23579
rect 1864 23547 1896 23579
rect 1936 23547 1968 23579
rect 2008 23547 2040 23579
rect 2080 23547 2112 23579
rect 2152 23547 2184 23579
rect 2224 23547 2256 23579
rect 2296 23547 2328 23579
rect 2368 23547 2400 23579
rect 2440 23547 2472 23579
rect 2512 23547 2544 23579
rect 2584 23547 2616 23579
rect 2656 23547 2688 23579
rect 2728 23547 2760 23579
rect 2800 23547 2832 23579
rect 2872 23547 2904 23579
rect 2944 23547 2976 23579
rect 3016 23547 3048 23579
rect 3088 23547 3120 23579
rect 3160 23547 3192 23579
rect 3232 23547 3264 23579
rect 3304 23547 3336 23579
rect 3376 23547 3408 23579
rect 3448 23547 3480 23579
rect 3520 23547 3552 23579
rect 3592 23547 3624 23579
rect 3664 23547 3696 23579
rect 3736 23547 3768 23579
rect 3808 23547 3840 23579
rect 3880 23547 3912 23579
rect 3952 23547 3984 23579
rect 4024 23547 4056 23579
rect 4096 23547 4128 23579
rect 4168 23547 4200 23579
rect 4240 23547 4272 23579
rect 4312 23547 4344 23579
rect 4384 23547 4416 23579
rect 4456 23547 4488 23579
rect 4528 23547 4560 23579
rect 4600 23547 4632 23579
rect 4672 23547 4704 23579
rect 4744 23547 4776 23579
rect 4816 23547 4848 23579
rect 4888 23547 4920 23579
rect 4960 23547 4992 23579
rect 5032 23547 5064 23579
rect 5104 23547 5136 23579
rect 5176 23547 5208 23579
rect 5248 23547 5280 23579
rect 5320 23547 5352 23579
rect 5392 23547 5424 23579
rect 5464 23547 5496 23579
rect 5536 23547 5568 23579
rect 5608 23547 5640 23579
rect 5680 23547 5712 23579
rect 5752 23547 5784 23579
rect 5824 23547 5856 23579
rect 5896 23547 5928 23579
rect 5968 23547 6000 23579
rect 6040 23547 6072 23579
rect 6112 23547 6144 23579
rect 6184 23547 6216 23579
rect 6256 23547 6288 23579
rect 6328 23547 6360 23579
rect 6400 23547 6432 23579
rect 6472 23547 6504 23579
rect 6544 23547 6576 23579
rect 6616 23547 6648 23579
rect 6688 23547 6720 23579
rect 6760 23547 6792 23579
rect 6832 23547 6864 23579
rect 6904 23547 6936 23579
rect 6976 23547 7008 23579
rect 7048 23547 7080 23579
rect 7120 23547 7152 23579
rect 7192 23547 7224 23579
rect 7264 23547 7296 23579
rect 7336 23547 7368 23579
rect 7408 23547 7440 23579
rect 7480 23547 7512 23579
rect 7552 23547 7584 23579
rect 7624 23547 7656 23579
rect 7696 23547 7728 23579
rect 7768 23547 7800 23579
rect 7840 23547 7872 23579
rect 7912 23547 7944 23579
rect 7984 23547 8016 23579
rect 8056 23547 8088 23579
rect 8128 23547 8160 23579
rect 8200 23547 8232 23579
rect 8272 23547 8304 23579
rect 8344 23547 8376 23579
rect 8416 23547 8448 23579
rect 8488 23547 8520 23579
rect 8560 23547 8592 23579
rect 8632 23547 8664 23579
rect 8704 23547 8736 23579
rect 8776 23547 8808 23579
rect 8848 23547 8880 23579
rect 8920 23547 8952 23579
rect 8992 23547 9024 23579
rect 9064 23547 9096 23579
rect 9136 23547 9168 23579
rect 9208 23547 9240 23579
rect 9280 23547 9312 23579
rect 9352 23547 9384 23579
rect 9424 23547 9456 23579
rect 9496 23547 9528 23579
rect 9568 23547 9600 23579
rect 9640 23547 9672 23579
rect 9712 23547 9744 23579
rect 9784 23547 9816 23579
rect 9856 23547 9888 23579
rect 9928 23547 9960 23579
rect 10000 23547 10032 23579
rect 10072 23547 10104 23579
rect 10144 23547 10176 23579
rect 10216 23547 10248 23579
rect 10288 23547 10320 23579
rect 10360 23547 10392 23579
rect 10432 23547 10464 23579
rect 10504 23547 10536 23579
rect 10576 23547 10608 23579
rect 10648 23547 10680 23579
rect 10720 23547 10752 23579
rect 10792 23547 10824 23579
rect 10864 23547 10896 23579
rect 10936 23547 10968 23579
rect 11008 23547 11040 23579
rect 11080 23547 11112 23579
rect 11152 23547 11184 23579
rect 11224 23547 11256 23579
rect 11296 23547 11328 23579
rect 11368 23547 11400 23579
rect 11440 23547 11472 23579
rect 11512 23547 11544 23579
rect 11584 23547 11616 23579
rect 11656 23547 11688 23579
rect 11728 23547 11760 23579
rect 11800 23547 11832 23579
rect 11872 23547 11904 23579
rect 11944 23547 11976 23579
rect 12016 23547 12048 23579
rect 12088 23547 12120 23579
rect 12160 23547 12192 23579
rect 12232 23547 12264 23579
rect 12304 23547 12336 23579
rect 12376 23547 12408 23579
rect 12448 23547 12480 23579
rect 12520 23547 12552 23579
rect 12592 23547 12624 23579
rect 12664 23547 12696 23579
rect 12736 23547 12768 23579
rect 12808 23547 12840 23579
rect 12880 23547 12912 23579
rect 12952 23547 12984 23579
rect 13024 23547 13056 23579
rect 13096 23547 13128 23579
rect 13168 23547 13200 23579
rect 13240 23547 13272 23579
rect 13312 23547 13344 23579
rect 13384 23547 13416 23579
rect 13456 23547 13488 23579
rect 13528 23547 13560 23579
rect 13600 23547 13632 23579
rect 13672 23547 13704 23579
rect 13744 23547 13776 23579
rect 13816 23547 13848 23579
rect 13888 23547 13920 23579
rect 13960 23547 13992 23579
rect 14032 23547 14064 23579
rect 14104 23547 14136 23579
rect 14176 23547 14208 23579
rect 14248 23547 14280 23579
rect 14320 23547 14352 23579
rect 14392 23547 14424 23579
rect 14464 23547 14496 23579
rect 14536 23547 14568 23579
rect 14608 23547 14640 23579
rect 14680 23547 14712 23579
rect 14752 23547 14784 23579
rect 14824 23547 14856 23579
rect 14896 23547 14928 23579
rect 14968 23547 15000 23579
rect 15040 23547 15072 23579
rect 15112 23547 15144 23579
rect 15184 23547 15216 23579
rect 15256 23547 15288 23579
rect 15328 23547 15360 23579
rect 15400 23547 15432 23579
rect 15472 23547 15504 23579
rect 15544 23547 15576 23579
rect 15616 23547 15648 23579
rect 15688 23547 15720 23579
rect 15760 23547 15792 23579
rect 15832 23547 15864 23579
rect 15904 23547 15936 23579
rect 64 23475 96 23507
rect 136 23475 168 23507
rect 208 23475 240 23507
rect 280 23475 312 23507
rect 352 23475 384 23507
rect 424 23475 456 23507
rect 496 23475 528 23507
rect 568 23475 600 23507
rect 640 23475 672 23507
rect 712 23475 744 23507
rect 784 23475 816 23507
rect 856 23475 888 23507
rect 928 23475 960 23507
rect 1000 23475 1032 23507
rect 1072 23475 1104 23507
rect 1144 23475 1176 23507
rect 1216 23475 1248 23507
rect 1288 23475 1320 23507
rect 1360 23475 1392 23507
rect 1432 23475 1464 23507
rect 1504 23475 1536 23507
rect 1576 23475 1608 23507
rect 1648 23475 1680 23507
rect 1720 23475 1752 23507
rect 1792 23475 1824 23507
rect 1864 23475 1896 23507
rect 1936 23475 1968 23507
rect 2008 23475 2040 23507
rect 2080 23475 2112 23507
rect 2152 23475 2184 23507
rect 2224 23475 2256 23507
rect 2296 23475 2328 23507
rect 2368 23475 2400 23507
rect 2440 23475 2472 23507
rect 2512 23475 2544 23507
rect 2584 23475 2616 23507
rect 2656 23475 2688 23507
rect 2728 23475 2760 23507
rect 2800 23475 2832 23507
rect 2872 23475 2904 23507
rect 2944 23475 2976 23507
rect 3016 23475 3048 23507
rect 3088 23475 3120 23507
rect 3160 23475 3192 23507
rect 3232 23475 3264 23507
rect 3304 23475 3336 23507
rect 3376 23475 3408 23507
rect 3448 23475 3480 23507
rect 3520 23475 3552 23507
rect 3592 23475 3624 23507
rect 3664 23475 3696 23507
rect 3736 23475 3768 23507
rect 3808 23475 3840 23507
rect 3880 23475 3912 23507
rect 3952 23475 3984 23507
rect 4024 23475 4056 23507
rect 4096 23475 4128 23507
rect 4168 23475 4200 23507
rect 4240 23475 4272 23507
rect 4312 23475 4344 23507
rect 4384 23475 4416 23507
rect 4456 23475 4488 23507
rect 4528 23475 4560 23507
rect 4600 23475 4632 23507
rect 4672 23475 4704 23507
rect 4744 23475 4776 23507
rect 4816 23475 4848 23507
rect 4888 23475 4920 23507
rect 4960 23475 4992 23507
rect 5032 23475 5064 23507
rect 5104 23475 5136 23507
rect 5176 23475 5208 23507
rect 5248 23475 5280 23507
rect 5320 23475 5352 23507
rect 5392 23475 5424 23507
rect 5464 23475 5496 23507
rect 5536 23475 5568 23507
rect 5608 23475 5640 23507
rect 5680 23475 5712 23507
rect 5752 23475 5784 23507
rect 5824 23475 5856 23507
rect 5896 23475 5928 23507
rect 5968 23475 6000 23507
rect 6040 23475 6072 23507
rect 6112 23475 6144 23507
rect 6184 23475 6216 23507
rect 6256 23475 6288 23507
rect 6328 23475 6360 23507
rect 6400 23475 6432 23507
rect 6472 23475 6504 23507
rect 6544 23475 6576 23507
rect 6616 23475 6648 23507
rect 6688 23475 6720 23507
rect 6760 23475 6792 23507
rect 6832 23475 6864 23507
rect 6904 23475 6936 23507
rect 6976 23475 7008 23507
rect 7048 23475 7080 23507
rect 7120 23475 7152 23507
rect 7192 23475 7224 23507
rect 7264 23475 7296 23507
rect 7336 23475 7368 23507
rect 7408 23475 7440 23507
rect 7480 23475 7512 23507
rect 7552 23475 7584 23507
rect 7624 23475 7656 23507
rect 7696 23475 7728 23507
rect 7768 23475 7800 23507
rect 7840 23475 7872 23507
rect 7912 23475 7944 23507
rect 7984 23475 8016 23507
rect 8056 23475 8088 23507
rect 8128 23475 8160 23507
rect 8200 23475 8232 23507
rect 8272 23475 8304 23507
rect 8344 23475 8376 23507
rect 8416 23475 8448 23507
rect 8488 23475 8520 23507
rect 8560 23475 8592 23507
rect 8632 23475 8664 23507
rect 8704 23475 8736 23507
rect 8776 23475 8808 23507
rect 8848 23475 8880 23507
rect 8920 23475 8952 23507
rect 8992 23475 9024 23507
rect 9064 23475 9096 23507
rect 9136 23475 9168 23507
rect 9208 23475 9240 23507
rect 9280 23475 9312 23507
rect 9352 23475 9384 23507
rect 9424 23475 9456 23507
rect 9496 23475 9528 23507
rect 9568 23475 9600 23507
rect 9640 23475 9672 23507
rect 9712 23475 9744 23507
rect 9784 23475 9816 23507
rect 9856 23475 9888 23507
rect 9928 23475 9960 23507
rect 10000 23475 10032 23507
rect 10072 23475 10104 23507
rect 10144 23475 10176 23507
rect 10216 23475 10248 23507
rect 10288 23475 10320 23507
rect 10360 23475 10392 23507
rect 10432 23475 10464 23507
rect 10504 23475 10536 23507
rect 10576 23475 10608 23507
rect 10648 23475 10680 23507
rect 10720 23475 10752 23507
rect 10792 23475 10824 23507
rect 10864 23475 10896 23507
rect 10936 23475 10968 23507
rect 11008 23475 11040 23507
rect 11080 23475 11112 23507
rect 11152 23475 11184 23507
rect 11224 23475 11256 23507
rect 11296 23475 11328 23507
rect 11368 23475 11400 23507
rect 11440 23475 11472 23507
rect 11512 23475 11544 23507
rect 11584 23475 11616 23507
rect 11656 23475 11688 23507
rect 11728 23475 11760 23507
rect 11800 23475 11832 23507
rect 11872 23475 11904 23507
rect 11944 23475 11976 23507
rect 12016 23475 12048 23507
rect 12088 23475 12120 23507
rect 12160 23475 12192 23507
rect 12232 23475 12264 23507
rect 12304 23475 12336 23507
rect 12376 23475 12408 23507
rect 12448 23475 12480 23507
rect 12520 23475 12552 23507
rect 12592 23475 12624 23507
rect 12664 23475 12696 23507
rect 12736 23475 12768 23507
rect 12808 23475 12840 23507
rect 12880 23475 12912 23507
rect 12952 23475 12984 23507
rect 13024 23475 13056 23507
rect 13096 23475 13128 23507
rect 13168 23475 13200 23507
rect 13240 23475 13272 23507
rect 13312 23475 13344 23507
rect 13384 23475 13416 23507
rect 13456 23475 13488 23507
rect 13528 23475 13560 23507
rect 13600 23475 13632 23507
rect 13672 23475 13704 23507
rect 13744 23475 13776 23507
rect 13816 23475 13848 23507
rect 13888 23475 13920 23507
rect 13960 23475 13992 23507
rect 14032 23475 14064 23507
rect 14104 23475 14136 23507
rect 14176 23475 14208 23507
rect 14248 23475 14280 23507
rect 14320 23475 14352 23507
rect 14392 23475 14424 23507
rect 14464 23475 14496 23507
rect 14536 23475 14568 23507
rect 14608 23475 14640 23507
rect 14680 23475 14712 23507
rect 14752 23475 14784 23507
rect 14824 23475 14856 23507
rect 14896 23475 14928 23507
rect 14968 23475 15000 23507
rect 15040 23475 15072 23507
rect 15112 23475 15144 23507
rect 15184 23475 15216 23507
rect 15256 23475 15288 23507
rect 15328 23475 15360 23507
rect 15400 23475 15432 23507
rect 15472 23475 15504 23507
rect 15544 23475 15576 23507
rect 15616 23475 15648 23507
rect 15688 23475 15720 23507
rect 15760 23475 15792 23507
rect 15832 23475 15864 23507
rect 15904 23475 15936 23507
rect 64 23403 96 23435
rect 136 23403 168 23435
rect 208 23403 240 23435
rect 280 23403 312 23435
rect 352 23403 384 23435
rect 424 23403 456 23435
rect 496 23403 528 23435
rect 568 23403 600 23435
rect 640 23403 672 23435
rect 712 23403 744 23435
rect 784 23403 816 23435
rect 856 23403 888 23435
rect 928 23403 960 23435
rect 1000 23403 1032 23435
rect 1072 23403 1104 23435
rect 1144 23403 1176 23435
rect 1216 23403 1248 23435
rect 1288 23403 1320 23435
rect 1360 23403 1392 23435
rect 1432 23403 1464 23435
rect 1504 23403 1536 23435
rect 1576 23403 1608 23435
rect 1648 23403 1680 23435
rect 1720 23403 1752 23435
rect 1792 23403 1824 23435
rect 1864 23403 1896 23435
rect 1936 23403 1968 23435
rect 2008 23403 2040 23435
rect 2080 23403 2112 23435
rect 2152 23403 2184 23435
rect 2224 23403 2256 23435
rect 2296 23403 2328 23435
rect 2368 23403 2400 23435
rect 2440 23403 2472 23435
rect 2512 23403 2544 23435
rect 2584 23403 2616 23435
rect 2656 23403 2688 23435
rect 2728 23403 2760 23435
rect 2800 23403 2832 23435
rect 2872 23403 2904 23435
rect 2944 23403 2976 23435
rect 3016 23403 3048 23435
rect 3088 23403 3120 23435
rect 3160 23403 3192 23435
rect 3232 23403 3264 23435
rect 3304 23403 3336 23435
rect 3376 23403 3408 23435
rect 3448 23403 3480 23435
rect 3520 23403 3552 23435
rect 3592 23403 3624 23435
rect 3664 23403 3696 23435
rect 3736 23403 3768 23435
rect 3808 23403 3840 23435
rect 3880 23403 3912 23435
rect 3952 23403 3984 23435
rect 4024 23403 4056 23435
rect 4096 23403 4128 23435
rect 4168 23403 4200 23435
rect 4240 23403 4272 23435
rect 4312 23403 4344 23435
rect 4384 23403 4416 23435
rect 4456 23403 4488 23435
rect 4528 23403 4560 23435
rect 4600 23403 4632 23435
rect 4672 23403 4704 23435
rect 4744 23403 4776 23435
rect 4816 23403 4848 23435
rect 4888 23403 4920 23435
rect 4960 23403 4992 23435
rect 5032 23403 5064 23435
rect 5104 23403 5136 23435
rect 5176 23403 5208 23435
rect 5248 23403 5280 23435
rect 5320 23403 5352 23435
rect 5392 23403 5424 23435
rect 5464 23403 5496 23435
rect 5536 23403 5568 23435
rect 5608 23403 5640 23435
rect 5680 23403 5712 23435
rect 5752 23403 5784 23435
rect 5824 23403 5856 23435
rect 5896 23403 5928 23435
rect 5968 23403 6000 23435
rect 6040 23403 6072 23435
rect 6112 23403 6144 23435
rect 6184 23403 6216 23435
rect 6256 23403 6288 23435
rect 6328 23403 6360 23435
rect 6400 23403 6432 23435
rect 6472 23403 6504 23435
rect 6544 23403 6576 23435
rect 6616 23403 6648 23435
rect 6688 23403 6720 23435
rect 6760 23403 6792 23435
rect 6832 23403 6864 23435
rect 6904 23403 6936 23435
rect 6976 23403 7008 23435
rect 7048 23403 7080 23435
rect 7120 23403 7152 23435
rect 7192 23403 7224 23435
rect 7264 23403 7296 23435
rect 7336 23403 7368 23435
rect 7408 23403 7440 23435
rect 7480 23403 7512 23435
rect 7552 23403 7584 23435
rect 7624 23403 7656 23435
rect 7696 23403 7728 23435
rect 7768 23403 7800 23435
rect 7840 23403 7872 23435
rect 7912 23403 7944 23435
rect 7984 23403 8016 23435
rect 8056 23403 8088 23435
rect 8128 23403 8160 23435
rect 8200 23403 8232 23435
rect 8272 23403 8304 23435
rect 8344 23403 8376 23435
rect 8416 23403 8448 23435
rect 8488 23403 8520 23435
rect 8560 23403 8592 23435
rect 8632 23403 8664 23435
rect 8704 23403 8736 23435
rect 8776 23403 8808 23435
rect 8848 23403 8880 23435
rect 8920 23403 8952 23435
rect 8992 23403 9024 23435
rect 9064 23403 9096 23435
rect 9136 23403 9168 23435
rect 9208 23403 9240 23435
rect 9280 23403 9312 23435
rect 9352 23403 9384 23435
rect 9424 23403 9456 23435
rect 9496 23403 9528 23435
rect 9568 23403 9600 23435
rect 9640 23403 9672 23435
rect 9712 23403 9744 23435
rect 9784 23403 9816 23435
rect 9856 23403 9888 23435
rect 9928 23403 9960 23435
rect 10000 23403 10032 23435
rect 10072 23403 10104 23435
rect 10144 23403 10176 23435
rect 10216 23403 10248 23435
rect 10288 23403 10320 23435
rect 10360 23403 10392 23435
rect 10432 23403 10464 23435
rect 10504 23403 10536 23435
rect 10576 23403 10608 23435
rect 10648 23403 10680 23435
rect 10720 23403 10752 23435
rect 10792 23403 10824 23435
rect 10864 23403 10896 23435
rect 10936 23403 10968 23435
rect 11008 23403 11040 23435
rect 11080 23403 11112 23435
rect 11152 23403 11184 23435
rect 11224 23403 11256 23435
rect 11296 23403 11328 23435
rect 11368 23403 11400 23435
rect 11440 23403 11472 23435
rect 11512 23403 11544 23435
rect 11584 23403 11616 23435
rect 11656 23403 11688 23435
rect 11728 23403 11760 23435
rect 11800 23403 11832 23435
rect 11872 23403 11904 23435
rect 11944 23403 11976 23435
rect 12016 23403 12048 23435
rect 12088 23403 12120 23435
rect 12160 23403 12192 23435
rect 12232 23403 12264 23435
rect 12304 23403 12336 23435
rect 12376 23403 12408 23435
rect 12448 23403 12480 23435
rect 12520 23403 12552 23435
rect 12592 23403 12624 23435
rect 12664 23403 12696 23435
rect 12736 23403 12768 23435
rect 12808 23403 12840 23435
rect 12880 23403 12912 23435
rect 12952 23403 12984 23435
rect 13024 23403 13056 23435
rect 13096 23403 13128 23435
rect 13168 23403 13200 23435
rect 13240 23403 13272 23435
rect 13312 23403 13344 23435
rect 13384 23403 13416 23435
rect 13456 23403 13488 23435
rect 13528 23403 13560 23435
rect 13600 23403 13632 23435
rect 13672 23403 13704 23435
rect 13744 23403 13776 23435
rect 13816 23403 13848 23435
rect 13888 23403 13920 23435
rect 13960 23403 13992 23435
rect 14032 23403 14064 23435
rect 14104 23403 14136 23435
rect 14176 23403 14208 23435
rect 14248 23403 14280 23435
rect 14320 23403 14352 23435
rect 14392 23403 14424 23435
rect 14464 23403 14496 23435
rect 14536 23403 14568 23435
rect 14608 23403 14640 23435
rect 14680 23403 14712 23435
rect 14752 23403 14784 23435
rect 14824 23403 14856 23435
rect 14896 23403 14928 23435
rect 14968 23403 15000 23435
rect 15040 23403 15072 23435
rect 15112 23403 15144 23435
rect 15184 23403 15216 23435
rect 15256 23403 15288 23435
rect 15328 23403 15360 23435
rect 15400 23403 15432 23435
rect 15472 23403 15504 23435
rect 15544 23403 15576 23435
rect 15616 23403 15648 23435
rect 15688 23403 15720 23435
rect 15760 23403 15792 23435
rect 15832 23403 15864 23435
rect 15904 23403 15936 23435
rect 64 23331 96 23363
rect 136 23331 168 23363
rect 208 23331 240 23363
rect 280 23331 312 23363
rect 352 23331 384 23363
rect 424 23331 456 23363
rect 496 23331 528 23363
rect 568 23331 600 23363
rect 640 23331 672 23363
rect 712 23331 744 23363
rect 784 23331 816 23363
rect 856 23331 888 23363
rect 928 23331 960 23363
rect 1000 23331 1032 23363
rect 1072 23331 1104 23363
rect 1144 23331 1176 23363
rect 1216 23331 1248 23363
rect 1288 23331 1320 23363
rect 1360 23331 1392 23363
rect 1432 23331 1464 23363
rect 1504 23331 1536 23363
rect 1576 23331 1608 23363
rect 1648 23331 1680 23363
rect 1720 23331 1752 23363
rect 1792 23331 1824 23363
rect 1864 23331 1896 23363
rect 1936 23331 1968 23363
rect 2008 23331 2040 23363
rect 2080 23331 2112 23363
rect 2152 23331 2184 23363
rect 2224 23331 2256 23363
rect 2296 23331 2328 23363
rect 2368 23331 2400 23363
rect 2440 23331 2472 23363
rect 2512 23331 2544 23363
rect 2584 23331 2616 23363
rect 2656 23331 2688 23363
rect 2728 23331 2760 23363
rect 2800 23331 2832 23363
rect 2872 23331 2904 23363
rect 2944 23331 2976 23363
rect 3016 23331 3048 23363
rect 3088 23331 3120 23363
rect 3160 23331 3192 23363
rect 3232 23331 3264 23363
rect 3304 23331 3336 23363
rect 3376 23331 3408 23363
rect 3448 23331 3480 23363
rect 3520 23331 3552 23363
rect 3592 23331 3624 23363
rect 3664 23331 3696 23363
rect 3736 23331 3768 23363
rect 3808 23331 3840 23363
rect 3880 23331 3912 23363
rect 3952 23331 3984 23363
rect 4024 23331 4056 23363
rect 4096 23331 4128 23363
rect 4168 23331 4200 23363
rect 4240 23331 4272 23363
rect 4312 23331 4344 23363
rect 4384 23331 4416 23363
rect 4456 23331 4488 23363
rect 4528 23331 4560 23363
rect 4600 23331 4632 23363
rect 4672 23331 4704 23363
rect 4744 23331 4776 23363
rect 4816 23331 4848 23363
rect 4888 23331 4920 23363
rect 4960 23331 4992 23363
rect 5032 23331 5064 23363
rect 5104 23331 5136 23363
rect 5176 23331 5208 23363
rect 5248 23331 5280 23363
rect 5320 23331 5352 23363
rect 5392 23331 5424 23363
rect 5464 23331 5496 23363
rect 5536 23331 5568 23363
rect 5608 23331 5640 23363
rect 5680 23331 5712 23363
rect 5752 23331 5784 23363
rect 5824 23331 5856 23363
rect 5896 23331 5928 23363
rect 5968 23331 6000 23363
rect 6040 23331 6072 23363
rect 6112 23331 6144 23363
rect 6184 23331 6216 23363
rect 6256 23331 6288 23363
rect 6328 23331 6360 23363
rect 6400 23331 6432 23363
rect 6472 23331 6504 23363
rect 6544 23331 6576 23363
rect 6616 23331 6648 23363
rect 6688 23331 6720 23363
rect 6760 23331 6792 23363
rect 6832 23331 6864 23363
rect 6904 23331 6936 23363
rect 6976 23331 7008 23363
rect 7048 23331 7080 23363
rect 7120 23331 7152 23363
rect 7192 23331 7224 23363
rect 7264 23331 7296 23363
rect 7336 23331 7368 23363
rect 7408 23331 7440 23363
rect 7480 23331 7512 23363
rect 7552 23331 7584 23363
rect 7624 23331 7656 23363
rect 7696 23331 7728 23363
rect 7768 23331 7800 23363
rect 7840 23331 7872 23363
rect 7912 23331 7944 23363
rect 7984 23331 8016 23363
rect 8056 23331 8088 23363
rect 8128 23331 8160 23363
rect 8200 23331 8232 23363
rect 8272 23331 8304 23363
rect 8344 23331 8376 23363
rect 8416 23331 8448 23363
rect 8488 23331 8520 23363
rect 8560 23331 8592 23363
rect 8632 23331 8664 23363
rect 8704 23331 8736 23363
rect 8776 23331 8808 23363
rect 8848 23331 8880 23363
rect 8920 23331 8952 23363
rect 8992 23331 9024 23363
rect 9064 23331 9096 23363
rect 9136 23331 9168 23363
rect 9208 23331 9240 23363
rect 9280 23331 9312 23363
rect 9352 23331 9384 23363
rect 9424 23331 9456 23363
rect 9496 23331 9528 23363
rect 9568 23331 9600 23363
rect 9640 23331 9672 23363
rect 9712 23331 9744 23363
rect 9784 23331 9816 23363
rect 9856 23331 9888 23363
rect 9928 23331 9960 23363
rect 10000 23331 10032 23363
rect 10072 23331 10104 23363
rect 10144 23331 10176 23363
rect 10216 23331 10248 23363
rect 10288 23331 10320 23363
rect 10360 23331 10392 23363
rect 10432 23331 10464 23363
rect 10504 23331 10536 23363
rect 10576 23331 10608 23363
rect 10648 23331 10680 23363
rect 10720 23331 10752 23363
rect 10792 23331 10824 23363
rect 10864 23331 10896 23363
rect 10936 23331 10968 23363
rect 11008 23331 11040 23363
rect 11080 23331 11112 23363
rect 11152 23331 11184 23363
rect 11224 23331 11256 23363
rect 11296 23331 11328 23363
rect 11368 23331 11400 23363
rect 11440 23331 11472 23363
rect 11512 23331 11544 23363
rect 11584 23331 11616 23363
rect 11656 23331 11688 23363
rect 11728 23331 11760 23363
rect 11800 23331 11832 23363
rect 11872 23331 11904 23363
rect 11944 23331 11976 23363
rect 12016 23331 12048 23363
rect 12088 23331 12120 23363
rect 12160 23331 12192 23363
rect 12232 23331 12264 23363
rect 12304 23331 12336 23363
rect 12376 23331 12408 23363
rect 12448 23331 12480 23363
rect 12520 23331 12552 23363
rect 12592 23331 12624 23363
rect 12664 23331 12696 23363
rect 12736 23331 12768 23363
rect 12808 23331 12840 23363
rect 12880 23331 12912 23363
rect 12952 23331 12984 23363
rect 13024 23331 13056 23363
rect 13096 23331 13128 23363
rect 13168 23331 13200 23363
rect 13240 23331 13272 23363
rect 13312 23331 13344 23363
rect 13384 23331 13416 23363
rect 13456 23331 13488 23363
rect 13528 23331 13560 23363
rect 13600 23331 13632 23363
rect 13672 23331 13704 23363
rect 13744 23331 13776 23363
rect 13816 23331 13848 23363
rect 13888 23331 13920 23363
rect 13960 23331 13992 23363
rect 14032 23331 14064 23363
rect 14104 23331 14136 23363
rect 14176 23331 14208 23363
rect 14248 23331 14280 23363
rect 14320 23331 14352 23363
rect 14392 23331 14424 23363
rect 14464 23331 14496 23363
rect 14536 23331 14568 23363
rect 14608 23331 14640 23363
rect 14680 23331 14712 23363
rect 14752 23331 14784 23363
rect 14824 23331 14856 23363
rect 14896 23331 14928 23363
rect 14968 23331 15000 23363
rect 15040 23331 15072 23363
rect 15112 23331 15144 23363
rect 15184 23331 15216 23363
rect 15256 23331 15288 23363
rect 15328 23331 15360 23363
rect 15400 23331 15432 23363
rect 15472 23331 15504 23363
rect 15544 23331 15576 23363
rect 15616 23331 15648 23363
rect 15688 23331 15720 23363
rect 15760 23331 15792 23363
rect 15832 23331 15864 23363
rect 15904 23331 15936 23363
rect 64 23259 96 23291
rect 136 23259 168 23291
rect 208 23259 240 23291
rect 280 23259 312 23291
rect 352 23259 384 23291
rect 424 23259 456 23291
rect 496 23259 528 23291
rect 568 23259 600 23291
rect 640 23259 672 23291
rect 712 23259 744 23291
rect 784 23259 816 23291
rect 856 23259 888 23291
rect 928 23259 960 23291
rect 1000 23259 1032 23291
rect 1072 23259 1104 23291
rect 1144 23259 1176 23291
rect 1216 23259 1248 23291
rect 1288 23259 1320 23291
rect 1360 23259 1392 23291
rect 1432 23259 1464 23291
rect 1504 23259 1536 23291
rect 1576 23259 1608 23291
rect 1648 23259 1680 23291
rect 1720 23259 1752 23291
rect 1792 23259 1824 23291
rect 1864 23259 1896 23291
rect 1936 23259 1968 23291
rect 2008 23259 2040 23291
rect 2080 23259 2112 23291
rect 2152 23259 2184 23291
rect 2224 23259 2256 23291
rect 2296 23259 2328 23291
rect 2368 23259 2400 23291
rect 2440 23259 2472 23291
rect 2512 23259 2544 23291
rect 2584 23259 2616 23291
rect 2656 23259 2688 23291
rect 2728 23259 2760 23291
rect 2800 23259 2832 23291
rect 2872 23259 2904 23291
rect 2944 23259 2976 23291
rect 3016 23259 3048 23291
rect 3088 23259 3120 23291
rect 3160 23259 3192 23291
rect 3232 23259 3264 23291
rect 3304 23259 3336 23291
rect 3376 23259 3408 23291
rect 3448 23259 3480 23291
rect 3520 23259 3552 23291
rect 3592 23259 3624 23291
rect 3664 23259 3696 23291
rect 3736 23259 3768 23291
rect 3808 23259 3840 23291
rect 3880 23259 3912 23291
rect 3952 23259 3984 23291
rect 4024 23259 4056 23291
rect 4096 23259 4128 23291
rect 4168 23259 4200 23291
rect 4240 23259 4272 23291
rect 4312 23259 4344 23291
rect 4384 23259 4416 23291
rect 4456 23259 4488 23291
rect 4528 23259 4560 23291
rect 4600 23259 4632 23291
rect 4672 23259 4704 23291
rect 4744 23259 4776 23291
rect 4816 23259 4848 23291
rect 4888 23259 4920 23291
rect 4960 23259 4992 23291
rect 5032 23259 5064 23291
rect 5104 23259 5136 23291
rect 5176 23259 5208 23291
rect 5248 23259 5280 23291
rect 5320 23259 5352 23291
rect 5392 23259 5424 23291
rect 5464 23259 5496 23291
rect 5536 23259 5568 23291
rect 5608 23259 5640 23291
rect 5680 23259 5712 23291
rect 5752 23259 5784 23291
rect 5824 23259 5856 23291
rect 5896 23259 5928 23291
rect 5968 23259 6000 23291
rect 6040 23259 6072 23291
rect 6112 23259 6144 23291
rect 6184 23259 6216 23291
rect 6256 23259 6288 23291
rect 6328 23259 6360 23291
rect 6400 23259 6432 23291
rect 6472 23259 6504 23291
rect 6544 23259 6576 23291
rect 6616 23259 6648 23291
rect 6688 23259 6720 23291
rect 6760 23259 6792 23291
rect 6832 23259 6864 23291
rect 6904 23259 6936 23291
rect 6976 23259 7008 23291
rect 7048 23259 7080 23291
rect 7120 23259 7152 23291
rect 7192 23259 7224 23291
rect 7264 23259 7296 23291
rect 7336 23259 7368 23291
rect 7408 23259 7440 23291
rect 7480 23259 7512 23291
rect 7552 23259 7584 23291
rect 7624 23259 7656 23291
rect 7696 23259 7728 23291
rect 7768 23259 7800 23291
rect 7840 23259 7872 23291
rect 7912 23259 7944 23291
rect 7984 23259 8016 23291
rect 8056 23259 8088 23291
rect 8128 23259 8160 23291
rect 8200 23259 8232 23291
rect 8272 23259 8304 23291
rect 8344 23259 8376 23291
rect 8416 23259 8448 23291
rect 8488 23259 8520 23291
rect 8560 23259 8592 23291
rect 8632 23259 8664 23291
rect 8704 23259 8736 23291
rect 8776 23259 8808 23291
rect 8848 23259 8880 23291
rect 8920 23259 8952 23291
rect 8992 23259 9024 23291
rect 9064 23259 9096 23291
rect 9136 23259 9168 23291
rect 9208 23259 9240 23291
rect 9280 23259 9312 23291
rect 9352 23259 9384 23291
rect 9424 23259 9456 23291
rect 9496 23259 9528 23291
rect 9568 23259 9600 23291
rect 9640 23259 9672 23291
rect 9712 23259 9744 23291
rect 9784 23259 9816 23291
rect 9856 23259 9888 23291
rect 9928 23259 9960 23291
rect 10000 23259 10032 23291
rect 10072 23259 10104 23291
rect 10144 23259 10176 23291
rect 10216 23259 10248 23291
rect 10288 23259 10320 23291
rect 10360 23259 10392 23291
rect 10432 23259 10464 23291
rect 10504 23259 10536 23291
rect 10576 23259 10608 23291
rect 10648 23259 10680 23291
rect 10720 23259 10752 23291
rect 10792 23259 10824 23291
rect 10864 23259 10896 23291
rect 10936 23259 10968 23291
rect 11008 23259 11040 23291
rect 11080 23259 11112 23291
rect 11152 23259 11184 23291
rect 11224 23259 11256 23291
rect 11296 23259 11328 23291
rect 11368 23259 11400 23291
rect 11440 23259 11472 23291
rect 11512 23259 11544 23291
rect 11584 23259 11616 23291
rect 11656 23259 11688 23291
rect 11728 23259 11760 23291
rect 11800 23259 11832 23291
rect 11872 23259 11904 23291
rect 11944 23259 11976 23291
rect 12016 23259 12048 23291
rect 12088 23259 12120 23291
rect 12160 23259 12192 23291
rect 12232 23259 12264 23291
rect 12304 23259 12336 23291
rect 12376 23259 12408 23291
rect 12448 23259 12480 23291
rect 12520 23259 12552 23291
rect 12592 23259 12624 23291
rect 12664 23259 12696 23291
rect 12736 23259 12768 23291
rect 12808 23259 12840 23291
rect 12880 23259 12912 23291
rect 12952 23259 12984 23291
rect 13024 23259 13056 23291
rect 13096 23259 13128 23291
rect 13168 23259 13200 23291
rect 13240 23259 13272 23291
rect 13312 23259 13344 23291
rect 13384 23259 13416 23291
rect 13456 23259 13488 23291
rect 13528 23259 13560 23291
rect 13600 23259 13632 23291
rect 13672 23259 13704 23291
rect 13744 23259 13776 23291
rect 13816 23259 13848 23291
rect 13888 23259 13920 23291
rect 13960 23259 13992 23291
rect 14032 23259 14064 23291
rect 14104 23259 14136 23291
rect 14176 23259 14208 23291
rect 14248 23259 14280 23291
rect 14320 23259 14352 23291
rect 14392 23259 14424 23291
rect 14464 23259 14496 23291
rect 14536 23259 14568 23291
rect 14608 23259 14640 23291
rect 14680 23259 14712 23291
rect 14752 23259 14784 23291
rect 14824 23259 14856 23291
rect 14896 23259 14928 23291
rect 14968 23259 15000 23291
rect 15040 23259 15072 23291
rect 15112 23259 15144 23291
rect 15184 23259 15216 23291
rect 15256 23259 15288 23291
rect 15328 23259 15360 23291
rect 15400 23259 15432 23291
rect 15472 23259 15504 23291
rect 15544 23259 15576 23291
rect 15616 23259 15648 23291
rect 15688 23259 15720 23291
rect 15760 23259 15792 23291
rect 15832 23259 15864 23291
rect 15904 23259 15936 23291
rect 64 23187 96 23219
rect 136 23187 168 23219
rect 208 23187 240 23219
rect 280 23187 312 23219
rect 352 23187 384 23219
rect 424 23187 456 23219
rect 496 23187 528 23219
rect 568 23187 600 23219
rect 640 23187 672 23219
rect 712 23187 744 23219
rect 784 23187 816 23219
rect 856 23187 888 23219
rect 928 23187 960 23219
rect 1000 23187 1032 23219
rect 1072 23187 1104 23219
rect 1144 23187 1176 23219
rect 1216 23187 1248 23219
rect 1288 23187 1320 23219
rect 1360 23187 1392 23219
rect 1432 23187 1464 23219
rect 1504 23187 1536 23219
rect 1576 23187 1608 23219
rect 1648 23187 1680 23219
rect 1720 23187 1752 23219
rect 1792 23187 1824 23219
rect 1864 23187 1896 23219
rect 1936 23187 1968 23219
rect 2008 23187 2040 23219
rect 2080 23187 2112 23219
rect 2152 23187 2184 23219
rect 2224 23187 2256 23219
rect 2296 23187 2328 23219
rect 2368 23187 2400 23219
rect 2440 23187 2472 23219
rect 2512 23187 2544 23219
rect 2584 23187 2616 23219
rect 2656 23187 2688 23219
rect 2728 23187 2760 23219
rect 2800 23187 2832 23219
rect 2872 23187 2904 23219
rect 2944 23187 2976 23219
rect 3016 23187 3048 23219
rect 3088 23187 3120 23219
rect 3160 23187 3192 23219
rect 3232 23187 3264 23219
rect 3304 23187 3336 23219
rect 3376 23187 3408 23219
rect 3448 23187 3480 23219
rect 3520 23187 3552 23219
rect 3592 23187 3624 23219
rect 3664 23187 3696 23219
rect 3736 23187 3768 23219
rect 3808 23187 3840 23219
rect 3880 23187 3912 23219
rect 3952 23187 3984 23219
rect 4024 23187 4056 23219
rect 4096 23187 4128 23219
rect 4168 23187 4200 23219
rect 4240 23187 4272 23219
rect 4312 23187 4344 23219
rect 4384 23187 4416 23219
rect 4456 23187 4488 23219
rect 4528 23187 4560 23219
rect 4600 23187 4632 23219
rect 4672 23187 4704 23219
rect 4744 23187 4776 23219
rect 4816 23187 4848 23219
rect 4888 23187 4920 23219
rect 4960 23187 4992 23219
rect 5032 23187 5064 23219
rect 5104 23187 5136 23219
rect 5176 23187 5208 23219
rect 5248 23187 5280 23219
rect 5320 23187 5352 23219
rect 5392 23187 5424 23219
rect 5464 23187 5496 23219
rect 5536 23187 5568 23219
rect 5608 23187 5640 23219
rect 5680 23187 5712 23219
rect 5752 23187 5784 23219
rect 5824 23187 5856 23219
rect 5896 23187 5928 23219
rect 5968 23187 6000 23219
rect 6040 23187 6072 23219
rect 6112 23187 6144 23219
rect 6184 23187 6216 23219
rect 6256 23187 6288 23219
rect 6328 23187 6360 23219
rect 6400 23187 6432 23219
rect 6472 23187 6504 23219
rect 6544 23187 6576 23219
rect 6616 23187 6648 23219
rect 6688 23187 6720 23219
rect 6760 23187 6792 23219
rect 6832 23187 6864 23219
rect 6904 23187 6936 23219
rect 6976 23187 7008 23219
rect 7048 23187 7080 23219
rect 7120 23187 7152 23219
rect 7192 23187 7224 23219
rect 7264 23187 7296 23219
rect 7336 23187 7368 23219
rect 7408 23187 7440 23219
rect 7480 23187 7512 23219
rect 7552 23187 7584 23219
rect 7624 23187 7656 23219
rect 7696 23187 7728 23219
rect 7768 23187 7800 23219
rect 7840 23187 7872 23219
rect 7912 23187 7944 23219
rect 7984 23187 8016 23219
rect 8056 23187 8088 23219
rect 8128 23187 8160 23219
rect 8200 23187 8232 23219
rect 8272 23187 8304 23219
rect 8344 23187 8376 23219
rect 8416 23187 8448 23219
rect 8488 23187 8520 23219
rect 8560 23187 8592 23219
rect 8632 23187 8664 23219
rect 8704 23187 8736 23219
rect 8776 23187 8808 23219
rect 8848 23187 8880 23219
rect 8920 23187 8952 23219
rect 8992 23187 9024 23219
rect 9064 23187 9096 23219
rect 9136 23187 9168 23219
rect 9208 23187 9240 23219
rect 9280 23187 9312 23219
rect 9352 23187 9384 23219
rect 9424 23187 9456 23219
rect 9496 23187 9528 23219
rect 9568 23187 9600 23219
rect 9640 23187 9672 23219
rect 9712 23187 9744 23219
rect 9784 23187 9816 23219
rect 9856 23187 9888 23219
rect 9928 23187 9960 23219
rect 10000 23187 10032 23219
rect 10072 23187 10104 23219
rect 10144 23187 10176 23219
rect 10216 23187 10248 23219
rect 10288 23187 10320 23219
rect 10360 23187 10392 23219
rect 10432 23187 10464 23219
rect 10504 23187 10536 23219
rect 10576 23187 10608 23219
rect 10648 23187 10680 23219
rect 10720 23187 10752 23219
rect 10792 23187 10824 23219
rect 10864 23187 10896 23219
rect 10936 23187 10968 23219
rect 11008 23187 11040 23219
rect 11080 23187 11112 23219
rect 11152 23187 11184 23219
rect 11224 23187 11256 23219
rect 11296 23187 11328 23219
rect 11368 23187 11400 23219
rect 11440 23187 11472 23219
rect 11512 23187 11544 23219
rect 11584 23187 11616 23219
rect 11656 23187 11688 23219
rect 11728 23187 11760 23219
rect 11800 23187 11832 23219
rect 11872 23187 11904 23219
rect 11944 23187 11976 23219
rect 12016 23187 12048 23219
rect 12088 23187 12120 23219
rect 12160 23187 12192 23219
rect 12232 23187 12264 23219
rect 12304 23187 12336 23219
rect 12376 23187 12408 23219
rect 12448 23187 12480 23219
rect 12520 23187 12552 23219
rect 12592 23187 12624 23219
rect 12664 23187 12696 23219
rect 12736 23187 12768 23219
rect 12808 23187 12840 23219
rect 12880 23187 12912 23219
rect 12952 23187 12984 23219
rect 13024 23187 13056 23219
rect 13096 23187 13128 23219
rect 13168 23187 13200 23219
rect 13240 23187 13272 23219
rect 13312 23187 13344 23219
rect 13384 23187 13416 23219
rect 13456 23187 13488 23219
rect 13528 23187 13560 23219
rect 13600 23187 13632 23219
rect 13672 23187 13704 23219
rect 13744 23187 13776 23219
rect 13816 23187 13848 23219
rect 13888 23187 13920 23219
rect 13960 23187 13992 23219
rect 14032 23187 14064 23219
rect 14104 23187 14136 23219
rect 14176 23187 14208 23219
rect 14248 23187 14280 23219
rect 14320 23187 14352 23219
rect 14392 23187 14424 23219
rect 14464 23187 14496 23219
rect 14536 23187 14568 23219
rect 14608 23187 14640 23219
rect 14680 23187 14712 23219
rect 14752 23187 14784 23219
rect 14824 23187 14856 23219
rect 14896 23187 14928 23219
rect 14968 23187 15000 23219
rect 15040 23187 15072 23219
rect 15112 23187 15144 23219
rect 15184 23187 15216 23219
rect 15256 23187 15288 23219
rect 15328 23187 15360 23219
rect 15400 23187 15432 23219
rect 15472 23187 15504 23219
rect 15544 23187 15576 23219
rect 15616 23187 15648 23219
rect 15688 23187 15720 23219
rect 15760 23187 15792 23219
rect 15832 23187 15864 23219
rect 15904 23187 15936 23219
rect 18 23021 50 23053
rect 18 22952 50 22984
rect 18 22883 50 22915
rect 18 22814 50 22846
rect 18 22745 50 22777
rect 18 22676 50 22708
rect 18 22607 50 22639
rect 18 22538 50 22570
rect 18 22469 50 22501
rect 18 22400 50 22432
rect 18 22331 50 22363
rect 18 22262 50 22294
rect 18 22193 50 22225
rect 18 22124 50 22156
rect 18 22055 50 22087
rect 18 21986 50 22018
rect 18 21917 50 21949
rect 18 21848 50 21880
rect 18 21779 50 21811
rect 18 21710 50 21742
rect 18 21641 50 21673
rect 18 21572 50 21604
rect 18 21503 50 21535
rect 18 21434 50 21466
rect 18 21365 50 21397
rect 18 21296 50 21328
rect 18 21227 50 21259
rect 18 21158 50 21190
rect 18 21089 50 21121
rect 18 21020 50 21052
rect 18 20951 50 20983
rect 18 20882 50 20914
rect 18 20813 50 20845
rect 18 20744 50 20776
rect 18 20675 50 20707
rect 18 20606 50 20638
rect 18 20537 50 20569
rect 18 20468 50 20500
rect 18 20399 50 20431
rect 18 20330 50 20362
rect 18 20261 50 20293
rect 18 20192 50 20224
rect 18 20123 50 20155
rect 18 20054 50 20086
rect 18 19985 50 20017
rect 18 19916 50 19948
rect 18 19847 50 19879
rect 18 19778 50 19810
rect 18 19709 50 19741
rect 18 19640 50 19672
rect 18 19571 50 19603
rect 18 19502 50 19534
rect 18 19433 50 19465
rect 18 19364 50 19396
rect 18 19295 50 19327
rect 18 19226 50 19258
rect 18 19157 50 19189
rect 18 19088 50 19120
rect 18 19019 50 19051
rect 18 18950 50 18982
rect 18 18881 50 18913
rect 18 18812 50 18844
rect 18 18743 50 18775
rect 18 18674 50 18706
rect 18 18605 50 18637
rect 18 18536 50 18568
rect 18 18467 50 18499
rect 18 18398 50 18430
rect 18 18329 50 18361
rect 18 18260 50 18292
rect 18 18191 50 18223
rect 18 18122 50 18154
rect 18 18053 50 18085
rect 18 17984 50 18016
rect 18 17915 50 17947
rect 18 17846 50 17878
rect 18 17777 50 17809
rect 18 17708 50 17740
rect 18 17639 50 17671
rect 18 17570 50 17602
rect 18 17502 50 17534
rect 15951 23010 15983 23042
rect 15951 22942 15983 22974
rect 15951 22874 15983 22906
rect 15951 22806 15983 22838
rect 15951 22738 15983 22770
rect 15951 22670 15983 22702
rect 15951 22602 15983 22634
rect 15951 22534 15983 22566
rect 15951 22466 15983 22498
rect 15951 22398 15983 22430
rect 15951 22330 15983 22362
rect 15951 22262 15983 22294
rect 15951 22194 15983 22226
rect 15951 22126 15983 22158
rect 15951 22058 15983 22090
rect 15951 21990 15983 22022
rect 15951 21922 15983 21954
rect 15951 21854 15983 21886
rect 15951 21786 15983 21818
rect 15951 21718 15983 21750
rect 15951 21650 15983 21682
rect 15951 21582 15983 21614
rect 15951 21514 15983 21546
rect 15951 21446 15983 21478
rect 15951 21378 15983 21410
rect 15951 21310 15983 21342
rect 15951 21242 15983 21274
rect 15951 21174 15983 21206
rect 15951 21106 15983 21138
rect 15951 21038 15983 21070
rect 15951 20970 15983 21002
rect 15951 20902 15983 20934
rect 15951 20834 15983 20866
rect 15951 20766 15983 20798
rect 15951 20698 15983 20730
rect 15951 20630 15983 20662
rect 15951 20562 15983 20594
rect 15951 20494 15983 20526
rect 15951 20426 15983 20458
rect 15951 20358 15983 20390
rect 15951 20290 15983 20322
rect 15951 20222 15983 20254
rect 15951 20154 15983 20186
rect 15951 20086 15983 20118
rect 15951 20018 15983 20050
rect 15951 19950 15983 19982
rect 15951 19882 15983 19914
rect 15951 19814 15983 19846
rect 15951 19746 15983 19778
rect 15951 19678 15983 19710
rect 15951 19610 15983 19642
rect 15951 19542 15983 19574
rect 15951 19474 15983 19506
rect 15951 19406 15983 19438
rect 15951 19338 15983 19370
rect 15951 19270 15983 19302
rect 15951 19202 15983 19234
rect 15951 19134 15983 19166
rect 15951 19066 15983 19098
rect 15951 18998 15983 19030
rect 15951 18930 15983 18962
rect 15951 18862 15983 18894
rect 15951 18794 15983 18826
rect 15951 18726 15983 18758
rect 15951 18658 15983 18690
rect 15951 18590 15983 18622
rect 15951 18522 15983 18554
rect 15951 18454 15983 18486
rect 15951 18386 15983 18418
rect 15951 18318 15983 18350
rect 15951 18250 15983 18282
rect 15951 18182 15983 18214
rect 15951 18114 15983 18146
rect 15951 18046 15983 18078
rect 15951 17978 15983 18010
rect 15951 17910 15983 17942
rect 15951 17842 15983 17874
rect 15951 17774 15983 17806
rect 15951 17706 15983 17738
rect 15951 17638 15983 17670
rect 15951 17570 15983 17602
rect 15951 17502 15983 17534
rect 0 31416 16000 31430
rect 0 31384 50 31416
rect 82 31384 118 31416
rect 150 31384 186 31416
rect 218 31384 254 31416
rect 286 31384 322 31416
rect 354 31384 390 31416
rect 422 31384 458 31416
rect 490 31384 526 31416
rect 558 31384 594 31416
rect 626 31384 662 31416
rect 694 31384 730 31416
rect 762 31384 798 31416
rect 830 31384 866 31416
rect 898 31384 934 31416
rect 966 31384 1002 31416
rect 1034 31384 1070 31416
rect 1102 31384 1138 31416
rect 1170 31384 1206 31416
rect 1238 31384 1274 31416
rect 1306 31384 1342 31416
rect 1374 31384 1410 31416
rect 1442 31384 1478 31416
rect 1510 31384 1546 31416
rect 1578 31384 1614 31416
rect 1646 31384 1682 31416
rect 1714 31384 1750 31416
rect 1782 31384 1818 31416
rect 1850 31384 1886 31416
rect 1918 31384 1954 31416
rect 1986 31384 2022 31416
rect 2054 31384 2090 31416
rect 2122 31384 2158 31416
rect 2190 31384 2226 31416
rect 2258 31384 2294 31416
rect 2326 31384 2362 31416
rect 2394 31384 2430 31416
rect 2462 31384 2498 31416
rect 2530 31384 2566 31416
rect 2598 31384 2634 31416
rect 2666 31384 2702 31416
rect 2734 31384 2770 31416
rect 2802 31384 2838 31416
rect 2870 31384 2906 31416
rect 2938 31384 2974 31416
rect 3006 31384 3042 31416
rect 3074 31384 3110 31416
rect 3142 31384 3178 31416
rect 3210 31384 3246 31416
rect 3278 31384 3314 31416
rect 3346 31384 3382 31416
rect 3414 31384 3450 31416
rect 3482 31384 3518 31416
rect 3550 31384 3586 31416
rect 3618 31384 3654 31416
rect 3686 31384 3722 31416
rect 3754 31384 3790 31416
rect 3822 31384 3858 31416
rect 3890 31384 3926 31416
rect 3958 31384 3994 31416
rect 4026 31384 4062 31416
rect 4094 31384 4130 31416
rect 4162 31384 4198 31416
rect 4230 31384 4266 31416
rect 4298 31384 4334 31416
rect 4366 31384 4402 31416
rect 4434 31384 4470 31416
rect 4502 31384 4538 31416
rect 4570 31384 4606 31416
rect 4638 31384 4674 31416
rect 4706 31384 4742 31416
rect 4774 31384 4810 31416
rect 4842 31384 4878 31416
rect 4910 31384 4946 31416
rect 4978 31384 5014 31416
rect 5046 31384 5082 31416
rect 5114 31384 5150 31416
rect 5182 31384 5218 31416
rect 5250 31384 5286 31416
rect 5318 31384 5354 31416
rect 5386 31384 5422 31416
rect 5454 31384 5490 31416
rect 5522 31384 5558 31416
rect 5590 31384 5626 31416
rect 5658 31384 5694 31416
rect 5726 31384 5762 31416
rect 5794 31384 5830 31416
rect 5862 31384 5898 31416
rect 5930 31384 5966 31416
rect 5998 31384 6034 31416
rect 6066 31384 6102 31416
rect 6134 31384 6170 31416
rect 6202 31384 6238 31416
rect 6270 31384 6306 31416
rect 6338 31384 6374 31416
rect 6406 31384 6442 31416
rect 6474 31384 6510 31416
rect 6542 31384 6578 31416
rect 6610 31384 6646 31416
rect 6678 31384 6714 31416
rect 6746 31384 6782 31416
rect 6814 31384 6850 31416
rect 6882 31384 6918 31416
rect 6950 31384 6986 31416
rect 7018 31384 7054 31416
rect 7086 31384 7122 31416
rect 7154 31384 7190 31416
rect 7222 31384 7258 31416
rect 7290 31384 7326 31416
rect 7358 31384 7394 31416
rect 7426 31384 7462 31416
rect 7494 31384 7530 31416
rect 7562 31384 7598 31416
rect 7630 31384 7666 31416
rect 7698 31384 7734 31416
rect 7766 31384 7802 31416
rect 7834 31384 7870 31416
rect 7902 31384 7938 31416
rect 7970 31384 8006 31416
rect 8038 31384 8074 31416
rect 8106 31384 8142 31416
rect 8174 31384 8210 31416
rect 8242 31384 8278 31416
rect 8310 31384 8346 31416
rect 8378 31384 8414 31416
rect 8446 31384 8482 31416
rect 8514 31384 8550 31416
rect 8582 31384 8618 31416
rect 8650 31384 8686 31416
rect 8718 31384 8754 31416
rect 8786 31384 8822 31416
rect 8854 31384 8890 31416
rect 8922 31384 8958 31416
rect 8990 31384 9026 31416
rect 9058 31384 9094 31416
rect 9126 31384 9162 31416
rect 9194 31384 9230 31416
rect 9262 31384 9298 31416
rect 9330 31384 9366 31416
rect 9398 31384 9434 31416
rect 9466 31384 9502 31416
rect 9534 31384 9570 31416
rect 9602 31384 9638 31416
rect 9670 31384 9706 31416
rect 9738 31384 9774 31416
rect 9806 31384 9842 31416
rect 9874 31384 9910 31416
rect 9942 31384 9978 31416
rect 10010 31384 10046 31416
rect 10078 31384 10114 31416
rect 10146 31384 10182 31416
rect 10214 31384 10250 31416
rect 10282 31384 10318 31416
rect 10350 31384 10386 31416
rect 10418 31384 10454 31416
rect 10486 31384 10522 31416
rect 10554 31384 10590 31416
rect 10622 31384 10658 31416
rect 10690 31384 10726 31416
rect 10758 31384 10794 31416
rect 10826 31384 10862 31416
rect 10894 31384 10930 31416
rect 10962 31384 10998 31416
rect 11030 31384 11066 31416
rect 11098 31384 11134 31416
rect 11166 31384 11202 31416
rect 11234 31384 11270 31416
rect 11302 31384 11338 31416
rect 11370 31384 11406 31416
rect 11438 31384 11474 31416
rect 11506 31384 11542 31416
rect 11574 31384 11610 31416
rect 11642 31384 11678 31416
rect 11710 31384 11746 31416
rect 11778 31384 11814 31416
rect 11846 31384 11882 31416
rect 11914 31384 11950 31416
rect 11982 31384 12018 31416
rect 12050 31384 12086 31416
rect 12118 31384 12154 31416
rect 12186 31384 12222 31416
rect 12254 31384 12290 31416
rect 12322 31384 12358 31416
rect 12390 31384 12426 31416
rect 12458 31384 12494 31416
rect 12526 31384 12562 31416
rect 12594 31384 12630 31416
rect 12662 31384 12698 31416
rect 12730 31384 12766 31416
rect 12798 31384 12834 31416
rect 12866 31384 12902 31416
rect 12934 31384 12970 31416
rect 13002 31384 13038 31416
rect 13070 31384 13106 31416
rect 13138 31384 13174 31416
rect 13206 31384 13242 31416
rect 13274 31384 13310 31416
rect 13342 31384 13378 31416
rect 13410 31384 13446 31416
rect 13478 31384 13514 31416
rect 13546 31384 13582 31416
rect 13614 31384 13650 31416
rect 13682 31384 13718 31416
rect 13750 31384 13786 31416
rect 13818 31384 13854 31416
rect 13886 31384 13922 31416
rect 13954 31384 13990 31416
rect 14022 31384 14058 31416
rect 14090 31384 14126 31416
rect 14158 31384 14194 31416
rect 14226 31384 14262 31416
rect 14294 31384 14330 31416
rect 14362 31384 14398 31416
rect 14430 31384 14466 31416
rect 14498 31384 14534 31416
rect 14566 31384 14602 31416
rect 14634 31384 14670 31416
rect 14702 31384 14738 31416
rect 14770 31384 14806 31416
rect 14838 31384 14874 31416
rect 14906 31384 14942 31416
rect 14974 31384 15010 31416
rect 15042 31384 15078 31416
rect 15110 31384 15146 31416
rect 15178 31384 15214 31416
rect 15246 31384 15282 31416
rect 15314 31384 15350 31416
rect 15382 31384 15442 31416
rect 15474 31384 15510 31416
rect 15542 31384 15578 31416
rect 15610 31384 15646 31416
rect 15678 31384 15714 31416
rect 15746 31384 15782 31416
rect 15814 31384 15850 31416
rect 15882 31384 15918 31416
rect 15950 31384 16000 31416
rect 0 31370 16000 31384
rect 0 27971 16000 28034
rect 0 27939 64 27971
rect 96 27939 136 27971
rect 168 27939 208 27971
rect 240 27939 280 27971
rect 312 27939 352 27971
rect 384 27939 424 27971
rect 456 27939 496 27971
rect 528 27939 568 27971
rect 600 27939 640 27971
rect 672 27939 712 27971
rect 744 27939 784 27971
rect 816 27939 856 27971
rect 888 27939 928 27971
rect 960 27939 1000 27971
rect 1032 27939 1072 27971
rect 1104 27939 1144 27971
rect 1176 27939 1216 27971
rect 1248 27939 1288 27971
rect 1320 27939 1360 27971
rect 1392 27939 1432 27971
rect 1464 27939 1504 27971
rect 1536 27939 1576 27971
rect 1608 27939 1648 27971
rect 1680 27939 1720 27971
rect 1752 27939 1792 27971
rect 1824 27939 1864 27971
rect 1896 27939 1936 27971
rect 1968 27939 2008 27971
rect 2040 27939 2080 27971
rect 2112 27939 2152 27971
rect 2184 27939 2224 27971
rect 2256 27939 2296 27971
rect 2328 27939 2368 27971
rect 2400 27939 2440 27971
rect 2472 27939 2512 27971
rect 2544 27939 2584 27971
rect 2616 27939 2656 27971
rect 2688 27939 2728 27971
rect 2760 27939 2800 27971
rect 2832 27939 2872 27971
rect 2904 27939 2944 27971
rect 2976 27939 3016 27971
rect 3048 27939 3088 27971
rect 3120 27939 3160 27971
rect 3192 27939 3232 27971
rect 3264 27939 3304 27971
rect 3336 27939 3376 27971
rect 3408 27939 3448 27971
rect 3480 27939 3520 27971
rect 3552 27939 3592 27971
rect 3624 27939 3664 27971
rect 3696 27939 3736 27971
rect 3768 27939 3808 27971
rect 3840 27939 3880 27971
rect 3912 27939 3952 27971
rect 3984 27939 4024 27971
rect 4056 27939 4096 27971
rect 4128 27939 4168 27971
rect 4200 27939 4240 27971
rect 4272 27939 4312 27971
rect 4344 27939 4384 27971
rect 4416 27939 4456 27971
rect 4488 27939 4528 27971
rect 4560 27939 4600 27971
rect 4632 27939 4672 27971
rect 4704 27939 4744 27971
rect 4776 27939 4816 27971
rect 4848 27939 4888 27971
rect 4920 27939 4960 27971
rect 4992 27939 5032 27971
rect 5064 27939 5104 27971
rect 5136 27939 5176 27971
rect 5208 27939 5248 27971
rect 5280 27939 5320 27971
rect 5352 27939 5392 27971
rect 5424 27939 5464 27971
rect 5496 27939 5536 27971
rect 5568 27939 5608 27971
rect 5640 27939 5680 27971
rect 5712 27939 5752 27971
rect 5784 27939 5824 27971
rect 5856 27939 5896 27971
rect 5928 27939 5968 27971
rect 6000 27939 6040 27971
rect 6072 27939 6112 27971
rect 6144 27939 6184 27971
rect 6216 27939 6256 27971
rect 6288 27939 6328 27971
rect 6360 27939 6400 27971
rect 6432 27939 6472 27971
rect 6504 27939 6544 27971
rect 6576 27939 6616 27971
rect 6648 27939 6688 27971
rect 6720 27939 6760 27971
rect 6792 27939 6832 27971
rect 6864 27939 6904 27971
rect 6936 27939 6976 27971
rect 7008 27939 7048 27971
rect 7080 27939 7120 27971
rect 7152 27939 7192 27971
rect 7224 27939 7264 27971
rect 7296 27939 7336 27971
rect 7368 27939 7408 27971
rect 7440 27939 7480 27971
rect 7512 27939 7552 27971
rect 7584 27939 7624 27971
rect 7656 27939 7696 27971
rect 7728 27939 7768 27971
rect 7800 27939 7840 27971
rect 7872 27939 7912 27971
rect 7944 27939 7984 27971
rect 8016 27939 8056 27971
rect 8088 27939 8128 27971
rect 8160 27939 8200 27971
rect 8232 27939 8272 27971
rect 8304 27939 8344 27971
rect 8376 27939 8416 27971
rect 8448 27939 8488 27971
rect 8520 27939 8560 27971
rect 8592 27939 8632 27971
rect 8664 27939 8704 27971
rect 8736 27939 8776 27971
rect 8808 27939 8848 27971
rect 8880 27939 8920 27971
rect 8952 27939 8992 27971
rect 9024 27939 9064 27971
rect 9096 27939 9136 27971
rect 9168 27939 9208 27971
rect 9240 27939 9280 27971
rect 9312 27939 9352 27971
rect 9384 27939 9424 27971
rect 9456 27939 9496 27971
rect 9528 27939 9568 27971
rect 9600 27939 9640 27971
rect 9672 27939 9712 27971
rect 9744 27939 9784 27971
rect 9816 27939 9856 27971
rect 9888 27939 9928 27971
rect 9960 27939 10000 27971
rect 10032 27939 10072 27971
rect 10104 27939 10144 27971
rect 10176 27939 10216 27971
rect 10248 27939 10288 27971
rect 10320 27939 10360 27971
rect 10392 27939 10432 27971
rect 10464 27939 10504 27971
rect 10536 27939 10576 27971
rect 10608 27939 10648 27971
rect 10680 27939 10720 27971
rect 10752 27939 10792 27971
rect 10824 27939 10864 27971
rect 10896 27939 10936 27971
rect 10968 27939 11008 27971
rect 11040 27939 11080 27971
rect 11112 27939 11152 27971
rect 11184 27939 11224 27971
rect 11256 27939 11296 27971
rect 11328 27939 11368 27971
rect 11400 27939 11440 27971
rect 11472 27939 11512 27971
rect 11544 27939 11584 27971
rect 11616 27939 11656 27971
rect 11688 27939 11728 27971
rect 11760 27939 11800 27971
rect 11832 27939 11872 27971
rect 11904 27939 11944 27971
rect 11976 27939 12016 27971
rect 12048 27939 12088 27971
rect 12120 27939 12160 27971
rect 12192 27939 12232 27971
rect 12264 27939 12304 27971
rect 12336 27939 12376 27971
rect 12408 27939 12448 27971
rect 12480 27939 12520 27971
rect 12552 27939 12592 27971
rect 12624 27939 12664 27971
rect 12696 27939 12736 27971
rect 12768 27939 12808 27971
rect 12840 27939 12880 27971
rect 12912 27939 12952 27971
rect 12984 27939 13024 27971
rect 13056 27939 13096 27971
rect 13128 27939 13168 27971
rect 13200 27939 13240 27971
rect 13272 27939 13312 27971
rect 13344 27939 13384 27971
rect 13416 27939 13456 27971
rect 13488 27939 13528 27971
rect 13560 27939 13600 27971
rect 13632 27939 13672 27971
rect 13704 27939 13744 27971
rect 13776 27939 13816 27971
rect 13848 27939 13888 27971
rect 13920 27939 13960 27971
rect 13992 27939 14032 27971
rect 14064 27939 14104 27971
rect 14136 27939 14176 27971
rect 14208 27939 14248 27971
rect 14280 27939 14320 27971
rect 14352 27939 14392 27971
rect 14424 27939 14464 27971
rect 14496 27939 14536 27971
rect 14568 27939 14608 27971
rect 14640 27939 14680 27971
rect 14712 27939 14752 27971
rect 14784 27939 14824 27971
rect 14856 27939 14896 27971
rect 14928 27939 14968 27971
rect 15000 27939 15040 27971
rect 15072 27939 15112 27971
rect 15144 27939 15184 27971
rect 15216 27939 15256 27971
rect 15288 27939 15328 27971
rect 15360 27939 15400 27971
rect 15432 27939 15472 27971
rect 15504 27939 15544 27971
rect 15576 27939 15616 27971
rect 15648 27939 15688 27971
rect 15720 27939 15760 27971
rect 15792 27939 15832 27971
rect 15864 27939 15904 27971
rect 15936 27939 16000 27971
rect 0 27899 16000 27939
rect 0 27867 64 27899
rect 96 27867 136 27899
rect 168 27867 208 27899
rect 240 27867 280 27899
rect 312 27867 352 27899
rect 384 27867 424 27899
rect 456 27867 496 27899
rect 528 27867 568 27899
rect 600 27867 640 27899
rect 672 27867 712 27899
rect 744 27867 784 27899
rect 816 27867 856 27899
rect 888 27867 928 27899
rect 960 27867 1000 27899
rect 1032 27867 1072 27899
rect 1104 27867 1144 27899
rect 1176 27867 1216 27899
rect 1248 27867 1288 27899
rect 1320 27867 1360 27899
rect 1392 27867 1432 27899
rect 1464 27867 1504 27899
rect 1536 27867 1576 27899
rect 1608 27867 1648 27899
rect 1680 27867 1720 27899
rect 1752 27867 1792 27899
rect 1824 27867 1864 27899
rect 1896 27867 1936 27899
rect 1968 27867 2008 27899
rect 2040 27867 2080 27899
rect 2112 27867 2152 27899
rect 2184 27867 2224 27899
rect 2256 27867 2296 27899
rect 2328 27867 2368 27899
rect 2400 27867 2440 27899
rect 2472 27867 2512 27899
rect 2544 27867 2584 27899
rect 2616 27867 2656 27899
rect 2688 27867 2728 27899
rect 2760 27867 2800 27899
rect 2832 27867 2872 27899
rect 2904 27867 2944 27899
rect 2976 27867 3016 27899
rect 3048 27867 3088 27899
rect 3120 27867 3160 27899
rect 3192 27867 3232 27899
rect 3264 27867 3304 27899
rect 3336 27867 3376 27899
rect 3408 27867 3448 27899
rect 3480 27867 3520 27899
rect 3552 27867 3592 27899
rect 3624 27867 3664 27899
rect 3696 27867 3736 27899
rect 3768 27867 3808 27899
rect 3840 27867 3880 27899
rect 3912 27867 3952 27899
rect 3984 27867 4024 27899
rect 4056 27867 4096 27899
rect 4128 27867 4168 27899
rect 4200 27867 4240 27899
rect 4272 27867 4312 27899
rect 4344 27867 4384 27899
rect 4416 27867 4456 27899
rect 4488 27867 4528 27899
rect 4560 27867 4600 27899
rect 4632 27867 4672 27899
rect 4704 27867 4744 27899
rect 4776 27867 4816 27899
rect 4848 27867 4888 27899
rect 4920 27867 4960 27899
rect 4992 27867 5032 27899
rect 5064 27867 5104 27899
rect 5136 27867 5176 27899
rect 5208 27867 5248 27899
rect 5280 27867 5320 27899
rect 5352 27867 5392 27899
rect 5424 27867 5464 27899
rect 5496 27867 5536 27899
rect 5568 27867 5608 27899
rect 5640 27867 5680 27899
rect 5712 27867 5752 27899
rect 5784 27867 5824 27899
rect 5856 27867 5896 27899
rect 5928 27867 5968 27899
rect 6000 27867 6040 27899
rect 6072 27867 6112 27899
rect 6144 27867 6184 27899
rect 6216 27867 6256 27899
rect 6288 27867 6328 27899
rect 6360 27867 6400 27899
rect 6432 27867 6472 27899
rect 6504 27867 6544 27899
rect 6576 27867 6616 27899
rect 6648 27867 6688 27899
rect 6720 27867 6760 27899
rect 6792 27867 6832 27899
rect 6864 27867 6904 27899
rect 6936 27867 6976 27899
rect 7008 27867 7048 27899
rect 7080 27867 7120 27899
rect 7152 27867 7192 27899
rect 7224 27867 7264 27899
rect 7296 27867 7336 27899
rect 7368 27867 7408 27899
rect 7440 27867 7480 27899
rect 7512 27867 7552 27899
rect 7584 27867 7624 27899
rect 7656 27867 7696 27899
rect 7728 27867 7768 27899
rect 7800 27867 7840 27899
rect 7872 27867 7912 27899
rect 7944 27867 7984 27899
rect 8016 27867 8056 27899
rect 8088 27867 8128 27899
rect 8160 27867 8200 27899
rect 8232 27867 8272 27899
rect 8304 27867 8344 27899
rect 8376 27867 8416 27899
rect 8448 27867 8488 27899
rect 8520 27867 8560 27899
rect 8592 27867 8632 27899
rect 8664 27867 8704 27899
rect 8736 27867 8776 27899
rect 8808 27867 8848 27899
rect 8880 27867 8920 27899
rect 8952 27867 8992 27899
rect 9024 27867 9064 27899
rect 9096 27867 9136 27899
rect 9168 27867 9208 27899
rect 9240 27867 9280 27899
rect 9312 27867 9352 27899
rect 9384 27867 9424 27899
rect 9456 27867 9496 27899
rect 9528 27867 9568 27899
rect 9600 27867 9640 27899
rect 9672 27867 9712 27899
rect 9744 27867 9784 27899
rect 9816 27867 9856 27899
rect 9888 27867 9928 27899
rect 9960 27867 10000 27899
rect 10032 27867 10072 27899
rect 10104 27867 10144 27899
rect 10176 27867 10216 27899
rect 10248 27867 10288 27899
rect 10320 27867 10360 27899
rect 10392 27867 10432 27899
rect 10464 27867 10504 27899
rect 10536 27867 10576 27899
rect 10608 27867 10648 27899
rect 10680 27867 10720 27899
rect 10752 27867 10792 27899
rect 10824 27867 10864 27899
rect 10896 27867 10936 27899
rect 10968 27867 11008 27899
rect 11040 27867 11080 27899
rect 11112 27867 11152 27899
rect 11184 27867 11224 27899
rect 11256 27867 11296 27899
rect 11328 27867 11368 27899
rect 11400 27867 11440 27899
rect 11472 27867 11512 27899
rect 11544 27867 11584 27899
rect 11616 27867 11656 27899
rect 11688 27867 11728 27899
rect 11760 27867 11800 27899
rect 11832 27867 11872 27899
rect 11904 27867 11944 27899
rect 11976 27867 12016 27899
rect 12048 27867 12088 27899
rect 12120 27867 12160 27899
rect 12192 27867 12232 27899
rect 12264 27867 12304 27899
rect 12336 27867 12376 27899
rect 12408 27867 12448 27899
rect 12480 27867 12520 27899
rect 12552 27867 12592 27899
rect 12624 27867 12664 27899
rect 12696 27867 12736 27899
rect 12768 27867 12808 27899
rect 12840 27867 12880 27899
rect 12912 27867 12952 27899
rect 12984 27867 13024 27899
rect 13056 27867 13096 27899
rect 13128 27867 13168 27899
rect 13200 27867 13240 27899
rect 13272 27867 13312 27899
rect 13344 27867 13384 27899
rect 13416 27867 13456 27899
rect 13488 27867 13528 27899
rect 13560 27867 13600 27899
rect 13632 27867 13672 27899
rect 13704 27867 13744 27899
rect 13776 27867 13816 27899
rect 13848 27867 13888 27899
rect 13920 27867 13960 27899
rect 13992 27867 14032 27899
rect 14064 27867 14104 27899
rect 14136 27867 14176 27899
rect 14208 27867 14248 27899
rect 14280 27867 14320 27899
rect 14352 27867 14392 27899
rect 14424 27867 14464 27899
rect 14496 27867 14536 27899
rect 14568 27867 14608 27899
rect 14640 27867 14680 27899
rect 14712 27867 14752 27899
rect 14784 27867 14824 27899
rect 14856 27867 14896 27899
rect 14928 27867 14968 27899
rect 15000 27867 15040 27899
rect 15072 27867 15112 27899
rect 15144 27867 15184 27899
rect 15216 27867 15256 27899
rect 15288 27867 15328 27899
rect 15360 27867 15400 27899
rect 15432 27867 15472 27899
rect 15504 27867 15544 27899
rect 15576 27867 15616 27899
rect 15648 27867 15688 27899
rect 15720 27867 15760 27899
rect 15792 27867 15832 27899
rect 15864 27867 15904 27899
rect 15936 27867 16000 27899
rect 0 27827 16000 27867
rect 0 27795 64 27827
rect 96 27795 136 27827
rect 168 27795 208 27827
rect 240 27795 280 27827
rect 312 27795 352 27827
rect 384 27795 424 27827
rect 456 27795 496 27827
rect 528 27795 568 27827
rect 600 27795 640 27827
rect 672 27795 712 27827
rect 744 27795 784 27827
rect 816 27795 856 27827
rect 888 27795 928 27827
rect 960 27795 1000 27827
rect 1032 27795 1072 27827
rect 1104 27795 1144 27827
rect 1176 27795 1216 27827
rect 1248 27795 1288 27827
rect 1320 27795 1360 27827
rect 1392 27795 1432 27827
rect 1464 27795 1504 27827
rect 1536 27795 1576 27827
rect 1608 27795 1648 27827
rect 1680 27795 1720 27827
rect 1752 27795 1792 27827
rect 1824 27795 1864 27827
rect 1896 27795 1936 27827
rect 1968 27795 2008 27827
rect 2040 27795 2080 27827
rect 2112 27795 2152 27827
rect 2184 27795 2224 27827
rect 2256 27795 2296 27827
rect 2328 27795 2368 27827
rect 2400 27795 2440 27827
rect 2472 27795 2512 27827
rect 2544 27795 2584 27827
rect 2616 27795 2656 27827
rect 2688 27795 2728 27827
rect 2760 27795 2800 27827
rect 2832 27795 2872 27827
rect 2904 27795 2944 27827
rect 2976 27795 3016 27827
rect 3048 27795 3088 27827
rect 3120 27795 3160 27827
rect 3192 27795 3232 27827
rect 3264 27795 3304 27827
rect 3336 27795 3376 27827
rect 3408 27795 3448 27827
rect 3480 27795 3520 27827
rect 3552 27795 3592 27827
rect 3624 27795 3664 27827
rect 3696 27795 3736 27827
rect 3768 27795 3808 27827
rect 3840 27795 3880 27827
rect 3912 27795 3952 27827
rect 3984 27795 4024 27827
rect 4056 27795 4096 27827
rect 4128 27795 4168 27827
rect 4200 27795 4240 27827
rect 4272 27795 4312 27827
rect 4344 27795 4384 27827
rect 4416 27795 4456 27827
rect 4488 27795 4528 27827
rect 4560 27795 4600 27827
rect 4632 27795 4672 27827
rect 4704 27795 4744 27827
rect 4776 27795 4816 27827
rect 4848 27795 4888 27827
rect 4920 27795 4960 27827
rect 4992 27795 5032 27827
rect 5064 27795 5104 27827
rect 5136 27795 5176 27827
rect 5208 27795 5248 27827
rect 5280 27795 5320 27827
rect 5352 27795 5392 27827
rect 5424 27795 5464 27827
rect 5496 27795 5536 27827
rect 5568 27795 5608 27827
rect 5640 27795 5680 27827
rect 5712 27795 5752 27827
rect 5784 27795 5824 27827
rect 5856 27795 5896 27827
rect 5928 27795 5968 27827
rect 6000 27795 6040 27827
rect 6072 27795 6112 27827
rect 6144 27795 6184 27827
rect 6216 27795 6256 27827
rect 6288 27795 6328 27827
rect 6360 27795 6400 27827
rect 6432 27795 6472 27827
rect 6504 27795 6544 27827
rect 6576 27795 6616 27827
rect 6648 27795 6688 27827
rect 6720 27795 6760 27827
rect 6792 27795 6832 27827
rect 6864 27795 6904 27827
rect 6936 27795 6976 27827
rect 7008 27795 7048 27827
rect 7080 27795 7120 27827
rect 7152 27795 7192 27827
rect 7224 27795 7264 27827
rect 7296 27795 7336 27827
rect 7368 27795 7408 27827
rect 7440 27795 7480 27827
rect 7512 27795 7552 27827
rect 7584 27795 7624 27827
rect 7656 27795 7696 27827
rect 7728 27795 7768 27827
rect 7800 27795 7840 27827
rect 7872 27795 7912 27827
rect 7944 27795 7984 27827
rect 8016 27795 8056 27827
rect 8088 27795 8128 27827
rect 8160 27795 8200 27827
rect 8232 27795 8272 27827
rect 8304 27795 8344 27827
rect 8376 27795 8416 27827
rect 8448 27795 8488 27827
rect 8520 27795 8560 27827
rect 8592 27795 8632 27827
rect 8664 27795 8704 27827
rect 8736 27795 8776 27827
rect 8808 27795 8848 27827
rect 8880 27795 8920 27827
rect 8952 27795 8992 27827
rect 9024 27795 9064 27827
rect 9096 27795 9136 27827
rect 9168 27795 9208 27827
rect 9240 27795 9280 27827
rect 9312 27795 9352 27827
rect 9384 27795 9424 27827
rect 9456 27795 9496 27827
rect 9528 27795 9568 27827
rect 9600 27795 9640 27827
rect 9672 27795 9712 27827
rect 9744 27795 9784 27827
rect 9816 27795 9856 27827
rect 9888 27795 9928 27827
rect 9960 27795 10000 27827
rect 10032 27795 10072 27827
rect 10104 27795 10144 27827
rect 10176 27795 10216 27827
rect 10248 27795 10288 27827
rect 10320 27795 10360 27827
rect 10392 27795 10432 27827
rect 10464 27795 10504 27827
rect 10536 27795 10576 27827
rect 10608 27795 10648 27827
rect 10680 27795 10720 27827
rect 10752 27795 10792 27827
rect 10824 27795 10864 27827
rect 10896 27795 10936 27827
rect 10968 27795 11008 27827
rect 11040 27795 11080 27827
rect 11112 27795 11152 27827
rect 11184 27795 11224 27827
rect 11256 27795 11296 27827
rect 11328 27795 11368 27827
rect 11400 27795 11440 27827
rect 11472 27795 11512 27827
rect 11544 27795 11584 27827
rect 11616 27795 11656 27827
rect 11688 27795 11728 27827
rect 11760 27795 11800 27827
rect 11832 27795 11872 27827
rect 11904 27795 11944 27827
rect 11976 27795 12016 27827
rect 12048 27795 12088 27827
rect 12120 27795 12160 27827
rect 12192 27795 12232 27827
rect 12264 27795 12304 27827
rect 12336 27795 12376 27827
rect 12408 27795 12448 27827
rect 12480 27795 12520 27827
rect 12552 27795 12592 27827
rect 12624 27795 12664 27827
rect 12696 27795 12736 27827
rect 12768 27795 12808 27827
rect 12840 27795 12880 27827
rect 12912 27795 12952 27827
rect 12984 27795 13024 27827
rect 13056 27795 13096 27827
rect 13128 27795 13168 27827
rect 13200 27795 13240 27827
rect 13272 27795 13312 27827
rect 13344 27795 13384 27827
rect 13416 27795 13456 27827
rect 13488 27795 13528 27827
rect 13560 27795 13600 27827
rect 13632 27795 13672 27827
rect 13704 27795 13744 27827
rect 13776 27795 13816 27827
rect 13848 27795 13888 27827
rect 13920 27795 13960 27827
rect 13992 27795 14032 27827
rect 14064 27795 14104 27827
rect 14136 27795 14176 27827
rect 14208 27795 14248 27827
rect 14280 27795 14320 27827
rect 14352 27795 14392 27827
rect 14424 27795 14464 27827
rect 14496 27795 14536 27827
rect 14568 27795 14608 27827
rect 14640 27795 14680 27827
rect 14712 27795 14752 27827
rect 14784 27795 14824 27827
rect 14856 27795 14896 27827
rect 14928 27795 14968 27827
rect 15000 27795 15040 27827
rect 15072 27795 15112 27827
rect 15144 27795 15184 27827
rect 15216 27795 15256 27827
rect 15288 27795 15328 27827
rect 15360 27795 15400 27827
rect 15432 27795 15472 27827
rect 15504 27795 15544 27827
rect 15576 27795 15616 27827
rect 15648 27795 15688 27827
rect 15720 27795 15760 27827
rect 15792 27795 15832 27827
rect 15864 27795 15904 27827
rect 15936 27795 16000 27827
rect 0 27755 16000 27795
rect 0 27723 64 27755
rect 96 27723 136 27755
rect 168 27723 208 27755
rect 240 27723 280 27755
rect 312 27723 352 27755
rect 384 27723 424 27755
rect 456 27723 496 27755
rect 528 27723 568 27755
rect 600 27723 640 27755
rect 672 27723 712 27755
rect 744 27723 784 27755
rect 816 27723 856 27755
rect 888 27723 928 27755
rect 960 27723 1000 27755
rect 1032 27723 1072 27755
rect 1104 27723 1144 27755
rect 1176 27723 1216 27755
rect 1248 27723 1288 27755
rect 1320 27723 1360 27755
rect 1392 27723 1432 27755
rect 1464 27723 1504 27755
rect 1536 27723 1576 27755
rect 1608 27723 1648 27755
rect 1680 27723 1720 27755
rect 1752 27723 1792 27755
rect 1824 27723 1864 27755
rect 1896 27723 1936 27755
rect 1968 27723 2008 27755
rect 2040 27723 2080 27755
rect 2112 27723 2152 27755
rect 2184 27723 2224 27755
rect 2256 27723 2296 27755
rect 2328 27723 2368 27755
rect 2400 27723 2440 27755
rect 2472 27723 2512 27755
rect 2544 27723 2584 27755
rect 2616 27723 2656 27755
rect 2688 27723 2728 27755
rect 2760 27723 2800 27755
rect 2832 27723 2872 27755
rect 2904 27723 2944 27755
rect 2976 27723 3016 27755
rect 3048 27723 3088 27755
rect 3120 27723 3160 27755
rect 3192 27723 3232 27755
rect 3264 27723 3304 27755
rect 3336 27723 3376 27755
rect 3408 27723 3448 27755
rect 3480 27723 3520 27755
rect 3552 27723 3592 27755
rect 3624 27723 3664 27755
rect 3696 27723 3736 27755
rect 3768 27723 3808 27755
rect 3840 27723 3880 27755
rect 3912 27723 3952 27755
rect 3984 27723 4024 27755
rect 4056 27723 4096 27755
rect 4128 27723 4168 27755
rect 4200 27723 4240 27755
rect 4272 27723 4312 27755
rect 4344 27723 4384 27755
rect 4416 27723 4456 27755
rect 4488 27723 4528 27755
rect 4560 27723 4600 27755
rect 4632 27723 4672 27755
rect 4704 27723 4744 27755
rect 4776 27723 4816 27755
rect 4848 27723 4888 27755
rect 4920 27723 4960 27755
rect 4992 27723 5032 27755
rect 5064 27723 5104 27755
rect 5136 27723 5176 27755
rect 5208 27723 5248 27755
rect 5280 27723 5320 27755
rect 5352 27723 5392 27755
rect 5424 27723 5464 27755
rect 5496 27723 5536 27755
rect 5568 27723 5608 27755
rect 5640 27723 5680 27755
rect 5712 27723 5752 27755
rect 5784 27723 5824 27755
rect 5856 27723 5896 27755
rect 5928 27723 5968 27755
rect 6000 27723 6040 27755
rect 6072 27723 6112 27755
rect 6144 27723 6184 27755
rect 6216 27723 6256 27755
rect 6288 27723 6328 27755
rect 6360 27723 6400 27755
rect 6432 27723 6472 27755
rect 6504 27723 6544 27755
rect 6576 27723 6616 27755
rect 6648 27723 6688 27755
rect 6720 27723 6760 27755
rect 6792 27723 6832 27755
rect 6864 27723 6904 27755
rect 6936 27723 6976 27755
rect 7008 27723 7048 27755
rect 7080 27723 7120 27755
rect 7152 27723 7192 27755
rect 7224 27723 7264 27755
rect 7296 27723 7336 27755
rect 7368 27723 7408 27755
rect 7440 27723 7480 27755
rect 7512 27723 7552 27755
rect 7584 27723 7624 27755
rect 7656 27723 7696 27755
rect 7728 27723 7768 27755
rect 7800 27723 7840 27755
rect 7872 27723 7912 27755
rect 7944 27723 7984 27755
rect 8016 27723 8056 27755
rect 8088 27723 8128 27755
rect 8160 27723 8200 27755
rect 8232 27723 8272 27755
rect 8304 27723 8344 27755
rect 8376 27723 8416 27755
rect 8448 27723 8488 27755
rect 8520 27723 8560 27755
rect 8592 27723 8632 27755
rect 8664 27723 8704 27755
rect 8736 27723 8776 27755
rect 8808 27723 8848 27755
rect 8880 27723 8920 27755
rect 8952 27723 8992 27755
rect 9024 27723 9064 27755
rect 9096 27723 9136 27755
rect 9168 27723 9208 27755
rect 9240 27723 9280 27755
rect 9312 27723 9352 27755
rect 9384 27723 9424 27755
rect 9456 27723 9496 27755
rect 9528 27723 9568 27755
rect 9600 27723 9640 27755
rect 9672 27723 9712 27755
rect 9744 27723 9784 27755
rect 9816 27723 9856 27755
rect 9888 27723 9928 27755
rect 9960 27723 10000 27755
rect 10032 27723 10072 27755
rect 10104 27723 10144 27755
rect 10176 27723 10216 27755
rect 10248 27723 10288 27755
rect 10320 27723 10360 27755
rect 10392 27723 10432 27755
rect 10464 27723 10504 27755
rect 10536 27723 10576 27755
rect 10608 27723 10648 27755
rect 10680 27723 10720 27755
rect 10752 27723 10792 27755
rect 10824 27723 10864 27755
rect 10896 27723 10936 27755
rect 10968 27723 11008 27755
rect 11040 27723 11080 27755
rect 11112 27723 11152 27755
rect 11184 27723 11224 27755
rect 11256 27723 11296 27755
rect 11328 27723 11368 27755
rect 11400 27723 11440 27755
rect 11472 27723 11512 27755
rect 11544 27723 11584 27755
rect 11616 27723 11656 27755
rect 11688 27723 11728 27755
rect 11760 27723 11800 27755
rect 11832 27723 11872 27755
rect 11904 27723 11944 27755
rect 11976 27723 12016 27755
rect 12048 27723 12088 27755
rect 12120 27723 12160 27755
rect 12192 27723 12232 27755
rect 12264 27723 12304 27755
rect 12336 27723 12376 27755
rect 12408 27723 12448 27755
rect 12480 27723 12520 27755
rect 12552 27723 12592 27755
rect 12624 27723 12664 27755
rect 12696 27723 12736 27755
rect 12768 27723 12808 27755
rect 12840 27723 12880 27755
rect 12912 27723 12952 27755
rect 12984 27723 13024 27755
rect 13056 27723 13096 27755
rect 13128 27723 13168 27755
rect 13200 27723 13240 27755
rect 13272 27723 13312 27755
rect 13344 27723 13384 27755
rect 13416 27723 13456 27755
rect 13488 27723 13528 27755
rect 13560 27723 13600 27755
rect 13632 27723 13672 27755
rect 13704 27723 13744 27755
rect 13776 27723 13816 27755
rect 13848 27723 13888 27755
rect 13920 27723 13960 27755
rect 13992 27723 14032 27755
rect 14064 27723 14104 27755
rect 14136 27723 14176 27755
rect 14208 27723 14248 27755
rect 14280 27723 14320 27755
rect 14352 27723 14392 27755
rect 14424 27723 14464 27755
rect 14496 27723 14536 27755
rect 14568 27723 14608 27755
rect 14640 27723 14680 27755
rect 14712 27723 14752 27755
rect 14784 27723 14824 27755
rect 14856 27723 14896 27755
rect 14928 27723 14968 27755
rect 15000 27723 15040 27755
rect 15072 27723 15112 27755
rect 15144 27723 15184 27755
rect 15216 27723 15256 27755
rect 15288 27723 15328 27755
rect 15360 27723 15400 27755
rect 15432 27723 15472 27755
rect 15504 27723 15544 27755
rect 15576 27723 15616 27755
rect 15648 27723 15688 27755
rect 15720 27723 15760 27755
rect 15792 27723 15832 27755
rect 15864 27723 15904 27755
rect 15936 27723 16000 27755
rect 0 27683 16000 27723
rect 0 27651 64 27683
rect 96 27651 136 27683
rect 168 27651 208 27683
rect 240 27651 280 27683
rect 312 27651 352 27683
rect 384 27651 424 27683
rect 456 27651 496 27683
rect 528 27651 568 27683
rect 600 27651 640 27683
rect 672 27651 712 27683
rect 744 27651 784 27683
rect 816 27651 856 27683
rect 888 27651 928 27683
rect 960 27651 1000 27683
rect 1032 27651 1072 27683
rect 1104 27651 1144 27683
rect 1176 27651 1216 27683
rect 1248 27651 1288 27683
rect 1320 27651 1360 27683
rect 1392 27651 1432 27683
rect 1464 27651 1504 27683
rect 1536 27651 1576 27683
rect 1608 27651 1648 27683
rect 1680 27651 1720 27683
rect 1752 27651 1792 27683
rect 1824 27651 1864 27683
rect 1896 27651 1936 27683
rect 1968 27651 2008 27683
rect 2040 27651 2080 27683
rect 2112 27651 2152 27683
rect 2184 27651 2224 27683
rect 2256 27651 2296 27683
rect 2328 27651 2368 27683
rect 2400 27651 2440 27683
rect 2472 27651 2512 27683
rect 2544 27651 2584 27683
rect 2616 27651 2656 27683
rect 2688 27651 2728 27683
rect 2760 27651 2800 27683
rect 2832 27651 2872 27683
rect 2904 27651 2944 27683
rect 2976 27651 3016 27683
rect 3048 27651 3088 27683
rect 3120 27651 3160 27683
rect 3192 27651 3232 27683
rect 3264 27651 3304 27683
rect 3336 27651 3376 27683
rect 3408 27651 3448 27683
rect 3480 27651 3520 27683
rect 3552 27651 3592 27683
rect 3624 27651 3664 27683
rect 3696 27651 3736 27683
rect 3768 27651 3808 27683
rect 3840 27651 3880 27683
rect 3912 27651 3952 27683
rect 3984 27651 4024 27683
rect 4056 27651 4096 27683
rect 4128 27651 4168 27683
rect 4200 27651 4240 27683
rect 4272 27651 4312 27683
rect 4344 27651 4384 27683
rect 4416 27651 4456 27683
rect 4488 27651 4528 27683
rect 4560 27651 4600 27683
rect 4632 27651 4672 27683
rect 4704 27651 4744 27683
rect 4776 27651 4816 27683
rect 4848 27651 4888 27683
rect 4920 27651 4960 27683
rect 4992 27651 5032 27683
rect 5064 27651 5104 27683
rect 5136 27651 5176 27683
rect 5208 27651 5248 27683
rect 5280 27651 5320 27683
rect 5352 27651 5392 27683
rect 5424 27651 5464 27683
rect 5496 27651 5536 27683
rect 5568 27651 5608 27683
rect 5640 27651 5680 27683
rect 5712 27651 5752 27683
rect 5784 27651 5824 27683
rect 5856 27651 5896 27683
rect 5928 27651 5968 27683
rect 6000 27651 6040 27683
rect 6072 27651 6112 27683
rect 6144 27651 6184 27683
rect 6216 27651 6256 27683
rect 6288 27651 6328 27683
rect 6360 27651 6400 27683
rect 6432 27651 6472 27683
rect 6504 27651 6544 27683
rect 6576 27651 6616 27683
rect 6648 27651 6688 27683
rect 6720 27651 6760 27683
rect 6792 27651 6832 27683
rect 6864 27651 6904 27683
rect 6936 27651 6976 27683
rect 7008 27651 7048 27683
rect 7080 27651 7120 27683
rect 7152 27651 7192 27683
rect 7224 27651 7264 27683
rect 7296 27651 7336 27683
rect 7368 27651 7408 27683
rect 7440 27651 7480 27683
rect 7512 27651 7552 27683
rect 7584 27651 7624 27683
rect 7656 27651 7696 27683
rect 7728 27651 7768 27683
rect 7800 27651 7840 27683
rect 7872 27651 7912 27683
rect 7944 27651 7984 27683
rect 8016 27651 8056 27683
rect 8088 27651 8128 27683
rect 8160 27651 8200 27683
rect 8232 27651 8272 27683
rect 8304 27651 8344 27683
rect 8376 27651 8416 27683
rect 8448 27651 8488 27683
rect 8520 27651 8560 27683
rect 8592 27651 8632 27683
rect 8664 27651 8704 27683
rect 8736 27651 8776 27683
rect 8808 27651 8848 27683
rect 8880 27651 8920 27683
rect 8952 27651 8992 27683
rect 9024 27651 9064 27683
rect 9096 27651 9136 27683
rect 9168 27651 9208 27683
rect 9240 27651 9280 27683
rect 9312 27651 9352 27683
rect 9384 27651 9424 27683
rect 9456 27651 9496 27683
rect 9528 27651 9568 27683
rect 9600 27651 9640 27683
rect 9672 27651 9712 27683
rect 9744 27651 9784 27683
rect 9816 27651 9856 27683
rect 9888 27651 9928 27683
rect 9960 27651 10000 27683
rect 10032 27651 10072 27683
rect 10104 27651 10144 27683
rect 10176 27651 10216 27683
rect 10248 27651 10288 27683
rect 10320 27651 10360 27683
rect 10392 27651 10432 27683
rect 10464 27651 10504 27683
rect 10536 27651 10576 27683
rect 10608 27651 10648 27683
rect 10680 27651 10720 27683
rect 10752 27651 10792 27683
rect 10824 27651 10864 27683
rect 10896 27651 10936 27683
rect 10968 27651 11008 27683
rect 11040 27651 11080 27683
rect 11112 27651 11152 27683
rect 11184 27651 11224 27683
rect 11256 27651 11296 27683
rect 11328 27651 11368 27683
rect 11400 27651 11440 27683
rect 11472 27651 11512 27683
rect 11544 27651 11584 27683
rect 11616 27651 11656 27683
rect 11688 27651 11728 27683
rect 11760 27651 11800 27683
rect 11832 27651 11872 27683
rect 11904 27651 11944 27683
rect 11976 27651 12016 27683
rect 12048 27651 12088 27683
rect 12120 27651 12160 27683
rect 12192 27651 12232 27683
rect 12264 27651 12304 27683
rect 12336 27651 12376 27683
rect 12408 27651 12448 27683
rect 12480 27651 12520 27683
rect 12552 27651 12592 27683
rect 12624 27651 12664 27683
rect 12696 27651 12736 27683
rect 12768 27651 12808 27683
rect 12840 27651 12880 27683
rect 12912 27651 12952 27683
rect 12984 27651 13024 27683
rect 13056 27651 13096 27683
rect 13128 27651 13168 27683
rect 13200 27651 13240 27683
rect 13272 27651 13312 27683
rect 13344 27651 13384 27683
rect 13416 27651 13456 27683
rect 13488 27651 13528 27683
rect 13560 27651 13600 27683
rect 13632 27651 13672 27683
rect 13704 27651 13744 27683
rect 13776 27651 13816 27683
rect 13848 27651 13888 27683
rect 13920 27651 13960 27683
rect 13992 27651 14032 27683
rect 14064 27651 14104 27683
rect 14136 27651 14176 27683
rect 14208 27651 14248 27683
rect 14280 27651 14320 27683
rect 14352 27651 14392 27683
rect 14424 27651 14464 27683
rect 14496 27651 14536 27683
rect 14568 27651 14608 27683
rect 14640 27651 14680 27683
rect 14712 27651 14752 27683
rect 14784 27651 14824 27683
rect 14856 27651 14896 27683
rect 14928 27651 14968 27683
rect 15000 27651 15040 27683
rect 15072 27651 15112 27683
rect 15144 27651 15184 27683
rect 15216 27651 15256 27683
rect 15288 27651 15328 27683
rect 15360 27651 15400 27683
rect 15432 27651 15472 27683
rect 15504 27651 15544 27683
rect 15576 27651 15616 27683
rect 15648 27651 15688 27683
rect 15720 27651 15760 27683
rect 15792 27651 15832 27683
rect 15864 27651 15904 27683
rect 15936 27651 16000 27683
rect 0 27611 16000 27651
rect 0 27579 64 27611
rect 96 27579 136 27611
rect 168 27579 208 27611
rect 240 27579 280 27611
rect 312 27579 352 27611
rect 384 27579 424 27611
rect 456 27579 496 27611
rect 528 27579 568 27611
rect 600 27579 640 27611
rect 672 27579 712 27611
rect 744 27579 784 27611
rect 816 27579 856 27611
rect 888 27579 928 27611
rect 960 27579 1000 27611
rect 1032 27579 1072 27611
rect 1104 27579 1144 27611
rect 1176 27579 1216 27611
rect 1248 27579 1288 27611
rect 1320 27579 1360 27611
rect 1392 27579 1432 27611
rect 1464 27579 1504 27611
rect 1536 27579 1576 27611
rect 1608 27579 1648 27611
rect 1680 27579 1720 27611
rect 1752 27579 1792 27611
rect 1824 27579 1864 27611
rect 1896 27579 1936 27611
rect 1968 27579 2008 27611
rect 2040 27579 2080 27611
rect 2112 27579 2152 27611
rect 2184 27579 2224 27611
rect 2256 27579 2296 27611
rect 2328 27579 2368 27611
rect 2400 27579 2440 27611
rect 2472 27579 2512 27611
rect 2544 27579 2584 27611
rect 2616 27579 2656 27611
rect 2688 27579 2728 27611
rect 2760 27579 2800 27611
rect 2832 27579 2872 27611
rect 2904 27579 2944 27611
rect 2976 27579 3016 27611
rect 3048 27579 3088 27611
rect 3120 27579 3160 27611
rect 3192 27579 3232 27611
rect 3264 27579 3304 27611
rect 3336 27579 3376 27611
rect 3408 27579 3448 27611
rect 3480 27579 3520 27611
rect 3552 27579 3592 27611
rect 3624 27579 3664 27611
rect 3696 27579 3736 27611
rect 3768 27579 3808 27611
rect 3840 27579 3880 27611
rect 3912 27579 3952 27611
rect 3984 27579 4024 27611
rect 4056 27579 4096 27611
rect 4128 27579 4168 27611
rect 4200 27579 4240 27611
rect 4272 27579 4312 27611
rect 4344 27579 4384 27611
rect 4416 27579 4456 27611
rect 4488 27579 4528 27611
rect 4560 27579 4600 27611
rect 4632 27579 4672 27611
rect 4704 27579 4744 27611
rect 4776 27579 4816 27611
rect 4848 27579 4888 27611
rect 4920 27579 4960 27611
rect 4992 27579 5032 27611
rect 5064 27579 5104 27611
rect 5136 27579 5176 27611
rect 5208 27579 5248 27611
rect 5280 27579 5320 27611
rect 5352 27579 5392 27611
rect 5424 27579 5464 27611
rect 5496 27579 5536 27611
rect 5568 27579 5608 27611
rect 5640 27579 5680 27611
rect 5712 27579 5752 27611
rect 5784 27579 5824 27611
rect 5856 27579 5896 27611
rect 5928 27579 5968 27611
rect 6000 27579 6040 27611
rect 6072 27579 6112 27611
rect 6144 27579 6184 27611
rect 6216 27579 6256 27611
rect 6288 27579 6328 27611
rect 6360 27579 6400 27611
rect 6432 27579 6472 27611
rect 6504 27579 6544 27611
rect 6576 27579 6616 27611
rect 6648 27579 6688 27611
rect 6720 27579 6760 27611
rect 6792 27579 6832 27611
rect 6864 27579 6904 27611
rect 6936 27579 6976 27611
rect 7008 27579 7048 27611
rect 7080 27579 7120 27611
rect 7152 27579 7192 27611
rect 7224 27579 7264 27611
rect 7296 27579 7336 27611
rect 7368 27579 7408 27611
rect 7440 27579 7480 27611
rect 7512 27579 7552 27611
rect 7584 27579 7624 27611
rect 7656 27579 7696 27611
rect 7728 27579 7768 27611
rect 7800 27579 7840 27611
rect 7872 27579 7912 27611
rect 7944 27579 7984 27611
rect 8016 27579 8056 27611
rect 8088 27579 8128 27611
rect 8160 27579 8200 27611
rect 8232 27579 8272 27611
rect 8304 27579 8344 27611
rect 8376 27579 8416 27611
rect 8448 27579 8488 27611
rect 8520 27579 8560 27611
rect 8592 27579 8632 27611
rect 8664 27579 8704 27611
rect 8736 27579 8776 27611
rect 8808 27579 8848 27611
rect 8880 27579 8920 27611
rect 8952 27579 8992 27611
rect 9024 27579 9064 27611
rect 9096 27579 9136 27611
rect 9168 27579 9208 27611
rect 9240 27579 9280 27611
rect 9312 27579 9352 27611
rect 9384 27579 9424 27611
rect 9456 27579 9496 27611
rect 9528 27579 9568 27611
rect 9600 27579 9640 27611
rect 9672 27579 9712 27611
rect 9744 27579 9784 27611
rect 9816 27579 9856 27611
rect 9888 27579 9928 27611
rect 9960 27579 10000 27611
rect 10032 27579 10072 27611
rect 10104 27579 10144 27611
rect 10176 27579 10216 27611
rect 10248 27579 10288 27611
rect 10320 27579 10360 27611
rect 10392 27579 10432 27611
rect 10464 27579 10504 27611
rect 10536 27579 10576 27611
rect 10608 27579 10648 27611
rect 10680 27579 10720 27611
rect 10752 27579 10792 27611
rect 10824 27579 10864 27611
rect 10896 27579 10936 27611
rect 10968 27579 11008 27611
rect 11040 27579 11080 27611
rect 11112 27579 11152 27611
rect 11184 27579 11224 27611
rect 11256 27579 11296 27611
rect 11328 27579 11368 27611
rect 11400 27579 11440 27611
rect 11472 27579 11512 27611
rect 11544 27579 11584 27611
rect 11616 27579 11656 27611
rect 11688 27579 11728 27611
rect 11760 27579 11800 27611
rect 11832 27579 11872 27611
rect 11904 27579 11944 27611
rect 11976 27579 12016 27611
rect 12048 27579 12088 27611
rect 12120 27579 12160 27611
rect 12192 27579 12232 27611
rect 12264 27579 12304 27611
rect 12336 27579 12376 27611
rect 12408 27579 12448 27611
rect 12480 27579 12520 27611
rect 12552 27579 12592 27611
rect 12624 27579 12664 27611
rect 12696 27579 12736 27611
rect 12768 27579 12808 27611
rect 12840 27579 12880 27611
rect 12912 27579 12952 27611
rect 12984 27579 13024 27611
rect 13056 27579 13096 27611
rect 13128 27579 13168 27611
rect 13200 27579 13240 27611
rect 13272 27579 13312 27611
rect 13344 27579 13384 27611
rect 13416 27579 13456 27611
rect 13488 27579 13528 27611
rect 13560 27579 13600 27611
rect 13632 27579 13672 27611
rect 13704 27579 13744 27611
rect 13776 27579 13816 27611
rect 13848 27579 13888 27611
rect 13920 27579 13960 27611
rect 13992 27579 14032 27611
rect 14064 27579 14104 27611
rect 14136 27579 14176 27611
rect 14208 27579 14248 27611
rect 14280 27579 14320 27611
rect 14352 27579 14392 27611
rect 14424 27579 14464 27611
rect 14496 27579 14536 27611
rect 14568 27579 14608 27611
rect 14640 27579 14680 27611
rect 14712 27579 14752 27611
rect 14784 27579 14824 27611
rect 14856 27579 14896 27611
rect 14928 27579 14968 27611
rect 15000 27579 15040 27611
rect 15072 27579 15112 27611
rect 15144 27579 15184 27611
rect 15216 27579 15256 27611
rect 15288 27579 15328 27611
rect 15360 27579 15400 27611
rect 15432 27579 15472 27611
rect 15504 27579 15544 27611
rect 15576 27579 15616 27611
rect 15648 27579 15688 27611
rect 15720 27579 15760 27611
rect 15792 27579 15832 27611
rect 15864 27579 15904 27611
rect 15936 27579 16000 27611
rect 0 27539 16000 27579
rect 0 27507 64 27539
rect 96 27507 136 27539
rect 168 27507 208 27539
rect 240 27507 280 27539
rect 312 27507 352 27539
rect 384 27507 424 27539
rect 456 27507 496 27539
rect 528 27507 568 27539
rect 600 27507 640 27539
rect 672 27507 712 27539
rect 744 27507 784 27539
rect 816 27507 856 27539
rect 888 27507 928 27539
rect 960 27507 1000 27539
rect 1032 27507 1072 27539
rect 1104 27507 1144 27539
rect 1176 27507 1216 27539
rect 1248 27507 1288 27539
rect 1320 27507 1360 27539
rect 1392 27507 1432 27539
rect 1464 27507 1504 27539
rect 1536 27507 1576 27539
rect 1608 27507 1648 27539
rect 1680 27507 1720 27539
rect 1752 27507 1792 27539
rect 1824 27507 1864 27539
rect 1896 27507 1936 27539
rect 1968 27507 2008 27539
rect 2040 27507 2080 27539
rect 2112 27507 2152 27539
rect 2184 27507 2224 27539
rect 2256 27507 2296 27539
rect 2328 27507 2368 27539
rect 2400 27507 2440 27539
rect 2472 27507 2512 27539
rect 2544 27507 2584 27539
rect 2616 27507 2656 27539
rect 2688 27507 2728 27539
rect 2760 27507 2800 27539
rect 2832 27507 2872 27539
rect 2904 27507 2944 27539
rect 2976 27507 3016 27539
rect 3048 27507 3088 27539
rect 3120 27507 3160 27539
rect 3192 27507 3232 27539
rect 3264 27507 3304 27539
rect 3336 27507 3376 27539
rect 3408 27507 3448 27539
rect 3480 27507 3520 27539
rect 3552 27507 3592 27539
rect 3624 27507 3664 27539
rect 3696 27507 3736 27539
rect 3768 27507 3808 27539
rect 3840 27507 3880 27539
rect 3912 27507 3952 27539
rect 3984 27507 4024 27539
rect 4056 27507 4096 27539
rect 4128 27507 4168 27539
rect 4200 27507 4240 27539
rect 4272 27507 4312 27539
rect 4344 27507 4384 27539
rect 4416 27507 4456 27539
rect 4488 27507 4528 27539
rect 4560 27507 4600 27539
rect 4632 27507 4672 27539
rect 4704 27507 4744 27539
rect 4776 27507 4816 27539
rect 4848 27507 4888 27539
rect 4920 27507 4960 27539
rect 4992 27507 5032 27539
rect 5064 27507 5104 27539
rect 5136 27507 5176 27539
rect 5208 27507 5248 27539
rect 5280 27507 5320 27539
rect 5352 27507 5392 27539
rect 5424 27507 5464 27539
rect 5496 27507 5536 27539
rect 5568 27507 5608 27539
rect 5640 27507 5680 27539
rect 5712 27507 5752 27539
rect 5784 27507 5824 27539
rect 5856 27507 5896 27539
rect 5928 27507 5968 27539
rect 6000 27507 6040 27539
rect 6072 27507 6112 27539
rect 6144 27507 6184 27539
rect 6216 27507 6256 27539
rect 6288 27507 6328 27539
rect 6360 27507 6400 27539
rect 6432 27507 6472 27539
rect 6504 27507 6544 27539
rect 6576 27507 6616 27539
rect 6648 27507 6688 27539
rect 6720 27507 6760 27539
rect 6792 27507 6832 27539
rect 6864 27507 6904 27539
rect 6936 27507 6976 27539
rect 7008 27507 7048 27539
rect 7080 27507 7120 27539
rect 7152 27507 7192 27539
rect 7224 27507 7264 27539
rect 7296 27507 7336 27539
rect 7368 27507 7408 27539
rect 7440 27507 7480 27539
rect 7512 27507 7552 27539
rect 7584 27507 7624 27539
rect 7656 27507 7696 27539
rect 7728 27507 7768 27539
rect 7800 27507 7840 27539
rect 7872 27507 7912 27539
rect 7944 27507 7984 27539
rect 8016 27507 8056 27539
rect 8088 27507 8128 27539
rect 8160 27507 8200 27539
rect 8232 27507 8272 27539
rect 8304 27507 8344 27539
rect 8376 27507 8416 27539
rect 8448 27507 8488 27539
rect 8520 27507 8560 27539
rect 8592 27507 8632 27539
rect 8664 27507 8704 27539
rect 8736 27507 8776 27539
rect 8808 27507 8848 27539
rect 8880 27507 8920 27539
rect 8952 27507 8992 27539
rect 9024 27507 9064 27539
rect 9096 27507 9136 27539
rect 9168 27507 9208 27539
rect 9240 27507 9280 27539
rect 9312 27507 9352 27539
rect 9384 27507 9424 27539
rect 9456 27507 9496 27539
rect 9528 27507 9568 27539
rect 9600 27507 9640 27539
rect 9672 27507 9712 27539
rect 9744 27507 9784 27539
rect 9816 27507 9856 27539
rect 9888 27507 9928 27539
rect 9960 27507 10000 27539
rect 10032 27507 10072 27539
rect 10104 27507 10144 27539
rect 10176 27507 10216 27539
rect 10248 27507 10288 27539
rect 10320 27507 10360 27539
rect 10392 27507 10432 27539
rect 10464 27507 10504 27539
rect 10536 27507 10576 27539
rect 10608 27507 10648 27539
rect 10680 27507 10720 27539
rect 10752 27507 10792 27539
rect 10824 27507 10864 27539
rect 10896 27507 10936 27539
rect 10968 27507 11008 27539
rect 11040 27507 11080 27539
rect 11112 27507 11152 27539
rect 11184 27507 11224 27539
rect 11256 27507 11296 27539
rect 11328 27507 11368 27539
rect 11400 27507 11440 27539
rect 11472 27507 11512 27539
rect 11544 27507 11584 27539
rect 11616 27507 11656 27539
rect 11688 27507 11728 27539
rect 11760 27507 11800 27539
rect 11832 27507 11872 27539
rect 11904 27507 11944 27539
rect 11976 27507 12016 27539
rect 12048 27507 12088 27539
rect 12120 27507 12160 27539
rect 12192 27507 12232 27539
rect 12264 27507 12304 27539
rect 12336 27507 12376 27539
rect 12408 27507 12448 27539
rect 12480 27507 12520 27539
rect 12552 27507 12592 27539
rect 12624 27507 12664 27539
rect 12696 27507 12736 27539
rect 12768 27507 12808 27539
rect 12840 27507 12880 27539
rect 12912 27507 12952 27539
rect 12984 27507 13024 27539
rect 13056 27507 13096 27539
rect 13128 27507 13168 27539
rect 13200 27507 13240 27539
rect 13272 27507 13312 27539
rect 13344 27507 13384 27539
rect 13416 27507 13456 27539
rect 13488 27507 13528 27539
rect 13560 27507 13600 27539
rect 13632 27507 13672 27539
rect 13704 27507 13744 27539
rect 13776 27507 13816 27539
rect 13848 27507 13888 27539
rect 13920 27507 13960 27539
rect 13992 27507 14032 27539
rect 14064 27507 14104 27539
rect 14136 27507 14176 27539
rect 14208 27507 14248 27539
rect 14280 27507 14320 27539
rect 14352 27507 14392 27539
rect 14424 27507 14464 27539
rect 14496 27507 14536 27539
rect 14568 27507 14608 27539
rect 14640 27507 14680 27539
rect 14712 27507 14752 27539
rect 14784 27507 14824 27539
rect 14856 27507 14896 27539
rect 14928 27507 14968 27539
rect 15000 27507 15040 27539
rect 15072 27507 15112 27539
rect 15144 27507 15184 27539
rect 15216 27507 15256 27539
rect 15288 27507 15328 27539
rect 15360 27507 15400 27539
rect 15432 27507 15472 27539
rect 15504 27507 15544 27539
rect 15576 27507 15616 27539
rect 15648 27507 15688 27539
rect 15720 27507 15760 27539
rect 15792 27507 15832 27539
rect 15864 27507 15904 27539
rect 15936 27507 16000 27539
rect 0 27467 16000 27507
rect 0 27435 64 27467
rect 96 27435 136 27467
rect 168 27435 208 27467
rect 240 27435 280 27467
rect 312 27435 352 27467
rect 384 27435 424 27467
rect 456 27435 496 27467
rect 528 27435 568 27467
rect 600 27435 640 27467
rect 672 27435 712 27467
rect 744 27435 784 27467
rect 816 27435 856 27467
rect 888 27435 928 27467
rect 960 27435 1000 27467
rect 1032 27435 1072 27467
rect 1104 27435 1144 27467
rect 1176 27435 1216 27467
rect 1248 27435 1288 27467
rect 1320 27435 1360 27467
rect 1392 27435 1432 27467
rect 1464 27435 1504 27467
rect 1536 27435 1576 27467
rect 1608 27435 1648 27467
rect 1680 27435 1720 27467
rect 1752 27435 1792 27467
rect 1824 27435 1864 27467
rect 1896 27435 1936 27467
rect 1968 27435 2008 27467
rect 2040 27435 2080 27467
rect 2112 27435 2152 27467
rect 2184 27435 2224 27467
rect 2256 27435 2296 27467
rect 2328 27435 2368 27467
rect 2400 27435 2440 27467
rect 2472 27435 2512 27467
rect 2544 27435 2584 27467
rect 2616 27435 2656 27467
rect 2688 27435 2728 27467
rect 2760 27435 2800 27467
rect 2832 27435 2872 27467
rect 2904 27435 2944 27467
rect 2976 27435 3016 27467
rect 3048 27435 3088 27467
rect 3120 27435 3160 27467
rect 3192 27435 3232 27467
rect 3264 27435 3304 27467
rect 3336 27435 3376 27467
rect 3408 27435 3448 27467
rect 3480 27435 3520 27467
rect 3552 27435 3592 27467
rect 3624 27435 3664 27467
rect 3696 27435 3736 27467
rect 3768 27435 3808 27467
rect 3840 27435 3880 27467
rect 3912 27435 3952 27467
rect 3984 27435 4024 27467
rect 4056 27435 4096 27467
rect 4128 27435 4168 27467
rect 4200 27435 4240 27467
rect 4272 27435 4312 27467
rect 4344 27435 4384 27467
rect 4416 27435 4456 27467
rect 4488 27435 4528 27467
rect 4560 27435 4600 27467
rect 4632 27435 4672 27467
rect 4704 27435 4744 27467
rect 4776 27435 4816 27467
rect 4848 27435 4888 27467
rect 4920 27435 4960 27467
rect 4992 27435 5032 27467
rect 5064 27435 5104 27467
rect 5136 27435 5176 27467
rect 5208 27435 5248 27467
rect 5280 27435 5320 27467
rect 5352 27435 5392 27467
rect 5424 27435 5464 27467
rect 5496 27435 5536 27467
rect 5568 27435 5608 27467
rect 5640 27435 5680 27467
rect 5712 27435 5752 27467
rect 5784 27435 5824 27467
rect 5856 27435 5896 27467
rect 5928 27435 5968 27467
rect 6000 27435 6040 27467
rect 6072 27435 6112 27467
rect 6144 27435 6184 27467
rect 6216 27435 6256 27467
rect 6288 27435 6328 27467
rect 6360 27435 6400 27467
rect 6432 27435 6472 27467
rect 6504 27435 6544 27467
rect 6576 27435 6616 27467
rect 6648 27435 6688 27467
rect 6720 27435 6760 27467
rect 6792 27435 6832 27467
rect 6864 27435 6904 27467
rect 6936 27435 6976 27467
rect 7008 27435 7048 27467
rect 7080 27435 7120 27467
rect 7152 27435 7192 27467
rect 7224 27435 7264 27467
rect 7296 27435 7336 27467
rect 7368 27435 7408 27467
rect 7440 27435 7480 27467
rect 7512 27435 7552 27467
rect 7584 27435 7624 27467
rect 7656 27435 7696 27467
rect 7728 27435 7768 27467
rect 7800 27435 7840 27467
rect 7872 27435 7912 27467
rect 7944 27435 7984 27467
rect 8016 27435 8056 27467
rect 8088 27435 8128 27467
rect 8160 27435 8200 27467
rect 8232 27435 8272 27467
rect 8304 27435 8344 27467
rect 8376 27435 8416 27467
rect 8448 27435 8488 27467
rect 8520 27435 8560 27467
rect 8592 27435 8632 27467
rect 8664 27435 8704 27467
rect 8736 27435 8776 27467
rect 8808 27435 8848 27467
rect 8880 27435 8920 27467
rect 8952 27435 8992 27467
rect 9024 27435 9064 27467
rect 9096 27435 9136 27467
rect 9168 27435 9208 27467
rect 9240 27435 9280 27467
rect 9312 27435 9352 27467
rect 9384 27435 9424 27467
rect 9456 27435 9496 27467
rect 9528 27435 9568 27467
rect 9600 27435 9640 27467
rect 9672 27435 9712 27467
rect 9744 27435 9784 27467
rect 9816 27435 9856 27467
rect 9888 27435 9928 27467
rect 9960 27435 10000 27467
rect 10032 27435 10072 27467
rect 10104 27435 10144 27467
rect 10176 27435 10216 27467
rect 10248 27435 10288 27467
rect 10320 27435 10360 27467
rect 10392 27435 10432 27467
rect 10464 27435 10504 27467
rect 10536 27435 10576 27467
rect 10608 27435 10648 27467
rect 10680 27435 10720 27467
rect 10752 27435 10792 27467
rect 10824 27435 10864 27467
rect 10896 27435 10936 27467
rect 10968 27435 11008 27467
rect 11040 27435 11080 27467
rect 11112 27435 11152 27467
rect 11184 27435 11224 27467
rect 11256 27435 11296 27467
rect 11328 27435 11368 27467
rect 11400 27435 11440 27467
rect 11472 27435 11512 27467
rect 11544 27435 11584 27467
rect 11616 27435 11656 27467
rect 11688 27435 11728 27467
rect 11760 27435 11800 27467
rect 11832 27435 11872 27467
rect 11904 27435 11944 27467
rect 11976 27435 12016 27467
rect 12048 27435 12088 27467
rect 12120 27435 12160 27467
rect 12192 27435 12232 27467
rect 12264 27435 12304 27467
rect 12336 27435 12376 27467
rect 12408 27435 12448 27467
rect 12480 27435 12520 27467
rect 12552 27435 12592 27467
rect 12624 27435 12664 27467
rect 12696 27435 12736 27467
rect 12768 27435 12808 27467
rect 12840 27435 12880 27467
rect 12912 27435 12952 27467
rect 12984 27435 13024 27467
rect 13056 27435 13096 27467
rect 13128 27435 13168 27467
rect 13200 27435 13240 27467
rect 13272 27435 13312 27467
rect 13344 27435 13384 27467
rect 13416 27435 13456 27467
rect 13488 27435 13528 27467
rect 13560 27435 13600 27467
rect 13632 27435 13672 27467
rect 13704 27435 13744 27467
rect 13776 27435 13816 27467
rect 13848 27435 13888 27467
rect 13920 27435 13960 27467
rect 13992 27435 14032 27467
rect 14064 27435 14104 27467
rect 14136 27435 14176 27467
rect 14208 27435 14248 27467
rect 14280 27435 14320 27467
rect 14352 27435 14392 27467
rect 14424 27435 14464 27467
rect 14496 27435 14536 27467
rect 14568 27435 14608 27467
rect 14640 27435 14680 27467
rect 14712 27435 14752 27467
rect 14784 27435 14824 27467
rect 14856 27435 14896 27467
rect 14928 27435 14968 27467
rect 15000 27435 15040 27467
rect 15072 27435 15112 27467
rect 15144 27435 15184 27467
rect 15216 27435 15256 27467
rect 15288 27435 15328 27467
rect 15360 27435 15400 27467
rect 15432 27435 15472 27467
rect 15504 27435 15544 27467
rect 15576 27435 15616 27467
rect 15648 27435 15688 27467
rect 15720 27435 15760 27467
rect 15792 27435 15832 27467
rect 15864 27435 15904 27467
rect 15936 27435 16000 27467
rect 0 27395 16000 27435
rect 0 27363 64 27395
rect 96 27363 136 27395
rect 168 27363 208 27395
rect 240 27363 280 27395
rect 312 27363 352 27395
rect 384 27363 424 27395
rect 456 27363 496 27395
rect 528 27363 568 27395
rect 600 27363 640 27395
rect 672 27363 712 27395
rect 744 27363 784 27395
rect 816 27363 856 27395
rect 888 27363 928 27395
rect 960 27363 1000 27395
rect 1032 27363 1072 27395
rect 1104 27363 1144 27395
rect 1176 27363 1216 27395
rect 1248 27363 1288 27395
rect 1320 27363 1360 27395
rect 1392 27363 1432 27395
rect 1464 27363 1504 27395
rect 1536 27363 1576 27395
rect 1608 27363 1648 27395
rect 1680 27363 1720 27395
rect 1752 27363 1792 27395
rect 1824 27363 1864 27395
rect 1896 27363 1936 27395
rect 1968 27363 2008 27395
rect 2040 27363 2080 27395
rect 2112 27363 2152 27395
rect 2184 27363 2224 27395
rect 2256 27363 2296 27395
rect 2328 27363 2368 27395
rect 2400 27363 2440 27395
rect 2472 27363 2512 27395
rect 2544 27363 2584 27395
rect 2616 27363 2656 27395
rect 2688 27363 2728 27395
rect 2760 27363 2800 27395
rect 2832 27363 2872 27395
rect 2904 27363 2944 27395
rect 2976 27363 3016 27395
rect 3048 27363 3088 27395
rect 3120 27363 3160 27395
rect 3192 27363 3232 27395
rect 3264 27363 3304 27395
rect 3336 27363 3376 27395
rect 3408 27363 3448 27395
rect 3480 27363 3520 27395
rect 3552 27363 3592 27395
rect 3624 27363 3664 27395
rect 3696 27363 3736 27395
rect 3768 27363 3808 27395
rect 3840 27363 3880 27395
rect 3912 27363 3952 27395
rect 3984 27363 4024 27395
rect 4056 27363 4096 27395
rect 4128 27363 4168 27395
rect 4200 27363 4240 27395
rect 4272 27363 4312 27395
rect 4344 27363 4384 27395
rect 4416 27363 4456 27395
rect 4488 27363 4528 27395
rect 4560 27363 4600 27395
rect 4632 27363 4672 27395
rect 4704 27363 4744 27395
rect 4776 27363 4816 27395
rect 4848 27363 4888 27395
rect 4920 27363 4960 27395
rect 4992 27363 5032 27395
rect 5064 27363 5104 27395
rect 5136 27363 5176 27395
rect 5208 27363 5248 27395
rect 5280 27363 5320 27395
rect 5352 27363 5392 27395
rect 5424 27363 5464 27395
rect 5496 27363 5536 27395
rect 5568 27363 5608 27395
rect 5640 27363 5680 27395
rect 5712 27363 5752 27395
rect 5784 27363 5824 27395
rect 5856 27363 5896 27395
rect 5928 27363 5968 27395
rect 6000 27363 6040 27395
rect 6072 27363 6112 27395
rect 6144 27363 6184 27395
rect 6216 27363 6256 27395
rect 6288 27363 6328 27395
rect 6360 27363 6400 27395
rect 6432 27363 6472 27395
rect 6504 27363 6544 27395
rect 6576 27363 6616 27395
rect 6648 27363 6688 27395
rect 6720 27363 6760 27395
rect 6792 27363 6832 27395
rect 6864 27363 6904 27395
rect 6936 27363 6976 27395
rect 7008 27363 7048 27395
rect 7080 27363 7120 27395
rect 7152 27363 7192 27395
rect 7224 27363 7264 27395
rect 7296 27363 7336 27395
rect 7368 27363 7408 27395
rect 7440 27363 7480 27395
rect 7512 27363 7552 27395
rect 7584 27363 7624 27395
rect 7656 27363 7696 27395
rect 7728 27363 7768 27395
rect 7800 27363 7840 27395
rect 7872 27363 7912 27395
rect 7944 27363 7984 27395
rect 8016 27363 8056 27395
rect 8088 27363 8128 27395
rect 8160 27363 8200 27395
rect 8232 27363 8272 27395
rect 8304 27363 8344 27395
rect 8376 27363 8416 27395
rect 8448 27363 8488 27395
rect 8520 27363 8560 27395
rect 8592 27363 8632 27395
rect 8664 27363 8704 27395
rect 8736 27363 8776 27395
rect 8808 27363 8848 27395
rect 8880 27363 8920 27395
rect 8952 27363 8992 27395
rect 9024 27363 9064 27395
rect 9096 27363 9136 27395
rect 9168 27363 9208 27395
rect 9240 27363 9280 27395
rect 9312 27363 9352 27395
rect 9384 27363 9424 27395
rect 9456 27363 9496 27395
rect 9528 27363 9568 27395
rect 9600 27363 9640 27395
rect 9672 27363 9712 27395
rect 9744 27363 9784 27395
rect 9816 27363 9856 27395
rect 9888 27363 9928 27395
rect 9960 27363 10000 27395
rect 10032 27363 10072 27395
rect 10104 27363 10144 27395
rect 10176 27363 10216 27395
rect 10248 27363 10288 27395
rect 10320 27363 10360 27395
rect 10392 27363 10432 27395
rect 10464 27363 10504 27395
rect 10536 27363 10576 27395
rect 10608 27363 10648 27395
rect 10680 27363 10720 27395
rect 10752 27363 10792 27395
rect 10824 27363 10864 27395
rect 10896 27363 10936 27395
rect 10968 27363 11008 27395
rect 11040 27363 11080 27395
rect 11112 27363 11152 27395
rect 11184 27363 11224 27395
rect 11256 27363 11296 27395
rect 11328 27363 11368 27395
rect 11400 27363 11440 27395
rect 11472 27363 11512 27395
rect 11544 27363 11584 27395
rect 11616 27363 11656 27395
rect 11688 27363 11728 27395
rect 11760 27363 11800 27395
rect 11832 27363 11872 27395
rect 11904 27363 11944 27395
rect 11976 27363 12016 27395
rect 12048 27363 12088 27395
rect 12120 27363 12160 27395
rect 12192 27363 12232 27395
rect 12264 27363 12304 27395
rect 12336 27363 12376 27395
rect 12408 27363 12448 27395
rect 12480 27363 12520 27395
rect 12552 27363 12592 27395
rect 12624 27363 12664 27395
rect 12696 27363 12736 27395
rect 12768 27363 12808 27395
rect 12840 27363 12880 27395
rect 12912 27363 12952 27395
rect 12984 27363 13024 27395
rect 13056 27363 13096 27395
rect 13128 27363 13168 27395
rect 13200 27363 13240 27395
rect 13272 27363 13312 27395
rect 13344 27363 13384 27395
rect 13416 27363 13456 27395
rect 13488 27363 13528 27395
rect 13560 27363 13600 27395
rect 13632 27363 13672 27395
rect 13704 27363 13744 27395
rect 13776 27363 13816 27395
rect 13848 27363 13888 27395
rect 13920 27363 13960 27395
rect 13992 27363 14032 27395
rect 14064 27363 14104 27395
rect 14136 27363 14176 27395
rect 14208 27363 14248 27395
rect 14280 27363 14320 27395
rect 14352 27363 14392 27395
rect 14424 27363 14464 27395
rect 14496 27363 14536 27395
rect 14568 27363 14608 27395
rect 14640 27363 14680 27395
rect 14712 27363 14752 27395
rect 14784 27363 14824 27395
rect 14856 27363 14896 27395
rect 14928 27363 14968 27395
rect 15000 27363 15040 27395
rect 15072 27363 15112 27395
rect 15144 27363 15184 27395
rect 15216 27363 15256 27395
rect 15288 27363 15328 27395
rect 15360 27363 15400 27395
rect 15432 27363 15472 27395
rect 15504 27363 15544 27395
rect 15576 27363 15616 27395
rect 15648 27363 15688 27395
rect 15720 27363 15760 27395
rect 15792 27363 15832 27395
rect 15864 27363 15904 27395
rect 15936 27363 16000 27395
rect 0 27323 16000 27363
rect 0 27291 64 27323
rect 96 27291 136 27323
rect 168 27291 208 27323
rect 240 27291 280 27323
rect 312 27291 352 27323
rect 384 27291 424 27323
rect 456 27291 496 27323
rect 528 27291 568 27323
rect 600 27291 640 27323
rect 672 27291 712 27323
rect 744 27291 784 27323
rect 816 27291 856 27323
rect 888 27291 928 27323
rect 960 27291 1000 27323
rect 1032 27291 1072 27323
rect 1104 27291 1144 27323
rect 1176 27291 1216 27323
rect 1248 27291 1288 27323
rect 1320 27291 1360 27323
rect 1392 27291 1432 27323
rect 1464 27291 1504 27323
rect 1536 27291 1576 27323
rect 1608 27291 1648 27323
rect 1680 27291 1720 27323
rect 1752 27291 1792 27323
rect 1824 27291 1864 27323
rect 1896 27291 1936 27323
rect 1968 27291 2008 27323
rect 2040 27291 2080 27323
rect 2112 27291 2152 27323
rect 2184 27291 2224 27323
rect 2256 27291 2296 27323
rect 2328 27291 2368 27323
rect 2400 27291 2440 27323
rect 2472 27291 2512 27323
rect 2544 27291 2584 27323
rect 2616 27291 2656 27323
rect 2688 27291 2728 27323
rect 2760 27291 2800 27323
rect 2832 27291 2872 27323
rect 2904 27291 2944 27323
rect 2976 27291 3016 27323
rect 3048 27291 3088 27323
rect 3120 27291 3160 27323
rect 3192 27291 3232 27323
rect 3264 27291 3304 27323
rect 3336 27291 3376 27323
rect 3408 27291 3448 27323
rect 3480 27291 3520 27323
rect 3552 27291 3592 27323
rect 3624 27291 3664 27323
rect 3696 27291 3736 27323
rect 3768 27291 3808 27323
rect 3840 27291 3880 27323
rect 3912 27291 3952 27323
rect 3984 27291 4024 27323
rect 4056 27291 4096 27323
rect 4128 27291 4168 27323
rect 4200 27291 4240 27323
rect 4272 27291 4312 27323
rect 4344 27291 4384 27323
rect 4416 27291 4456 27323
rect 4488 27291 4528 27323
rect 4560 27291 4600 27323
rect 4632 27291 4672 27323
rect 4704 27291 4744 27323
rect 4776 27291 4816 27323
rect 4848 27291 4888 27323
rect 4920 27291 4960 27323
rect 4992 27291 5032 27323
rect 5064 27291 5104 27323
rect 5136 27291 5176 27323
rect 5208 27291 5248 27323
rect 5280 27291 5320 27323
rect 5352 27291 5392 27323
rect 5424 27291 5464 27323
rect 5496 27291 5536 27323
rect 5568 27291 5608 27323
rect 5640 27291 5680 27323
rect 5712 27291 5752 27323
rect 5784 27291 5824 27323
rect 5856 27291 5896 27323
rect 5928 27291 5968 27323
rect 6000 27291 6040 27323
rect 6072 27291 6112 27323
rect 6144 27291 6184 27323
rect 6216 27291 6256 27323
rect 6288 27291 6328 27323
rect 6360 27291 6400 27323
rect 6432 27291 6472 27323
rect 6504 27291 6544 27323
rect 6576 27291 6616 27323
rect 6648 27291 6688 27323
rect 6720 27291 6760 27323
rect 6792 27291 6832 27323
rect 6864 27291 6904 27323
rect 6936 27291 6976 27323
rect 7008 27291 7048 27323
rect 7080 27291 7120 27323
rect 7152 27291 7192 27323
rect 7224 27291 7264 27323
rect 7296 27291 7336 27323
rect 7368 27291 7408 27323
rect 7440 27291 7480 27323
rect 7512 27291 7552 27323
rect 7584 27291 7624 27323
rect 7656 27291 7696 27323
rect 7728 27291 7768 27323
rect 7800 27291 7840 27323
rect 7872 27291 7912 27323
rect 7944 27291 7984 27323
rect 8016 27291 8056 27323
rect 8088 27291 8128 27323
rect 8160 27291 8200 27323
rect 8232 27291 8272 27323
rect 8304 27291 8344 27323
rect 8376 27291 8416 27323
rect 8448 27291 8488 27323
rect 8520 27291 8560 27323
rect 8592 27291 8632 27323
rect 8664 27291 8704 27323
rect 8736 27291 8776 27323
rect 8808 27291 8848 27323
rect 8880 27291 8920 27323
rect 8952 27291 8992 27323
rect 9024 27291 9064 27323
rect 9096 27291 9136 27323
rect 9168 27291 9208 27323
rect 9240 27291 9280 27323
rect 9312 27291 9352 27323
rect 9384 27291 9424 27323
rect 9456 27291 9496 27323
rect 9528 27291 9568 27323
rect 9600 27291 9640 27323
rect 9672 27291 9712 27323
rect 9744 27291 9784 27323
rect 9816 27291 9856 27323
rect 9888 27291 9928 27323
rect 9960 27291 10000 27323
rect 10032 27291 10072 27323
rect 10104 27291 10144 27323
rect 10176 27291 10216 27323
rect 10248 27291 10288 27323
rect 10320 27291 10360 27323
rect 10392 27291 10432 27323
rect 10464 27291 10504 27323
rect 10536 27291 10576 27323
rect 10608 27291 10648 27323
rect 10680 27291 10720 27323
rect 10752 27291 10792 27323
rect 10824 27291 10864 27323
rect 10896 27291 10936 27323
rect 10968 27291 11008 27323
rect 11040 27291 11080 27323
rect 11112 27291 11152 27323
rect 11184 27291 11224 27323
rect 11256 27291 11296 27323
rect 11328 27291 11368 27323
rect 11400 27291 11440 27323
rect 11472 27291 11512 27323
rect 11544 27291 11584 27323
rect 11616 27291 11656 27323
rect 11688 27291 11728 27323
rect 11760 27291 11800 27323
rect 11832 27291 11872 27323
rect 11904 27291 11944 27323
rect 11976 27291 12016 27323
rect 12048 27291 12088 27323
rect 12120 27291 12160 27323
rect 12192 27291 12232 27323
rect 12264 27291 12304 27323
rect 12336 27291 12376 27323
rect 12408 27291 12448 27323
rect 12480 27291 12520 27323
rect 12552 27291 12592 27323
rect 12624 27291 12664 27323
rect 12696 27291 12736 27323
rect 12768 27291 12808 27323
rect 12840 27291 12880 27323
rect 12912 27291 12952 27323
rect 12984 27291 13024 27323
rect 13056 27291 13096 27323
rect 13128 27291 13168 27323
rect 13200 27291 13240 27323
rect 13272 27291 13312 27323
rect 13344 27291 13384 27323
rect 13416 27291 13456 27323
rect 13488 27291 13528 27323
rect 13560 27291 13600 27323
rect 13632 27291 13672 27323
rect 13704 27291 13744 27323
rect 13776 27291 13816 27323
rect 13848 27291 13888 27323
rect 13920 27291 13960 27323
rect 13992 27291 14032 27323
rect 14064 27291 14104 27323
rect 14136 27291 14176 27323
rect 14208 27291 14248 27323
rect 14280 27291 14320 27323
rect 14352 27291 14392 27323
rect 14424 27291 14464 27323
rect 14496 27291 14536 27323
rect 14568 27291 14608 27323
rect 14640 27291 14680 27323
rect 14712 27291 14752 27323
rect 14784 27291 14824 27323
rect 14856 27291 14896 27323
rect 14928 27291 14968 27323
rect 15000 27291 15040 27323
rect 15072 27291 15112 27323
rect 15144 27291 15184 27323
rect 15216 27291 15256 27323
rect 15288 27291 15328 27323
rect 15360 27291 15400 27323
rect 15432 27291 15472 27323
rect 15504 27291 15544 27323
rect 15576 27291 15616 27323
rect 15648 27291 15688 27323
rect 15720 27291 15760 27323
rect 15792 27291 15832 27323
rect 15864 27291 15904 27323
rect 15936 27291 16000 27323
rect 0 27251 16000 27291
rect 0 27219 64 27251
rect 96 27219 136 27251
rect 168 27219 208 27251
rect 240 27219 280 27251
rect 312 27219 352 27251
rect 384 27219 424 27251
rect 456 27219 496 27251
rect 528 27219 568 27251
rect 600 27219 640 27251
rect 672 27219 712 27251
rect 744 27219 784 27251
rect 816 27219 856 27251
rect 888 27219 928 27251
rect 960 27219 1000 27251
rect 1032 27219 1072 27251
rect 1104 27219 1144 27251
rect 1176 27219 1216 27251
rect 1248 27219 1288 27251
rect 1320 27219 1360 27251
rect 1392 27219 1432 27251
rect 1464 27219 1504 27251
rect 1536 27219 1576 27251
rect 1608 27219 1648 27251
rect 1680 27219 1720 27251
rect 1752 27219 1792 27251
rect 1824 27219 1864 27251
rect 1896 27219 1936 27251
rect 1968 27219 2008 27251
rect 2040 27219 2080 27251
rect 2112 27219 2152 27251
rect 2184 27219 2224 27251
rect 2256 27219 2296 27251
rect 2328 27219 2368 27251
rect 2400 27219 2440 27251
rect 2472 27219 2512 27251
rect 2544 27219 2584 27251
rect 2616 27219 2656 27251
rect 2688 27219 2728 27251
rect 2760 27219 2800 27251
rect 2832 27219 2872 27251
rect 2904 27219 2944 27251
rect 2976 27219 3016 27251
rect 3048 27219 3088 27251
rect 3120 27219 3160 27251
rect 3192 27219 3232 27251
rect 3264 27219 3304 27251
rect 3336 27219 3376 27251
rect 3408 27219 3448 27251
rect 3480 27219 3520 27251
rect 3552 27219 3592 27251
rect 3624 27219 3664 27251
rect 3696 27219 3736 27251
rect 3768 27219 3808 27251
rect 3840 27219 3880 27251
rect 3912 27219 3952 27251
rect 3984 27219 4024 27251
rect 4056 27219 4096 27251
rect 4128 27219 4168 27251
rect 4200 27219 4240 27251
rect 4272 27219 4312 27251
rect 4344 27219 4384 27251
rect 4416 27219 4456 27251
rect 4488 27219 4528 27251
rect 4560 27219 4600 27251
rect 4632 27219 4672 27251
rect 4704 27219 4744 27251
rect 4776 27219 4816 27251
rect 4848 27219 4888 27251
rect 4920 27219 4960 27251
rect 4992 27219 5032 27251
rect 5064 27219 5104 27251
rect 5136 27219 5176 27251
rect 5208 27219 5248 27251
rect 5280 27219 5320 27251
rect 5352 27219 5392 27251
rect 5424 27219 5464 27251
rect 5496 27219 5536 27251
rect 5568 27219 5608 27251
rect 5640 27219 5680 27251
rect 5712 27219 5752 27251
rect 5784 27219 5824 27251
rect 5856 27219 5896 27251
rect 5928 27219 5968 27251
rect 6000 27219 6040 27251
rect 6072 27219 6112 27251
rect 6144 27219 6184 27251
rect 6216 27219 6256 27251
rect 6288 27219 6328 27251
rect 6360 27219 6400 27251
rect 6432 27219 6472 27251
rect 6504 27219 6544 27251
rect 6576 27219 6616 27251
rect 6648 27219 6688 27251
rect 6720 27219 6760 27251
rect 6792 27219 6832 27251
rect 6864 27219 6904 27251
rect 6936 27219 6976 27251
rect 7008 27219 7048 27251
rect 7080 27219 7120 27251
rect 7152 27219 7192 27251
rect 7224 27219 7264 27251
rect 7296 27219 7336 27251
rect 7368 27219 7408 27251
rect 7440 27219 7480 27251
rect 7512 27219 7552 27251
rect 7584 27219 7624 27251
rect 7656 27219 7696 27251
rect 7728 27219 7768 27251
rect 7800 27219 7840 27251
rect 7872 27219 7912 27251
rect 7944 27219 7984 27251
rect 8016 27219 8056 27251
rect 8088 27219 8128 27251
rect 8160 27219 8200 27251
rect 8232 27219 8272 27251
rect 8304 27219 8344 27251
rect 8376 27219 8416 27251
rect 8448 27219 8488 27251
rect 8520 27219 8560 27251
rect 8592 27219 8632 27251
rect 8664 27219 8704 27251
rect 8736 27219 8776 27251
rect 8808 27219 8848 27251
rect 8880 27219 8920 27251
rect 8952 27219 8992 27251
rect 9024 27219 9064 27251
rect 9096 27219 9136 27251
rect 9168 27219 9208 27251
rect 9240 27219 9280 27251
rect 9312 27219 9352 27251
rect 9384 27219 9424 27251
rect 9456 27219 9496 27251
rect 9528 27219 9568 27251
rect 9600 27219 9640 27251
rect 9672 27219 9712 27251
rect 9744 27219 9784 27251
rect 9816 27219 9856 27251
rect 9888 27219 9928 27251
rect 9960 27219 10000 27251
rect 10032 27219 10072 27251
rect 10104 27219 10144 27251
rect 10176 27219 10216 27251
rect 10248 27219 10288 27251
rect 10320 27219 10360 27251
rect 10392 27219 10432 27251
rect 10464 27219 10504 27251
rect 10536 27219 10576 27251
rect 10608 27219 10648 27251
rect 10680 27219 10720 27251
rect 10752 27219 10792 27251
rect 10824 27219 10864 27251
rect 10896 27219 10936 27251
rect 10968 27219 11008 27251
rect 11040 27219 11080 27251
rect 11112 27219 11152 27251
rect 11184 27219 11224 27251
rect 11256 27219 11296 27251
rect 11328 27219 11368 27251
rect 11400 27219 11440 27251
rect 11472 27219 11512 27251
rect 11544 27219 11584 27251
rect 11616 27219 11656 27251
rect 11688 27219 11728 27251
rect 11760 27219 11800 27251
rect 11832 27219 11872 27251
rect 11904 27219 11944 27251
rect 11976 27219 12016 27251
rect 12048 27219 12088 27251
rect 12120 27219 12160 27251
rect 12192 27219 12232 27251
rect 12264 27219 12304 27251
rect 12336 27219 12376 27251
rect 12408 27219 12448 27251
rect 12480 27219 12520 27251
rect 12552 27219 12592 27251
rect 12624 27219 12664 27251
rect 12696 27219 12736 27251
rect 12768 27219 12808 27251
rect 12840 27219 12880 27251
rect 12912 27219 12952 27251
rect 12984 27219 13024 27251
rect 13056 27219 13096 27251
rect 13128 27219 13168 27251
rect 13200 27219 13240 27251
rect 13272 27219 13312 27251
rect 13344 27219 13384 27251
rect 13416 27219 13456 27251
rect 13488 27219 13528 27251
rect 13560 27219 13600 27251
rect 13632 27219 13672 27251
rect 13704 27219 13744 27251
rect 13776 27219 13816 27251
rect 13848 27219 13888 27251
rect 13920 27219 13960 27251
rect 13992 27219 14032 27251
rect 14064 27219 14104 27251
rect 14136 27219 14176 27251
rect 14208 27219 14248 27251
rect 14280 27219 14320 27251
rect 14352 27219 14392 27251
rect 14424 27219 14464 27251
rect 14496 27219 14536 27251
rect 14568 27219 14608 27251
rect 14640 27219 14680 27251
rect 14712 27219 14752 27251
rect 14784 27219 14824 27251
rect 14856 27219 14896 27251
rect 14928 27219 14968 27251
rect 15000 27219 15040 27251
rect 15072 27219 15112 27251
rect 15144 27219 15184 27251
rect 15216 27219 15256 27251
rect 15288 27219 15328 27251
rect 15360 27219 15400 27251
rect 15432 27219 15472 27251
rect 15504 27219 15544 27251
rect 15576 27219 15616 27251
rect 15648 27219 15688 27251
rect 15720 27219 15760 27251
rect 15792 27219 15832 27251
rect 15864 27219 15904 27251
rect 15936 27219 16000 27251
rect 0 27179 16000 27219
rect 0 27147 64 27179
rect 96 27147 136 27179
rect 168 27147 208 27179
rect 240 27147 280 27179
rect 312 27147 352 27179
rect 384 27147 424 27179
rect 456 27147 496 27179
rect 528 27147 568 27179
rect 600 27147 640 27179
rect 672 27147 712 27179
rect 744 27147 784 27179
rect 816 27147 856 27179
rect 888 27147 928 27179
rect 960 27147 1000 27179
rect 1032 27147 1072 27179
rect 1104 27147 1144 27179
rect 1176 27147 1216 27179
rect 1248 27147 1288 27179
rect 1320 27147 1360 27179
rect 1392 27147 1432 27179
rect 1464 27147 1504 27179
rect 1536 27147 1576 27179
rect 1608 27147 1648 27179
rect 1680 27147 1720 27179
rect 1752 27147 1792 27179
rect 1824 27147 1864 27179
rect 1896 27147 1936 27179
rect 1968 27147 2008 27179
rect 2040 27147 2080 27179
rect 2112 27147 2152 27179
rect 2184 27147 2224 27179
rect 2256 27147 2296 27179
rect 2328 27147 2368 27179
rect 2400 27147 2440 27179
rect 2472 27147 2512 27179
rect 2544 27147 2584 27179
rect 2616 27147 2656 27179
rect 2688 27147 2728 27179
rect 2760 27147 2800 27179
rect 2832 27147 2872 27179
rect 2904 27147 2944 27179
rect 2976 27147 3016 27179
rect 3048 27147 3088 27179
rect 3120 27147 3160 27179
rect 3192 27147 3232 27179
rect 3264 27147 3304 27179
rect 3336 27147 3376 27179
rect 3408 27147 3448 27179
rect 3480 27147 3520 27179
rect 3552 27147 3592 27179
rect 3624 27147 3664 27179
rect 3696 27147 3736 27179
rect 3768 27147 3808 27179
rect 3840 27147 3880 27179
rect 3912 27147 3952 27179
rect 3984 27147 4024 27179
rect 4056 27147 4096 27179
rect 4128 27147 4168 27179
rect 4200 27147 4240 27179
rect 4272 27147 4312 27179
rect 4344 27147 4384 27179
rect 4416 27147 4456 27179
rect 4488 27147 4528 27179
rect 4560 27147 4600 27179
rect 4632 27147 4672 27179
rect 4704 27147 4744 27179
rect 4776 27147 4816 27179
rect 4848 27147 4888 27179
rect 4920 27147 4960 27179
rect 4992 27147 5032 27179
rect 5064 27147 5104 27179
rect 5136 27147 5176 27179
rect 5208 27147 5248 27179
rect 5280 27147 5320 27179
rect 5352 27147 5392 27179
rect 5424 27147 5464 27179
rect 5496 27147 5536 27179
rect 5568 27147 5608 27179
rect 5640 27147 5680 27179
rect 5712 27147 5752 27179
rect 5784 27147 5824 27179
rect 5856 27147 5896 27179
rect 5928 27147 5968 27179
rect 6000 27147 6040 27179
rect 6072 27147 6112 27179
rect 6144 27147 6184 27179
rect 6216 27147 6256 27179
rect 6288 27147 6328 27179
rect 6360 27147 6400 27179
rect 6432 27147 6472 27179
rect 6504 27147 6544 27179
rect 6576 27147 6616 27179
rect 6648 27147 6688 27179
rect 6720 27147 6760 27179
rect 6792 27147 6832 27179
rect 6864 27147 6904 27179
rect 6936 27147 6976 27179
rect 7008 27147 7048 27179
rect 7080 27147 7120 27179
rect 7152 27147 7192 27179
rect 7224 27147 7264 27179
rect 7296 27147 7336 27179
rect 7368 27147 7408 27179
rect 7440 27147 7480 27179
rect 7512 27147 7552 27179
rect 7584 27147 7624 27179
rect 7656 27147 7696 27179
rect 7728 27147 7768 27179
rect 7800 27147 7840 27179
rect 7872 27147 7912 27179
rect 7944 27147 7984 27179
rect 8016 27147 8056 27179
rect 8088 27147 8128 27179
rect 8160 27147 8200 27179
rect 8232 27147 8272 27179
rect 8304 27147 8344 27179
rect 8376 27147 8416 27179
rect 8448 27147 8488 27179
rect 8520 27147 8560 27179
rect 8592 27147 8632 27179
rect 8664 27147 8704 27179
rect 8736 27147 8776 27179
rect 8808 27147 8848 27179
rect 8880 27147 8920 27179
rect 8952 27147 8992 27179
rect 9024 27147 9064 27179
rect 9096 27147 9136 27179
rect 9168 27147 9208 27179
rect 9240 27147 9280 27179
rect 9312 27147 9352 27179
rect 9384 27147 9424 27179
rect 9456 27147 9496 27179
rect 9528 27147 9568 27179
rect 9600 27147 9640 27179
rect 9672 27147 9712 27179
rect 9744 27147 9784 27179
rect 9816 27147 9856 27179
rect 9888 27147 9928 27179
rect 9960 27147 10000 27179
rect 10032 27147 10072 27179
rect 10104 27147 10144 27179
rect 10176 27147 10216 27179
rect 10248 27147 10288 27179
rect 10320 27147 10360 27179
rect 10392 27147 10432 27179
rect 10464 27147 10504 27179
rect 10536 27147 10576 27179
rect 10608 27147 10648 27179
rect 10680 27147 10720 27179
rect 10752 27147 10792 27179
rect 10824 27147 10864 27179
rect 10896 27147 10936 27179
rect 10968 27147 11008 27179
rect 11040 27147 11080 27179
rect 11112 27147 11152 27179
rect 11184 27147 11224 27179
rect 11256 27147 11296 27179
rect 11328 27147 11368 27179
rect 11400 27147 11440 27179
rect 11472 27147 11512 27179
rect 11544 27147 11584 27179
rect 11616 27147 11656 27179
rect 11688 27147 11728 27179
rect 11760 27147 11800 27179
rect 11832 27147 11872 27179
rect 11904 27147 11944 27179
rect 11976 27147 12016 27179
rect 12048 27147 12088 27179
rect 12120 27147 12160 27179
rect 12192 27147 12232 27179
rect 12264 27147 12304 27179
rect 12336 27147 12376 27179
rect 12408 27147 12448 27179
rect 12480 27147 12520 27179
rect 12552 27147 12592 27179
rect 12624 27147 12664 27179
rect 12696 27147 12736 27179
rect 12768 27147 12808 27179
rect 12840 27147 12880 27179
rect 12912 27147 12952 27179
rect 12984 27147 13024 27179
rect 13056 27147 13096 27179
rect 13128 27147 13168 27179
rect 13200 27147 13240 27179
rect 13272 27147 13312 27179
rect 13344 27147 13384 27179
rect 13416 27147 13456 27179
rect 13488 27147 13528 27179
rect 13560 27147 13600 27179
rect 13632 27147 13672 27179
rect 13704 27147 13744 27179
rect 13776 27147 13816 27179
rect 13848 27147 13888 27179
rect 13920 27147 13960 27179
rect 13992 27147 14032 27179
rect 14064 27147 14104 27179
rect 14136 27147 14176 27179
rect 14208 27147 14248 27179
rect 14280 27147 14320 27179
rect 14352 27147 14392 27179
rect 14424 27147 14464 27179
rect 14496 27147 14536 27179
rect 14568 27147 14608 27179
rect 14640 27147 14680 27179
rect 14712 27147 14752 27179
rect 14784 27147 14824 27179
rect 14856 27147 14896 27179
rect 14928 27147 14968 27179
rect 15000 27147 15040 27179
rect 15072 27147 15112 27179
rect 15144 27147 15184 27179
rect 15216 27147 15256 27179
rect 15288 27147 15328 27179
rect 15360 27147 15400 27179
rect 15432 27147 15472 27179
rect 15504 27147 15544 27179
rect 15576 27147 15616 27179
rect 15648 27147 15688 27179
rect 15720 27147 15760 27179
rect 15792 27147 15832 27179
rect 15864 27147 15904 27179
rect 15936 27147 16000 27179
rect 0 27107 16000 27147
rect 0 27075 64 27107
rect 96 27075 136 27107
rect 168 27075 208 27107
rect 240 27075 280 27107
rect 312 27075 352 27107
rect 384 27075 424 27107
rect 456 27075 496 27107
rect 528 27075 568 27107
rect 600 27075 640 27107
rect 672 27075 712 27107
rect 744 27075 784 27107
rect 816 27075 856 27107
rect 888 27075 928 27107
rect 960 27075 1000 27107
rect 1032 27075 1072 27107
rect 1104 27075 1144 27107
rect 1176 27075 1216 27107
rect 1248 27075 1288 27107
rect 1320 27075 1360 27107
rect 1392 27075 1432 27107
rect 1464 27075 1504 27107
rect 1536 27075 1576 27107
rect 1608 27075 1648 27107
rect 1680 27075 1720 27107
rect 1752 27075 1792 27107
rect 1824 27075 1864 27107
rect 1896 27075 1936 27107
rect 1968 27075 2008 27107
rect 2040 27075 2080 27107
rect 2112 27075 2152 27107
rect 2184 27075 2224 27107
rect 2256 27075 2296 27107
rect 2328 27075 2368 27107
rect 2400 27075 2440 27107
rect 2472 27075 2512 27107
rect 2544 27075 2584 27107
rect 2616 27075 2656 27107
rect 2688 27075 2728 27107
rect 2760 27075 2800 27107
rect 2832 27075 2872 27107
rect 2904 27075 2944 27107
rect 2976 27075 3016 27107
rect 3048 27075 3088 27107
rect 3120 27075 3160 27107
rect 3192 27075 3232 27107
rect 3264 27075 3304 27107
rect 3336 27075 3376 27107
rect 3408 27075 3448 27107
rect 3480 27075 3520 27107
rect 3552 27075 3592 27107
rect 3624 27075 3664 27107
rect 3696 27075 3736 27107
rect 3768 27075 3808 27107
rect 3840 27075 3880 27107
rect 3912 27075 3952 27107
rect 3984 27075 4024 27107
rect 4056 27075 4096 27107
rect 4128 27075 4168 27107
rect 4200 27075 4240 27107
rect 4272 27075 4312 27107
rect 4344 27075 4384 27107
rect 4416 27075 4456 27107
rect 4488 27075 4528 27107
rect 4560 27075 4600 27107
rect 4632 27075 4672 27107
rect 4704 27075 4744 27107
rect 4776 27075 4816 27107
rect 4848 27075 4888 27107
rect 4920 27075 4960 27107
rect 4992 27075 5032 27107
rect 5064 27075 5104 27107
rect 5136 27075 5176 27107
rect 5208 27075 5248 27107
rect 5280 27075 5320 27107
rect 5352 27075 5392 27107
rect 5424 27075 5464 27107
rect 5496 27075 5536 27107
rect 5568 27075 5608 27107
rect 5640 27075 5680 27107
rect 5712 27075 5752 27107
rect 5784 27075 5824 27107
rect 5856 27075 5896 27107
rect 5928 27075 5968 27107
rect 6000 27075 6040 27107
rect 6072 27075 6112 27107
rect 6144 27075 6184 27107
rect 6216 27075 6256 27107
rect 6288 27075 6328 27107
rect 6360 27075 6400 27107
rect 6432 27075 6472 27107
rect 6504 27075 6544 27107
rect 6576 27075 6616 27107
rect 6648 27075 6688 27107
rect 6720 27075 6760 27107
rect 6792 27075 6832 27107
rect 6864 27075 6904 27107
rect 6936 27075 6976 27107
rect 7008 27075 7048 27107
rect 7080 27075 7120 27107
rect 7152 27075 7192 27107
rect 7224 27075 7264 27107
rect 7296 27075 7336 27107
rect 7368 27075 7408 27107
rect 7440 27075 7480 27107
rect 7512 27075 7552 27107
rect 7584 27075 7624 27107
rect 7656 27075 7696 27107
rect 7728 27075 7768 27107
rect 7800 27075 7840 27107
rect 7872 27075 7912 27107
rect 7944 27075 7984 27107
rect 8016 27075 8056 27107
rect 8088 27075 8128 27107
rect 8160 27075 8200 27107
rect 8232 27075 8272 27107
rect 8304 27075 8344 27107
rect 8376 27075 8416 27107
rect 8448 27075 8488 27107
rect 8520 27075 8560 27107
rect 8592 27075 8632 27107
rect 8664 27075 8704 27107
rect 8736 27075 8776 27107
rect 8808 27075 8848 27107
rect 8880 27075 8920 27107
rect 8952 27075 8992 27107
rect 9024 27075 9064 27107
rect 9096 27075 9136 27107
rect 9168 27075 9208 27107
rect 9240 27075 9280 27107
rect 9312 27075 9352 27107
rect 9384 27075 9424 27107
rect 9456 27075 9496 27107
rect 9528 27075 9568 27107
rect 9600 27075 9640 27107
rect 9672 27075 9712 27107
rect 9744 27075 9784 27107
rect 9816 27075 9856 27107
rect 9888 27075 9928 27107
rect 9960 27075 10000 27107
rect 10032 27075 10072 27107
rect 10104 27075 10144 27107
rect 10176 27075 10216 27107
rect 10248 27075 10288 27107
rect 10320 27075 10360 27107
rect 10392 27075 10432 27107
rect 10464 27075 10504 27107
rect 10536 27075 10576 27107
rect 10608 27075 10648 27107
rect 10680 27075 10720 27107
rect 10752 27075 10792 27107
rect 10824 27075 10864 27107
rect 10896 27075 10936 27107
rect 10968 27075 11008 27107
rect 11040 27075 11080 27107
rect 11112 27075 11152 27107
rect 11184 27075 11224 27107
rect 11256 27075 11296 27107
rect 11328 27075 11368 27107
rect 11400 27075 11440 27107
rect 11472 27075 11512 27107
rect 11544 27075 11584 27107
rect 11616 27075 11656 27107
rect 11688 27075 11728 27107
rect 11760 27075 11800 27107
rect 11832 27075 11872 27107
rect 11904 27075 11944 27107
rect 11976 27075 12016 27107
rect 12048 27075 12088 27107
rect 12120 27075 12160 27107
rect 12192 27075 12232 27107
rect 12264 27075 12304 27107
rect 12336 27075 12376 27107
rect 12408 27075 12448 27107
rect 12480 27075 12520 27107
rect 12552 27075 12592 27107
rect 12624 27075 12664 27107
rect 12696 27075 12736 27107
rect 12768 27075 12808 27107
rect 12840 27075 12880 27107
rect 12912 27075 12952 27107
rect 12984 27075 13024 27107
rect 13056 27075 13096 27107
rect 13128 27075 13168 27107
rect 13200 27075 13240 27107
rect 13272 27075 13312 27107
rect 13344 27075 13384 27107
rect 13416 27075 13456 27107
rect 13488 27075 13528 27107
rect 13560 27075 13600 27107
rect 13632 27075 13672 27107
rect 13704 27075 13744 27107
rect 13776 27075 13816 27107
rect 13848 27075 13888 27107
rect 13920 27075 13960 27107
rect 13992 27075 14032 27107
rect 14064 27075 14104 27107
rect 14136 27075 14176 27107
rect 14208 27075 14248 27107
rect 14280 27075 14320 27107
rect 14352 27075 14392 27107
rect 14424 27075 14464 27107
rect 14496 27075 14536 27107
rect 14568 27075 14608 27107
rect 14640 27075 14680 27107
rect 14712 27075 14752 27107
rect 14784 27075 14824 27107
rect 14856 27075 14896 27107
rect 14928 27075 14968 27107
rect 15000 27075 15040 27107
rect 15072 27075 15112 27107
rect 15144 27075 15184 27107
rect 15216 27075 15256 27107
rect 15288 27075 15328 27107
rect 15360 27075 15400 27107
rect 15432 27075 15472 27107
rect 15504 27075 15544 27107
rect 15576 27075 15616 27107
rect 15648 27075 15688 27107
rect 15720 27075 15760 27107
rect 15792 27075 15832 27107
rect 15864 27075 15904 27107
rect 15936 27075 16000 27107
rect 0 27035 16000 27075
rect 0 27003 64 27035
rect 96 27003 136 27035
rect 168 27003 208 27035
rect 240 27003 280 27035
rect 312 27003 352 27035
rect 384 27003 424 27035
rect 456 27003 496 27035
rect 528 27003 568 27035
rect 600 27003 640 27035
rect 672 27003 712 27035
rect 744 27003 784 27035
rect 816 27003 856 27035
rect 888 27003 928 27035
rect 960 27003 1000 27035
rect 1032 27003 1072 27035
rect 1104 27003 1144 27035
rect 1176 27003 1216 27035
rect 1248 27003 1288 27035
rect 1320 27003 1360 27035
rect 1392 27003 1432 27035
rect 1464 27003 1504 27035
rect 1536 27003 1576 27035
rect 1608 27003 1648 27035
rect 1680 27003 1720 27035
rect 1752 27003 1792 27035
rect 1824 27003 1864 27035
rect 1896 27003 1936 27035
rect 1968 27003 2008 27035
rect 2040 27003 2080 27035
rect 2112 27003 2152 27035
rect 2184 27003 2224 27035
rect 2256 27003 2296 27035
rect 2328 27003 2368 27035
rect 2400 27003 2440 27035
rect 2472 27003 2512 27035
rect 2544 27003 2584 27035
rect 2616 27003 2656 27035
rect 2688 27003 2728 27035
rect 2760 27003 2800 27035
rect 2832 27003 2872 27035
rect 2904 27003 2944 27035
rect 2976 27003 3016 27035
rect 3048 27003 3088 27035
rect 3120 27003 3160 27035
rect 3192 27003 3232 27035
rect 3264 27003 3304 27035
rect 3336 27003 3376 27035
rect 3408 27003 3448 27035
rect 3480 27003 3520 27035
rect 3552 27003 3592 27035
rect 3624 27003 3664 27035
rect 3696 27003 3736 27035
rect 3768 27003 3808 27035
rect 3840 27003 3880 27035
rect 3912 27003 3952 27035
rect 3984 27003 4024 27035
rect 4056 27003 4096 27035
rect 4128 27003 4168 27035
rect 4200 27003 4240 27035
rect 4272 27003 4312 27035
rect 4344 27003 4384 27035
rect 4416 27003 4456 27035
rect 4488 27003 4528 27035
rect 4560 27003 4600 27035
rect 4632 27003 4672 27035
rect 4704 27003 4744 27035
rect 4776 27003 4816 27035
rect 4848 27003 4888 27035
rect 4920 27003 4960 27035
rect 4992 27003 5032 27035
rect 5064 27003 5104 27035
rect 5136 27003 5176 27035
rect 5208 27003 5248 27035
rect 5280 27003 5320 27035
rect 5352 27003 5392 27035
rect 5424 27003 5464 27035
rect 5496 27003 5536 27035
rect 5568 27003 5608 27035
rect 5640 27003 5680 27035
rect 5712 27003 5752 27035
rect 5784 27003 5824 27035
rect 5856 27003 5896 27035
rect 5928 27003 5968 27035
rect 6000 27003 6040 27035
rect 6072 27003 6112 27035
rect 6144 27003 6184 27035
rect 6216 27003 6256 27035
rect 6288 27003 6328 27035
rect 6360 27003 6400 27035
rect 6432 27003 6472 27035
rect 6504 27003 6544 27035
rect 6576 27003 6616 27035
rect 6648 27003 6688 27035
rect 6720 27003 6760 27035
rect 6792 27003 6832 27035
rect 6864 27003 6904 27035
rect 6936 27003 6976 27035
rect 7008 27003 7048 27035
rect 7080 27003 7120 27035
rect 7152 27003 7192 27035
rect 7224 27003 7264 27035
rect 7296 27003 7336 27035
rect 7368 27003 7408 27035
rect 7440 27003 7480 27035
rect 7512 27003 7552 27035
rect 7584 27003 7624 27035
rect 7656 27003 7696 27035
rect 7728 27003 7768 27035
rect 7800 27003 7840 27035
rect 7872 27003 7912 27035
rect 7944 27003 7984 27035
rect 8016 27003 8056 27035
rect 8088 27003 8128 27035
rect 8160 27003 8200 27035
rect 8232 27003 8272 27035
rect 8304 27003 8344 27035
rect 8376 27003 8416 27035
rect 8448 27003 8488 27035
rect 8520 27003 8560 27035
rect 8592 27003 8632 27035
rect 8664 27003 8704 27035
rect 8736 27003 8776 27035
rect 8808 27003 8848 27035
rect 8880 27003 8920 27035
rect 8952 27003 8992 27035
rect 9024 27003 9064 27035
rect 9096 27003 9136 27035
rect 9168 27003 9208 27035
rect 9240 27003 9280 27035
rect 9312 27003 9352 27035
rect 9384 27003 9424 27035
rect 9456 27003 9496 27035
rect 9528 27003 9568 27035
rect 9600 27003 9640 27035
rect 9672 27003 9712 27035
rect 9744 27003 9784 27035
rect 9816 27003 9856 27035
rect 9888 27003 9928 27035
rect 9960 27003 10000 27035
rect 10032 27003 10072 27035
rect 10104 27003 10144 27035
rect 10176 27003 10216 27035
rect 10248 27003 10288 27035
rect 10320 27003 10360 27035
rect 10392 27003 10432 27035
rect 10464 27003 10504 27035
rect 10536 27003 10576 27035
rect 10608 27003 10648 27035
rect 10680 27003 10720 27035
rect 10752 27003 10792 27035
rect 10824 27003 10864 27035
rect 10896 27003 10936 27035
rect 10968 27003 11008 27035
rect 11040 27003 11080 27035
rect 11112 27003 11152 27035
rect 11184 27003 11224 27035
rect 11256 27003 11296 27035
rect 11328 27003 11368 27035
rect 11400 27003 11440 27035
rect 11472 27003 11512 27035
rect 11544 27003 11584 27035
rect 11616 27003 11656 27035
rect 11688 27003 11728 27035
rect 11760 27003 11800 27035
rect 11832 27003 11872 27035
rect 11904 27003 11944 27035
rect 11976 27003 12016 27035
rect 12048 27003 12088 27035
rect 12120 27003 12160 27035
rect 12192 27003 12232 27035
rect 12264 27003 12304 27035
rect 12336 27003 12376 27035
rect 12408 27003 12448 27035
rect 12480 27003 12520 27035
rect 12552 27003 12592 27035
rect 12624 27003 12664 27035
rect 12696 27003 12736 27035
rect 12768 27003 12808 27035
rect 12840 27003 12880 27035
rect 12912 27003 12952 27035
rect 12984 27003 13024 27035
rect 13056 27003 13096 27035
rect 13128 27003 13168 27035
rect 13200 27003 13240 27035
rect 13272 27003 13312 27035
rect 13344 27003 13384 27035
rect 13416 27003 13456 27035
rect 13488 27003 13528 27035
rect 13560 27003 13600 27035
rect 13632 27003 13672 27035
rect 13704 27003 13744 27035
rect 13776 27003 13816 27035
rect 13848 27003 13888 27035
rect 13920 27003 13960 27035
rect 13992 27003 14032 27035
rect 14064 27003 14104 27035
rect 14136 27003 14176 27035
rect 14208 27003 14248 27035
rect 14280 27003 14320 27035
rect 14352 27003 14392 27035
rect 14424 27003 14464 27035
rect 14496 27003 14536 27035
rect 14568 27003 14608 27035
rect 14640 27003 14680 27035
rect 14712 27003 14752 27035
rect 14784 27003 14824 27035
rect 14856 27003 14896 27035
rect 14928 27003 14968 27035
rect 15000 27003 15040 27035
rect 15072 27003 15112 27035
rect 15144 27003 15184 27035
rect 15216 27003 15256 27035
rect 15288 27003 15328 27035
rect 15360 27003 15400 27035
rect 15432 27003 15472 27035
rect 15504 27003 15544 27035
rect 15576 27003 15616 27035
rect 15648 27003 15688 27035
rect 15720 27003 15760 27035
rect 15792 27003 15832 27035
rect 15864 27003 15904 27035
rect 15936 27003 16000 27035
rect 0 26963 16000 27003
rect 0 26931 64 26963
rect 96 26931 136 26963
rect 168 26931 208 26963
rect 240 26931 280 26963
rect 312 26931 352 26963
rect 384 26931 424 26963
rect 456 26931 496 26963
rect 528 26931 568 26963
rect 600 26931 640 26963
rect 672 26931 712 26963
rect 744 26931 784 26963
rect 816 26931 856 26963
rect 888 26931 928 26963
rect 960 26931 1000 26963
rect 1032 26931 1072 26963
rect 1104 26931 1144 26963
rect 1176 26931 1216 26963
rect 1248 26931 1288 26963
rect 1320 26931 1360 26963
rect 1392 26931 1432 26963
rect 1464 26931 1504 26963
rect 1536 26931 1576 26963
rect 1608 26931 1648 26963
rect 1680 26931 1720 26963
rect 1752 26931 1792 26963
rect 1824 26931 1864 26963
rect 1896 26931 1936 26963
rect 1968 26931 2008 26963
rect 2040 26931 2080 26963
rect 2112 26931 2152 26963
rect 2184 26931 2224 26963
rect 2256 26931 2296 26963
rect 2328 26931 2368 26963
rect 2400 26931 2440 26963
rect 2472 26931 2512 26963
rect 2544 26931 2584 26963
rect 2616 26931 2656 26963
rect 2688 26931 2728 26963
rect 2760 26931 2800 26963
rect 2832 26931 2872 26963
rect 2904 26931 2944 26963
rect 2976 26931 3016 26963
rect 3048 26931 3088 26963
rect 3120 26931 3160 26963
rect 3192 26931 3232 26963
rect 3264 26931 3304 26963
rect 3336 26931 3376 26963
rect 3408 26931 3448 26963
rect 3480 26931 3520 26963
rect 3552 26931 3592 26963
rect 3624 26931 3664 26963
rect 3696 26931 3736 26963
rect 3768 26931 3808 26963
rect 3840 26931 3880 26963
rect 3912 26931 3952 26963
rect 3984 26931 4024 26963
rect 4056 26931 4096 26963
rect 4128 26931 4168 26963
rect 4200 26931 4240 26963
rect 4272 26931 4312 26963
rect 4344 26931 4384 26963
rect 4416 26931 4456 26963
rect 4488 26931 4528 26963
rect 4560 26931 4600 26963
rect 4632 26931 4672 26963
rect 4704 26931 4744 26963
rect 4776 26931 4816 26963
rect 4848 26931 4888 26963
rect 4920 26931 4960 26963
rect 4992 26931 5032 26963
rect 5064 26931 5104 26963
rect 5136 26931 5176 26963
rect 5208 26931 5248 26963
rect 5280 26931 5320 26963
rect 5352 26931 5392 26963
rect 5424 26931 5464 26963
rect 5496 26931 5536 26963
rect 5568 26931 5608 26963
rect 5640 26931 5680 26963
rect 5712 26931 5752 26963
rect 5784 26931 5824 26963
rect 5856 26931 5896 26963
rect 5928 26931 5968 26963
rect 6000 26931 6040 26963
rect 6072 26931 6112 26963
rect 6144 26931 6184 26963
rect 6216 26931 6256 26963
rect 6288 26931 6328 26963
rect 6360 26931 6400 26963
rect 6432 26931 6472 26963
rect 6504 26931 6544 26963
rect 6576 26931 6616 26963
rect 6648 26931 6688 26963
rect 6720 26931 6760 26963
rect 6792 26931 6832 26963
rect 6864 26931 6904 26963
rect 6936 26931 6976 26963
rect 7008 26931 7048 26963
rect 7080 26931 7120 26963
rect 7152 26931 7192 26963
rect 7224 26931 7264 26963
rect 7296 26931 7336 26963
rect 7368 26931 7408 26963
rect 7440 26931 7480 26963
rect 7512 26931 7552 26963
rect 7584 26931 7624 26963
rect 7656 26931 7696 26963
rect 7728 26931 7768 26963
rect 7800 26931 7840 26963
rect 7872 26931 7912 26963
rect 7944 26931 7984 26963
rect 8016 26931 8056 26963
rect 8088 26931 8128 26963
rect 8160 26931 8200 26963
rect 8232 26931 8272 26963
rect 8304 26931 8344 26963
rect 8376 26931 8416 26963
rect 8448 26931 8488 26963
rect 8520 26931 8560 26963
rect 8592 26931 8632 26963
rect 8664 26931 8704 26963
rect 8736 26931 8776 26963
rect 8808 26931 8848 26963
rect 8880 26931 8920 26963
rect 8952 26931 8992 26963
rect 9024 26931 9064 26963
rect 9096 26931 9136 26963
rect 9168 26931 9208 26963
rect 9240 26931 9280 26963
rect 9312 26931 9352 26963
rect 9384 26931 9424 26963
rect 9456 26931 9496 26963
rect 9528 26931 9568 26963
rect 9600 26931 9640 26963
rect 9672 26931 9712 26963
rect 9744 26931 9784 26963
rect 9816 26931 9856 26963
rect 9888 26931 9928 26963
rect 9960 26931 10000 26963
rect 10032 26931 10072 26963
rect 10104 26931 10144 26963
rect 10176 26931 10216 26963
rect 10248 26931 10288 26963
rect 10320 26931 10360 26963
rect 10392 26931 10432 26963
rect 10464 26931 10504 26963
rect 10536 26931 10576 26963
rect 10608 26931 10648 26963
rect 10680 26931 10720 26963
rect 10752 26931 10792 26963
rect 10824 26931 10864 26963
rect 10896 26931 10936 26963
rect 10968 26931 11008 26963
rect 11040 26931 11080 26963
rect 11112 26931 11152 26963
rect 11184 26931 11224 26963
rect 11256 26931 11296 26963
rect 11328 26931 11368 26963
rect 11400 26931 11440 26963
rect 11472 26931 11512 26963
rect 11544 26931 11584 26963
rect 11616 26931 11656 26963
rect 11688 26931 11728 26963
rect 11760 26931 11800 26963
rect 11832 26931 11872 26963
rect 11904 26931 11944 26963
rect 11976 26931 12016 26963
rect 12048 26931 12088 26963
rect 12120 26931 12160 26963
rect 12192 26931 12232 26963
rect 12264 26931 12304 26963
rect 12336 26931 12376 26963
rect 12408 26931 12448 26963
rect 12480 26931 12520 26963
rect 12552 26931 12592 26963
rect 12624 26931 12664 26963
rect 12696 26931 12736 26963
rect 12768 26931 12808 26963
rect 12840 26931 12880 26963
rect 12912 26931 12952 26963
rect 12984 26931 13024 26963
rect 13056 26931 13096 26963
rect 13128 26931 13168 26963
rect 13200 26931 13240 26963
rect 13272 26931 13312 26963
rect 13344 26931 13384 26963
rect 13416 26931 13456 26963
rect 13488 26931 13528 26963
rect 13560 26931 13600 26963
rect 13632 26931 13672 26963
rect 13704 26931 13744 26963
rect 13776 26931 13816 26963
rect 13848 26931 13888 26963
rect 13920 26931 13960 26963
rect 13992 26931 14032 26963
rect 14064 26931 14104 26963
rect 14136 26931 14176 26963
rect 14208 26931 14248 26963
rect 14280 26931 14320 26963
rect 14352 26931 14392 26963
rect 14424 26931 14464 26963
rect 14496 26931 14536 26963
rect 14568 26931 14608 26963
rect 14640 26931 14680 26963
rect 14712 26931 14752 26963
rect 14784 26931 14824 26963
rect 14856 26931 14896 26963
rect 14928 26931 14968 26963
rect 15000 26931 15040 26963
rect 15072 26931 15112 26963
rect 15144 26931 15184 26963
rect 15216 26931 15256 26963
rect 15288 26931 15328 26963
rect 15360 26931 15400 26963
rect 15432 26931 15472 26963
rect 15504 26931 15544 26963
rect 15576 26931 15616 26963
rect 15648 26931 15688 26963
rect 15720 26931 15760 26963
rect 15792 26931 15832 26963
rect 15864 26931 15904 26963
rect 15936 26931 16000 26963
rect 0 26891 16000 26931
rect 0 26859 64 26891
rect 96 26859 136 26891
rect 168 26859 208 26891
rect 240 26859 280 26891
rect 312 26859 352 26891
rect 384 26859 424 26891
rect 456 26859 496 26891
rect 528 26859 568 26891
rect 600 26859 640 26891
rect 672 26859 712 26891
rect 744 26859 784 26891
rect 816 26859 856 26891
rect 888 26859 928 26891
rect 960 26859 1000 26891
rect 1032 26859 1072 26891
rect 1104 26859 1144 26891
rect 1176 26859 1216 26891
rect 1248 26859 1288 26891
rect 1320 26859 1360 26891
rect 1392 26859 1432 26891
rect 1464 26859 1504 26891
rect 1536 26859 1576 26891
rect 1608 26859 1648 26891
rect 1680 26859 1720 26891
rect 1752 26859 1792 26891
rect 1824 26859 1864 26891
rect 1896 26859 1936 26891
rect 1968 26859 2008 26891
rect 2040 26859 2080 26891
rect 2112 26859 2152 26891
rect 2184 26859 2224 26891
rect 2256 26859 2296 26891
rect 2328 26859 2368 26891
rect 2400 26859 2440 26891
rect 2472 26859 2512 26891
rect 2544 26859 2584 26891
rect 2616 26859 2656 26891
rect 2688 26859 2728 26891
rect 2760 26859 2800 26891
rect 2832 26859 2872 26891
rect 2904 26859 2944 26891
rect 2976 26859 3016 26891
rect 3048 26859 3088 26891
rect 3120 26859 3160 26891
rect 3192 26859 3232 26891
rect 3264 26859 3304 26891
rect 3336 26859 3376 26891
rect 3408 26859 3448 26891
rect 3480 26859 3520 26891
rect 3552 26859 3592 26891
rect 3624 26859 3664 26891
rect 3696 26859 3736 26891
rect 3768 26859 3808 26891
rect 3840 26859 3880 26891
rect 3912 26859 3952 26891
rect 3984 26859 4024 26891
rect 4056 26859 4096 26891
rect 4128 26859 4168 26891
rect 4200 26859 4240 26891
rect 4272 26859 4312 26891
rect 4344 26859 4384 26891
rect 4416 26859 4456 26891
rect 4488 26859 4528 26891
rect 4560 26859 4600 26891
rect 4632 26859 4672 26891
rect 4704 26859 4744 26891
rect 4776 26859 4816 26891
rect 4848 26859 4888 26891
rect 4920 26859 4960 26891
rect 4992 26859 5032 26891
rect 5064 26859 5104 26891
rect 5136 26859 5176 26891
rect 5208 26859 5248 26891
rect 5280 26859 5320 26891
rect 5352 26859 5392 26891
rect 5424 26859 5464 26891
rect 5496 26859 5536 26891
rect 5568 26859 5608 26891
rect 5640 26859 5680 26891
rect 5712 26859 5752 26891
rect 5784 26859 5824 26891
rect 5856 26859 5896 26891
rect 5928 26859 5968 26891
rect 6000 26859 6040 26891
rect 6072 26859 6112 26891
rect 6144 26859 6184 26891
rect 6216 26859 6256 26891
rect 6288 26859 6328 26891
rect 6360 26859 6400 26891
rect 6432 26859 6472 26891
rect 6504 26859 6544 26891
rect 6576 26859 6616 26891
rect 6648 26859 6688 26891
rect 6720 26859 6760 26891
rect 6792 26859 6832 26891
rect 6864 26859 6904 26891
rect 6936 26859 6976 26891
rect 7008 26859 7048 26891
rect 7080 26859 7120 26891
rect 7152 26859 7192 26891
rect 7224 26859 7264 26891
rect 7296 26859 7336 26891
rect 7368 26859 7408 26891
rect 7440 26859 7480 26891
rect 7512 26859 7552 26891
rect 7584 26859 7624 26891
rect 7656 26859 7696 26891
rect 7728 26859 7768 26891
rect 7800 26859 7840 26891
rect 7872 26859 7912 26891
rect 7944 26859 7984 26891
rect 8016 26859 8056 26891
rect 8088 26859 8128 26891
rect 8160 26859 8200 26891
rect 8232 26859 8272 26891
rect 8304 26859 8344 26891
rect 8376 26859 8416 26891
rect 8448 26859 8488 26891
rect 8520 26859 8560 26891
rect 8592 26859 8632 26891
rect 8664 26859 8704 26891
rect 8736 26859 8776 26891
rect 8808 26859 8848 26891
rect 8880 26859 8920 26891
rect 8952 26859 8992 26891
rect 9024 26859 9064 26891
rect 9096 26859 9136 26891
rect 9168 26859 9208 26891
rect 9240 26859 9280 26891
rect 9312 26859 9352 26891
rect 9384 26859 9424 26891
rect 9456 26859 9496 26891
rect 9528 26859 9568 26891
rect 9600 26859 9640 26891
rect 9672 26859 9712 26891
rect 9744 26859 9784 26891
rect 9816 26859 9856 26891
rect 9888 26859 9928 26891
rect 9960 26859 10000 26891
rect 10032 26859 10072 26891
rect 10104 26859 10144 26891
rect 10176 26859 10216 26891
rect 10248 26859 10288 26891
rect 10320 26859 10360 26891
rect 10392 26859 10432 26891
rect 10464 26859 10504 26891
rect 10536 26859 10576 26891
rect 10608 26859 10648 26891
rect 10680 26859 10720 26891
rect 10752 26859 10792 26891
rect 10824 26859 10864 26891
rect 10896 26859 10936 26891
rect 10968 26859 11008 26891
rect 11040 26859 11080 26891
rect 11112 26859 11152 26891
rect 11184 26859 11224 26891
rect 11256 26859 11296 26891
rect 11328 26859 11368 26891
rect 11400 26859 11440 26891
rect 11472 26859 11512 26891
rect 11544 26859 11584 26891
rect 11616 26859 11656 26891
rect 11688 26859 11728 26891
rect 11760 26859 11800 26891
rect 11832 26859 11872 26891
rect 11904 26859 11944 26891
rect 11976 26859 12016 26891
rect 12048 26859 12088 26891
rect 12120 26859 12160 26891
rect 12192 26859 12232 26891
rect 12264 26859 12304 26891
rect 12336 26859 12376 26891
rect 12408 26859 12448 26891
rect 12480 26859 12520 26891
rect 12552 26859 12592 26891
rect 12624 26859 12664 26891
rect 12696 26859 12736 26891
rect 12768 26859 12808 26891
rect 12840 26859 12880 26891
rect 12912 26859 12952 26891
rect 12984 26859 13024 26891
rect 13056 26859 13096 26891
rect 13128 26859 13168 26891
rect 13200 26859 13240 26891
rect 13272 26859 13312 26891
rect 13344 26859 13384 26891
rect 13416 26859 13456 26891
rect 13488 26859 13528 26891
rect 13560 26859 13600 26891
rect 13632 26859 13672 26891
rect 13704 26859 13744 26891
rect 13776 26859 13816 26891
rect 13848 26859 13888 26891
rect 13920 26859 13960 26891
rect 13992 26859 14032 26891
rect 14064 26859 14104 26891
rect 14136 26859 14176 26891
rect 14208 26859 14248 26891
rect 14280 26859 14320 26891
rect 14352 26859 14392 26891
rect 14424 26859 14464 26891
rect 14496 26859 14536 26891
rect 14568 26859 14608 26891
rect 14640 26859 14680 26891
rect 14712 26859 14752 26891
rect 14784 26859 14824 26891
rect 14856 26859 14896 26891
rect 14928 26859 14968 26891
rect 15000 26859 15040 26891
rect 15072 26859 15112 26891
rect 15144 26859 15184 26891
rect 15216 26859 15256 26891
rect 15288 26859 15328 26891
rect 15360 26859 15400 26891
rect 15432 26859 15472 26891
rect 15504 26859 15544 26891
rect 15576 26859 15616 26891
rect 15648 26859 15688 26891
rect 15720 26859 15760 26891
rect 15792 26859 15832 26891
rect 15864 26859 15904 26891
rect 15936 26859 16000 26891
rect 0 26819 16000 26859
rect 0 26787 64 26819
rect 96 26787 136 26819
rect 168 26787 208 26819
rect 240 26787 280 26819
rect 312 26787 352 26819
rect 384 26787 424 26819
rect 456 26787 496 26819
rect 528 26787 568 26819
rect 600 26787 640 26819
rect 672 26787 712 26819
rect 744 26787 784 26819
rect 816 26787 856 26819
rect 888 26787 928 26819
rect 960 26787 1000 26819
rect 1032 26787 1072 26819
rect 1104 26787 1144 26819
rect 1176 26787 1216 26819
rect 1248 26787 1288 26819
rect 1320 26787 1360 26819
rect 1392 26787 1432 26819
rect 1464 26787 1504 26819
rect 1536 26787 1576 26819
rect 1608 26787 1648 26819
rect 1680 26787 1720 26819
rect 1752 26787 1792 26819
rect 1824 26787 1864 26819
rect 1896 26787 1936 26819
rect 1968 26787 2008 26819
rect 2040 26787 2080 26819
rect 2112 26787 2152 26819
rect 2184 26787 2224 26819
rect 2256 26787 2296 26819
rect 2328 26787 2368 26819
rect 2400 26787 2440 26819
rect 2472 26787 2512 26819
rect 2544 26787 2584 26819
rect 2616 26787 2656 26819
rect 2688 26787 2728 26819
rect 2760 26787 2800 26819
rect 2832 26787 2872 26819
rect 2904 26787 2944 26819
rect 2976 26787 3016 26819
rect 3048 26787 3088 26819
rect 3120 26787 3160 26819
rect 3192 26787 3232 26819
rect 3264 26787 3304 26819
rect 3336 26787 3376 26819
rect 3408 26787 3448 26819
rect 3480 26787 3520 26819
rect 3552 26787 3592 26819
rect 3624 26787 3664 26819
rect 3696 26787 3736 26819
rect 3768 26787 3808 26819
rect 3840 26787 3880 26819
rect 3912 26787 3952 26819
rect 3984 26787 4024 26819
rect 4056 26787 4096 26819
rect 4128 26787 4168 26819
rect 4200 26787 4240 26819
rect 4272 26787 4312 26819
rect 4344 26787 4384 26819
rect 4416 26787 4456 26819
rect 4488 26787 4528 26819
rect 4560 26787 4600 26819
rect 4632 26787 4672 26819
rect 4704 26787 4744 26819
rect 4776 26787 4816 26819
rect 4848 26787 4888 26819
rect 4920 26787 4960 26819
rect 4992 26787 5032 26819
rect 5064 26787 5104 26819
rect 5136 26787 5176 26819
rect 5208 26787 5248 26819
rect 5280 26787 5320 26819
rect 5352 26787 5392 26819
rect 5424 26787 5464 26819
rect 5496 26787 5536 26819
rect 5568 26787 5608 26819
rect 5640 26787 5680 26819
rect 5712 26787 5752 26819
rect 5784 26787 5824 26819
rect 5856 26787 5896 26819
rect 5928 26787 5968 26819
rect 6000 26787 6040 26819
rect 6072 26787 6112 26819
rect 6144 26787 6184 26819
rect 6216 26787 6256 26819
rect 6288 26787 6328 26819
rect 6360 26787 6400 26819
rect 6432 26787 6472 26819
rect 6504 26787 6544 26819
rect 6576 26787 6616 26819
rect 6648 26787 6688 26819
rect 6720 26787 6760 26819
rect 6792 26787 6832 26819
rect 6864 26787 6904 26819
rect 6936 26787 6976 26819
rect 7008 26787 7048 26819
rect 7080 26787 7120 26819
rect 7152 26787 7192 26819
rect 7224 26787 7264 26819
rect 7296 26787 7336 26819
rect 7368 26787 7408 26819
rect 7440 26787 7480 26819
rect 7512 26787 7552 26819
rect 7584 26787 7624 26819
rect 7656 26787 7696 26819
rect 7728 26787 7768 26819
rect 7800 26787 7840 26819
rect 7872 26787 7912 26819
rect 7944 26787 7984 26819
rect 8016 26787 8056 26819
rect 8088 26787 8128 26819
rect 8160 26787 8200 26819
rect 8232 26787 8272 26819
rect 8304 26787 8344 26819
rect 8376 26787 8416 26819
rect 8448 26787 8488 26819
rect 8520 26787 8560 26819
rect 8592 26787 8632 26819
rect 8664 26787 8704 26819
rect 8736 26787 8776 26819
rect 8808 26787 8848 26819
rect 8880 26787 8920 26819
rect 8952 26787 8992 26819
rect 9024 26787 9064 26819
rect 9096 26787 9136 26819
rect 9168 26787 9208 26819
rect 9240 26787 9280 26819
rect 9312 26787 9352 26819
rect 9384 26787 9424 26819
rect 9456 26787 9496 26819
rect 9528 26787 9568 26819
rect 9600 26787 9640 26819
rect 9672 26787 9712 26819
rect 9744 26787 9784 26819
rect 9816 26787 9856 26819
rect 9888 26787 9928 26819
rect 9960 26787 10000 26819
rect 10032 26787 10072 26819
rect 10104 26787 10144 26819
rect 10176 26787 10216 26819
rect 10248 26787 10288 26819
rect 10320 26787 10360 26819
rect 10392 26787 10432 26819
rect 10464 26787 10504 26819
rect 10536 26787 10576 26819
rect 10608 26787 10648 26819
rect 10680 26787 10720 26819
rect 10752 26787 10792 26819
rect 10824 26787 10864 26819
rect 10896 26787 10936 26819
rect 10968 26787 11008 26819
rect 11040 26787 11080 26819
rect 11112 26787 11152 26819
rect 11184 26787 11224 26819
rect 11256 26787 11296 26819
rect 11328 26787 11368 26819
rect 11400 26787 11440 26819
rect 11472 26787 11512 26819
rect 11544 26787 11584 26819
rect 11616 26787 11656 26819
rect 11688 26787 11728 26819
rect 11760 26787 11800 26819
rect 11832 26787 11872 26819
rect 11904 26787 11944 26819
rect 11976 26787 12016 26819
rect 12048 26787 12088 26819
rect 12120 26787 12160 26819
rect 12192 26787 12232 26819
rect 12264 26787 12304 26819
rect 12336 26787 12376 26819
rect 12408 26787 12448 26819
rect 12480 26787 12520 26819
rect 12552 26787 12592 26819
rect 12624 26787 12664 26819
rect 12696 26787 12736 26819
rect 12768 26787 12808 26819
rect 12840 26787 12880 26819
rect 12912 26787 12952 26819
rect 12984 26787 13024 26819
rect 13056 26787 13096 26819
rect 13128 26787 13168 26819
rect 13200 26787 13240 26819
rect 13272 26787 13312 26819
rect 13344 26787 13384 26819
rect 13416 26787 13456 26819
rect 13488 26787 13528 26819
rect 13560 26787 13600 26819
rect 13632 26787 13672 26819
rect 13704 26787 13744 26819
rect 13776 26787 13816 26819
rect 13848 26787 13888 26819
rect 13920 26787 13960 26819
rect 13992 26787 14032 26819
rect 14064 26787 14104 26819
rect 14136 26787 14176 26819
rect 14208 26787 14248 26819
rect 14280 26787 14320 26819
rect 14352 26787 14392 26819
rect 14424 26787 14464 26819
rect 14496 26787 14536 26819
rect 14568 26787 14608 26819
rect 14640 26787 14680 26819
rect 14712 26787 14752 26819
rect 14784 26787 14824 26819
rect 14856 26787 14896 26819
rect 14928 26787 14968 26819
rect 15000 26787 15040 26819
rect 15072 26787 15112 26819
rect 15144 26787 15184 26819
rect 15216 26787 15256 26819
rect 15288 26787 15328 26819
rect 15360 26787 15400 26819
rect 15432 26787 15472 26819
rect 15504 26787 15544 26819
rect 15576 26787 15616 26819
rect 15648 26787 15688 26819
rect 15720 26787 15760 26819
rect 15792 26787 15832 26819
rect 15864 26787 15904 26819
rect 15936 26787 16000 26819
rect 0 26747 16000 26787
rect 0 26715 64 26747
rect 96 26715 136 26747
rect 168 26715 208 26747
rect 240 26715 280 26747
rect 312 26715 352 26747
rect 384 26715 424 26747
rect 456 26715 496 26747
rect 528 26715 568 26747
rect 600 26715 640 26747
rect 672 26715 712 26747
rect 744 26715 784 26747
rect 816 26715 856 26747
rect 888 26715 928 26747
rect 960 26715 1000 26747
rect 1032 26715 1072 26747
rect 1104 26715 1144 26747
rect 1176 26715 1216 26747
rect 1248 26715 1288 26747
rect 1320 26715 1360 26747
rect 1392 26715 1432 26747
rect 1464 26715 1504 26747
rect 1536 26715 1576 26747
rect 1608 26715 1648 26747
rect 1680 26715 1720 26747
rect 1752 26715 1792 26747
rect 1824 26715 1864 26747
rect 1896 26715 1936 26747
rect 1968 26715 2008 26747
rect 2040 26715 2080 26747
rect 2112 26715 2152 26747
rect 2184 26715 2224 26747
rect 2256 26715 2296 26747
rect 2328 26715 2368 26747
rect 2400 26715 2440 26747
rect 2472 26715 2512 26747
rect 2544 26715 2584 26747
rect 2616 26715 2656 26747
rect 2688 26715 2728 26747
rect 2760 26715 2800 26747
rect 2832 26715 2872 26747
rect 2904 26715 2944 26747
rect 2976 26715 3016 26747
rect 3048 26715 3088 26747
rect 3120 26715 3160 26747
rect 3192 26715 3232 26747
rect 3264 26715 3304 26747
rect 3336 26715 3376 26747
rect 3408 26715 3448 26747
rect 3480 26715 3520 26747
rect 3552 26715 3592 26747
rect 3624 26715 3664 26747
rect 3696 26715 3736 26747
rect 3768 26715 3808 26747
rect 3840 26715 3880 26747
rect 3912 26715 3952 26747
rect 3984 26715 4024 26747
rect 4056 26715 4096 26747
rect 4128 26715 4168 26747
rect 4200 26715 4240 26747
rect 4272 26715 4312 26747
rect 4344 26715 4384 26747
rect 4416 26715 4456 26747
rect 4488 26715 4528 26747
rect 4560 26715 4600 26747
rect 4632 26715 4672 26747
rect 4704 26715 4744 26747
rect 4776 26715 4816 26747
rect 4848 26715 4888 26747
rect 4920 26715 4960 26747
rect 4992 26715 5032 26747
rect 5064 26715 5104 26747
rect 5136 26715 5176 26747
rect 5208 26715 5248 26747
rect 5280 26715 5320 26747
rect 5352 26715 5392 26747
rect 5424 26715 5464 26747
rect 5496 26715 5536 26747
rect 5568 26715 5608 26747
rect 5640 26715 5680 26747
rect 5712 26715 5752 26747
rect 5784 26715 5824 26747
rect 5856 26715 5896 26747
rect 5928 26715 5968 26747
rect 6000 26715 6040 26747
rect 6072 26715 6112 26747
rect 6144 26715 6184 26747
rect 6216 26715 6256 26747
rect 6288 26715 6328 26747
rect 6360 26715 6400 26747
rect 6432 26715 6472 26747
rect 6504 26715 6544 26747
rect 6576 26715 6616 26747
rect 6648 26715 6688 26747
rect 6720 26715 6760 26747
rect 6792 26715 6832 26747
rect 6864 26715 6904 26747
rect 6936 26715 6976 26747
rect 7008 26715 7048 26747
rect 7080 26715 7120 26747
rect 7152 26715 7192 26747
rect 7224 26715 7264 26747
rect 7296 26715 7336 26747
rect 7368 26715 7408 26747
rect 7440 26715 7480 26747
rect 7512 26715 7552 26747
rect 7584 26715 7624 26747
rect 7656 26715 7696 26747
rect 7728 26715 7768 26747
rect 7800 26715 7840 26747
rect 7872 26715 7912 26747
rect 7944 26715 7984 26747
rect 8016 26715 8056 26747
rect 8088 26715 8128 26747
rect 8160 26715 8200 26747
rect 8232 26715 8272 26747
rect 8304 26715 8344 26747
rect 8376 26715 8416 26747
rect 8448 26715 8488 26747
rect 8520 26715 8560 26747
rect 8592 26715 8632 26747
rect 8664 26715 8704 26747
rect 8736 26715 8776 26747
rect 8808 26715 8848 26747
rect 8880 26715 8920 26747
rect 8952 26715 8992 26747
rect 9024 26715 9064 26747
rect 9096 26715 9136 26747
rect 9168 26715 9208 26747
rect 9240 26715 9280 26747
rect 9312 26715 9352 26747
rect 9384 26715 9424 26747
rect 9456 26715 9496 26747
rect 9528 26715 9568 26747
rect 9600 26715 9640 26747
rect 9672 26715 9712 26747
rect 9744 26715 9784 26747
rect 9816 26715 9856 26747
rect 9888 26715 9928 26747
rect 9960 26715 10000 26747
rect 10032 26715 10072 26747
rect 10104 26715 10144 26747
rect 10176 26715 10216 26747
rect 10248 26715 10288 26747
rect 10320 26715 10360 26747
rect 10392 26715 10432 26747
rect 10464 26715 10504 26747
rect 10536 26715 10576 26747
rect 10608 26715 10648 26747
rect 10680 26715 10720 26747
rect 10752 26715 10792 26747
rect 10824 26715 10864 26747
rect 10896 26715 10936 26747
rect 10968 26715 11008 26747
rect 11040 26715 11080 26747
rect 11112 26715 11152 26747
rect 11184 26715 11224 26747
rect 11256 26715 11296 26747
rect 11328 26715 11368 26747
rect 11400 26715 11440 26747
rect 11472 26715 11512 26747
rect 11544 26715 11584 26747
rect 11616 26715 11656 26747
rect 11688 26715 11728 26747
rect 11760 26715 11800 26747
rect 11832 26715 11872 26747
rect 11904 26715 11944 26747
rect 11976 26715 12016 26747
rect 12048 26715 12088 26747
rect 12120 26715 12160 26747
rect 12192 26715 12232 26747
rect 12264 26715 12304 26747
rect 12336 26715 12376 26747
rect 12408 26715 12448 26747
rect 12480 26715 12520 26747
rect 12552 26715 12592 26747
rect 12624 26715 12664 26747
rect 12696 26715 12736 26747
rect 12768 26715 12808 26747
rect 12840 26715 12880 26747
rect 12912 26715 12952 26747
rect 12984 26715 13024 26747
rect 13056 26715 13096 26747
rect 13128 26715 13168 26747
rect 13200 26715 13240 26747
rect 13272 26715 13312 26747
rect 13344 26715 13384 26747
rect 13416 26715 13456 26747
rect 13488 26715 13528 26747
rect 13560 26715 13600 26747
rect 13632 26715 13672 26747
rect 13704 26715 13744 26747
rect 13776 26715 13816 26747
rect 13848 26715 13888 26747
rect 13920 26715 13960 26747
rect 13992 26715 14032 26747
rect 14064 26715 14104 26747
rect 14136 26715 14176 26747
rect 14208 26715 14248 26747
rect 14280 26715 14320 26747
rect 14352 26715 14392 26747
rect 14424 26715 14464 26747
rect 14496 26715 14536 26747
rect 14568 26715 14608 26747
rect 14640 26715 14680 26747
rect 14712 26715 14752 26747
rect 14784 26715 14824 26747
rect 14856 26715 14896 26747
rect 14928 26715 14968 26747
rect 15000 26715 15040 26747
rect 15072 26715 15112 26747
rect 15144 26715 15184 26747
rect 15216 26715 15256 26747
rect 15288 26715 15328 26747
rect 15360 26715 15400 26747
rect 15432 26715 15472 26747
rect 15504 26715 15544 26747
rect 15576 26715 15616 26747
rect 15648 26715 15688 26747
rect 15720 26715 15760 26747
rect 15792 26715 15832 26747
rect 15864 26715 15904 26747
rect 15936 26715 16000 26747
rect 0 26675 16000 26715
rect 0 26643 64 26675
rect 96 26643 136 26675
rect 168 26643 208 26675
rect 240 26643 280 26675
rect 312 26643 352 26675
rect 384 26643 424 26675
rect 456 26643 496 26675
rect 528 26643 568 26675
rect 600 26643 640 26675
rect 672 26643 712 26675
rect 744 26643 784 26675
rect 816 26643 856 26675
rect 888 26643 928 26675
rect 960 26643 1000 26675
rect 1032 26643 1072 26675
rect 1104 26643 1144 26675
rect 1176 26643 1216 26675
rect 1248 26643 1288 26675
rect 1320 26643 1360 26675
rect 1392 26643 1432 26675
rect 1464 26643 1504 26675
rect 1536 26643 1576 26675
rect 1608 26643 1648 26675
rect 1680 26643 1720 26675
rect 1752 26643 1792 26675
rect 1824 26643 1864 26675
rect 1896 26643 1936 26675
rect 1968 26643 2008 26675
rect 2040 26643 2080 26675
rect 2112 26643 2152 26675
rect 2184 26643 2224 26675
rect 2256 26643 2296 26675
rect 2328 26643 2368 26675
rect 2400 26643 2440 26675
rect 2472 26643 2512 26675
rect 2544 26643 2584 26675
rect 2616 26643 2656 26675
rect 2688 26643 2728 26675
rect 2760 26643 2800 26675
rect 2832 26643 2872 26675
rect 2904 26643 2944 26675
rect 2976 26643 3016 26675
rect 3048 26643 3088 26675
rect 3120 26643 3160 26675
rect 3192 26643 3232 26675
rect 3264 26643 3304 26675
rect 3336 26643 3376 26675
rect 3408 26643 3448 26675
rect 3480 26643 3520 26675
rect 3552 26643 3592 26675
rect 3624 26643 3664 26675
rect 3696 26643 3736 26675
rect 3768 26643 3808 26675
rect 3840 26643 3880 26675
rect 3912 26643 3952 26675
rect 3984 26643 4024 26675
rect 4056 26643 4096 26675
rect 4128 26643 4168 26675
rect 4200 26643 4240 26675
rect 4272 26643 4312 26675
rect 4344 26643 4384 26675
rect 4416 26643 4456 26675
rect 4488 26643 4528 26675
rect 4560 26643 4600 26675
rect 4632 26643 4672 26675
rect 4704 26643 4744 26675
rect 4776 26643 4816 26675
rect 4848 26643 4888 26675
rect 4920 26643 4960 26675
rect 4992 26643 5032 26675
rect 5064 26643 5104 26675
rect 5136 26643 5176 26675
rect 5208 26643 5248 26675
rect 5280 26643 5320 26675
rect 5352 26643 5392 26675
rect 5424 26643 5464 26675
rect 5496 26643 5536 26675
rect 5568 26643 5608 26675
rect 5640 26643 5680 26675
rect 5712 26643 5752 26675
rect 5784 26643 5824 26675
rect 5856 26643 5896 26675
rect 5928 26643 5968 26675
rect 6000 26643 6040 26675
rect 6072 26643 6112 26675
rect 6144 26643 6184 26675
rect 6216 26643 6256 26675
rect 6288 26643 6328 26675
rect 6360 26643 6400 26675
rect 6432 26643 6472 26675
rect 6504 26643 6544 26675
rect 6576 26643 6616 26675
rect 6648 26643 6688 26675
rect 6720 26643 6760 26675
rect 6792 26643 6832 26675
rect 6864 26643 6904 26675
rect 6936 26643 6976 26675
rect 7008 26643 7048 26675
rect 7080 26643 7120 26675
rect 7152 26643 7192 26675
rect 7224 26643 7264 26675
rect 7296 26643 7336 26675
rect 7368 26643 7408 26675
rect 7440 26643 7480 26675
rect 7512 26643 7552 26675
rect 7584 26643 7624 26675
rect 7656 26643 7696 26675
rect 7728 26643 7768 26675
rect 7800 26643 7840 26675
rect 7872 26643 7912 26675
rect 7944 26643 7984 26675
rect 8016 26643 8056 26675
rect 8088 26643 8128 26675
rect 8160 26643 8200 26675
rect 8232 26643 8272 26675
rect 8304 26643 8344 26675
rect 8376 26643 8416 26675
rect 8448 26643 8488 26675
rect 8520 26643 8560 26675
rect 8592 26643 8632 26675
rect 8664 26643 8704 26675
rect 8736 26643 8776 26675
rect 8808 26643 8848 26675
rect 8880 26643 8920 26675
rect 8952 26643 8992 26675
rect 9024 26643 9064 26675
rect 9096 26643 9136 26675
rect 9168 26643 9208 26675
rect 9240 26643 9280 26675
rect 9312 26643 9352 26675
rect 9384 26643 9424 26675
rect 9456 26643 9496 26675
rect 9528 26643 9568 26675
rect 9600 26643 9640 26675
rect 9672 26643 9712 26675
rect 9744 26643 9784 26675
rect 9816 26643 9856 26675
rect 9888 26643 9928 26675
rect 9960 26643 10000 26675
rect 10032 26643 10072 26675
rect 10104 26643 10144 26675
rect 10176 26643 10216 26675
rect 10248 26643 10288 26675
rect 10320 26643 10360 26675
rect 10392 26643 10432 26675
rect 10464 26643 10504 26675
rect 10536 26643 10576 26675
rect 10608 26643 10648 26675
rect 10680 26643 10720 26675
rect 10752 26643 10792 26675
rect 10824 26643 10864 26675
rect 10896 26643 10936 26675
rect 10968 26643 11008 26675
rect 11040 26643 11080 26675
rect 11112 26643 11152 26675
rect 11184 26643 11224 26675
rect 11256 26643 11296 26675
rect 11328 26643 11368 26675
rect 11400 26643 11440 26675
rect 11472 26643 11512 26675
rect 11544 26643 11584 26675
rect 11616 26643 11656 26675
rect 11688 26643 11728 26675
rect 11760 26643 11800 26675
rect 11832 26643 11872 26675
rect 11904 26643 11944 26675
rect 11976 26643 12016 26675
rect 12048 26643 12088 26675
rect 12120 26643 12160 26675
rect 12192 26643 12232 26675
rect 12264 26643 12304 26675
rect 12336 26643 12376 26675
rect 12408 26643 12448 26675
rect 12480 26643 12520 26675
rect 12552 26643 12592 26675
rect 12624 26643 12664 26675
rect 12696 26643 12736 26675
rect 12768 26643 12808 26675
rect 12840 26643 12880 26675
rect 12912 26643 12952 26675
rect 12984 26643 13024 26675
rect 13056 26643 13096 26675
rect 13128 26643 13168 26675
rect 13200 26643 13240 26675
rect 13272 26643 13312 26675
rect 13344 26643 13384 26675
rect 13416 26643 13456 26675
rect 13488 26643 13528 26675
rect 13560 26643 13600 26675
rect 13632 26643 13672 26675
rect 13704 26643 13744 26675
rect 13776 26643 13816 26675
rect 13848 26643 13888 26675
rect 13920 26643 13960 26675
rect 13992 26643 14032 26675
rect 14064 26643 14104 26675
rect 14136 26643 14176 26675
rect 14208 26643 14248 26675
rect 14280 26643 14320 26675
rect 14352 26643 14392 26675
rect 14424 26643 14464 26675
rect 14496 26643 14536 26675
rect 14568 26643 14608 26675
rect 14640 26643 14680 26675
rect 14712 26643 14752 26675
rect 14784 26643 14824 26675
rect 14856 26643 14896 26675
rect 14928 26643 14968 26675
rect 15000 26643 15040 26675
rect 15072 26643 15112 26675
rect 15144 26643 15184 26675
rect 15216 26643 15256 26675
rect 15288 26643 15328 26675
rect 15360 26643 15400 26675
rect 15432 26643 15472 26675
rect 15504 26643 15544 26675
rect 15576 26643 15616 26675
rect 15648 26643 15688 26675
rect 15720 26643 15760 26675
rect 15792 26643 15832 26675
rect 15864 26643 15904 26675
rect 15936 26643 16000 26675
rect 0 26603 16000 26643
rect 0 26571 64 26603
rect 96 26571 136 26603
rect 168 26571 208 26603
rect 240 26571 280 26603
rect 312 26571 352 26603
rect 384 26571 424 26603
rect 456 26571 496 26603
rect 528 26571 568 26603
rect 600 26571 640 26603
rect 672 26571 712 26603
rect 744 26571 784 26603
rect 816 26571 856 26603
rect 888 26571 928 26603
rect 960 26571 1000 26603
rect 1032 26571 1072 26603
rect 1104 26571 1144 26603
rect 1176 26571 1216 26603
rect 1248 26571 1288 26603
rect 1320 26571 1360 26603
rect 1392 26571 1432 26603
rect 1464 26571 1504 26603
rect 1536 26571 1576 26603
rect 1608 26571 1648 26603
rect 1680 26571 1720 26603
rect 1752 26571 1792 26603
rect 1824 26571 1864 26603
rect 1896 26571 1936 26603
rect 1968 26571 2008 26603
rect 2040 26571 2080 26603
rect 2112 26571 2152 26603
rect 2184 26571 2224 26603
rect 2256 26571 2296 26603
rect 2328 26571 2368 26603
rect 2400 26571 2440 26603
rect 2472 26571 2512 26603
rect 2544 26571 2584 26603
rect 2616 26571 2656 26603
rect 2688 26571 2728 26603
rect 2760 26571 2800 26603
rect 2832 26571 2872 26603
rect 2904 26571 2944 26603
rect 2976 26571 3016 26603
rect 3048 26571 3088 26603
rect 3120 26571 3160 26603
rect 3192 26571 3232 26603
rect 3264 26571 3304 26603
rect 3336 26571 3376 26603
rect 3408 26571 3448 26603
rect 3480 26571 3520 26603
rect 3552 26571 3592 26603
rect 3624 26571 3664 26603
rect 3696 26571 3736 26603
rect 3768 26571 3808 26603
rect 3840 26571 3880 26603
rect 3912 26571 3952 26603
rect 3984 26571 4024 26603
rect 4056 26571 4096 26603
rect 4128 26571 4168 26603
rect 4200 26571 4240 26603
rect 4272 26571 4312 26603
rect 4344 26571 4384 26603
rect 4416 26571 4456 26603
rect 4488 26571 4528 26603
rect 4560 26571 4600 26603
rect 4632 26571 4672 26603
rect 4704 26571 4744 26603
rect 4776 26571 4816 26603
rect 4848 26571 4888 26603
rect 4920 26571 4960 26603
rect 4992 26571 5032 26603
rect 5064 26571 5104 26603
rect 5136 26571 5176 26603
rect 5208 26571 5248 26603
rect 5280 26571 5320 26603
rect 5352 26571 5392 26603
rect 5424 26571 5464 26603
rect 5496 26571 5536 26603
rect 5568 26571 5608 26603
rect 5640 26571 5680 26603
rect 5712 26571 5752 26603
rect 5784 26571 5824 26603
rect 5856 26571 5896 26603
rect 5928 26571 5968 26603
rect 6000 26571 6040 26603
rect 6072 26571 6112 26603
rect 6144 26571 6184 26603
rect 6216 26571 6256 26603
rect 6288 26571 6328 26603
rect 6360 26571 6400 26603
rect 6432 26571 6472 26603
rect 6504 26571 6544 26603
rect 6576 26571 6616 26603
rect 6648 26571 6688 26603
rect 6720 26571 6760 26603
rect 6792 26571 6832 26603
rect 6864 26571 6904 26603
rect 6936 26571 6976 26603
rect 7008 26571 7048 26603
rect 7080 26571 7120 26603
rect 7152 26571 7192 26603
rect 7224 26571 7264 26603
rect 7296 26571 7336 26603
rect 7368 26571 7408 26603
rect 7440 26571 7480 26603
rect 7512 26571 7552 26603
rect 7584 26571 7624 26603
rect 7656 26571 7696 26603
rect 7728 26571 7768 26603
rect 7800 26571 7840 26603
rect 7872 26571 7912 26603
rect 7944 26571 7984 26603
rect 8016 26571 8056 26603
rect 8088 26571 8128 26603
rect 8160 26571 8200 26603
rect 8232 26571 8272 26603
rect 8304 26571 8344 26603
rect 8376 26571 8416 26603
rect 8448 26571 8488 26603
rect 8520 26571 8560 26603
rect 8592 26571 8632 26603
rect 8664 26571 8704 26603
rect 8736 26571 8776 26603
rect 8808 26571 8848 26603
rect 8880 26571 8920 26603
rect 8952 26571 8992 26603
rect 9024 26571 9064 26603
rect 9096 26571 9136 26603
rect 9168 26571 9208 26603
rect 9240 26571 9280 26603
rect 9312 26571 9352 26603
rect 9384 26571 9424 26603
rect 9456 26571 9496 26603
rect 9528 26571 9568 26603
rect 9600 26571 9640 26603
rect 9672 26571 9712 26603
rect 9744 26571 9784 26603
rect 9816 26571 9856 26603
rect 9888 26571 9928 26603
rect 9960 26571 10000 26603
rect 10032 26571 10072 26603
rect 10104 26571 10144 26603
rect 10176 26571 10216 26603
rect 10248 26571 10288 26603
rect 10320 26571 10360 26603
rect 10392 26571 10432 26603
rect 10464 26571 10504 26603
rect 10536 26571 10576 26603
rect 10608 26571 10648 26603
rect 10680 26571 10720 26603
rect 10752 26571 10792 26603
rect 10824 26571 10864 26603
rect 10896 26571 10936 26603
rect 10968 26571 11008 26603
rect 11040 26571 11080 26603
rect 11112 26571 11152 26603
rect 11184 26571 11224 26603
rect 11256 26571 11296 26603
rect 11328 26571 11368 26603
rect 11400 26571 11440 26603
rect 11472 26571 11512 26603
rect 11544 26571 11584 26603
rect 11616 26571 11656 26603
rect 11688 26571 11728 26603
rect 11760 26571 11800 26603
rect 11832 26571 11872 26603
rect 11904 26571 11944 26603
rect 11976 26571 12016 26603
rect 12048 26571 12088 26603
rect 12120 26571 12160 26603
rect 12192 26571 12232 26603
rect 12264 26571 12304 26603
rect 12336 26571 12376 26603
rect 12408 26571 12448 26603
rect 12480 26571 12520 26603
rect 12552 26571 12592 26603
rect 12624 26571 12664 26603
rect 12696 26571 12736 26603
rect 12768 26571 12808 26603
rect 12840 26571 12880 26603
rect 12912 26571 12952 26603
rect 12984 26571 13024 26603
rect 13056 26571 13096 26603
rect 13128 26571 13168 26603
rect 13200 26571 13240 26603
rect 13272 26571 13312 26603
rect 13344 26571 13384 26603
rect 13416 26571 13456 26603
rect 13488 26571 13528 26603
rect 13560 26571 13600 26603
rect 13632 26571 13672 26603
rect 13704 26571 13744 26603
rect 13776 26571 13816 26603
rect 13848 26571 13888 26603
rect 13920 26571 13960 26603
rect 13992 26571 14032 26603
rect 14064 26571 14104 26603
rect 14136 26571 14176 26603
rect 14208 26571 14248 26603
rect 14280 26571 14320 26603
rect 14352 26571 14392 26603
rect 14424 26571 14464 26603
rect 14496 26571 14536 26603
rect 14568 26571 14608 26603
rect 14640 26571 14680 26603
rect 14712 26571 14752 26603
rect 14784 26571 14824 26603
rect 14856 26571 14896 26603
rect 14928 26571 14968 26603
rect 15000 26571 15040 26603
rect 15072 26571 15112 26603
rect 15144 26571 15184 26603
rect 15216 26571 15256 26603
rect 15288 26571 15328 26603
rect 15360 26571 15400 26603
rect 15432 26571 15472 26603
rect 15504 26571 15544 26603
rect 15576 26571 15616 26603
rect 15648 26571 15688 26603
rect 15720 26571 15760 26603
rect 15792 26571 15832 26603
rect 15864 26571 15904 26603
rect 15936 26571 16000 26603
rect 0 26531 16000 26571
rect 0 26499 64 26531
rect 96 26499 136 26531
rect 168 26499 208 26531
rect 240 26499 280 26531
rect 312 26499 352 26531
rect 384 26499 424 26531
rect 456 26499 496 26531
rect 528 26499 568 26531
rect 600 26499 640 26531
rect 672 26499 712 26531
rect 744 26499 784 26531
rect 816 26499 856 26531
rect 888 26499 928 26531
rect 960 26499 1000 26531
rect 1032 26499 1072 26531
rect 1104 26499 1144 26531
rect 1176 26499 1216 26531
rect 1248 26499 1288 26531
rect 1320 26499 1360 26531
rect 1392 26499 1432 26531
rect 1464 26499 1504 26531
rect 1536 26499 1576 26531
rect 1608 26499 1648 26531
rect 1680 26499 1720 26531
rect 1752 26499 1792 26531
rect 1824 26499 1864 26531
rect 1896 26499 1936 26531
rect 1968 26499 2008 26531
rect 2040 26499 2080 26531
rect 2112 26499 2152 26531
rect 2184 26499 2224 26531
rect 2256 26499 2296 26531
rect 2328 26499 2368 26531
rect 2400 26499 2440 26531
rect 2472 26499 2512 26531
rect 2544 26499 2584 26531
rect 2616 26499 2656 26531
rect 2688 26499 2728 26531
rect 2760 26499 2800 26531
rect 2832 26499 2872 26531
rect 2904 26499 2944 26531
rect 2976 26499 3016 26531
rect 3048 26499 3088 26531
rect 3120 26499 3160 26531
rect 3192 26499 3232 26531
rect 3264 26499 3304 26531
rect 3336 26499 3376 26531
rect 3408 26499 3448 26531
rect 3480 26499 3520 26531
rect 3552 26499 3592 26531
rect 3624 26499 3664 26531
rect 3696 26499 3736 26531
rect 3768 26499 3808 26531
rect 3840 26499 3880 26531
rect 3912 26499 3952 26531
rect 3984 26499 4024 26531
rect 4056 26499 4096 26531
rect 4128 26499 4168 26531
rect 4200 26499 4240 26531
rect 4272 26499 4312 26531
rect 4344 26499 4384 26531
rect 4416 26499 4456 26531
rect 4488 26499 4528 26531
rect 4560 26499 4600 26531
rect 4632 26499 4672 26531
rect 4704 26499 4744 26531
rect 4776 26499 4816 26531
rect 4848 26499 4888 26531
rect 4920 26499 4960 26531
rect 4992 26499 5032 26531
rect 5064 26499 5104 26531
rect 5136 26499 5176 26531
rect 5208 26499 5248 26531
rect 5280 26499 5320 26531
rect 5352 26499 5392 26531
rect 5424 26499 5464 26531
rect 5496 26499 5536 26531
rect 5568 26499 5608 26531
rect 5640 26499 5680 26531
rect 5712 26499 5752 26531
rect 5784 26499 5824 26531
rect 5856 26499 5896 26531
rect 5928 26499 5968 26531
rect 6000 26499 6040 26531
rect 6072 26499 6112 26531
rect 6144 26499 6184 26531
rect 6216 26499 6256 26531
rect 6288 26499 6328 26531
rect 6360 26499 6400 26531
rect 6432 26499 6472 26531
rect 6504 26499 6544 26531
rect 6576 26499 6616 26531
rect 6648 26499 6688 26531
rect 6720 26499 6760 26531
rect 6792 26499 6832 26531
rect 6864 26499 6904 26531
rect 6936 26499 6976 26531
rect 7008 26499 7048 26531
rect 7080 26499 7120 26531
rect 7152 26499 7192 26531
rect 7224 26499 7264 26531
rect 7296 26499 7336 26531
rect 7368 26499 7408 26531
rect 7440 26499 7480 26531
rect 7512 26499 7552 26531
rect 7584 26499 7624 26531
rect 7656 26499 7696 26531
rect 7728 26499 7768 26531
rect 7800 26499 7840 26531
rect 7872 26499 7912 26531
rect 7944 26499 7984 26531
rect 8016 26499 8056 26531
rect 8088 26499 8128 26531
rect 8160 26499 8200 26531
rect 8232 26499 8272 26531
rect 8304 26499 8344 26531
rect 8376 26499 8416 26531
rect 8448 26499 8488 26531
rect 8520 26499 8560 26531
rect 8592 26499 8632 26531
rect 8664 26499 8704 26531
rect 8736 26499 8776 26531
rect 8808 26499 8848 26531
rect 8880 26499 8920 26531
rect 8952 26499 8992 26531
rect 9024 26499 9064 26531
rect 9096 26499 9136 26531
rect 9168 26499 9208 26531
rect 9240 26499 9280 26531
rect 9312 26499 9352 26531
rect 9384 26499 9424 26531
rect 9456 26499 9496 26531
rect 9528 26499 9568 26531
rect 9600 26499 9640 26531
rect 9672 26499 9712 26531
rect 9744 26499 9784 26531
rect 9816 26499 9856 26531
rect 9888 26499 9928 26531
rect 9960 26499 10000 26531
rect 10032 26499 10072 26531
rect 10104 26499 10144 26531
rect 10176 26499 10216 26531
rect 10248 26499 10288 26531
rect 10320 26499 10360 26531
rect 10392 26499 10432 26531
rect 10464 26499 10504 26531
rect 10536 26499 10576 26531
rect 10608 26499 10648 26531
rect 10680 26499 10720 26531
rect 10752 26499 10792 26531
rect 10824 26499 10864 26531
rect 10896 26499 10936 26531
rect 10968 26499 11008 26531
rect 11040 26499 11080 26531
rect 11112 26499 11152 26531
rect 11184 26499 11224 26531
rect 11256 26499 11296 26531
rect 11328 26499 11368 26531
rect 11400 26499 11440 26531
rect 11472 26499 11512 26531
rect 11544 26499 11584 26531
rect 11616 26499 11656 26531
rect 11688 26499 11728 26531
rect 11760 26499 11800 26531
rect 11832 26499 11872 26531
rect 11904 26499 11944 26531
rect 11976 26499 12016 26531
rect 12048 26499 12088 26531
rect 12120 26499 12160 26531
rect 12192 26499 12232 26531
rect 12264 26499 12304 26531
rect 12336 26499 12376 26531
rect 12408 26499 12448 26531
rect 12480 26499 12520 26531
rect 12552 26499 12592 26531
rect 12624 26499 12664 26531
rect 12696 26499 12736 26531
rect 12768 26499 12808 26531
rect 12840 26499 12880 26531
rect 12912 26499 12952 26531
rect 12984 26499 13024 26531
rect 13056 26499 13096 26531
rect 13128 26499 13168 26531
rect 13200 26499 13240 26531
rect 13272 26499 13312 26531
rect 13344 26499 13384 26531
rect 13416 26499 13456 26531
rect 13488 26499 13528 26531
rect 13560 26499 13600 26531
rect 13632 26499 13672 26531
rect 13704 26499 13744 26531
rect 13776 26499 13816 26531
rect 13848 26499 13888 26531
rect 13920 26499 13960 26531
rect 13992 26499 14032 26531
rect 14064 26499 14104 26531
rect 14136 26499 14176 26531
rect 14208 26499 14248 26531
rect 14280 26499 14320 26531
rect 14352 26499 14392 26531
rect 14424 26499 14464 26531
rect 14496 26499 14536 26531
rect 14568 26499 14608 26531
rect 14640 26499 14680 26531
rect 14712 26499 14752 26531
rect 14784 26499 14824 26531
rect 14856 26499 14896 26531
rect 14928 26499 14968 26531
rect 15000 26499 15040 26531
rect 15072 26499 15112 26531
rect 15144 26499 15184 26531
rect 15216 26499 15256 26531
rect 15288 26499 15328 26531
rect 15360 26499 15400 26531
rect 15432 26499 15472 26531
rect 15504 26499 15544 26531
rect 15576 26499 15616 26531
rect 15648 26499 15688 26531
rect 15720 26499 15760 26531
rect 15792 26499 15832 26531
rect 15864 26499 15904 26531
rect 15936 26499 16000 26531
rect 0 26459 16000 26499
rect 0 26427 64 26459
rect 96 26427 136 26459
rect 168 26427 208 26459
rect 240 26427 280 26459
rect 312 26427 352 26459
rect 384 26427 424 26459
rect 456 26427 496 26459
rect 528 26427 568 26459
rect 600 26427 640 26459
rect 672 26427 712 26459
rect 744 26427 784 26459
rect 816 26427 856 26459
rect 888 26427 928 26459
rect 960 26427 1000 26459
rect 1032 26427 1072 26459
rect 1104 26427 1144 26459
rect 1176 26427 1216 26459
rect 1248 26427 1288 26459
rect 1320 26427 1360 26459
rect 1392 26427 1432 26459
rect 1464 26427 1504 26459
rect 1536 26427 1576 26459
rect 1608 26427 1648 26459
rect 1680 26427 1720 26459
rect 1752 26427 1792 26459
rect 1824 26427 1864 26459
rect 1896 26427 1936 26459
rect 1968 26427 2008 26459
rect 2040 26427 2080 26459
rect 2112 26427 2152 26459
rect 2184 26427 2224 26459
rect 2256 26427 2296 26459
rect 2328 26427 2368 26459
rect 2400 26427 2440 26459
rect 2472 26427 2512 26459
rect 2544 26427 2584 26459
rect 2616 26427 2656 26459
rect 2688 26427 2728 26459
rect 2760 26427 2800 26459
rect 2832 26427 2872 26459
rect 2904 26427 2944 26459
rect 2976 26427 3016 26459
rect 3048 26427 3088 26459
rect 3120 26427 3160 26459
rect 3192 26427 3232 26459
rect 3264 26427 3304 26459
rect 3336 26427 3376 26459
rect 3408 26427 3448 26459
rect 3480 26427 3520 26459
rect 3552 26427 3592 26459
rect 3624 26427 3664 26459
rect 3696 26427 3736 26459
rect 3768 26427 3808 26459
rect 3840 26427 3880 26459
rect 3912 26427 3952 26459
rect 3984 26427 4024 26459
rect 4056 26427 4096 26459
rect 4128 26427 4168 26459
rect 4200 26427 4240 26459
rect 4272 26427 4312 26459
rect 4344 26427 4384 26459
rect 4416 26427 4456 26459
rect 4488 26427 4528 26459
rect 4560 26427 4600 26459
rect 4632 26427 4672 26459
rect 4704 26427 4744 26459
rect 4776 26427 4816 26459
rect 4848 26427 4888 26459
rect 4920 26427 4960 26459
rect 4992 26427 5032 26459
rect 5064 26427 5104 26459
rect 5136 26427 5176 26459
rect 5208 26427 5248 26459
rect 5280 26427 5320 26459
rect 5352 26427 5392 26459
rect 5424 26427 5464 26459
rect 5496 26427 5536 26459
rect 5568 26427 5608 26459
rect 5640 26427 5680 26459
rect 5712 26427 5752 26459
rect 5784 26427 5824 26459
rect 5856 26427 5896 26459
rect 5928 26427 5968 26459
rect 6000 26427 6040 26459
rect 6072 26427 6112 26459
rect 6144 26427 6184 26459
rect 6216 26427 6256 26459
rect 6288 26427 6328 26459
rect 6360 26427 6400 26459
rect 6432 26427 6472 26459
rect 6504 26427 6544 26459
rect 6576 26427 6616 26459
rect 6648 26427 6688 26459
rect 6720 26427 6760 26459
rect 6792 26427 6832 26459
rect 6864 26427 6904 26459
rect 6936 26427 6976 26459
rect 7008 26427 7048 26459
rect 7080 26427 7120 26459
rect 7152 26427 7192 26459
rect 7224 26427 7264 26459
rect 7296 26427 7336 26459
rect 7368 26427 7408 26459
rect 7440 26427 7480 26459
rect 7512 26427 7552 26459
rect 7584 26427 7624 26459
rect 7656 26427 7696 26459
rect 7728 26427 7768 26459
rect 7800 26427 7840 26459
rect 7872 26427 7912 26459
rect 7944 26427 7984 26459
rect 8016 26427 8056 26459
rect 8088 26427 8128 26459
rect 8160 26427 8200 26459
rect 8232 26427 8272 26459
rect 8304 26427 8344 26459
rect 8376 26427 8416 26459
rect 8448 26427 8488 26459
rect 8520 26427 8560 26459
rect 8592 26427 8632 26459
rect 8664 26427 8704 26459
rect 8736 26427 8776 26459
rect 8808 26427 8848 26459
rect 8880 26427 8920 26459
rect 8952 26427 8992 26459
rect 9024 26427 9064 26459
rect 9096 26427 9136 26459
rect 9168 26427 9208 26459
rect 9240 26427 9280 26459
rect 9312 26427 9352 26459
rect 9384 26427 9424 26459
rect 9456 26427 9496 26459
rect 9528 26427 9568 26459
rect 9600 26427 9640 26459
rect 9672 26427 9712 26459
rect 9744 26427 9784 26459
rect 9816 26427 9856 26459
rect 9888 26427 9928 26459
rect 9960 26427 10000 26459
rect 10032 26427 10072 26459
rect 10104 26427 10144 26459
rect 10176 26427 10216 26459
rect 10248 26427 10288 26459
rect 10320 26427 10360 26459
rect 10392 26427 10432 26459
rect 10464 26427 10504 26459
rect 10536 26427 10576 26459
rect 10608 26427 10648 26459
rect 10680 26427 10720 26459
rect 10752 26427 10792 26459
rect 10824 26427 10864 26459
rect 10896 26427 10936 26459
rect 10968 26427 11008 26459
rect 11040 26427 11080 26459
rect 11112 26427 11152 26459
rect 11184 26427 11224 26459
rect 11256 26427 11296 26459
rect 11328 26427 11368 26459
rect 11400 26427 11440 26459
rect 11472 26427 11512 26459
rect 11544 26427 11584 26459
rect 11616 26427 11656 26459
rect 11688 26427 11728 26459
rect 11760 26427 11800 26459
rect 11832 26427 11872 26459
rect 11904 26427 11944 26459
rect 11976 26427 12016 26459
rect 12048 26427 12088 26459
rect 12120 26427 12160 26459
rect 12192 26427 12232 26459
rect 12264 26427 12304 26459
rect 12336 26427 12376 26459
rect 12408 26427 12448 26459
rect 12480 26427 12520 26459
rect 12552 26427 12592 26459
rect 12624 26427 12664 26459
rect 12696 26427 12736 26459
rect 12768 26427 12808 26459
rect 12840 26427 12880 26459
rect 12912 26427 12952 26459
rect 12984 26427 13024 26459
rect 13056 26427 13096 26459
rect 13128 26427 13168 26459
rect 13200 26427 13240 26459
rect 13272 26427 13312 26459
rect 13344 26427 13384 26459
rect 13416 26427 13456 26459
rect 13488 26427 13528 26459
rect 13560 26427 13600 26459
rect 13632 26427 13672 26459
rect 13704 26427 13744 26459
rect 13776 26427 13816 26459
rect 13848 26427 13888 26459
rect 13920 26427 13960 26459
rect 13992 26427 14032 26459
rect 14064 26427 14104 26459
rect 14136 26427 14176 26459
rect 14208 26427 14248 26459
rect 14280 26427 14320 26459
rect 14352 26427 14392 26459
rect 14424 26427 14464 26459
rect 14496 26427 14536 26459
rect 14568 26427 14608 26459
rect 14640 26427 14680 26459
rect 14712 26427 14752 26459
rect 14784 26427 14824 26459
rect 14856 26427 14896 26459
rect 14928 26427 14968 26459
rect 15000 26427 15040 26459
rect 15072 26427 15112 26459
rect 15144 26427 15184 26459
rect 15216 26427 15256 26459
rect 15288 26427 15328 26459
rect 15360 26427 15400 26459
rect 15432 26427 15472 26459
rect 15504 26427 15544 26459
rect 15576 26427 15616 26459
rect 15648 26427 15688 26459
rect 15720 26427 15760 26459
rect 15792 26427 15832 26459
rect 15864 26427 15904 26459
rect 15936 26427 16000 26459
rect 0 26387 16000 26427
rect 0 26355 64 26387
rect 96 26355 136 26387
rect 168 26355 208 26387
rect 240 26355 280 26387
rect 312 26355 352 26387
rect 384 26355 424 26387
rect 456 26355 496 26387
rect 528 26355 568 26387
rect 600 26355 640 26387
rect 672 26355 712 26387
rect 744 26355 784 26387
rect 816 26355 856 26387
rect 888 26355 928 26387
rect 960 26355 1000 26387
rect 1032 26355 1072 26387
rect 1104 26355 1144 26387
rect 1176 26355 1216 26387
rect 1248 26355 1288 26387
rect 1320 26355 1360 26387
rect 1392 26355 1432 26387
rect 1464 26355 1504 26387
rect 1536 26355 1576 26387
rect 1608 26355 1648 26387
rect 1680 26355 1720 26387
rect 1752 26355 1792 26387
rect 1824 26355 1864 26387
rect 1896 26355 1936 26387
rect 1968 26355 2008 26387
rect 2040 26355 2080 26387
rect 2112 26355 2152 26387
rect 2184 26355 2224 26387
rect 2256 26355 2296 26387
rect 2328 26355 2368 26387
rect 2400 26355 2440 26387
rect 2472 26355 2512 26387
rect 2544 26355 2584 26387
rect 2616 26355 2656 26387
rect 2688 26355 2728 26387
rect 2760 26355 2800 26387
rect 2832 26355 2872 26387
rect 2904 26355 2944 26387
rect 2976 26355 3016 26387
rect 3048 26355 3088 26387
rect 3120 26355 3160 26387
rect 3192 26355 3232 26387
rect 3264 26355 3304 26387
rect 3336 26355 3376 26387
rect 3408 26355 3448 26387
rect 3480 26355 3520 26387
rect 3552 26355 3592 26387
rect 3624 26355 3664 26387
rect 3696 26355 3736 26387
rect 3768 26355 3808 26387
rect 3840 26355 3880 26387
rect 3912 26355 3952 26387
rect 3984 26355 4024 26387
rect 4056 26355 4096 26387
rect 4128 26355 4168 26387
rect 4200 26355 4240 26387
rect 4272 26355 4312 26387
rect 4344 26355 4384 26387
rect 4416 26355 4456 26387
rect 4488 26355 4528 26387
rect 4560 26355 4600 26387
rect 4632 26355 4672 26387
rect 4704 26355 4744 26387
rect 4776 26355 4816 26387
rect 4848 26355 4888 26387
rect 4920 26355 4960 26387
rect 4992 26355 5032 26387
rect 5064 26355 5104 26387
rect 5136 26355 5176 26387
rect 5208 26355 5248 26387
rect 5280 26355 5320 26387
rect 5352 26355 5392 26387
rect 5424 26355 5464 26387
rect 5496 26355 5536 26387
rect 5568 26355 5608 26387
rect 5640 26355 5680 26387
rect 5712 26355 5752 26387
rect 5784 26355 5824 26387
rect 5856 26355 5896 26387
rect 5928 26355 5968 26387
rect 6000 26355 6040 26387
rect 6072 26355 6112 26387
rect 6144 26355 6184 26387
rect 6216 26355 6256 26387
rect 6288 26355 6328 26387
rect 6360 26355 6400 26387
rect 6432 26355 6472 26387
rect 6504 26355 6544 26387
rect 6576 26355 6616 26387
rect 6648 26355 6688 26387
rect 6720 26355 6760 26387
rect 6792 26355 6832 26387
rect 6864 26355 6904 26387
rect 6936 26355 6976 26387
rect 7008 26355 7048 26387
rect 7080 26355 7120 26387
rect 7152 26355 7192 26387
rect 7224 26355 7264 26387
rect 7296 26355 7336 26387
rect 7368 26355 7408 26387
rect 7440 26355 7480 26387
rect 7512 26355 7552 26387
rect 7584 26355 7624 26387
rect 7656 26355 7696 26387
rect 7728 26355 7768 26387
rect 7800 26355 7840 26387
rect 7872 26355 7912 26387
rect 7944 26355 7984 26387
rect 8016 26355 8056 26387
rect 8088 26355 8128 26387
rect 8160 26355 8200 26387
rect 8232 26355 8272 26387
rect 8304 26355 8344 26387
rect 8376 26355 8416 26387
rect 8448 26355 8488 26387
rect 8520 26355 8560 26387
rect 8592 26355 8632 26387
rect 8664 26355 8704 26387
rect 8736 26355 8776 26387
rect 8808 26355 8848 26387
rect 8880 26355 8920 26387
rect 8952 26355 8992 26387
rect 9024 26355 9064 26387
rect 9096 26355 9136 26387
rect 9168 26355 9208 26387
rect 9240 26355 9280 26387
rect 9312 26355 9352 26387
rect 9384 26355 9424 26387
rect 9456 26355 9496 26387
rect 9528 26355 9568 26387
rect 9600 26355 9640 26387
rect 9672 26355 9712 26387
rect 9744 26355 9784 26387
rect 9816 26355 9856 26387
rect 9888 26355 9928 26387
rect 9960 26355 10000 26387
rect 10032 26355 10072 26387
rect 10104 26355 10144 26387
rect 10176 26355 10216 26387
rect 10248 26355 10288 26387
rect 10320 26355 10360 26387
rect 10392 26355 10432 26387
rect 10464 26355 10504 26387
rect 10536 26355 10576 26387
rect 10608 26355 10648 26387
rect 10680 26355 10720 26387
rect 10752 26355 10792 26387
rect 10824 26355 10864 26387
rect 10896 26355 10936 26387
rect 10968 26355 11008 26387
rect 11040 26355 11080 26387
rect 11112 26355 11152 26387
rect 11184 26355 11224 26387
rect 11256 26355 11296 26387
rect 11328 26355 11368 26387
rect 11400 26355 11440 26387
rect 11472 26355 11512 26387
rect 11544 26355 11584 26387
rect 11616 26355 11656 26387
rect 11688 26355 11728 26387
rect 11760 26355 11800 26387
rect 11832 26355 11872 26387
rect 11904 26355 11944 26387
rect 11976 26355 12016 26387
rect 12048 26355 12088 26387
rect 12120 26355 12160 26387
rect 12192 26355 12232 26387
rect 12264 26355 12304 26387
rect 12336 26355 12376 26387
rect 12408 26355 12448 26387
rect 12480 26355 12520 26387
rect 12552 26355 12592 26387
rect 12624 26355 12664 26387
rect 12696 26355 12736 26387
rect 12768 26355 12808 26387
rect 12840 26355 12880 26387
rect 12912 26355 12952 26387
rect 12984 26355 13024 26387
rect 13056 26355 13096 26387
rect 13128 26355 13168 26387
rect 13200 26355 13240 26387
rect 13272 26355 13312 26387
rect 13344 26355 13384 26387
rect 13416 26355 13456 26387
rect 13488 26355 13528 26387
rect 13560 26355 13600 26387
rect 13632 26355 13672 26387
rect 13704 26355 13744 26387
rect 13776 26355 13816 26387
rect 13848 26355 13888 26387
rect 13920 26355 13960 26387
rect 13992 26355 14032 26387
rect 14064 26355 14104 26387
rect 14136 26355 14176 26387
rect 14208 26355 14248 26387
rect 14280 26355 14320 26387
rect 14352 26355 14392 26387
rect 14424 26355 14464 26387
rect 14496 26355 14536 26387
rect 14568 26355 14608 26387
rect 14640 26355 14680 26387
rect 14712 26355 14752 26387
rect 14784 26355 14824 26387
rect 14856 26355 14896 26387
rect 14928 26355 14968 26387
rect 15000 26355 15040 26387
rect 15072 26355 15112 26387
rect 15144 26355 15184 26387
rect 15216 26355 15256 26387
rect 15288 26355 15328 26387
rect 15360 26355 15400 26387
rect 15432 26355 15472 26387
rect 15504 26355 15544 26387
rect 15576 26355 15616 26387
rect 15648 26355 15688 26387
rect 15720 26355 15760 26387
rect 15792 26355 15832 26387
rect 15864 26355 15904 26387
rect 15936 26355 16000 26387
rect 0 26315 16000 26355
rect 0 26283 64 26315
rect 96 26283 136 26315
rect 168 26283 208 26315
rect 240 26283 280 26315
rect 312 26283 352 26315
rect 384 26283 424 26315
rect 456 26283 496 26315
rect 528 26283 568 26315
rect 600 26283 640 26315
rect 672 26283 712 26315
rect 744 26283 784 26315
rect 816 26283 856 26315
rect 888 26283 928 26315
rect 960 26283 1000 26315
rect 1032 26283 1072 26315
rect 1104 26283 1144 26315
rect 1176 26283 1216 26315
rect 1248 26283 1288 26315
rect 1320 26283 1360 26315
rect 1392 26283 1432 26315
rect 1464 26283 1504 26315
rect 1536 26283 1576 26315
rect 1608 26283 1648 26315
rect 1680 26283 1720 26315
rect 1752 26283 1792 26315
rect 1824 26283 1864 26315
rect 1896 26283 1936 26315
rect 1968 26283 2008 26315
rect 2040 26283 2080 26315
rect 2112 26283 2152 26315
rect 2184 26283 2224 26315
rect 2256 26283 2296 26315
rect 2328 26283 2368 26315
rect 2400 26283 2440 26315
rect 2472 26283 2512 26315
rect 2544 26283 2584 26315
rect 2616 26283 2656 26315
rect 2688 26283 2728 26315
rect 2760 26283 2800 26315
rect 2832 26283 2872 26315
rect 2904 26283 2944 26315
rect 2976 26283 3016 26315
rect 3048 26283 3088 26315
rect 3120 26283 3160 26315
rect 3192 26283 3232 26315
rect 3264 26283 3304 26315
rect 3336 26283 3376 26315
rect 3408 26283 3448 26315
rect 3480 26283 3520 26315
rect 3552 26283 3592 26315
rect 3624 26283 3664 26315
rect 3696 26283 3736 26315
rect 3768 26283 3808 26315
rect 3840 26283 3880 26315
rect 3912 26283 3952 26315
rect 3984 26283 4024 26315
rect 4056 26283 4096 26315
rect 4128 26283 4168 26315
rect 4200 26283 4240 26315
rect 4272 26283 4312 26315
rect 4344 26283 4384 26315
rect 4416 26283 4456 26315
rect 4488 26283 4528 26315
rect 4560 26283 4600 26315
rect 4632 26283 4672 26315
rect 4704 26283 4744 26315
rect 4776 26283 4816 26315
rect 4848 26283 4888 26315
rect 4920 26283 4960 26315
rect 4992 26283 5032 26315
rect 5064 26283 5104 26315
rect 5136 26283 5176 26315
rect 5208 26283 5248 26315
rect 5280 26283 5320 26315
rect 5352 26283 5392 26315
rect 5424 26283 5464 26315
rect 5496 26283 5536 26315
rect 5568 26283 5608 26315
rect 5640 26283 5680 26315
rect 5712 26283 5752 26315
rect 5784 26283 5824 26315
rect 5856 26283 5896 26315
rect 5928 26283 5968 26315
rect 6000 26283 6040 26315
rect 6072 26283 6112 26315
rect 6144 26283 6184 26315
rect 6216 26283 6256 26315
rect 6288 26283 6328 26315
rect 6360 26283 6400 26315
rect 6432 26283 6472 26315
rect 6504 26283 6544 26315
rect 6576 26283 6616 26315
rect 6648 26283 6688 26315
rect 6720 26283 6760 26315
rect 6792 26283 6832 26315
rect 6864 26283 6904 26315
rect 6936 26283 6976 26315
rect 7008 26283 7048 26315
rect 7080 26283 7120 26315
rect 7152 26283 7192 26315
rect 7224 26283 7264 26315
rect 7296 26283 7336 26315
rect 7368 26283 7408 26315
rect 7440 26283 7480 26315
rect 7512 26283 7552 26315
rect 7584 26283 7624 26315
rect 7656 26283 7696 26315
rect 7728 26283 7768 26315
rect 7800 26283 7840 26315
rect 7872 26283 7912 26315
rect 7944 26283 7984 26315
rect 8016 26283 8056 26315
rect 8088 26283 8128 26315
rect 8160 26283 8200 26315
rect 8232 26283 8272 26315
rect 8304 26283 8344 26315
rect 8376 26283 8416 26315
rect 8448 26283 8488 26315
rect 8520 26283 8560 26315
rect 8592 26283 8632 26315
rect 8664 26283 8704 26315
rect 8736 26283 8776 26315
rect 8808 26283 8848 26315
rect 8880 26283 8920 26315
rect 8952 26283 8992 26315
rect 9024 26283 9064 26315
rect 9096 26283 9136 26315
rect 9168 26283 9208 26315
rect 9240 26283 9280 26315
rect 9312 26283 9352 26315
rect 9384 26283 9424 26315
rect 9456 26283 9496 26315
rect 9528 26283 9568 26315
rect 9600 26283 9640 26315
rect 9672 26283 9712 26315
rect 9744 26283 9784 26315
rect 9816 26283 9856 26315
rect 9888 26283 9928 26315
rect 9960 26283 10000 26315
rect 10032 26283 10072 26315
rect 10104 26283 10144 26315
rect 10176 26283 10216 26315
rect 10248 26283 10288 26315
rect 10320 26283 10360 26315
rect 10392 26283 10432 26315
rect 10464 26283 10504 26315
rect 10536 26283 10576 26315
rect 10608 26283 10648 26315
rect 10680 26283 10720 26315
rect 10752 26283 10792 26315
rect 10824 26283 10864 26315
rect 10896 26283 10936 26315
rect 10968 26283 11008 26315
rect 11040 26283 11080 26315
rect 11112 26283 11152 26315
rect 11184 26283 11224 26315
rect 11256 26283 11296 26315
rect 11328 26283 11368 26315
rect 11400 26283 11440 26315
rect 11472 26283 11512 26315
rect 11544 26283 11584 26315
rect 11616 26283 11656 26315
rect 11688 26283 11728 26315
rect 11760 26283 11800 26315
rect 11832 26283 11872 26315
rect 11904 26283 11944 26315
rect 11976 26283 12016 26315
rect 12048 26283 12088 26315
rect 12120 26283 12160 26315
rect 12192 26283 12232 26315
rect 12264 26283 12304 26315
rect 12336 26283 12376 26315
rect 12408 26283 12448 26315
rect 12480 26283 12520 26315
rect 12552 26283 12592 26315
rect 12624 26283 12664 26315
rect 12696 26283 12736 26315
rect 12768 26283 12808 26315
rect 12840 26283 12880 26315
rect 12912 26283 12952 26315
rect 12984 26283 13024 26315
rect 13056 26283 13096 26315
rect 13128 26283 13168 26315
rect 13200 26283 13240 26315
rect 13272 26283 13312 26315
rect 13344 26283 13384 26315
rect 13416 26283 13456 26315
rect 13488 26283 13528 26315
rect 13560 26283 13600 26315
rect 13632 26283 13672 26315
rect 13704 26283 13744 26315
rect 13776 26283 13816 26315
rect 13848 26283 13888 26315
rect 13920 26283 13960 26315
rect 13992 26283 14032 26315
rect 14064 26283 14104 26315
rect 14136 26283 14176 26315
rect 14208 26283 14248 26315
rect 14280 26283 14320 26315
rect 14352 26283 14392 26315
rect 14424 26283 14464 26315
rect 14496 26283 14536 26315
rect 14568 26283 14608 26315
rect 14640 26283 14680 26315
rect 14712 26283 14752 26315
rect 14784 26283 14824 26315
rect 14856 26283 14896 26315
rect 14928 26283 14968 26315
rect 15000 26283 15040 26315
rect 15072 26283 15112 26315
rect 15144 26283 15184 26315
rect 15216 26283 15256 26315
rect 15288 26283 15328 26315
rect 15360 26283 15400 26315
rect 15432 26283 15472 26315
rect 15504 26283 15544 26315
rect 15576 26283 15616 26315
rect 15648 26283 15688 26315
rect 15720 26283 15760 26315
rect 15792 26283 15832 26315
rect 15864 26283 15904 26315
rect 15936 26283 16000 26315
rect 0 26243 16000 26283
rect 0 26211 64 26243
rect 96 26211 136 26243
rect 168 26211 208 26243
rect 240 26211 280 26243
rect 312 26211 352 26243
rect 384 26211 424 26243
rect 456 26211 496 26243
rect 528 26211 568 26243
rect 600 26211 640 26243
rect 672 26211 712 26243
rect 744 26211 784 26243
rect 816 26211 856 26243
rect 888 26211 928 26243
rect 960 26211 1000 26243
rect 1032 26211 1072 26243
rect 1104 26211 1144 26243
rect 1176 26211 1216 26243
rect 1248 26211 1288 26243
rect 1320 26211 1360 26243
rect 1392 26211 1432 26243
rect 1464 26211 1504 26243
rect 1536 26211 1576 26243
rect 1608 26211 1648 26243
rect 1680 26211 1720 26243
rect 1752 26211 1792 26243
rect 1824 26211 1864 26243
rect 1896 26211 1936 26243
rect 1968 26211 2008 26243
rect 2040 26211 2080 26243
rect 2112 26211 2152 26243
rect 2184 26211 2224 26243
rect 2256 26211 2296 26243
rect 2328 26211 2368 26243
rect 2400 26211 2440 26243
rect 2472 26211 2512 26243
rect 2544 26211 2584 26243
rect 2616 26211 2656 26243
rect 2688 26211 2728 26243
rect 2760 26211 2800 26243
rect 2832 26211 2872 26243
rect 2904 26211 2944 26243
rect 2976 26211 3016 26243
rect 3048 26211 3088 26243
rect 3120 26211 3160 26243
rect 3192 26211 3232 26243
rect 3264 26211 3304 26243
rect 3336 26211 3376 26243
rect 3408 26211 3448 26243
rect 3480 26211 3520 26243
rect 3552 26211 3592 26243
rect 3624 26211 3664 26243
rect 3696 26211 3736 26243
rect 3768 26211 3808 26243
rect 3840 26211 3880 26243
rect 3912 26211 3952 26243
rect 3984 26211 4024 26243
rect 4056 26211 4096 26243
rect 4128 26211 4168 26243
rect 4200 26211 4240 26243
rect 4272 26211 4312 26243
rect 4344 26211 4384 26243
rect 4416 26211 4456 26243
rect 4488 26211 4528 26243
rect 4560 26211 4600 26243
rect 4632 26211 4672 26243
rect 4704 26211 4744 26243
rect 4776 26211 4816 26243
rect 4848 26211 4888 26243
rect 4920 26211 4960 26243
rect 4992 26211 5032 26243
rect 5064 26211 5104 26243
rect 5136 26211 5176 26243
rect 5208 26211 5248 26243
rect 5280 26211 5320 26243
rect 5352 26211 5392 26243
rect 5424 26211 5464 26243
rect 5496 26211 5536 26243
rect 5568 26211 5608 26243
rect 5640 26211 5680 26243
rect 5712 26211 5752 26243
rect 5784 26211 5824 26243
rect 5856 26211 5896 26243
rect 5928 26211 5968 26243
rect 6000 26211 6040 26243
rect 6072 26211 6112 26243
rect 6144 26211 6184 26243
rect 6216 26211 6256 26243
rect 6288 26211 6328 26243
rect 6360 26211 6400 26243
rect 6432 26211 6472 26243
rect 6504 26211 6544 26243
rect 6576 26211 6616 26243
rect 6648 26211 6688 26243
rect 6720 26211 6760 26243
rect 6792 26211 6832 26243
rect 6864 26211 6904 26243
rect 6936 26211 6976 26243
rect 7008 26211 7048 26243
rect 7080 26211 7120 26243
rect 7152 26211 7192 26243
rect 7224 26211 7264 26243
rect 7296 26211 7336 26243
rect 7368 26211 7408 26243
rect 7440 26211 7480 26243
rect 7512 26211 7552 26243
rect 7584 26211 7624 26243
rect 7656 26211 7696 26243
rect 7728 26211 7768 26243
rect 7800 26211 7840 26243
rect 7872 26211 7912 26243
rect 7944 26211 7984 26243
rect 8016 26211 8056 26243
rect 8088 26211 8128 26243
rect 8160 26211 8200 26243
rect 8232 26211 8272 26243
rect 8304 26211 8344 26243
rect 8376 26211 8416 26243
rect 8448 26211 8488 26243
rect 8520 26211 8560 26243
rect 8592 26211 8632 26243
rect 8664 26211 8704 26243
rect 8736 26211 8776 26243
rect 8808 26211 8848 26243
rect 8880 26211 8920 26243
rect 8952 26211 8992 26243
rect 9024 26211 9064 26243
rect 9096 26211 9136 26243
rect 9168 26211 9208 26243
rect 9240 26211 9280 26243
rect 9312 26211 9352 26243
rect 9384 26211 9424 26243
rect 9456 26211 9496 26243
rect 9528 26211 9568 26243
rect 9600 26211 9640 26243
rect 9672 26211 9712 26243
rect 9744 26211 9784 26243
rect 9816 26211 9856 26243
rect 9888 26211 9928 26243
rect 9960 26211 10000 26243
rect 10032 26211 10072 26243
rect 10104 26211 10144 26243
rect 10176 26211 10216 26243
rect 10248 26211 10288 26243
rect 10320 26211 10360 26243
rect 10392 26211 10432 26243
rect 10464 26211 10504 26243
rect 10536 26211 10576 26243
rect 10608 26211 10648 26243
rect 10680 26211 10720 26243
rect 10752 26211 10792 26243
rect 10824 26211 10864 26243
rect 10896 26211 10936 26243
rect 10968 26211 11008 26243
rect 11040 26211 11080 26243
rect 11112 26211 11152 26243
rect 11184 26211 11224 26243
rect 11256 26211 11296 26243
rect 11328 26211 11368 26243
rect 11400 26211 11440 26243
rect 11472 26211 11512 26243
rect 11544 26211 11584 26243
rect 11616 26211 11656 26243
rect 11688 26211 11728 26243
rect 11760 26211 11800 26243
rect 11832 26211 11872 26243
rect 11904 26211 11944 26243
rect 11976 26211 12016 26243
rect 12048 26211 12088 26243
rect 12120 26211 12160 26243
rect 12192 26211 12232 26243
rect 12264 26211 12304 26243
rect 12336 26211 12376 26243
rect 12408 26211 12448 26243
rect 12480 26211 12520 26243
rect 12552 26211 12592 26243
rect 12624 26211 12664 26243
rect 12696 26211 12736 26243
rect 12768 26211 12808 26243
rect 12840 26211 12880 26243
rect 12912 26211 12952 26243
rect 12984 26211 13024 26243
rect 13056 26211 13096 26243
rect 13128 26211 13168 26243
rect 13200 26211 13240 26243
rect 13272 26211 13312 26243
rect 13344 26211 13384 26243
rect 13416 26211 13456 26243
rect 13488 26211 13528 26243
rect 13560 26211 13600 26243
rect 13632 26211 13672 26243
rect 13704 26211 13744 26243
rect 13776 26211 13816 26243
rect 13848 26211 13888 26243
rect 13920 26211 13960 26243
rect 13992 26211 14032 26243
rect 14064 26211 14104 26243
rect 14136 26211 14176 26243
rect 14208 26211 14248 26243
rect 14280 26211 14320 26243
rect 14352 26211 14392 26243
rect 14424 26211 14464 26243
rect 14496 26211 14536 26243
rect 14568 26211 14608 26243
rect 14640 26211 14680 26243
rect 14712 26211 14752 26243
rect 14784 26211 14824 26243
rect 14856 26211 14896 26243
rect 14928 26211 14968 26243
rect 15000 26211 15040 26243
rect 15072 26211 15112 26243
rect 15144 26211 15184 26243
rect 15216 26211 15256 26243
rect 15288 26211 15328 26243
rect 15360 26211 15400 26243
rect 15432 26211 15472 26243
rect 15504 26211 15544 26243
rect 15576 26211 15616 26243
rect 15648 26211 15688 26243
rect 15720 26211 15760 26243
rect 15792 26211 15832 26243
rect 15864 26211 15904 26243
rect 15936 26211 16000 26243
rect 0 26171 16000 26211
rect 0 26139 64 26171
rect 96 26139 136 26171
rect 168 26139 208 26171
rect 240 26139 280 26171
rect 312 26139 352 26171
rect 384 26139 424 26171
rect 456 26139 496 26171
rect 528 26139 568 26171
rect 600 26139 640 26171
rect 672 26139 712 26171
rect 744 26139 784 26171
rect 816 26139 856 26171
rect 888 26139 928 26171
rect 960 26139 1000 26171
rect 1032 26139 1072 26171
rect 1104 26139 1144 26171
rect 1176 26139 1216 26171
rect 1248 26139 1288 26171
rect 1320 26139 1360 26171
rect 1392 26139 1432 26171
rect 1464 26139 1504 26171
rect 1536 26139 1576 26171
rect 1608 26139 1648 26171
rect 1680 26139 1720 26171
rect 1752 26139 1792 26171
rect 1824 26139 1864 26171
rect 1896 26139 1936 26171
rect 1968 26139 2008 26171
rect 2040 26139 2080 26171
rect 2112 26139 2152 26171
rect 2184 26139 2224 26171
rect 2256 26139 2296 26171
rect 2328 26139 2368 26171
rect 2400 26139 2440 26171
rect 2472 26139 2512 26171
rect 2544 26139 2584 26171
rect 2616 26139 2656 26171
rect 2688 26139 2728 26171
rect 2760 26139 2800 26171
rect 2832 26139 2872 26171
rect 2904 26139 2944 26171
rect 2976 26139 3016 26171
rect 3048 26139 3088 26171
rect 3120 26139 3160 26171
rect 3192 26139 3232 26171
rect 3264 26139 3304 26171
rect 3336 26139 3376 26171
rect 3408 26139 3448 26171
rect 3480 26139 3520 26171
rect 3552 26139 3592 26171
rect 3624 26139 3664 26171
rect 3696 26139 3736 26171
rect 3768 26139 3808 26171
rect 3840 26139 3880 26171
rect 3912 26139 3952 26171
rect 3984 26139 4024 26171
rect 4056 26139 4096 26171
rect 4128 26139 4168 26171
rect 4200 26139 4240 26171
rect 4272 26139 4312 26171
rect 4344 26139 4384 26171
rect 4416 26139 4456 26171
rect 4488 26139 4528 26171
rect 4560 26139 4600 26171
rect 4632 26139 4672 26171
rect 4704 26139 4744 26171
rect 4776 26139 4816 26171
rect 4848 26139 4888 26171
rect 4920 26139 4960 26171
rect 4992 26139 5032 26171
rect 5064 26139 5104 26171
rect 5136 26139 5176 26171
rect 5208 26139 5248 26171
rect 5280 26139 5320 26171
rect 5352 26139 5392 26171
rect 5424 26139 5464 26171
rect 5496 26139 5536 26171
rect 5568 26139 5608 26171
rect 5640 26139 5680 26171
rect 5712 26139 5752 26171
rect 5784 26139 5824 26171
rect 5856 26139 5896 26171
rect 5928 26139 5968 26171
rect 6000 26139 6040 26171
rect 6072 26139 6112 26171
rect 6144 26139 6184 26171
rect 6216 26139 6256 26171
rect 6288 26139 6328 26171
rect 6360 26139 6400 26171
rect 6432 26139 6472 26171
rect 6504 26139 6544 26171
rect 6576 26139 6616 26171
rect 6648 26139 6688 26171
rect 6720 26139 6760 26171
rect 6792 26139 6832 26171
rect 6864 26139 6904 26171
rect 6936 26139 6976 26171
rect 7008 26139 7048 26171
rect 7080 26139 7120 26171
rect 7152 26139 7192 26171
rect 7224 26139 7264 26171
rect 7296 26139 7336 26171
rect 7368 26139 7408 26171
rect 7440 26139 7480 26171
rect 7512 26139 7552 26171
rect 7584 26139 7624 26171
rect 7656 26139 7696 26171
rect 7728 26139 7768 26171
rect 7800 26139 7840 26171
rect 7872 26139 7912 26171
rect 7944 26139 7984 26171
rect 8016 26139 8056 26171
rect 8088 26139 8128 26171
rect 8160 26139 8200 26171
rect 8232 26139 8272 26171
rect 8304 26139 8344 26171
rect 8376 26139 8416 26171
rect 8448 26139 8488 26171
rect 8520 26139 8560 26171
rect 8592 26139 8632 26171
rect 8664 26139 8704 26171
rect 8736 26139 8776 26171
rect 8808 26139 8848 26171
rect 8880 26139 8920 26171
rect 8952 26139 8992 26171
rect 9024 26139 9064 26171
rect 9096 26139 9136 26171
rect 9168 26139 9208 26171
rect 9240 26139 9280 26171
rect 9312 26139 9352 26171
rect 9384 26139 9424 26171
rect 9456 26139 9496 26171
rect 9528 26139 9568 26171
rect 9600 26139 9640 26171
rect 9672 26139 9712 26171
rect 9744 26139 9784 26171
rect 9816 26139 9856 26171
rect 9888 26139 9928 26171
rect 9960 26139 10000 26171
rect 10032 26139 10072 26171
rect 10104 26139 10144 26171
rect 10176 26139 10216 26171
rect 10248 26139 10288 26171
rect 10320 26139 10360 26171
rect 10392 26139 10432 26171
rect 10464 26139 10504 26171
rect 10536 26139 10576 26171
rect 10608 26139 10648 26171
rect 10680 26139 10720 26171
rect 10752 26139 10792 26171
rect 10824 26139 10864 26171
rect 10896 26139 10936 26171
rect 10968 26139 11008 26171
rect 11040 26139 11080 26171
rect 11112 26139 11152 26171
rect 11184 26139 11224 26171
rect 11256 26139 11296 26171
rect 11328 26139 11368 26171
rect 11400 26139 11440 26171
rect 11472 26139 11512 26171
rect 11544 26139 11584 26171
rect 11616 26139 11656 26171
rect 11688 26139 11728 26171
rect 11760 26139 11800 26171
rect 11832 26139 11872 26171
rect 11904 26139 11944 26171
rect 11976 26139 12016 26171
rect 12048 26139 12088 26171
rect 12120 26139 12160 26171
rect 12192 26139 12232 26171
rect 12264 26139 12304 26171
rect 12336 26139 12376 26171
rect 12408 26139 12448 26171
rect 12480 26139 12520 26171
rect 12552 26139 12592 26171
rect 12624 26139 12664 26171
rect 12696 26139 12736 26171
rect 12768 26139 12808 26171
rect 12840 26139 12880 26171
rect 12912 26139 12952 26171
rect 12984 26139 13024 26171
rect 13056 26139 13096 26171
rect 13128 26139 13168 26171
rect 13200 26139 13240 26171
rect 13272 26139 13312 26171
rect 13344 26139 13384 26171
rect 13416 26139 13456 26171
rect 13488 26139 13528 26171
rect 13560 26139 13600 26171
rect 13632 26139 13672 26171
rect 13704 26139 13744 26171
rect 13776 26139 13816 26171
rect 13848 26139 13888 26171
rect 13920 26139 13960 26171
rect 13992 26139 14032 26171
rect 14064 26139 14104 26171
rect 14136 26139 14176 26171
rect 14208 26139 14248 26171
rect 14280 26139 14320 26171
rect 14352 26139 14392 26171
rect 14424 26139 14464 26171
rect 14496 26139 14536 26171
rect 14568 26139 14608 26171
rect 14640 26139 14680 26171
rect 14712 26139 14752 26171
rect 14784 26139 14824 26171
rect 14856 26139 14896 26171
rect 14928 26139 14968 26171
rect 15000 26139 15040 26171
rect 15072 26139 15112 26171
rect 15144 26139 15184 26171
rect 15216 26139 15256 26171
rect 15288 26139 15328 26171
rect 15360 26139 15400 26171
rect 15432 26139 15472 26171
rect 15504 26139 15544 26171
rect 15576 26139 15616 26171
rect 15648 26139 15688 26171
rect 15720 26139 15760 26171
rect 15792 26139 15832 26171
rect 15864 26139 15904 26171
rect 15936 26139 16000 26171
rect 0 26099 16000 26139
rect 0 26067 64 26099
rect 96 26067 136 26099
rect 168 26067 208 26099
rect 240 26067 280 26099
rect 312 26067 352 26099
rect 384 26067 424 26099
rect 456 26067 496 26099
rect 528 26067 568 26099
rect 600 26067 640 26099
rect 672 26067 712 26099
rect 744 26067 784 26099
rect 816 26067 856 26099
rect 888 26067 928 26099
rect 960 26067 1000 26099
rect 1032 26067 1072 26099
rect 1104 26067 1144 26099
rect 1176 26067 1216 26099
rect 1248 26067 1288 26099
rect 1320 26067 1360 26099
rect 1392 26067 1432 26099
rect 1464 26067 1504 26099
rect 1536 26067 1576 26099
rect 1608 26067 1648 26099
rect 1680 26067 1720 26099
rect 1752 26067 1792 26099
rect 1824 26067 1864 26099
rect 1896 26067 1936 26099
rect 1968 26067 2008 26099
rect 2040 26067 2080 26099
rect 2112 26067 2152 26099
rect 2184 26067 2224 26099
rect 2256 26067 2296 26099
rect 2328 26067 2368 26099
rect 2400 26067 2440 26099
rect 2472 26067 2512 26099
rect 2544 26067 2584 26099
rect 2616 26067 2656 26099
rect 2688 26067 2728 26099
rect 2760 26067 2800 26099
rect 2832 26067 2872 26099
rect 2904 26067 2944 26099
rect 2976 26067 3016 26099
rect 3048 26067 3088 26099
rect 3120 26067 3160 26099
rect 3192 26067 3232 26099
rect 3264 26067 3304 26099
rect 3336 26067 3376 26099
rect 3408 26067 3448 26099
rect 3480 26067 3520 26099
rect 3552 26067 3592 26099
rect 3624 26067 3664 26099
rect 3696 26067 3736 26099
rect 3768 26067 3808 26099
rect 3840 26067 3880 26099
rect 3912 26067 3952 26099
rect 3984 26067 4024 26099
rect 4056 26067 4096 26099
rect 4128 26067 4168 26099
rect 4200 26067 4240 26099
rect 4272 26067 4312 26099
rect 4344 26067 4384 26099
rect 4416 26067 4456 26099
rect 4488 26067 4528 26099
rect 4560 26067 4600 26099
rect 4632 26067 4672 26099
rect 4704 26067 4744 26099
rect 4776 26067 4816 26099
rect 4848 26067 4888 26099
rect 4920 26067 4960 26099
rect 4992 26067 5032 26099
rect 5064 26067 5104 26099
rect 5136 26067 5176 26099
rect 5208 26067 5248 26099
rect 5280 26067 5320 26099
rect 5352 26067 5392 26099
rect 5424 26067 5464 26099
rect 5496 26067 5536 26099
rect 5568 26067 5608 26099
rect 5640 26067 5680 26099
rect 5712 26067 5752 26099
rect 5784 26067 5824 26099
rect 5856 26067 5896 26099
rect 5928 26067 5968 26099
rect 6000 26067 6040 26099
rect 6072 26067 6112 26099
rect 6144 26067 6184 26099
rect 6216 26067 6256 26099
rect 6288 26067 6328 26099
rect 6360 26067 6400 26099
rect 6432 26067 6472 26099
rect 6504 26067 6544 26099
rect 6576 26067 6616 26099
rect 6648 26067 6688 26099
rect 6720 26067 6760 26099
rect 6792 26067 6832 26099
rect 6864 26067 6904 26099
rect 6936 26067 6976 26099
rect 7008 26067 7048 26099
rect 7080 26067 7120 26099
rect 7152 26067 7192 26099
rect 7224 26067 7264 26099
rect 7296 26067 7336 26099
rect 7368 26067 7408 26099
rect 7440 26067 7480 26099
rect 7512 26067 7552 26099
rect 7584 26067 7624 26099
rect 7656 26067 7696 26099
rect 7728 26067 7768 26099
rect 7800 26067 7840 26099
rect 7872 26067 7912 26099
rect 7944 26067 7984 26099
rect 8016 26067 8056 26099
rect 8088 26067 8128 26099
rect 8160 26067 8200 26099
rect 8232 26067 8272 26099
rect 8304 26067 8344 26099
rect 8376 26067 8416 26099
rect 8448 26067 8488 26099
rect 8520 26067 8560 26099
rect 8592 26067 8632 26099
rect 8664 26067 8704 26099
rect 8736 26067 8776 26099
rect 8808 26067 8848 26099
rect 8880 26067 8920 26099
rect 8952 26067 8992 26099
rect 9024 26067 9064 26099
rect 9096 26067 9136 26099
rect 9168 26067 9208 26099
rect 9240 26067 9280 26099
rect 9312 26067 9352 26099
rect 9384 26067 9424 26099
rect 9456 26067 9496 26099
rect 9528 26067 9568 26099
rect 9600 26067 9640 26099
rect 9672 26067 9712 26099
rect 9744 26067 9784 26099
rect 9816 26067 9856 26099
rect 9888 26067 9928 26099
rect 9960 26067 10000 26099
rect 10032 26067 10072 26099
rect 10104 26067 10144 26099
rect 10176 26067 10216 26099
rect 10248 26067 10288 26099
rect 10320 26067 10360 26099
rect 10392 26067 10432 26099
rect 10464 26067 10504 26099
rect 10536 26067 10576 26099
rect 10608 26067 10648 26099
rect 10680 26067 10720 26099
rect 10752 26067 10792 26099
rect 10824 26067 10864 26099
rect 10896 26067 10936 26099
rect 10968 26067 11008 26099
rect 11040 26067 11080 26099
rect 11112 26067 11152 26099
rect 11184 26067 11224 26099
rect 11256 26067 11296 26099
rect 11328 26067 11368 26099
rect 11400 26067 11440 26099
rect 11472 26067 11512 26099
rect 11544 26067 11584 26099
rect 11616 26067 11656 26099
rect 11688 26067 11728 26099
rect 11760 26067 11800 26099
rect 11832 26067 11872 26099
rect 11904 26067 11944 26099
rect 11976 26067 12016 26099
rect 12048 26067 12088 26099
rect 12120 26067 12160 26099
rect 12192 26067 12232 26099
rect 12264 26067 12304 26099
rect 12336 26067 12376 26099
rect 12408 26067 12448 26099
rect 12480 26067 12520 26099
rect 12552 26067 12592 26099
rect 12624 26067 12664 26099
rect 12696 26067 12736 26099
rect 12768 26067 12808 26099
rect 12840 26067 12880 26099
rect 12912 26067 12952 26099
rect 12984 26067 13024 26099
rect 13056 26067 13096 26099
rect 13128 26067 13168 26099
rect 13200 26067 13240 26099
rect 13272 26067 13312 26099
rect 13344 26067 13384 26099
rect 13416 26067 13456 26099
rect 13488 26067 13528 26099
rect 13560 26067 13600 26099
rect 13632 26067 13672 26099
rect 13704 26067 13744 26099
rect 13776 26067 13816 26099
rect 13848 26067 13888 26099
rect 13920 26067 13960 26099
rect 13992 26067 14032 26099
rect 14064 26067 14104 26099
rect 14136 26067 14176 26099
rect 14208 26067 14248 26099
rect 14280 26067 14320 26099
rect 14352 26067 14392 26099
rect 14424 26067 14464 26099
rect 14496 26067 14536 26099
rect 14568 26067 14608 26099
rect 14640 26067 14680 26099
rect 14712 26067 14752 26099
rect 14784 26067 14824 26099
rect 14856 26067 14896 26099
rect 14928 26067 14968 26099
rect 15000 26067 15040 26099
rect 15072 26067 15112 26099
rect 15144 26067 15184 26099
rect 15216 26067 15256 26099
rect 15288 26067 15328 26099
rect 15360 26067 15400 26099
rect 15432 26067 15472 26099
rect 15504 26067 15544 26099
rect 15576 26067 15616 26099
rect 15648 26067 15688 26099
rect 15720 26067 15760 26099
rect 15792 26067 15832 26099
rect 15864 26067 15904 26099
rect 15936 26067 16000 26099
rect 0 26027 16000 26067
rect 0 25995 64 26027
rect 96 25995 136 26027
rect 168 25995 208 26027
rect 240 25995 280 26027
rect 312 25995 352 26027
rect 384 25995 424 26027
rect 456 25995 496 26027
rect 528 25995 568 26027
rect 600 25995 640 26027
rect 672 25995 712 26027
rect 744 25995 784 26027
rect 816 25995 856 26027
rect 888 25995 928 26027
rect 960 25995 1000 26027
rect 1032 25995 1072 26027
rect 1104 25995 1144 26027
rect 1176 25995 1216 26027
rect 1248 25995 1288 26027
rect 1320 25995 1360 26027
rect 1392 25995 1432 26027
rect 1464 25995 1504 26027
rect 1536 25995 1576 26027
rect 1608 25995 1648 26027
rect 1680 25995 1720 26027
rect 1752 25995 1792 26027
rect 1824 25995 1864 26027
rect 1896 25995 1936 26027
rect 1968 25995 2008 26027
rect 2040 25995 2080 26027
rect 2112 25995 2152 26027
rect 2184 25995 2224 26027
rect 2256 25995 2296 26027
rect 2328 25995 2368 26027
rect 2400 25995 2440 26027
rect 2472 25995 2512 26027
rect 2544 25995 2584 26027
rect 2616 25995 2656 26027
rect 2688 25995 2728 26027
rect 2760 25995 2800 26027
rect 2832 25995 2872 26027
rect 2904 25995 2944 26027
rect 2976 25995 3016 26027
rect 3048 25995 3088 26027
rect 3120 25995 3160 26027
rect 3192 25995 3232 26027
rect 3264 25995 3304 26027
rect 3336 25995 3376 26027
rect 3408 25995 3448 26027
rect 3480 25995 3520 26027
rect 3552 25995 3592 26027
rect 3624 25995 3664 26027
rect 3696 25995 3736 26027
rect 3768 25995 3808 26027
rect 3840 25995 3880 26027
rect 3912 25995 3952 26027
rect 3984 25995 4024 26027
rect 4056 25995 4096 26027
rect 4128 25995 4168 26027
rect 4200 25995 4240 26027
rect 4272 25995 4312 26027
rect 4344 25995 4384 26027
rect 4416 25995 4456 26027
rect 4488 25995 4528 26027
rect 4560 25995 4600 26027
rect 4632 25995 4672 26027
rect 4704 25995 4744 26027
rect 4776 25995 4816 26027
rect 4848 25995 4888 26027
rect 4920 25995 4960 26027
rect 4992 25995 5032 26027
rect 5064 25995 5104 26027
rect 5136 25995 5176 26027
rect 5208 25995 5248 26027
rect 5280 25995 5320 26027
rect 5352 25995 5392 26027
rect 5424 25995 5464 26027
rect 5496 25995 5536 26027
rect 5568 25995 5608 26027
rect 5640 25995 5680 26027
rect 5712 25995 5752 26027
rect 5784 25995 5824 26027
rect 5856 25995 5896 26027
rect 5928 25995 5968 26027
rect 6000 25995 6040 26027
rect 6072 25995 6112 26027
rect 6144 25995 6184 26027
rect 6216 25995 6256 26027
rect 6288 25995 6328 26027
rect 6360 25995 6400 26027
rect 6432 25995 6472 26027
rect 6504 25995 6544 26027
rect 6576 25995 6616 26027
rect 6648 25995 6688 26027
rect 6720 25995 6760 26027
rect 6792 25995 6832 26027
rect 6864 25995 6904 26027
rect 6936 25995 6976 26027
rect 7008 25995 7048 26027
rect 7080 25995 7120 26027
rect 7152 25995 7192 26027
rect 7224 25995 7264 26027
rect 7296 25995 7336 26027
rect 7368 25995 7408 26027
rect 7440 25995 7480 26027
rect 7512 25995 7552 26027
rect 7584 25995 7624 26027
rect 7656 25995 7696 26027
rect 7728 25995 7768 26027
rect 7800 25995 7840 26027
rect 7872 25995 7912 26027
rect 7944 25995 7984 26027
rect 8016 25995 8056 26027
rect 8088 25995 8128 26027
rect 8160 25995 8200 26027
rect 8232 25995 8272 26027
rect 8304 25995 8344 26027
rect 8376 25995 8416 26027
rect 8448 25995 8488 26027
rect 8520 25995 8560 26027
rect 8592 25995 8632 26027
rect 8664 25995 8704 26027
rect 8736 25995 8776 26027
rect 8808 25995 8848 26027
rect 8880 25995 8920 26027
rect 8952 25995 8992 26027
rect 9024 25995 9064 26027
rect 9096 25995 9136 26027
rect 9168 25995 9208 26027
rect 9240 25995 9280 26027
rect 9312 25995 9352 26027
rect 9384 25995 9424 26027
rect 9456 25995 9496 26027
rect 9528 25995 9568 26027
rect 9600 25995 9640 26027
rect 9672 25995 9712 26027
rect 9744 25995 9784 26027
rect 9816 25995 9856 26027
rect 9888 25995 9928 26027
rect 9960 25995 10000 26027
rect 10032 25995 10072 26027
rect 10104 25995 10144 26027
rect 10176 25995 10216 26027
rect 10248 25995 10288 26027
rect 10320 25995 10360 26027
rect 10392 25995 10432 26027
rect 10464 25995 10504 26027
rect 10536 25995 10576 26027
rect 10608 25995 10648 26027
rect 10680 25995 10720 26027
rect 10752 25995 10792 26027
rect 10824 25995 10864 26027
rect 10896 25995 10936 26027
rect 10968 25995 11008 26027
rect 11040 25995 11080 26027
rect 11112 25995 11152 26027
rect 11184 25995 11224 26027
rect 11256 25995 11296 26027
rect 11328 25995 11368 26027
rect 11400 25995 11440 26027
rect 11472 25995 11512 26027
rect 11544 25995 11584 26027
rect 11616 25995 11656 26027
rect 11688 25995 11728 26027
rect 11760 25995 11800 26027
rect 11832 25995 11872 26027
rect 11904 25995 11944 26027
rect 11976 25995 12016 26027
rect 12048 25995 12088 26027
rect 12120 25995 12160 26027
rect 12192 25995 12232 26027
rect 12264 25995 12304 26027
rect 12336 25995 12376 26027
rect 12408 25995 12448 26027
rect 12480 25995 12520 26027
rect 12552 25995 12592 26027
rect 12624 25995 12664 26027
rect 12696 25995 12736 26027
rect 12768 25995 12808 26027
rect 12840 25995 12880 26027
rect 12912 25995 12952 26027
rect 12984 25995 13024 26027
rect 13056 25995 13096 26027
rect 13128 25995 13168 26027
rect 13200 25995 13240 26027
rect 13272 25995 13312 26027
rect 13344 25995 13384 26027
rect 13416 25995 13456 26027
rect 13488 25995 13528 26027
rect 13560 25995 13600 26027
rect 13632 25995 13672 26027
rect 13704 25995 13744 26027
rect 13776 25995 13816 26027
rect 13848 25995 13888 26027
rect 13920 25995 13960 26027
rect 13992 25995 14032 26027
rect 14064 25995 14104 26027
rect 14136 25995 14176 26027
rect 14208 25995 14248 26027
rect 14280 25995 14320 26027
rect 14352 25995 14392 26027
rect 14424 25995 14464 26027
rect 14496 25995 14536 26027
rect 14568 25995 14608 26027
rect 14640 25995 14680 26027
rect 14712 25995 14752 26027
rect 14784 25995 14824 26027
rect 14856 25995 14896 26027
rect 14928 25995 14968 26027
rect 15000 25995 15040 26027
rect 15072 25995 15112 26027
rect 15144 25995 15184 26027
rect 15216 25995 15256 26027
rect 15288 25995 15328 26027
rect 15360 25995 15400 26027
rect 15432 25995 15472 26027
rect 15504 25995 15544 26027
rect 15576 25995 15616 26027
rect 15648 25995 15688 26027
rect 15720 25995 15760 26027
rect 15792 25995 15832 26027
rect 15864 25995 15904 26027
rect 15936 25995 16000 26027
rect 0 25955 16000 25995
rect 0 25923 64 25955
rect 96 25923 136 25955
rect 168 25923 208 25955
rect 240 25923 280 25955
rect 312 25923 352 25955
rect 384 25923 424 25955
rect 456 25923 496 25955
rect 528 25923 568 25955
rect 600 25923 640 25955
rect 672 25923 712 25955
rect 744 25923 784 25955
rect 816 25923 856 25955
rect 888 25923 928 25955
rect 960 25923 1000 25955
rect 1032 25923 1072 25955
rect 1104 25923 1144 25955
rect 1176 25923 1216 25955
rect 1248 25923 1288 25955
rect 1320 25923 1360 25955
rect 1392 25923 1432 25955
rect 1464 25923 1504 25955
rect 1536 25923 1576 25955
rect 1608 25923 1648 25955
rect 1680 25923 1720 25955
rect 1752 25923 1792 25955
rect 1824 25923 1864 25955
rect 1896 25923 1936 25955
rect 1968 25923 2008 25955
rect 2040 25923 2080 25955
rect 2112 25923 2152 25955
rect 2184 25923 2224 25955
rect 2256 25923 2296 25955
rect 2328 25923 2368 25955
rect 2400 25923 2440 25955
rect 2472 25923 2512 25955
rect 2544 25923 2584 25955
rect 2616 25923 2656 25955
rect 2688 25923 2728 25955
rect 2760 25923 2800 25955
rect 2832 25923 2872 25955
rect 2904 25923 2944 25955
rect 2976 25923 3016 25955
rect 3048 25923 3088 25955
rect 3120 25923 3160 25955
rect 3192 25923 3232 25955
rect 3264 25923 3304 25955
rect 3336 25923 3376 25955
rect 3408 25923 3448 25955
rect 3480 25923 3520 25955
rect 3552 25923 3592 25955
rect 3624 25923 3664 25955
rect 3696 25923 3736 25955
rect 3768 25923 3808 25955
rect 3840 25923 3880 25955
rect 3912 25923 3952 25955
rect 3984 25923 4024 25955
rect 4056 25923 4096 25955
rect 4128 25923 4168 25955
rect 4200 25923 4240 25955
rect 4272 25923 4312 25955
rect 4344 25923 4384 25955
rect 4416 25923 4456 25955
rect 4488 25923 4528 25955
rect 4560 25923 4600 25955
rect 4632 25923 4672 25955
rect 4704 25923 4744 25955
rect 4776 25923 4816 25955
rect 4848 25923 4888 25955
rect 4920 25923 4960 25955
rect 4992 25923 5032 25955
rect 5064 25923 5104 25955
rect 5136 25923 5176 25955
rect 5208 25923 5248 25955
rect 5280 25923 5320 25955
rect 5352 25923 5392 25955
rect 5424 25923 5464 25955
rect 5496 25923 5536 25955
rect 5568 25923 5608 25955
rect 5640 25923 5680 25955
rect 5712 25923 5752 25955
rect 5784 25923 5824 25955
rect 5856 25923 5896 25955
rect 5928 25923 5968 25955
rect 6000 25923 6040 25955
rect 6072 25923 6112 25955
rect 6144 25923 6184 25955
rect 6216 25923 6256 25955
rect 6288 25923 6328 25955
rect 6360 25923 6400 25955
rect 6432 25923 6472 25955
rect 6504 25923 6544 25955
rect 6576 25923 6616 25955
rect 6648 25923 6688 25955
rect 6720 25923 6760 25955
rect 6792 25923 6832 25955
rect 6864 25923 6904 25955
rect 6936 25923 6976 25955
rect 7008 25923 7048 25955
rect 7080 25923 7120 25955
rect 7152 25923 7192 25955
rect 7224 25923 7264 25955
rect 7296 25923 7336 25955
rect 7368 25923 7408 25955
rect 7440 25923 7480 25955
rect 7512 25923 7552 25955
rect 7584 25923 7624 25955
rect 7656 25923 7696 25955
rect 7728 25923 7768 25955
rect 7800 25923 7840 25955
rect 7872 25923 7912 25955
rect 7944 25923 7984 25955
rect 8016 25923 8056 25955
rect 8088 25923 8128 25955
rect 8160 25923 8200 25955
rect 8232 25923 8272 25955
rect 8304 25923 8344 25955
rect 8376 25923 8416 25955
rect 8448 25923 8488 25955
rect 8520 25923 8560 25955
rect 8592 25923 8632 25955
rect 8664 25923 8704 25955
rect 8736 25923 8776 25955
rect 8808 25923 8848 25955
rect 8880 25923 8920 25955
rect 8952 25923 8992 25955
rect 9024 25923 9064 25955
rect 9096 25923 9136 25955
rect 9168 25923 9208 25955
rect 9240 25923 9280 25955
rect 9312 25923 9352 25955
rect 9384 25923 9424 25955
rect 9456 25923 9496 25955
rect 9528 25923 9568 25955
rect 9600 25923 9640 25955
rect 9672 25923 9712 25955
rect 9744 25923 9784 25955
rect 9816 25923 9856 25955
rect 9888 25923 9928 25955
rect 9960 25923 10000 25955
rect 10032 25923 10072 25955
rect 10104 25923 10144 25955
rect 10176 25923 10216 25955
rect 10248 25923 10288 25955
rect 10320 25923 10360 25955
rect 10392 25923 10432 25955
rect 10464 25923 10504 25955
rect 10536 25923 10576 25955
rect 10608 25923 10648 25955
rect 10680 25923 10720 25955
rect 10752 25923 10792 25955
rect 10824 25923 10864 25955
rect 10896 25923 10936 25955
rect 10968 25923 11008 25955
rect 11040 25923 11080 25955
rect 11112 25923 11152 25955
rect 11184 25923 11224 25955
rect 11256 25923 11296 25955
rect 11328 25923 11368 25955
rect 11400 25923 11440 25955
rect 11472 25923 11512 25955
rect 11544 25923 11584 25955
rect 11616 25923 11656 25955
rect 11688 25923 11728 25955
rect 11760 25923 11800 25955
rect 11832 25923 11872 25955
rect 11904 25923 11944 25955
rect 11976 25923 12016 25955
rect 12048 25923 12088 25955
rect 12120 25923 12160 25955
rect 12192 25923 12232 25955
rect 12264 25923 12304 25955
rect 12336 25923 12376 25955
rect 12408 25923 12448 25955
rect 12480 25923 12520 25955
rect 12552 25923 12592 25955
rect 12624 25923 12664 25955
rect 12696 25923 12736 25955
rect 12768 25923 12808 25955
rect 12840 25923 12880 25955
rect 12912 25923 12952 25955
rect 12984 25923 13024 25955
rect 13056 25923 13096 25955
rect 13128 25923 13168 25955
rect 13200 25923 13240 25955
rect 13272 25923 13312 25955
rect 13344 25923 13384 25955
rect 13416 25923 13456 25955
rect 13488 25923 13528 25955
rect 13560 25923 13600 25955
rect 13632 25923 13672 25955
rect 13704 25923 13744 25955
rect 13776 25923 13816 25955
rect 13848 25923 13888 25955
rect 13920 25923 13960 25955
rect 13992 25923 14032 25955
rect 14064 25923 14104 25955
rect 14136 25923 14176 25955
rect 14208 25923 14248 25955
rect 14280 25923 14320 25955
rect 14352 25923 14392 25955
rect 14424 25923 14464 25955
rect 14496 25923 14536 25955
rect 14568 25923 14608 25955
rect 14640 25923 14680 25955
rect 14712 25923 14752 25955
rect 14784 25923 14824 25955
rect 14856 25923 14896 25955
rect 14928 25923 14968 25955
rect 15000 25923 15040 25955
rect 15072 25923 15112 25955
rect 15144 25923 15184 25955
rect 15216 25923 15256 25955
rect 15288 25923 15328 25955
rect 15360 25923 15400 25955
rect 15432 25923 15472 25955
rect 15504 25923 15544 25955
rect 15576 25923 15616 25955
rect 15648 25923 15688 25955
rect 15720 25923 15760 25955
rect 15792 25923 15832 25955
rect 15864 25923 15904 25955
rect 15936 25923 16000 25955
rect 0 25883 16000 25923
rect 0 25851 64 25883
rect 96 25851 136 25883
rect 168 25851 208 25883
rect 240 25851 280 25883
rect 312 25851 352 25883
rect 384 25851 424 25883
rect 456 25851 496 25883
rect 528 25851 568 25883
rect 600 25851 640 25883
rect 672 25851 712 25883
rect 744 25851 784 25883
rect 816 25851 856 25883
rect 888 25851 928 25883
rect 960 25851 1000 25883
rect 1032 25851 1072 25883
rect 1104 25851 1144 25883
rect 1176 25851 1216 25883
rect 1248 25851 1288 25883
rect 1320 25851 1360 25883
rect 1392 25851 1432 25883
rect 1464 25851 1504 25883
rect 1536 25851 1576 25883
rect 1608 25851 1648 25883
rect 1680 25851 1720 25883
rect 1752 25851 1792 25883
rect 1824 25851 1864 25883
rect 1896 25851 1936 25883
rect 1968 25851 2008 25883
rect 2040 25851 2080 25883
rect 2112 25851 2152 25883
rect 2184 25851 2224 25883
rect 2256 25851 2296 25883
rect 2328 25851 2368 25883
rect 2400 25851 2440 25883
rect 2472 25851 2512 25883
rect 2544 25851 2584 25883
rect 2616 25851 2656 25883
rect 2688 25851 2728 25883
rect 2760 25851 2800 25883
rect 2832 25851 2872 25883
rect 2904 25851 2944 25883
rect 2976 25851 3016 25883
rect 3048 25851 3088 25883
rect 3120 25851 3160 25883
rect 3192 25851 3232 25883
rect 3264 25851 3304 25883
rect 3336 25851 3376 25883
rect 3408 25851 3448 25883
rect 3480 25851 3520 25883
rect 3552 25851 3592 25883
rect 3624 25851 3664 25883
rect 3696 25851 3736 25883
rect 3768 25851 3808 25883
rect 3840 25851 3880 25883
rect 3912 25851 3952 25883
rect 3984 25851 4024 25883
rect 4056 25851 4096 25883
rect 4128 25851 4168 25883
rect 4200 25851 4240 25883
rect 4272 25851 4312 25883
rect 4344 25851 4384 25883
rect 4416 25851 4456 25883
rect 4488 25851 4528 25883
rect 4560 25851 4600 25883
rect 4632 25851 4672 25883
rect 4704 25851 4744 25883
rect 4776 25851 4816 25883
rect 4848 25851 4888 25883
rect 4920 25851 4960 25883
rect 4992 25851 5032 25883
rect 5064 25851 5104 25883
rect 5136 25851 5176 25883
rect 5208 25851 5248 25883
rect 5280 25851 5320 25883
rect 5352 25851 5392 25883
rect 5424 25851 5464 25883
rect 5496 25851 5536 25883
rect 5568 25851 5608 25883
rect 5640 25851 5680 25883
rect 5712 25851 5752 25883
rect 5784 25851 5824 25883
rect 5856 25851 5896 25883
rect 5928 25851 5968 25883
rect 6000 25851 6040 25883
rect 6072 25851 6112 25883
rect 6144 25851 6184 25883
rect 6216 25851 6256 25883
rect 6288 25851 6328 25883
rect 6360 25851 6400 25883
rect 6432 25851 6472 25883
rect 6504 25851 6544 25883
rect 6576 25851 6616 25883
rect 6648 25851 6688 25883
rect 6720 25851 6760 25883
rect 6792 25851 6832 25883
rect 6864 25851 6904 25883
rect 6936 25851 6976 25883
rect 7008 25851 7048 25883
rect 7080 25851 7120 25883
rect 7152 25851 7192 25883
rect 7224 25851 7264 25883
rect 7296 25851 7336 25883
rect 7368 25851 7408 25883
rect 7440 25851 7480 25883
rect 7512 25851 7552 25883
rect 7584 25851 7624 25883
rect 7656 25851 7696 25883
rect 7728 25851 7768 25883
rect 7800 25851 7840 25883
rect 7872 25851 7912 25883
rect 7944 25851 7984 25883
rect 8016 25851 8056 25883
rect 8088 25851 8128 25883
rect 8160 25851 8200 25883
rect 8232 25851 8272 25883
rect 8304 25851 8344 25883
rect 8376 25851 8416 25883
rect 8448 25851 8488 25883
rect 8520 25851 8560 25883
rect 8592 25851 8632 25883
rect 8664 25851 8704 25883
rect 8736 25851 8776 25883
rect 8808 25851 8848 25883
rect 8880 25851 8920 25883
rect 8952 25851 8992 25883
rect 9024 25851 9064 25883
rect 9096 25851 9136 25883
rect 9168 25851 9208 25883
rect 9240 25851 9280 25883
rect 9312 25851 9352 25883
rect 9384 25851 9424 25883
rect 9456 25851 9496 25883
rect 9528 25851 9568 25883
rect 9600 25851 9640 25883
rect 9672 25851 9712 25883
rect 9744 25851 9784 25883
rect 9816 25851 9856 25883
rect 9888 25851 9928 25883
rect 9960 25851 10000 25883
rect 10032 25851 10072 25883
rect 10104 25851 10144 25883
rect 10176 25851 10216 25883
rect 10248 25851 10288 25883
rect 10320 25851 10360 25883
rect 10392 25851 10432 25883
rect 10464 25851 10504 25883
rect 10536 25851 10576 25883
rect 10608 25851 10648 25883
rect 10680 25851 10720 25883
rect 10752 25851 10792 25883
rect 10824 25851 10864 25883
rect 10896 25851 10936 25883
rect 10968 25851 11008 25883
rect 11040 25851 11080 25883
rect 11112 25851 11152 25883
rect 11184 25851 11224 25883
rect 11256 25851 11296 25883
rect 11328 25851 11368 25883
rect 11400 25851 11440 25883
rect 11472 25851 11512 25883
rect 11544 25851 11584 25883
rect 11616 25851 11656 25883
rect 11688 25851 11728 25883
rect 11760 25851 11800 25883
rect 11832 25851 11872 25883
rect 11904 25851 11944 25883
rect 11976 25851 12016 25883
rect 12048 25851 12088 25883
rect 12120 25851 12160 25883
rect 12192 25851 12232 25883
rect 12264 25851 12304 25883
rect 12336 25851 12376 25883
rect 12408 25851 12448 25883
rect 12480 25851 12520 25883
rect 12552 25851 12592 25883
rect 12624 25851 12664 25883
rect 12696 25851 12736 25883
rect 12768 25851 12808 25883
rect 12840 25851 12880 25883
rect 12912 25851 12952 25883
rect 12984 25851 13024 25883
rect 13056 25851 13096 25883
rect 13128 25851 13168 25883
rect 13200 25851 13240 25883
rect 13272 25851 13312 25883
rect 13344 25851 13384 25883
rect 13416 25851 13456 25883
rect 13488 25851 13528 25883
rect 13560 25851 13600 25883
rect 13632 25851 13672 25883
rect 13704 25851 13744 25883
rect 13776 25851 13816 25883
rect 13848 25851 13888 25883
rect 13920 25851 13960 25883
rect 13992 25851 14032 25883
rect 14064 25851 14104 25883
rect 14136 25851 14176 25883
rect 14208 25851 14248 25883
rect 14280 25851 14320 25883
rect 14352 25851 14392 25883
rect 14424 25851 14464 25883
rect 14496 25851 14536 25883
rect 14568 25851 14608 25883
rect 14640 25851 14680 25883
rect 14712 25851 14752 25883
rect 14784 25851 14824 25883
rect 14856 25851 14896 25883
rect 14928 25851 14968 25883
rect 15000 25851 15040 25883
rect 15072 25851 15112 25883
rect 15144 25851 15184 25883
rect 15216 25851 15256 25883
rect 15288 25851 15328 25883
rect 15360 25851 15400 25883
rect 15432 25851 15472 25883
rect 15504 25851 15544 25883
rect 15576 25851 15616 25883
rect 15648 25851 15688 25883
rect 15720 25851 15760 25883
rect 15792 25851 15832 25883
rect 15864 25851 15904 25883
rect 15936 25851 16000 25883
rect 0 25811 16000 25851
rect 0 25779 64 25811
rect 96 25779 136 25811
rect 168 25779 208 25811
rect 240 25779 280 25811
rect 312 25779 352 25811
rect 384 25779 424 25811
rect 456 25779 496 25811
rect 528 25779 568 25811
rect 600 25779 640 25811
rect 672 25779 712 25811
rect 744 25779 784 25811
rect 816 25779 856 25811
rect 888 25779 928 25811
rect 960 25779 1000 25811
rect 1032 25779 1072 25811
rect 1104 25779 1144 25811
rect 1176 25779 1216 25811
rect 1248 25779 1288 25811
rect 1320 25779 1360 25811
rect 1392 25779 1432 25811
rect 1464 25779 1504 25811
rect 1536 25779 1576 25811
rect 1608 25779 1648 25811
rect 1680 25779 1720 25811
rect 1752 25779 1792 25811
rect 1824 25779 1864 25811
rect 1896 25779 1936 25811
rect 1968 25779 2008 25811
rect 2040 25779 2080 25811
rect 2112 25779 2152 25811
rect 2184 25779 2224 25811
rect 2256 25779 2296 25811
rect 2328 25779 2368 25811
rect 2400 25779 2440 25811
rect 2472 25779 2512 25811
rect 2544 25779 2584 25811
rect 2616 25779 2656 25811
rect 2688 25779 2728 25811
rect 2760 25779 2800 25811
rect 2832 25779 2872 25811
rect 2904 25779 2944 25811
rect 2976 25779 3016 25811
rect 3048 25779 3088 25811
rect 3120 25779 3160 25811
rect 3192 25779 3232 25811
rect 3264 25779 3304 25811
rect 3336 25779 3376 25811
rect 3408 25779 3448 25811
rect 3480 25779 3520 25811
rect 3552 25779 3592 25811
rect 3624 25779 3664 25811
rect 3696 25779 3736 25811
rect 3768 25779 3808 25811
rect 3840 25779 3880 25811
rect 3912 25779 3952 25811
rect 3984 25779 4024 25811
rect 4056 25779 4096 25811
rect 4128 25779 4168 25811
rect 4200 25779 4240 25811
rect 4272 25779 4312 25811
rect 4344 25779 4384 25811
rect 4416 25779 4456 25811
rect 4488 25779 4528 25811
rect 4560 25779 4600 25811
rect 4632 25779 4672 25811
rect 4704 25779 4744 25811
rect 4776 25779 4816 25811
rect 4848 25779 4888 25811
rect 4920 25779 4960 25811
rect 4992 25779 5032 25811
rect 5064 25779 5104 25811
rect 5136 25779 5176 25811
rect 5208 25779 5248 25811
rect 5280 25779 5320 25811
rect 5352 25779 5392 25811
rect 5424 25779 5464 25811
rect 5496 25779 5536 25811
rect 5568 25779 5608 25811
rect 5640 25779 5680 25811
rect 5712 25779 5752 25811
rect 5784 25779 5824 25811
rect 5856 25779 5896 25811
rect 5928 25779 5968 25811
rect 6000 25779 6040 25811
rect 6072 25779 6112 25811
rect 6144 25779 6184 25811
rect 6216 25779 6256 25811
rect 6288 25779 6328 25811
rect 6360 25779 6400 25811
rect 6432 25779 6472 25811
rect 6504 25779 6544 25811
rect 6576 25779 6616 25811
rect 6648 25779 6688 25811
rect 6720 25779 6760 25811
rect 6792 25779 6832 25811
rect 6864 25779 6904 25811
rect 6936 25779 6976 25811
rect 7008 25779 7048 25811
rect 7080 25779 7120 25811
rect 7152 25779 7192 25811
rect 7224 25779 7264 25811
rect 7296 25779 7336 25811
rect 7368 25779 7408 25811
rect 7440 25779 7480 25811
rect 7512 25779 7552 25811
rect 7584 25779 7624 25811
rect 7656 25779 7696 25811
rect 7728 25779 7768 25811
rect 7800 25779 7840 25811
rect 7872 25779 7912 25811
rect 7944 25779 7984 25811
rect 8016 25779 8056 25811
rect 8088 25779 8128 25811
rect 8160 25779 8200 25811
rect 8232 25779 8272 25811
rect 8304 25779 8344 25811
rect 8376 25779 8416 25811
rect 8448 25779 8488 25811
rect 8520 25779 8560 25811
rect 8592 25779 8632 25811
rect 8664 25779 8704 25811
rect 8736 25779 8776 25811
rect 8808 25779 8848 25811
rect 8880 25779 8920 25811
rect 8952 25779 8992 25811
rect 9024 25779 9064 25811
rect 9096 25779 9136 25811
rect 9168 25779 9208 25811
rect 9240 25779 9280 25811
rect 9312 25779 9352 25811
rect 9384 25779 9424 25811
rect 9456 25779 9496 25811
rect 9528 25779 9568 25811
rect 9600 25779 9640 25811
rect 9672 25779 9712 25811
rect 9744 25779 9784 25811
rect 9816 25779 9856 25811
rect 9888 25779 9928 25811
rect 9960 25779 10000 25811
rect 10032 25779 10072 25811
rect 10104 25779 10144 25811
rect 10176 25779 10216 25811
rect 10248 25779 10288 25811
rect 10320 25779 10360 25811
rect 10392 25779 10432 25811
rect 10464 25779 10504 25811
rect 10536 25779 10576 25811
rect 10608 25779 10648 25811
rect 10680 25779 10720 25811
rect 10752 25779 10792 25811
rect 10824 25779 10864 25811
rect 10896 25779 10936 25811
rect 10968 25779 11008 25811
rect 11040 25779 11080 25811
rect 11112 25779 11152 25811
rect 11184 25779 11224 25811
rect 11256 25779 11296 25811
rect 11328 25779 11368 25811
rect 11400 25779 11440 25811
rect 11472 25779 11512 25811
rect 11544 25779 11584 25811
rect 11616 25779 11656 25811
rect 11688 25779 11728 25811
rect 11760 25779 11800 25811
rect 11832 25779 11872 25811
rect 11904 25779 11944 25811
rect 11976 25779 12016 25811
rect 12048 25779 12088 25811
rect 12120 25779 12160 25811
rect 12192 25779 12232 25811
rect 12264 25779 12304 25811
rect 12336 25779 12376 25811
rect 12408 25779 12448 25811
rect 12480 25779 12520 25811
rect 12552 25779 12592 25811
rect 12624 25779 12664 25811
rect 12696 25779 12736 25811
rect 12768 25779 12808 25811
rect 12840 25779 12880 25811
rect 12912 25779 12952 25811
rect 12984 25779 13024 25811
rect 13056 25779 13096 25811
rect 13128 25779 13168 25811
rect 13200 25779 13240 25811
rect 13272 25779 13312 25811
rect 13344 25779 13384 25811
rect 13416 25779 13456 25811
rect 13488 25779 13528 25811
rect 13560 25779 13600 25811
rect 13632 25779 13672 25811
rect 13704 25779 13744 25811
rect 13776 25779 13816 25811
rect 13848 25779 13888 25811
rect 13920 25779 13960 25811
rect 13992 25779 14032 25811
rect 14064 25779 14104 25811
rect 14136 25779 14176 25811
rect 14208 25779 14248 25811
rect 14280 25779 14320 25811
rect 14352 25779 14392 25811
rect 14424 25779 14464 25811
rect 14496 25779 14536 25811
rect 14568 25779 14608 25811
rect 14640 25779 14680 25811
rect 14712 25779 14752 25811
rect 14784 25779 14824 25811
rect 14856 25779 14896 25811
rect 14928 25779 14968 25811
rect 15000 25779 15040 25811
rect 15072 25779 15112 25811
rect 15144 25779 15184 25811
rect 15216 25779 15256 25811
rect 15288 25779 15328 25811
rect 15360 25779 15400 25811
rect 15432 25779 15472 25811
rect 15504 25779 15544 25811
rect 15576 25779 15616 25811
rect 15648 25779 15688 25811
rect 15720 25779 15760 25811
rect 15792 25779 15832 25811
rect 15864 25779 15904 25811
rect 15936 25779 16000 25811
rect 0 25739 16000 25779
rect 0 25707 64 25739
rect 96 25707 136 25739
rect 168 25707 208 25739
rect 240 25707 280 25739
rect 312 25707 352 25739
rect 384 25707 424 25739
rect 456 25707 496 25739
rect 528 25707 568 25739
rect 600 25707 640 25739
rect 672 25707 712 25739
rect 744 25707 784 25739
rect 816 25707 856 25739
rect 888 25707 928 25739
rect 960 25707 1000 25739
rect 1032 25707 1072 25739
rect 1104 25707 1144 25739
rect 1176 25707 1216 25739
rect 1248 25707 1288 25739
rect 1320 25707 1360 25739
rect 1392 25707 1432 25739
rect 1464 25707 1504 25739
rect 1536 25707 1576 25739
rect 1608 25707 1648 25739
rect 1680 25707 1720 25739
rect 1752 25707 1792 25739
rect 1824 25707 1864 25739
rect 1896 25707 1936 25739
rect 1968 25707 2008 25739
rect 2040 25707 2080 25739
rect 2112 25707 2152 25739
rect 2184 25707 2224 25739
rect 2256 25707 2296 25739
rect 2328 25707 2368 25739
rect 2400 25707 2440 25739
rect 2472 25707 2512 25739
rect 2544 25707 2584 25739
rect 2616 25707 2656 25739
rect 2688 25707 2728 25739
rect 2760 25707 2800 25739
rect 2832 25707 2872 25739
rect 2904 25707 2944 25739
rect 2976 25707 3016 25739
rect 3048 25707 3088 25739
rect 3120 25707 3160 25739
rect 3192 25707 3232 25739
rect 3264 25707 3304 25739
rect 3336 25707 3376 25739
rect 3408 25707 3448 25739
rect 3480 25707 3520 25739
rect 3552 25707 3592 25739
rect 3624 25707 3664 25739
rect 3696 25707 3736 25739
rect 3768 25707 3808 25739
rect 3840 25707 3880 25739
rect 3912 25707 3952 25739
rect 3984 25707 4024 25739
rect 4056 25707 4096 25739
rect 4128 25707 4168 25739
rect 4200 25707 4240 25739
rect 4272 25707 4312 25739
rect 4344 25707 4384 25739
rect 4416 25707 4456 25739
rect 4488 25707 4528 25739
rect 4560 25707 4600 25739
rect 4632 25707 4672 25739
rect 4704 25707 4744 25739
rect 4776 25707 4816 25739
rect 4848 25707 4888 25739
rect 4920 25707 4960 25739
rect 4992 25707 5032 25739
rect 5064 25707 5104 25739
rect 5136 25707 5176 25739
rect 5208 25707 5248 25739
rect 5280 25707 5320 25739
rect 5352 25707 5392 25739
rect 5424 25707 5464 25739
rect 5496 25707 5536 25739
rect 5568 25707 5608 25739
rect 5640 25707 5680 25739
rect 5712 25707 5752 25739
rect 5784 25707 5824 25739
rect 5856 25707 5896 25739
rect 5928 25707 5968 25739
rect 6000 25707 6040 25739
rect 6072 25707 6112 25739
rect 6144 25707 6184 25739
rect 6216 25707 6256 25739
rect 6288 25707 6328 25739
rect 6360 25707 6400 25739
rect 6432 25707 6472 25739
rect 6504 25707 6544 25739
rect 6576 25707 6616 25739
rect 6648 25707 6688 25739
rect 6720 25707 6760 25739
rect 6792 25707 6832 25739
rect 6864 25707 6904 25739
rect 6936 25707 6976 25739
rect 7008 25707 7048 25739
rect 7080 25707 7120 25739
rect 7152 25707 7192 25739
rect 7224 25707 7264 25739
rect 7296 25707 7336 25739
rect 7368 25707 7408 25739
rect 7440 25707 7480 25739
rect 7512 25707 7552 25739
rect 7584 25707 7624 25739
rect 7656 25707 7696 25739
rect 7728 25707 7768 25739
rect 7800 25707 7840 25739
rect 7872 25707 7912 25739
rect 7944 25707 7984 25739
rect 8016 25707 8056 25739
rect 8088 25707 8128 25739
rect 8160 25707 8200 25739
rect 8232 25707 8272 25739
rect 8304 25707 8344 25739
rect 8376 25707 8416 25739
rect 8448 25707 8488 25739
rect 8520 25707 8560 25739
rect 8592 25707 8632 25739
rect 8664 25707 8704 25739
rect 8736 25707 8776 25739
rect 8808 25707 8848 25739
rect 8880 25707 8920 25739
rect 8952 25707 8992 25739
rect 9024 25707 9064 25739
rect 9096 25707 9136 25739
rect 9168 25707 9208 25739
rect 9240 25707 9280 25739
rect 9312 25707 9352 25739
rect 9384 25707 9424 25739
rect 9456 25707 9496 25739
rect 9528 25707 9568 25739
rect 9600 25707 9640 25739
rect 9672 25707 9712 25739
rect 9744 25707 9784 25739
rect 9816 25707 9856 25739
rect 9888 25707 9928 25739
rect 9960 25707 10000 25739
rect 10032 25707 10072 25739
rect 10104 25707 10144 25739
rect 10176 25707 10216 25739
rect 10248 25707 10288 25739
rect 10320 25707 10360 25739
rect 10392 25707 10432 25739
rect 10464 25707 10504 25739
rect 10536 25707 10576 25739
rect 10608 25707 10648 25739
rect 10680 25707 10720 25739
rect 10752 25707 10792 25739
rect 10824 25707 10864 25739
rect 10896 25707 10936 25739
rect 10968 25707 11008 25739
rect 11040 25707 11080 25739
rect 11112 25707 11152 25739
rect 11184 25707 11224 25739
rect 11256 25707 11296 25739
rect 11328 25707 11368 25739
rect 11400 25707 11440 25739
rect 11472 25707 11512 25739
rect 11544 25707 11584 25739
rect 11616 25707 11656 25739
rect 11688 25707 11728 25739
rect 11760 25707 11800 25739
rect 11832 25707 11872 25739
rect 11904 25707 11944 25739
rect 11976 25707 12016 25739
rect 12048 25707 12088 25739
rect 12120 25707 12160 25739
rect 12192 25707 12232 25739
rect 12264 25707 12304 25739
rect 12336 25707 12376 25739
rect 12408 25707 12448 25739
rect 12480 25707 12520 25739
rect 12552 25707 12592 25739
rect 12624 25707 12664 25739
rect 12696 25707 12736 25739
rect 12768 25707 12808 25739
rect 12840 25707 12880 25739
rect 12912 25707 12952 25739
rect 12984 25707 13024 25739
rect 13056 25707 13096 25739
rect 13128 25707 13168 25739
rect 13200 25707 13240 25739
rect 13272 25707 13312 25739
rect 13344 25707 13384 25739
rect 13416 25707 13456 25739
rect 13488 25707 13528 25739
rect 13560 25707 13600 25739
rect 13632 25707 13672 25739
rect 13704 25707 13744 25739
rect 13776 25707 13816 25739
rect 13848 25707 13888 25739
rect 13920 25707 13960 25739
rect 13992 25707 14032 25739
rect 14064 25707 14104 25739
rect 14136 25707 14176 25739
rect 14208 25707 14248 25739
rect 14280 25707 14320 25739
rect 14352 25707 14392 25739
rect 14424 25707 14464 25739
rect 14496 25707 14536 25739
rect 14568 25707 14608 25739
rect 14640 25707 14680 25739
rect 14712 25707 14752 25739
rect 14784 25707 14824 25739
rect 14856 25707 14896 25739
rect 14928 25707 14968 25739
rect 15000 25707 15040 25739
rect 15072 25707 15112 25739
rect 15144 25707 15184 25739
rect 15216 25707 15256 25739
rect 15288 25707 15328 25739
rect 15360 25707 15400 25739
rect 15432 25707 15472 25739
rect 15504 25707 15544 25739
rect 15576 25707 15616 25739
rect 15648 25707 15688 25739
rect 15720 25707 15760 25739
rect 15792 25707 15832 25739
rect 15864 25707 15904 25739
rect 15936 25707 16000 25739
rect 0 25667 16000 25707
rect 0 25635 64 25667
rect 96 25635 136 25667
rect 168 25635 208 25667
rect 240 25635 280 25667
rect 312 25635 352 25667
rect 384 25635 424 25667
rect 456 25635 496 25667
rect 528 25635 568 25667
rect 600 25635 640 25667
rect 672 25635 712 25667
rect 744 25635 784 25667
rect 816 25635 856 25667
rect 888 25635 928 25667
rect 960 25635 1000 25667
rect 1032 25635 1072 25667
rect 1104 25635 1144 25667
rect 1176 25635 1216 25667
rect 1248 25635 1288 25667
rect 1320 25635 1360 25667
rect 1392 25635 1432 25667
rect 1464 25635 1504 25667
rect 1536 25635 1576 25667
rect 1608 25635 1648 25667
rect 1680 25635 1720 25667
rect 1752 25635 1792 25667
rect 1824 25635 1864 25667
rect 1896 25635 1936 25667
rect 1968 25635 2008 25667
rect 2040 25635 2080 25667
rect 2112 25635 2152 25667
rect 2184 25635 2224 25667
rect 2256 25635 2296 25667
rect 2328 25635 2368 25667
rect 2400 25635 2440 25667
rect 2472 25635 2512 25667
rect 2544 25635 2584 25667
rect 2616 25635 2656 25667
rect 2688 25635 2728 25667
rect 2760 25635 2800 25667
rect 2832 25635 2872 25667
rect 2904 25635 2944 25667
rect 2976 25635 3016 25667
rect 3048 25635 3088 25667
rect 3120 25635 3160 25667
rect 3192 25635 3232 25667
rect 3264 25635 3304 25667
rect 3336 25635 3376 25667
rect 3408 25635 3448 25667
rect 3480 25635 3520 25667
rect 3552 25635 3592 25667
rect 3624 25635 3664 25667
rect 3696 25635 3736 25667
rect 3768 25635 3808 25667
rect 3840 25635 3880 25667
rect 3912 25635 3952 25667
rect 3984 25635 4024 25667
rect 4056 25635 4096 25667
rect 4128 25635 4168 25667
rect 4200 25635 4240 25667
rect 4272 25635 4312 25667
rect 4344 25635 4384 25667
rect 4416 25635 4456 25667
rect 4488 25635 4528 25667
rect 4560 25635 4600 25667
rect 4632 25635 4672 25667
rect 4704 25635 4744 25667
rect 4776 25635 4816 25667
rect 4848 25635 4888 25667
rect 4920 25635 4960 25667
rect 4992 25635 5032 25667
rect 5064 25635 5104 25667
rect 5136 25635 5176 25667
rect 5208 25635 5248 25667
rect 5280 25635 5320 25667
rect 5352 25635 5392 25667
rect 5424 25635 5464 25667
rect 5496 25635 5536 25667
rect 5568 25635 5608 25667
rect 5640 25635 5680 25667
rect 5712 25635 5752 25667
rect 5784 25635 5824 25667
rect 5856 25635 5896 25667
rect 5928 25635 5968 25667
rect 6000 25635 6040 25667
rect 6072 25635 6112 25667
rect 6144 25635 6184 25667
rect 6216 25635 6256 25667
rect 6288 25635 6328 25667
rect 6360 25635 6400 25667
rect 6432 25635 6472 25667
rect 6504 25635 6544 25667
rect 6576 25635 6616 25667
rect 6648 25635 6688 25667
rect 6720 25635 6760 25667
rect 6792 25635 6832 25667
rect 6864 25635 6904 25667
rect 6936 25635 6976 25667
rect 7008 25635 7048 25667
rect 7080 25635 7120 25667
rect 7152 25635 7192 25667
rect 7224 25635 7264 25667
rect 7296 25635 7336 25667
rect 7368 25635 7408 25667
rect 7440 25635 7480 25667
rect 7512 25635 7552 25667
rect 7584 25635 7624 25667
rect 7656 25635 7696 25667
rect 7728 25635 7768 25667
rect 7800 25635 7840 25667
rect 7872 25635 7912 25667
rect 7944 25635 7984 25667
rect 8016 25635 8056 25667
rect 8088 25635 8128 25667
rect 8160 25635 8200 25667
rect 8232 25635 8272 25667
rect 8304 25635 8344 25667
rect 8376 25635 8416 25667
rect 8448 25635 8488 25667
rect 8520 25635 8560 25667
rect 8592 25635 8632 25667
rect 8664 25635 8704 25667
rect 8736 25635 8776 25667
rect 8808 25635 8848 25667
rect 8880 25635 8920 25667
rect 8952 25635 8992 25667
rect 9024 25635 9064 25667
rect 9096 25635 9136 25667
rect 9168 25635 9208 25667
rect 9240 25635 9280 25667
rect 9312 25635 9352 25667
rect 9384 25635 9424 25667
rect 9456 25635 9496 25667
rect 9528 25635 9568 25667
rect 9600 25635 9640 25667
rect 9672 25635 9712 25667
rect 9744 25635 9784 25667
rect 9816 25635 9856 25667
rect 9888 25635 9928 25667
rect 9960 25635 10000 25667
rect 10032 25635 10072 25667
rect 10104 25635 10144 25667
rect 10176 25635 10216 25667
rect 10248 25635 10288 25667
rect 10320 25635 10360 25667
rect 10392 25635 10432 25667
rect 10464 25635 10504 25667
rect 10536 25635 10576 25667
rect 10608 25635 10648 25667
rect 10680 25635 10720 25667
rect 10752 25635 10792 25667
rect 10824 25635 10864 25667
rect 10896 25635 10936 25667
rect 10968 25635 11008 25667
rect 11040 25635 11080 25667
rect 11112 25635 11152 25667
rect 11184 25635 11224 25667
rect 11256 25635 11296 25667
rect 11328 25635 11368 25667
rect 11400 25635 11440 25667
rect 11472 25635 11512 25667
rect 11544 25635 11584 25667
rect 11616 25635 11656 25667
rect 11688 25635 11728 25667
rect 11760 25635 11800 25667
rect 11832 25635 11872 25667
rect 11904 25635 11944 25667
rect 11976 25635 12016 25667
rect 12048 25635 12088 25667
rect 12120 25635 12160 25667
rect 12192 25635 12232 25667
rect 12264 25635 12304 25667
rect 12336 25635 12376 25667
rect 12408 25635 12448 25667
rect 12480 25635 12520 25667
rect 12552 25635 12592 25667
rect 12624 25635 12664 25667
rect 12696 25635 12736 25667
rect 12768 25635 12808 25667
rect 12840 25635 12880 25667
rect 12912 25635 12952 25667
rect 12984 25635 13024 25667
rect 13056 25635 13096 25667
rect 13128 25635 13168 25667
rect 13200 25635 13240 25667
rect 13272 25635 13312 25667
rect 13344 25635 13384 25667
rect 13416 25635 13456 25667
rect 13488 25635 13528 25667
rect 13560 25635 13600 25667
rect 13632 25635 13672 25667
rect 13704 25635 13744 25667
rect 13776 25635 13816 25667
rect 13848 25635 13888 25667
rect 13920 25635 13960 25667
rect 13992 25635 14032 25667
rect 14064 25635 14104 25667
rect 14136 25635 14176 25667
rect 14208 25635 14248 25667
rect 14280 25635 14320 25667
rect 14352 25635 14392 25667
rect 14424 25635 14464 25667
rect 14496 25635 14536 25667
rect 14568 25635 14608 25667
rect 14640 25635 14680 25667
rect 14712 25635 14752 25667
rect 14784 25635 14824 25667
rect 14856 25635 14896 25667
rect 14928 25635 14968 25667
rect 15000 25635 15040 25667
rect 15072 25635 15112 25667
rect 15144 25635 15184 25667
rect 15216 25635 15256 25667
rect 15288 25635 15328 25667
rect 15360 25635 15400 25667
rect 15432 25635 15472 25667
rect 15504 25635 15544 25667
rect 15576 25635 15616 25667
rect 15648 25635 15688 25667
rect 15720 25635 15760 25667
rect 15792 25635 15832 25667
rect 15864 25635 15904 25667
rect 15936 25635 16000 25667
rect 0 25595 16000 25635
rect 0 25563 64 25595
rect 96 25563 136 25595
rect 168 25563 208 25595
rect 240 25563 280 25595
rect 312 25563 352 25595
rect 384 25563 424 25595
rect 456 25563 496 25595
rect 528 25563 568 25595
rect 600 25563 640 25595
rect 672 25563 712 25595
rect 744 25563 784 25595
rect 816 25563 856 25595
rect 888 25563 928 25595
rect 960 25563 1000 25595
rect 1032 25563 1072 25595
rect 1104 25563 1144 25595
rect 1176 25563 1216 25595
rect 1248 25563 1288 25595
rect 1320 25563 1360 25595
rect 1392 25563 1432 25595
rect 1464 25563 1504 25595
rect 1536 25563 1576 25595
rect 1608 25563 1648 25595
rect 1680 25563 1720 25595
rect 1752 25563 1792 25595
rect 1824 25563 1864 25595
rect 1896 25563 1936 25595
rect 1968 25563 2008 25595
rect 2040 25563 2080 25595
rect 2112 25563 2152 25595
rect 2184 25563 2224 25595
rect 2256 25563 2296 25595
rect 2328 25563 2368 25595
rect 2400 25563 2440 25595
rect 2472 25563 2512 25595
rect 2544 25563 2584 25595
rect 2616 25563 2656 25595
rect 2688 25563 2728 25595
rect 2760 25563 2800 25595
rect 2832 25563 2872 25595
rect 2904 25563 2944 25595
rect 2976 25563 3016 25595
rect 3048 25563 3088 25595
rect 3120 25563 3160 25595
rect 3192 25563 3232 25595
rect 3264 25563 3304 25595
rect 3336 25563 3376 25595
rect 3408 25563 3448 25595
rect 3480 25563 3520 25595
rect 3552 25563 3592 25595
rect 3624 25563 3664 25595
rect 3696 25563 3736 25595
rect 3768 25563 3808 25595
rect 3840 25563 3880 25595
rect 3912 25563 3952 25595
rect 3984 25563 4024 25595
rect 4056 25563 4096 25595
rect 4128 25563 4168 25595
rect 4200 25563 4240 25595
rect 4272 25563 4312 25595
rect 4344 25563 4384 25595
rect 4416 25563 4456 25595
rect 4488 25563 4528 25595
rect 4560 25563 4600 25595
rect 4632 25563 4672 25595
rect 4704 25563 4744 25595
rect 4776 25563 4816 25595
rect 4848 25563 4888 25595
rect 4920 25563 4960 25595
rect 4992 25563 5032 25595
rect 5064 25563 5104 25595
rect 5136 25563 5176 25595
rect 5208 25563 5248 25595
rect 5280 25563 5320 25595
rect 5352 25563 5392 25595
rect 5424 25563 5464 25595
rect 5496 25563 5536 25595
rect 5568 25563 5608 25595
rect 5640 25563 5680 25595
rect 5712 25563 5752 25595
rect 5784 25563 5824 25595
rect 5856 25563 5896 25595
rect 5928 25563 5968 25595
rect 6000 25563 6040 25595
rect 6072 25563 6112 25595
rect 6144 25563 6184 25595
rect 6216 25563 6256 25595
rect 6288 25563 6328 25595
rect 6360 25563 6400 25595
rect 6432 25563 6472 25595
rect 6504 25563 6544 25595
rect 6576 25563 6616 25595
rect 6648 25563 6688 25595
rect 6720 25563 6760 25595
rect 6792 25563 6832 25595
rect 6864 25563 6904 25595
rect 6936 25563 6976 25595
rect 7008 25563 7048 25595
rect 7080 25563 7120 25595
rect 7152 25563 7192 25595
rect 7224 25563 7264 25595
rect 7296 25563 7336 25595
rect 7368 25563 7408 25595
rect 7440 25563 7480 25595
rect 7512 25563 7552 25595
rect 7584 25563 7624 25595
rect 7656 25563 7696 25595
rect 7728 25563 7768 25595
rect 7800 25563 7840 25595
rect 7872 25563 7912 25595
rect 7944 25563 7984 25595
rect 8016 25563 8056 25595
rect 8088 25563 8128 25595
rect 8160 25563 8200 25595
rect 8232 25563 8272 25595
rect 8304 25563 8344 25595
rect 8376 25563 8416 25595
rect 8448 25563 8488 25595
rect 8520 25563 8560 25595
rect 8592 25563 8632 25595
rect 8664 25563 8704 25595
rect 8736 25563 8776 25595
rect 8808 25563 8848 25595
rect 8880 25563 8920 25595
rect 8952 25563 8992 25595
rect 9024 25563 9064 25595
rect 9096 25563 9136 25595
rect 9168 25563 9208 25595
rect 9240 25563 9280 25595
rect 9312 25563 9352 25595
rect 9384 25563 9424 25595
rect 9456 25563 9496 25595
rect 9528 25563 9568 25595
rect 9600 25563 9640 25595
rect 9672 25563 9712 25595
rect 9744 25563 9784 25595
rect 9816 25563 9856 25595
rect 9888 25563 9928 25595
rect 9960 25563 10000 25595
rect 10032 25563 10072 25595
rect 10104 25563 10144 25595
rect 10176 25563 10216 25595
rect 10248 25563 10288 25595
rect 10320 25563 10360 25595
rect 10392 25563 10432 25595
rect 10464 25563 10504 25595
rect 10536 25563 10576 25595
rect 10608 25563 10648 25595
rect 10680 25563 10720 25595
rect 10752 25563 10792 25595
rect 10824 25563 10864 25595
rect 10896 25563 10936 25595
rect 10968 25563 11008 25595
rect 11040 25563 11080 25595
rect 11112 25563 11152 25595
rect 11184 25563 11224 25595
rect 11256 25563 11296 25595
rect 11328 25563 11368 25595
rect 11400 25563 11440 25595
rect 11472 25563 11512 25595
rect 11544 25563 11584 25595
rect 11616 25563 11656 25595
rect 11688 25563 11728 25595
rect 11760 25563 11800 25595
rect 11832 25563 11872 25595
rect 11904 25563 11944 25595
rect 11976 25563 12016 25595
rect 12048 25563 12088 25595
rect 12120 25563 12160 25595
rect 12192 25563 12232 25595
rect 12264 25563 12304 25595
rect 12336 25563 12376 25595
rect 12408 25563 12448 25595
rect 12480 25563 12520 25595
rect 12552 25563 12592 25595
rect 12624 25563 12664 25595
rect 12696 25563 12736 25595
rect 12768 25563 12808 25595
rect 12840 25563 12880 25595
rect 12912 25563 12952 25595
rect 12984 25563 13024 25595
rect 13056 25563 13096 25595
rect 13128 25563 13168 25595
rect 13200 25563 13240 25595
rect 13272 25563 13312 25595
rect 13344 25563 13384 25595
rect 13416 25563 13456 25595
rect 13488 25563 13528 25595
rect 13560 25563 13600 25595
rect 13632 25563 13672 25595
rect 13704 25563 13744 25595
rect 13776 25563 13816 25595
rect 13848 25563 13888 25595
rect 13920 25563 13960 25595
rect 13992 25563 14032 25595
rect 14064 25563 14104 25595
rect 14136 25563 14176 25595
rect 14208 25563 14248 25595
rect 14280 25563 14320 25595
rect 14352 25563 14392 25595
rect 14424 25563 14464 25595
rect 14496 25563 14536 25595
rect 14568 25563 14608 25595
rect 14640 25563 14680 25595
rect 14712 25563 14752 25595
rect 14784 25563 14824 25595
rect 14856 25563 14896 25595
rect 14928 25563 14968 25595
rect 15000 25563 15040 25595
rect 15072 25563 15112 25595
rect 15144 25563 15184 25595
rect 15216 25563 15256 25595
rect 15288 25563 15328 25595
rect 15360 25563 15400 25595
rect 15432 25563 15472 25595
rect 15504 25563 15544 25595
rect 15576 25563 15616 25595
rect 15648 25563 15688 25595
rect 15720 25563 15760 25595
rect 15792 25563 15832 25595
rect 15864 25563 15904 25595
rect 15936 25563 16000 25595
rect 0 25523 16000 25563
rect 0 25491 64 25523
rect 96 25491 136 25523
rect 168 25491 208 25523
rect 240 25491 280 25523
rect 312 25491 352 25523
rect 384 25491 424 25523
rect 456 25491 496 25523
rect 528 25491 568 25523
rect 600 25491 640 25523
rect 672 25491 712 25523
rect 744 25491 784 25523
rect 816 25491 856 25523
rect 888 25491 928 25523
rect 960 25491 1000 25523
rect 1032 25491 1072 25523
rect 1104 25491 1144 25523
rect 1176 25491 1216 25523
rect 1248 25491 1288 25523
rect 1320 25491 1360 25523
rect 1392 25491 1432 25523
rect 1464 25491 1504 25523
rect 1536 25491 1576 25523
rect 1608 25491 1648 25523
rect 1680 25491 1720 25523
rect 1752 25491 1792 25523
rect 1824 25491 1864 25523
rect 1896 25491 1936 25523
rect 1968 25491 2008 25523
rect 2040 25491 2080 25523
rect 2112 25491 2152 25523
rect 2184 25491 2224 25523
rect 2256 25491 2296 25523
rect 2328 25491 2368 25523
rect 2400 25491 2440 25523
rect 2472 25491 2512 25523
rect 2544 25491 2584 25523
rect 2616 25491 2656 25523
rect 2688 25491 2728 25523
rect 2760 25491 2800 25523
rect 2832 25491 2872 25523
rect 2904 25491 2944 25523
rect 2976 25491 3016 25523
rect 3048 25491 3088 25523
rect 3120 25491 3160 25523
rect 3192 25491 3232 25523
rect 3264 25491 3304 25523
rect 3336 25491 3376 25523
rect 3408 25491 3448 25523
rect 3480 25491 3520 25523
rect 3552 25491 3592 25523
rect 3624 25491 3664 25523
rect 3696 25491 3736 25523
rect 3768 25491 3808 25523
rect 3840 25491 3880 25523
rect 3912 25491 3952 25523
rect 3984 25491 4024 25523
rect 4056 25491 4096 25523
rect 4128 25491 4168 25523
rect 4200 25491 4240 25523
rect 4272 25491 4312 25523
rect 4344 25491 4384 25523
rect 4416 25491 4456 25523
rect 4488 25491 4528 25523
rect 4560 25491 4600 25523
rect 4632 25491 4672 25523
rect 4704 25491 4744 25523
rect 4776 25491 4816 25523
rect 4848 25491 4888 25523
rect 4920 25491 4960 25523
rect 4992 25491 5032 25523
rect 5064 25491 5104 25523
rect 5136 25491 5176 25523
rect 5208 25491 5248 25523
rect 5280 25491 5320 25523
rect 5352 25491 5392 25523
rect 5424 25491 5464 25523
rect 5496 25491 5536 25523
rect 5568 25491 5608 25523
rect 5640 25491 5680 25523
rect 5712 25491 5752 25523
rect 5784 25491 5824 25523
rect 5856 25491 5896 25523
rect 5928 25491 5968 25523
rect 6000 25491 6040 25523
rect 6072 25491 6112 25523
rect 6144 25491 6184 25523
rect 6216 25491 6256 25523
rect 6288 25491 6328 25523
rect 6360 25491 6400 25523
rect 6432 25491 6472 25523
rect 6504 25491 6544 25523
rect 6576 25491 6616 25523
rect 6648 25491 6688 25523
rect 6720 25491 6760 25523
rect 6792 25491 6832 25523
rect 6864 25491 6904 25523
rect 6936 25491 6976 25523
rect 7008 25491 7048 25523
rect 7080 25491 7120 25523
rect 7152 25491 7192 25523
rect 7224 25491 7264 25523
rect 7296 25491 7336 25523
rect 7368 25491 7408 25523
rect 7440 25491 7480 25523
rect 7512 25491 7552 25523
rect 7584 25491 7624 25523
rect 7656 25491 7696 25523
rect 7728 25491 7768 25523
rect 7800 25491 7840 25523
rect 7872 25491 7912 25523
rect 7944 25491 7984 25523
rect 8016 25491 8056 25523
rect 8088 25491 8128 25523
rect 8160 25491 8200 25523
rect 8232 25491 8272 25523
rect 8304 25491 8344 25523
rect 8376 25491 8416 25523
rect 8448 25491 8488 25523
rect 8520 25491 8560 25523
rect 8592 25491 8632 25523
rect 8664 25491 8704 25523
rect 8736 25491 8776 25523
rect 8808 25491 8848 25523
rect 8880 25491 8920 25523
rect 8952 25491 8992 25523
rect 9024 25491 9064 25523
rect 9096 25491 9136 25523
rect 9168 25491 9208 25523
rect 9240 25491 9280 25523
rect 9312 25491 9352 25523
rect 9384 25491 9424 25523
rect 9456 25491 9496 25523
rect 9528 25491 9568 25523
rect 9600 25491 9640 25523
rect 9672 25491 9712 25523
rect 9744 25491 9784 25523
rect 9816 25491 9856 25523
rect 9888 25491 9928 25523
rect 9960 25491 10000 25523
rect 10032 25491 10072 25523
rect 10104 25491 10144 25523
rect 10176 25491 10216 25523
rect 10248 25491 10288 25523
rect 10320 25491 10360 25523
rect 10392 25491 10432 25523
rect 10464 25491 10504 25523
rect 10536 25491 10576 25523
rect 10608 25491 10648 25523
rect 10680 25491 10720 25523
rect 10752 25491 10792 25523
rect 10824 25491 10864 25523
rect 10896 25491 10936 25523
rect 10968 25491 11008 25523
rect 11040 25491 11080 25523
rect 11112 25491 11152 25523
rect 11184 25491 11224 25523
rect 11256 25491 11296 25523
rect 11328 25491 11368 25523
rect 11400 25491 11440 25523
rect 11472 25491 11512 25523
rect 11544 25491 11584 25523
rect 11616 25491 11656 25523
rect 11688 25491 11728 25523
rect 11760 25491 11800 25523
rect 11832 25491 11872 25523
rect 11904 25491 11944 25523
rect 11976 25491 12016 25523
rect 12048 25491 12088 25523
rect 12120 25491 12160 25523
rect 12192 25491 12232 25523
rect 12264 25491 12304 25523
rect 12336 25491 12376 25523
rect 12408 25491 12448 25523
rect 12480 25491 12520 25523
rect 12552 25491 12592 25523
rect 12624 25491 12664 25523
rect 12696 25491 12736 25523
rect 12768 25491 12808 25523
rect 12840 25491 12880 25523
rect 12912 25491 12952 25523
rect 12984 25491 13024 25523
rect 13056 25491 13096 25523
rect 13128 25491 13168 25523
rect 13200 25491 13240 25523
rect 13272 25491 13312 25523
rect 13344 25491 13384 25523
rect 13416 25491 13456 25523
rect 13488 25491 13528 25523
rect 13560 25491 13600 25523
rect 13632 25491 13672 25523
rect 13704 25491 13744 25523
rect 13776 25491 13816 25523
rect 13848 25491 13888 25523
rect 13920 25491 13960 25523
rect 13992 25491 14032 25523
rect 14064 25491 14104 25523
rect 14136 25491 14176 25523
rect 14208 25491 14248 25523
rect 14280 25491 14320 25523
rect 14352 25491 14392 25523
rect 14424 25491 14464 25523
rect 14496 25491 14536 25523
rect 14568 25491 14608 25523
rect 14640 25491 14680 25523
rect 14712 25491 14752 25523
rect 14784 25491 14824 25523
rect 14856 25491 14896 25523
rect 14928 25491 14968 25523
rect 15000 25491 15040 25523
rect 15072 25491 15112 25523
rect 15144 25491 15184 25523
rect 15216 25491 15256 25523
rect 15288 25491 15328 25523
rect 15360 25491 15400 25523
rect 15432 25491 15472 25523
rect 15504 25491 15544 25523
rect 15576 25491 15616 25523
rect 15648 25491 15688 25523
rect 15720 25491 15760 25523
rect 15792 25491 15832 25523
rect 15864 25491 15904 25523
rect 15936 25491 16000 25523
rect 0 25451 16000 25491
rect 0 25419 64 25451
rect 96 25419 136 25451
rect 168 25419 208 25451
rect 240 25419 280 25451
rect 312 25419 352 25451
rect 384 25419 424 25451
rect 456 25419 496 25451
rect 528 25419 568 25451
rect 600 25419 640 25451
rect 672 25419 712 25451
rect 744 25419 784 25451
rect 816 25419 856 25451
rect 888 25419 928 25451
rect 960 25419 1000 25451
rect 1032 25419 1072 25451
rect 1104 25419 1144 25451
rect 1176 25419 1216 25451
rect 1248 25419 1288 25451
rect 1320 25419 1360 25451
rect 1392 25419 1432 25451
rect 1464 25419 1504 25451
rect 1536 25419 1576 25451
rect 1608 25419 1648 25451
rect 1680 25419 1720 25451
rect 1752 25419 1792 25451
rect 1824 25419 1864 25451
rect 1896 25419 1936 25451
rect 1968 25419 2008 25451
rect 2040 25419 2080 25451
rect 2112 25419 2152 25451
rect 2184 25419 2224 25451
rect 2256 25419 2296 25451
rect 2328 25419 2368 25451
rect 2400 25419 2440 25451
rect 2472 25419 2512 25451
rect 2544 25419 2584 25451
rect 2616 25419 2656 25451
rect 2688 25419 2728 25451
rect 2760 25419 2800 25451
rect 2832 25419 2872 25451
rect 2904 25419 2944 25451
rect 2976 25419 3016 25451
rect 3048 25419 3088 25451
rect 3120 25419 3160 25451
rect 3192 25419 3232 25451
rect 3264 25419 3304 25451
rect 3336 25419 3376 25451
rect 3408 25419 3448 25451
rect 3480 25419 3520 25451
rect 3552 25419 3592 25451
rect 3624 25419 3664 25451
rect 3696 25419 3736 25451
rect 3768 25419 3808 25451
rect 3840 25419 3880 25451
rect 3912 25419 3952 25451
rect 3984 25419 4024 25451
rect 4056 25419 4096 25451
rect 4128 25419 4168 25451
rect 4200 25419 4240 25451
rect 4272 25419 4312 25451
rect 4344 25419 4384 25451
rect 4416 25419 4456 25451
rect 4488 25419 4528 25451
rect 4560 25419 4600 25451
rect 4632 25419 4672 25451
rect 4704 25419 4744 25451
rect 4776 25419 4816 25451
rect 4848 25419 4888 25451
rect 4920 25419 4960 25451
rect 4992 25419 5032 25451
rect 5064 25419 5104 25451
rect 5136 25419 5176 25451
rect 5208 25419 5248 25451
rect 5280 25419 5320 25451
rect 5352 25419 5392 25451
rect 5424 25419 5464 25451
rect 5496 25419 5536 25451
rect 5568 25419 5608 25451
rect 5640 25419 5680 25451
rect 5712 25419 5752 25451
rect 5784 25419 5824 25451
rect 5856 25419 5896 25451
rect 5928 25419 5968 25451
rect 6000 25419 6040 25451
rect 6072 25419 6112 25451
rect 6144 25419 6184 25451
rect 6216 25419 6256 25451
rect 6288 25419 6328 25451
rect 6360 25419 6400 25451
rect 6432 25419 6472 25451
rect 6504 25419 6544 25451
rect 6576 25419 6616 25451
rect 6648 25419 6688 25451
rect 6720 25419 6760 25451
rect 6792 25419 6832 25451
rect 6864 25419 6904 25451
rect 6936 25419 6976 25451
rect 7008 25419 7048 25451
rect 7080 25419 7120 25451
rect 7152 25419 7192 25451
rect 7224 25419 7264 25451
rect 7296 25419 7336 25451
rect 7368 25419 7408 25451
rect 7440 25419 7480 25451
rect 7512 25419 7552 25451
rect 7584 25419 7624 25451
rect 7656 25419 7696 25451
rect 7728 25419 7768 25451
rect 7800 25419 7840 25451
rect 7872 25419 7912 25451
rect 7944 25419 7984 25451
rect 8016 25419 8056 25451
rect 8088 25419 8128 25451
rect 8160 25419 8200 25451
rect 8232 25419 8272 25451
rect 8304 25419 8344 25451
rect 8376 25419 8416 25451
rect 8448 25419 8488 25451
rect 8520 25419 8560 25451
rect 8592 25419 8632 25451
rect 8664 25419 8704 25451
rect 8736 25419 8776 25451
rect 8808 25419 8848 25451
rect 8880 25419 8920 25451
rect 8952 25419 8992 25451
rect 9024 25419 9064 25451
rect 9096 25419 9136 25451
rect 9168 25419 9208 25451
rect 9240 25419 9280 25451
rect 9312 25419 9352 25451
rect 9384 25419 9424 25451
rect 9456 25419 9496 25451
rect 9528 25419 9568 25451
rect 9600 25419 9640 25451
rect 9672 25419 9712 25451
rect 9744 25419 9784 25451
rect 9816 25419 9856 25451
rect 9888 25419 9928 25451
rect 9960 25419 10000 25451
rect 10032 25419 10072 25451
rect 10104 25419 10144 25451
rect 10176 25419 10216 25451
rect 10248 25419 10288 25451
rect 10320 25419 10360 25451
rect 10392 25419 10432 25451
rect 10464 25419 10504 25451
rect 10536 25419 10576 25451
rect 10608 25419 10648 25451
rect 10680 25419 10720 25451
rect 10752 25419 10792 25451
rect 10824 25419 10864 25451
rect 10896 25419 10936 25451
rect 10968 25419 11008 25451
rect 11040 25419 11080 25451
rect 11112 25419 11152 25451
rect 11184 25419 11224 25451
rect 11256 25419 11296 25451
rect 11328 25419 11368 25451
rect 11400 25419 11440 25451
rect 11472 25419 11512 25451
rect 11544 25419 11584 25451
rect 11616 25419 11656 25451
rect 11688 25419 11728 25451
rect 11760 25419 11800 25451
rect 11832 25419 11872 25451
rect 11904 25419 11944 25451
rect 11976 25419 12016 25451
rect 12048 25419 12088 25451
rect 12120 25419 12160 25451
rect 12192 25419 12232 25451
rect 12264 25419 12304 25451
rect 12336 25419 12376 25451
rect 12408 25419 12448 25451
rect 12480 25419 12520 25451
rect 12552 25419 12592 25451
rect 12624 25419 12664 25451
rect 12696 25419 12736 25451
rect 12768 25419 12808 25451
rect 12840 25419 12880 25451
rect 12912 25419 12952 25451
rect 12984 25419 13024 25451
rect 13056 25419 13096 25451
rect 13128 25419 13168 25451
rect 13200 25419 13240 25451
rect 13272 25419 13312 25451
rect 13344 25419 13384 25451
rect 13416 25419 13456 25451
rect 13488 25419 13528 25451
rect 13560 25419 13600 25451
rect 13632 25419 13672 25451
rect 13704 25419 13744 25451
rect 13776 25419 13816 25451
rect 13848 25419 13888 25451
rect 13920 25419 13960 25451
rect 13992 25419 14032 25451
rect 14064 25419 14104 25451
rect 14136 25419 14176 25451
rect 14208 25419 14248 25451
rect 14280 25419 14320 25451
rect 14352 25419 14392 25451
rect 14424 25419 14464 25451
rect 14496 25419 14536 25451
rect 14568 25419 14608 25451
rect 14640 25419 14680 25451
rect 14712 25419 14752 25451
rect 14784 25419 14824 25451
rect 14856 25419 14896 25451
rect 14928 25419 14968 25451
rect 15000 25419 15040 25451
rect 15072 25419 15112 25451
rect 15144 25419 15184 25451
rect 15216 25419 15256 25451
rect 15288 25419 15328 25451
rect 15360 25419 15400 25451
rect 15432 25419 15472 25451
rect 15504 25419 15544 25451
rect 15576 25419 15616 25451
rect 15648 25419 15688 25451
rect 15720 25419 15760 25451
rect 15792 25419 15832 25451
rect 15864 25419 15904 25451
rect 15936 25419 16000 25451
rect 0 25379 16000 25419
rect 0 25347 64 25379
rect 96 25347 136 25379
rect 168 25347 208 25379
rect 240 25347 280 25379
rect 312 25347 352 25379
rect 384 25347 424 25379
rect 456 25347 496 25379
rect 528 25347 568 25379
rect 600 25347 640 25379
rect 672 25347 712 25379
rect 744 25347 784 25379
rect 816 25347 856 25379
rect 888 25347 928 25379
rect 960 25347 1000 25379
rect 1032 25347 1072 25379
rect 1104 25347 1144 25379
rect 1176 25347 1216 25379
rect 1248 25347 1288 25379
rect 1320 25347 1360 25379
rect 1392 25347 1432 25379
rect 1464 25347 1504 25379
rect 1536 25347 1576 25379
rect 1608 25347 1648 25379
rect 1680 25347 1720 25379
rect 1752 25347 1792 25379
rect 1824 25347 1864 25379
rect 1896 25347 1936 25379
rect 1968 25347 2008 25379
rect 2040 25347 2080 25379
rect 2112 25347 2152 25379
rect 2184 25347 2224 25379
rect 2256 25347 2296 25379
rect 2328 25347 2368 25379
rect 2400 25347 2440 25379
rect 2472 25347 2512 25379
rect 2544 25347 2584 25379
rect 2616 25347 2656 25379
rect 2688 25347 2728 25379
rect 2760 25347 2800 25379
rect 2832 25347 2872 25379
rect 2904 25347 2944 25379
rect 2976 25347 3016 25379
rect 3048 25347 3088 25379
rect 3120 25347 3160 25379
rect 3192 25347 3232 25379
rect 3264 25347 3304 25379
rect 3336 25347 3376 25379
rect 3408 25347 3448 25379
rect 3480 25347 3520 25379
rect 3552 25347 3592 25379
rect 3624 25347 3664 25379
rect 3696 25347 3736 25379
rect 3768 25347 3808 25379
rect 3840 25347 3880 25379
rect 3912 25347 3952 25379
rect 3984 25347 4024 25379
rect 4056 25347 4096 25379
rect 4128 25347 4168 25379
rect 4200 25347 4240 25379
rect 4272 25347 4312 25379
rect 4344 25347 4384 25379
rect 4416 25347 4456 25379
rect 4488 25347 4528 25379
rect 4560 25347 4600 25379
rect 4632 25347 4672 25379
rect 4704 25347 4744 25379
rect 4776 25347 4816 25379
rect 4848 25347 4888 25379
rect 4920 25347 4960 25379
rect 4992 25347 5032 25379
rect 5064 25347 5104 25379
rect 5136 25347 5176 25379
rect 5208 25347 5248 25379
rect 5280 25347 5320 25379
rect 5352 25347 5392 25379
rect 5424 25347 5464 25379
rect 5496 25347 5536 25379
rect 5568 25347 5608 25379
rect 5640 25347 5680 25379
rect 5712 25347 5752 25379
rect 5784 25347 5824 25379
rect 5856 25347 5896 25379
rect 5928 25347 5968 25379
rect 6000 25347 6040 25379
rect 6072 25347 6112 25379
rect 6144 25347 6184 25379
rect 6216 25347 6256 25379
rect 6288 25347 6328 25379
rect 6360 25347 6400 25379
rect 6432 25347 6472 25379
rect 6504 25347 6544 25379
rect 6576 25347 6616 25379
rect 6648 25347 6688 25379
rect 6720 25347 6760 25379
rect 6792 25347 6832 25379
rect 6864 25347 6904 25379
rect 6936 25347 6976 25379
rect 7008 25347 7048 25379
rect 7080 25347 7120 25379
rect 7152 25347 7192 25379
rect 7224 25347 7264 25379
rect 7296 25347 7336 25379
rect 7368 25347 7408 25379
rect 7440 25347 7480 25379
rect 7512 25347 7552 25379
rect 7584 25347 7624 25379
rect 7656 25347 7696 25379
rect 7728 25347 7768 25379
rect 7800 25347 7840 25379
rect 7872 25347 7912 25379
rect 7944 25347 7984 25379
rect 8016 25347 8056 25379
rect 8088 25347 8128 25379
rect 8160 25347 8200 25379
rect 8232 25347 8272 25379
rect 8304 25347 8344 25379
rect 8376 25347 8416 25379
rect 8448 25347 8488 25379
rect 8520 25347 8560 25379
rect 8592 25347 8632 25379
rect 8664 25347 8704 25379
rect 8736 25347 8776 25379
rect 8808 25347 8848 25379
rect 8880 25347 8920 25379
rect 8952 25347 8992 25379
rect 9024 25347 9064 25379
rect 9096 25347 9136 25379
rect 9168 25347 9208 25379
rect 9240 25347 9280 25379
rect 9312 25347 9352 25379
rect 9384 25347 9424 25379
rect 9456 25347 9496 25379
rect 9528 25347 9568 25379
rect 9600 25347 9640 25379
rect 9672 25347 9712 25379
rect 9744 25347 9784 25379
rect 9816 25347 9856 25379
rect 9888 25347 9928 25379
rect 9960 25347 10000 25379
rect 10032 25347 10072 25379
rect 10104 25347 10144 25379
rect 10176 25347 10216 25379
rect 10248 25347 10288 25379
rect 10320 25347 10360 25379
rect 10392 25347 10432 25379
rect 10464 25347 10504 25379
rect 10536 25347 10576 25379
rect 10608 25347 10648 25379
rect 10680 25347 10720 25379
rect 10752 25347 10792 25379
rect 10824 25347 10864 25379
rect 10896 25347 10936 25379
rect 10968 25347 11008 25379
rect 11040 25347 11080 25379
rect 11112 25347 11152 25379
rect 11184 25347 11224 25379
rect 11256 25347 11296 25379
rect 11328 25347 11368 25379
rect 11400 25347 11440 25379
rect 11472 25347 11512 25379
rect 11544 25347 11584 25379
rect 11616 25347 11656 25379
rect 11688 25347 11728 25379
rect 11760 25347 11800 25379
rect 11832 25347 11872 25379
rect 11904 25347 11944 25379
rect 11976 25347 12016 25379
rect 12048 25347 12088 25379
rect 12120 25347 12160 25379
rect 12192 25347 12232 25379
rect 12264 25347 12304 25379
rect 12336 25347 12376 25379
rect 12408 25347 12448 25379
rect 12480 25347 12520 25379
rect 12552 25347 12592 25379
rect 12624 25347 12664 25379
rect 12696 25347 12736 25379
rect 12768 25347 12808 25379
rect 12840 25347 12880 25379
rect 12912 25347 12952 25379
rect 12984 25347 13024 25379
rect 13056 25347 13096 25379
rect 13128 25347 13168 25379
rect 13200 25347 13240 25379
rect 13272 25347 13312 25379
rect 13344 25347 13384 25379
rect 13416 25347 13456 25379
rect 13488 25347 13528 25379
rect 13560 25347 13600 25379
rect 13632 25347 13672 25379
rect 13704 25347 13744 25379
rect 13776 25347 13816 25379
rect 13848 25347 13888 25379
rect 13920 25347 13960 25379
rect 13992 25347 14032 25379
rect 14064 25347 14104 25379
rect 14136 25347 14176 25379
rect 14208 25347 14248 25379
rect 14280 25347 14320 25379
rect 14352 25347 14392 25379
rect 14424 25347 14464 25379
rect 14496 25347 14536 25379
rect 14568 25347 14608 25379
rect 14640 25347 14680 25379
rect 14712 25347 14752 25379
rect 14784 25347 14824 25379
rect 14856 25347 14896 25379
rect 14928 25347 14968 25379
rect 15000 25347 15040 25379
rect 15072 25347 15112 25379
rect 15144 25347 15184 25379
rect 15216 25347 15256 25379
rect 15288 25347 15328 25379
rect 15360 25347 15400 25379
rect 15432 25347 15472 25379
rect 15504 25347 15544 25379
rect 15576 25347 15616 25379
rect 15648 25347 15688 25379
rect 15720 25347 15760 25379
rect 15792 25347 15832 25379
rect 15864 25347 15904 25379
rect 15936 25347 16000 25379
rect 0 25307 16000 25347
rect 0 25275 64 25307
rect 96 25275 136 25307
rect 168 25275 208 25307
rect 240 25275 280 25307
rect 312 25275 352 25307
rect 384 25275 424 25307
rect 456 25275 496 25307
rect 528 25275 568 25307
rect 600 25275 640 25307
rect 672 25275 712 25307
rect 744 25275 784 25307
rect 816 25275 856 25307
rect 888 25275 928 25307
rect 960 25275 1000 25307
rect 1032 25275 1072 25307
rect 1104 25275 1144 25307
rect 1176 25275 1216 25307
rect 1248 25275 1288 25307
rect 1320 25275 1360 25307
rect 1392 25275 1432 25307
rect 1464 25275 1504 25307
rect 1536 25275 1576 25307
rect 1608 25275 1648 25307
rect 1680 25275 1720 25307
rect 1752 25275 1792 25307
rect 1824 25275 1864 25307
rect 1896 25275 1936 25307
rect 1968 25275 2008 25307
rect 2040 25275 2080 25307
rect 2112 25275 2152 25307
rect 2184 25275 2224 25307
rect 2256 25275 2296 25307
rect 2328 25275 2368 25307
rect 2400 25275 2440 25307
rect 2472 25275 2512 25307
rect 2544 25275 2584 25307
rect 2616 25275 2656 25307
rect 2688 25275 2728 25307
rect 2760 25275 2800 25307
rect 2832 25275 2872 25307
rect 2904 25275 2944 25307
rect 2976 25275 3016 25307
rect 3048 25275 3088 25307
rect 3120 25275 3160 25307
rect 3192 25275 3232 25307
rect 3264 25275 3304 25307
rect 3336 25275 3376 25307
rect 3408 25275 3448 25307
rect 3480 25275 3520 25307
rect 3552 25275 3592 25307
rect 3624 25275 3664 25307
rect 3696 25275 3736 25307
rect 3768 25275 3808 25307
rect 3840 25275 3880 25307
rect 3912 25275 3952 25307
rect 3984 25275 4024 25307
rect 4056 25275 4096 25307
rect 4128 25275 4168 25307
rect 4200 25275 4240 25307
rect 4272 25275 4312 25307
rect 4344 25275 4384 25307
rect 4416 25275 4456 25307
rect 4488 25275 4528 25307
rect 4560 25275 4600 25307
rect 4632 25275 4672 25307
rect 4704 25275 4744 25307
rect 4776 25275 4816 25307
rect 4848 25275 4888 25307
rect 4920 25275 4960 25307
rect 4992 25275 5032 25307
rect 5064 25275 5104 25307
rect 5136 25275 5176 25307
rect 5208 25275 5248 25307
rect 5280 25275 5320 25307
rect 5352 25275 5392 25307
rect 5424 25275 5464 25307
rect 5496 25275 5536 25307
rect 5568 25275 5608 25307
rect 5640 25275 5680 25307
rect 5712 25275 5752 25307
rect 5784 25275 5824 25307
rect 5856 25275 5896 25307
rect 5928 25275 5968 25307
rect 6000 25275 6040 25307
rect 6072 25275 6112 25307
rect 6144 25275 6184 25307
rect 6216 25275 6256 25307
rect 6288 25275 6328 25307
rect 6360 25275 6400 25307
rect 6432 25275 6472 25307
rect 6504 25275 6544 25307
rect 6576 25275 6616 25307
rect 6648 25275 6688 25307
rect 6720 25275 6760 25307
rect 6792 25275 6832 25307
rect 6864 25275 6904 25307
rect 6936 25275 6976 25307
rect 7008 25275 7048 25307
rect 7080 25275 7120 25307
rect 7152 25275 7192 25307
rect 7224 25275 7264 25307
rect 7296 25275 7336 25307
rect 7368 25275 7408 25307
rect 7440 25275 7480 25307
rect 7512 25275 7552 25307
rect 7584 25275 7624 25307
rect 7656 25275 7696 25307
rect 7728 25275 7768 25307
rect 7800 25275 7840 25307
rect 7872 25275 7912 25307
rect 7944 25275 7984 25307
rect 8016 25275 8056 25307
rect 8088 25275 8128 25307
rect 8160 25275 8200 25307
rect 8232 25275 8272 25307
rect 8304 25275 8344 25307
rect 8376 25275 8416 25307
rect 8448 25275 8488 25307
rect 8520 25275 8560 25307
rect 8592 25275 8632 25307
rect 8664 25275 8704 25307
rect 8736 25275 8776 25307
rect 8808 25275 8848 25307
rect 8880 25275 8920 25307
rect 8952 25275 8992 25307
rect 9024 25275 9064 25307
rect 9096 25275 9136 25307
rect 9168 25275 9208 25307
rect 9240 25275 9280 25307
rect 9312 25275 9352 25307
rect 9384 25275 9424 25307
rect 9456 25275 9496 25307
rect 9528 25275 9568 25307
rect 9600 25275 9640 25307
rect 9672 25275 9712 25307
rect 9744 25275 9784 25307
rect 9816 25275 9856 25307
rect 9888 25275 9928 25307
rect 9960 25275 10000 25307
rect 10032 25275 10072 25307
rect 10104 25275 10144 25307
rect 10176 25275 10216 25307
rect 10248 25275 10288 25307
rect 10320 25275 10360 25307
rect 10392 25275 10432 25307
rect 10464 25275 10504 25307
rect 10536 25275 10576 25307
rect 10608 25275 10648 25307
rect 10680 25275 10720 25307
rect 10752 25275 10792 25307
rect 10824 25275 10864 25307
rect 10896 25275 10936 25307
rect 10968 25275 11008 25307
rect 11040 25275 11080 25307
rect 11112 25275 11152 25307
rect 11184 25275 11224 25307
rect 11256 25275 11296 25307
rect 11328 25275 11368 25307
rect 11400 25275 11440 25307
rect 11472 25275 11512 25307
rect 11544 25275 11584 25307
rect 11616 25275 11656 25307
rect 11688 25275 11728 25307
rect 11760 25275 11800 25307
rect 11832 25275 11872 25307
rect 11904 25275 11944 25307
rect 11976 25275 12016 25307
rect 12048 25275 12088 25307
rect 12120 25275 12160 25307
rect 12192 25275 12232 25307
rect 12264 25275 12304 25307
rect 12336 25275 12376 25307
rect 12408 25275 12448 25307
rect 12480 25275 12520 25307
rect 12552 25275 12592 25307
rect 12624 25275 12664 25307
rect 12696 25275 12736 25307
rect 12768 25275 12808 25307
rect 12840 25275 12880 25307
rect 12912 25275 12952 25307
rect 12984 25275 13024 25307
rect 13056 25275 13096 25307
rect 13128 25275 13168 25307
rect 13200 25275 13240 25307
rect 13272 25275 13312 25307
rect 13344 25275 13384 25307
rect 13416 25275 13456 25307
rect 13488 25275 13528 25307
rect 13560 25275 13600 25307
rect 13632 25275 13672 25307
rect 13704 25275 13744 25307
rect 13776 25275 13816 25307
rect 13848 25275 13888 25307
rect 13920 25275 13960 25307
rect 13992 25275 14032 25307
rect 14064 25275 14104 25307
rect 14136 25275 14176 25307
rect 14208 25275 14248 25307
rect 14280 25275 14320 25307
rect 14352 25275 14392 25307
rect 14424 25275 14464 25307
rect 14496 25275 14536 25307
rect 14568 25275 14608 25307
rect 14640 25275 14680 25307
rect 14712 25275 14752 25307
rect 14784 25275 14824 25307
rect 14856 25275 14896 25307
rect 14928 25275 14968 25307
rect 15000 25275 15040 25307
rect 15072 25275 15112 25307
rect 15144 25275 15184 25307
rect 15216 25275 15256 25307
rect 15288 25275 15328 25307
rect 15360 25275 15400 25307
rect 15432 25275 15472 25307
rect 15504 25275 15544 25307
rect 15576 25275 15616 25307
rect 15648 25275 15688 25307
rect 15720 25275 15760 25307
rect 15792 25275 15832 25307
rect 15864 25275 15904 25307
rect 15936 25275 16000 25307
rect 0 25235 16000 25275
rect 0 25203 64 25235
rect 96 25203 136 25235
rect 168 25203 208 25235
rect 240 25203 280 25235
rect 312 25203 352 25235
rect 384 25203 424 25235
rect 456 25203 496 25235
rect 528 25203 568 25235
rect 600 25203 640 25235
rect 672 25203 712 25235
rect 744 25203 784 25235
rect 816 25203 856 25235
rect 888 25203 928 25235
rect 960 25203 1000 25235
rect 1032 25203 1072 25235
rect 1104 25203 1144 25235
rect 1176 25203 1216 25235
rect 1248 25203 1288 25235
rect 1320 25203 1360 25235
rect 1392 25203 1432 25235
rect 1464 25203 1504 25235
rect 1536 25203 1576 25235
rect 1608 25203 1648 25235
rect 1680 25203 1720 25235
rect 1752 25203 1792 25235
rect 1824 25203 1864 25235
rect 1896 25203 1936 25235
rect 1968 25203 2008 25235
rect 2040 25203 2080 25235
rect 2112 25203 2152 25235
rect 2184 25203 2224 25235
rect 2256 25203 2296 25235
rect 2328 25203 2368 25235
rect 2400 25203 2440 25235
rect 2472 25203 2512 25235
rect 2544 25203 2584 25235
rect 2616 25203 2656 25235
rect 2688 25203 2728 25235
rect 2760 25203 2800 25235
rect 2832 25203 2872 25235
rect 2904 25203 2944 25235
rect 2976 25203 3016 25235
rect 3048 25203 3088 25235
rect 3120 25203 3160 25235
rect 3192 25203 3232 25235
rect 3264 25203 3304 25235
rect 3336 25203 3376 25235
rect 3408 25203 3448 25235
rect 3480 25203 3520 25235
rect 3552 25203 3592 25235
rect 3624 25203 3664 25235
rect 3696 25203 3736 25235
rect 3768 25203 3808 25235
rect 3840 25203 3880 25235
rect 3912 25203 3952 25235
rect 3984 25203 4024 25235
rect 4056 25203 4096 25235
rect 4128 25203 4168 25235
rect 4200 25203 4240 25235
rect 4272 25203 4312 25235
rect 4344 25203 4384 25235
rect 4416 25203 4456 25235
rect 4488 25203 4528 25235
rect 4560 25203 4600 25235
rect 4632 25203 4672 25235
rect 4704 25203 4744 25235
rect 4776 25203 4816 25235
rect 4848 25203 4888 25235
rect 4920 25203 4960 25235
rect 4992 25203 5032 25235
rect 5064 25203 5104 25235
rect 5136 25203 5176 25235
rect 5208 25203 5248 25235
rect 5280 25203 5320 25235
rect 5352 25203 5392 25235
rect 5424 25203 5464 25235
rect 5496 25203 5536 25235
rect 5568 25203 5608 25235
rect 5640 25203 5680 25235
rect 5712 25203 5752 25235
rect 5784 25203 5824 25235
rect 5856 25203 5896 25235
rect 5928 25203 5968 25235
rect 6000 25203 6040 25235
rect 6072 25203 6112 25235
rect 6144 25203 6184 25235
rect 6216 25203 6256 25235
rect 6288 25203 6328 25235
rect 6360 25203 6400 25235
rect 6432 25203 6472 25235
rect 6504 25203 6544 25235
rect 6576 25203 6616 25235
rect 6648 25203 6688 25235
rect 6720 25203 6760 25235
rect 6792 25203 6832 25235
rect 6864 25203 6904 25235
rect 6936 25203 6976 25235
rect 7008 25203 7048 25235
rect 7080 25203 7120 25235
rect 7152 25203 7192 25235
rect 7224 25203 7264 25235
rect 7296 25203 7336 25235
rect 7368 25203 7408 25235
rect 7440 25203 7480 25235
rect 7512 25203 7552 25235
rect 7584 25203 7624 25235
rect 7656 25203 7696 25235
rect 7728 25203 7768 25235
rect 7800 25203 7840 25235
rect 7872 25203 7912 25235
rect 7944 25203 7984 25235
rect 8016 25203 8056 25235
rect 8088 25203 8128 25235
rect 8160 25203 8200 25235
rect 8232 25203 8272 25235
rect 8304 25203 8344 25235
rect 8376 25203 8416 25235
rect 8448 25203 8488 25235
rect 8520 25203 8560 25235
rect 8592 25203 8632 25235
rect 8664 25203 8704 25235
rect 8736 25203 8776 25235
rect 8808 25203 8848 25235
rect 8880 25203 8920 25235
rect 8952 25203 8992 25235
rect 9024 25203 9064 25235
rect 9096 25203 9136 25235
rect 9168 25203 9208 25235
rect 9240 25203 9280 25235
rect 9312 25203 9352 25235
rect 9384 25203 9424 25235
rect 9456 25203 9496 25235
rect 9528 25203 9568 25235
rect 9600 25203 9640 25235
rect 9672 25203 9712 25235
rect 9744 25203 9784 25235
rect 9816 25203 9856 25235
rect 9888 25203 9928 25235
rect 9960 25203 10000 25235
rect 10032 25203 10072 25235
rect 10104 25203 10144 25235
rect 10176 25203 10216 25235
rect 10248 25203 10288 25235
rect 10320 25203 10360 25235
rect 10392 25203 10432 25235
rect 10464 25203 10504 25235
rect 10536 25203 10576 25235
rect 10608 25203 10648 25235
rect 10680 25203 10720 25235
rect 10752 25203 10792 25235
rect 10824 25203 10864 25235
rect 10896 25203 10936 25235
rect 10968 25203 11008 25235
rect 11040 25203 11080 25235
rect 11112 25203 11152 25235
rect 11184 25203 11224 25235
rect 11256 25203 11296 25235
rect 11328 25203 11368 25235
rect 11400 25203 11440 25235
rect 11472 25203 11512 25235
rect 11544 25203 11584 25235
rect 11616 25203 11656 25235
rect 11688 25203 11728 25235
rect 11760 25203 11800 25235
rect 11832 25203 11872 25235
rect 11904 25203 11944 25235
rect 11976 25203 12016 25235
rect 12048 25203 12088 25235
rect 12120 25203 12160 25235
rect 12192 25203 12232 25235
rect 12264 25203 12304 25235
rect 12336 25203 12376 25235
rect 12408 25203 12448 25235
rect 12480 25203 12520 25235
rect 12552 25203 12592 25235
rect 12624 25203 12664 25235
rect 12696 25203 12736 25235
rect 12768 25203 12808 25235
rect 12840 25203 12880 25235
rect 12912 25203 12952 25235
rect 12984 25203 13024 25235
rect 13056 25203 13096 25235
rect 13128 25203 13168 25235
rect 13200 25203 13240 25235
rect 13272 25203 13312 25235
rect 13344 25203 13384 25235
rect 13416 25203 13456 25235
rect 13488 25203 13528 25235
rect 13560 25203 13600 25235
rect 13632 25203 13672 25235
rect 13704 25203 13744 25235
rect 13776 25203 13816 25235
rect 13848 25203 13888 25235
rect 13920 25203 13960 25235
rect 13992 25203 14032 25235
rect 14064 25203 14104 25235
rect 14136 25203 14176 25235
rect 14208 25203 14248 25235
rect 14280 25203 14320 25235
rect 14352 25203 14392 25235
rect 14424 25203 14464 25235
rect 14496 25203 14536 25235
rect 14568 25203 14608 25235
rect 14640 25203 14680 25235
rect 14712 25203 14752 25235
rect 14784 25203 14824 25235
rect 14856 25203 14896 25235
rect 14928 25203 14968 25235
rect 15000 25203 15040 25235
rect 15072 25203 15112 25235
rect 15144 25203 15184 25235
rect 15216 25203 15256 25235
rect 15288 25203 15328 25235
rect 15360 25203 15400 25235
rect 15432 25203 15472 25235
rect 15504 25203 15544 25235
rect 15576 25203 15616 25235
rect 15648 25203 15688 25235
rect 15720 25203 15760 25235
rect 15792 25203 15832 25235
rect 15864 25203 15904 25235
rect 15936 25203 16000 25235
rect 0 25163 16000 25203
rect 0 25131 64 25163
rect 96 25131 136 25163
rect 168 25131 208 25163
rect 240 25131 280 25163
rect 312 25131 352 25163
rect 384 25131 424 25163
rect 456 25131 496 25163
rect 528 25131 568 25163
rect 600 25131 640 25163
rect 672 25131 712 25163
rect 744 25131 784 25163
rect 816 25131 856 25163
rect 888 25131 928 25163
rect 960 25131 1000 25163
rect 1032 25131 1072 25163
rect 1104 25131 1144 25163
rect 1176 25131 1216 25163
rect 1248 25131 1288 25163
rect 1320 25131 1360 25163
rect 1392 25131 1432 25163
rect 1464 25131 1504 25163
rect 1536 25131 1576 25163
rect 1608 25131 1648 25163
rect 1680 25131 1720 25163
rect 1752 25131 1792 25163
rect 1824 25131 1864 25163
rect 1896 25131 1936 25163
rect 1968 25131 2008 25163
rect 2040 25131 2080 25163
rect 2112 25131 2152 25163
rect 2184 25131 2224 25163
rect 2256 25131 2296 25163
rect 2328 25131 2368 25163
rect 2400 25131 2440 25163
rect 2472 25131 2512 25163
rect 2544 25131 2584 25163
rect 2616 25131 2656 25163
rect 2688 25131 2728 25163
rect 2760 25131 2800 25163
rect 2832 25131 2872 25163
rect 2904 25131 2944 25163
rect 2976 25131 3016 25163
rect 3048 25131 3088 25163
rect 3120 25131 3160 25163
rect 3192 25131 3232 25163
rect 3264 25131 3304 25163
rect 3336 25131 3376 25163
rect 3408 25131 3448 25163
rect 3480 25131 3520 25163
rect 3552 25131 3592 25163
rect 3624 25131 3664 25163
rect 3696 25131 3736 25163
rect 3768 25131 3808 25163
rect 3840 25131 3880 25163
rect 3912 25131 3952 25163
rect 3984 25131 4024 25163
rect 4056 25131 4096 25163
rect 4128 25131 4168 25163
rect 4200 25131 4240 25163
rect 4272 25131 4312 25163
rect 4344 25131 4384 25163
rect 4416 25131 4456 25163
rect 4488 25131 4528 25163
rect 4560 25131 4600 25163
rect 4632 25131 4672 25163
rect 4704 25131 4744 25163
rect 4776 25131 4816 25163
rect 4848 25131 4888 25163
rect 4920 25131 4960 25163
rect 4992 25131 5032 25163
rect 5064 25131 5104 25163
rect 5136 25131 5176 25163
rect 5208 25131 5248 25163
rect 5280 25131 5320 25163
rect 5352 25131 5392 25163
rect 5424 25131 5464 25163
rect 5496 25131 5536 25163
rect 5568 25131 5608 25163
rect 5640 25131 5680 25163
rect 5712 25131 5752 25163
rect 5784 25131 5824 25163
rect 5856 25131 5896 25163
rect 5928 25131 5968 25163
rect 6000 25131 6040 25163
rect 6072 25131 6112 25163
rect 6144 25131 6184 25163
rect 6216 25131 6256 25163
rect 6288 25131 6328 25163
rect 6360 25131 6400 25163
rect 6432 25131 6472 25163
rect 6504 25131 6544 25163
rect 6576 25131 6616 25163
rect 6648 25131 6688 25163
rect 6720 25131 6760 25163
rect 6792 25131 6832 25163
rect 6864 25131 6904 25163
rect 6936 25131 6976 25163
rect 7008 25131 7048 25163
rect 7080 25131 7120 25163
rect 7152 25131 7192 25163
rect 7224 25131 7264 25163
rect 7296 25131 7336 25163
rect 7368 25131 7408 25163
rect 7440 25131 7480 25163
rect 7512 25131 7552 25163
rect 7584 25131 7624 25163
rect 7656 25131 7696 25163
rect 7728 25131 7768 25163
rect 7800 25131 7840 25163
rect 7872 25131 7912 25163
rect 7944 25131 7984 25163
rect 8016 25131 8056 25163
rect 8088 25131 8128 25163
rect 8160 25131 8200 25163
rect 8232 25131 8272 25163
rect 8304 25131 8344 25163
rect 8376 25131 8416 25163
rect 8448 25131 8488 25163
rect 8520 25131 8560 25163
rect 8592 25131 8632 25163
rect 8664 25131 8704 25163
rect 8736 25131 8776 25163
rect 8808 25131 8848 25163
rect 8880 25131 8920 25163
rect 8952 25131 8992 25163
rect 9024 25131 9064 25163
rect 9096 25131 9136 25163
rect 9168 25131 9208 25163
rect 9240 25131 9280 25163
rect 9312 25131 9352 25163
rect 9384 25131 9424 25163
rect 9456 25131 9496 25163
rect 9528 25131 9568 25163
rect 9600 25131 9640 25163
rect 9672 25131 9712 25163
rect 9744 25131 9784 25163
rect 9816 25131 9856 25163
rect 9888 25131 9928 25163
rect 9960 25131 10000 25163
rect 10032 25131 10072 25163
rect 10104 25131 10144 25163
rect 10176 25131 10216 25163
rect 10248 25131 10288 25163
rect 10320 25131 10360 25163
rect 10392 25131 10432 25163
rect 10464 25131 10504 25163
rect 10536 25131 10576 25163
rect 10608 25131 10648 25163
rect 10680 25131 10720 25163
rect 10752 25131 10792 25163
rect 10824 25131 10864 25163
rect 10896 25131 10936 25163
rect 10968 25131 11008 25163
rect 11040 25131 11080 25163
rect 11112 25131 11152 25163
rect 11184 25131 11224 25163
rect 11256 25131 11296 25163
rect 11328 25131 11368 25163
rect 11400 25131 11440 25163
rect 11472 25131 11512 25163
rect 11544 25131 11584 25163
rect 11616 25131 11656 25163
rect 11688 25131 11728 25163
rect 11760 25131 11800 25163
rect 11832 25131 11872 25163
rect 11904 25131 11944 25163
rect 11976 25131 12016 25163
rect 12048 25131 12088 25163
rect 12120 25131 12160 25163
rect 12192 25131 12232 25163
rect 12264 25131 12304 25163
rect 12336 25131 12376 25163
rect 12408 25131 12448 25163
rect 12480 25131 12520 25163
rect 12552 25131 12592 25163
rect 12624 25131 12664 25163
rect 12696 25131 12736 25163
rect 12768 25131 12808 25163
rect 12840 25131 12880 25163
rect 12912 25131 12952 25163
rect 12984 25131 13024 25163
rect 13056 25131 13096 25163
rect 13128 25131 13168 25163
rect 13200 25131 13240 25163
rect 13272 25131 13312 25163
rect 13344 25131 13384 25163
rect 13416 25131 13456 25163
rect 13488 25131 13528 25163
rect 13560 25131 13600 25163
rect 13632 25131 13672 25163
rect 13704 25131 13744 25163
rect 13776 25131 13816 25163
rect 13848 25131 13888 25163
rect 13920 25131 13960 25163
rect 13992 25131 14032 25163
rect 14064 25131 14104 25163
rect 14136 25131 14176 25163
rect 14208 25131 14248 25163
rect 14280 25131 14320 25163
rect 14352 25131 14392 25163
rect 14424 25131 14464 25163
rect 14496 25131 14536 25163
rect 14568 25131 14608 25163
rect 14640 25131 14680 25163
rect 14712 25131 14752 25163
rect 14784 25131 14824 25163
rect 14856 25131 14896 25163
rect 14928 25131 14968 25163
rect 15000 25131 15040 25163
rect 15072 25131 15112 25163
rect 15144 25131 15184 25163
rect 15216 25131 15256 25163
rect 15288 25131 15328 25163
rect 15360 25131 15400 25163
rect 15432 25131 15472 25163
rect 15504 25131 15544 25163
rect 15576 25131 15616 25163
rect 15648 25131 15688 25163
rect 15720 25131 15760 25163
rect 15792 25131 15832 25163
rect 15864 25131 15904 25163
rect 15936 25131 16000 25163
rect 0 25091 16000 25131
rect 0 25059 64 25091
rect 96 25059 136 25091
rect 168 25059 208 25091
rect 240 25059 280 25091
rect 312 25059 352 25091
rect 384 25059 424 25091
rect 456 25059 496 25091
rect 528 25059 568 25091
rect 600 25059 640 25091
rect 672 25059 712 25091
rect 744 25059 784 25091
rect 816 25059 856 25091
rect 888 25059 928 25091
rect 960 25059 1000 25091
rect 1032 25059 1072 25091
rect 1104 25059 1144 25091
rect 1176 25059 1216 25091
rect 1248 25059 1288 25091
rect 1320 25059 1360 25091
rect 1392 25059 1432 25091
rect 1464 25059 1504 25091
rect 1536 25059 1576 25091
rect 1608 25059 1648 25091
rect 1680 25059 1720 25091
rect 1752 25059 1792 25091
rect 1824 25059 1864 25091
rect 1896 25059 1936 25091
rect 1968 25059 2008 25091
rect 2040 25059 2080 25091
rect 2112 25059 2152 25091
rect 2184 25059 2224 25091
rect 2256 25059 2296 25091
rect 2328 25059 2368 25091
rect 2400 25059 2440 25091
rect 2472 25059 2512 25091
rect 2544 25059 2584 25091
rect 2616 25059 2656 25091
rect 2688 25059 2728 25091
rect 2760 25059 2800 25091
rect 2832 25059 2872 25091
rect 2904 25059 2944 25091
rect 2976 25059 3016 25091
rect 3048 25059 3088 25091
rect 3120 25059 3160 25091
rect 3192 25059 3232 25091
rect 3264 25059 3304 25091
rect 3336 25059 3376 25091
rect 3408 25059 3448 25091
rect 3480 25059 3520 25091
rect 3552 25059 3592 25091
rect 3624 25059 3664 25091
rect 3696 25059 3736 25091
rect 3768 25059 3808 25091
rect 3840 25059 3880 25091
rect 3912 25059 3952 25091
rect 3984 25059 4024 25091
rect 4056 25059 4096 25091
rect 4128 25059 4168 25091
rect 4200 25059 4240 25091
rect 4272 25059 4312 25091
rect 4344 25059 4384 25091
rect 4416 25059 4456 25091
rect 4488 25059 4528 25091
rect 4560 25059 4600 25091
rect 4632 25059 4672 25091
rect 4704 25059 4744 25091
rect 4776 25059 4816 25091
rect 4848 25059 4888 25091
rect 4920 25059 4960 25091
rect 4992 25059 5032 25091
rect 5064 25059 5104 25091
rect 5136 25059 5176 25091
rect 5208 25059 5248 25091
rect 5280 25059 5320 25091
rect 5352 25059 5392 25091
rect 5424 25059 5464 25091
rect 5496 25059 5536 25091
rect 5568 25059 5608 25091
rect 5640 25059 5680 25091
rect 5712 25059 5752 25091
rect 5784 25059 5824 25091
rect 5856 25059 5896 25091
rect 5928 25059 5968 25091
rect 6000 25059 6040 25091
rect 6072 25059 6112 25091
rect 6144 25059 6184 25091
rect 6216 25059 6256 25091
rect 6288 25059 6328 25091
rect 6360 25059 6400 25091
rect 6432 25059 6472 25091
rect 6504 25059 6544 25091
rect 6576 25059 6616 25091
rect 6648 25059 6688 25091
rect 6720 25059 6760 25091
rect 6792 25059 6832 25091
rect 6864 25059 6904 25091
rect 6936 25059 6976 25091
rect 7008 25059 7048 25091
rect 7080 25059 7120 25091
rect 7152 25059 7192 25091
rect 7224 25059 7264 25091
rect 7296 25059 7336 25091
rect 7368 25059 7408 25091
rect 7440 25059 7480 25091
rect 7512 25059 7552 25091
rect 7584 25059 7624 25091
rect 7656 25059 7696 25091
rect 7728 25059 7768 25091
rect 7800 25059 7840 25091
rect 7872 25059 7912 25091
rect 7944 25059 7984 25091
rect 8016 25059 8056 25091
rect 8088 25059 8128 25091
rect 8160 25059 8200 25091
rect 8232 25059 8272 25091
rect 8304 25059 8344 25091
rect 8376 25059 8416 25091
rect 8448 25059 8488 25091
rect 8520 25059 8560 25091
rect 8592 25059 8632 25091
rect 8664 25059 8704 25091
rect 8736 25059 8776 25091
rect 8808 25059 8848 25091
rect 8880 25059 8920 25091
rect 8952 25059 8992 25091
rect 9024 25059 9064 25091
rect 9096 25059 9136 25091
rect 9168 25059 9208 25091
rect 9240 25059 9280 25091
rect 9312 25059 9352 25091
rect 9384 25059 9424 25091
rect 9456 25059 9496 25091
rect 9528 25059 9568 25091
rect 9600 25059 9640 25091
rect 9672 25059 9712 25091
rect 9744 25059 9784 25091
rect 9816 25059 9856 25091
rect 9888 25059 9928 25091
rect 9960 25059 10000 25091
rect 10032 25059 10072 25091
rect 10104 25059 10144 25091
rect 10176 25059 10216 25091
rect 10248 25059 10288 25091
rect 10320 25059 10360 25091
rect 10392 25059 10432 25091
rect 10464 25059 10504 25091
rect 10536 25059 10576 25091
rect 10608 25059 10648 25091
rect 10680 25059 10720 25091
rect 10752 25059 10792 25091
rect 10824 25059 10864 25091
rect 10896 25059 10936 25091
rect 10968 25059 11008 25091
rect 11040 25059 11080 25091
rect 11112 25059 11152 25091
rect 11184 25059 11224 25091
rect 11256 25059 11296 25091
rect 11328 25059 11368 25091
rect 11400 25059 11440 25091
rect 11472 25059 11512 25091
rect 11544 25059 11584 25091
rect 11616 25059 11656 25091
rect 11688 25059 11728 25091
rect 11760 25059 11800 25091
rect 11832 25059 11872 25091
rect 11904 25059 11944 25091
rect 11976 25059 12016 25091
rect 12048 25059 12088 25091
rect 12120 25059 12160 25091
rect 12192 25059 12232 25091
rect 12264 25059 12304 25091
rect 12336 25059 12376 25091
rect 12408 25059 12448 25091
rect 12480 25059 12520 25091
rect 12552 25059 12592 25091
rect 12624 25059 12664 25091
rect 12696 25059 12736 25091
rect 12768 25059 12808 25091
rect 12840 25059 12880 25091
rect 12912 25059 12952 25091
rect 12984 25059 13024 25091
rect 13056 25059 13096 25091
rect 13128 25059 13168 25091
rect 13200 25059 13240 25091
rect 13272 25059 13312 25091
rect 13344 25059 13384 25091
rect 13416 25059 13456 25091
rect 13488 25059 13528 25091
rect 13560 25059 13600 25091
rect 13632 25059 13672 25091
rect 13704 25059 13744 25091
rect 13776 25059 13816 25091
rect 13848 25059 13888 25091
rect 13920 25059 13960 25091
rect 13992 25059 14032 25091
rect 14064 25059 14104 25091
rect 14136 25059 14176 25091
rect 14208 25059 14248 25091
rect 14280 25059 14320 25091
rect 14352 25059 14392 25091
rect 14424 25059 14464 25091
rect 14496 25059 14536 25091
rect 14568 25059 14608 25091
rect 14640 25059 14680 25091
rect 14712 25059 14752 25091
rect 14784 25059 14824 25091
rect 14856 25059 14896 25091
rect 14928 25059 14968 25091
rect 15000 25059 15040 25091
rect 15072 25059 15112 25091
rect 15144 25059 15184 25091
rect 15216 25059 15256 25091
rect 15288 25059 15328 25091
rect 15360 25059 15400 25091
rect 15432 25059 15472 25091
rect 15504 25059 15544 25091
rect 15576 25059 15616 25091
rect 15648 25059 15688 25091
rect 15720 25059 15760 25091
rect 15792 25059 15832 25091
rect 15864 25059 15904 25091
rect 15936 25059 16000 25091
rect 0 25019 16000 25059
rect 0 24987 64 25019
rect 96 24987 136 25019
rect 168 24987 208 25019
rect 240 24987 280 25019
rect 312 24987 352 25019
rect 384 24987 424 25019
rect 456 24987 496 25019
rect 528 24987 568 25019
rect 600 24987 640 25019
rect 672 24987 712 25019
rect 744 24987 784 25019
rect 816 24987 856 25019
rect 888 24987 928 25019
rect 960 24987 1000 25019
rect 1032 24987 1072 25019
rect 1104 24987 1144 25019
rect 1176 24987 1216 25019
rect 1248 24987 1288 25019
rect 1320 24987 1360 25019
rect 1392 24987 1432 25019
rect 1464 24987 1504 25019
rect 1536 24987 1576 25019
rect 1608 24987 1648 25019
rect 1680 24987 1720 25019
rect 1752 24987 1792 25019
rect 1824 24987 1864 25019
rect 1896 24987 1936 25019
rect 1968 24987 2008 25019
rect 2040 24987 2080 25019
rect 2112 24987 2152 25019
rect 2184 24987 2224 25019
rect 2256 24987 2296 25019
rect 2328 24987 2368 25019
rect 2400 24987 2440 25019
rect 2472 24987 2512 25019
rect 2544 24987 2584 25019
rect 2616 24987 2656 25019
rect 2688 24987 2728 25019
rect 2760 24987 2800 25019
rect 2832 24987 2872 25019
rect 2904 24987 2944 25019
rect 2976 24987 3016 25019
rect 3048 24987 3088 25019
rect 3120 24987 3160 25019
rect 3192 24987 3232 25019
rect 3264 24987 3304 25019
rect 3336 24987 3376 25019
rect 3408 24987 3448 25019
rect 3480 24987 3520 25019
rect 3552 24987 3592 25019
rect 3624 24987 3664 25019
rect 3696 24987 3736 25019
rect 3768 24987 3808 25019
rect 3840 24987 3880 25019
rect 3912 24987 3952 25019
rect 3984 24987 4024 25019
rect 4056 24987 4096 25019
rect 4128 24987 4168 25019
rect 4200 24987 4240 25019
rect 4272 24987 4312 25019
rect 4344 24987 4384 25019
rect 4416 24987 4456 25019
rect 4488 24987 4528 25019
rect 4560 24987 4600 25019
rect 4632 24987 4672 25019
rect 4704 24987 4744 25019
rect 4776 24987 4816 25019
rect 4848 24987 4888 25019
rect 4920 24987 4960 25019
rect 4992 24987 5032 25019
rect 5064 24987 5104 25019
rect 5136 24987 5176 25019
rect 5208 24987 5248 25019
rect 5280 24987 5320 25019
rect 5352 24987 5392 25019
rect 5424 24987 5464 25019
rect 5496 24987 5536 25019
rect 5568 24987 5608 25019
rect 5640 24987 5680 25019
rect 5712 24987 5752 25019
rect 5784 24987 5824 25019
rect 5856 24987 5896 25019
rect 5928 24987 5968 25019
rect 6000 24987 6040 25019
rect 6072 24987 6112 25019
rect 6144 24987 6184 25019
rect 6216 24987 6256 25019
rect 6288 24987 6328 25019
rect 6360 24987 6400 25019
rect 6432 24987 6472 25019
rect 6504 24987 6544 25019
rect 6576 24987 6616 25019
rect 6648 24987 6688 25019
rect 6720 24987 6760 25019
rect 6792 24987 6832 25019
rect 6864 24987 6904 25019
rect 6936 24987 6976 25019
rect 7008 24987 7048 25019
rect 7080 24987 7120 25019
rect 7152 24987 7192 25019
rect 7224 24987 7264 25019
rect 7296 24987 7336 25019
rect 7368 24987 7408 25019
rect 7440 24987 7480 25019
rect 7512 24987 7552 25019
rect 7584 24987 7624 25019
rect 7656 24987 7696 25019
rect 7728 24987 7768 25019
rect 7800 24987 7840 25019
rect 7872 24987 7912 25019
rect 7944 24987 7984 25019
rect 8016 24987 8056 25019
rect 8088 24987 8128 25019
rect 8160 24987 8200 25019
rect 8232 24987 8272 25019
rect 8304 24987 8344 25019
rect 8376 24987 8416 25019
rect 8448 24987 8488 25019
rect 8520 24987 8560 25019
rect 8592 24987 8632 25019
rect 8664 24987 8704 25019
rect 8736 24987 8776 25019
rect 8808 24987 8848 25019
rect 8880 24987 8920 25019
rect 8952 24987 8992 25019
rect 9024 24987 9064 25019
rect 9096 24987 9136 25019
rect 9168 24987 9208 25019
rect 9240 24987 9280 25019
rect 9312 24987 9352 25019
rect 9384 24987 9424 25019
rect 9456 24987 9496 25019
rect 9528 24987 9568 25019
rect 9600 24987 9640 25019
rect 9672 24987 9712 25019
rect 9744 24987 9784 25019
rect 9816 24987 9856 25019
rect 9888 24987 9928 25019
rect 9960 24987 10000 25019
rect 10032 24987 10072 25019
rect 10104 24987 10144 25019
rect 10176 24987 10216 25019
rect 10248 24987 10288 25019
rect 10320 24987 10360 25019
rect 10392 24987 10432 25019
rect 10464 24987 10504 25019
rect 10536 24987 10576 25019
rect 10608 24987 10648 25019
rect 10680 24987 10720 25019
rect 10752 24987 10792 25019
rect 10824 24987 10864 25019
rect 10896 24987 10936 25019
rect 10968 24987 11008 25019
rect 11040 24987 11080 25019
rect 11112 24987 11152 25019
rect 11184 24987 11224 25019
rect 11256 24987 11296 25019
rect 11328 24987 11368 25019
rect 11400 24987 11440 25019
rect 11472 24987 11512 25019
rect 11544 24987 11584 25019
rect 11616 24987 11656 25019
rect 11688 24987 11728 25019
rect 11760 24987 11800 25019
rect 11832 24987 11872 25019
rect 11904 24987 11944 25019
rect 11976 24987 12016 25019
rect 12048 24987 12088 25019
rect 12120 24987 12160 25019
rect 12192 24987 12232 25019
rect 12264 24987 12304 25019
rect 12336 24987 12376 25019
rect 12408 24987 12448 25019
rect 12480 24987 12520 25019
rect 12552 24987 12592 25019
rect 12624 24987 12664 25019
rect 12696 24987 12736 25019
rect 12768 24987 12808 25019
rect 12840 24987 12880 25019
rect 12912 24987 12952 25019
rect 12984 24987 13024 25019
rect 13056 24987 13096 25019
rect 13128 24987 13168 25019
rect 13200 24987 13240 25019
rect 13272 24987 13312 25019
rect 13344 24987 13384 25019
rect 13416 24987 13456 25019
rect 13488 24987 13528 25019
rect 13560 24987 13600 25019
rect 13632 24987 13672 25019
rect 13704 24987 13744 25019
rect 13776 24987 13816 25019
rect 13848 24987 13888 25019
rect 13920 24987 13960 25019
rect 13992 24987 14032 25019
rect 14064 24987 14104 25019
rect 14136 24987 14176 25019
rect 14208 24987 14248 25019
rect 14280 24987 14320 25019
rect 14352 24987 14392 25019
rect 14424 24987 14464 25019
rect 14496 24987 14536 25019
rect 14568 24987 14608 25019
rect 14640 24987 14680 25019
rect 14712 24987 14752 25019
rect 14784 24987 14824 25019
rect 14856 24987 14896 25019
rect 14928 24987 14968 25019
rect 15000 24987 15040 25019
rect 15072 24987 15112 25019
rect 15144 24987 15184 25019
rect 15216 24987 15256 25019
rect 15288 24987 15328 25019
rect 15360 24987 15400 25019
rect 15432 24987 15472 25019
rect 15504 24987 15544 25019
rect 15576 24987 15616 25019
rect 15648 24987 15688 25019
rect 15720 24987 15760 25019
rect 15792 24987 15832 25019
rect 15864 24987 15904 25019
rect 15936 24987 16000 25019
rect 0 24947 16000 24987
rect 0 24915 64 24947
rect 96 24915 136 24947
rect 168 24915 208 24947
rect 240 24915 280 24947
rect 312 24915 352 24947
rect 384 24915 424 24947
rect 456 24915 496 24947
rect 528 24915 568 24947
rect 600 24915 640 24947
rect 672 24915 712 24947
rect 744 24915 784 24947
rect 816 24915 856 24947
rect 888 24915 928 24947
rect 960 24915 1000 24947
rect 1032 24915 1072 24947
rect 1104 24915 1144 24947
rect 1176 24915 1216 24947
rect 1248 24915 1288 24947
rect 1320 24915 1360 24947
rect 1392 24915 1432 24947
rect 1464 24915 1504 24947
rect 1536 24915 1576 24947
rect 1608 24915 1648 24947
rect 1680 24915 1720 24947
rect 1752 24915 1792 24947
rect 1824 24915 1864 24947
rect 1896 24915 1936 24947
rect 1968 24915 2008 24947
rect 2040 24915 2080 24947
rect 2112 24915 2152 24947
rect 2184 24915 2224 24947
rect 2256 24915 2296 24947
rect 2328 24915 2368 24947
rect 2400 24915 2440 24947
rect 2472 24915 2512 24947
rect 2544 24915 2584 24947
rect 2616 24915 2656 24947
rect 2688 24915 2728 24947
rect 2760 24915 2800 24947
rect 2832 24915 2872 24947
rect 2904 24915 2944 24947
rect 2976 24915 3016 24947
rect 3048 24915 3088 24947
rect 3120 24915 3160 24947
rect 3192 24915 3232 24947
rect 3264 24915 3304 24947
rect 3336 24915 3376 24947
rect 3408 24915 3448 24947
rect 3480 24915 3520 24947
rect 3552 24915 3592 24947
rect 3624 24915 3664 24947
rect 3696 24915 3736 24947
rect 3768 24915 3808 24947
rect 3840 24915 3880 24947
rect 3912 24915 3952 24947
rect 3984 24915 4024 24947
rect 4056 24915 4096 24947
rect 4128 24915 4168 24947
rect 4200 24915 4240 24947
rect 4272 24915 4312 24947
rect 4344 24915 4384 24947
rect 4416 24915 4456 24947
rect 4488 24915 4528 24947
rect 4560 24915 4600 24947
rect 4632 24915 4672 24947
rect 4704 24915 4744 24947
rect 4776 24915 4816 24947
rect 4848 24915 4888 24947
rect 4920 24915 4960 24947
rect 4992 24915 5032 24947
rect 5064 24915 5104 24947
rect 5136 24915 5176 24947
rect 5208 24915 5248 24947
rect 5280 24915 5320 24947
rect 5352 24915 5392 24947
rect 5424 24915 5464 24947
rect 5496 24915 5536 24947
rect 5568 24915 5608 24947
rect 5640 24915 5680 24947
rect 5712 24915 5752 24947
rect 5784 24915 5824 24947
rect 5856 24915 5896 24947
rect 5928 24915 5968 24947
rect 6000 24915 6040 24947
rect 6072 24915 6112 24947
rect 6144 24915 6184 24947
rect 6216 24915 6256 24947
rect 6288 24915 6328 24947
rect 6360 24915 6400 24947
rect 6432 24915 6472 24947
rect 6504 24915 6544 24947
rect 6576 24915 6616 24947
rect 6648 24915 6688 24947
rect 6720 24915 6760 24947
rect 6792 24915 6832 24947
rect 6864 24915 6904 24947
rect 6936 24915 6976 24947
rect 7008 24915 7048 24947
rect 7080 24915 7120 24947
rect 7152 24915 7192 24947
rect 7224 24915 7264 24947
rect 7296 24915 7336 24947
rect 7368 24915 7408 24947
rect 7440 24915 7480 24947
rect 7512 24915 7552 24947
rect 7584 24915 7624 24947
rect 7656 24915 7696 24947
rect 7728 24915 7768 24947
rect 7800 24915 7840 24947
rect 7872 24915 7912 24947
rect 7944 24915 7984 24947
rect 8016 24915 8056 24947
rect 8088 24915 8128 24947
rect 8160 24915 8200 24947
rect 8232 24915 8272 24947
rect 8304 24915 8344 24947
rect 8376 24915 8416 24947
rect 8448 24915 8488 24947
rect 8520 24915 8560 24947
rect 8592 24915 8632 24947
rect 8664 24915 8704 24947
rect 8736 24915 8776 24947
rect 8808 24915 8848 24947
rect 8880 24915 8920 24947
rect 8952 24915 8992 24947
rect 9024 24915 9064 24947
rect 9096 24915 9136 24947
rect 9168 24915 9208 24947
rect 9240 24915 9280 24947
rect 9312 24915 9352 24947
rect 9384 24915 9424 24947
rect 9456 24915 9496 24947
rect 9528 24915 9568 24947
rect 9600 24915 9640 24947
rect 9672 24915 9712 24947
rect 9744 24915 9784 24947
rect 9816 24915 9856 24947
rect 9888 24915 9928 24947
rect 9960 24915 10000 24947
rect 10032 24915 10072 24947
rect 10104 24915 10144 24947
rect 10176 24915 10216 24947
rect 10248 24915 10288 24947
rect 10320 24915 10360 24947
rect 10392 24915 10432 24947
rect 10464 24915 10504 24947
rect 10536 24915 10576 24947
rect 10608 24915 10648 24947
rect 10680 24915 10720 24947
rect 10752 24915 10792 24947
rect 10824 24915 10864 24947
rect 10896 24915 10936 24947
rect 10968 24915 11008 24947
rect 11040 24915 11080 24947
rect 11112 24915 11152 24947
rect 11184 24915 11224 24947
rect 11256 24915 11296 24947
rect 11328 24915 11368 24947
rect 11400 24915 11440 24947
rect 11472 24915 11512 24947
rect 11544 24915 11584 24947
rect 11616 24915 11656 24947
rect 11688 24915 11728 24947
rect 11760 24915 11800 24947
rect 11832 24915 11872 24947
rect 11904 24915 11944 24947
rect 11976 24915 12016 24947
rect 12048 24915 12088 24947
rect 12120 24915 12160 24947
rect 12192 24915 12232 24947
rect 12264 24915 12304 24947
rect 12336 24915 12376 24947
rect 12408 24915 12448 24947
rect 12480 24915 12520 24947
rect 12552 24915 12592 24947
rect 12624 24915 12664 24947
rect 12696 24915 12736 24947
rect 12768 24915 12808 24947
rect 12840 24915 12880 24947
rect 12912 24915 12952 24947
rect 12984 24915 13024 24947
rect 13056 24915 13096 24947
rect 13128 24915 13168 24947
rect 13200 24915 13240 24947
rect 13272 24915 13312 24947
rect 13344 24915 13384 24947
rect 13416 24915 13456 24947
rect 13488 24915 13528 24947
rect 13560 24915 13600 24947
rect 13632 24915 13672 24947
rect 13704 24915 13744 24947
rect 13776 24915 13816 24947
rect 13848 24915 13888 24947
rect 13920 24915 13960 24947
rect 13992 24915 14032 24947
rect 14064 24915 14104 24947
rect 14136 24915 14176 24947
rect 14208 24915 14248 24947
rect 14280 24915 14320 24947
rect 14352 24915 14392 24947
rect 14424 24915 14464 24947
rect 14496 24915 14536 24947
rect 14568 24915 14608 24947
rect 14640 24915 14680 24947
rect 14712 24915 14752 24947
rect 14784 24915 14824 24947
rect 14856 24915 14896 24947
rect 14928 24915 14968 24947
rect 15000 24915 15040 24947
rect 15072 24915 15112 24947
rect 15144 24915 15184 24947
rect 15216 24915 15256 24947
rect 15288 24915 15328 24947
rect 15360 24915 15400 24947
rect 15432 24915 15472 24947
rect 15504 24915 15544 24947
rect 15576 24915 15616 24947
rect 15648 24915 15688 24947
rect 15720 24915 15760 24947
rect 15792 24915 15832 24947
rect 15864 24915 15904 24947
rect 15936 24915 16000 24947
rect 0 24875 16000 24915
rect 0 24843 64 24875
rect 96 24843 136 24875
rect 168 24843 208 24875
rect 240 24843 280 24875
rect 312 24843 352 24875
rect 384 24843 424 24875
rect 456 24843 496 24875
rect 528 24843 568 24875
rect 600 24843 640 24875
rect 672 24843 712 24875
rect 744 24843 784 24875
rect 816 24843 856 24875
rect 888 24843 928 24875
rect 960 24843 1000 24875
rect 1032 24843 1072 24875
rect 1104 24843 1144 24875
rect 1176 24843 1216 24875
rect 1248 24843 1288 24875
rect 1320 24843 1360 24875
rect 1392 24843 1432 24875
rect 1464 24843 1504 24875
rect 1536 24843 1576 24875
rect 1608 24843 1648 24875
rect 1680 24843 1720 24875
rect 1752 24843 1792 24875
rect 1824 24843 1864 24875
rect 1896 24843 1936 24875
rect 1968 24843 2008 24875
rect 2040 24843 2080 24875
rect 2112 24843 2152 24875
rect 2184 24843 2224 24875
rect 2256 24843 2296 24875
rect 2328 24843 2368 24875
rect 2400 24843 2440 24875
rect 2472 24843 2512 24875
rect 2544 24843 2584 24875
rect 2616 24843 2656 24875
rect 2688 24843 2728 24875
rect 2760 24843 2800 24875
rect 2832 24843 2872 24875
rect 2904 24843 2944 24875
rect 2976 24843 3016 24875
rect 3048 24843 3088 24875
rect 3120 24843 3160 24875
rect 3192 24843 3232 24875
rect 3264 24843 3304 24875
rect 3336 24843 3376 24875
rect 3408 24843 3448 24875
rect 3480 24843 3520 24875
rect 3552 24843 3592 24875
rect 3624 24843 3664 24875
rect 3696 24843 3736 24875
rect 3768 24843 3808 24875
rect 3840 24843 3880 24875
rect 3912 24843 3952 24875
rect 3984 24843 4024 24875
rect 4056 24843 4096 24875
rect 4128 24843 4168 24875
rect 4200 24843 4240 24875
rect 4272 24843 4312 24875
rect 4344 24843 4384 24875
rect 4416 24843 4456 24875
rect 4488 24843 4528 24875
rect 4560 24843 4600 24875
rect 4632 24843 4672 24875
rect 4704 24843 4744 24875
rect 4776 24843 4816 24875
rect 4848 24843 4888 24875
rect 4920 24843 4960 24875
rect 4992 24843 5032 24875
rect 5064 24843 5104 24875
rect 5136 24843 5176 24875
rect 5208 24843 5248 24875
rect 5280 24843 5320 24875
rect 5352 24843 5392 24875
rect 5424 24843 5464 24875
rect 5496 24843 5536 24875
rect 5568 24843 5608 24875
rect 5640 24843 5680 24875
rect 5712 24843 5752 24875
rect 5784 24843 5824 24875
rect 5856 24843 5896 24875
rect 5928 24843 5968 24875
rect 6000 24843 6040 24875
rect 6072 24843 6112 24875
rect 6144 24843 6184 24875
rect 6216 24843 6256 24875
rect 6288 24843 6328 24875
rect 6360 24843 6400 24875
rect 6432 24843 6472 24875
rect 6504 24843 6544 24875
rect 6576 24843 6616 24875
rect 6648 24843 6688 24875
rect 6720 24843 6760 24875
rect 6792 24843 6832 24875
rect 6864 24843 6904 24875
rect 6936 24843 6976 24875
rect 7008 24843 7048 24875
rect 7080 24843 7120 24875
rect 7152 24843 7192 24875
rect 7224 24843 7264 24875
rect 7296 24843 7336 24875
rect 7368 24843 7408 24875
rect 7440 24843 7480 24875
rect 7512 24843 7552 24875
rect 7584 24843 7624 24875
rect 7656 24843 7696 24875
rect 7728 24843 7768 24875
rect 7800 24843 7840 24875
rect 7872 24843 7912 24875
rect 7944 24843 7984 24875
rect 8016 24843 8056 24875
rect 8088 24843 8128 24875
rect 8160 24843 8200 24875
rect 8232 24843 8272 24875
rect 8304 24843 8344 24875
rect 8376 24843 8416 24875
rect 8448 24843 8488 24875
rect 8520 24843 8560 24875
rect 8592 24843 8632 24875
rect 8664 24843 8704 24875
rect 8736 24843 8776 24875
rect 8808 24843 8848 24875
rect 8880 24843 8920 24875
rect 8952 24843 8992 24875
rect 9024 24843 9064 24875
rect 9096 24843 9136 24875
rect 9168 24843 9208 24875
rect 9240 24843 9280 24875
rect 9312 24843 9352 24875
rect 9384 24843 9424 24875
rect 9456 24843 9496 24875
rect 9528 24843 9568 24875
rect 9600 24843 9640 24875
rect 9672 24843 9712 24875
rect 9744 24843 9784 24875
rect 9816 24843 9856 24875
rect 9888 24843 9928 24875
rect 9960 24843 10000 24875
rect 10032 24843 10072 24875
rect 10104 24843 10144 24875
rect 10176 24843 10216 24875
rect 10248 24843 10288 24875
rect 10320 24843 10360 24875
rect 10392 24843 10432 24875
rect 10464 24843 10504 24875
rect 10536 24843 10576 24875
rect 10608 24843 10648 24875
rect 10680 24843 10720 24875
rect 10752 24843 10792 24875
rect 10824 24843 10864 24875
rect 10896 24843 10936 24875
rect 10968 24843 11008 24875
rect 11040 24843 11080 24875
rect 11112 24843 11152 24875
rect 11184 24843 11224 24875
rect 11256 24843 11296 24875
rect 11328 24843 11368 24875
rect 11400 24843 11440 24875
rect 11472 24843 11512 24875
rect 11544 24843 11584 24875
rect 11616 24843 11656 24875
rect 11688 24843 11728 24875
rect 11760 24843 11800 24875
rect 11832 24843 11872 24875
rect 11904 24843 11944 24875
rect 11976 24843 12016 24875
rect 12048 24843 12088 24875
rect 12120 24843 12160 24875
rect 12192 24843 12232 24875
rect 12264 24843 12304 24875
rect 12336 24843 12376 24875
rect 12408 24843 12448 24875
rect 12480 24843 12520 24875
rect 12552 24843 12592 24875
rect 12624 24843 12664 24875
rect 12696 24843 12736 24875
rect 12768 24843 12808 24875
rect 12840 24843 12880 24875
rect 12912 24843 12952 24875
rect 12984 24843 13024 24875
rect 13056 24843 13096 24875
rect 13128 24843 13168 24875
rect 13200 24843 13240 24875
rect 13272 24843 13312 24875
rect 13344 24843 13384 24875
rect 13416 24843 13456 24875
rect 13488 24843 13528 24875
rect 13560 24843 13600 24875
rect 13632 24843 13672 24875
rect 13704 24843 13744 24875
rect 13776 24843 13816 24875
rect 13848 24843 13888 24875
rect 13920 24843 13960 24875
rect 13992 24843 14032 24875
rect 14064 24843 14104 24875
rect 14136 24843 14176 24875
rect 14208 24843 14248 24875
rect 14280 24843 14320 24875
rect 14352 24843 14392 24875
rect 14424 24843 14464 24875
rect 14496 24843 14536 24875
rect 14568 24843 14608 24875
rect 14640 24843 14680 24875
rect 14712 24843 14752 24875
rect 14784 24843 14824 24875
rect 14856 24843 14896 24875
rect 14928 24843 14968 24875
rect 15000 24843 15040 24875
rect 15072 24843 15112 24875
rect 15144 24843 15184 24875
rect 15216 24843 15256 24875
rect 15288 24843 15328 24875
rect 15360 24843 15400 24875
rect 15432 24843 15472 24875
rect 15504 24843 15544 24875
rect 15576 24843 15616 24875
rect 15648 24843 15688 24875
rect 15720 24843 15760 24875
rect 15792 24843 15832 24875
rect 15864 24843 15904 24875
rect 15936 24843 16000 24875
rect 0 24803 16000 24843
rect 0 24771 64 24803
rect 96 24771 136 24803
rect 168 24771 208 24803
rect 240 24771 280 24803
rect 312 24771 352 24803
rect 384 24771 424 24803
rect 456 24771 496 24803
rect 528 24771 568 24803
rect 600 24771 640 24803
rect 672 24771 712 24803
rect 744 24771 784 24803
rect 816 24771 856 24803
rect 888 24771 928 24803
rect 960 24771 1000 24803
rect 1032 24771 1072 24803
rect 1104 24771 1144 24803
rect 1176 24771 1216 24803
rect 1248 24771 1288 24803
rect 1320 24771 1360 24803
rect 1392 24771 1432 24803
rect 1464 24771 1504 24803
rect 1536 24771 1576 24803
rect 1608 24771 1648 24803
rect 1680 24771 1720 24803
rect 1752 24771 1792 24803
rect 1824 24771 1864 24803
rect 1896 24771 1936 24803
rect 1968 24771 2008 24803
rect 2040 24771 2080 24803
rect 2112 24771 2152 24803
rect 2184 24771 2224 24803
rect 2256 24771 2296 24803
rect 2328 24771 2368 24803
rect 2400 24771 2440 24803
rect 2472 24771 2512 24803
rect 2544 24771 2584 24803
rect 2616 24771 2656 24803
rect 2688 24771 2728 24803
rect 2760 24771 2800 24803
rect 2832 24771 2872 24803
rect 2904 24771 2944 24803
rect 2976 24771 3016 24803
rect 3048 24771 3088 24803
rect 3120 24771 3160 24803
rect 3192 24771 3232 24803
rect 3264 24771 3304 24803
rect 3336 24771 3376 24803
rect 3408 24771 3448 24803
rect 3480 24771 3520 24803
rect 3552 24771 3592 24803
rect 3624 24771 3664 24803
rect 3696 24771 3736 24803
rect 3768 24771 3808 24803
rect 3840 24771 3880 24803
rect 3912 24771 3952 24803
rect 3984 24771 4024 24803
rect 4056 24771 4096 24803
rect 4128 24771 4168 24803
rect 4200 24771 4240 24803
rect 4272 24771 4312 24803
rect 4344 24771 4384 24803
rect 4416 24771 4456 24803
rect 4488 24771 4528 24803
rect 4560 24771 4600 24803
rect 4632 24771 4672 24803
rect 4704 24771 4744 24803
rect 4776 24771 4816 24803
rect 4848 24771 4888 24803
rect 4920 24771 4960 24803
rect 4992 24771 5032 24803
rect 5064 24771 5104 24803
rect 5136 24771 5176 24803
rect 5208 24771 5248 24803
rect 5280 24771 5320 24803
rect 5352 24771 5392 24803
rect 5424 24771 5464 24803
rect 5496 24771 5536 24803
rect 5568 24771 5608 24803
rect 5640 24771 5680 24803
rect 5712 24771 5752 24803
rect 5784 24771 5824 24803
rect 5856 24771 5896 24803
rect 5928 24771 5968 24803
rect 6000 24771 6040 24803
rect 6072 24771 6112 24803
rect 6144 24771 6184 24803
rect 6216 24771 6256 24803
rect 6288 24771 6328 24803
rect 6360 24771 6400 24803
rect 6432 24771 6472 24803
rect 6504 24771 6544 24803
rect 6576 24771 6616 24803
rect 6648 24771 6688 24803
rect 6720 24771 6760 24803
rect 6792 24771 6832 24803
rect 6864 24771 6904 24803
rect 6936 24771 6976 24803
rect 7008 24771 7048 24803
rect 7080 24771 7120 24803
rect 7152 24771 7192 24803
rect 7224 24771 7264 24803
rect 7296 24771 7336 24803
rect 7368 24771 7408 24803
rect 7440 24771 7480 24803
rect 7512 24771 7552 24803
rect 7584 24771 7624 24803
rect 7656 24771 7696 24803
rect 7728 24771 7768 24803
rect 7800 24771 7840 24803
rect 7872 24771 7912 24803
rect 7944 24771 7984 24803
rect 8016 24771 8056 24803
rect 8088 24771 8128 24803
rect 8160 24771 8200 24803
rect 8232 24771 8272 24803
rect 8304 24771 8344 24803
rect 8376 24771 8416 24803
rect 8448 24771 8488 24803
rect 8520 24771 8560 24803
rect 8592 24771 8632 24803
rect 8664 24771 8704 24803
rect 8736 24771 8776 24803
rect 8808 24771 8848 24803
rect 8880 24771 8920 24803
rect 8952 24771 8992 24803
rect 9024 24771 9064 24803
rect 9096 24771 9136 24803
rect 9168 24771 9208 24803
rect 9240 24771 9280 24803
rect 9312 24771 9352 24803
rect 9384 24771 9424 24803
rect 9456 24771 9496 24803
rect 9528 24771 9568 24803
rect 9600 24771 9640 24803
rect 9672 24771 9712 24803
rect 9744 24771 9784 24803
rect 9816 24771 9856 24803
rect 9888 24771 9928 24803
rect 9960 24771 10000 24803
rect 10032 24771 10072 24803
rect 10104 24771 10144 24803
rect 10176 24771 10216 24803
rect 10248 24771 10288 24803
rect 10320 24771 10360 24803
rect 10392 24771 10432 24803
rect 10464 24771 10504 24803
rect 10536 24771 10576 24803
rect 10608 24771 10648 24803
rect 10680 24771 10720 24803
rect 10752 24771 10792 24803
rect 10824 24771 10864 24803
rect 10896 24771 10936 24803
rect 10968 24771 11008 24803
rect 11040 24771 11080 24803
rect 11112 24771 11152 24803
rect 11184 24771 11224 24803
rect 11256 24771 11296 24803
rect 11328 24771 11368 24803
rect 11400 24771 11440 24803
rect 11472 24771 11512 24803
rect 11544 24771 11584 24803
rect 11616 24771 11656 24803
rect 11688 24771 11728 24803
rect 11760 24771 11800 24803
rect 11832 24771 11872 24803
rect 11904 24771 11944 24803
rect 11976 24771 12016 24803
rect 12048 24771 12088 24803
rect 12120 24771 12160 24803
rect 12192 24771 12232 24803
rect 12264 24771 12304 24803
rect 12336 24771 12376 24803
rect 12408 24771 12448 24803
rect 12480 24771 12520 24803
rect 12552 24771 12592 24803
rect 12624 24771 12664 24803
rect 12696 24771 12736 24803
rect 12768 24771 12808 24803
rect 12840 24771 12880 24803
rect 12912 24771 12952 24803
rect 12984 24771 13024 24803
rect 13056 24771 13096 24803
rect 13128 24771 13168 24803
rect 13200 24771 13240 24803
rect 13272 24771 13312 24803
rect 13344 24771 13384 24803
rect 13416 24771 13456 24803
rect 13488 24771 13528 24803
rect 13560 24771 13600 24803
rect 13632 24771 13672 24803
rect 13704 24771 13744 24803
rect 13776 24771 13816 24803
rect 13848 24771 13888 24803
rect 13920 24771 13960 24803
rect 13992 24771 14032 24803
rect 14064 24771 14104 24803
rect 14136 24771 14176 24803
rect 14208 24771 14248 24803
rect 14280 24771 14320 24803
rect 14352 24771 14392 24803
rect 14424 24771 14464 24803
rect 14496 24771 14536 24803
rect 14568 24771 14608 24803
rect 14640 24771 14680 24803
rect 14712 24771 14752 24803
rect 14784 24771 14824 24803
rect 14856 24771 14896 24803
rect 14928 24771 14968 24803
rect 15000 24771 15040 24803
rect 15072 24771 15112 24803
rect 15144 24771 15184 24803
rect 15216 24771 15256 24803
rect 15288 24771 15328 24803
rect 15360 24771 15400 24803
rect 15432 24771 15472 24803
rect 15504 24771 15544 24803
rect 15576 24771 15616 24803
rect 15648 24771 15688 24803
rect 15720 24771 15760 24803
rect 15792 24771 15832 24803
rect 15864 24771 15904 24803
rect 15936 24771 16000 24803
rect 0 24731 16000 24771
rect 0 24699 64 24731
rect 96 24699 136 24731
rect 168 24699 208 24731
rect 240 24699 280 24731
rect 312 24699 352 24731
rect 384 24699 424 24731
rect 456 24699 496 24731
rect 528 24699 568 24731
rect 600 24699 640 24731
rect 672 24699 712 24731
rect 744 24699 784 24731
rect 816 24699 856 24731
rect 888 24699 928 24731
rect 960 24699 1000 24731
rect 1032 24699 1072 24731
rect 1104 24699 1144 24731
rect 1176 24699 1216 24731
rect 1248 24699 1288 24731
rect 1320 24699 1360 24731
rect 1392 24699 1432 24731
rect 1464 24699 1504 24731
rect 1536 24699 1576 24731
rect 1608 24699 1648 24731
rect 1680 24699 1720 24731
rect 1752 24699 1792 24731
rect 1824 24699 1864 24731
rect 1896 24699 1936 24731
rect 1968 24699 2008 24731
rect 2040 24699 2080 24731
rect 2112 24699 2152 24731
rect 2184 24699 2224 24731
rect 2256 24699 2296 24731
rect 2328 24699 2368 24731
rect 2400 24699 2440 24731
rect 2472 24699 2512 24731
rect 2544 24699 2584 24731
rect 2616 24699 2656 24731
rect 2688 24699 2728 24731
rect 2760 24699 2800 24731
rect 2832 24699 2872 24731
rect 2904 24699 2944 24731
rect 2976 24699 3016 24731
rect 3048 24699 3088 24731
rect 3120 24699 3160 24731
rect 3192 24699 3232 24731
rect 3264 24699 3304 24731
rect 3336 24699 3376 24731
rect 3408 24699 3448 24731
rect 3480 24699 3520 24731
rect 3552 24699 3592 24731
rect 3624 24699 3664 24731
rect 3696 24699 3736 24731
rect 3768 24699 3808 24731
rect 3840 24699 3880 24731
rect 3912 24699 3952 24731
rect 3984 24699 4024 24731
rect 4056 24699 4096 24731
rect 4128 24699 4168 24731
rect 4200 24699 4240 24731
rect 4272 24699 4312 24731
rect 4344 24699 4384 24731
rect 4416 24699 4456 24731
rect 4488 24699 4528 24731
rect 4560 24699 4600 24731
rect 4632 24699 4672 24731
rect 4704 24699 4744 24731
rect 4776 24699 4816 24731
rect 4848 24699 4888 24731
rect 4920 24699 4960 24731
rect 4992 24699 5032 24731
rect 5064 24699 5104 24731
rect 5136 24699 5176 24731
rect 5208 24699 5248 24731
rect 5280 24699 5320 24731
rect 5352 24699 5392 24731
rect 5424 24699 5464 24731
rect 5496 24699 5536 24731
rect 5568 24699 5608 24731
rect 5640 24699 5680 24731
rect 5712 24699 5752 24731
rect 5784 24699 5824 24731
rect 5856 24699 5896 24731
rect 5928 24699 5968 24731
rect 6000 24699 6040 24731
rect 6072 24699 6112 24731
rect 6144 24699 6184 24731
rect 6216 24699 6256 24731
rect 6288 24699 6328 24731
rect 6360 24699 6400 24731
rect 6432 24699 6472 24731
rect 6504 24699 6544 24731
rect 6576 24699 6616 24731
rect 6648 24699 6688 24731
rect 6720 24699 6760 24731
rect 6792 24699 6832 24731
rect 6864 24699 6904 24731
rect 6936 24699 6976 24731
rect 7008 24699 7048 24731
rect 7080 24699 7120 24731
rect 7152 24699 7192 24731
rect 7224 24699 7264 24731
rect 7296 24699 7336 24731
rect 7368 24699 7408 24731
rect 7440 24699 7480 24731
rect 7512 24699 7552 24731
rect 7584 24699 7624 24731
rect 7656 24699 7696 24731
rect 7728 24699 7768 24731
rect 7800 24699 7840 24731
rect 7872 24699 7912 24731
rect 7944 24699 7984 24731
rect 8016 24699 8056 24731
rect 8088 24699 8128 24731
rect 8160 24699 8200 24731
rect 8232 24699 8272 24731
rect 8304 24699 8344 24731
rect 8376 24699 8416 24731
rect 8448 24699 8488 24731
rect 8520 24699 8560 24731
rect 8592 24699 8632 24731
rect 8664 24699 8704 24731
rect 8736 24699 8776 24731
rect 8808 24699 8848 24731
rect 8880 24699 8920 24731
rect 8952 24699 8992 24731
rect 9024 24699 9064 24731
rect 9096 24699 9136 24731
rect 9168 24699 9208 24731
rect 9240 24699 9280 24731
rect 9312 24699 9352 24731
rect 9384 24699 9424 24731
rect 9456 24699 9496 24731
rect 9528 24699 9568 24731
rect 9600 24699 9640 24731
rect 9672 24699 9712 24731
rect 9744 24699 9784 24731
rect 9816 24699 9856 24731
rect 9888 24699 9928 24731
rect 9960 24699 10000 24731
rect 10032 24699 10072 24731
rect 10104 24699 10144 24731
rect 10176 24699 10216 24731
rect 10248 24699 10288 24731
rect 10320 24699 10360 24731
rect 10392 24699 10432 24731
rect 10464 24699 10504 24731
rect 10536 24699 10576 24731
rect 10608 24699 10648 24731
rect 10680 24699 10720 24731
rect 10752 24699 10792 24731
rect 10824 24699 10864 24731
rect 10896 24699 10936 24731
rect 10968 24699 11008 24731
rect 11040 24699 11080 24731
rect 11112 24699 11152 24731
rect 11184 24699 11224 24731
rect 11256 24699 11296 24731
rect 11328 24699 11368 24731
rect 11400 24699 11440 24731
rect 11472 24699 11512 24731
rect 11544 24699 11584 24731
rect 11616 24699 11656 24731
rect 11688 24699 11728 24731
rect 11760 24699 11800 24731
rect 11832 24699 11872 24731
rect 11904 24699 11944 24731
rect 11976 24699 12016 24731
rect 12048 24699 12088 24731
rect 12120 24699 12160 24731
rect 12192 24699 12232 24731
rect 12264 24699 12304 24731
rect 12336 24699 12376 24731
rect 12408 24699 12448 24731
rect 12480 24699 12520 24731
rect 12552 24699 12592 24731
rect 12624 24699 12664 24731
rect 12696 24699 12736 24731
rect 12768 24699 12808 24731
rect 12840 24699 12880 24731
rect 12912 24699 12952 24731
rect 12984 24699 13024 24731
rect 13056 24699 13096 24731
rect 13128 24699 13168 24731
rect 13200 24699 13240 24731
rect 13272 24699 13312 24731
rect 13344 24699 13384 24731
rect 13416 24699 13456 24731
rect 13488 24699 13528 24731
rect 13560 24699 13600 24731
rect 13632 24699 13672 24731
rect 13704 24699 13744 24731
rect 13776 24699 13816 24731
rect 13848 24699 13888 24731
rect 13920 24699 13960 24731
rect 13992 24699 14032 24731
rect 14064 24699 14104 24731
rect 14136 24699 14176 24731
rect 14208 24699 14248 24731
rect 14280 24699 14320 24731
rect 14352 24699 14392 24731
rect 14424 24699 14464 24731
rect 14496 24699 14536 24731
rect 14568 24699 14608 24731
rect 14640 24699 14680 24731
rect 14712 24699 14752 24731
rect 14784 24699 14824 24731
rect 14856 24699 14896 24731
rect 14928 24699 14968 24731
rect 15000 24699 15040 24731
rect 15072 24699 15112 24731
rect 15144 24699 15184 24731
rect 15216 24699 15256 24731
rect 15288 24699 15328 24731
rect 15360 24699 15400 24731
rect 15432 24699 15472 24731
rect 15504 24699 15544 24731
rect 15576 24699 15616 24731
rect 15648 24699 15688 24731
rect 15720 24699 15760 24731
rect 15792 24699 15832 24731
rect 15864 24699 15904 24731
rect 15936 24699 16000 24731
rect 0 24659 16000 24699
rect 0 24627 64 24659
rect 96 24627 136 24659
rect 168 24627 208 24659
rect 240 24627 280 24659
rect 312 24627 352 24659
rect 384 24627 424 24659
rect 456 24627 496 24659
rect 528 24627 568 24659
rect 600 24627 640 24659
rect 672 24627 712 24659
rect 744 24627 784 24659
rect 816 24627 856 24659
rect 888 24627 928 24659
rect 960 24627 1000 24659
rect 1032 24627 1072 24659
rect 1104 24627 1144 24659
rect 1176 24627 1216 24659
rect 1248 24627 1288 24659
rect 1320 24627 1360 24659
rect 1392 24627 1432 24659
rect 1464 24627 1504 24659
rect 1536 24627 1576 24659
rect 1608 24627 1648 24659
rect 1680 24627 1720 24659
rect 1752 24627 1792 24659
rect 1824 24627 1864 24659
rect 1896 24627 1936 24659
rect 1968 24627 2008 24659
rect 2040 24627 2080 24659
rect 2112 24627 2152 24659
rect 2184 24627 2224 24659
rect 2256 24627 2296 24659
rect 2328 24627 2368 24659
rect 2400 24627 2440 24659
rect 2472 24627 2512 24659
rect 2544 24627 2584 24659
rect 2616 24627 2656 24659
rect 2688 24627 2728 24659
rect 2760 24627 2800 24659
rect 2832 24627 2872 24659
rect 2904 24627 2944 24659
rect 2976 24627 3016 24659
rect 3048 24627 3088 24659
rect 3120 24627 3160 24659
rect 3192 24627 3232 24659
rect 3264 24627 3304 24659
rect 3336 24627 3376 24659
rect 3408 24627 3448 24659
rect 3480 24627 3520 24659
rect 3552 24627 3592 24659
rect 3624 24627 3664 24659
rect 3696 24627 3736 24659
rect 3768 24627 3808 24659
rect 3840 24627 3880 24659
rect 3912 24627 3952 24659
rect 3984 24627 4024 24659
rect 4056 24627 4096 24659
rect 4128 24627 4168 24659
rect 4200 24627 4240 24659
rect 4272 24627 4312 24659
rect 4344 24627 4384 24659
rect 4416 24627 4456 24659
rect 4488 24627 4528 24659
rect 4560 24627 4600 24659
rect 4632 24627 4672 24659
rect 4704 24627 4744 24659
rect 4776 24627 4816 24659
rect 4848 24627 4888 24659
rect 4920 24627 4960 24659
rect 4992 24627 5032 24659
rect 5064 24627 5104 24659
rect 5136 24627 5176 24659
rect 5208 24627 5248 24659
rect 5280 24627 5320 24659
rect 5352 24627 5392 24659
rect 5424 24627 5464 24659
rect 5496 24627 5536 24659
rect 5568 24627 5608 24659
rect 5640 24627 5680 24659
rect 5712 24627 5752 24659
rect 5784 24627 5824 24659
rect 5856 24627 5896 24659
rect 5928 24627 5968 24659
rect 6000 24627 6040 24659
rect 6072 24627 6112 24659
rect 6144 24627 6184 24659
rect 6216 24627 6256 24659
rect 6288 24627 6328 24659
rect 6360 24627 6400 24659
rect 6432 24627 6472 24659
rect 6504 24627 6544 24659
rect 6576 24627 6616 24659
rect 6648 24627 6688 24659
rect 6720 24627 6760 24659
rect 6792 24627 6832 24659
rect 6864 24627 6904 24659
rect 6936 24627 6976 24659
rect 7008 24627 7048 24659
rect 7080 24627 7120 24659
rect 7152 24627 7192 24659
rect 7224 24627 7264 24659
rect 7296 24627 7336 24659
rect 7368 24627 7408 24659
rect 7440 24627 7480 24659
rect 7512 24627 7552 24659
rect 7584 24627 7624 24659
rect 7656 24627 7696 24659
rect 7728 24627 7768 24659
rect 7800 24627 7840 24659
rect 7872 24627 7912 24659
rect 7944 24627 7984 24659
rect 8016 24627 8056 24659
rect 8088 24627 8128 24659
rect 8160 24627 8200 24659
rect 8232 24627 8272 24659
rect 8304 24627 8344 24659
rect 8376 24627 8416 24659
rect 8448 24627 8488 24659
rect 8520 24627 8560 24659
rect 8592 24627 8632 24659
rect 8664 24627 8704 24659
rect 8736 24627 8776 24659
rect 8808 24627 8848 24659
rect 8880 24627 8920 24659
rect 8952 24627 8992 24659
rect 9024 24627 9064 24659
rect 9096 24627 9136 24659
rect 9168 24627 9208 24659
rect 9240 24627 9280 24659
rect 9312 24627 9352 24659
rect 9384 24627 9424 24659
rect 9456 24627 9496 24659
rect 9528 24627 9568 24659
rect 9600 24627 9640 24659
rect 9672 24627 9712 24659
rect 9744 24627 9784 24659
rect 9816 24627 9856 24659
rect 9888 24627 9928 24659
rect 9960 24627 10000 24659
rect 10032 24627 10072 24659
rect 10104 24627 10144 24659
rect 10176 24627 10216 24659
rect 10248 24627 10288 24659
rect 10320 24627 10360 24659
rect 10392 24627 10432 24659
rect 10464 24627 10504 24659
rect 10536 24627 10576 24659
rect 10608 24627 10648 24659
rect 10680 24627 10720 24659
rect 10752 24627 10792 24659
rect 10824 24627 10864 24659
rect 10896 24627 10936 24659
rect 10968 24627 11008 24659
rect 11040 24627 11080 24659
rect 11112 24627 11152 24659
rect 11184 24627 11224 24659
rect 11256 24627 11296 24659
rect 11328 24627 11368 24659
rect 11400 24627 11440 24659
rect 11472 24627 11512 24659
rect 11544 24627 11584 24659
rect 11616 24627 11656 24659
rect 11688 24627 11728 24659
rect 11760 24627 11800 24659
rect 11832 24627 11872 24659
rect 11904 24627 11944 24659
rect 11976 24627 12016 24659
rect 12048 24627 12088 24659
rect 12120 24627 12160 24659
rect 12192 24627 12232 24659
rect 12264 24627 12304 24659
rect 12336 24627 12376 24659
rect 12408 24627 12448 24659
rect 12480 24627 12520 24659
rect 12552 24627 12592 24659
rect 12624 24627 12664 24659
rect 12696 24627 12736 24659
rect 12768 24627 12808 24659
rect 12840 24627 12880 24659
rect 12912 24627 12952 24659
rect 12984 24627 13024 24659
rect 13056 24627 13096 24659
rect 13128 24627 13168 24659
rect 13200 24627 13240 24659
rect 13272 24627 13312 24659
rect 13344 24627 13384 24659
rect 13416 24627 13456 24659
rect 13488 24627 13528 24659
rect 13560 24627 13600 24659
rect 13632 24627 13672 24659
rect 13704 24627 13744 24659
rect 13776 24627 13816 24659
rect 13848 24627 13888 24659
rect 13920 24627 13960 24659
rect 13992 24627 14032 24659
rect 14064 24627 14104 24659
rect 14136 24627 14176 24659
rect 14208 24627 14248 24659
rect 14280 24627 14320 24659
rect 14352 24627 14392 24659
rect 14424 24627 14464 24659
rect 14496 24627 14536 24659
rect 14568 24627 14608 24659
rect 14640 24627 14680 24659
rect 14712 24627 14752 24659
rect 14784 24627 14824 24659
rect 14856 24627 14896 24659
rect 14928 24627 14968 24659
rect 15000 24627 15040 24659
rect 15072 24627 15112 24659
rect 15144 24627 15184 24659
rect 15216 24627 15256 24659
rect 15288 24627 15328 24659
rect 15360 24627 15400 24659
rect 15432 24627 15472 24659
rect 15504 24627 15544 24659
rect 15576 24627 15616 24659
rect 15648 24627 15688 24659
rect 15720 24627 15760 24659
rect 15792 24627 15832 24659
rect 15864 24627 15904 24659
rect 15936 24627 16000 24659
rect 0 24587 16000 24627
rect 0 24555 64 24587
rect 96 24555 136 24587
rect 168 24555 208 24587
rect 240 24555 280 24587
rect 312 24555 352 24587
rect 384 24555 424 24587
rect 456 24555 496 24587
rect 528 24555 568 24587
rect 600 24555 640 24587
rect 672 24555 712 24587
rect 744 24555 784 24587
rect 816 24555 856 24587
rect 888 24555 928 24587
rect 960 24555 1000 24587
rect 1032 24555 1072 24587
rect 1104 24555 1144 24587
rect 1176 24555 1216 24587
rect 1248 24555 1288 24587
rect 1320 24555 1360 24587
rect 1392 24555 1432 24587
rect 1464 24555 1504 24587
rect 1536 24555 1576 24587
rect 1608 24555 1648 24587
rect 1680 24555 1720 24587
rect 1752 24555 1792 24587
rect 1824 24555 1864 24587
rect 1896 24555 1936 24587
rect 1968 24555 2008 24587
rect 2040 24555 2080 24587
rect 2112 24555 2152 24587
rect 2184 24555 2224 24587
rect 2256 24555 2296 24587
rect 2328 24555 2368 24587
rect 2400 24555 2440 24587
rect 2472 24555 2512 24587
rect 2544 24555 2584 24587
rect 2616 24555 2656 24587
rect 2688 24555 2728 24587
rect 2760 24555 2800 24587
rect 2832 24555 2872 24587
rect 2904 24555 2944 24587
rect 2976 24555 3016 24587
rect 3048 24555 3088 24587
rect 3120 24555 3160 24587
rect 3192 24555 3232 24587
rect 3264 24555 3304 24587
rect 3336 24555 3376 24587
rect 3408 24555 3448 24587
rect 3480 24555 3520 24587
rect 3552 24555 3592 24587
rect 3624 24555 3664 24587
rect 3696 24555 3736 24587
rect 3768 24555 3808 24587
rect 3840 24555 3880 24587
rect 3912 24555 3952 24587
rect 3984 24555 4024 24587
rect 4056 24555 4096 24587
rect 4128 24555 4168 24587
rect 4200 24555 4240 24587
rect 4272 24555 4312 24587
rect 4344 24555 4384 24587
rect 4416 24555 4456 24587
rect 4488 24555 4528 24587
rect 4560 24555 4600 24587
rect 4632 24555 4672 24587
rect 4704 24555 4744 24587
rect 4776 24555 4816 24587
rect 4848 24555 4888 24587
rect 4920 24555 4960 24587
rect 4992 24555 5032 24587
rect 5064 24555 5104 24587
rect 5136 24555 5176 24587
rect 5208 24555 5248 24587
rect 5280 24555 5320 24587
rect 5352 24555 5392 24587
rect 5424 24555 5464 24587
rect 5496 24555 5536 24587
rect 5568 24555 5608 24587
rect 5640 24555 5680 24587
rect 5712 24555 5752 24587
rect 5784 24555 5824 24587
rect 5856 24555 5896 24587
rect 5928 24555 5968 24587
rect 6000 24555 6040 24587
rect 6072 24555 6112 24587
rect 6144 24555 6184 24587
rect 6216 24555 6256 24587
rect 6288 24555 6328 24587
rect 6360 24555 6400 24587
rect 6432 24555 6472 24587
rect 6504 24555 6544 24587
rect 6576 24555 6616 24587
rect 6648 24555 6688 24587
rect 6720 24555 6760 24587
rect 6792 24555 6832 24587
rect 6864 24555 6904 24587
rect 6936 24555 6976 24587
rect 7008 24555 7048 24587
rect 7080 24555 7120 24587
rect 7152 24555 7192 24587
rect 7224 24555 7264 24587
rect 7296 24555 7336 24587
rect 7368 24555 7408 24587
rect 7440 24555 7480 24587
rect 7512 24555 7552 24587
rect 7584 24555 7624 24587
rect 7656 24555 7696 24587
rect 7728 24555 7768 24587
rect 7800 24555 7840 24587
rect 7872 24555 7912 24587
rect 7944 24555 7984 24587
rect 8016 24555 8056 24587
rect 8088 24555 8128 24587
rect 8160 24555 8200 24587
rect 8232 24555 8272 24587
rect 8304 24555 8344 24587
rect 8376 24555 8416 24587
rect 8448 24555 8488 24587
rect 8520 24555 8560 24587
rect 8592 24555 8632 24587
rect 8664 24555 8704 24587
rect 8736 24555 8776 24587
rect 8808 24555 8848 24587
rect 8880 24555 8920 24587
rect 8952 24555 8992 24587
rect 9024 24555 9064 24587
rect 9096 24555 9136 24587
rect 9168 24555 9208 24587
rect 9240 24555 9280 24587
rect 9312 24555 9352 24587
rect 9384 24555 9424 24587
rect 9456 24555 9496 24587
rect 9528 24555 9568 24587
rect 9600 24555 9640 24587
rect 9672 24555 9712 24587
rect 9744 24555 9784 24587
rect 9816 24555 9856 24587
rect 9888 24555 9928 24587
rect 9960 24555 10000 24587
rect 10032 24555 10072 24587
rect 10104 24555 10144 24587
rect 10176 24555 10216 24587
rect 10248 24555 10288 24587
rect 10320 24555 10360 24587
rect 10392 24555 10432 24587
rect 10464 24555 10504 24587
rect 10536 24555 10576 24587
rect 10608 24555 10648 24587
rect 10680 24555 10720 24587
rect 10752 24555 10792 24587
rect 10824 24555 10864 24587
rect 10896 24555 10936 24587
rect 10968 24555 11008 24587
rect 11040 24555 11080 24587
rect 11112 24555 11152 24587
rect 11184 24555 11224 24587
rect 11256 24555 11296 24587
rect 11328 24555 11368 24587
rect 11400 24555 11440 24587
rect 11472 24555 11512 24587
rect 11544 24555 11584 24587
rect 11616 24555 11656 24587
rect 11688 24555 11728 24587
rect 11760 24555 11800 24587
rect 11832 24555 11872 24587
rect 11904 24555 11944 24587
rect 11976 24555 12016 24587
rect 12048 24555 12088 24587
rect 12120 24555 12160 24587
rect 12192 24555 12232 24587
rect 12264 24555 12304 24587
rect 12336 24555 12376 24587
rect 12408 24555 12448 24587
rect 12480 24555 12520 24587
rect 12552 24555 12592 24587
rect 12624 24555 12664 24587
rect 12696 24555 12736 24587
rect 12768 24555 12808 24587
rect 12840 24555 12880 24587
rect 12912 24555 12952 24587
rect 12984 24555 13024 24587
rect 13056 24555 13096 24587
rect 13128 24555 13168 24587
rect 13200 24555 13240 24587
rect 13272 24555 13312 24587
rect 13344 24555 13384 24587
rect 13416 24555 13456 24587
rect 13488 24555 13528 24587
rect 13560 24555 13600 24587
rect 13632 24555 13672 24587
rect 13704 24555 13744 24587
rect 13776 24555 13816 24587
rect 13848 24555 13888 24587
rect 13920 24555 13960 24587
rect 13992 24555 14032 24587
rect 14064 24555 14104 24587
rect 14136 24555 14176 24587
rect 14208 24555 14248 24587
rect 14280 24555 14320 24587
rect 14352 24555 14392 24587
rect 14424 24555 14464 24587
rect 14496 24555 14536 24587
rect 14568 24555 14608 24587
rect 14640 24555 14680 24587
rect 14712 24555 14752 24587
rect 14784 24555 14824 24587
rect 14856 24555 14896 24587
rect 14928 24555 14968 24587
rect 15000 24555 15040 24587
rect 15072 24555 15112 24587
rect 15144 24555 15184 24587
rect 15216 24555 15256 24587
rect 15288 24555 15328 24587
rect 15360 24555 15400 24587
rect 15432 24555 15472 24587
rect 15504 24555 15544 24587
rect 15576 24555 15616 24587
rect 15648 24555 15688 24587
rect 15720 24555 15760 24587
rect 15792 24555 15832 24587
rect 15864 24555 15904 24587
rect 15936 24555 16000 24587
rect 0 24515 16000 24555
rect 0 24483 64 24515
rect 96 24483 136 24515
rect 168 24483 208 24515
rect 240 24483 280 24515
rect 312 24483 352 24515
rect 384 24483 424 24515
rect 456 24483 496 24515
rect 528 24483 568 24515
rect 600 24483 640 24515
rect 672 24483 712 24515
rect 744 24483 784 24515
rect 816 24483 856 24515
rect 888 24483 928 24515
rect 960 24483 1000 24515
rect 1032 24483 1072 24515
rect 1104 24483 1144 24515
rect 1176 24483 1216 24515
rect 1248 24483 1288 24515
rect 1320 24483 1360 24515
rect 1392 24483 1432 24515
rect 1464 24483 1504 24515
rect 1536 24483 1576 24515
rect 1608 24483 1648 24515
rect 1680 24483 1720 24515
rect 1752 24483 1792 24515
rect 1824 24483 1864 24515
rect 1896 24483 1936 24515
rect 1968 24483 2008 24515
rect 2040 24483 2080 24515
rect 2112 24483 2152 24515
rect 2184 24483 2224 24515
rect 2256 24483 2296 24515
rect 2328 24483 2368 24515
rect 2400 24483 2440 24515
rect 2472 24483 2512 24515
rect 2544 24483 2584 24515
rect 2616 24483 2656 24515
rect 2688 24483 2728 24515
rect 2760 24483 2800 24515
rect 2832 24483 2872 24515
rect 2904 24483 2944 24515
rect 2976 24483 3016 24515
rect 3048 24483 3088 24515
rect 3120 24483 3160 24515
rect 3192 24483 3232 24515
rect 3264 24483 3304 24515
rect 3336 24483 3376 24515
rect 3408 24483 3448 24515
rect 3480 24483 3520 24515
rect 3552 24483 3592 24515
rect 3624 24483 3664 24515
rect 3696 24483 3736 24515
rect 3768 24483 3808 24515
rect 3840 24483 3880 24515
rect 3912 24483 3952 24515
rect 3984 24483 4024 24515
rect 4056 24483 4096 24515
rect 4128 24483 4168 24515
rect 4200 24483 4240 24515
rect 4272 24483 4312 24515
rect 4344 24483 4384 24515
rect 4416 24483 4456 24515
rect 4488 24483 4528 24515
rect 4560 24483 4600 24515
rect 4632 24483 4672 24515
rect 4704 24483 4744 24515
rect 4776 24483 4816 24515
rect 4848 24483 4888 24515
rect 4920 24483 4960 24515
rect 4992 24483 5032 24515
rect 5064 24483 5104 24515
rect 5136 24483 5176 24515
rect 5208 24483 5248 24515
rect 5280 24483 5320 24515
rect 5352 24483 5392 24515
rect 5424 24483 5464 24515
rect 5496 24483 5536 24515
rect 5568 24483 5608 24515
rect 5640 24483 5680 24515
rect 5712 24483 5752 24515
rect 5784 24483 5824 24515
rect 5856 24483 5896 24515
rect 5928 24483 5968 24515
rect 6000 24483 6040 24515
rect 6072 24483 6112 24515
rect 6144 24483 6184 24515
rect 6216 24483 6256 24515
rect 6288 24483 6328 24515
rect 6360 24483 6400 24515
rect 6432 24483 6472 24515
rect 6504 24483 6544 24515
rect 6576 24483 6616 24515
rect 6648 24483 6688 24515
rect 6720 24483 6760 24515
rect 6792 24483 6832 24515
rect 6864 24483 6904 24515
rect 6936 24483 6976 24515
rect 7008 24483 7048 24515
rect 7080 24483 7120 24515
rect 7152 24483 7192 24515
rect 7224 24483 7264 24515
rect 7296 24483 7336 24515
rect 7368 24483 7408 24515
rect 7440 24483 7480 24515
rect 7512 24483 7552 24515
rect 7584 24483 7624 24515
rect 7656 24483 7696 24515
rect 7728 24483 7768 24515
rect 7800 24483 7840 24515
rect 7872 24483 7912 24515
rect 7944 24483 7984 24515
rect 8016 24483 8056 24515
rect 8088 24483 8128 24515
rect 8160 24483 8200 24515
rect 8232 24483 8272 24515
rect 8304 24483 8344 24515
rect 8376 24483 8416 24515
rect 8448 24483 8488 24515
rect 8520 24483 8560 24515
rect 8592 24483 8632 24515
rect 8664 24483 8704 24515
rect 8736 24483 8776 24515
rect 8808 24483 8848 24515
rect 8880 24483 8920 24515
rect 8952 24483 8992 24515
rect 9024 24483 9064 24515
rect 9096 24483 9136 24515
rect 9168 24483 9208 24515
rect 9240 24483 9280 24515
rect 9312 24483 9352 24515
rect 9384 24483 9424 24515
rect 9456 24483 9496 24515
rect 9528 24483 9568 24515
rect 9600 24483 9640 24515
rect 9672 24483 9712 24515
rect 9744 24483 9784 24515
rect 9816 24483 9856 24515
rect 9888 24483 9928 24515
rect 9960 24483 10000 24515
rect 10032 24483 10072 24515
rect 10104 24483 10144 24515
rect 10176 24483 10216 24515
rect 10248 24483 10288 24515
rect 10320 24483 10360 24515
rect 10392 24483 10432 24515
rect 10464 24483 10504 24515
rect 10536 24483 10576 24515
rect 10608 24483 10648 24515
rect 10680 24483 10720 24515
rect 10752 24483 10792 24515
rect 10824 24483 10864 24515
rect 10896 24483 10936 24515
rect 10968 24483 11008 24515
rect 11040 24483 11080 24515
rect 11112 24483 11152 24515
rect 11184 24483 11224 24515
rect 11256 24483 11296 24515
rect 11328 24483 11368 24515
rect 11400 24483 11440 24515
rect 11472 24483 11512 24515
rect 11544 24483 11584 24515
rect 11616 24483 11656 24515
rect 11688 24483 11728 24515
rect 11760 24483 11800 24515
rect 11832 24483 11872 24515
rect 11904 24483 11944 24515
rect 11976 24483 12016 24515
rect 12048 24483 12088 24515
rect 12120 24483 12160 24515
rect 12192 24483 12232 24515
rect 12264 24483 12304 24515
rect 12336 24483 12376 24515
rect 12408 24483 12448 24515
rect 12480 24483 12520 24515
rect 12552 24483 12592 24515
rect 12624 24483 12664 24515
rect 12696 24483 12736 24515
rect 12768 24483 12808 24515
rect 12840 24483 12880 24515
rect 12912 24483 12952 24515
rect 12984 24483 13024 24515
rect 13056 24483 13096 24515
rect 13128 24483 13168 24515
rect 13200 24483 13240 24515
rect 13272 24483 13312 24515
rect 13344 24483 13384 24515
rect 13416 24483 13456 24515
rect 13488 24483 13528 24515
rect 13560 24483 13600 24515
rect 13632 24483 13672 24515
rect 13704 24483 13744 24515
rect 13776 24483 13816 24515
rect 13848 24483 13888 24515
rect 13920 24483 13960 24515
rect 13992 24483 14032 24515
rect 14064 24483 14104 24515
rect 14136 24483 14176 24515
rect 14208 24483 14248 24515
rect 14280 24483 14320 24515
rect 14352 24483 14392 24515
rect 14424 24483 14464 24515
rect 14496 24483 14536 24515
rect 14568 24483 14608 24515
rect 14640 24483 14680 24515
rect 14712 24483 14752 24515
rect 14784 24483 14824 24515
rect 14856 24483 14896 24515
rect 14928 24483 14968 24515
rect 15000 24483 15040 24515
rect 15072 24483 15112 24515
rect 15144 24483 15184 24515
rect 15216 24483 15256 24515
rect 15288 24483 15328 24515
rect 15360 24483 15400 24515
rect 15432 24483 15472 24515
rect 15504 24483 15544 24515
rect 15576 24483 15616 24515
rect 15648 24483 15688 24515
rect 15720 24483 15760 24515
rect 15792 24483 15832 24515
rect 15864 24483 15904 24515
rect 15936 24483 16000 24515
rect 0 24443 16000 24483
rect 0 24411 64 24443
rect 96 24411 136 24443
rect 168 24411 208 24443
rect 240 24411 280 24443
rect 312 24411 352 24443
rect 384 24411 424 24443
rect 456 24411 496 24443
rect 528 24411 568 24443
rect 600 24411 640 24443
rect 672 24411 712 24443
rect 744 24411 784 24443
rect 816 24411 856 24443
rect 888 24411 928 24443
rect 960 24411 1000 24443
rect 1032 24411 1072 24443
rect 1104 24411 1144 24443
rect 1176 24411 1216 24443
rect 1248 24411 1288 24443
rect 1320 24411 1360 24443
rect 1392 24411 1432 24443
rect 1464 24411 1504 24443
rect 1536 24411 1576 24443
rect 1608 24411 1648 24443
rect 1680 24411 1720 24443
rect 1752 24411 1792 24443
rect 1824 24411 1864 24443
rect 1896 24411 1936 24443
rect 1968 24411 2008 24443
rect 2040 24411 2080 24443
rect 2112 24411 2152 24443
rect 2184 24411 2224 24443
rect 2256 24411 2296 24443
rect 2328 24411 2368 24443
rect 2400 24411 2440 24443
rect 2472 24411 2512 24443
rect 2544 24411 2584 24443
rect 2616 24411 2656 24443
rect 2688 24411 2728 24443
rect 2760 24411 2800 24443
rect 2832 24411 2872 24443
rect 2904 24411 2944 24443
rect 2976 24411 3016 24443
rect 3048 24411 3088 24443
rect 3120 24411 3160 24443
rect 3192 24411 3232 24443
rect 3264 24411 3304 24443
rect 3336 24411 3376 24443
rect 3408 24411 3448 24443
rect 3480 24411 3520 24443
rect 3552 24411 3592 24443
rect 3624 24411 3664 24443
rect 3696 24411 3736 24443
rect 3768 24411 3808 24443
rect 3840 24411 3880 24443
rect 3912 24411 3952 24443
rect 3984 24411 4024 24443
rect 4056 24411 4096 24443
rect 4128 24411 4168 24443
rect 4200 24411 4240 24443
rect 4272 24411 4312 24443
rect 4344 24411 4384 24443
rect 4416 24411 4456 24443
rect 4488 24411 4528 24443
rect 4560 24411 4600 24443
rect 4632 24411 4672 24443
rect 4704 24411 4744 24443
rect 4776 24411 4816 24443
rect 4848 24411 4888 24443
rect 4920 24411 4960 24443
rect 4992 24411 5032 24443
rect 5064 24411 5104 24443
rect 5136 24411 5176 24443
rect 5208 24411 5248 24443
rect 5280 24411 5320 24443
rect 5352 24411 5392 24443
rect 5424 24411 5464 24443
rect 5496 24411 5536 24443
rect 5568 24411 5608 24443
rect 5640 24411 5680 24443
rect 5712 24411 5752 24443
rect 5784 24411 5824 24443
rect 5856 24411 5896 24443
rect 5928 24411 5968 24443
rect 6000 24411 6040 24443
rect 6072 24411 6112 24443
rect 6144 24411 6184 24443
rect 6216 24411 6256 24443
rect 6288 24411 6328 24443
rect 6360 24411 6400 24443
rect 6432 24411 6472 24443
rect 6504 24411 6544 24443
rect 6576 24411 6616 24443
rect 6648 24411 6688 24443
rect 6720 24411 6760 24443
rect 6792 24411 6832 24443
rect 6864 24411 6904 24443
rect 6936 24411 6976 24443
rect 7008 24411 7048 24443
rect 7080 24411 7120 24443
rect 7152 24411 7192 24443
rect 7224 24411 7264 24443
rect 7296 24411 7336 24443
rect 7368 24411 7408 24443
rect 7440 24411 7480 24443
rect 7512 24411 7552 24443
rect 7584 24411 7624 24443
rect 7656 24411 7696 24443
rect 7728 24411 7768 24443
rect 7800 24411 7840 24443
rect 7872 24411 7912 24443
rect 7944 24411 7984 24443
rect 8016 24411 8056 24443
rect 8088 24411 8128 24443
rect 8160 24411 8200 24443
rect 8232 24411 8272 24443
rect 8304 24411 8344 24443
rect 8376 24411 8416 24443
rect 8448 24411 8488 24443
rect 8520 24411 8560 24443
rect 8592 24411 8632 24443
rect 8664 24411 8704 24443
rect 8736 24411 8776 24443
rect 8808 24411 8848 24443
rect 8880 24411 8920 24443
rect 8952 24411 8992 24443
rect 9024 24411 9064 24443
rect 9096 24411 9136 24443
rect 9168 24411 9208 24443
rect 9240 24411 9280 24443
rect 9312 24411 9352 24443
rect 9384 24411 9424 24443
rect 9456 24411 9496 24443
rect 9528 24411 9568 24443
rect 9600 24411 9640 24443
rect 9672 24411 9712 24443
rect 9744 24411 9784 24443
rect 9816 24411 9856 24443
rect 9888 24411 9928 24443
rect 9960 24411 10000 24443
rect 10032 24411 10072 24443
rect 10104 24411 10144 24443
rect 10176 24411 10216 24443
rect 10248 24411 10288 24443
rect 10320 24411 10360 24443
rect 10392 24411 10432 24443
rect 10464 24411 10504 24443
rect 10536 24411 10576 24443
rect 10608 24411 10648 24443
rect 10680 24411 10720 24443
rect 10752 24411 10792 24443
rect 10824 24411 10864 24443
rect 10896 24411 10936 24443
rect 10968 24411 11008 24443
rect 11040 24411 11080 24443
rect 11112 24411 11152 24443
rect 11184 24411 11224 24443
rect 11256 24411 11296 24443
rect 11328 24411 11368 24443
rect 11400 24411 11440 24443
rect 11472 24411 11512 24443
rect 11544 24411 11584 24443
rect 11616 24411 11656 24443
rect 11688 24411 11728 24443
rect 11760 24411 11800 24443
rect 11832 24411 11872 24443
rect 11904 24411 11944 24443
rect 11976 24411 12016 24443
rect 12048 24411 12088 24443
rect 12120 24411 12160 24443
rect 12192 24411 12232 24443
rect 12264 24411 12304 24443
rect 12336 24411 12376 24443
rect 12408 24411 12448 24443
rect 12480 24411 12520 24443
rect 12552 24411 12592 24443
rect 12624 24411 12664 24443
rect 12696 24411 12736 24443
rect 12768 24411 12808 24443
rect 12840 24411 12880 24443
rect 12912 24411 12952 24443
rect 12984 24411 13024 24443
rect 13056 24411 13096 24443
rect 13128 24411 13168 24443
rect 13200 24411 13240 24443
rect 13272 24411 13312 24443
rect 13344 24411 13384 24443
rect 13416 24411 13456 24443
rect 13488 24411 13528 24443
rect 13560 24411 13600 24443
rect 13632 24411 13672 24443
rect 13704 24411 13744 24443
rect 13776 24411 13816 24443
rect 13848 24411 13888 24443
rect 13920 24411 13960 24443
rect 13992 24411 14032 24443
rect 14064 24411 14104 24443
rect 14136 24411 14176 24443
rect 14208 24411 14248 24443
rect 14280 24411 14320 24443
rect 14352 24411 14392 24443
rect 14424 24411 14464 24443
rect 14496 24411 14536 24443
rect 14568 24411 14608 24443
rect 14640 24411 14680 24443
rect 14712 24411 14752 24443
rect 14784 24411 14824 24443
rect 14856 24411 14896 24443
rect 14928 24411 14968 24443
rect 15000 24411 15040 24443
rect 15072 24411 15112 24443
rect 15144 24411 15184 24443
rect 15216 24411 15256 24443
rect 15288 24411 15328 24443
rect 15360 24411 15400 24443
rect 15432 24411 15472 24443
rect 15504 24411 15544 24443
rect 15576 24411 15616 24443
rect 15648 24411 15688 24443
rect 15720 24411 15760 24443
rect 15792 24411 15832 24443
rect 15864 24411 15904 24443
rect 15936 24411 16000 24443
rect 0 24371 16000 24411
rect 0 24339 64 24371
rect 96 24339 136 24371
rect 168 24339 208 24371
rect 240 24339 280 24371
rect 312 24339 352 24371
rect 384 24339 424 24371
rect 456 24339 496 24371
rect 528 24339 568 24371
rect 600 24339 640 24371
rect 672 24339 712 24371
rect 744 24339 784 24371
rect 816 24339 856 24371
rect 888 24339 928 24371
rect 960 24339 1000 24371
rect 1032 24339 1072 24371
rect 1104 24339 1144 24371
rect 1176 24339 1216 24371
rect 1248 24339 1288 24371
rect 1320 24339 1360 24371
rect 1392 24339 1432 24371
rect 1464 24339 1504 24371
rect 1536 24339 1576 24371
rect 1608 24339 1648 24371
rect 1680 24339 1720 24371
rect 1752 24339 1792 24371
rect 1824 24339 1864 24371
rect 1896 24339 1936 24371
rect 1968 24339 2008 24371
rect 2040 24339 2080 24371
rect 2112 24339 2152 24371
rect 2184 24339 2224 24371
rect 2256 24339 2296 24371
rect 2328 24339 2368 24371
rect 2400 24339 2440 24371
rect 2472 24339 2512 24371
rect 2544 24339 2584 24371
rect 2616 24339 2656 24371
rect 2688 24339 2728 24371
rect 2760 24339 2800 24371
rect 2832 24339 2872 24371
rect 2904 24339 2944 24371
rect 2976 24339 3016 24371
rect 3048 24339 3088 24371
rect 3120 24339 3160 24371
rect 3192 24339 3232 24371
rect 3264 24339 3304 24371
rect 3336 24339 3376 24371
rect 3408 24339 3448 24371
rect 3480 24339 3520 24371
rect 3552 24339 3592 24371
rect 3624 24339 3664 24371
rect 3696 24339 3736 24371
rect 3768 24339 3808 24371
rect 3840 24339 3880 24371
rect 3912 24339 3952 24371
rect 3984 24339 4024 24371
rect 4056 24339 4096 24371
rect 4128 24339 4168 24371
rect 4200 24339 4240 24371
rect 4272 24339 4312 24371
rect 4344 24339 4384 24371
rect 4416 24339 4456 24371
rect 4488 24339 4528 24371
rect 4560 24339 4600 24371
rect 4632 24339 4672 24371
rect 4704 24339 4744 24371
rect 4776 24339 4816 24371
rect 4848 24339 4888 24371
rect 4920 24339 4960 24371
rect 4992 24339 5032 24371
rect 5064 24339 5104 24371
rect 5136 24339 5176 24371
rect 5208 24339 5248 24371
rect 5280 24339 5320 24371
rect 5352 24339 5392 24371
rect 5424 24339 5464 24371
rect 5496 24339 5536 24371
rect 5568 24339 5608 24371
rect 5640 24339 5680 24371
rect 5712 24339 5752 24371
rect 5784 24339 5824 24371
rect 5856 24339 5896 24371
rect 5928 24339 5968 24371
rect 6000 24339 6040 24371
rect 6072 24339 6112 24371
rect 6144 24339 6184 24371
rect 6216 24339 6256 24371
rect 6288 24339 6328 24371
rect 6360 24339 6400 24371
rect 6432 24339 6472 24371
rect 6504 24339 6544 24371
rect 6576 24339 6616 24371
rect 6648 24339 6688 24371
rect 6720 24339 6760 24371
rect 6792 24339 6832 24371
rect 6864 24339 6904 24371
rect 6936 24339 6976 24371
rect 7008 24339 7048 24371
rect 7080 24339 7120 24371
rect 7152 24339 7192 24371
rect 7224 24339 7264 24371
rect 7296 24339 7336 24371
rect 7368 24339 7408 24371
rect 7440 24339 7480 24371
rect 7512 24339 7552 24371
rect 7584 24339 7624 24371
rect 7656 24339 7696 24371
rect 7728 24339 7768 24371
rect 7800 24339 7840 24371
rect 7872 24339 7912 24371
rect 7944 24339 7984 24371
rect 8016 24339 8056 24371
rect 8088 24339 8128 24371
rect 8160 24339 8200 24371
rect 8232 24339 8272 24371
rect 8304 24339 8344 24371
rect 8376 24339 8416 24371
rect 8448 24339 8488 24371
rect 8520 24339 8560 24371
rect 8592 24339 8632 24371
rect 8664 24339 8704 24371
rect 8736 24339 8776 24371
rect 8808 24339 8848 24371
rect 8880 24339 8920 24371
rect 8952 24339 8992 24371
rect 9024 24339 9064 24371
rect 9096 24339 9136 24371
rect 9168 24339 9208 24371
rect 9240 24339 9280 24371
rect 9312 24339 9352 24371
rect 9384 24339 9424 24371
rect 9456 24339 9496 24371
rect 9528 24339 9568 24371
rect 9600 24339 9640 24371
rect 9672 24339 9712 24371
rect 9744 24339 9784 24371
rect 9816 24339 9856 24371
rect 9888 24339 9928 24371
rect 9960 24339 10000 24371
rect 10032 24339 10072 24371
rect 10104 24339 10144 24371
rect 10176 24339 10216 24371
rect 10248 24339 10288 24371
rect 10320 24339 10360 24371
rect 10392 24339 10432 24371
rect 10464 24339 10504 24371
rect 10536 24339 10576 24371
rect 10608 24339 10648 24371
rect 10680 24339 10720 24371
rect 10752 24339 10792 24371
rect 10824 24339 10864 24371
rect 10896 24339 10936 24371
rect 10968 24339 11008 24371
rect 11040 24339 11080 24371
rect 11112 24339 11152 24371
rect 11184 24339 11224 24371
rect 11256 24339 11296 24371
rect 11328 24339 11368 24371
rect 11400 24339 11440 24371
rect 11472 24339 11512 24371
rect 11544 24339 11584 24371
rect 11616 24339 11656 24371
rect 11688 24339 11728 24371
rect 11760 24339 11800 24371
rect 11832 24339 11872 24371
rect 11904 24339 11944 24371
rect 11976 24339 12016 24371
rect 12048 24339 12088 24371
rect 12120 24339 12160 24371
rect 12192 24339 12232 24371
rect 12264 24339 12304 24371
rect 12336 24339 12376 24371
rect 12408 24339 12448 24371
rect 12480 24339 12520 24371
rect 12552 24339 12592 24371
rect 12624 24339 12664 24371
rect 12696 24339 12736 24371
rect 12768 24339 12808 24371
rect 12840 24339 12880 24371
rect 12912 24339 12952 24371
rect 12984 24339 13024 24371
rect 13056 24339 13096 24371
rect 13128 24339 13168 24371
rect 13200 24339 13240 24371
rect 13272 24339 13312 24371
rect 13344 24339 13384 24371
rect 13416 24339 13456 24371
rect 13488 24339 13528 24371
rect 13560 24339 13600 24371
rect 13632 24339 13672 24371
rect 13704 24339 13744 24371
rect 13776 24339 13816 24371
rect 13848 24339 13888 24371
rect 13920 24339 13960 24371
rect 13992 24339 14032 24371
rect 14064 24339 14104 24371
rect 14136 24339 14176 24371
rect 14208 24339 14248 24371
rect 14280 24339 14320 24371
rect 14352 24339 14392 24371
rect 14424 24339 14464 24371
rect 14496 24339 14536 24371
rect 14568 24339 14608 24371
rect 14640 24339 14680 24371
rect 14712 24339 14752 24371
rect 14784 24339 14824 24371
rect 14856 24339 14896 24371
rect 14928 24339 14968 24371
rect 15000 24339 15040 24371
rect 15072 24339 15112 24371
rect 15144 24339 15184 24371
rect 15216 24339 15256 24371
rect 15288 24339 15328 24371
rect 15360 24339 15400 24371
rect 15432 24339 15472 24371
rect 15504 24339 15544 24371
rect 15576 24339 15616 24371
rect 15648 24339 15688 24371
rect 15720 24339 15760 24371
rect 15792 24339 15832 24371
rect 15864 24339 15904 24371
rect 15936 24339 16000 24371
rect 0 24299 16000 24339
rect 0 24267 64 24299
rect 96 24267 136 24299
rect 168 24267 208 24299
rect 240 24267 280 24299
rect 312 24267 352 24299
rect 384 24267 424 24299
rect 456 24267 496 24299
rect 528 24267 568 24299
rect 600 24267 640 24299
rect 672 24267 712 24299
rect 744 24267 784 24299
rect 816 24267 856 24299
rect 888 24267 928 24299
rect 960 24267 1000 24299
rect 1032 24267 1072 24299
rect 1104 24267 1144 24299
rect 1176 24267 1216 24299
rect 1248 24267 1288 24299
rect 1320 24267 1360 24299
rect 1392 24267 1432 24299
rect 1464 24267 1504 24299
rect 1536 24267 1576 24299
rect 1608 24267 1648 24299
rect 1680 24267 1720 24299
rect 1752 24267 1792 24299
rect 1824 24267 1864 24299
rect 1896 24267 1936 24299
rect 1968 24267 2008 24299
rect 2040 24267 2080 24299
rect 2112 24267 2152 24299
rect 2184 24267 2224 24299
rect 2256 24267 2296 24299
rect 2328 24267 2368 24299
rect 2400 24267 2440 24299
rect 2472 24267 2512 24299
rect 2544 24267 2584 24299
rect 2616 24267 2656 24299
rect 2688 24267 2728 24299
rect 2760 24267 2800 24299
rect 2832 24267 2872 24299
rect 2904 24267 2944 24299
rect 2976 24267 3016 24299
rect 3048 24267 3088 24299
rect 3120 24267 3160 24299
rect 3192 24267 3232 24299
rect 3264 24267 3304 24299
rect 3336 24267 3376 24299
rect 3408 24267 3448 24299
rect 3480 24267 3520 24299
rect 3552 24267 3592 24299
rect 3624 24267 3664 24299
rect 3696 24267 3736 24299
rect 3768 24267 3808 24299
rect 3840 24267 3880 24299
rect 3912 24267 3952 24299
rect 3984 24267 4024 24299
rect 4056 24267 4096 24299
rect 4128 24267 4168 24299
rect 4200 24267 4240 24299
rect 4272 24267 4312 24299
rect 4344 24267 4384 24299
rect 4416 24267 4456 24299
rect 4488 24267 4528 24299
rect 4560 24267 4600 24299
rect 4632 24267 4672 24299
rect 4704 24267 4744 24299
rect 4776 24267 4816 24299
rect 4848 24267 4888 24299
rect 4920 24267 4960 24299
rect 4992 24267 5032 24299
rect 5064 24267 5104 24299
rect 5136 24267 5176 24299
rect 5208 24267 5248 24299
rect 5280 24267 5320 24299
rect 5352 24267 5392 24299
rect 5424 24267 5464 24299
rect 5496 24267 5536 24299
rect 5568 24267 5608 24299
rect 5640 24267 5680 24299
rect 5712 24267 5752 24299
rect 5784 24267 5824 24299
rect 5856 24267 5896 24299
rect 5928 24267 5968 24299
rect 6000 24267 6040 24299
rect 6072 24267 6112 24299
rect 6144 24267 6184 24299
rect 6216 24267 6256 24299
rect 6288 24267 6328 24299
rect 6360 24267 6400 24299
rect 6432 24267 6472 24299
rect 6504 24267 6544 24299
rect 6576 24267 6616 24299
rect 6648 24267 6688 24299
rect 6720 24267 6760 24299
rect 6792 24267 6832 24299
rect 6864 24267 6904 24299
rect 6936 24267 6976 24299
rect 7008 24267 7048 24299
rect 7080 24267 7120 24299
rect 7152 24267 7192 24299
rect 7224 24267 7264 24299
rect 7296 24267 7336 24299
rect 7368 24267 7408 24299
rect 7440 24267 7480 24299
rect 7512 24267 7552 24299
rect 7584 24267 7624 24299
rect 7656 24267 7696 24299
rect 7728 24267 7768 24299
rect 7800 24267 7840 24299
rect 7872 24267 7912 24299
rect 7944 24267 7984 24299
rect 8016 24267 8056 24299
rect 8088 24267 8128 24299
rect 8160 24267 8200 24299
rect 8232 24267 8272 24299
rect 8304 24267 8344 24299
rect 8376 24267 8416 24299
rect 8448 24267 8488 24299
rect 8520 24267 8560 24299
rect 8592 24267 8632 24299
rect 8664 24267 8704 24299
rect 8736 24267 8776 24299
rect 8808 24267 8848 24299
rect 8880 24267 8920 24299
rect 8952 24267 8992 24299
rect 9024 24267 9064 24299
rect 9096 24267 9136 24299
rect 9168 24267 9208 24299
rect 9240 24267 9280 24299
rect 9312 24267 9352 24299
rect 9384 24267 9424 24299
rect 9456 24267 9496 24299
rect 9528 24267 9568 24299
rect 9600 24267 9640 24299
rect 9672 24267 9712 24299
rect 9744 24267 9784 24299
rect 9816 24267 9856 24299
rect 9888 24267 9928 24299
rect 9960 24267 10000 24299
rect 10032 24267 10072 24299
rect 10104 24267 10144 24299
rect 10176 24267 10216 24299
rect 10248 24267 10288 24299
rect 10320 24267 10360 24299
rect 10392 24267 10432 24299
rect 10464 24267 10504 24299
rect 10536 24267 10576 24299
rect 10608 24267 10648 24299
rect 10680 24267 10720 24299
rect 10752 24267 10792 24299
rect 10824 24267 10864 24299
rect 10896 24267 10936 24299
rect 10968 24267 11008 24299
rect 11040 24267 11080 24299
rect 11112 24267 11152 24299
rect 11184 24267 11224 24299
rect 11256 24267 11296 24299
rect 11328 24267 11368 24299
rect 11400 24267 11440 24299
rect 11472 24267 11512 24299
rect 11544 24267 11584 24299
rect 11616 24267 11656 24299
rect 11688 24267 11728 24299
rect 11760 24267 11800 24299
rect 11832 24267 11872 24299
rect 11904 24267 11944 24299
rect 11976 24267 12016 24299
rect 12048 24267 12088 24299
rect 12120 24267 12160 24299
rect 12192 24267 12232 24299
rect 12264 24267 12304 24299
rect 12336 24267 12376 24299
rect 12408 24267 12448 24299
rect 12480 24267 12520 24299
rect 12552 24267 12592 24299
rect 12624 24267 12664 24299
rect 12696 24267 12736 24299
rect 12768 24267 12808 24299
rect 12840 24267 12880 24299
rect 12912 24267 12952 24299
rect 12984 24267 13024 24299
rect 13056 24267 13096 24299
rect 13128 24267 13168 24299
rect 13200 24267 13240 24299
rect 13272 24267 13312 24299
rect 13344 24267 13384 24299
rect 13416 24267 13456 24299
rect 13488 24267 13528 24299
rect 13560 24267 13600 24299
rect 13632 24267 13672 24299
rect 13704 24267 13744 24299
rect 13776 24267 13816 24299
rect 13848 24267 13888 24299
rect 13920 24267 13960 24299
rect 13992 24267 14032 24299
rect 14064 24267 14104 24299
rect 14136 24267 14176 24299
rect 14208 24267 14248 24299
rect 14280 24267 14320 24299
rect 14352 24267 14392 24299
rect 14424 24267 14464 24299
rect 14496 24267 14536 24299
rect 14568 24267 14608 24299
rect 14640 24267 14680 24299
rect 14712 24267 14752 24299
rect 14784 24267 14824 24299
rect 14856 24267 14896 24299
rect 14928 24267 14968 24299
rect 15000 24267 15040 24299
rect 15072 24267 15112 24299
rect 15144 24267 15184 24299
rect 15216 24267 15256 24299
rect 15288 24267 15328 24299
rect 15360 24267 15400 24299
rect 15432 24267 15472 24299
rect 15504 24267 15544 24299
rect 15576 24267 15616 24299
rect 15648 24267 15688 24299
rect 15720 24267 15760 24299
rect 15792 24267 15832 24299
rect 15864 24267 15904 24299
rect 15936 24267 16000 24299
rect 0 24227 16000 24267
rect 0 24195 64 24227
rect 96 24195 136 24227
rect 168 24195 208 24227
rect 240 24195 280 24227
rect 312 24195 352 24227
rect 384 24195 424 24227
rect 456 24195 496 24227
rect 528 24195 568 24227
rect 600 24195 640 24227
rect 672 24195 712 24227
rect 744 24195 784 24227
rect 816 24195 856 24227
rect 888 24195 928 24227
rect 960 24195 1000 24227
rect 1032 24195 1072 24227
rect 1104 24195 1144 24227
rect 1176 24195 1216 24227
rect 1248 24195 1288 24227
rect 1320 24195 1360 24227
rect 1392 24195 1432 24227
rect 1464 24195 1504 24227
rect 1536 24195 1576 24227
rect 1608 24195 1648 24227
rect 1680 24195 1720 24227
rect 1752 24195 1792 24227
rect 1824 24195 1864 24227
rect 1896 24195 1936 24227
rect 1968 24195 2008 24227
rect 2040 24195 2080 24227
rect 2112 24195 2152 24227
rect 2184 24195 2224 24227
rect 2256 24195 2296 24227
rect 2328 24195 2368 24227
rect 2400 24195 2440 24227
rect 2472 24195 2512 24227
rect 2544 24195 2584 24227
rect 2616 24195 2656 24227
rect 2688 24195 2728 24227
rect 2760 24195 2800 24227
rect 2832 24195 2872 24227
rect 2904 24195 2944 24227
rect 2976 24195 3016 24227
rect 3048 24195 3088 24227
rect 3120 24195 3160 24227
rect 3192 24195 3232 24227
rect 3264 24195 3304 24227
rect 3336 24195 3376 24227
rect 3408 24195 3448 24227
rect 3480 24195 3520 24227
rect 3552 24195 3592 24227
rect 3624 24195 3664 24227
rect 3696 24195 3736 24227
rect 3768 24195 3808 24227
rect 3840 24195 3880 24227
rect 3912 24195 3952 24227
rect 3984 24195 4024 24227
rect 4056 24195 4096 24227
rect 4128 24195 4168 24227
rect 4200 24195 4240 24227
rect 4272 24195 4312 24227
rect 4344 24195 4384 24227
rect 4416 24195 4456 24227
rect 4488 24195 4528 24227
rect 4560 24195 4600 24227
rect 4632 24195 4672 24227
rect 4704 24195 4744 24227
rect 4776 24195 4816 24227
rect 4848 24195 4888 24227
rect 4920 24195 4960 24227
rect 4992 24195 5032 24227
rect 5064 24195 5104 24227
rect 5136 24195 5176 24227
rect 5208 24195 5248 24227
rect 5280 24195 5320 24227
rect 5352 24195 5392 24227
rect 5424 24195 5464 24227
rect 5496 24195 5536 24227
rect 5568 24195 5608 24227
rect 5640 24195 5680 24227
rect 5712 24195 5752 24227
rect 5784 24195 5824 24227
rect 5856 24195 5896 24227
rect 5928 24195 5968 24227
rect 6000 24195 6040 24227
rect 6072 24195 6112 24227
rect 6144 24195 6184 24227
rect 6216 24195 6256 24227
rect 6288 24195 6328 24227
rect 6360 24195 6400 24227
rect 6432 24195 6472 24227
rect 6504 24195 6544 24227
rect 6576 24195 6616 24227
rect 6648 24195 6688 24227
rect 6720 24195 6760 24227
rect 6792 24195 6832 24227
rect 6864 24195 6904 24227
rect 6936 24195 6976 24227
rect 7008 24195 7048 24227
rect 7080 24195 7120 24227
rect 7152 24195 7192 24227
rect 7224 24195 7264 24227
rect 7296 24195 7336 24227
rect 7368 24195 7408 24227
rect 7440 24195 7480 24227
rect 7512 24195 7552 24227
rect 7584 24195 7624 24227
rect 7656 24195 7696 24227
rect 7728 24195 7768 24227
rect 7800 24195 7840 24227
rect 7872 24195 7912 24227
rect 7944 24195 7984 24227
rect 8016 24195 8056 24227
rect 8088 24195 8128 24227
rect 8160 24195 8200 24227
rect 8232 24195 8272 24227
rect 8304 24195 8344 24227
rect 8376 24195 8416 24227
rect 8448 24195 8488 24227
rect 8520 24195 8560 24227
rect 8592 24195 8632 24227
rect 8664 24195 8704 24227
rect 8736 24195 8776 24227
rect 8808 24195 8848 24227
rect 8880 24195 8920 24227
rect 8952 24195 8992 24227
rect 9024 24195 9064 24227
rect 9096 24195 9136 24227
rect 9168 24195 9208 24227
rect 9240 24195 9280 24227
rect 9312 24195 9352 24227
rect 9384 24195 9424 24227
rect 9456 24195 9496 24227
rect 9528 24195 9568 24227
rect 9600 24195 9640 24227
rect 9672 24195 9712 24227
rect 9744 24195 9784 24227
rect 9816 24195 9856 24227
rect 9888 24195 9928 24227
rect 9960 24195 10000 24227
rect 10032 24195 10072 24227
rect 10104 24195 10144 24227
rect 10176 24195 10216 24227
rect 10248 24195 10288 24227
rect 10320 24195 10360 24227
rect 10392 24195 10432 24227
rect 10464 24195 10504 24227
rect 10536 24195 10576 24227
rect 10608 24195 10648 24227
rect 10680 24195 10720 24227
rect 10752 24195 10792 24227
rect 10824 24195 10864 24227
rect 10896 24195 10936 24227
rect 10968 24195 11008 24227
rect 11040 24195 11080 24227
rect 11112 24195 11152 24227
rect 11184 24195 11224 24227
rect 11256 24195 11296 24227
rect 11328 24195 11368 24227
rect 11400 24195 11440 24227
rect 11472 24195 11512 24227
rect 11544 24195 11584 24227
rect 11616 24195 11656 24227
rect 11688 24195 11728 24227
rect 11760 24195 11800 24227
rect 11832 24195 11872 24227
rect 11904 24195 11944 24227
rect 11976 24195 12016 24227
rect 12048 24195 12088 24227
rect 12120 24195 12160 24227
rect 12192 24195 12232 24227
rect 12264 24195 12304 24227
rect 12336 24195 12376 24227
rect 12408 24195 12448 24227
rect 12480 24195 12520 24227
rect 12552 24195 12592 24227
rect 12624 24195 12664 24227
rect 12696 24195 12736 24227
rect 12768 24195 12808 24227
rect 12840 24195 12880 24227
rect 12912 24195 12952 24227
rect 12984 24195 13024 24227
rect 13056 24195 13096 24227
rect 13128 24195 13168 24227
rect 13200 24195 13240 24227
rect 13272 24195 13312 24227
rect 13344 24195 13384 24227
rect 13416 24195 13456 24227
rect 13488 24195 13528 24227
rect 13560 24195 13600 24227
rect 13632 24195 13672 24227
rect 13704 24195 13744 24227
rect 13776 24195 13816 24227
rect 13848 24195 13888 24227
rect 13920 24195 13960 24227
rect 13992 24195 14032 24227
rect 14064 24195 14104 24227
rect 14136 24195 14176 24227
rect 14208 24195 14248 24227
rect 14280 24195 14320 24227
rect 14352 24195 14392 24227
rect 14424 24195 14464 24227
rect 14496 24195 14536 24227
rect 14568 24195 14608 24227
rect 14640 24195 14680 24227
rect 14712 24195 14752 24227
rect 14784 24195 14824 24227
rect 14856 24195 14896 24227
rect 14928 24195 14968 24227
rect 15000 24195 15040 24227
rect 15072 24195 15112 24227
rect 15144 24195 15184 24227
rect 15216 24195 15256 24227
rect 15288 24195 15328 24227
rect 15360 24195 15400 24227
rect 15432 24195 15472 24227
rect 15504 24195 15544 24227
rect 15576 24195 15616 24227
rect 15648 24195 15688 24227
rect 15720 24195 15760 24227
rect 15792 24195 15832 24227
rect 15864 24195 15904 24227
rect 15936 24195 16000 24227
rect 0 24155 16000 24195
rect 0 24123 64 24155
rect 96 24123 136 24155
rect 168 24123 208 24155
rect 240 24123 280 24155
rect 312 24123 352 24155
rect 384 24123 424 24155
rect 456 24123 496 24155
rect 528 24123 568 24155
rect 600 24123 640 24155
rect 672 24123 712 24155
rect 744 24123 784 24155
rect 816 24123 856 24155
rect 888 24123 928 24155
rect 960 24123 1000 24155
rect 1032 24123 1072 24155
rect 1104 24123 1144 24155
rect 1176 24123 1216 24155
rect 1248 24123 1288 24155
rect 1320 24123 1360 24155
rect 1392 24123 1432 24155
rect 1464 24123 1504 24155
rect 1536 24123 1576 24155
rect 1608 24123 1648 24155
rect 1680 24123 1720 24155
rect 1752 24123 1792 24155
rect 1824 24123 1864 24155
rect 1896 24123 1936 24155
rect 1968 24123 2008 24155
rect 2040 24123 2080 24155
rect 2112 24123 2152 24155
rect 2184 24123 2224 24155
rect 2256 24123 2296 24155
rect 2328 24123 2368 24155
rect 2400 24123 2440 24155
rect 2472 24123 2512 24155
rect 2544 24123 2584 24155
rect 2616 24123 2656 24155
rect 2688 24123 2728 24155
rect 2760 24123 2800 24155
rect 2832 24123 2872 24155
rect 2904 24123 2944 24155
rect 2976 24123 3016 24155
rect 3048 24123 3088 24155
rect 3120 24123 3160 24155
rect 3192 24123 3232 24155
rect 3264 24123 3304 24155
rect 3336 24123 3376 24155
rect 3408 24123 3448 24155
rect 3480 24123 3520 24155
rect 3552 24123 3592 24155
rect 3624 24123 3664 24155
rect 3696 24123 3736 24155
rect 3768 24123 3808 24155
rect 3840 24123 3880 24155
rect 3912 24123 3952 24155
rect 3984 24123 4024 24155
rect 4056 24123 4096 24155
rect 4128 24123 4168 24155
rect 4200 24123 4240 24155
rect 4272 24123 4312 24155
rect 4344 24123 4384 24155
rect 4416 24123 4456 24155
rect 4488 24123 4528 24155
rect 4560 24123 4600 24155
rect 4632 24123 4672 24155
rect 4704 24123 4744 24155
rect 4776 24123 4816 24155
rect 4848 24123 4888 24155
rect 4920 24123 4960 24155
rect 4992 24123 5032 24155
rect 5064 24123 5104 24155
rect 5136 24123 5176 24155
rect 5208 24123 5248 24155
rect 5280 24123 5320 24155
rect 5352 24123 5392 24155
rect 5424 24123 5464 24155
rect 5496 24123 5536 24155
rect 5568 24123 5608 24155
rect 5640 24123 5680 24155
rect 5712 24123 5752 24155
rect 5784 24123 5824 24155
rect 5856 24123 5896 24155
rect 5928 24123 5968 24155
rect 6000 24123 6040 24155
rect 6072 24123 6112 24155
rect 6144 24123 6184 24155
rect 6216 24123 6256 24155
rect 6288 24123 6328 24155
rect 6360 24123 6400 24155
rect 6432 24123 6472 24155
rect 6504 24123 6544 24155
rect 6576 24123 6616 24155
rect 6648 24123 6688 24155
rect 6720 24123 6760 24155
rect 6792 24123 6832 24155
rect 6864 24123 6904 24155
rect 6936 24123 6976 24155
rect 7008 24123 7048 24155
rect 7080 24123 7120 24155
rect 7152 24123 7192 24155
rect 7224 24123 7264 24155
rect 7296 24123 7336 24155
rect 7368 24123 7408 24155
rect 7440 24123 7480 24155
rect 7512 24123 7552 24155
rect 7584 24123 7624 24155
rect 7656 24123 7696 24155
rect 7728 24123 7768 24155
rect 7800 24123 7840 24155
rect 7872 24123 7912 24155
rect 7944 24123 7984 24155
rect 8016 24123 8056 24155
rect 8088 24123 8128 24155
rect 8160 24123 8200 24155
rect 8232 24123 8272 24155
rect 8304 24123 8344 24155
rect 8376 24123 8416 24155
rect 8448 24123 8488 24155
rect 8520 24123 8560 24155
rect 8592 24123 8632 24155
rect 8664 24123 8704 24155
rect 8736 24123 8776 24155
rect 8808 24123 8848 24155
rect 8880 24123 8920 24155
rect 8952 24123 8992 24155
rect 9024 24123 9064 24155
rect 9096 24123 9136 24155
rect 9168 24123 9208 24155
rect 9240 24123 9280 24155
rect 9312 24123 9352 24155
rect 9384 24123 9424 24155
rect 9456 24123 9496 24155
rect 9528 24123 9568 24155
rect 9600 24123 9640 24155
rect 9672 24123 9712 24155
rect 9744 24123 9784 24155
rect 9816 24123 9856 24155
rect 9888 24123 9928 24155
rect 9960 24123 10000 24155
rect 10032 24123 10072 24155
rect 10104 24123 10144 24155
rect 10176 24123 10216 24155
rect 10248 24123 10288 24155
rect 10320 24123 10360 24155
rect 10392 24123 10432 24155
rect 10464 24123 10504 24155
rect 10536 24123 10576 24155
rect 10608 24123 10648 24155
rect 10680 24123 10720 24155
rect 10752 24123 10792 24155
rect 10824 24123 10864 24155
rect 10896 24123 10936 24155
rect 10968 24123 11008 24155
rect 11040 24123 11080 24155
rect 11112 24123 11152 24155
rect 11184 24123 11224 24155
rect 11256 24123 11296 24155
rect 11328 24123 11368 24155
rect 11400 24123 11440 24155
rect 11472 24123 11512 24155
rect 11544 24123 11584 24155
rect 11616 24123 11656 24155
rect 11688 24123 11728 24155
rect 11760 24123 11800 24155
rect 11832 24123 11872 24155
rect 11904 24123 11944 24155
rect 11976 24123 12016 24155
rect 12048 24123 12088 24155
rect 12120 24123 12160 24155
rect 12192 24123 12232 24155
rect 12264 24123 12304 24155
rect 12336 24123 12376 24155
rect 12408 24123 12448 24155
rect 12480 24123 12520 24155
rect 12552 24123 12592 24155
rect 12624 24123 12664 24155
rect 12696 24123 12736 24155
rect 12768 24123 12808 24155
rect 12840 24123 12880 24155
rect 12912 24123 12952 24155
rect 12984 24123 13024 24155
rect 13056 24123 13096 24155
rect 13128 24123 13168 24155
rect 13200 24123 13240 24155
rect 13272 24123 13312 24155
rect 13344 24123 13384 24155
rect 13416 24123 13456 24155
rect 13488 24123 13528 24155
rect 13560 24123 13600 24155
rect 13632 24123 13672 24155
rect 13704 24123 13744 24155
rect 13776 24123 13816 24155
rect 13848 24123 13888 24155
rect 13920 24123 13960 24155
rect 13992 24123 14032 24155
rect 14064 24123 14104 24155
rect 14136 24123 14176 24155
rect 14208 24123 14248 24155
rect 14280 24123 14320 24155
rect 14352 24123 14392 24155
rect 14424 24123 14464 24155
rect 14496 24123 14536 24155
rect 14568 24123 14608 24155
rect 14640 24123 14680 24155
rect 14712 24123 14752 24155
rect 14784 24123 14824 24155
rect 14856 24123 14896 24155
rect 14928 24123 14968 24155
rect 15000 24123 15040 24155
rect 15072 24123 15112 24155
rect 15144 24123 15184 24155
rect 15216 24123 15256 24155
rect 15288 24123 15328 24155
rect 15360 24123 15400 24155
rect 15432 24123 15472 24155
rect 15504 24123 15544 24155
rect 15576 24123 15616 24155
rect 15648 24123 15688 24155
rect 15720 24123 15760 24155
rect 15792 24123 15832 24155
rect 15864 24123 15904 24155
rect 15936 24123 16000 24155
rect 0 24083 16000 24123
rect 0 24051 64 24083
rect 96 24051 136 24083
rect 168 24051 208 24083
rect 240 24051 280 24083
rect 312 24051 352 24083
rect 384 24051 424 24083
rect 456 24051 496 24083
rect 528 24051 568 24083
rect 600 24051 640 24083
rect 672 24051 712 24083
rect 744 24051 784 24083
rect 816 24051 856 24083
rect 888 24051 928 24083
rect 960 24051 1000 24083
rect 1032 24051 1072 24083
rect 1104 24051 1144 24083
rect 1176 24051 1216 24083
rect 1248 24051 1288 24083
rect 1320 24051 1360 24083
rect 1392 24051 1432 24083
rect 1464 24051 1504 24083
rect 1536 24051 1576 24083
rect 1608 24051 1648 24083
rect 1680 24051 1720 24083
rect 1752 24051 1792 24083
rect 1824 24051 1864 24083
rect 1896 24051 1936 24083
rect 1968 24051 2008 24083
rect 2040 24051 2080 24083
rect 2112 24051 2152 24083
rect 2184 24051 2224 24083
rect 2256 24051 2296 24083
rect 2328 24051 2368 24083
rect 2400 24051 2440 24083
rect 2472 24051 2512 24083
rect 2544 24051 2584 24083
rect 2616 24051 2656 24083
rect 2688 24051 2728 24083
rect 2760 24051 2800 24083
rect 2832 24051 2872 24083
rect 2904 24051 2944 24083
rect 2976 24051 3016 24083
rect 3048 24051 3088 24083
rect 3120 24051 3160 24083
rect 3192 24051 3232 24083
rect 3264 24051 3304 24083
rect 3336 24051 3376 24083
rect 3408 24051 3448 24083
rect 3480 24051 3520 24083
rect 3552 24051 3592 24083
rect 3624 24051 3664 24083
rect 3696 24051 3736 24083
rect 3768 24051 3808 24083
rect 3840 24051 3880 24083
rect 3912 24051 3952 24083
rect 3984 24051 4024 24083
rect 4056 24051 4096 24083
rect 4128 24051 4168 24083
rect 4200 24051 4240 24083
rect 4272 24051 4312 24083
rect 4344 24051 4384 24083
rect 4416 24051 4456 24083
rect 4488 24051 4528 24083
rect 4560 24051 4600 24083
rect 4632 24051 4672 24083
rect 4704 24051 4744 24083
rect 4776 24051 4816 24083
rect 4848 24051 4888 24083
rect 4920 24051 4960 24083
rect 4992 24051 5032 24083
rect 5064 24051 5104 24083
rect 5136 24051 5176 24083
rect 5208 24051 5248 24083
rect 5280 24051 5320 24083
rect 5352 24051 5392 24083
rect 5424 24051 5464 24083
rect 5496 24051 5536 24083
rect 5568 24051 5608 24083
rect 5640 24051 5680 24083
rect 5712 24051 5752 24083
rect 5784 24051 5824 24083
rect 5856 24051 5896 24083
rect 5928 24051 5968 24083
rect 6000 24051 6040 24083
rect 6072 24051 6112 24083
rect 6144 24051 6184 24083
rect 6216 24051 6256 24083
rect 6288 24051 6328 24083
rect 6360 24051 6400 24083
rect 6432 24051 6472 24083
rect 6504 24051 6544 24083
rect 6576 24051 6616 24083
rect 6648 24051 6688 24083
rect 6720 24051 6760 24083
rect 6792 24051 6832 24083
rect 6864 24051 6904 24083
rect 6936 24051 6976 24083
rect 7008 24051 7048 24083
rect 7080 24051 7120 24083
rect 7152 24051 7192 24083
rect 7224 24051 7264 24083
rect 7296 24051 7336 24083
rect 7368 24051 7408 24083
rect 7440 24051 7480 24083
rect 7512 24051 7552 24083
rect 7584 24051 7624 24083
rect 7656 24051 7696 24083
rect 7728 24051 7768 24083
rect 7800 24051 7840 24083
rect 7872 24051 7912 24083
rect 7944 24051 7984 24083
rect 8016 24051 8056 24083
rect 8088 24051 8128 24083
rect 8160 24051 8200 24083
rect 8232 24051 8272 24083
rect 8304 24051 8344 24083
rect 8376 24051 8416 24083
rect 8448 24051 8488 24083
rect 8520 24051 8560 24083
rect 8592 24051 8632 24083
rect 8664 24051 8704 24083
rect 8736 24051 8776 24083
rect 8808 24051 8848 24083
rect 8880 24051 8920 24083
rect 8952 24051 8992 24083
rect 9024 24051 9064 24083
rect 9096 24051 9136 24083
rect 9168 24051 9208 24083
rect 9240 24051 9280 24083
rect 9312 24051 9352 24083
rect 9384 24051 9424 24083
rect 9456 24051 9496 24083
rect 9528 24051 9568 24083
rect 9600 24051 9640 24083
rect 9672 24051 9712 24083
rect 9744 24051 9784 24083
rect 9816 24051 9856 24083
rect 9888 24051 9928 24083
rect 9960 24051 10000 24083
rect 10032 24051 10072 24083
rect 10104 24051 10144 24083
rect 10176 24051 10216 24083
rect 10248 24051 10288 24083
rect 10320 24051 10360 24083
rect 10392 24051 10432 24083
rect 10464 24051 10504 24083
rect 10536 24051 10576 24083
rect 10608 24051 10648 24083
rect 10680 24051 10720 24083
rect 10752 24051 10792 24083
rect 10824 24051 10864 24083
rect 10896 24051 10936 24083
rect 10968 24051 11008 24083
rect 11040 24051 11080 24083
rect 11112 24051 11152 24083
rect 11184 24051 11224 24083
rect 11256 24051 11296 24083
rect 11328 24051 11368 24083
rect 11400 24051 11440 24083
rect 11472 24051 11512 24083
rect 11544 24051 11584 24083
rect 11616 24051 11656 24083
rect 11688 24051 11728 24083
rect 11760 24051 11800 24083
rect 11832 24051 11872 24083
rect 11904 24051 11944 24083
rect 11976 24051 12016 24083
rect 12048 24051 12088 24083
rect 12120 24051 12160 24083
rect 12192 24051 12232 24083
rect 12264 24051 12304 24083
rect 12336 24051 12376 24083
rect 12408 24051 12448 24083
rect 12480 24051 12520 24083
rect 12552 24051 12592 24083
rect 12624 24051 12664 24083
rect 12696 24051 12736 24083
rect 12768 24051 12808 24083
rect 12840 24051 12880 24083
rect 12912 24051 12952 24083
rect 12984 24051 13024 24083
rect 13056 24051 13096 24083
rect 13128 24051 13168 24083
rect 13200 24051 13240 24083
rect 13272 24051 13312 24083
rect 13344 24051 13384 24083
rect 13416 24051 13456 24083
rect 13488 24051 13528 24083
rect 13560 24051 13600 24083
rect 13632 24051 13672 24083
rect 13704 24051 13744 24083
rect 13776 24051 13816 24083
rect 13848 24051 13888 24083
rect 13920 24051 13960 24083
rect 13992 24051 14032 24083
rect 14064 24051 14104 24083
rect 14136 24051 14176 24083
rect 14208 24051 14248 24083
rect 14280 24051 14320 24083
rect 14352 24051 14392 24083
rect 14424 24051 14464 24083
rect 14496 24051 14536 24083
rect 14568 24051 14608 24083
rect 14640 24051 14680 24083
rect 14712 24051 14752 24083
rect 14784 24051 14824 24083
rect 14856 24051 14896 24083
rect 14928 24051 14968 24083
rect 15000 24051 15040 24083
rect 15072 24051 15112 24083
rect 15144 24051 15184 24083
rect 15216 24051 15256 24083
rect 15288 24051 15328 24083
rect 15360 24051 15400 24083
rect 15432 24051 15472 24083
rect 15504 24051 15544 24083
rect 15576 24051 15616 24083
rect 15648 24051 15688 24083
rect 15720 24051 15760 24083
rect 15792 24051 15832 24083
rect 15864 24051 15904 24083
rect 15936 24051 16000 24083
rect 0 24011 16000 24051
rect 0 23979 64 24011
rect 96 23979 136 24011
rect 168 23979 208 24011
rect 240 23979 280 24011
rect 312 23979 352 24011
rect 384 23979 424 24011
rect 456 23979 496 24011
rect 528 23979 568 24011
rect 600 23979 640 24011
rect 672 23979 712 24011
rect 744 23979 784 24011
rect 816 23979 856 24011
rect 888 23979 928 24011
rect 960 23979 1000 24011
rect 1032 23979 1072 24011
rect 1104 23979 1144 24011
rect 1176 23979 1216 24011
rect 1248 23979 1288 24011
rect 1320 23979 1360 24011
rect 1392 23979 1432 24011
rect 1464 23979 1504 24011
rect 1536 23979 1576 24011
rect 1608 23979 1648 24011
rect 1680 23979 1720 24011
rect 1752 23979 1792 24011
rect 1824 23979 1864 24011
rect 1896 23979 1936 24011
rect 1968 23979 2008 24011
rect 2040 23979 2080 24011
rect 2112 23979 2152 24011
rect 2184 23979 2224 24011
rect 2256 23979 2296 24011
rect 2328 23979 2368 24011
rect 2400 23979 2440 24011
rect 2472 23979 2512 24011
rect 2544 23979 2584 24011
rect 2616 23979 2656 24011
rect 2688 23979 2728 24011
rect 2760 23979 2800 24011
rect 2832 23979 2872 24011
rect 2904 23979 2944 24011
rect 2976 23979 3016 24011
rect 3048 23979 3088 24011
rect 3120 23979 3160 24011
rect 3192 23979 3232 24011
rect 3264 23979 3304 24011
rect 3336 23979 3376 24011
rect 3408 23979 3448 24011
rect 3480 23979 3520 24011
rect 3552 23979 3592 24011
rect 3624 23979 3664 24011
rect 3696 23979 3736 24011
rect 3768 23979 3808 24011
rect 3840 23979 3880 24011
rect 3912 23979 3952 24011
rect 3984 23979 4024 24011
rect 4056 23979 4096 24011
rect 4128 23979 4168 24011
rect 4200 23979 4240 24011
rect 4272 23979 4312 24011
rect 4344 23979 4384 24011
rect 4416 23979 4456 24011
rect 4488 23979 4528 24011
rect 4560 23979 4600 24011
rect 4632 23979 4672 24011
rect 4704 23979 4744 24011
rect 4776 23979 4816 24011
rect 4848 23979 4888 24011
rect 4920 23979 4960 24011
rect 4992 23979 5032 24011
rect 5064 23979 5104 24011
rect 5136 23979 5176 24011
rect 5208 23979 5248 24011
rect 5280 23979 5320 24011
rect 5352 23979 5392 24011
rect 5424 23979 5464 24011
rect 5496 23979 5536 24011
rect 5568 23979 5608 24011
rect 5640 23979 5680 24011
rect 5712 23979 5752 24011
rect 5784 23979 5824 24011
rect 5856 23979 5896 24011
rect 5928 23979 5968 24011
rect 6000 23979 6040 24011
rect 6072 23979 6112 24011
rect 6144 23979 6184 24011
rect 6216 23979 6256 24011
rect 6288 23979 6328 24011
rect 6360 23979 6400 24011
rect 6432 23979 6472 24011
rect 6504 23979 6544 24011
rect 6576 23979 6616 24011
rect 6648 23979 6688 24011
rect 6720 23979 6760 24011
rect 6792 23979 6832 24011
rect 6864 23979 6904 24011
rect 6936 23979 6976 24011
rect 7008 23979 7048 24011
rect 7080 23979 7120 24011
rect 7152 23979 7192 24011
rect 7224 23979 7264 24011
rect 7296 23979 7336 24011
rect 7368 23979 7408 24011
rect 7440 23979 7480 24011
rect 7512 23979 7552 24011
rect 7584 23979 7624 24011
rect 7656 23979 7696 24011
rect 7728 23979 7768 24011
rect 7800 23979 7840 24011
rect 7872 23979 7912 24011
rect 7944 23979 7984 24011
rect 8016 23979 8056 24011
rect 8088 23979 8128 24011
rect 8160 23979 8200 24011
rect 8232 23979 8272 24011
rect 8304 23979 8344 24011
rect 8376 23979 8416 24011
rect 8448 23979 8488 24011
rect 8520 23979 8560 24011
rect 8592 23979 8632 24011
rect 8664 23979 8704 24011
rect 8736 23979 8776 24011
rect 8808 23979 8848 24011
rect 8880 23979 8920 24011
rect 8952 23979 8992 24011
rect 9024 23979 9064 24011
rect 9096 23979 9136 24011
rect 9168 23979 9208 24011
rect 9240 23979 9280 24011
rect 9312 23979 9352 24011
rect 9384 23979 9424 24011
rect 9456 23979 9496 24011
rect 9528 23979 9568 24011
rect 9600 23979 9640 24011
rect 9672 23979 9712 24011
rect 9744 23979 9784 24011
rect 9816 23979 9856 24011
rect 9888 23979 9928 24011
rect 9960 23979 10000 24011
rect 10032 23979 10072 24011
rect 10104 23979 10144 24011
rect 10176 23979 10216 24011
rect 10248 23979 10288 24011
rect 10320 23979 10360 24011
rect 10392 23979 10432 24011
rect 10464 23979 10504 24011
rect 10536 23979 10576 24011
rect 10608 23979 10648 24011
rect 10680 23979 10720 24011
rect 10752 23979 10792 24011
rect 10824 23979 10864 24011
rect 10896 23979 10936 24011
rect 10968 23979 11008 24011
rect 11040 23979 11080 24011
rect 11112 23979 11152 24011
rect 11184 23979 11224 24011
rect 11256 23979 11296 24011
rect 11328 23979 11368 24011
rect 11400 23979 11440 24011
rect 11472 23979 11512 24011
rect 11544 23979 11584 24011
rect 11616 23979 11656 24011
rect 11688 23979 11728 24011
rect 11760 23979 11800 24011
rect 11832 23979 11872 24011
rect 11904 23979 11944 24011
rect 11976 23979 12016 24011
rect 12048 23979 12088 24011
rect 12120 23979 12160 24011
rect 12192 23979 12232 24011
rect 12264 23979 12304 24011
rect 12336 23979 12376 24011
rect 12408 23979 12448 24011
rect 12480 23979 12520 24011
rect 12552 23979 12592 24011
rect 12624 23979 12664 24011
rect 12696 23979 12736 24011
rect 12768 23979 12808 24011
rect 12840 23979 12880 24011
rect 12912 23979 12952 24011
rect 12984 23979 13024 24011
rect 13056 23979 13096 24011
rect 13128 23979 13168 24011
rect 13200 23979 13240 24011
rect 13272 23979 13312 24011
rect 13344 23979 13384 24011
rect 13416 23979 13456 24011
rect 13488 23979 13528 24011
rect 13560 23979 13600 24011
rect 13632 23979 13672 24011
rect 13704 23979 13744 24011
rect 13776 23979 13816 24011
rect 13848 23979 13888 24011
rect 13920 23979 13960 24011
rect 13992 23979 14032 24011
rect 14064 23979 14104 24011
rect 14136 23979 14176 24011
rect 14208 23979 14248 24011
rect 14280 23979 14320 24011
rect 14352 23979 14392 24011
rect 14424 23979 14464 24011
rect 14496 23979 14536 24011
rect 14568 23979 14608 24011
rect 14640 23979 14680 24011
rect 14712 23979 14752 24011
rect 14784 23979 14824 24011
rect 14856 23979 14896 24011
rect 14928 23979 14968 24011
rect 15000 23979 15040 24011
rect 15072 23979 15112 24011
rect 15144 23979 15184 24011
rect 15216 23979 15256 24011
rect 15288 23979 15328 24011
rect 15360 23979 15400 24011
rect 15432 23979 15472 24011
rect 15504 23979 15544 24011
rect 15576 23979 15616 24011
rect 15648 23979 15688 24011
rect 15720 23979 15760 24011
rect 15792 23979 15832 24011
rect 15864 23979 15904 24011
rect 15936 23979 16000 24011
rect 0 23939 16000 23979
rect 0 23907 64 23939
rect 96 23907 136 23939
rect 168 23907 208 23939
rect 240 23907 280 23939
rect 312 23907 352 23939
rect 384 23907 424 23939
rect 456 23907 496 23939
rect 528 23907 568 23939
rect 600 23907 640 23939
rect 672 23907 712 23939
rect 744 23907 784 23939
rect 816 23907 856 23939
rect 888 23907 928 23939
rect 960 23907 1000 23939
rect 1032 23907 1072 23939
rect 1104 23907 1144 23939
rect 1176 23907 1216 23939
rect 1248 23907 1288 23939
rect 1320 23907 1360 23939
rect 1392 23907 1432 23939
rect 1464 23907 1504 23939
rect 1536 23907 1576 23939
rect 1608 23907 1648 23939
rect 1680 23907 1720 23939
rect 1752 23907 1792 23939
rect 1824 23907 1864 23939
rect 1896 23907 1936 23939
rect 1968 23907 2008 23939
rect 2040 23907 2080 23939
rect 2112 23907 2152 23939
rect 2184 23907 2224 23939
rect 2256 23907 2296 23939
rect 2328 23907 2368 23939
rect 2400 23907 2440 23939
rect 2472 23907 2512 23939
rect 2544 23907 2584 23939
rect 2616 23907 2656 23939
rect 2688 23907 2728 23939
rect 2760 23907 2800 23939
rect 2832 23907 2872 23939
rect 2904 23907 2944 23939
rect 2976 23907 3016 23939
rect 3048 23907 3088 23939
rect 3120 23907 3160 23939
rect 3192 23907 3232 23939
rect 3264 23907 3304 23939
rect 3336 23907 3376 23939
rect 3408 23907 3448 23939
rect 3480 23907 3520 23939
rect 3552 23907 3592 23939
rect 3624 23907 3664 23939
rect 3696 23907 3736 23939
rect 3768 23907 3808 23939
rect 3840 23907 3880 23939
rect 3912 23907 3952 23939
rect 3984 23907 4024 23939
rect 4056 23907 4096 23939
rect 4128 23907 4168 23939
rect 4200 23907 4240 23939
rect 4272 23907 4312 23939
rect 4344 23907 4384 23939
rect 4416 23907 4456 23939
rect 4488 23907 4528 23939
rect 4560 23907 4600 23939
rect 4632 23907 4672 23939
rect 4704 23907 4744 23939
rect 4776 23907 4816 23939
rect 4848 23907 4888 23939
rect 4920 23907 4960 23939
rect 4992 23907 5032 23939
rect 5064 23907 5104 23939
rect 5136 23907 5176 23939
rect 5208 23907 5248 23939
rect 5280 23907 5320 23939
rect 5352 23907 5392 23939
rect 5424 23907 5464 23939
rect 5496 23907 5536 23939
rect 5568 23907 5608 23939
rect 5640 23907 5680 23939
rect 5712 23907 5752 23939
rect 5784 23907 5824 23939
rect 5856 23907 5896 23939
rect 5928 23907 5968 23939
rect 6000 23907 6040 23939
rect 6072 23907 6112 23939
rect 6144 23907 6184 23939
rect 6216 23907 6256 23939
rect 6288 23907 6328 23939
rect 6360 23907 6400 23939
rect 6432 23907 6472 23939
rect 6504 23907 6544 23939
rect 6576 23907 6616 23939
rect 6648 23907 6688 23939
rect 6720 23907 6760 23939
rect 6792 23907 6832 23939
rect 6864 23907 6904 23939
rect 6936 23907 6976 23939
rect 7008 23907 7048 23939
rect 7080 23907 7120 23939
rect 7152 23907 7192 23939
rect 7224 23907 7264 23939
rect 7296 23907 7336 23939
rect 7368 23907 7408 23939
rect 7440 23907 7480 23939
rect 7512 23907 7552 23939
rect 7584 23907 7624 23939
rect 7656 23907 7696 23939
rect 7728 23907 7768 23939
rect 7800 23907 7840 23939
rect 7872 23907 7912 23939
rect 7944 23907 7984 23939
rect 8016 23907 8056 23939
rect 8088 23907 8128 23939
rect 8160 23907 8200 23939
rect 8232 23907 8272 23939
rect 8304 23907 8344 23939
rect 8376 23907 8416 23939
rect 8448 23907 8488 23939
rect 8520 23907 8560 23939
rect 8592 23907 8632 23939
rect 8664 23907 8704 23939
rect 8736 23907 8776 23939
rect 8808 23907 8848 23939
rect 8880 23907 8920 23939
rect 8952 23907 8992 23939
rect 9024 23907 9064 23939
rect 9096 23907 9136 23939
rect 9168 23907 9208 23939
rect 9240 23907 9280 23939
rect 9312 23907 9352 23939
rect 9384 23907 9424 23939
rect 9456 23907 9496 23939
rect 9528 23907 9568 23939
rect 9600 23907 9640 23939
rect 9672 23907 9712 23939
rect 9744 23907 9784 23939
rect 9816 23907 9856 23939
rect 9888 23907 9928 23939
rect 9960 23907 10000 23939
rect 10032 23907 10072 23939
rect 10104 23907 10144 23939
rect 10176 23907 10216 23939
rect 10248 23907 10288 23939
rect 10320 23907 10360 23939
rect 10392 23907 10432 23939
rect 10464 23907 10504 23939
rect 10536 23907 10576 23939
rect 10608 23907 10648 23939
rect 10680 23907 10720 23939
rect 10752 23907 10792 23939
rect 10824 23907 10864 23939
rect 10896 23907 10936 23939
rect 10968 23907 11008 23939
rect 11040 23907 11080 23939
rect 11112 23907 11152 23939
rect 11184 23907 11224 23939
rect 11256 23907 11296 23939
rect 11328 23907 11368 23939
rect 11400 23907 11440 23939
rect 11472 23907 11512 23939
rect 11544 23907 11584 23939
rect 11616 23907 11656 23939
rect 11688 23907 11728 23939
rect 11760 23907 11800 23939
rect 11832 23907 11872 23939
rect 11904 23907 11944 23939
rect 11976 23907 12016 23939
rect 12048 23907 12088 23939
rect 12120 23907 12160 23939
rect 12192 23907 12232 23939
rect 12264 23907 12304 23939
rect 12336 23907 12376 23939
rect 12408 23907 12448 23939
rect 12480 23907 12520 23939
rect 12552 23907 12592 23939
rect 12624 23907 12664 23939
rect 12696 23907 12736 23939
rect 12768 23907 12808 23939
rect 12840 23907 12880 23939
rect 12912 23907 12952 23939
rect 12984 23907 13024 23939
rect 13056 23907 13096 23939
rect 13128 23907 13168 23939
rect 13200 23907 13240 23939
rect 13272 23907 13312 23939
rect 13344 23907 13384 23939
rect 13416 23907 13456 23939
rect 13488 23907 13528 23939
rect 13560 23907 13600 23939
rect 13632 23907 13672 23939
rect 13704 23907 13744 23939
rect 13776 23907 13816 23939
rect 13848 23907 13888 23939
rect 13920 23907 13960 23939
rect 13992 23907 14032 23939
rect 14064 23907 14104 23939
rect 14136 23907 14176 23939
rect 14208 23907 14248 23939
rect 14280 23907 14320 23939
rect 14352 23907 14392 23939
rect 14424 23907 14464 23939
rect 14496 23907 14536 23939
rect 14568 23907 14608 23939
rect 14640 23907 14680 23939
rect 14712 23907 14752 23939
rect 14784 23907 14824 23939
rect 14856 23907 14896 23939
rect 14928 23907 14968 23939
rect 15000 23907 15040 23939
rect 15072 23907 15112 23939
rect 15144 23907 15184 23939
rect 15216 23907 15256 23939
rect 15288 23907 15328 23939
rect 15360 23907 15400 23939
rect 15432 23907 15472 23939
rect 15504 23907 15544 23939
rect 15576 23907 15616 23939
rect 15648 23907 15688 23939
rect 15720 23907 15760 23939
rect 15792 23907 15832 23939
rect 15864 23907 15904 23939
rect 15936 23907 16000 23939
rect 0 23867 16000 23907
rect 0 23835 64 23867
rect 96 23835 136 23867
rect 168 23835 208 23867
rect 240 23835 280 23867
rect 312 23835 352 23867
rect 384 23835 424 23867
rect 456 23835 496 23867
rect 528 23835 568 23867
rect 600 23835 640 23867
rect 672 23835 712 23867
rect 744 23835 784 23867
rect 816 23835 856 23867
rect 888 23835 928 23867
rect 960 23835 1000 23867
rect 1032 23835 1072 23867
rect 1104 23835 1144 23867
rect 1176 23835 1216 23867
rect 1248 23835 1288 23867
rect 1320 23835 1360 23867
rect 1392 23835 1432 23867
rect 1464 23835 1504 23867
rect 1536 23835 1576 23867
rect 1608 23835 1648 23867
rect 1680 23835 1720 23867
rect 1752 23835 1792 23867
rect 1824 23835 1864 23867
rect 1896 23835 1936 23867
rect 1968 23835 2008 23867
rect 2040 23835 2080 23867
rect 2112 23835 2152 23867
rect 2184 23835 2224 23867
rect 2256 23835 2296 23867
rect 2328 23835 2368 23867
rect 2400 23835 2440 23867
rect 2472 23835 2512 23867
rect 2544 23835 2584 23867
rect 2616 23835 2656 23867
rect 2688 23835 2728 23867
rect 2760 23835 2800 23867
rect 2832 23835 2872 23867
rect 2904 23835 2944 23867
rect 2976 23835 3016 23867
rect 3048 23835 3088 23867
rect 3120 23835 3160 23867
rect 3192 23835 3232 23867
rect 3264 23835 3304 23867
rect 3336 23835 3376 23867
rect 3408 23835 3448 23867
rect 3480 23835 3520 23867
rect 3552 23835 3592 23867
rect 3624 23835 3664 23867
rect 3696 23835 3736 23867
rect 3768 23835 3808 23867
rect 3840 23835 3880 23867
rect 3912 23835 3952 23867
rect 3984 23835 4024 23867
rect 4056 23835 4096 23867
rect 4128 23835 4168 23867
rect 4200 23835 4240 23867
rect 4272 23835 4312 23867
rect 4344 23835 4384 23867
rect 4416 23835 4456 23867
rect 4488 23835 4528 23867
rect 4560 23835 4600 23867
rect 4632 23835 4672 23867
rect 4704 23835 4744 23867
rect 4776 23835 4816 23867
rect 4848 23835 4888 23867
rect 4920 23835 4960 23867
rect 4992 23835 5032 23867
rect 5064 23835 5104 23867
rect 5136 23835 5176 23867
rect 5208 23835 5248 23867
rect 5280 23835 5320 23867
rect 5352 23835 5392 23867
rect 5424 23835 5464 23867
rect 5496 23835 5536 23867
rect 5568 23835 5608 23867
rect 5640 23835 5680 23867
rect 5712 23835 5752 23867
rect 5784 23835 5824 23867
rect 5856 23835 5896 23867
rect 5928 23835 5968 23867
rect 6000 23835 6040 23867
rect 6072 23835 6112 23867
rect 6144 23835 6184 23867
rect 6216 23835 6256 23867
rect 6288 23835 6328 23867
rect 6360 23835 6400 23867
rect 6432 23835 6472 23867
rect 6504 23835 6544 23867
rect 6576 23835 6616 23867
rect 6648 23835 6688 23867
rect 6720 23835 6760 23867
rect 6792 23835 6832 23867
rect 6864 23835 6904 23867
rect 6936 23835 6976 23867
rect 7008 23835 7048 23867
rect 7080 23835 7120 23867
rect 7152 23835 7192 23867
rect 7224 23835 7264 23867
rect 7296 23835 7336 23867
rect 7368 23835 7408 23867
rect 7440 23835 7480 23867
rect 7512 23835 7552 23867
rect 7584 23835 7624 23867
rect 7656 23835 7696 23867
rect 7728 23835 7768 23867
rect 7800 23835 7840 23867
rect 7872 23835 7912 23867
rect 7944 23835 7984 23867
rect 8016 23835 8056 23867
rect 8088 23835 8128 23867
rect 8160 23835 8200 23867
rect 8232 23835 8272 23867
rect 8304 23835 8344 23867
rect 8376 23835 8416 23867
rect 8448 23835 8488 23867
rect 8520 23835 8560 23867
rect 8592 23835 8632 23867
rect 8664 23835 8704 23867
rect 8736 23835 8776 23867
rect 8808 23835 8848 23867
rect 8880 23835 8920 23867
rect 8952 23835 8992 23867
rect 9024 23835 9064 23867
rect 9096 23835 9136 23867
rect 9168 23835 9208 23867
rect 9240 23835 9280 23867
rect 9312 23835 9352 23867
rect 9384 23835 9424 23867
rect 9456 23835 9496 23867
rect 9528 23835 9568 23867
rect 9600 23835 9640 23867
rect 9672 23835 9712 23867
rect 9744 23835 9784 23867
rect 9816 23835 9856 23867
rect 9888 23835 9928 23867
rect 9960 23835 10000 23867
rect 10032 23835 10072 23867
rect 10104 23835 10144 23867
rect 10176 23835 10216 23867
rect 10248 23835 10288 23867
rect 10320 23835 10360 23867
rect 10392 23835 10432 23867
rect 10464 23835 10504 23867
rect 10536 23835 10576 23867
rect 10608 23835 10648 23867
rect 10680 23835 10720 23867
rect 10752 23835 10792 23867
rect 10824 23835 10864 23867
rect 10896 23835 10936 23867
rect 10968 23835 11008 23867
rect 11040 23835 11080 23867
rect 11112 23835 11152 23867
rect 11184 23835 11224 23867
rect 11256 23835 11296 23867
rect 11328 23835 11368 23867
rect 11400 23835 11440 23867
rect 11472 23835 11512 23867
rect 11544 23835 11584 23867
rect 11616 23835 11656 23867
rect 11688 23835 11728 23867
rect 11760 23835 11800 23867
rect 11832 23835 11872 23867
rect 11904 23835 11944 23867
rect 11976 23835 12016 23867
rect 12048 23835 12088 23867
rect 12120 23835 12160 23867
rect 12192 23835 12232 23867
rect 12264 23835 12304 23867
rect 12336 23835 12376 23867
rect 12408 23835 12448 23867
rect 12480 23835 12520 23867
rect 12552 23835 12592 23867
rect 12624 23835 12664 23867
rect 12696 23835 12736 23867
rect 12768 23835 12808 23867
rect 12840 23835 12880 23867
rect 12912 23835 12952 23867
rect 12984 23835 13024 23867
rect 13056 23835 13096 23867
rect 13128 23835 13168 23867
rect 13200 23835 13240 23867
rect 13272 23835 13312 23867
rect 13344 23835 13384 23867
rect 13416 23835 13456 23867
rect 13488 23835 13528 23867
rect 13560 23835 13600 23867
rect 13632 23835 13672 23867
rect 13704 23835 13744 23867
rect 13776 23835 13816 23867
rect 13848 23835 13888 23867
rect 13920 23835 13960 23867
rect 13992 23835 14032 23867
rect 14064 23835 14104 23867
rect 14136 23835 14176 23867
rect 14208 23835 14248 23867
rect 14280 23835 14320 23867
rect 14352 23835 14392 23867
rect 14424 23835 14464 23867
rect 14496 23835 14536 23867
rect 14568 23835 14608 23867
rect 14640 23835 14680 23867
rect 14712 23835 14752 23867
rect 14784 23835 14824 23867
rect 14856 23835 14896 23867
rect 14928 23835 14968 23867
rect 15000 23835 15040 23867
rect 15072 23835 15112 23867
rect 15144 23835 15184 23867
rect 15216 23835 15256 23867
rect 15288 23835 15328 23867
rect 15360 23835 15400 23867
rect 15432 23835 15472 23867
rect 15504 23835 15544 23867
rect 15576 23835 15616 23867
rect 15648 23835 15688 23867
rect 15720 23835 15760 23867
rect 15792 23835 15832 23867
rect 15864 23835 15904 23867
rect 15936 23835 16000 23867
rect 0 23795 16000 23835
rect 0 23763 64 23795
rect 96 23763 136 23795
rect 168 23763 208 23795
rect 240 23763 280 23795
rect 312 23763 352 23795
rect 384 23763 424 23795
rect 456 23763 496 23795
rect 528 23763 568 23795
rect 600 23763 640 23795
rect 672 23763 712 23795
rect 744 23763 784 23795
rect 816 23763 856 23795
rect 888 23763 928 23795
rect 960 23763 1000 23795
rect 1032 23763 1072 23795
rect 1104 23763 1144 23795
rect 1176 23763 1216 23795
rect 1248 23763 1288 23795
rect 1320 23763 1360 23795
rect 1392 23763 1432 23795
rect 1464 23763 1504 23795
rect 1536 23763 1576 23795
rect 1608 23763 1648 23795
rect 1680 23763 1720 23795
rect 1752 23763 1792 23795
rect 1824 23763 1864 23795
rect 1896 23763 1936 23795
rect 1968 23763 2008 23795
rect 2040 23763 2080 23795
rect 2112 23763 2152 23795
rect 2184 23763 2224 23795
rect 2256 23763 2296 23795
rect 2328 23763 2368 23795
rect 2400 23763 2440 23795
rect 2472 23763 2512 23795
rect 2544 23763 2584 23795
rect 2616 23763 2656 23795
rect 2688 23763 2728 23795
rect 2760 23763 2800 23795
rect 2832 23763 2872 23795
rect 2904 23763 2944 23795
rect 2976 23763 3016 23795
rect 3048 23763 3088 23795
rect 3120 23763 3160 23795
rect 3192 23763 3232 23795
rect 3264 23763 3304 23795
rect 3336 23763 3376 23795
rect 3408 23763 3448 23795
rect 3480 23763 3520 23795
rect 3552 23763 3592 23795
rect 3624 23763 3664 23795
rect 3696 23763 3736 23795
rect 3768 23763 3808 23795
rect 3840 23763 3880 23795
rect 3912 23763 3952 23795
rect 3984 23763 4024 23795
rect 4056 23763 4096 23795
rect 4128 23763 4168 23795
rect 4200 23763 4240 23795
rect 4272 23763 4312 23795
rect 4344 23763 4384 23795
rect 4416 23763 4456 23795
rect 4488 23763 4528 23795
rect 4560 23763 4600 23795
rect 4632 23763 4672 23795
rect 4704 23763 4744 23795
rect 4776 23763 4816 23795
rect 4848 23763 4888 23795
rect 4920 23763 4960 23795
rect 4992 23763 5032 23795
rect 5064 23763 5104 23795
rect 5136 23763 5176 23795
rect 5208 23763 5248 23795
rect 5280 23763 5320 23795
rect 5352 23763 5392 23795
rect 5424 23763 5464 23795
rect 5496 23763 5536 23795
rect 5568 23763 5608 23795
rect 5640 23763 5680 23795
rect 5712 23763 5752 23795
rect 5784 23763 5824 23795
rect 5856 23763 5896 23795
rect 5928 23763 5968 23795
rect 6000 23763 6040 23795
rect 6072 23763 6112 23795
rect 6144 23763 6184 23795
rect 6216 23763 6256 23795
rect 6288 23763 6328 23795
rect 6360 23763 6400 23795
rect 6432 23763 6472 23795
rect 6504 23763 6544 23795
rect 6576 23763 6616 23795
rect 6648 23763 6688 23795
rect 6720 23763 6760 23795
rect 6792 23763 6832 23795
rect 6864 23763 6904 23795
rect 6936 23763 6976 23795
rect 7008 23763 7048 23795
rect 7080 23763 7120 23795
rect 7152 23763 7192 23795
rect 7224 23763 7264 23795
rect 7296 23763 7336 23795
rect 7368 23763 7408 23795
rect 7440 23763 7480 23795
rect 7512 23763 7552 23795
rect 7584 23763 7624 23795
rect 7656 23763 7696 23795
rect 7728 23763 7768 23795
rect 7800 23763 7840 23795
rect 7872 23763 7912 23795
rect 7944 23763 7984 23795
rect 8016 23763 8056 23795
rect 8088 23763 8128 23795
rect 8160 23763 8200 23795
rect 8232 23763 8272 23795
rect 8304 23763 8344 23795
rect 8376 23763 8416 23795
rect 8448 23763 8488 23795
rect 8520 23763 8560 23795
rect 8592 23763 8632 23795
rect 8664 23763 8704 23795
rect 8736 23763 8776 23795
rect 8808 23763 8848 23795
rect 8880 23763 8920 23795
rect 8952 23763 8992 23795
rect 9024 23763 9064 23795
rect 9096 23763 9136 23795
rect 9168 23763 9208 23795
rect 9240 23763 9280 23795
rect 9312 23763 9352 23795
rect 9384 23763 9424 23795
rect 9456 23763 9496 23795
rect 9528 23763 9568 23795
rect 9600 23763 9640 23795
rect 9672 23763 9712 23795
rect 9744 23763 9784 23795
rect 9816 23763 9856 23795
rect 9888 23763 9928 23795
rect 9960 23763 10000 23795
rect 10032 23763 10072 23795
rect 10104 23763 10144 23795
rect 10176 23763 10216 23795
rect 10248 23763 10288 23795
rect 10320 23763 10360 23795
rect 10392 23763 10432 23795
rect 10464 23763 10504 23795
rect 10536 23763 10576 23795
rect 10608 23763 10648 23795
rect 10680 23763 10720 23795
rect 10752 23763 10792 23795
rect 10824 23763 10864 23795
rect 10896 23763 10936 23795
rect 10968 23763 11008 23795
rect 11040 23763 11080 23795
rect 11112 23763 11152 23795
rect 11184 23763 11224 23795
rect 11256 23763 11296 23795
rect 11328 23763 11368 23795
rect 11400 23763 11440 23795
rect 11472 23763 11512 23795
rect 11544 23763 11584 23795
rect 11616 23763 11656 23795
rect 11688 23763 11728 23795
rect 11760 23763 11800 23795
rect 11832 23763 11872 23795
rect 11904 23763 11944 23795
rect 11976 23763 12016 23795
rect 12048 23763 12088 23795
rect 12120 23763 12160 23795
rect 12192 23763 12232 23795
rect 12264 23763 12304 23795
rect 12336 23763 12376 23795
rect 12408 23763 12448 23795
rect 12480 23763 12520 23795
rect 12552 23763 12592 23795
rect 12624 23763 12664 23795
rect 12696 23763 12736 23795
rect 12768 23763 12808 23795
rect 12840 23763 12880 23795
rect 12912 23763 12952 23795
rect 12984 23763 13024 23795
rect 13056 23763 13096 23795
rect 13128 23763 13168 23795
rect 13200 23763 13240 23795
rect 13272 23763 13312 23795
rect 13344 23763 13384 23795
rect 13416 23763 13456 23795
rect 13488 23763 13528 23795
rect 13560 23763 13600 23795
rect 13632 23763 13672 23795
rect 13704 23763 13744 23795
rect 13776 23763 13816 23795
rect 13848 23763 13888 23795
rect 13920 23763 13960 23795
rect 13992 23763 14032 23795
rect 14064 23763 14104 23795
rect 14136 23763 14176 23795
rect 14208 23763 14248 23795
rect 14280 23763 14320 23795
rect 14352 23763 14392 23795
rect 14424 23763 14464 23795
rect 14496 23763 14536 23795
rect 14568 23763 14608 23795
rect 14640 23763 14680 23795
rect 14712 23763 14752 23795
rect 14784 23763 14824 23795
rect 14856 23763 14896 23795
rect 14928 23763 14968 23795
rect 15000 23763 15040 23795
rect 15072 23763 15112 23795
rect 15144 23763 15184 23795
rect 15216 23763 15256 23795
rect 15288 23763 15328 23795
rect 15360 23763 15400 23795
rect 15432 23763 15472 23795
rect 15504 23763 15544 23795
rect 15576 23763 15616 23795
rect 15648 23763 15688 23795
rect 15720 23763 15760 23795
rect 15792 23763 15832 23795
rect 15864 23763 15904 23795
rect 15936 23763 16000 23795
rect 0 23723 16000 23763
rect 0 23691 64 23723
rect 96 23691 136 23723
rect 168 23691 208 23723
rect 240 23691 280 23723
rect 312 23691 352 23723
rect 384 23691 424 23723
rect 456 23691 496 23723
rect 528 23691 568 23723
rect 600 23691 640 23723
rect 672 23691 712 23723
rect 744 23691 784 23723
rect 816 23691 856 23723
rect 888 23691 928 23723
rect 960 23691 1000 23723
rect 1032 23691 1072 23723
rect 1104 23691 1144 23723
rect 1176 23691 1216 23723
rect 1248 23691 1288 23723
rect 1320 23691 1360 23723
rect 1392 23691 1432 23723
rect 1464 23691 1504 23723
rect 1536 23691 1576 23723
rect 1608 23691 1648 23723
rect 1680 23691 1720 23723
rect 1752 23691 1792 23723
rect 1824 23691 1864 23723
rect 1896 23691 1936 23723
rect 1968 23691 2008 23723
rect 2040 23691 2080 23723
rect 2112 23691 2152 23723
rect 2184 23691 2224 23723
rect 2256 23691 2296 23723
rect 2328 23691 2368 23723
rect 2400 23691 2440 23723
rect 2472 23691 2512 23723
rect 2544 23691 2584 23723
rect 2616 23691 2656 23723
rect 2688 23691 2728 23723
rect 2760 23691 2800 23723
rect 2832 23691 2872 23723
rect 2904 23691 2944 23723
rect 2976 23691 3016 23723
rect 3048 23691 3088 23723
rect 3120 23691 3160 23723
rect 3192 23691 3232 23723
rect 3264 23691 3304 23723
rect 3336 23691 3376 23723
rect 3408 23691 3448 23723
rect 3480 23691 3520 23723
rect 3552 23691 3592 23723
rect 3624 23691 3664 23723
rect 3696 23691 3736 23723
rect 3768 23691 3808 23723
rect 3840 23691 3880 23723
rect 3912 23691 3952 23723
rect 3984 23691 4024 23723
rect 4056 23691 4096 23723
rect 4128 23691 4168 23723
rect 4200 23691 4240 23723
rect 4272 23691 4312 23723
rect 4344 23691 4384 23723
rect 4416 23691 4456 23723
rect 4488 23691 4528 23723
rect 4560 23691 4600 23723
rect 4632 23691 4672 23723
rect 4704 23691 4744 23723
rect 4776 23691 4816 23723
rect 4848 23691 4888 23723
rect 4920 23691 4960 23723
rect 4992 23691 5032 23723
rect 5064 23691 5104 23723
rect 5136 23691 5176 23723
rect 5208 23691 5248 23723
rect 5280 23691 5320 23723
rect 5352 23691 5392 23723
rect 5424 23691 5464 23723
rect 5496 23691 5536 23723
rect 5568 23691 5608 23723
rect 5640 23691 5680 23723
rect 5712 23691 5752 23723
rect 5784 23691 5824 23723
rect 5856 23691 5896 23723
rect 5928 23691 5968 23723
rect 6000 23691 6040 23723
rect 6072 23691 6112 23723
rect 6144 23691 6184 23723
rect 6216 23691 6256 23723
rect 6288 23691 6328 23723
rect 6360 23691 6400 23723
rect 6432 23691 6472 23723
rect 6504 23691 6544 23723
rect 6576 23691 6616 23723
rect 6648 23691 6688 23723
rect 6720 23691 6760 23723
rect 6792 23691 6832 23723
rect 6864 23691 6904 23723
rect 6936 23691 6976 23723
rect 7008 23691 7048 23723
rect 7080 23691 7120 23723
rect 7152 23691 7192 23723
rect 7224 23691 7264 23723
rect 7296 23691 7336 23723
rect 7368 23691 7408 23723
rect 7440 23691 7480 23723
rect 7512 23691 7552 23723
rect 7584 23691 7624 23723
rect 7656 23691 7696 23723
rect 7728 23691 7768 23723
rect 7800 23691 7840 23723
rect 7872 23691 7912 23723
rect 7944 23691 7984 23723
rect 8016 23691 8056 23723
rect 8088 23691 8128 23723
rect 8160 23691 8200 23723
rect 8232 23691 8272 23723
rect 8304 23691 8344 23723
rect 8376 23691 8416 23723
rect 8448 23691 8488 23723
rect 8520 23691 8560 23723
rect 8592 23691 8632 23723
rect 8664 23691 8704 23723
rect 8736 23691 8776 23723
rect 8808 23691 8848 23723
rect 8880 23691 8920 23723
rect 8952 23691 8992 23723
rect 9024 23691 9064 23723
rect 9096 23691 9136 23723
rect 9168 23691 9208 23723
rect 9240 23691 9280 23723
rect 9312 23691 9352 23723
rect 9384 23691 9424 23723
rect 9456 23691 9496 23723
rect 9528 23691 9568 23723
rect 9600 23691 9640 23723
rect 9672 23691 9712 23723
rect 9744 23691 9784 23723
rect 9816 23691 9856 23723
rect 9888 23691 9928 23723
rect 9960 23691 10000 23723
rect 10032 23691 10072 23723
rect 10104 23691 10144 23723
rect 10176 23691 10216 23723
rect 10248 23691 10288 23723
rect 10320 23691 10360 23723
rect 10392 23691 10432 23723
rect 10464 23691 10504 23723
rect 10536 23691 10576 23723
rect 10608 23691 10648 23723
rect 10680 23691 10720 23723
rect 10752 23691 10792 23723
rect 10824 23691 10864 23723
rect 10896 23691 10936 23723
rect 10968 23691 11008 23723
rect 11040 23691 11080 23723
rect 11112 23691 11152 23723
rect 11184 23691 11224 23723
rect 11256 23691 11296 23723
rect 11328 23691 11368 23723
rect 11400 23691 11440 23723
rect 11472 23691 11512 23723
rect 11544 23691 11584 23723
rect 11616 23691 11656 23723
rect 11688 23691 11728 23723
rect 11760 23691 11800 23723
rect 11832 23691 11872 23723
rect 11904 23691 11944 23723
rect 11976 23691 12016 23723
rect 12048 23691 12088 23723
rect 12120 23691 12160 23723
rect 12192 23691 12232 23723
rect 12264 23691 12304 23723
rect 12336 23691 12376 23723
rect 12408 23691 12448 23723
rect 12480 23691 12520 23723
rect 12552 23691 12592 23723
rect 12624 23691 12664 23723
rect 12696 23691 12736 23723
rect 12768 23691 12808 23723
rect 12840 23691 12880 23723
rect 12912 23691 12952 23723
rect 12984 23691 13024 23723
rect 13056 23691 13096 23723
rect 13128 23691 13168 23723
rect 13200 23691 13240 23723
rect 13272 23691 13312 23723
rect 13344 23691 13384 23723
rect 13416 23691 13456 23723
rect 13488 23691 13528 23723
rect 13560 23691 13600 23723
rect 13632 23691 13672 23723
rect 13704 23691 13744 23723
rect 13776 23691 13816 23723
rect 13848 23691 13888 23723
rect 13920 23691 13960 23723
rect 13992 23691 14032 23723
rect 14064 23691 14104 23723
rect 14136 23691 14176 23723
rect 14208 23691 14248 23723
rect 14280 23691 14320 23723
rect 14352 23691 14392 23723
rect 14424 23691 14464 23723
rect 14496 23691 14536 23723
rect 14568 23691 14608 23723
rect 14640 23691 14680 23723
rect 14712 23691 14752 23723
rect 14784 23691 14824 23723
rect 14856 23691 14896 23723
rect 14928 23691 14968 23723
rect 15000 23691 15040 23723
rect 15072 23691 15112 23723
rect 15144 23691 15184 23723
rect 15216 23691 15256 23723
rect 15288 23691 15328 23723
rect 15360 23691 15400 23723
rect 15432 23691 15472 23723
rect 15504 23691 15544 23723
rect 15576 23691 15616 23723
rect 15648 23691 15688 23723
rect 15720 23691 15760 23723
rect 15792 23691 15832 23723
rect 15864 23691 15904 23723
rect 15936 23691 16000 23723
rect 0 23651 16000 23691
rect 0 23619 64 23651
rect 96 23619 136 23651
rect 168 23619 208 23651
rect 240 23619 280 23651
rect 312 23619 352 23651
rect 384 23619 424 23651
rect 456 23619 496 23651
rect 528 23619 568 23651
rect 600 23619 640 23651
rect 672 23619 712 23651
rect 744 23619 784 23651
rect 816 23619 856 23651
rect 888 23619 928 23651
rect 960 23619 1000 23651
rect 1032 23619 1072 23651
rect 1104 23619 1144 23651
rect 1176 23619 1216 23651
rect 1248 23619 1288 23651
rect 1320 23619 1360 23651
rect 1392 23619 1432 23651
rect 1464 23619 1504 23651
rect 1536 23619 1576 23651
rect 1608 23619 1648 23651
rect 1680 23619 1720 23651
rect 1752 23619 1792 23651
rect 1824 23619 1864 23651
rect 1896 23619 1936 23651
rect 1968 23619 2008 23651
rect 2040 23619 2080 23651
rect 2112 23619 2152 23651
rect 2184 23619 2224 23651
rect 2256 23619 2296 23651
rect 2328 23619 2368 23651
rect 2400 23619 2440 23651
rect 2472 23619 2512 23651
rect 2544 23619 2584 23651
rect 2616 23619 2656 23651
rect 2688 23619 2728 23651
rect 2760 23619 2800 23651
rect 2832 23619 2872 23651
rect 2904 23619 2944 23651
rect 2976 23619 3016 23651
rect 3048 23619 3088 23651
rect 3120 23619 3160 23651
rect 3192 23619 3232 23651
rect 3264 23619 3304 23651
rect 3336 23619 3376 23651
rect 3408 23619 3448 23651
rect 3480 23619 3520 23651
rect 3552 23619 3592 23651
rect 3624 23619 3664 23651
rect 3696 23619 3736 23651
rect 3768 23619 3808 23651
rect 3840 23619 3880 23651
rect 3912 23619 3952 23651
rect 3984 23619 4024 23651
rect 4056 23619 4096 23651
rect 4128 23619 4168 23651
rect 4200 23619 4240 23651
rect 4272 23619 4312 23651
rect 4344 23619 4384 23651
rect 4416 23619 4456 23651
rect 4488 23619 4528 23651
rect 4560 23619 4600 23651
rect 4632 23619 4672 23651
rect 4704 23619 4744 23651
rect 4776 23619 4816 23651
rect 4848 23619 4888 23651
rect 4920 23619 4960 23651
rect 4992 23619 5032 23651
rect 5064 23619 5104 23651
rect 5136 23619 5176 23651
rect 5208 23619 5248 23651
rect 5280 23619 5320 23651
rect 5352 23619 5392 23651
rect 5424 23619 5464 23651
rect 5496 23619 5536 23651
rect 5568 23619 5608 23651
rect 5640 23619 5680 23651
rect 5712 23619 5752 23651
rect 5784 23619 5824 23651
rect 5856 23619 5896 23651
rect 5928 23619 5968 23651
rect 6000 23619 6040 23651
rect 6072 23619 6112 23651
rect 6144 23619 6184 23651
rect 6216 23619 6256 23651
rect 6288 23619 6328 23651
rect 6360 23619 6400 23651
rect 6432 23619 6472 23651
rect 6504 23619 6544 23651
rect 6576 23619 6616 23651
rect 6648 23619 6688 23651
rect 6720 23619 6760 23651
rect 6792 23619 6832 23651
rect 6864 23619 6904 23651
rect 6936 23619 6976 23651
rect 7008 23619 7048 23651
rect 7080 23619 7120 23651
rect 7152 23619 7192 23651
rect 7224 23619 7264 23651
rect 7296 23619 7336 23651
rect 7368 23619 7408 23651
rect 7440 23619 7480 23651
rect 7512 23619 7552 23651
rect 7584 23619 7624 23651
rect 7656 23619 7696 23651
rect 7728 23619 7768 23651
rect 7800 23619 7840 23651
rect 7872 23619 7912 23651
rect 7944 23619 7984 23651
rect 8016 23619 8056 23651
rect 8088 23619 8128 23651
rect 8160 23619 8200 23651
rect 8232 23619 8272 23651
rect 8304 23619 8344 23651
rect 8376 23619 8416 23651
rect 8448 23619 8488 23651
rect 8520 23619 8560 23651
rect 8592 23619 8632 23651
rect 8664 23619 8704 23651
rect 8736 23619 8776 23651
rect 8808 23619 8848 23651
rect 8880 23619 8920 23651
rect 8952 23619 8992 23651
rect 9024 23619 9064 23651
rect 9096 23619 9136 23651
rect 9168 23619 9208 23651
rect 9240 23619 9280 23651
rect 9312 23619 9352 23651
rect 9384 23619 9424 23651
rect 9456 23619 9496 23651
rect 9528 23619 9568 23651
rect 9600 23619 9640 23651
rect 9672 23619 9712 23651
rect 9744 23619 9784 23651
rect 9816 23619 9856 23651
rect 9888 23619 9928 23651
rect 9960 23619 10000 23651
rect 10032 23619 10072 23651
rect 10104 23619 10144 23651
rect 10176 23619 10216 23651
rect 10248 23619 10288 23651
rect 10320 23619 10360 23651
rect 10392 23619 10432 23651
rect 10464 23619 10504 23651
rect 10536 23619 10576 23651
rect 10608 23619 10648 23651
rect 10680 23619 10720 23651
rect 10752 23619 10792 23651
rect 10824 23619 10864 23651
rect 10896 23619 10936 23651
rect 10968 23619 11008 23651
rect 11040 23619 11080 23651
rect 11112 23619 11152 23651
rect 11184 23619 11224 23651
rect 11256 23619 11296 23651
rect 11328 23619 11368 23651
rect 11400 23619 11440 23651
rect 11472 23619 11512 23651
rect 11544 23619 11584 23651
rect 11616 23619 11656 23651
rect 11688 23619 11728 23651
rect 11760 23619 11800 23651
rect 11832 23619 11872 23651
rect 11904 23619 11944 23651
rect 11976 23619 12016 23651
rect 12048 23619 12088 23651
rect 12120 23619 12160 23651
rect 12192 23619 12232 23651
rect 12264 23619 12304 23651
rect 12336 23619 12376 23651
rect 12408 23619 12448 23651
rect 12480 23619 12520 23651
rect 12552 23619 12592 23651
rect 12624 23619 12664 23651
rect 12696 23619 12736 23651
rect 12768 23619 12808 23651
rect 12840 23619 12880 23651
rect 12912 23619 12952 23651
rect 12984 23619 13024 23651
rect 13056 23619 13096 23651
rect 13128 23619 13168 23651
rect 13200 23619 13240 23651
rect 13272 23619 13312 23651
rect 13344 23619 13384 23651
rect 13416 23619 13456 23651
rect 13488 23619 13528 23651
rect 13560 23619 13600 23651
rect 13632 23619 13672 23651
rect 13704 23619 13744 23651
rect 13776 23619 13816 23651
rect 13848 23619 13888 23651
rect 13920 23619 13960 23651
rect 13992 23619 14032 23651
rect 14064 23619 14104 23651
rect 14136 23619 14176 23651
rect 14208 23619 14248 23651
rect 14280 23619 14320 23651
rect 14352 23619 14392 23651
rect 14424 23619 14464 23651
rect 14496 23619 14536 23651
rect 14568 23619 14608 23651
rect 14640 23619 14680 23651
rect 14712 23619 14752 23651
rect 14784 23619 14824 23651
rect 14856 23619 14896 23651
rect 14928 23619 14968 23651
rect 15000 23619 15040 23651
rect 15072 23619 15112 23651
rect 15144 23619 15184 23651
rect 15216 23619 15256 23651
rect 15288 23619 15328 23651
rect 15360 23619 15400 23651
rect 15432 23619 15472 23651
rect 15504 23619 15544 23651
rect 15576 23619 15616 23651
rect 15648 23619 15688 23651
rect 15720 23619 15760 23651
rect 15792 23619 15832 23651
rect 15864 23619 15904 23651
rect 15936 23619 16000 23651
rect 0 23579 16000 23619
rect 0 23547 64 23579
rect 96 23547 136 23579
rect 168 23547 208 23579
rect 240 23547 280 23579
rect 312 23547 352 23579
rect 384 23547 424 23579
rect 456 23547 496 23579
rect 528 23547 568 23579
rect 600 23547 640 23579
rect 672 23547 712 23579
rect 744 23547 784 23579
rect 816 23547 856 23579
rect 888 23547 928 23579
rect 960 23547 1000 23579
rect 1032 23547 1072 23579
rect 1104 23547 1144 23579
rect 1176 23547 1216 23579
rect 1248 23547 1288 23579
rect 1320 23547 1360 23579
rect 1392 23547 1432 23579
rect 1464 23547 1504 23579
rect 1536 23547 1576 23579
rect 1608 23547 1648 23579
rect 1680 23547 1720 23579
rect 1752 23547 1792 23579
rect 1824 23547 1864 23579
rect 1896 23547 1936 23579
rect 1968 23547 2008 23579
rect 2040 23547 2080 23579
rect 2112 23547 2152 23579
rect 2184 23547 2224 23579
rect 2256 23547 2296 23579
rect 2328 23547 2368 23579
rect 2400 23547 2440 23579
rect 2472 23547 2512 23579
rect 2544 23547 2584 23579
rect 2616 23547 2656 23579
rect 2688 23547 2728 23579
rect 2760 23547 2800 23579
rect 2832 23547 2872 23579
rect 2904 23547 2944 23579
rect 2976 23547 3016 23579
rect 3048 23547 3088 23579
rect 3120 23547 3160 23579
rect 3192 23547 3232 23579
rect 3264 23547 3304 23579
rect 3336 23547 3376 23579
rect 3408 23547 3448 23579
rect 3480 23547 3520 23579
rect 3552 23547 3592 23579
rect 3624 23547 3664 23579
rect 3696 23547 3736 23579
rect 3768 23547 3808 23579
rect 3840 23547 3880 23579
rect 3912 23547 3952 23579
rect 3984 23547 4024 23579
rect 4056 23547 4096 23579
rect 4128 23547 4168 23579
rect 4200 23547 4240 23579
rect 4272 23547 4312 23579
rect 4344 23547 4384 23579
rect 4416 23547 4456 23579
rect 4488 23547 4528 23579
rect 4560 23547 4600 23579
rect 4632 23547 4672 23579
rect 4704 23547 4744 23579
rect 4776 23547 4816 23579
rect 4848 23547 4888 23579
rect 4920 23547 4960 23579
rect 4992 23547 5032 23579
rect 5064 23547 5104 23579
rect 5136 23547 5176 23579
rect 5208 23547 5248 23579
rect 5280 23547 5320 23579
rect 5352 23547 5392 23579
rect 5424 23547 5464 23579
rect 5496 23547 5536 23579
rect 5568 23547 5608 23579
rect 5640 23547 5680 23579
rect 5712 23547 5752 23579
rect 5784 23547 5824 23579
rect 5856 23547 5896 23579
rect 5928 23547 5968 23579
rect 6000 23547 6040 23579
rect 6072 23547 6112 23579
rect 6144 23547 6184 23579
rect 6216 23547 6256 23579
rect 6288 23547 6328 23579
rect 6360 23547 6400 23579
rect 6432 23547 6472 23579
rect 6504 23547 6544 23579
rect 6576 23547 6616 23579
rect 6648 23547 6688 23579
rect 6720 23547 6760 23579
rect 6792 23547 6832 23579
rect 6864 23547 6904 23579
rect 6936 23547 6976 23579
rect 7008 23547 7048 23579
rect 7080 23547 7120 23579
rect 7152 23547 7192 23579
rect 7224 23547 7264 23579
rect 7296 23547 7336 23579
rect 7368 23547 7408 23579
rect 7440 23547 7480 23579
rect 7512 23547 7552 23579
rect 7584 23547 7624 23579
rect 7656 23547 7696 23579
rect 7728 23547 7768 23579
rect 7800 23547 7840 23579
rect 7872 23547 7912 23579
rect 7944 23547 7984 23579
rect 8016 23547 8056 23579
rect 8088 23547 8128 23579
rect 8160 23547 8200 23579
rect 8232 23547 8272 23579
rect 8304 23547 8344 23579
rect 8376 23547 8416 23579
rect 8448 23547 8488 23579
rect 8520 23547 8560 23579
rect 8592 23547 8632 23579
rect 8664 23547 8704 23579
rect 8736 23547 8776 23579
rect 8808 23547 8848 23579
rect 8880 23547 8920 23579
rect 8952 23547 8992 23579
rect 9024 23547 9064 23579
rect 9096 23547 9136 23579
rect 9168 23547 9208 23579
rect 9240 23547 9280 23579
rect 9312 23547 9352 23579
rect 9384 23547 9424 23579
rect 9456 23547 9496 23579
rect 9528 23547 9568 23579
rect 9600 23547 9640 23579
rect 9672 23547 9712 23579
rect 9744 23547 9784 23579
rect 9816 23547 9856 23579
rect 9888 23547 9928 23579
rect 9960 23547 10000 23579
rect 10032 23547 10072 23579
rect 10104 23547 10144 23579
rect 10176 23547 10216 23579
rect 10248 23547 10288 23579
rect 10320 23547 10360 23579
rect 10392 23547 10432 23579
rect 10464 23547 10504 23579
rect 10536 23547 10576 23579
rect 10608 23547 10648 23579
rect 10680 23547 10720 23579
rect 10752 23547 10792 23579
rect 10824 23547 10864 23579
rect 10896 23547 10936 23579
rect 10968 23547 11008 23579
rect 11040 23547 11080 23579
rect 11112 23547 11152 23579
rect 11184 23547 11224 23579
rect 11256 23547 11296 23579
rect 11328 23547 11368 23579
rect 11400 23547 11440 23579
rect 11472 23547 11512 23579
rect 11544 23547 11584 23579
rect 11616 23547 11656 23579
rect 11688 23547 11728 23579
rect 11760 23547 11800 23579
rect 11832 23547 11872 23579
rect 11904 23547 11944 23579
rect 11976 23547 12016 23579
rect 12048 23547 12088 23579
rect 12120 23547 12160 23579
rect 12192 23547 12232 23579
rect 12264 23547 12304 23579
rect 12336 23547 12376 23579
rect 12408 23547 12448 23579
rect 12480 23547 12520 23579
rect 12552 23547 12592 23579
rect 12624 23547 12664 23579
rect 12696 23547 12736 23579
rect 12768 23547 12808 23579
rect 12840 23547 12880 23579
rect 12912 23547 12952 23579
rect 12984 23547 13024 23579
rect 13056 23547 13096 23579
rect 13128 23547 13168 23579
rect 13200 23547 13240 23579
rect 13272 23547 13312 23579
rect 13344 23547 13384 23579
rect 13416 23547 13456 23579
rect 13488 23547 13528 23579
rect 13560 23547 13600 23579
rect 13632 23547 13672 23579
rect 13704 23547 13744 23579
rect 13776 23547 13816 23579
rect 13848 23547 13888 23579
rect 13920 23547 13960 23579
rect 13992 23547 14032 23579
rect 14064 23547 14104 23579
rect 14136 23547 14176 23579
rect 14208 23547 14248 23579
rect 14280 23547 14320 23579
rect 14352 23547 14392 23579
rect 14424 23547 14464 23579
rect 14496 23547 14536 23579
rect 14568 23547 14608 23579
rect 14640 23547 14680 23579
rect 14712 23547 14752 23579
rect 14784 23547 14824 23579
rect 14856 23547 14896 23579
rect 14928 23547 14968 23579
rect 15000 23547 15040 23579
rect 15072 23547 15112 23579
rect 15144 23547 15184 23579
rect 15216 23547 15256 23579
rect 15288 23547 15328 23579
rect 15360 23547 15400 23579
rect 15432 23547 15472 23579
rect 15504 23547 15544 23579
rect 15576 23547 15616 23579
rect 15648 23547 15688 23579
rect 15720 23547 15760 23579
rect 15792 23547 15832 23579
rect 15864 23547 15904 23579
rect 15936 23547 16000 23579
rect 0 23507 16000 23547
rect 0 23475 64 23507
rect 96 23475 136 23507
rect 168 23475 208 23507
rect 240 23475 280 23507
rect 312 23475 352 23507
rect 384 23475 424 23507
rect 456 23475 496 23507
rect 528 23475 568 23507
rect 600 23475 640 23507
rect 672 23475 712 23507
rect 744 23475 784 23507
rect 816 23475 856 23507
rect 888 23475 928 23507
rect 960 23475 1000 23507
rect 1032 23475 1072 23507
rect 1104 23475 1144 23507
rect 1176 23475 1216 23507
rect 1248 23475 1288 23507
rect 1320 23475 1360 23507
rect 1392 23475 1432 23507
rect 1464 23475 1504 23507
rect 1536 23475 1576 23507
rect 1608 23475 1648 23507
rect 1680 23475 1720 23507
rect 1752 23475 1792 23507
rect 1824 23475 1864 23507
rect 1896 23475 1936 23507
rect 1968 23475 2008 23507
rect 2040 23475 2080 23507
rect 2112 23475 2152 23507
rect 2184 23475 2224 23507
rect 2256 23475 2296 23507
rect 2328 23475 2368 23507
rect 2400 23475 2440 23507
rect 2472 23475 2512 23507
rect 2544 23475 2584 23507
rect 2616 23475 2656 23507
rect 2688 23475 2728 23507
rect 2760 23475 2800 23507
rect 2832 23475 2872 23507
rect 2904 23475 2944 23507
rect 2976 23475 3016 23507
rect 3048 23475 3088 23507
rect 3120 23475 3160 23507
rect 3192 23475 3232 23507
rect 3264 23475 3304 23507
rect 3336 23475 3376 23507
rect 3408 23475 3448 23507
rect 3480 23475 3520 23507
rect 3552 23475 3592 23507
rect 3624 23475 3664 23507
rect 3696 23475 3736 23507
rect 3768 23475 3808 23507
rect 3840 23475 3880 23507
rect 3912 23475 3952 23507
rect 3984 23475 4024 23507
rect 4056 23475 4096 23507
rect 4128 23475 4168 23507
rect 4200 23475 4240 23507
rect 4272 23475 4312 23507
rect 4344 23475 4384 23507
rect 4416 23475 4456 23507
rect 4488 23475 4528 23507
rect 4560 23475 4600 23507
rect 4632 23475 4672 23507
rect 4704 23475 4744 23507
rect 4776 23475 4816 23507
rect 4848 23475 4888 23507
rect 4920 23475 4960 23507
rect 4992 23475 5032 23507
rect 5064 23475 5104 23507
rect 5136 23475 5176 23507
rect 5208 23475 5248 23507
rect 5280 23475 5320 23507
rect 5352 23475 5392 23507
rect 5424 23475 5464 23507
rect 5496 23475 5536 23507
rect 5568 23475 5608 23507
rect 5640 23475 5680 23507
rect 5712 23475 5752 23507
rect 5784 23475 5824 23507
rect 5856 23475 5896 23507
rect 5928 23475 5968 23507
rect 6000 23475 6040 23507
rect 6072 23475 6112 23507
rect 6144 23475 6184 23507
rect 6216 23475 6256 23507
rect 6288 23475 6328 23507
rect 6360 23475 6400 23507
rect 6432 23475 6472 23507
rect 6504 23475 6544 23507
rect 6576 23475 6616 23507
rect 6648 23475 6688 23507
rect 6720 23475 6760 23507
rect 6792 23475 6832 23507
rect 6864 23475 6904 23507
rect 6936 23475 6976 23507
rect 7008 23475 7048 23507
rect 7080 23475 7120 23507
rect 7152 23475 7192 23507
rect 7224 23475 7264 23507
rect 7296 23475 7336 23507
rect 7368 23475 7408 23507
rect 7440 23475 7480 23507
rect 7512 23475 7552 23507
rect 7584 23475 7624 23507
rect 7656 23475 7696 23507
rect 7728 23475 7768 23507
rect 7800 23475 7840 23507
rect 7872 23475 7912 23507
rect 7944 23475 7984 23507
rect 8016 23475 8056 23507
rect 8088 23475 8128 23507
rect 8160 23475 8200 23507
rect 8232 23475 8272 23507
rect 8304 23475 8344 23507
rect 8376 23475 8416 23507
rect 8448 23475 8488 23507
rect 8520 23475 8560 23507
rect 8592 23475 8632 23507
rect 8664 23475 8704 23507
rect 8736 23475 8776 23507
rect 8808 23475 8848 23507
rect 8880 23475 8920 23507
rect 8952 23475 8992 23507
rect 9024 23475 9064 23507
rect 9096 23475 9136 23507
rect 9168 23475 9208 23507
rect 9240 23475 9280 23507
rect 9312 23475 9352 23507
rect 9384 23475 9424 23507
rect 9456 23475 9496 23507
rect 9528 23475 9568 23507
rect 9600 23475 9640 23507
rect 9672 23475 9712 23507
rect 9744 23475 9784 23507
rect 9816 23475 9856 23507
rect 9888 23475 9928 23507
rect 9960 23475 10000 23507
rect 10032 23475 10072 23507
rect 10104 23475 10144 23507
rect 10176 23475 10216 23507
rect 10248 23475 10288 23507
rect 10320 23475 10360 23507
rect 10392 23475 10432 23507
rect 10464 23475 10504 23507
rect 10536 23475 10576 23507
rect 10608 23475 10648 23507
rect 10680 23475 10720 23507
rect 10752 23475 10792 23507
rect 10824 23475 10864 23507
rect 10896 23475 10936 23507
rect 10968 23475 11008 23507
rect 11040 23475 11080 23507
rect 11112 23475 11152 23507
rect 11184 23475 11224 23507
rect 11256 23475 11296 23507
rect 11328 23475 11368 23507
rect 11400 23475 11440 23507
rect 11472 23475 11512 23507
rect 11544 23475 11584 23507
rect 11616 23475 11656 23507
rect 11688 23475 11728 23507
rect 11760 23475 11800 23507
rect 11832 23475 11872 23507
rect 11904 23475 11944 23507
rect 11976 23475 12016 23507
rect 12048 23475 12088 23507
rect 12120 23475 12160 23507
rect 12192 23475 12232 23507
rect 12264 23475 12304 23507
rect 12336 23475 12376 23507
rect 12408 23475 12448 23507
rect 12480 23475 12520 23507
rect 12552 23475 12592 23507
rect 12624 23475 12664 23507
rect 12696 23475 12736 23507
rect 12768 23475 12808 23507
rect 12840 23475 12880 23507
rect 12912 23475 12952 23507
rect 12984 23475 13024 23507
rect 13056 23475 13096 23507
rect 13128 23475 13168 23507
rect 13200 23475 13240 23507
rect 13272 23475 13312 23507
rect 13344 23475 13384 23507
rect 13416 23475 13456 23507
rect 13488 23475 13528 23507
rect 13560 23475 13600 23507
rect 13632 23475 13672 23507
rect 13704 23475 13744 23507
rect 13776 23475 13816 23507
rect 13848 23475 13888 23507
rect 13920 23475 13960 23507
rect 13992 23475 14032 23507
rect 14064 23475 14104 23507
rect 14136 23475 14176 23507
rect 14208 23475 14248 23507
rect 14280 23475 14320 23507
rect 14352 23475 14392 23507
rect 14424 23475 14464 23507
rect 14496 23475 14536 23507
rect 14568 23475 14608 23507
rect 14640 23475 14680 23507
rect 14712 23475 14752 23507
rect 14784 23475 14824 23507
rect 14856 23475 14896 23507
rect 14928 23475 14968 23507
rect 15000 23475 15040 23507
rect 15072 23475 15112 23507
rect 15144 23475 15184 23507
rect 15216 23475 15256 23507
rect 15288 23475 15328 23507
rect 15360 23475 15400 23507
rect 15432 23475 15472 23507
rect 15504 23475 15544 23507
rect 15576 23475 15616 23507
rect 15648 23475 15688 23507
rect 15720 23475 15760 23507
rect 15792 23475 15832 23507
rect 15864 23475 15904 23507
rect 15936 23475 16000 23507
rect 0 23435 16000 23475
rect 0 23403 64 23435
rect 96 23403 136 23435
rect 168 23403 208 23435
rect 240 23403 280 23435
rect 312 23403 352 23435
rect 384 23403 424 23435
rect 456 23403 496 23435
rect 528 23403 568 23435
rect 600 23403 640 23435
rect 672 23403 712 23435
rect 744 23403 784 23435
rect 816 23403 856 23435
rect 888 23403 928 23435
rect 960 23403 1000 23435
rect 1032 23403 1072 23435
rect 1104 23403 1144 23435
rect 1176 23403 1216 23435
rect 1248 23403 1288 23435
rect 1320 23403 1360 23435
rect 1392 23403 1432 23435
rect 1464 23403 1504 23435
rect 1536 23403 1576 23435
rect 1608 23403 1648 23435
rect 1680 23403 1720 23435
rect 1752 23403 1792 23435
rect 1824 23403 1864 23435
rect 1896 23403 1936 23435
rect 1968 23403 2008 23435
rect 2040 23403 2080 23435
rect 2112 23403 2152 23435
rect 2184 23403 2224 23435
rect 2256 23403 2296 23435
rect 2328 23403 2368 23435
rect 2400 23403 2440 23435
rect 2472 23403 2512 23435
rect 2544 23403 2584 23435
rect 2616 23403 2656 23435
rect 2688 23403 2728 23435
rect 2760 23403 2800 23435
rect 2832 23403 2872 23435
rect 2904 23403 2944 23435
rect 2976 23403 3016 23435
rect 3048 23403 3088 23435
rect 3120 23403 3160 23435
rect 3192 23403 3232 23435
rect 3264 23403 3304 23435
rect 3336 23403 3376 23435
rect 3408 23403 3448 23435
rect 3480 23403 3520 23435
rect 3552 23403 3592 23435
rect 3624 23403 3664 23435
rect 3696 23403 3736 23435
rect 3768 23403 3808 23435
rect 3840 23403 3880 23435
rect 3912 23403 3952 23435
rect 3984 23403 4024 23435
rect 4056 23403 4096 23435
rect 4128 23403 4168 23435
rect 4200 23403 4240 23435
rect 4272 23403 4312 23435
rect 4344 23403 4384 23435
rect 4416 23403 4456 23435
rect 4488 23403 4528 23435
rect 4560 23403 4600 23435
rect 4632 23403 4672 23435
rect 4704 23403 4744 23435
rect 4776 23403 4816 23435
rect 4848 23403 4888 23435
rect 4920 23403 4960 23435
rect 4992 23403 5032 23435
rect 5064 23403 5104 23435
rect 5136 23403 5176 23435
rect 5208 23403 5248 23435
rect 5280 23403 5320 23435
rect 5352 23403 5392 23435
rect 5424 23403 5464 23435
rect 5496 23403 5536 23435
rect 5568 23403 5608 23435
rect 5640 23403 5680 23435
rect 5712 23403 5752 23435
rect 5784 23403 5824 23435
rect 5856 23403 5896 23435
rect 5928 23403 5968 23435
rect 6000 23403 6040 23435
rect 6072 23403 6112 23435
rect 6144 23403 6184 23435
rect 6216 23403 6256 23435
rect 6288 23403 6328 23435
rect 6360 23403 6400 23435
rect 6432 23403 6472 23435
rect 6504 23403 6544 23435
rect 6576 23403 6616 23435
rect 6648 23403 6688 23435
rect 6720 23403 6760 23435
rect 6792 23403 6832 23435
rect 6864 23403 6904 23435
rect 6936 23403 6976 23435
rect 7008 23403 7048 23435
rect 7080 23403 7120 23435
rect 7152 23403 7192 23435
rect 7224 23403 7264 23435
rect 7296 23403 7336 23435
rect 7368 23403 7408 23435
rect 7440 23403 7480 23435
rect 7512 23403 7552 23435
rect 7584 23403 7624 23435
rect 7656 23403 7696 23435
rect 7728 23403 7768 23435
rect 7800 23403 7840 23435
rect 7872 23403 7912 23435
rect 7944 23403 7984 23435
rect 8016 23403 8056 23435
rect 8088 23403 8128 23435
rect 8160 23403 8200 23435
rect 8232 23403 8272 23435
rect 8304 23403 8344 23435
rect 8376 23403 8416 23435
rect 8448 23403 8488 23435
rect 8520 23403 8560 23435
rect 8592 23403 8632 23435
rect 8664 23403 8704 23435
rect 8736 23403 8776 23435
rect 8808 23403 8848 23435
rect 8880 23403 8920 23435
rect 8952 23403 8992 23435
rect 9024 23403 9064 23435
rect 9096 23403 9136 23435
rect 9168 23403 9208 23435
rect 9240 23403 9280 23435
rect 9312 23403 9352 23435
rect 9384 23403 9424 23435
rect 9456 23403 9496 23435
rect 9528 23403 9568 23435
rect 9600 23403 9640 23435
rect 9672 23403 9712 23435
rect 9744 23403 9784 23435
rect 9816 23403 9856 23435
rect 9888 23403 9928 23435
rect 9960 23403 10000 23435
rect 10032 23403 10072 23435
rect 10104 23403 10144 23435
rect 10176 23403 10216 23435
rect 10248 23403 10288 23435
rect 10320 23403 10360 23435
rect 10392 23403 10432 23435
rect 10464 23403 10504 23435
rect 10536 23403 10576 23435
rect 10608 23403 10648 23435
rect 10680 23403 10720 23435
rect 10752 23403 10792 23435
rect 10824 23403 10864 23435
rect 10896 23403 10936 23435
rect 10968 23403 11008 23435
rect 11040 23403 11080 23435
rect 11112 23403 11152 23435
rect 11184 23403 11224 23435
rect 11256 23403 11296 23435
rect 11328 23403 11368 23435
rect 11400 23403 11440 23435
rect 11472 23403 11512 23435
rect 11544 23403 11584 23435
rect 11616 23403 11656 23435
rect 11688 23403 11728 23435
rect 11760 23403 11800 23435
rect 11832 23403 11872 23435
rect 11904 23403 11944 23435
rect 11976 23403 12016 23435
rect 12048 23403 12088 23435
rect 12120 23403 12160 23435
rect 12192 23403 12232 23435
rect 12264 23403 12304 23435
rect 12336 23403 12376 23435
rect 12408 23403 12448 23435
rect 12480 23403 12520 23435
rect 12552 23403 12592 23435
rect 12624 23403 12664 23435
rect 12696 23403 12736 23435
rect 12768 23403 12808 23435
rect 12840 23403 12880 23435
rect 12912 23403 12952 23435
rect 12984 23403 13024 23435
rect 13056 23403 13096 23435
rect 13128 23403 13168 23435
rect 13200 23403 13240 23435
rect 13272 23403 13312 23435
rect 13344 23403 13384 23435
rect 13416 23403 13456 23435
rect 13488 23403 13528 23435
rect 13560 23403 13600 23435
rect 13632 23403 13672 23435
rect 13704 23403 13744 23435
rect 13776 23403 13816 23435
rect 13848 23403 13888 23435
rect 13920 23403 13960 23435
rect 13992 23403 14032 23435
rect 14064 23403 14104 23435
rect 14136 23403 14176 23435
rect 14208 23403 14248 23435
rect 14280 23403 14320 23435
rect 14352 23403 14392 23435
rect 14424 23403 14464 23435
rect 14496 23403 14536 23435
rect 14568 23403 14608 23435
rect 14640 23403 14680 23435
rect 14712 23403 14752 23435
rect 14784 23403 14824 23435
rect 14856 23403 14896 23435
rect 14928 23403 14968 23435
rect 15000 23403 15040 23435
rect 15072 23403 15112 23435
rect 15144 23403 15184 23435
rect 15216 23403 15256 23435
rect 15288 23403 15328 23435
rect 15360 23403 15400 23435
rect 15432 23403 15472 23435
rect 15504 23403 15544 23435
rect 15576 23403 15616 23435
rect 15648 23403 15688 23435
rect 15720 23403 15760 23435
rect 15792 23403 15832 23435
rect 15864 23403 15904 23435
rect 15936 23403 16000 23435
rect 0 23363 16000 23403
rect 0 23331 64 23363
rect 96 23331 136 23363
rect 168 23331 208 23363
rect 240 23331 280 23363
rect 312 23331 352 23363
rect 384 23331 424 23363
rect 456 23331 496 23363
rect 528 23331 568 23363
rect 600 23331 640 23363
rect 672 23331 712 23363
rect 744 23331 784 23363
rect 816 23331 856 23363
rect 888 23331 928 23363
rect 960 23331 1000 23363
rect 1032 23331 1072 23363
rect 1104 23331 1144 23363
rect 1176 23331 1216 23363
rect 1248 23331 1288 23363
rect 1320 23331 1360 23363
rect 1392 23331 1432 23363
rect 1464 23331 1504 23363
rect 1536 23331 1576 23363
rect 1608 23331 1648 23363
rect 1680 23331 1720 23363
rect 1752 23331 1792 23363
rect 1824 23331 1864 23363
rect 1896 23331 1936 23363
rect 1968 23331 2008 23363
rect 2040 23331 2080 23363
rect 2112 23331 2152 23363
rect 2184 23331 2224 23363
rect 2256 23331 2296 23363
rect 2328 23331 2368 23363
rect 2400 23331 2440 23363
rect 2472 23331 2512 23363
rect 2544 23331 2584 23363
rect 2616 23331 2656 23363
rect 2688 23331 2728 23363
rect 2760 23331 2800 23363
rect 2832 23331 2872 23363
rect 2904 23331 2944 23363
rect 2976 23331 3016 23363
rect 3048 23331 3088 23363
rect 3120 23331 3160 23363
rect 3192 23331 3232 23363
rect 3264 23331 3304 23363
rect 3336 23331 3376 23363
rect 3408 23331 3448 23363
rect 3480 23331 3520 23363
rect 3552 23331 3592 23363
rect 3624 23331 3664 23363
rect 3696 23331 3736 23363
rect 3768 23331 3808 23363
rect 3840 23331 3880 23363
rect 3912 23331 3952 23363
rect 3984 23331 4024 23363
rect 4056 23331 4096 23363
rect 4128 23331 4168 23363
rect 4200 23331 4240 23363
rect 4272 23331 4312 23363
rect 4344 23331 4384 23363
rect 4416 23331 4456 23363
rect 4488 23331 4528 23363
rect 4560 23331 4600 23363
rect 4632 23331 4672 23363
rect 4704 23331 4744 23363
rect 4776 23331 4816 23363
rect 4848 23331 4888 23363
rect 4920 23331 4960 23363
rect 4992 23331 5032 23363
rect 5064 23331 5104 23363
rect 5136 23331 5176 23363
rect 5208 23331 5248 23363
rect 5280 23331 5320 23363
rect 5352 23331 5392 23363
rect 5424 23331 5464 23363
rect 5496 23331 5536 23363
rect 5568 23331 5608 23363
rect 5640 23331 5680 23363
rect 5712 23331 5752 23363
rect 5784 23331 5824 23363
rect 5856 23331 5896 23363
rect 5928 23331 5968 23363
rect 6000 23331 6040 23363
rect 6072 23331 6112 23363
rect 6144 23331 6184 23363
rect 6216 23331 6256 23363
rect 6288 23331 6328 23363
rect 6360 23331 6400 23363
rect 6432 23331 6472 23363
rect 6504 23331 6544 23363
rect 6576 23331 6616 23363
rect 6648 23331 6688 23363
rect 6720 23331 6760 23363
rect 6792 23331 6832 23363
rect 6864 23331 6904 23363
rect 6936 23331 6976 23363
rect 7008 23331 7048 23363
rect 7080 23331 7120 23363
rect 7152 23331 7192 23363
rect 7224 23331 7264 23363
rect 7296 23331 7336 23363
rect 7368 23331 7408 23363
rect 7440 23331 7480 23363
rect 7512 23331 7552 23363
rect 7584 23331 7624 23363
rect 7656 23331 7696 23363
rect 7728 23331 7768 23363
rect 7800 23331 7840 23363
rect 7872 23331 7912 23363
rect 7944 23331 7984 23363
rect 8016 23331 8056 23363
rect 8088 23331 8128 23363
rect 8160 23331 8200 23363
rect 8232 23331 8272 23363
rect 8304 23331 8344 23363
rect 8376 23331 8416 23363
rect 8448 23331 8488 23363
rect 8520 23331 8560 23363
rect 8592 23331 8632 23363
rect 8664 23331 8704 23363
rect 8736 23331 8776 23363
rect 8808 23331 8848 23363
rect 8880 23331 8920 23363
rect 8952 23331 8992 23363
rect 9024 23331 9064 23363
rect 9096 23331 9136 23363
rect 9168 23331 9208 23363
rect 9240 23331 9280 23363
rect 9312 23331 9352 23363
rect 9384 23331 9424 23363
rect 9456 23331 9496 23363
rect 9528 23331 9568 23363
rect 9600 23331 9640 23363
rect 9672 23331 9712 23363
rect 9744 23331 9784 23363
rect 9816 23331 9856 23363
rect 9888 23331 9928 23363
rect 9960 23331 10000 23363
rect 10032 23331 10072 23363
rect 10104 23331 10144 23363
rect 10176 23331 10216 23363
rect 10248 23331 10288 23363
rect 10320 23331 10360 23363
rect 10392 23331 10432 23363
rect 10464 23331 10504 23363
rect 10536 23331 10576 23363
rect 10608 23331 10648 23363
rect 10680 23331 10720 23363
rect 10752 23331 10792 23363
rect 10824 23331 10864 23363
rect 10896 23331 10936 23363
rect 10968 23331 11008 23363
rect 11040 23331 11080 23363
rect 11112 23331 11152 23363
rect 11184 23331 11224 23363
rect 11256 23331 11296 23363
rect 11328 23331 11368 23363
rect 11400 23331 11440 23363
rect 11472 23331 11512 23363
rect 11544 23331 11584 23363
rect 11616 23331 11656 23363
rect 11688 23331 11728 23363
rect 11760 23331 11800 23363
rect 11832 23331 11872 23363
rect 11904 23331 11944 23363
rect 11976 23331 12016 23363
rect 12048 23331 12088 23363
rect 12120 23331 12160 23363
rect 12192 23331 12232 23363
rect 12264 23331 12304 23363
rect 12336 23331 12376 23363
rect 12408 23331 12448 23363
rect 12480 23331 12520 23363
rect 12552 23331 12592 23363
rect 12624 23331 12664 23363
rect 12696 23331 12736 23363
rect 12768 23331 12808 23363
rect 12840 23331 12880 23363
rect 12912 23331 12952 23363
rect 12984 23331 13024 23363
rect 13056 23331 13096 23363
rect 13128 23331 13168 23363
rect 13200 23331 13240 23363
rect 13272 23331 13312 23363
rect 13344 23331 13384 23363
rect 13416 23331 13456 23363
rect 13488 23331 13528 23363
rect 13560 23331 13600 23363
rect 13632 23331 13672 23363
rect 13704 23331 13744 23363
rect 13776 23331 13816 23363
rect 13848 23331 13888 23363
rect 13920 23331 13960 23363
rect 13992 23331 14032 23363
rect 14064 23331 14104 23363
rect 14136 23331 14176 23363
rect 14208 23331 14248 23363
rect 14280 23331 14320 23363
rect 14352 23331 14392 23363
rect 14424 23331 14464 23363
rect 14496 23331 14536 23363
rect 14568 23331 14608 23363
rect 14640 23331 14680 23363
rect 14712 23331 14752 23363
rect 14784 23331 14824 23363
rect 14856 23331 14896 23363
rect 14928 23331 14968 23363
rect 15000 23331 15040 23363
rect 15072 23331 15112 23363
rect 15144 23331 15184 23363
rect 15216 23331 15256 23363
rect 15288 23331 15328 23363
rect 15360 23331 15400 23363
rect 15432 23331 15472 23363
rect 15504 23331 15544 23363
rect 15576 23331 15616 23363
rect 15648 23331 15688 23363
rect 15720 23331 15760 23363
rect 15792 23331 15832 23363
rect 15864 23331 15904 23363
rect 15936 23331 16000 23363
rect 0 23291 16000 23331
rect 0 23259 64 23291
rect 96 23259 136 23291
rect 168 23259 208 23291
rect 240 23259 280 23291
rect 312 23259 352 23291
rect 384 23259 424 23291
rect 456 23259 496 23291
rect 528 23259 568 23291
rect 600 23259 640 23291
rect 672 23259 712 23291
rect 744 23259 784 23291
rect 816 23259 856 23291
rect 888 23259 928 23291
rect 960 23259 1000 23291
rect 1032 23259 1072 23291
rect 1104 23259 1144 23291
rect 1176 23259 1216 23291
rect 1248 23259 1288 23291
rect 1320 23259 1360 23291
rect 1392 23259 1432 23291
rect 1464 23259 1504 23291
rect 1536 23259 1576 23291
rect 1608 23259 1648 23291
rect 1680 23259 1720 23291
rect 1752 23259 1792 23291
rect 1824 23259 1864 23291
rect 1896 23259 1936 23291
rect 1968 23259 2008 23291
rect 2040 23259 2080 23291
rect 2112 23259 2152 23291
rect 2184 23259 2224 23291
rect 2256 23259 2296 23291
rect 2328 23259 2368 23291
rect 2400 23259 2440 23291
rect 2472 23259 2512 23291
rect 2544 23259 2584 23291
rect 2616 23259 2656 23291
rect 2688 23259 2728 23291
rect 2760 23259 2800 23291
rect 2832 23259 2872 23291
rect 2904 23259 2944 23291
rect 2976 23259 3016 23291
rect 3048 23259 3088 23291
rect 3120 23259 3160 23291
rect 3192 23259 3232 23291
rect 3264 23259 3304 23291
rect 3336 23259 3376 23291
rect 3408 23259 3448 23291
rect 3480 23259 3520 23291
rect 3552 23259 3592 23291
rect 3624 23259 3664 23291
rect 3696 23259 3736 23291
rect 3768 23259 3808 23291
rect 3840 23259 3880 23291
rect 3912 23259 3952 23291
rect 3984 23259 4024 23291
rect 4056 23259 4096 23291
rect 4128 23259 4168 23291
rect 4200 23259 4240 23291
rect 4272 23259 4312 23291
rect 4344 23259 4384 23291
rect 4416 23259 4456 23291
rect 4488 23259 4528 23291
rect 4560 23259 4600 23291
rect 4632 23259 4672 23291
rect 4704 23259 4744 23291
rect 4776 23259 4816 23291
rect 4848 23259 4888 23291
rect 4920 23259 4960 23291
rect 4992 23259 5032 23291
rect 5064 23259 5104 23291
rect 5136 23259 5176 23291
rect 5208 23259 5248 23291
rect 5280 23259 5320 23291
rect 5352 23259 5392 23291
rect 5424 23259 5464 23291
rect 5496 23259 5536 23291
rect 5568 23259 5608 23291
rect 5640 23259 5680 23291
rect 5712 23259 5752 23291
rect 5784 23259 5824 23291
rect 5856 23259 5896 23291
rect 5928 23259 5968 23291
rect 6000 23259 6040 23291
rect 6072 23259 6112 23291
rect 6144 23259 6184 23291
rect 6216 23259 6256 23291
rect 6288 23259 6328 23291
rect 6360 23259 6400 23291
rect 6432 23259 6472 23291
rect 6504 23259 6544 23291
rect 6576 23259 6616 23291
rect 6648 23259 6688 23291
rect 6720 23259 6760 23291
rect 6792 23259 6832 23291
rect 6864 23259 6904 23291
rect 6936 23259 6976 23291
rect 7008 23259 7048 23291
rect 7080 23259 7120 23291
rect 7152 23259 7192 23291
rect 7224 23259 7264 23291
rect 7296 23259 7336 23291
rect 7368 23259 7408 23291
rect 7440 23259 7480 23291
rect 7512 23259 7552 23291
rect 7584 23259 7624 23291
rect 7656 23259 7696 23291
rect 7728 23259 7768 23291
rect 7800 23259 7840 23291
rect 7872 23259 7912 23291
rect 7944 23259 7984 23291
rect 8016 23259 8056 23291
rect 8088 23259 8128 23291
rect 8160 23259 8200 23291
rect 8232 23259 8272 23291
rect 8304 23259 8344 23291
rect 8376 23259 8416 23291
rect 8448 23259 8488 23291
rect 8520 23259 8560 23291
rect 8592 23259 8632 23291
rect 8664 23259 8704 23291
rect 8736 23259 8776 23291
rect 8808 23259 8848 23291
rect 8880 23259 8920 23291
rect 8952 23259 8992 23291
rect 9024 23259 9064 23291
rect 9096 23259 9136 23291
rect 9168 23259 9208 23291
rect 9240 23259 9280 23291
rect 9312 23259 9352 23291
rect 9384 23259 9424 23291
rect 9456 23259 9496 23291
rect 9528 23259 9568 23291
rect 9600 23259 9640 23291
rect 9672 23259 9712 23291
rect 9744 23259 9784 23291
rect 9816 23259 9856 23291
rect 9888 23259 9928 23291
rect 9960 23259 10000 23291
rect 10032 23259 10072 23291
rect 10104 23259 10144 23291
rect 10176 23259 10216 23291
rect 10248 23259 10288 23291
rect 10320 23259 10360 23291
rect 10392 23259 10432 23291
rect 10464 23259 10504 23291
rect 10536 23259 10576 23291
rect 10608 23259 10648 23291
rect 10680 23259 10720 23291
rect 10752 23259 10792 23291
rect 10824 23259 10864 23291
rect 10896 23259 10936 23291
rect 10968 23259 11008 23291
rect 11040 23259 11080 23291
rect 11112 23259 11152 23291
rect 11184 23259 11224 23291
rect 11256 23259 11296 23291
rect 11328 23259 11368 23291
rect 11400 23259 11440 23291
rect 11472 23259 11512 23291
rect 11544 23259 11584 23291
rect 11616 23259 11656 23291
rect 11688 23259 11728 23291
rect 11760 23259 11800 23291
rect 11832 23259 11872 23291
rect 11904 23259 11944 23291
rect 11976 23259 12016 23291
rect 12048 23259 12088 23291
rect 12120 23259 12160 23291
rect 12192 23259 12232 23291
rect 12264 23259 12304 23291
rect 12336 23259 12376 23291
rect 12408 23259 12448 23291
rect 12480 23259 12520 23291
rect 12552 23259 12592 23291
rect 12624 23259 12664 23291
rect 12696 23259 12736 23291
rect 12768 23259 12808 23291
rect 12840 23259 12880 23291
rect 12912 23259 12952 23291
rect 12984 23259 13024 23291
rect 13056 23259 13096 23291
rect 13128 23259 13168 23291
rect 13200 23259 13240 23291
rect 13272 23259 13312 23291
rect 13344 23259 13384 23291
rect 13416 23259 13456 23291
rect 13488 23259 13528 23291
rect 13560 23259 13600 23291
rect 13632 23259 13672 23291
rect 13704 23259 13744 23291
rect 13776 23259 13816 23291
rect 13848 23259 13888 23291
rect 13920 23259 13960 23291
rect 13992 23259 14032 23291
rect 14064 23259 14104 23291
rect 14136 23259 14176 23291
rect 14208 23259 14248 23291
rect 14280 23259 14320 23291
rect 14352 23259 14392 23291
rect 14424 23259 14464 23291
rect 14496 23259 14536 23291
rect 14568 23259 14608 23291
rect 14640 23259 14680 23291
rect 14712 23259 14752 23291
rect 14784 23259 14824 23291
rect 14856 23259 14896 23291
rect 14928 23259 14968 23291
rect 15000 23259 15040 23291
rect 15072 23259 15112 23291
rect 15144 23259 15184 23291
rect 15216 23259 15256 23291
rect 15288 23259 15328 23291
rect 15360 23259 15400 23291
rect 15432 23259 15472 23291
rect 15504 23259 15544 23291
rect 15576 23259 15616 23291
rect 15648 23259 15688 23291
rect 15720 23259 15760 23291
rect 15792 23259 15832 23291
rect 15864 23259 15904 23291
rect 15936 23259 16000 23291
rect 0 23219 16000 23259
rect 0 23187 64 23219
rect 96 23187 136 23219
rect 168 23187 208 23219
rect 240 23187 280 23219
rect 312 23187 352 23219
rect 384 23187 424 23219
rect 456 23187 496 23219
rect 528 23187 568 23219
rect 600 23187 640 23219
rect 672 23187 712 23219
rect 744 23187 784 23219
rect 816 23187 856 23219
rect 888 23187 928 23219
rect 960 23187 1000 23219
rect 1032 23187 1072 23219
rect 1104 23187 1144 23219
rect 1176 23187 1216 23219
rect 1248 23187 1288 23219
rect 1320 23187 1360 23219
rect 1392 23187 1432 23219
rect 1464 23187 1504 23219
rect 1536 23187 1576 23219
rect 1608 23187 1648 23219
rect 1680 23187 1720 23219
rect 1752 23187 1792 23219
rect 1824 23187 1864 23219
rect 1896 23187 1936 23219
rect 1968 23187 2008 23219
rect 2040 23187 2080 23219
rect 2112 23187 2152 23219
rect 2184 23187 2224 23219
rect 2256 23187 2296 23219
rect 2328 23187 2368 23219
rect 2400 23187 2440 23219
rect 2472 23187 2512 23219
rect 2544 23187 2584 23219
rect 2616 23187 2656 23219
rect 2688 23187 2728 23219
rect 2760 23187 2800 23219
rect 2832 23187 2872 23219
rect 2904 23187 2944 23219
rect 2976 23187 3016 23219
rect 3048 23187 3088 23219
rect 3120 23187 3160 23219
rect 3192 23187 3232 23219
rect 3264 23187 3304 23219
rect 3336 23187 3376 23219
rect 3408 23187 3448 23219
rect 3480 23187 3520 23219
rect 3552 23187 3592 23219
rect 3624 23187 3664 23219
rect 3696 23187 3736 23219
rect 3768 23187 3808 23219
rect 3840 23187 3880 23219
rect 3912 23187 3952 23219
rect 3984 23187 4024 23219
rect 4056 23187 4096 23219
rect 4128 23187 4168 23219
rect 4200 23187 4240 23219
rect 4272 23187 4312 23219
rect 4344 23187 4384 23219
rect 4416 23187 4456 23219
rect 4488 23187 4528 23219
rect 4560 23187 4600 23219
rect 4632 23187 4672 23219
rect 4704 23187 4744 23219
rect 4776 23187 4816 23219
rect 4848 23187 4888 23219
rect 4920 23187 4960 23219
rect 4992 23187 5032 23219
rect 5064 23187 5104 23219
rect 5136 23187 5176 23219
rect 5208 23187 5248 23219
rect 5280 23187 5320 23219
rect 5352 23187 5392 23219
rect 5424 23187 5464 23219
rect 5496 23187 5536 23219
rect 5568 23187 5608 23219
rect 5640 23187 5680 23219
rect 5712 23187 5752 23219
rect 5784 23187 5824 23219
rect 5856 23187 5896 23219
rect 5928 23187 5968 23219
rect 6000 23187 6040 23219
rect 6072 23187 6112 23219
rect 6144 23187 6184 23219
rect 6216 23187 6256 23219
rect 6288 23187 6328 23219
rect 6360 23187 6400 23219
rect 6432 23187 6472 23219
rect 6504 23187 6544 23219
rect 6576 23187 6616 23219
rect 6648 23187 6688 23219
rect 6720 23187 6760 23219
rect 6792 23187 6832 23219
rect 6864 23187 6904 23219
rect 6936 23187 6976 23219
rect 7008 23187 7048 23219
rect 7080 23187 7120 23219
rect 7152 23187 7192 23219
rect 7224 23187 7264 23219
rect 7296 23187 7336 23219
rect 7368 23187 7408 23219
rect 7440 23187 7480 23219
rect 7512 23187 7552 23219
rect 7584 23187 7624 23219
rect 7656 23187 7696 23219
rect 7728 23187 7768 23219
rect 7800 23187 7840 23219
rect 7872 23187 7912 23219
rect 7944 23187 7984 23219
rect 8016 23187 8056 23219
rect 8088 23187 8128 23219
rect 8160 23187 8200 23219
rect 8232 23187 8272 23219
rect 8304 23187 8344 23219
rect 8376 23187 8416 23219
rect 8448 23187 8488 23219
rect 8520 23187 8560 23219
rect 8592 23187 8632 23219
rect 8664 23187 8704 23219
rect 8736 23187 8776 23219
rect 8808 23187 8848 23219
rect 8880 23187 8920 23219
rect 8952 23187 8992 23219
rect 9024 23187 9064 23219
rect 9096 23187 9136 23219
rect 9168 23187 9208 23219
rect 9240 23187 9280 23219
rect 9312 23187 9352 23219
rect 9384 23187 9424 23219
rect 9456 23187 9496 23219
rect 9528 23187 9568 23219
rect 9600 23187 9640 23219
rect 9672 23187 9712 23219
rect 9744 23187 9784 23219
rect 9816 23187 9856 23219
rect 9888 23187 9928 23219
rect 9960 23187 10000 23219
rect 10032 23187 10072 23219
rect 10104 23187 10144 23219
rect 10176 23187 10216 23219
rect 10248 23187 10288 23219
rect 10320 23187 10360 23219
rect 10392 23187 10432 23219
rect 10464 23187 10504 23219
rect 10536 23187 10576 23219
rect 10608 23187 10648 23219
rect 10680 23187 10720 23219
rect 10752 23187 10792 23219
rect 10824 23187 10864 23219
rect 10896 23187 10936 23219
rect 10968 23187 11008 23219
rect 11040 23187 11080 23219
rect 11112 23187 11152 23219
rect 11184 23187 11224 23219
rect 11256 23187 11296 23219
rect 11328 23187 11368 23219
rect 11400 23187 11440 23219
rect 11472 23187 11512 23219
rect 11544 23187 11584 23219
rect 11616 23187 11656 23219
rect 11688 23187 11728 23219
rect 11760 23187 11800 23219
rect 11832 23187 11872 23219
rect 11904 23187 11944 23219
rect 11976 23187 12016 23219
rect 12048 23187 12088 23219
rect 12120 23187 12160 23219
rect 12192 23187 12232 23219
rect 12264 23187 12304 23219
rect 12336 23187 12376 23219
rect 12408 23187 12448 23219
rect 12480 23187 12520 23219
rect 12552 23187 12592 23219
rect 12624 23187 12664 23219
rect 12696 23187 12736 23219
rect 12768 23187 12808 23219
rect 12840 23187 12880 23219
rect 12912 23187 12952 23219
rect 12984 23187 13024 23219
rect 13056 23187 13096 23219
rect 13128 23187 13168 23219
rect 13200 23187 13240 23219
rect 13272 23187 13312 23219
rect 13344 23187 13384 23219
rect 13416 23187 13456 23219
rect 13488 23187 13528 23219
rect 13560 23187 13600 23219
rect 13632 23187 13672 23219
rect 13704 23187 13744 23219
rect 13776 23187 13816 23219
rect 13848 23187 13888 23219
rect 13920 23187 13960 23219
rect 13992 23187 14032 23219
rect 14064 23187 14104 23219
rect 14136 23187 14176 23219
rect 14208 23187 14248 23219
rect 14280 23187 14320 23219
rect 14352 23187 14392 23219
rect 14424 23187 14464 23219
rect 14496 23187 14536 23219
rect 14568 23187 14608 23219
rect 14640 23187 14680 23219
rect 14712 23187 14752 23219
rect 14784 23187 14824 23219
rect 14856 23187 14896 23219
rect 14928 23187 14968 23219
rect 15000 23187 15040 23219
rect 15072 23187 15112 23219
rect 15144 23187 15184 23219
rect 15216 23187 15256 23219
rect 15288 23187 15328 23219
rect 15360 23187 15400 23219
rect 15432 23187 15472 23219
rect 15504 23187 15544 23219
rect 15576 23187 15616 23219
rect 15648 23187 15688 23219
rect 15720 23187 15760 23219
rect 15792 23187 15832 23219
rect 15864 23187 15904 23219
rect 15936 23187 16000 23219
rect 0 23124 16000 23187
rect 0 23121 68 23124
rect 0 23089 18 23121
rect 50 23089 68 23121
rect 0 23053 68 23089
rect 0 23021 18 23053
rect 50 23021 68 23053
rect 0 22984 68 23021
rect 0 22952 18 22984
rect 50 22952 68 22984
rect 0 22915 68 22952
rect 0 22883 18 22915
rect 50 22883 68 22915
rect 0 22846 68 22883
rect 0 22814 18 22846
rect 50 22814 68 22846
rect 0 22777 68 22814
rect 0 22745 18 22777
rect 50 22745 68 22777
rect 0 22708 68 22745
rect 0 22676 18 22708
rect 50 22676 68 22708
rect 0 22639 68 22676
rect 0 22607 18 22639
rect 50 22607 68 22639
rect 0 22570 68 22607
rect 0 22538 18 22570
rect 50 22538 68 22570
rect 0 22501 68 22538
rect 0 22469 18 22501
rect 50 22469 68 22501
rect 0 22432 68 22469
rect 0 22400 18 22432
rect 50 22400 68 22432
rect 0 22363 68 22400
rect 0 22331 18 22363
rect 50 22331 68 22363
rect 0 22294 68 22331
rect 0 22262 18 22294
rect 50 22262 68 22294
rect 0 22225 68 22262
rect 0 22193 18 22225
rect 50 22193 68 22225
rect 0 22156 68 22193
rect 0 22124 18 22156
rect 50 22124 68 22156
rect 0 22087 68 22124
rect 0 22055 18 22087
rect 50 22055 68 22087
rect 0 22018 68 22055
rect 0 21986 18 22018
rect 50 21986 68 22018
rect 0 21949 68 21986
rect 0 21917 18 21949
rect 50 21917 68 21949
rect 0 21880 68 21917
rect 0 21848 18 21880
rect 50 21848 68 21880
rect 0 21811 68 21848
rect 0 21779 18 21811
rect 50 21779 68 21811
rect 0 21742 68 21779
rect 0 21710 18 21742
rect 50 21710 68 21742
rect 0 21673 68 21710
rect 0 21641 18 21673
rect 50 21641 68 21673
rect 0 21604 68 21641
rect 0 21572 18 21604
rect 50 21572 68 21604
rect 0 21535 68 21572
rect 0 21503 18 21535
rect 50 21503 68 21535
rect 0 21466 68 21503
rect 0 21434 18 21466
rect 50 21434 68 21466
rect 0 21397 68 21434
rect 0 21365 18 21397
rect 50 21365 68 21397
rect 0 21328 68 21365
rect 0 21296 18 21328
rect 50 21296 68 21328
rect 0 21259 68 21296
rect 0 21227 18 21259
rect 50 21227 68 21259
rect 0 21190 68 21227
rect 0 21158 18 21190
rect 50 21158 68 21190
rect 0 21121 68 21158
rect 0 21089 18 21121
rect 50 21089 68 21121
rect 0 21052 68 21089
rect 0 21020 18 21052
rect 50 21020 68 21052
rect 0 20983 68 21020
rect 0 20951 18 20983
rect 50 20951 68 20983
rect 0 20914 68 20951
rect 0 20882 18 20914
rect 50 20882 68 20914
rect 0 20845 68 20882
rect 0 20813 18 20845
rect 50 20813 68 20845
rect 0 20776 68 20813
rect 0 20744 18 20776
rect 50 20744 68 20776
rect 0 20707 68 20744
rect 0 20675 18 20707
rect 50 20675 68 20707
rect 0 20638 68 20675
rect 0 20606 18 20638
rect 50 20606 68 20638
rect 0 20569 68 20606
rect 0 20537 18 20569
rect 50 20537 68 20569
rect 0 20500 68 20537
rect 0 20468 18 20500
rect 50 20468 68 20500
rect 0 20431 68 20468
rect 0 20399 18 20431
rect 50 20399 68 20431
rect 0 20362 68 20399
rect 0 20330 18 20362
rect 50 20330 68 20362
rect 0 20293 68 20330
rect 0 20261 18 20293
rect 50 20261 68 20293
rect 0 20224 68 20261
rect 0 20192 18 20224
rect 50 20192 68 20224
rect 0 20155 68 20192
rect 0 20123 18 20155
rect 50 20123 68 20155
rect 0 20086 68 20123
rect 0 20054 18 20086
rect 50 20054 68 20086
rect 0 20017 68 20054
rect 0 19985 18 20017
rect 50 19985 68 20017
rect 0 19948 68 19985
rect 0 19916 18 19948
rect 50 19916 68 19948
rect 0 19879 68 19916
rect 0 19847 18 19879
rect 50 19847 68 19879
rect 0 19810 68 19847
rect 0 19778 18 19810
rect 50 19778 68 19810
rect 0 19741 68 19778
rect 0 19709 18 19741
rect 50 19709 68 19741
rect 0 19672 68 19709
rect 0 19640 18 19672
rect 50 19640 68 19672
rect 0 19603 68 19640
rect 0 19571 18 19603
rect 50 19571 68 19603
rect 0 19534 68 19571
rect 0 19502 18 19534
rect 50 19502 68 19534
rect 0 19465 68 19502
rect 0 19433 18 19465
rect 50 19433 68 19465
rect 0 19396 68 19433
rect 0 19364 18 19396
rect 50 19364 68 19396
rect 0 19327 68 19364
rect 0 19295 18 19327
rect 50 19295 68 19327
rect 0 19258 68 19295
rect 0 19226 18 19258
rect 50 19226 68 19258
rect 0 19189 68 19226
rect 0 19157 18 19189
rect 50 19157 68 19189
rect 0 19120 68 19157
rect 0 19088 18 19120
rect 50 19088 68 19120
rect 0 19051 68 19088
rect 0 19019 18 19051
rect 50 19019 68 19051
rect 0 18982 68 19019
rect 0 18950 18 18982
rect 50 18950 68 18982
rect 0 18913 68 18950
rect 0 18881 18 18913
rect 50 18881 68 18913
rect 0 18844 68 18881
rect 0 18812 18 18844
rect 50 18812 68 18844
rect 0 18775 68 18812
rect 0 18743 18 18775
rect 50 18743 68 18775
rect 0 18706 68 18743
rect 0 18674 18 18706
rect 50 18674 68 18706
rect 0 18637 68 18674
rect 0 18605 18 18637
rect 50 18605 68 18637
rect 0 18568 68 18605
rect 0 18536 18 18568
rect 50 18536 68 18568
rect 0 18499 68 18536
rect 0 18467 18 18499
rect 50 18467 68 18499
rect 0 18430 68 18467
rect 0 18398 18 18430
rect 50 18398 68 18430
rect 0 18361 68 18398
rect 0 18329 18 18361
rect 50 18329 68 18361
rect 0 18292 68 18329
rect 0 18260 18 18292
rect 50 18260 68 18292
rect 0 18223 68 18260
rect 0 18191 18 18223
rect 50 18191 68 18223
rect 0 18154 68 18191
rect 0 18122 18 18154
rect 50 18122 68 18154
rect 0 18085 68 18122
rect 0 18053 18 18085
rect 50 18053 68 18085
rect 0 18016 68 18053
rect 0 17984 18 18016
rect 50 17984 68 18016
rect 0 17947 68 17984
rect 0 17915 18 17947
rect 50 17915 68 17947
rect 0 17878 68 17915
rect 0 17846 18 17878
rect 50 17846 68 17878
rect 0 17809 68 17846
rect 0 17777 18 17809
rect 50 17777 68 17809
rect 0 17740 68 17777
rect 0 17708 18 17740
rect 50 17708 68 17740
rect 0 17671 68 17708
rect 0 17639 18 17671
rect 50 17639 68 17671
rect 0 17602 68 17639
rect 0 17570 18 17602
rect 50 17570 68 17602
rect 0 17534 68 17570
rect 0 17502 18 17534
rect 50 17502 68 17534
rect 0 13000 68 17502
rect 15934 23110 16000 23124
rect 15934 23078 15951 23110
rect 15983 23078 16000 23110
rect 15934 23042 16000 23078
rect 15934 23010 15951 23042
rect 15983 23010 16000 23042
rect 15934 22974 16000 23010
rect 15934 22942 15951 22974
rect 15983 22942 16000 22974
rect 15934 22906 16000 22942
rect 15934 22874 15951 22906
rect 15983 22874 16000 22906
rect 15934 22838 16000 22874
rect 15934 22806 15951 22838
rect 15983 22806 16000 22838
rect 15934 22770 16000 22806
rect 15934 22738 15951 22770
rect 15983 22738 16000 22770
rect 15934 22702 16000 22738
rect 15934 22670 15951 22702
rect 15983 22670 16000 22702
rect 15934 22634 16000 22670
rect 15934 22602 15951 22634
rect 15983 22602 16000 22634
rect 15934 22566 16000 22602
rect 15934 22534 15951 22566
rect 15983 22534 16000 22566
rect 15934 22498 16000 22534
rect 15934 22466 15951 22498
rect 15983 22466 16000 22498
rect 15934 22430 16000 22466
rect 15934 22398 15951 22430
rect 15983 22398 16000 22430
rect 15934 22362 16000 22398
rect 15934 22330 15951 22362
rect 15983 22330 16000 22362
rect 15934 22294 16000 22330
rect 15934 22262 15951 22294
rect 15983 22262 16000 22294
rect 15934 22226 16000 22262
rect 15934 22194 15951 22226
rect 15983 22194 16000 22226
rect 15934 22158 16000 22194
rect 15934 22126 15951 22158
rect 15983 22126 16000 22158
rect 15934 22090 16000 22126
rect 15934 22058 15951 22090
rect 15983 22058 16000 22090
rect 15934 22022 16000 22058
rect 15934 21990 15951 22022
rect 15983 21990 16000 22022
rect 15934 21954 16000 21990
rect 15934 21922 15951 21954
rect 15983 21922 16000 21954
rect 15934 21886 16000 21922
rect 15934 21854 15951 21886
rect 15983 21854 16000 21886
rect 15934 21818 16000 21854
rect 15934 21786 15951 21818
rect 15983 21786 16000 21818
rect 15934 21750 16000 21786
rect 15934 21718 15951 21750
rect 15983 21718 16000 21750
rect 15934 21682 16000 21718
rect 15934 21650 15951 21682
rect 15983 21650 16000 21682
rect 15934 21614 16000 21650
rect 15934 21582 15951 21614
rect 15983 21582 16000 21614
rect 15934 21546 16000 21582
rect 15934 21514 15951 21546
rect 15983 21514 16000 21546
rect 15934 21478 16000 21514
rect 15934 21446 15951 21478
rect 15983 21446 16000 21478
rect 15934 21410 16000 21446
rect 15934 21378 15951 21410
rect 15983 21378 16000 21410
rect 15934 21342 16000 21378
rect 15934 21310 15951 21342
rect 15983 21310 16000 21342
rect 15934 21274 16000 21310
rect 15934 21242 15951 21274
rect 15983 21242 16000 21274
rect 15934 21206 16000 21242
rect 15934 21174 15951 21206
rect 15983 21174 16000 21206
rect 15934 21138 16000 21174
rect 15934 21106 15951 21138
rect 15983 21106 16000 21138
rect 15934 21070 16000 21106
rect 15934 21038 15951 21070
rect 15983 21038 16000 21070
rect 15934 21002 16000 21038
rect 15934 20970 15951 21002
rect 15983 20970 16000 21002
rect 15934 20934 16000 20970
rect 15934 20902 15951 20934
rect 15983 20902 16000 20934
rect 15934 20866 16000 20902
rect 15934 20834 15951 20866
rect 15983 20834 16000 20866
rect 15934 20798 16000 20834
rect 15934 20766 15951 20798
rect 15983 20766 16000 20798
rect 15934 20730 16000 20766
rect 15934 20698 15951 20730
rect 15983 20698 16000 20730
rect 15934 20662 16000 20698
rect 15934 20630 15951 20662
rect 15983 20630 16000 20662
rect 15934 20594 16000 20630
rect 15934 20562 15951 20594
rect 15983 20562 16000 20594
rect 15934 20526 16000 20562
rect 15934 20494 15951 20526
rect 15983 20494 16000 20526
rect 15934 20458 16000 20494
rect 15934 20426 15951 20458
rect 15983 20426 16000 20458
rect 15934 20390 16000 20426
rect 15934 20358 15951 20390
rect 15983 20358 16000 20390
rect 15934 20322 16000 20358
rect 15934 20290 15951 20322
rect 15983 20290 16000 20322
rect 15934 20254 16000 20290
rect 15934 20222 15951 20254
rect 15983 20222 16000 20254
rect 15934 20186 16000 20222
rect 15934 20154 15951 20186
rect 15983 20154 16000 20186
rect 15934 20118 16000 20154
rect 15934 20086 15951 20118
rect 15983 20086 16000 20118
rect 15934 20050 16000 20086
rect 15934 20018 15951 20050
rect 15983 20018 16000 20050
rect 15934 19982 16000 20018
rect 15934 19950 15951 19982
rect 15983 19950 16000 19982
rect 15934 19914 16000 19950
rect 15934 19882 15951 19914
rect 15983 19882 16000 19914
rect 15934 19846 16000 19882
rect 15934 19814 15951 19846
rect 15983 19814 16000 19846
rect 15934 19778 16000 19814
rect 15934 19746 15951 19778
rect 15983 19746 16000 19778
rect 15934 19710 16000 19746
rect 15934 19678 15951 19710
rect 15983 19678 16000 19710
rect 15934 19642 16000 19678
rect 15934 19610 15951 19642
rect 15983 19610 16000 19642
rect 15934 19574 16000 19610
rect 15934 19542 15951 19574
rect 15983 19542 16000 19574
rect 15934 19506 16000 19542
rect 15934 19474 15951 19506
rect 15983 19474 16000 19506
rect 15934 19438 16000 19474
rect 15934 19406 15951 19438
rect 15983 19406 16000 19438
rect 15934 19370 16000 19406
rect 15934 19338 15951 19370
rect 15983 19338 16000 19370
rect 15934 19302 16000 19338
rect 15934 19270 15951 19302
rect 15983 19270 16000 19302
rect 15934 19234 16000 19270
rect 15934 19202 15951 19234
rect 15983 19202 16000 19234
rect 15934 19166 16000 19202
rect 15934 19134 15951 19166
rect 15983 19134 16000 19166
rect 15934 19098 16000 19134
rect 15934 19066 15951 19098
rect 15983 19066 16000 19098
rect 15934 19030 16000 19066
rect 15934 18998 15951 19030
rect 15983 18998 16000 19030
rect 15934 18962 16000 18998
rect 15934 18930 15951 18962
rect 15983 18930 16000 18962
rect 15934 18894 16000 18930
rect 15934 18862 15951 18894
rect 15983 18862 16000 18894
rect 15934 18826 16000 18862
rect 15934 18794 15951 18826
rect 15983 18794 16000 18826
rect 15934 18758 16000 18794
rect 15934 18726 15951 18758
rect 15983 18726 16000 18758
rect 15934 18690 16000 18726
rect 15934 18658 15951 18690
rect 15983 18658 16000 18690
rect 15934 18622 16000 18658
rect 15934 18590 15951 18622
rect 15983 18590 16000 18622
rect 15934 18554 16000 18590
rect 15934 18522 15951 18554
rect 15983 18522 16000 18554
rect 15934 18486 16000 18522
rect 15934 18454 15951 18486
rect 15983 18454 16000 18486
rect 15934 18418 16000 18454
rect 15934 18386 15951 18418
rect 15983 18386 16000 18418
rect 15934 18350 16000 18386
rect 15934 18318 15951 18350
rect 15983 18318 16000 18350
rect 15934 18282 16000 18318
rect 15934 18250 15951 18282
rect 15983 18250 16000 18282
rect 15934 18214 16000 18250
rect 15934 18182 15951 18214
rect 15983 18182 16000 18214
rect 15934 18146 16000 18182
rect 15934 18114 15951 18146
rect 15983 18114 16000 18146
rect 15934 18078 16000 18114
rect 15934 18046 15951 18078
rect 15983 18046 16000 18078
rect 15934 18010 16000 18046
rect 15934 17978 15951 18010
rect 15983 17978 16000 18010
rect 15934 17942 16000 17978
rect 15934 17910 15951 17942
rect 15983 17910 16000 17942
rect 15934 17874 16000 17910
rect 15934 17842 15951 17874
rect 15983 17842 16000 17874
rect 15934 17806 16000 17842
rect 15934 17774 15951 17806
rect 15983 17774 16000 17806
rect 15934 17738 16000 17774
rect 15934 17706 15951 17738
rect 15983 17706 16000 17738
rect 15934 17670 16000 17706
rect 15934 17638 15951 17670
rect 15983 17638 16000 17670
rect 15934 17602 16000 17638
rect 15934 17570 15951 17602
rect 15983 17570 16000 17602
rect 15934 17534 16000 17570
rect 15934 17502 15951 17534
rect 15983 17502 16000 17534
rect 15934 13000 16000 17502
<< nsubdiff >>
rect 118 33384 150 33416
rect 186 33384 218 33416
rect 254 33384 286 33416
rect 322 33384 354 33416
rect 390 33384 422 33416
rect 458 33384 490 33416
rect 526 33384 558 33416
rect 594 33384 626 33416
rect 662 33384 694 33416
rect 730 33384 762 33416
rect 798 33384 830 33416
rect 866 33384 898 33416
rect 934 33384 966 33416
rect 1002 33384 1034 33416
rect 1070 33384 1102 33416
rect 1138 33384 1170 33416
rect 1206 33384 1238 33416
rect 1274 33384 1306 33416
rect 1342 33384 1374 33416
rect 1410 33384 1442 33416
rect 1478 33384 1510 33416
rect 1546 33384 1578 33416
rect 1614 33384 1646 33416
rect 1682 33384 1714 33416
rect 1750 33384 1782 33416
rect 1818 33384 1850 33416
rect 1886 33384 1918 33416
rect 1954 33384 1986 33416
rect 2022 33384 2054 33416
rect 2090 33384 2122 33416
rect 2158 33384 2190 33416
rect 2226 33384 2258 33416
rect 2294 33384 2326 33416
rect 2362 33384 2394 33416
rect 2430 33384 2462 33416
rect 2498 33384 2530 33416
rect 2566 33384 2598 33416
rect 2634 33384 2666 33416
rect 2702 33384 2734 33416
rect 2770 33384 2802 33416
rect 2838 33384 2870 33416
rect 2906 33384 2938 33416
rect 2974 33384 3006 33416
rect 3042 33384 3074 33416
rect 3110 33384 3142 33416
rect 3178 33384 3210 33416
rect 3246 33384 3278 33416
rect 3314 33384 3346 33416
rect 3382 33384 3414 33416
rect 3450 33384 3482 33416
rect 3518 33384 3550 33416
rect 3586 33384 3618 33416
rect 3654 33384 3686 33416
rect 3722 33384 3754 33416
rect 3790 33384 3822 33416
rect 3858 33384 3890 33416
rect 3926 33384 3958 33416
rect 3994 33384 4026 33416
rect 4062 33384 4094 33416
rect 4130 33384 4162 33416
rect 4198 33384 4230 33416
rect 4266 33384 4298 33416
rect 4334 33384 4366 33416
rect 4402 33384 4434 33416
rect 4470 33384 4502 33416
rect 4538 33384 4570 33416
rect 4606 33384 4638 33416
rect 4674 33384 4706 33416
rect 4742 33384 4774 33416
rect 4810 33384 4842 33416
rect 4878 33384 4910 33416
rect 4946 33384 4978 33416
rect 5014 33384 5046 33416
rect 5082 33384 5114 33416
rect 5150 33384 5182 33416
rect 5218 33384 5250 33416
rect 5286 33384 5318 33416
rect 5354 33384 5386 33416
rect 5422 33384 5454 33416
rect 5490 33384 5522 33416
rect 5558 33384 5590 33416
rect 5626 33384 5658 33416
rect 5694 33384 5726 33416
rect 5762 33384 5794 33416
rect 5830 33384 5862 33416
rect 5898 33384 5930 33416
rect 5966 33384 5998 33416
rect 6034 33384 6066 33416
rect 6102 33384 6134 33416
rect 6170 33384 6202 33416
rect 6238 33384 6270 33416
rect 6306 33384 6338 33416
rect 6374 33384 6406 33416
rect 6442 33384 6474 33416
rect 6510 33384 6542 33416
rect 6578 33384 6610 33416
rect 6646 33384 6678 33416
rect 6714 33384 6746 33416
rect 6782 33384 6814 33416
rect 6850 33384 6882 33416
rect 6918 33384 6950 33416
rect 6986 33384 7018 33416
rect 7054 33384 7086 33416
rect 7122 33384 7154 33416
rect 7190 33384 7222 33416
rect 7258 33384 7290 33416
rect 7326 33384 7358 33416
rect 7394 33384 7426 33416
rect 7462 33384 7494 33416
rect 7530 33384 7562 33416
rect 7598 33384 7630 33416
rect 7666 33384 7698 33416
rect 7734 33384 7766 33416
rect 7802 33384 7834 33416
rect 7870 33384 7902 33416
rect 7938 33384 7970 33416
rect 8006 33384 8038 33416
rect 8074 33384 8106 33416
rect 8142 33384 8174 33416
rect 8210 33384 8242 33416
rect 8278 33384 8310 33416
rect 8346 33384 8378 33416
rect 8414 33384 8446 33416
rect 8482 33384 8514 33416
rect 8550 33384 8582 33416
rect 8618 33384 8650 33416
rect 8686 33384 8718 33416
rect 8754 33384 8786 33416
rect 8822 33384 8854 33416
rect 8890 33384 8922 33416
rect 8958 33384 8990 33416
rect 9026 33384 9058 33416
rect 9094 33384 9126 33416
rect 9162 33384 9194 33416
rect 9230 33384 9262 33416
rect 9298 33384 9330 33416
rect 9366 33384 9398 33416
rect 9434 33384 9466 33416
rect 9502 33384 9534 33416
rect 9570 33384 9602 33416
rect 9638 33384 9670 33416
rect 9706 33384 9738 33416
rect 9774 33384 9806 33416
rect 9842 33384 9874 33416
rect 9910 33384 9942 33416
rect 9978 33384 10010 33416
rect 10046 33384 10078 33416
rect 10114 33384 10146 33416
rect 10182 33384 10214 33416
rect 10250 33384 10282 33416
rect 10318 33384 10350 33416
rect 10386 33384 10418 33416
rect 10454 33384 10486 33416
rect 10522 33384 10554 33416
rect 10590 33384 10622 33416
rect 10658 33384 10690 33416
rect 10726 33384 10758 33416
rect 10794 33384 10826 33416
rect 10862 33384 10894 33416
rect 10930 33384 10962 33416
rect 10998 33384 11030 33416
rect 11066 33384 11098 33416
rect 11134 33384 11166 33416
rect 11202 33384 11234 33416
rect 11270 33384 11302 33416
rect 11338 33384 11370 33416
rect 11406 33384 11438 33416
rect 11474 33384 11506 33416
rect 11542 33384 11574 33416
rect 11610 33384 11642 33416
rect 11678 33384 11710 33416
rect 11746 33384 11778 33416
rect 11814 33384 11846 33416
rect 11882 33384 11914 33416
rect 11950 33384 11982 33416
rect 12018 33384 12050 33416
rect 12086 33384 12118 33416
rect 12154 33384 12186 33416
rect 12222 33384 12254 33416
rect 12290 33384 12322 33416
rect 12358 33384 12390 33416
rect 12426 33384 12458 33416
rect 12494 33384 12526 33416
rect 12562 33384 12594 33416
rect 12630 33384 12662 33416
rect 12698 33384 12730 33416
rect 12766 33384 12798 33416
rect 12834 33384 12866 33416
rect 12902 33384 12934 33416
rect 12970 33384 13002 33416
rect 13038 33384 13070 33416
rect 13106 33384 13138 33416
rect 13174 33384 13206 33416
rect 13242 33384 13274 33416
rect 13310 33384 13342 33416
rect 13378 33384 13410 33416
rect 13446 33384 13478 33416
rect 13514 33384 13546 33416
rect 13582 33384 13614 33416
rect 13650 33384 13682 33416
rect 13718 33384 13750 33416
rect 13786 33384 13818 33416
rect 13854 33384 13886 33416
rect 13922 33384 13954 33416
rect 13990 33384 14022 33416
rect 14058 33384 14090 33416
rect 14126 33384 14158 33416
rect 14194 33384 14226 33416
rect 14262 33384 14294 33416
rect 14330 33384 14362 33416
rect 14398 33384 14430 33416
rect 14466 33384 14498 33416
rect 14534 33384 14566 33416
rect 14602 33384 14634 33416
rect 14670 33384 14702 33416
rect 14738 33384 14770 33416
rect 14806 33384 14838 33416
rect 14874 33384 14906 33416
rect 14942 33384 14974 33416
rect 15010 33384 15042 33416
rect 15078 33384 15110 33416
rect 15146 33384 15178 33416
rect 15214 33384 15246 33416
rect 15282 33384 15314 33416
rect 15350 33384 15382 33416
rect 15442 33384 15474 33416
rect 15510 33384 15542 33416
rect 15578 33384 15610 33416
rect 15646 33384 15678 33416
rect 15714 33384 15746 33416
rect 15782 33384 15814 33416
rect 15850 33384 15882 33416
rect 15918 33384 15950 33416
rect 118 29684 150 29716
rect 186 29684 218 29716
rect 254 29684 286 29716
rect 322 29684 354 29716
rect 390 29684 422 29716
rect 458 29684 490 29716
rect 526 29684 558 29716
rect 594 29684 626 29716
rect 662 29684 694 29716
rect 730 29684 762 29716
rect 798 29684 830 29716
rect 866 29684 898 29716
rect 934 29684 966 29716
rect 1002 29684 1034 29716
rect 1070 29684 1102 29716
rect 1138 29684 1170 29716
rect 1206 29684 1238 29716
rect 1274 29684 1306 29716
rect 1342 29684 1374 29716
rect 1410 29684 1442 29716
rect 1478 29684 1510 29716
rect 1546 29684 1578 29716
rect 1614 29684 1646 29716
rect 1682 29684 1714 29716
rect 1750 29684 1782 29716
rect 1818 29684 1850 29716
rect 1886 29684 1918 29716
rect 1954 29684 1986 29716
rect 2022 29684 2054 29716
rect 2090 29684 2122 29716
rect 2158 29684 2190 29716
rect 2226 29684 2258 29716
rect 2294 29684 2326 29716
rect 2362 29684 2394 29716
rect 2430 29684 2462 29716
rect 2498 29684 2530 29716
rect 2566 29684 2598 29716
rect 2634 29684 2666 29716
rect 2702 29684 2734 29716
rect 2770 29684 2802 29716
rect 2838 29684 2870 29716
rect 2906 29684 2938 29716
rect 2974 29684 3006 29716
rect 3042 29684 3074 29716
rect 3110 29684 3142 29716
rect 3178 29684 3210 29716
rect 3246 29684 3278 29716
rect 3314 29684 3346 29716
rect 3382 29684 3414 29716
rect 3450 29684 3482 29716
rect 3518 29684 3550 29716
rect 3586 29684 3618 29716
rect 3654 29684 3686 29716
rect 3722 29684 3754 29716
rect 3790 29684 3822 29716
rect 3858 29684 3890 29716
rect 3926 29684 3958 29716
rect 3994 29684 4026 29716
rect 4062 29684 4094 29716
rect 4130 29684 4162 29716
rect 4198 29684 4230 29716
rect 4266 29684 4298 29716
rect 4334 29684 4366 29716
rect 4402 29684 4434 29716
rect 4470 29684 4502 29716
rect 4538 29684 4570 29716
rect 4606 29684 4638 29716
rect 4674 29684 4706 29716
rect 4742 29684 4774 29716
rect 4810 29684 4842 29716
rect 4878 29684 4910 29716
rect 4946 29684 4978 29716
rect 5014 29684 5046 29716
rect 5082 29684 5114 29716
rect 5150 29684 5182 29716
rect 5218 29684 5250 29716
rect 5286 29684 5318 29716
rect 5354 29684 5386 29716
rect 5422 29684 5454 29716
rect 5490 29684 5522 29716
rect 5558 29684 5590 29716
rect 5626 29684 5658 29716
rect 5694 29684 5726 29716
rect 5762 29684 5794 29716
rect 5830 29684 5862 29716
rect 5898 29684 5930 29716
rect 5966 29684 5998 29716
rect 6034 29684 6066 29716
rect 6102 29684 6134 29716
rect 6170 29684 6202 29716
rect 6238 29684 6270 29716
rect 6306 29684 6338 29716
rect 6374 29684 6406 29716
rect 6442 29684 6474 29716
rect 6510 29684 6542 29716
rect 6578 29684 6610 29716
rect 6646 29684 6678 29716
rect 6714 29684 6746 29716
rect 6782 29684 6814 29716
rect 6850 29684 6882 29716
rect 6918 29684 6950 29716
rect 6986 29684 7018 29716
rect 7054 29684 7086 29716
rect 7122 29684 7154 29716
rect 7190 29684 7222 29716
rect 7258 29684 7290 29716
rect 7326 29684 7358 29716
rect 7394 29684 7426 29716
rect 7462 29684 7494 29716
rect 7530 29684 7562 29716
rect 7598 29684 7630 29716
rect 7666 29684 7698 29716
rect 7734 29684 7766 29716
rect 7802 29684 7834 29716
rect 7870 29684 7902 29716
rect 7938 29684 7970 29716
rect 8006 29684 8038 29716
rect 8074 29684 8106 29716
rect 8142 29684 8174 29716
rect 8210 29684 8242 29716
rect 8278 29684 8310 29716
rect 8346 29684 8378 29716
rect 8414 29684 8446 29716
rect 8482 29684 8514 29716
rect 8550 29684 8582 29716
rect 8618 29684 8650 29716
rect 8686 29684 8718 29716
rect 8754 29684 8786 29716
rect 8822 29684 8854 29716
rect 8890 29684 8922 29716
rect 8958 29684 8990 29716
rect 9026 29684 9058 29716
rect 9094 29684 9126 29716
rect 9162 29684 9194 29716
rect 9230 29684 9262 29716
rect 9298 29684 9330 29716
rect 9366 29684 9398 29716
rect 9434 29684 9466 29716
rect 9502 29684 9534 29716
rect 9570 29684 9602 29716
rect 9638 29684 9670 29716
rect 9706 29684 9738 29716
rect 9774 29684 9806 29716
rect 9842 29684 9874 29716
rect 9910 29684 9942 29716
rect 9978 29684 10010 29716
rect 10046 29684 10078 29716
rect 10114 29684 10146 29716
rect 10182 29684 10214 29716
rect 10250 29684 10282 29716
rect 10318 29684 10350 29716
rect 10386 29684 10418 29716
rect 10454 29684 10486 29716
rect 10522 29684 10554 29716
rect 10590 29684 10622 29716
rect 10658 29684 10690 29716
rect 10726 29684 10758 29716
rect 10794 29684 10826 29716
rect 10862 29684 10894 29716
rect 10930 29684 10962 29716
rect 10998 29684 11030 29716
rect 11066 29684 11098 29716
rect 11134 29684 11166 29716
rect 11202 29684 11234 29716
rect 11270 29684 11302 29716
rect 11338 29684 11370 29716
rect 11406 29684 11438 29716
rect 11474 29684 11506 29716
rect 11542 29684 11574 29716
rect 11610 29684 11642 29716
rect 11678 29684 11710 29716
rect 11746 29684 11778 29716
rect 11814 29684 11846 29716
rect 11882 29684 11914 29716
rect 11950 29684 11982 29716
rect 12018 29684 12050 29716
rect 12086 29684 12118 29716
rect 12154 29684 12186 29716
rect 12222 29684 12254 29716
rect 12290 29684 12322 29716
rect 12358 29684 12390 29716
rect 12426 29684 12458 29716
rect 12494 29684 12526 29716
rect 12562 29684 12594 29716
rect 12630 29684 12662 29716
rect 12698 29684 12730 29716
rect 12766 29684 12798 29716
rect 12834 29684 12866 29716
rect 12902 29684 12934 29716
rect 12970 29684 13002 29716
rect 13038 29684 13070 29716
rect 13106 29684 13138 29716
rect 13174 29684 13206 29716
rect 13242 29684 13274 29716
rect 13310 29684 13342 29716
rect 13378 29684 13410 29716
rect 13446 29684 13478 29716
rect 13514 29684 13546 29716
rect 13582 29684 13614 29716
rect 13650 29684 13682 29716
rect 13718 29684 13750 29716
rect 13786 29684 13818 29716
rect 13854 29684 13886 29716
rect 13922 29684 13954 29716
rect 13990 29684 14022 29716
rect 14058 29684 14090 29716
rect 14126 29684 14158 29716
rect 14194 29684 14226 29716
rect 14262 29684 14294 29716
rect 14330 29684 14362 29716
rect 14398 29684 14430 29716
rect 14466 29684 14498 29716
rect 14534 29684 14566 29716
rect 14602 29684 14634 29716
rect 14670 29684 14702 29716
rect 14738 29684 14770 29716
rect 14806 29684 14838 29716
rect 14874 29684 14906 29716
rect 14942 29684 14974 29716
rect 15010 29684 15042 29716
rect 15078 29684 15110 29716
rect 15146 29684 15178 29716
rect 15214 29684 15246 29716
rect 15282 29684 15314 29716
rect 15350 29684 15382 29716
rect 15442 29684 15474 29716
rect 15510 29684 15542 29716
rect 15578 29684 15610 29716
rect 15646 29684 15678 29716
rect 15714 29684 15746 29716
rect 15782 29684 15814 29716
rect 15850 29684 15882 29716
rect 15918 29684 15950 29716
rect 96 12658 128 12690
rect 164 12658 196 12690
rect 232 12658 264 12690
rect 300 12658 332 12690
rect 368 12658 400 12690
rect 436 12658 468 12690
rect 504 12658 536 12690
rect 572 12658 604 12690
rect 640 12658 672 12690
rect 708 12658 740 12690
rect 776 12658 808 12690
rect 844 12658 876 12690
rect 912 12658 944 12690
rect 980 12658 1012 12690
rect 1048 12658 1080 12690
rect 1116 12658 1148 12690
rect 1184 12658 1216 12690
rect 1252 12658 1284 12690
rect 1320 12658 1352 12690
rect 1388 12658 1420 12690
rect 1456 12658 1488 12690
rect 1524 12658 1556 12690
rect 1592 12658 1624 12690
rect 1660 12658 1692 12690
rect 1728 12658 1760 12690
rect 1796 12658 1828 12690
rect 1864 12658 1896 12690
rect 1932 12658 1964 12690
rect 2000 12658 2032 12690
rect 2068 12658 2100 12690
rect 2136 12658 2168 12690
rect 2204 12658 2236 12690
rect 2272 12658 2304 12690
rect 2340 12658 2372 12690
rect 2408 12658 2440 12690
rect 2476 12658 2508 12690
rect 2544 12658 2576 12690
rect 2612 12658 2644 12690
rect 2680 12658 2712 12690
rect 2748 12658 2780 12690
rect 2816 12658 2848 12690
rect 2884 12658 2916 12690
rect 2952 12658 2984 12690
rect 3020 12658 3052 12690
rect 3088 12658 3120 12690
rect 3156 12658 3188 12690
rect 3224 12658 3256 12690
rect 3292 12658 3324 12690
rect 3360 12658 3392 12690
rect 3428 12658 3460 12690
rect 3496 12658 3528 12690
rect 3564 12658 3596 12690
rect 3632 12658 3664 12690
rect 3700 12658 3732 12690
rect 3768 12658 3800 12690
rect 3836 12658 3868 12690
rect 3904 12658 3936 12690
rect 3972 12658 4004 12690
rect 4040 12658 4072 12690
rect 4108 12658 4140 12690
rect 4176 12658 4208 12690
rect 4244 12658 4276 12690
rect 4312 12658 4344 12690
rect 4380 12658 4412 12690
rect 4448 12658 4480 12690
rect 4516 12658 4548 12690
rect 4584 12658 4616 12690
rect 4652 12658 4684 12690
rect 4720 12658 4752 12690
rect 4788 12658 4820 12690
rect 4856 12658 4888 12690
rect 4924 12658 4956 12690
rect 4992 12658 5024 12690
rect 5060 12658 5092 12690
rect 5128 12658 5160 12690
rect 5196 12658 5228 12690
rect 5264 12658 5296 12690
rect 5332 12658 5364 12690
rect 5400 12658 5432 12690
rect 5468 12658 5500 12690
rect 5536 12658 5568 12690
rect 5604 12658 5636 12690
rect 5672 12658 5704 12690
rect 5740 12658 5772 12690
rect 5808 12658 5840 12690
rect 5876 12658 5908 12690
rect 5944 12658 5976 12690
rect 6012 12658 6044 12690
rect 6080 12658 6112 12690
rect 6148 12658 6180 12690
rect 6216 12658 6248 12690
rect 6284 12658 6316 12690
rect 6352 12658 6384 12690
rect 6420 12658 6452 12690
rect 6488 12658 6520 12690
rect 6556 12658 6588 12690
rect 6624 12658 6656 12690
rect 6692 12658 6724 12690
rect 6760 12658 6792 12690
rect 6828 12658 6860 12690
rect 6896 12658 6928 12690
rect 6964 12658 6996 12690
rect 7032 12658 7064 12690
rect 7100 12658 7132 12690
rect 7168 12658 7200 12690
rect 7236 12658 7268 12690
rect 7304 12658 7336 12690
rect 7372 12658 7404 12690
rect 7440 12658 7472 12690
rect 7508 12658 7540 12690
rect 7576 12658 7608 12690
rect 7644 12658 7676 12690
rect 7712 12658 7744 12690
rect 7780 12658 7812 12690
rect 7848 12658 7880 12690
rect 7916 12658 7948 12690
rect 7984 12658 8016 12690
rect 8052 12658 8084 12690
rect 8120 12658 8152 12690
rect 8188 12658 8220 12690
rect 8256 12658 8288 12690
rect 8324 12658 8356 12690
rect 8392 12658 8424 12690
rect 8460 12658 8492 12690
rect 8528 12658 8560 12690
rect 8596 12658 8628 12690
rect 8664 12658 8696 12690
rect 8732 12658 8764 12690
rect 8800 12658 8832 12690
rect 8868 12658 8900 12690
rect 8936 12658 8968 12690
rect 9004 12658 9036 12690
rect 9072 12658 9104 12690
rect 9140 12658 9172 12690
rect 9208 12658 9240 12690
rect 9276 12658 9308 12690
rect 9344 12658 9376 12690
rect 9412 12658 9444 12690
rect 9480 12658 9512 12690
rect 9548 12658 9580 12690
rect 9616 12658 9648 12690
rect 9684 12658 9716 12690
rect 9752 12658 9784 12690
rect 9820 12658 9852 12690
rect 9888 12658 9920 12690
rect 9956 12658 9988 12690
rect 10024 12658 10056 12690
rect 10092 12658 10124 12690
rect 10160 12658 10192 12690
rect 10228 12658 10260 12690
rect 10296 12658 10328 12690
rect 10364 12658 10396 12690
rect 10432 12658 10464 12690
rect 10500 12658 10532 12690
rect 10568 12658 10600 12690
rect 10636 12658 10668 12690
rect 10704 12658 10736 12690
rect 10772 12658 10804 12690
rect 10840 12658 10872 12690
rect 10908 12658 10940 12690
rect 10976 12658 11008 12690
rect 11044 12658 11076 12690
rect 11112 12658 11144 12690
rect 11180 12658 11212 12690
rect 11248 12658 11280 12690
rect 11316 12658 11348 12690
rect 11384 12658 11416 12690
rect 11452 12658 11484 12690
rect 11520 12658 11552 12690
rect 11588 12658 11620 12690
rect 11656 12658 11688 12690
rect 11724 12658 11756 12690
rect 11792 12658 11824 12690
rect 11860 12658 11892 12690
rect 11928 12658 11960 12690
rect 11996 12658 12028 12690
rect 12064 12658 12096 12690
rect 12132 12658 12164 12690
rect 12200 12658 12232 12690
rect 12268 12658 12300 12690
rect 12336 12658 12368 12690
rect 12404 12658 12436 12690
rect 12472 12658 12504 12690
rect 12540 12658 12572 12690
rect 12608 12658 12640 12690
rect 12676 12658 12708 12690
rect 12744 12658 12776 12690
rect 12812 12658 12844 12690
rect 12880 12658 12912 12690
rect 12948 12658 12980 12690
rect 13016 12658 13048 12690
rect 13084 12658 13116 12690
rect 13152 12658 13184 12690
rect 13220 12658 13252 12690
rect 13288 12658 13320 12690
rect 13356 12658 13388 12690
rect 13424 12658 13456 12690
rect 13492 12658 13524 12690
rect 13560 12658 13592 12690
rect 13628 12658 13660 12690
rect 13696 12658 13728 12690
rect 13764 12658 13796 12690
rect 13832 12658 13864 12690
rect 13900 12658 13932 12690
rect 13968 12658 14000 12690
rect 14036 12658 14068 12690
rect 14104 12658 14136 12690
rect 14172 12658 14204 12690
rect 14240 12658 14272 12690
rect 14308 12658 14340 12690
rect 14376 12658 14408 12690
rect 14444 12658 14476 12690
rect 14512 12658 14544 12690
rect 14580 12658 14612 12690
rect 14648 12658 14680 12690
rect 14716 12658 14748 12690
rect 14784 12658 14816 12690
rect 14852 12658 14884 12690
rect 14920 12658 14952 12690
rect 14988 12658 15020 12690
rect 15056 12658 15088 12690
rect 15124 12658 15156 12690
rect 15192 12658 15224 12690
rect 15260 12658 15292 12690
rect 15328 12658 15360 12690
rect 15396 12658 15428 12690
rect 15464 12658 15496 12690
rect 15532 12658 15564 12690
rect 15600 12658 15632 12690
rect 15668 12658 15700 12690
rect 15736 12658 15768 12690
rect 15804 12658 15836 12690
rect 15872 12658 15904 12690
rect 15940 12658 15972 12690
rect 18 12474 50 12506
rect 18 12406 50 12438
rect 18 12338 50 12370
rect 18 12270 50 12302
rect 18 12202 50 12234
rect 18 12134 50 12166
rect 18 12066 50 12098
rect 18 11998 50 12030
rect 18 11930 50 11962
rect 18 11862 50 11894
rect 18 11794 50 11826
rect 18 11726 50 11758
rect 18 11658 50 11690
rect 18 11590 50 11622
rect 18 11522 50 11554
rect 18 11454 50 11486
rect 18 11386 50 11418
rect 18 11318 50 11350
rect 18 11250 50 11282
rect 18 11182 50 11214
rect 18 11114 50 11146
rect 18 11046 50 11078
rect 18 10978 50 11010
rect 18 10910 50 10942
rect 18 10842 50 10874
rect 18 10774 50 10806
rect 18 10706 50 10738
rect 18 10638 50 10670
rect 18 10570 50 10602
rect 18 10502 50 10534
rect 18 10434 50 10466
rect 18 10366 50 10398
rect 18 10298 50 10330
rect 18 10230 50 10262
rect 18 10162 50 10194
rect 18 10094 50 10126
rect 18 10026 50 10058
rect 18 9958 50 9990
rect 18 9890 50 9922
rect 18 9822 50 9854
rect 18 9754 50 9786
rect 18 9686 50 9718
rect 18 9618 50 9650
rect 18 9550 50 9582
rect 18 9482 50 9514
rect 18 9414 50 9446
rect 18 9346 50 9378
rect 18 9278 50 9310
rect 18 9210 50 9242
rect 18 9142 50 9174
rect 18 9074 50 9106
rect 18 9006 50 9038
rect 18 8938 50 8970
rect 18 8870 50 8902
rect 18 8802 50 8834
rect 18 8734 50 8766
rect 18 8666 50 8698
rect 18 8598 50 8630
rect 18 8530 50 8562
rect 18 8462 50 8494
rect 18 8394 50 8426
rect 18 8326 50 8358
rect 18 8258 50 8290
rect 18 8190 50 8222
rect 18 8122 50 8154
rect 18 8054 50 8086
rect 18 7986 50 8018
rect 18 7918 50 7950
rect 18 7850 50 7882
rect 18 7782 50 7814
rect 18 7714 50 7746
rect 18 7646 50 7678
rect 18 7578 50 7610
rect 18 7510 50 7542
rect 18 7442 50 7474
rect 18 7374 50 7406
rect 18 7306 50 7338
rect 18 7238 50 7270
rect 18 7170 50 7202
rect 18 7102 50 7134
rect 18 7034 50 7066
rect 18 6966 50 6998
rect 18 6898 50 6930
rect 18 6830 50 6862
rect 18 6762 50 6794
rect 18 6694 50 6726
rect 18 6626 50 6658
rect 18 6558 50 6590
rect 18 6490 50 6522
rect 18 6422 50 6454
rect 18 6354 50 6386
rect 18 6286 50 6318
rect 18 6218 50 6250
rect 15950 12474 15982 12506
rect 15950 12406 15982 12438
rect 15950 12338 15982 12370
rect 15950 12270 15982 12302
rect 15950 12202 15982 12234
rect 15950 12134 15982 12166
rect 15950 12066 15982 12098
rect 15950 11998 15982 12030
rect 15950 11930 15982 11962
rect 15950 11862 15982 11894
rect 15950 11794 15982 11826
rect 15950 11726 15982 11758
rect 15950 11658 15982 11690
rect 15950 11590 15982 11622
rect 15950 11522 15982 11554
rect 15950 11454 15982 11486
rect 15950 11386 15982 11418
rect 15950 11318 15982 11350
rect 15950 11250 15982 11282
rect 15950 11182 15982 11214
rect 15950 11114 15982 11146
rect 15950 11046 15982 11078
rect 15950 10978 15982 11010
rect 15950 10910 15982 10942
rect 15950 10842 15982 10874
rect 15950 10774 15982 10806
rect 15950 10706 15982 10738
rect 15950 10638 15982 10670
rect 15950 10570 15982 10602
rect 15950 10502 15982 10534
rect 15950 10434 15982 10466
rect 15950 10366 15982 10398
rect 15950 10298 15982 10330
rect 15950 10230 15982 10262
rect 15950 10162 15982 10194
rect 15950 10094 15982 10126
rect 15950 10026 15982 10058
rect 15950 9958 15982 9990
rect 15950 9890 15982 9922
rect 15950 9822 15982 9854
rect 15950 9754 15982 9786
rect 15950 9686 15982 9718
rect 15950 9618 15982 9650
rect 15950 9550 15982 9582
rect 15950 9482 15982 9514
rect 15950 9414 15982 9446
rect 15950 9346 15982 9378
rect 15950 9278 15982 9310
rect 15950 9210 15982 9242
rect 15950 9142 15982 9174
rect 15950 9074 15982 9106
rect 15950 9006 15982 9038
rect 15950 8938 15982 8970
rect 15950 8870 15982 8902
rect 15950 8802 15982 8834
rect 15950 8734 15982 8766
rect 15950 8666 15982 8698
rect 15950 8598 15982 8630
rect 15950 8530 15982 8562
rect 15950 8462 15982 8494
rect 15950 8394 15982 8426
rect 15950 8326 15982 8358
rect 15950 8258 15982 8290
rect 15950 8190 15982 8222
rect 15950 8122 15982 8154
rect 15950 8054 15982 8086
rect 15950 7986 15982 8018
rect 15950 7918 15982 7950
rect 15950 7850 15982 7882
rect 15950 7782 15982 7814
rect 15950 7714 15982 7746
rect 15950 7646 15982 7678
rect 15950 7578 15982 7610
rect 15950 7510 15982 7542
rect 15950 7442 15982 7474
rect 15950 7374 15982 7406
rect 15950 7306 15982 7338
rect 15950 7238 15982 7270
rect 15950 7170 15982 7202
rect 15950 7102 15982 7134
rect 15950 7034 15982 7066
rect 15950 6966 15982 6998
rect 15950 6898 15982 6930
rect 15950 6830 15982 6862
rect 15950 6762 15982 6794
rect 15950 6694 15982 6726
rect 15950 6626 15982 6658
rect 15950 6558 15982 6590
rect 15950 6490 15982 6522
rect 15950 6422 15982 6454
rect 15950 6354 15982 6386
rect 15950 6286 15982 6318
rect 15950 6218 15982 6250
rect 96 6102 128 6134
rect 164 6102 196 6134
rect 232 6102 264 6134
rect 300 6102 332 6134
rect 368 6102 400 6134
rect 436 6102 468 6134
rect 504 6102 536 6134
rect 572 6102 604 6134
rect 640 6102 672 6134
rect 708 6102 740 6134
rect 776 6102 808 6134
rect 844 6102 876 6134
rect 912 6102 944 6134
rect 980 6102 1012 6134
rect 1048 6102 1080 6134
rect 1116 6102 1148 6134
rect 1184 6102 1216 6134
rect 1252 6102 1284 6134
rect 1320 6102 1352 6134
rect 1388 6102 1420 6134
rect 1456 6102 1488 6134
rect 1524 6102 1556 6134
rect 1592 6102 1624 6134
rect 1660 6102 1692 6134
rect 1728 6102 1760 6134
rect 1796 6102 1828 6134
rect 1864 6102 1896 6134
rect 1932 6102 1964 6134
rect 2000 6102 2032 6134
rect 2068 6102 2100 6134
rect 2136 6102 2168 6134
rect 2204 6102 2236 6134
rect 2272 6102 2304 6134
rect 2340 6102 2372 6134
rect 2408 6102 2440 6134
rect 2476 6102 2508 6134
rect 2544 6102 2576 6134
rect 2612 6102 2644 6134
rect 2680 6102 2712 6134
rect 2748 6102 2780 6134
rect 2816 6102 2848 6134
rect 2884 6102 2916 6134
rect 2952 6102 2984 6134
rect 3020 6102 3052 6134
rect 3088 6102 3120 6134
rect 3156 6102 3188 6134
rect 3224 6102 3256 6134
rect 3292 6102 3324 6134
rect 3360 6102 3392 6134
rect 3428 6102 3460 6134
rect 3496 6102 3528 6134
rect 3564 6102 3596 6134
rect 3632 6102 3664 6134
rect 3700 6102 3732 6134
rect 3768 6102 3800 6134
rect 3836 6102 3868 6134
rect 3904 6102 3936 6134
rect 3972 6102 4004 6134
rect 4040 6102 4072 6134
rect 4108 6102 4140 6134
rect 4176 6102 4208 6134
rect 4244 6102 4276 6134
rect 4312 6102 4344 6134
rect 4380 6102 4412 6134
rect 4448 6102 4480 6134
rect 4516 6102 4548 6134
rect 4584 6102 4616 6134
rect 4652 6102 4684 6134
rect 4720 6102 4752 6134
rect 4788 6102 4820 6134
rect 4856 6102 4888 6134
rect 4924 6102 4956 6134
rect 4992 6102 5024 6134
rect 5060 6102 5092 6134
rect 5128 6102 5160 6134
rect 5196 6102 5228 6134
rect 5264 6102 5296 6134
rect 5332 6102 5364 6134
rect 5400 6102 5432 6134
rect 5468 6102 5500 6134
rect 5536 6102 5568 6134
rect 5604 6102 5636 6134
rect 5672 6102 5704 6134
rect 5740 6102 5772 6134
rect 5808 6102 5840 6134
rect 5876 6102 5908 6134
rect 5944 6102 5976 6134
rect 6012 6102 6044 6134
rect 6080 6102 6112 6134
rect 6148 6102 6180 6134
rect 6216 6102 6248 6134
rect 6284 6102 6316 6134
rect 6352 6102 6384 6134
rect 6420 6102 6452 6134
rect 6488 6102 6520 6134
rect 6556 6102 6588 6134
rect 6624 6102 6656 6134
rect 6692 6102 6724 6134
rect 6760 6102 6792 6134
rect 6828 6102 6860 6134
rect 6896 6102 6928 6134
rect 6964 6102 6996 6134
rect 7032 6102 7064 6134
rect 7100 6102 7132 6134
rect 7168 6102 7200 6134
rect 7236 6102 7268 6134
rect 7304 6102 7336 6134
rect 7372 6102 7404 6134
rect 7440 6102 7472 6134
rect 7508 6102 7540 6134
rect 7576 6102 7608 6134
rect 7644 6102 7676 6134
rect 7712 6102 7744 6134
rect 7780 6102 7812 6134
rect 7848 6102 7880 6134
rect 7916 6102 7948 6134
rect 7984 6102 8016 6134
rect 8052 6102 8084 6134
rect 8120 6102 8152 6134
rect 8188 6102 8220 6134
rect 8256 6102 8288 6134
rect 8324 6102 8356 6134
rect 8392 6102 8424 6134
rect 8460 6102 8492 6134
rect 8528 6102 8560 6134
rect 8596 6102 8628 6134
rect 8664 6102 8696 6134
rect 8732 6102 8764 6134
rect 8800 6102 8832 6134
rect 8868 6102 8900 6134
rect 8936 6102 8968 6134
rect 9004 6102 9036 6134
rect 9072 6102 9104 6134
rect 9140 6102 9172 6134
rect 9208 6102 9240 6134
rect 9276 6102 9308 6134
rect 9344 6102 9376 6134
rect 9412 6102 9444 6134
rect 9480 6102 9512 6134
rect 9548 6102 9580 6134
rect 9616 6102 9648 6134
rect 9684 6102 9716 6134
rect 9752 6102 9784 6134
rect 9820 6102 9852 6134
rect 9888 6102 9920 6134
rect 9956 6102 9988 6134
rect 10024 6102 10056 6134
rect 10092 6102 10124 6134
rect 10160 6102 10192 6134
rect 10228 6102 10260 6134
rect 10296 6102 10328 6134
rect 10364 6102 10396 6134
rect 10432 6102 10464 6134
rect 10500 6102 10532 6134
rect 10568 6102 10600 6134
rect 10636 6102 10668 6134
rect 10704 6102 10736 6134
rect 10772 6102 10804 6134
rect 10840 6102 10872 6134
rect 10908 6102 10940 6134
rect 10976 6102 11008 6134
rect 11044 6102 11076 6134
rect 11112 6102 11144 6134
rect 11180 6102 11212 6134
rect 11248 6102 11280 6134
rect 11316 6102 11348 6134
rect 11384 6102 11416 6134
rect 11452 6102 11484 6134
rect 11520 6102 11552 6134
rect 11588 6102 11620 6134
rect 11656 6102 11688 6134
rect 11724 6102 11756 6134
rect 11792 6102 11824 6134
rect 11860 6102 11892 6134
rect 11928 6102 11960 6134
rect 11996 6102 12028 6134
rect 12064 6102 12096 6134
rect 12132 6102 12164 6134
rect 12200 6102 12232 6134
rect 12268 6102 12300 6134
rect 12336 6102 12368 6134
rect 12404 6102 12436 6134
rect 12472 6102 12504 6134
rect 12540 6102 12572 6134
rect 12608 6102 12640 6134
rect 12676 6102 12708 6134
rect 12744 6102 12776 6134
rect 12812 6102 12844 6134
rect 12880 6102 12912 6134
rect 12948 6102 12980 6134
rect 13016 6102 13048 6134
rect 13084 6102 13116 6134
rect 13152 6102 13184 6134
rect 13220 6102 13252 6134
rect 13288 6102 13320 6134
rect 13356 6102 13388 6134
rect 13424 6102 13456 6134
rect 13492 6102 13524 6134
rect 13560 6102 13592 6134
rect 13628 6102 13660 6134
rect 13696 6102 13728 6134
rect 13764 6102 13796 6134
rect 13832 6102 13864 6134
rect 13900 6102 13932 6134
rect 13968 6102 14000 6134
rect 14036 6102 14068 6134
rect 14104 6102 14136 6134
rect 14172 6102 14204 6134
rect 14240 6102 14272 6134
rect 14308 6102 14340 6134
rect 14376 6102 14408 6134
rect 14444 6102 14476 6134
rect 14512 6102 14544 6134
rect 14580 6102 14612 6134
rect 14648 6102 14680 6134
rect 14716 6102 14748 6134
rect 14784 6102 14816 6134
rect 14852 6102 14884 6134
rect 14920 6102 14952 6134
rect 14988 6102 15020 6134
rect 15056 6102 15088 6134
rect 15124 6102 15156 6134
rect 15192 6102 15224 6134
rect 15260 6102 15292 6134
rect 15328 6102 15360 6134
rect 15396 6102 15428 6134
rect 15464 6102 15496 6134
rect 15532 6102 15564 6134
rect 15600 6102 15632 6134
rect 15668 6102 15700 6134
rect 15736 6102 15768 6134
rect 15804 6102 15836 6134
rect 15872 6102 15904 6134
rect 15940 6102 15972 6134
rect 0 33416 16000 33430
rect 0 33384 50 33416
rect 82 33384 118 33416
rect 150 33384 186 33416
rect 218 33384 254 33416
rect 286 33384 322 33416
rect 354 33384 390 33416
rect 422 33384 458 33416
rect 490 33384 526 33416
rect 558 33384 594 33416
rect 626 33384 662 33416
rect 694 33384 730 33416
rect 762 33384 798 33416
rect 830 33384 866 33416
rect 898 33384 934 33416
rect 966 33384 1002 33416
rect 1034 33384 1070 33416
rect 1102 33384 1138 33416
rect 1170 33384 1206 33416
rect 1238 33384 1274 33416
rect 1306 33384 1342 33416
rect 1374 33384 1410 33416
rect 1442 33384 1478 33416
rect 1510 33384 1546 33416
rect 1578 33384 1614 33416
rect 1646 33384 1682 33416
rect 1714 33384 1750 33416
rect 1782 33384 1818 33416
rect 1850 33384 1886 33416
rect 1918 33384 1954 33416
rect 1986 33384 2022 33416
rect 2054 33384 2090 33416
rect 2122 33384 2158 33416
rect 2190 33384 2226 33416
rect 2258 33384 2294 33416
rect 2326 33384 2362 33416
rect 2394 33384 2430 33416
rect 2462 33384 2498 33416
rect 2530 33384 2566 33416
rect 2598 33384 2634 33416
rect 2666 33384 2702 33416
rect 2734 33384 2770 33416
rect 2802 33384 2838 33416
rect 2870 33384 2906 33416
rect 2938 33384 2974 33416
rect 3006 33384 3042 33416
rect 3074 33384 3110 33416
rect 3142 33384 3178 33416
rect 3210 33384 3246 33416
rect 3278 33384 3314 33416
rect 3346 33384 3382 33416
rect 3414 33384 3450 33416
rect 3482 33384 3518 33416
rect 3550 33384 3586 33416
rect 3618 33384 3654 33416
rect 3686 33384 3722 33416
rect 3754 33384 3790 33416
rect 3822 33384 3858 33416
rect 3890 33384 3926 33416
rect 3958 33384 3994 33416
rect 4026 33384 4062 33416
rect 4094 33384 4130 33416
rect 4162 33384 4198 33416
rect 4230 33384 4266 33416
rect 4298 33384 4334 33416
rect 4366 33384 4402 33416
rect 4434 33384 4470 33416
rect 4502 33384 4538 33416
rect 4570 33384 4606 33416
rect 4638 33384 4674 33416
rect 4706 33384 4742 33416
rect 4774 33384 4810 33416
rect 4842 33384 4878 33416
rect 4910 33384 4946 33416
rect 4978 33384 5014 33416
rect 5046 33384 5082 33416
rect 5114 33384 5150 33416
rect 5182 33384 5218 33416
rect 5250 33384 5286 33416
rect 5318 33384 5354 33416
rect 5386 33384 5422 33416
rect 5454 33384 5490 33416
rect 5522 33384 5558 33416
rect 5590 33384 5626 33416
rect 5658 33384 5694 33416
rect 5726 33384 5762 33416
rect 5794 33384 5830 33416
rect 5862 33384 5898 33416
rect 5930 33384 5966 33416
rect 5998 33384 6034 33416
rect 6066 33384 6102 33416
rect 6134 33384 6170 33416
rect 6202 33384 6238 33416
rect 6270 33384 6306 33416
rect 6338 33384 6374 33416
rect 6406 33384 6442 33416
rect 6474 33384 6510 33416
rect 6542 33384 6578 33416
rect 6610 33384 6646 33416
rect 6678 33384 6714 33416
rect 6746 33384 6782 33416
rect 6814 33384 6850 33416
rect 6882 33384 6918 33416
rect 6950 33384 6986 33416
rect 7018 33384 7054 33416
rect 7086 33384 7122 33416
rect 7154 33384 7190 33416
rect 7222 33384 7258 33416
rect 7290 33384 7326 33416
rect 7358 33384 7394 33416
rect 7426 33384 7462 33416
rect 7494 33384 7530 33416
rect 7562 33384 7598 33416
rect 7630 33384 7666 33416
rect 7698 33384 7734 33416
rect 7766 33384 7802 33416
rect 7834 33384 7870 33416
rect 7902 33384 7938 33416
rect 7970 33384 8006 33416
rect 8038 33384 8074 33416
rect 8106 33384 8142 33416
rect 8174 33384 8210 33416
rect 8242 33384 8278 33416
rect 8310 33384 8346 33416
rect 8378 33384 8414 33416
rect 8446 33384 8482 33416
rect 8514 33384 8550 33416
rect 8582 33384 8618 33416
rect 8650 33384 8686 33416
rect 8718 33384 8754 33416
rect 8786 33384 8822 33416
rect 8854 33384 8890 33416
rect 8922 33384 8958 33416
rect 8990 33384 9026 33416
rect 9058 33384 9094 33416
rect 9126 33384 9162 33416
rect 9194 33384 9230 33416
rect 9262 33384 9298 33416
rect 9330 33384 9366 33416
rect 9398 33384 9434 33416
rect 9466 33384 9502 33416
rect 9534 33384 9570 33416
rect 9602 33384 9638 33416
rect 9670 33384 9706 33416
rect 9738 33384 9774 33416
rect 9806 33384 9842 33416
rect 9874 33384 9910 33416
rect 9942 33384 9978 33416
rect 10010 33384 10046 33416
rect 10078 33384 10114 33416
rect 10146 33384 10182 33416
rect 10214 33384 10250 33416
rect 10282 33384 10318 33416
rect 10350 33384 10386 33416
rect 10418 33384 10454 33416
rect 10486 33384 10522 33416
rect 10554 33384 10590 33416
rect 10622 33384 10658 33416
rect 10690 33384 10726 33416
rect 10758 33384 10794 33416
rect 10826 33384 10862 33416
rect 10894 33384 10930 33416
rect 10962 33384 10998 33416
rect 11030 33384 11066 33416
rect 11098 33384 11134 33416
rect 11166 33384 11202 33416
rect 11234 33384 11270 33416
rect 11302 33384 11338 33416
rect 11370 33384 11406 33416
rect 11438 33384 11474 33416
rect 11506 33384 11542 33416
rect 11574 33384 11610 33416
rect 11642 33384 11678 33416
rect 11710 33384 11746 33416
rect 11778 33384 11814 33416
rect 11846 33384 11882 33416
rect 11914 33384 11950 33416
rect 11982 33384 12018 33416
rect 12050 33384 12086 33416
rect 12118 33384 12154 33416
rect 12186 33384 12222 33416
rect 12254 33384 12290 33416
rect 12322 33384 12358 33416
rect 12390 33384 12426 33416
rect 12458 33384 12494 33416
rect 12526 33384 12562 33416
rect 12594 33384 12630 33416
rect 12662 33384 12698 33416
rect 12730 33384 12766 33416
rect 12798 33384 12834 33416
rect 12866 33384 12902 33416
rect 12934 33384 12970 33416
rect 13002 33384 13038 33416
rect 13070 33384 13106 33416
rect 13138 33384 13174 33416
rect 13206 33384 13242 33416
rect 13274 33384 13310 33416
rect 13342 33384 13378 33416
rect 13410 33384 13446 33416
rect 13478 33384 13514 33416
rect 13546 33384 13582 33416
rect 13614 33384 13650 33416
rect 13682 33384 13718 33416
rect 13750 33384 13786 33416
rect 13818 33384 13854 33416
rect 13886 33384 13922 33416
rect 13954 33384 13990 33416
rect 14022 33384 14058 33416
rect 14090 33384 14126 33416
rect 14158 33384 14194 33416
rect 14226 33384 14262 33416
rect 14294 33384 14330 33416
rect 14362 33384 14398 33416
rect 14430 33384 14466 33416
rect 14498 33384 14534 33416
rect 14566 33384 14602 33416
rect 14634 33384 14670 33416
rect 14702 33384 14738 33416
rect 14770 33384 14806 33416
rect 14838 33384 14874 33416
rect 14906 33384 14942 33416
rect 14974 33384 15010 33416
rect 15042 33384 15078 33416
rect 15110 33384 15146 33416
rect 15178 33384 15214 33416
rect 15246 33384 15282 33416
rect 15314 33384 15350 33416
rect 15382 33384 15442 33416
rect 15474 33384 15510 33416
rect 15542 33384 15578 33416
rect 15610 33384 15646 33416
rect 15678 33384 15714 33416
rect 15746 33384 15782 33416
rect 15814 33384 15850 33416
rect 15882 33384 15918 33416
rect 15950 33384 16000 33416
rect 0 33370 16000 33384
rect 0 29716 16000 29730
rect 0 29684 50 29716
rect 82 29684 118 29716
rect 150 29684 186 29716
rect 218 29684 254 29716
rect 286 29684 322 29716
rect 354 29684 390 29716
rect 422 29684 458 29716
rect 490 29684 526 29716
rect 558 29684 594 29716
rect 626 29684 662 29716
rect 694 29684 730 29716
rect 762 29684 798 29716
rect 830 29684 866 29716
rect 898 29684 934 29716
rect 966 29684 1002 29716
rect 1034 29684 1070 29716
rect 1102 29684 1138 29716
rect 1170 29684 1206 29716
rect 1238 29684 1274 29716
rect 1306 29684 1342 29716
rect 1374 29684 1410 29716
rect 1442 29684 1478 29716
rect 1510 29684 1546 29716
rect 1578 29684 1614 29716
rect 1646 29684 1682 29716
rect 1714 29684 1750 29716
rect 1782 29684 1818 29716
rect 1850 29684 1886 29716
rect 1918 29684 1954 29716
rect 1986 29684 2022 29716
rect 2054 29684 2090 29716
rect 2122 29684 2158 29716
rect 2190 29684 2226 29716
rect 2258 29684 2294 29716
rect 2326 29684 2362 29716
rect 2394 29684 2430 29716
rect 2462 29684 2498 29716
rect 2530 29684 2566 29716
rect 2598 29684 2634 29716
rect 2666 29684 2702 29716
rect 2734 29684 2770 29716
rect 2802 29684 2838 29716
rect 2870 29684 2906 29716
rect 2938 29684 2974 29716
rect 3006 29684 3042 29716
rect 3074 29684 3110 29716
rect 3142 29684 3178 29716
rect 3210 29684 3246 29716
rect 3278 29684 3314 29716
rect 3346 29684 3382 29716
rect 3414 29684 3450 29716
rect 3482 29684 3518 29716
rect 3550 29684 3586 29716
rect 3618 29684 3654 29716
rect 3686 29684 3722 29716
rect 3754 29684 3790 29716
rect 3822 29684 3858 29716
rect 3890 29684 3926 29716
rect 3958 29684 3994 29716
rect 4026 29684 4062 29716
rect 4094 29684 4130 29716
rect 4162 29684 4198 29716
rect 4230 29684 4266 29716
rect 4298 29684 4334 29716
rect 4366 29684 4402 29716
rect 4434 29684 4470 29716
rect 4502 29684 4538 29716
rect 4570 29684 4606 29716
rect 4638 29684 4674 29716
rect 4706 29684 4742 29716
rect 4774 29684 4810 29716
rect 4842 29684 4878 29716
rect 4910 29684 4946 29716
rect 4978 29684 5014 29716
rect 5046 29684 5082 29716
rect 5114 29684 5150 29716
rect 5182 29684 5218 29716
rect 5250 29684 5286 29716
rect 5318 29684 5354 29716
rect 5386 29684 5422 29716
rect 5454 29684 5490 29716
rect 5522 29684 5558 29716
rect 5590 29684 5626 29716
rect 5658 29684 5694 29716
rect 5726 29684 5762 29716
rect 5794 29684 5830 29716
rect 5862 29684 5898 29716
rect 5930 29684 5966 29716
rect 5998 29684 6034 29716
rect 6066 29684 6102 29716
rect 6134 29684 6170 29716
rect 6202 29684 6238 29716
rect 6270 29684 6306 29716
rect 6338 29684 6374 29716
rect 6406 29684 6442 29716
rect 6474 29684 6510 29716
rect 6542 29684 6578 29716
rect 6610 29684 6646 29716
rect 6678 29684 6714 29716
rect 6746 29684 6782 29716
rect 6814 29684 6850 29716
rect 6882 29684 6918 29716
rect 6950 29684 6986 29716
rect 7018 29684 7054 29716
rect 7086 29684 7122 29716
rect 7154 29684 7190 29716
rect 7222 29684 7258 29716
rect 7290 29684 7326 29716
rect 7358 29684 7394 29716
rect 7426 29684 7462 29716
rect 7494 29684 7530 29716
rect 7562 29684 7598 29716
rect 7630 29684 7666 29716
rect 7698 29684 7734 29716
rect 7766 29684 7802 29716
rect 7834 29684 7870 29716
rect 7902 29684 7938 29716
rect 7970 29684 8006 29716
rect 8038 29684 8074 29716
rect 8106 29684 8142 29716
rect 8174 29684 8210 29716
rect 8242 29684 8278 29716
rect 8310 29684 8346 29716
rect 8378 29684 8414 29716
rect 8446 29684 8482 29716
rect 8514 29684 8550 29716
rect 8582 29684 8618 29716
rect 8650 29684 8686 29716
rect 8718 29684 8754 29716
rect 8786 29684 8822 29716
rect 8854 29684 8890 29716
rect 8922 29684 8958 29716
rect 8990 29684 9026 29716
rect 9058 29684 9094 29716
rect 9126 29684 9162 29716
rect 9194 29684 9230 29716
rect 9262 29684 9298 29716
rect 9330 29684 9366 29716
rect 9398 29684 9434 29716
rect 9466 29684 9502 29716
rect 9534 29684 9570 29716
rect 9602 29684 9638 29716
rect 9670 29684 9706 29716
rect 9738 29684 9774 29716
rect 9806 29684 9842 29716
rect 9874 29684 9910 29716
rect 9942 29684 9978 29716
rect 10010 29684 10046 29716
rect 10078 29684 10114 29716
rect 10146 29684 10182 29716
rect 10214 29684 10250 29716
rect 10282 29684 10318 29716
rect 10350 29684 10386 29716
rect 10418 29684 10454 29716
rect 10486 29684 10522 29716
rect 10554 29684 10590 29716
rect 10622 29684 10658 29716
rect 10690 29684 10726 29716
rect 10758 29684 10794 29716
rect 10826 29684 10862 29716
rect 10894 29684 10930 29716
rect 10962 29684 10998 29716
rect 11030 29684 11066 29716
rect 11098 29684 11134 29716
rect 11166 29684 11202 29716
rect 11234 29684 11270 29716
rect 11302 29684 11338 29716
rect 11370 29684 11406 29716
rect 11438 29684 11474 29716
rect 11506 29684 11542 29716
rect 11574 29684 11610 29716
rect 11642 29684 11678 29716
rect 11710 29684 11746 29716
rect 11778 29684 11814 29716
rect 11846 29684 11882 29716
rect 11914 29684 11950 29716
rect 11982 29684 12018 29716
rect 12050 29684 12086 29716
rect 12118 29684 12154 29716
rect 12186 29684 12222 29716
rect 12254 29684 12290 29716
rect 12322 29684 12358 29716
rect 12390 29684 12426 29716
rect 12458 29684 12494 29716
rect 12526 29684 12562 29716
rect 12594 29684 12630 29716
rect 12662 29684 12698 29716
rect 12730 29684 12766 29716
rect 12798 29684 12834 29716
rect 12866 29684 12902 29716
rect 12934 29684 12970 29716
rect 13002 29684 13038 29716
rect 13070 29684 13106 29716
rect 13138 29684 13174 29716
rect 13206 29684 13242 29716
rect 13274 29684 13310 29716
rect 13342 29684 13378 29716
rect 13410 29684 13446 29716
rect 13478 29684 13514 29716
rect 13546 29684 13582 29716
rect 13614 29684 13650 29716
rect 13682 29684 13718 29716
rect 13750 29684 13786 29716
rect 13818 29684 13854 29716
rect 13886 29684 13922 29716
rect 13954 29684 13990 29716
rect 14022 29684 14058 29716
rect 14090 29684 14126 29716
rect 14158 29684 14194 29716
rect 14226 29684 14262 29716
rect 14294 29684 14330 29716
rect 14362 29684 14398 29716
rect 14430 29684 14466 29716
rect 14498 29684 14534 29716
rect 14566 29684 14602 29716
rect 14634 29684 14670 29716
rect 14702 29684 14738 29716
rect 14770 29684 14806 29716
rect 14838 29684 14874 29716
rect 14906 29684 14942 29716
rect 14974 29684 15010 29716
rect 15042 29684 15078 29716
rect 15110 29684 15146 29716
rect 15178 29684 15214 29716
rect 15246 29684 15282 29716
rect 15314 29684 15350 29716
rect 15382 29684 15442 29716
rect 15474 29684 15510 29716
rect 15542 29684 15578 29716
rect 15610 29684 15646 29716
rect 15678 29684 15714 29716
rect 15746 29684 15782 29716
rect 15814 29684 15850 29716
rect 15882 29684 15918 29716
rect 15950 29684 16000 29716
rect 0 29670 16000 29684
rect 0 12690 16000 12708
rect 0 12658 28 12690
rect 60 12658 96 12690
rect 128 12658 164 12690
rect 196 12658 232 12690
rect 264 12658 300 12690
rect 332 12658 368 12690
rect 400 12658 436 12690
rect 468 12658 504 12690
rect 536 12658 572 12690
rect 604 12658 640 12690
rect 672 12658 708 12690
rect 740 12658 776 12690
rect 808 12658 844 12690
rect 876 12658 912 12690
rect 944 12658 980 12690
rect 1012 12658 1048 12690
rect 1080 12658 1116 12690
rect 1148 12658 1184 12690
rect 1216 12658 1252 12690
rect 1284 12658 1320 12690
rect 1352 12658 1388 12690
rect 1420 12658 1456 12690
rect 1488 12658 1524 12690
rect 1556 12658 1592 12690
rect 1624 12658 1660 12690
rect 1692 12658 1728 12690
rect 1760 12658 1796 12690
rect 1828 12658 1864 12690
rect 1896 12658 1932 12690
rect 1964 12658 2000 12690
rect 2032 12658 2068 12690
rect 2100 12658 2136 12690
rect 2168 12658 2204 12690
rect 2236 12658 2272 12690
rect 2304 12658 2340 12690
rect 2372 12658 2408 12690
rect 2440 12658 2476 12690
rect 2508 12658 2544 12690
rect 2576 12658 2612 12690
rect 2644 12658 2680 12690
rect 2712 12658 2748 12690
rect 2780 12658 2816 12690
rect 2848 12658 2884 12690
rect 2916 12658 2952 12690
rect 2984 12658 3020 12690
rect 3052 12658 3088 12690
rect 3120 12658 3156 12690
rect 3188 12658 3224 12690
rect 3256 12658 3292 12690
rect 3324 12658 3360 12690
rect 3392 12658 3428 12690
rect 3460 12658 3496 12690
rect 3528 12658 3564 12690
rect 3596 12658 3632 12690
rect 3664 12658 3700 12690
rect 3732 12658 3768 12690
rect 3800 12658 3836 12690
rect 3868 12658 3904 12690
rect 3936 12658 3972 12690
rect 4004 12658 4040 12690
rect 4072 12658 4108 12690
rect 4140 12658 4176 12690
rect 4208 12658 4244 12690
rect 4276 12658 4312 12690
rect 4344 12658 4380 12690
rect 4412 12658 4448 12690
rect 4480 12658 4516 12690
rect 4548 12658 4584 12690
rect 4616 12658 4652 12690
rect 4684 12658 4720 12690
rect 4752 12658 4788 12690
rect 4820 12658 4856 12690
rect 4888 12658 4924 12690
rect 4956 12658 4992 12690
rect 5024 12658 5060 12690
rect 5092 12658 5128 12690
rect 5160 12658 5196 12690
rect 5228 12658 5264 12690
rect 5296 12658 5332 12690
rect 5364 12658 5400 12690
rect 5432 12658 5468 12690
rect 5500 12658 5536 12690
rect 5568 12658 5604 12690
rect 5636 12658 5672 12690
rect 5704 12658 5740 12690
rect 5772 12658 5808 12690
rect 5840 12658 5876 12690
rect 5908 12658 5944 12690
rect 5976 12658 6012 12690
rect 6044 12658 6080 12690
rect 6112 12658 6148 12690
rect 6180 12658 6216 12690
rect 6248 12658 6284 12690
rect 6316 12658 6352 12690
rect 6384 12658 6420 12690
rect 6452 12658 6488 12690
rect 6520 12658 6556 12690
rect 6588 12658 6624 12690
rect 6656 12658 6692 12690
rect 6724 12658 6760 12690
rect 6792 12658 6828 12690
rect 6860 12658 6896 12690
rect 6928 12658 6964 12690
rect 6996 12658 7032 12690
rect 7064 12658 7100 12690
rect 7132 12658 7168 12690
rect 7200 12658 7236 12690
rect 7268 12658 7304 12690
rect 7336 12658 7372 12690
rect 7404 12658 7440 12690
rect 7472 12658 7508 12690
rect 7540 12658 7576 12690
rect 7608 12658 7644 12690
rect 7676 12658 7712 12690
rect 7744 12658 7780 12690
rect 7812 12658 7848 12690
rect 7880 12658 7916 12690
rect 7948 12658 7984 12690
rect 8016 12658 8052 12690
rect 8084 12658 8120 12690
rect 8152 12658 8188 12690
rect 8220 12658 8256 12690
rect 8288 12658 8324 12690
rect 8356 12658 8392 12690
rect 8424 12658 8460 12690
rect 8492 12658 8528 12690
rect 8560 12658 8596 12690
rect 8628 12658 8664 12690
rect 8696 12658 8732 12690
rect 8764 12658 8800 12690
rect 8832 12658 8868 12690
rect 8900 12658 8936 12690
rect 8968 12658 9004 12690
rect 9036 12658 9072 12690
rect 9104 12658 9140 12690
rect 9172 12658 9208 12690
rect 9240 12658 9276 12690
rect 9308 12658 9344 12690
rect 9376 12658 9412 12690
rect 9444 12658 9480 12690
rect 9512 12658 9548 12690
rect 9580 12658 9616 12690
rect 9648 12658 9684 12690
rect 9716 12658 9752 12690
rect 9784 12658 9820 12690
rect 9852 12658 9888 12690
rect 9920 12658 9956 12690
rect 9988 12658 10024 12690
rect 10056 12658 10092 12690
rect 10124 12658 10160 12690
rect 10192 12658 10228 12690
rect 10260 12658 10296 12690
rect 10328 12658 10364 12690
rect 10396 12658 10432 12690
rect 10464 12658 10500 12690
rect 10532 12658 10568 12690
rect 10600 12658 10636 12690
rect 10668 12658 10704 12690
rect 10736 12658 10772 12690
rect 10804 12658 10840 12690
rect 10872 12658 10908 12690
rect 10940 12658 10976 12690
rect 11008 12658 11044 12690
rect 11076 12658 11112 12690
rect 11144 12658 11180 12690
rect 11212 12658 11248 12690
rect 11280 12658 11316 12690
rect 11348 12658 11384 12690
rect 11416 12658 11452 12690
rect 11484 12658 11520 12690
rect 11552 12658 11588 12690
rect 11620 12658 11656 12690
rect 11688 12658 11724 12690
rect 11756 12658 11792 12690
rect 11824 12658 11860 12690
rect 11892 12658 11928 12690
rect 11960 12658 11996 12690
rect 12028 12658 12064 12690
rect 12096 12658 12132 12690
rect 12164 12658 12200 12690
rect 12232 12658 12268 12690
rect 12300 12658 12336 12690
rect 12368 12658 12404 12690
rect 12436 12658 12472 12690
rect 12504 12658 12540 12690
rect 12572 12658 12608 12690
rect 12640 12658 12676 12690
rect 12708 12658 12744 12690
rect 12776 12658 12812 12690
rect 12844 12658 12880 12690
rect 12912 12658 12948 12690
rect 12980 12658 13016 12690
rect 13048 12658 13084 12690
rect 13116 12658 13152 12690
rect 13184 12658 13220 12690
rect 13252 12658 13288 12690
rect 13320 12658 13356 12690
rect 13388 12658 13424 12690
rect 13456 12658 13492 12690
rect 13524 12658 13560 12690
rect 13592 12658 13628 12690
rect 13660 12658 13696 12690
rect 13728 12658 13764 12690
rect 13796 12658 13832 12690
rect 13864 12658 13900 12690
rect 13932 12658 13968 12690
rect 14000 12658 14036 12690
rect 14068 12658 14104 12690
rect 14136 12658 14172 12690
rect 14204 12658 14240 12690
rect 14272 12658 14308 12690
rect 14340 12658 14376 12690
rect 14408 12658 14444 12690
rect 14476 12658 14512 12690
rect 14544 12658 14580 12690
rect 14612 12658 14648 12690
rect 14680 12658 14716 12690
rect 14748 12658 14784 12690
rect 14816 12658 14852 12690
rect 14884 12658 14920 12690
rect 14952 12658 14988 12690
rect 15020 12658 15056 12690
rect 15088 12658 15124 12690
rect 15156 12658 15192 12690
rect 15224 12658 15260 12690
rect 15292 12658 15328 12690
rect 15360 12658 15396 12690
rect 15428 12658 15464 12690
rect 15496 12658 15532 12690
rect 15564 12658 15600 12690
rect 15632 12658 15668 12690
rect 15700 12658 15736 12690
rect 15768 12658 15804 12690
rect 15836 12658 15872 12690
rect 15904 12658 15940 12690
rect 15972 12658 16000 12690
rect 0 12640 16000 12658
rect 0 12574 68 12640
rect 0 12542 18 12574
rect 50 12542 68 12574
rect 0 12506 68 12542
rect 0 12474 18 12506
rect 50 12474 68 12506
rect 0 12438 68 12474
rect 0 12406 18 12438
rect 50 12406 68 12438
rect 0 12370 68 12406
rect 0 12338 18 12370
rect 50 12338 68 12370
rect 0 12302 68 12338
rect 0 12270 18 12302
rect 50 12270 68 12302
rect 0 12234 68 12270
rect 0 12202 18 12234
rect 50 12202 68 12234
rect 0 12166 68 12202
rect 0 12134 18 12166
rect 50 12134 68 12166
rect 0 12098 68 12134
rect 0 12066 18 12098
rect 50 12066 68 12098
rect 0 12030 68 12066
rect 0 11998 18 12030
rect 50 11998 68 12030
rect 0 11962 68 11998
rect 0 11930 18 11962
rect 50 11930 68 11962
rect 0 11894 68 11930
rect 0 11862 18 11894
rect 50 11862 68 11894
rect 0 11826 68 11862
rect 0 11794 18 11826
rect 50 11794 68 11826
rect 0 11758 68 11794
rect 0 11726 18 11758
rect 50 11726 68 11758
rect 0 11690 68 11726
rect 0 11658 18 11690
rect 50 11658 68 11690
rect 0 11622 68 11658
rect 0 11590 18 11622
rect 50 11590 68 11622
rect 0 11554 68 11590
rect 0 11522 18 11554
rect 50 11522 68 11554
rect 0 11486 68 11522
rect 0 11454 18 11486
rect 50 11454 68 11486
rect 0 11418 68 11454
rect 0 11386 18 11418
rect 50 11386 68 11418
rect 0 11350 68 11386
rect 0 11318 18 11350
rect 50 11318 68 11350
rect 0 11282 68 11318
rect 0 11250 18 11282
rect 50 11250 68 11282
rect 0 11214 68 11250
rect 0 11182 18 11214
rect 50 11182 68 11214
rect 0 11146 68 11182
rect 0 11114 18 11146
rect 50 11114 68 11146
rect 0 11078 68 11114
rect 0 11046 18 11078
rect 50 11046 68 11078
rect 0 11010 68 11046
rect 0 10978 18 11010
rect 50 10978 68 11010
rect 0 10942 68 10978
rect 0 10910 18 10942
rect 50 10910 68 10942
rect 0 10874 68 10910
rect 0 10842 18 10874
rect 50 10842 68 10874
rect 0 10806 68 10842
rect 0 10774 18 10806
rect 50 10774 68 10806
rect 0 10738 68 10774
rect 0 10706 18 10738
rect 50 10706 68 10738
rect 0 10670 68 10706
rect 0 10638 18 10670
rect 50 10638 68 10670
rect 0 10602 68 10638
rect 0 10570 18 10602
rect 50 10570 68 10602
rect 0 10534 68 10570
rect 0 10502 18 10534
rect 50 10502 68 10534
rect 0 10466 68 10502
rect 0 10434 18 10466
rect 50 10434 68 10466
rect 0 10398 68 10434
rect 0 10366 18 10398
rect 50 10366 68 10398
rect 0 10330 68 10366
rect 0 10298 18 10330
rect 50 10298 68 10330
rect 0 10262 68 10298
rect 0 10230 18 10262
rect 50 10230 68 10262
rect 0 10194 68 10230
rect 0 10162 18 10194
rect 50 10162 68 10194
rect 0 10126 68 10162
rect 0 10094 18 10126
rect 50 10094 68 10126
rect 0 10058 68 10094
rect 0 10026 18 10058
rect 50 10026 68 10058
rect 0 9990 68 10026
rect 0 9958 18 9990
rect 50 9958 68 9990
rect 0 9922 68 9958
rect 0 9890 18 9922
rect 50 9890 68 9922
rect 0 9854 68 9890
rect 0 9822 18 9854
rect 50 9822 68 9854
rect 0 9786 68 9822
rect 0 9754 18 9786
rect 50 9754 68 9786
rect 0 9718 68 9754
rect 0 9686 18 9718
rect 50 9686 68 9718
rect 0 9650 68 9686
rect 0 9618 18 9650
rect 50 9618 68 9650
rect 0 9582 68 9618
rect 0 9550 18 9582
rect 50 9550 68 9582
rect 0 9514 68 9550
rect 0 9482 18 9514
rect 50 9482 68 9514
rect 0 9446 68 9482
rect 0 9414 18 9446
rect 50 9414 68 9446
rect 0 9378 68 9414
rect 0 9346 18 9378
rect 50 9346 68 9378
rect 0 9310 68 9346
rect 0 9278 18 9310
rect 50 9278 68 9310
rect 0 9242 68 9278
rect 0 9210 18 9242
rect 50 9210 68 9242
rect 0 9174 68 9210
rect 0 9142 18 9174
rect 50 9142 68 9174
rect 0 9106 68 9142
rect 0 9074 18 9106
rect 50 9074 68 9106
rect 0 9038 68 9074
rect 0 9006 18 9038
rect 50 9006 68 9038
rect 0 8970 68 9006
rect 0 8938 18 8970
rect 50 8938 68 8970
rect 0 8902 68 8938
rect 0 8870 18 8902
rect 50 8870 68 8902
rect 0 8834 68 8870
rect 0 8802 18 8834
rect 50 8802 68 8834
rect 0 8766 68 8802
rect 0 8734 18 8766
rect 50 8734 68 8766
rect 0 8698 68 8734
rect 0 8666 18 8698
rect 50 8666 68 8698
rect 0 8630 68 8666
rect 0 8598 18 8630
rect 50 8598 68 8630
rect 0 8562 68 8598
rect 0 8530 18 8562
rect 50 8530 68 8562
rect 0 8494 68 8530
rect 0 8462 18 8494
rect 50 8462 68 8494
rect 0 8426 68 8462
rect 0 8394 18 8426
rect 50 8394 68 8426
rect 0 8358 68 8394
rect 0 8326 18 8358
rect 50 8326 68 8358
rect 0 8290 68 8326
rect 0 8258 18 8290
rect 50 8258 68 8290
rect 0 8222 68 8258
rect 0 8190 18 8222
rect 50 8190 68 8222
rect 0 8154 68 8190
rect 0 8122 18 8154
rect 50 8122 68 8154
rect 0 8086 68 8122
rect 0 8054 18 8086
rect 50 8054 68 8086
rect 0 8018 68 8054
rect 0 7986 18 8018
rect 50 7986 68 8018
rect 0 7950 68 7986
rect 0 7918 18 7950
rect 50 7918 68 7950
rect 0 7882 68 7918
rect 0 7850 18 7882
rect 50 7850 68 7882
rect 0 7814 68 7850
rect 0 7782 18 7814
rect 50 7782 68 7814
rect 0 7746 68 7782
rect 0 7714 18 7746
rect 50 7714 68 7746
rect 0 7678 68 7714
rect 0 7646 18 7678
rect 50 7646 68 7678
rect 0 7610 68 7646
rect 0 7578 18 7610
rect 50 7578 68 7610
rect 0 7542 68 7578
rect 0 7510 18 7542
rect 50 7510 68 7542
rect 0 7474 68 7510
rect 0 7442 18 7474
rect 50 7442 68 7474
rect 0 7406 68 7442
rect 0 7374 18 7406
rect 50 7374 68 7406
rect 0 7338 68 7374
rect 0 7306 18 7338
rect 50 7306 68 7338
rect 0 7270 68 7306
rect 0 7238 18 7270
rect 50 7238 68 7270
rect 0 7202 68 7238
rect 0 7170 18 7202
rect 50 7170 68 7202
rect 0 7134 68 7170
rect 0 7102 18 7134
rect 50 7102 68 7134
rect 0 7066 68 7102
rect 0 7034 18 7066
rect 50 7034 68 7066
rect 0 6998 68 7034
rect 0 6966 18 6998
rect 50 6966 68 6998
rect 0 6930 68 6966
rect 0 6898 18 6930
rect 50 6898 68 6930
rect 0 6862 68 6898
rect 0 6830 18 6862
rect 50 6830 68 6862
rect 0 6794 68 6830
rect 0 6762 18 6794
rect 50 6762 68 6794
rect 0 6726 68 6762
rect 0 6694 18 6726
rect 50 6694 68 6726
rect 0 6658 68 6694
rect 0 6626 18 6658
rect 50 6626 68 6658
rect 0 6590 68 6626
rect 0 6558 18 6590
rect 50 6558 68 6590
rect 0 6522 68 6558
rect 0 6490 18 6522
rect 50 6490 68 6522
rect 0 6454 68 6490
rect 0 6422 18 6454
rect 50 6422 68 6454
rect 0 6386 68 6422
rect 0 6354 18 6386
rect 50 6354 68 6386
rect 0 6318 68 6354
rect 0 6286 18 6318
rect 50 6286 68 6318
rect 0 6250 68 6286
rect 0 6218 18 6250
rect 50 6218 68 6250
rect 0 6152 68 6218
rect 15932 12574 16000 12640
rect 15932 12542 15950 12574
rect 15982 12542 16000 12574
rect 15932 12506 16000 12542
rect 15932 12474 15950 12506
rect 15982 12474 16000 12506
rect 15932 12438 16000 12474
rect 15932 12406 15950 12438
rect 15982 12406 16000 12438
rect 15932 12370 16000 12406
rect 15932 12338 15950 12370
rect 15982 12338 16000 12370
rect 15932 12302 16000 12338
rect 15932 12270 15950 12302
rect 15982 12270 16000 12302
rect 15932 12234 16000 12270
rect 15932 12202 15950 12234
rect 15982 12202 16000 12234
rect 15932 12166 16000 12202
rect 15932 12134 15950 12166
rect 15982 12134 16000 12166
rect 15932 12098 16000 12134
rect 15932 12066 15950 12098
rect 15982 12066 16000 12098
rect 15932 12030 16000 12066
rect 15932 11998 15950 12030
rect 15982 11998 16000 12030
rect 15932 11962 16000 11998
rect 15932 11930 15950 11962
rect 15982 11930 16000 11962
rect 15932 11894 16000 11930
rect 15932 11862 15950 11894
rect 15982 11862 16000 11894
rect 15932 11826 16000 11862
rect 15932 11794 15950 11826
rect 15982 11794 16000 11826
rect 15932 11758 16000 11794
rect 15932 11726 15950 11758
rect 15982 11726 16000 11758
rect 15932 11690 16000 11726
rect 15932 11658 15950 11690
rect 15982 11658 16000 11690
rect 15932 11622 16000 11658
rect 15932 11590 15950 11622
rect 15982 11590 16000 11622
rect 15932 11554 16000 11590
rect 15932 11522 15950 11554
rect 15982 11522 16000 11554
rect 15932 11486 16000 11522
rect 15932 11454 15950 11486
rect 15982 11454 16000 11486
rect 15932 11418 16000 11454
rect 15932 11386 15950 11418
rect 15982 11386 16000 11418
rect 15932 11350 16000 11386
rect 15932 11318 15950 11350
rect 15982 11318 16000 11350
rect 15932 11282 16000 11318
rect 15932 11250 15950 11282
rect 15982 11250 16000 11282
rect 15932 11214 16000 11250
rect 15932 11182 15950 11214
rect 15982 11182 16000 11214
rect 15932 11146 16000 11182
rect 15932 11114 15950 11146
rect 15982 11114 16000 11146
rect 15932 11078 16000 11114
rect 15932 11046 15950 11078
rect 15982 11046 16000 11078
rect 15932 11010 16000 11046
rect 15932 10978 15950 11010
rect 15982 10978 16000 11010
rect 15932 10942 16000 10978
rect 15932 10910 15950 10942
rect 15982 10910 16000 10942
rect 15932 10874 16000 10910
rect 15932 10842 15950 10874
rect 15982 10842 16000 10874
rect 15932 10806 16000 10842
rect 15932 10774 15950 10806
rect 15982 10774 16000 10806
rect 15932 10738 16000 10774
rect 15932 10706 15950 10738
rect 15982 10706 16000 10738
rect 15932 10670 16000 10706
rect 15932 10638 15950 10670
rect 15982 10638 16000 10670
rect 15932 10602 16000 10638
rect 15932 10570 15950 10602
rect 15982 10570 16000 10602
rect 15932 10534 16000 10570
rect 15932 10502 15950 10534
rect 15982 10502 16000 10534
rect 15932 10466 16000 10502
rect 15932 10434 15950 10466
rect 15982 10434 16000 10466
rect 15932 10398 16000 10434
rect 15932 10366 15950 10398
rect 15982 10366 16000 10398
rect 15932 10330 16000 10366
rect 15932 10298 15950 10330
rect 15982 10298 16000 10330
rect 15932 10262 16000 10298
rect 15932 10230 15950 10262
rect 15982 10230 16000 10262
rect 15932 10194 16000 10230
rect 15932 10162 15950 10194
rect 15982 10162 16000 10194
rect 15932 10126 16000 10162
rect 15932 10094 15950 10126
rect 15982 10094 16000 10126
rect 15932 10058 16000 10094
rect 15932 10026 15950 10058
rect 15982 10026 16000 10058
rect 15932 9990 16000 10026
rect 15932 9958 15950 9990
rect 15982 9958 16000 9990
rect 15932 9922 16000 9958
rect 15932 9890 15950 9922
rect 15982 9890 16000 9922
rect 15932 9854 16000 9890
rect 15932 9822 15950 9854
rect 15982 9822 16000 9854
rect 15932 9786 16000 9822
rect 15932 9754 15950 9786
rect 15982 9754 16000 9786
rect 15932 9718 16000 9754
rect 15932 9686 15950 9718
rect 15982 9686 16000 9718
rect 15932 9650 16000 9686
rect 15932 9618 15950 9650
rect 15982 9618 16000 9650
rect 15932 9582 16000 9618
rect 15932 9550 15950 9582
rect 15982 9550 16000 9582
rect 15932 9514 16000 9550
rect 15932 9482 15950 9514
rect 15982 9482 16000 9514
rect 15932 9446 16000 9482
rect 15932 9414 15950 9446
rect 15982 9414 16000 9446
rect 15932 9378 16000 9414
rect 15932 9346 15950 9378
rect 15982 9346 16000 9378
rect 15932 9310 16000 9346
rect 15932 9278 15950 9310
rect 15982 9278 16000 9310
rect 15932 9242 16000 9278
rect 15932 9210 15950 9242
rect 15982 9210 16000 9242
rect 15932 9174 16000 9210
rect 15932 9142 15950 9174
rect 15982 9142 16000 9174
rect 15932 9106 16000 9142
rect 15932 9074 15950 9106
rect 15982 9074 16000 9106
rect 15932 9038 16000 9074
rect 15932 9006 15950 9038
rect 15982 9006 16000 9038
rect 15932 8970 16000 9006
rect 15932 8938 15950 8970
rect 15982 8938 16000 8970
rect 15932 8902 16000 8938
rect 15932 8870 15950 8902
rect 15982 8870 16000 8902
rect 15932 8834 16000 8870
rect 15932 8802 15950 8834
rect 15982 8802 16000 8834
rect 15932 8766 16000 8802
rect 15932 8734 15950 8766
rect 15982 8734 16000 8766
rect 15932 8698 16000 8734
rect 15932 8666 15950 8698
rect 15982 8666 16000 8698
rect 15932 8630 16000 8666
rect 15932 8598 15950 8630
rect 15982 8598 16000 8630
rect 15932 8562 16000 8598
rect 15932 8530 15950 8562
rect 15982 8530 16000 8562
rect 15932 8494 16000 8530
rect 15932 8462 15950 8494
rect 15982 8462 16000 8494
rect 15932 8426 16000 8462
rect 15932 8394 15950 8426
rect 15982 8394 16000 8426
rect 15932 8358 16000 8394
rect 15932 8326 15950 8358
rect 15982 8326 16000 8358
rect 15932 8290 16000 8326
rect 15932 8258 15950 8290
rect 15982 8258 16000 8290
rect 15932 8222 16000 8258
rect 15932 8190 15950 8222
rect 15982 8190 16000 8222
rect 15932 8154 16000 8190
rect 15932 8122 15950 8154
rect 15982 8122 16000 8154
rect 15932 8086 16000 8122
rect 15932 8054 15950 8086
rect 15982 8054 16000 8086
rect 15932 8018 16000 8054
rect 15932 7986 15950 8018
rect 15982 7986 16000 8018
rect 15932 7950 16000 7986
rect 15932 7918 15950 7950
rect 15982 7918 16000 7950
rect 15932 7882 16000 7918
rect 15932 7850 15950 7882
rect 15982 7850 16000 7882
rect 15932 7814 16000 7850
rect 15932 7782 15950 7814
rect 15982 7782 16000 7814
rect 15932 7746 16000 7782
rect 15932 7714 15950 7746
rect 15982 7714 16000 7746
rect 15932 7678 16000 7714
rect 15932 7646 15950 7678
rect 15982 7646 16000 7678
rect 15932 7610 16000 7646
rect 15932 7578 15950 7610
rect 15982 7578 16000 7610
rect 15932 7542 16000 7578
rect 15932 7510 15950 7542
rect 15982 7510 16000 7542
rect 15932 7474 16000 7510
rect 15932 7442 15950 7474
rect 15982 7442 16000 7474
rect 15932 7406 16000 7442
rect 15932 7374 15950 7406
rect 15982 7374 16000 7406
rect 15932 7338 16000 7374
rect 15932 7306 15950 7338
rect 15982 7306 16000 7338
rect 15932 7270 16000 7306
rect 15932 7238 15950 7270
rect 15982 7238 16000 7270
rect 15932 7202 16000 7238
rect 15932 7170 15950 7202
rect 15982 7170 16000 7202
rect 15932 7134 16000 7170
rect 15932 7102 15950 7134
rect 15982 7102 16000 7134
rect 15932 7066 16000 7102
rect 15932 7034 15950 7066
rect 15982 7034 16000 7066
rect 15932 6998 16000 7034
rect 15932 6966 15950 6998
rect 15982 6966 16000 6998
rect 15932 6930 16000 6966
rect 15932 6898 15950 6930
rect 15982 6898 16000 6930
rect 15932 6862 16000 6898
rect 15932 6830 15950 6862
rect 15982 6830 16000 6862
rect 15932 6794 16000 6830
rect 15932 6762 15950 6794
rect 15982 6762 16000 6794
rect 15932 6726 16000 6762
rect 15932 6694 15950 6726
rect 15982 6694 16000 6726
rect 15932 6658 16000 6694
rect 15932 6626 15950 6658
rect 15982 6626 16000 6658
rect 15932 6590 16000 6626
rect 15932 6558 15950 6590
rect 15982 6558 16000 6590
rect 15932 6522 16000 6558
rect 15932 6490 15950 6522
rect 15982 6490 16000 6522
rect 15932 6454 16000 6490
rect 15932 6422 15950 6454
rect 15982 6422 16000 6454
rect 15932 6386 16000 6422
rect 15932 6354 15950 6386
rect 15982 6354 16000 6386
rect 15932 6318 16000 6354
rect 15932 6286 15950 6318
rect 15982 6286 16000 6318
rect 15932 6250 16000 6286
rect 15932 6218 15950 6250
rect 15982 6218 16000 6250
rect 15932 6152 16000 6218
rect 0 6134 16000 6152
rect 0 6102 28 6134
rect 60 6102 96 6134
rect 128 6102 164 6134
rect 196 6102 232 6134
rect 264 6102 300 6134
rect 332 6102 368 6134
rect 400 6102 436 6134
rect 468 6102 504 6134
rect 536 6102 572 6134
rect 604 6102 640 6134
rect 672 6102 708 6134
rect 740 6102 776 6134
rect 808 6102 844 6134
rect 876 6102 912 6134
rect 944 6102 980 6134
rect 1012 6102 1048 6134
rect 1080 6102 1116 6134
rect 1148 6102 1184 6134
rect 1216 6102 1252 6134
rect 1284 6102 1320 6134
rect 1352 6102 1388 6134
rect 1420 6102 1456 6134
rect 1488 6102 1524 6134
rect 1556 6102 1592 6134
rect 1624 6102 1660 6134
rect 1692 6102 1728 6134
rect 1760 6102 1796 6134
rect 1828 6102 1864 6134
rect 1896 6102 1932 6134
rect 1964 6102 2000 6134
rect 2032 6102 2068 6134
rect 2100 6102 2136 6134
rect 2168 6102 2204 6134
rect 2236 6102 2272 6134
rect 2304 6102 2340 6134
rect 2372 6102 2408 6134
rect 2440 6102 2476 6134
rect 2508 6102 2544 6134
rect 2576 6102 2612 6134
rect 2644 6102 2680 6134
rect 2712 6102 2748 6134
rect 2780 6102 2816 6134
rect 2848 6102 2884 6134
rect 2916 6102 2952 6134
rect 2984 6102 3020 6134
rect 3052 6102 3088 6134
rect 3120 6102 3156 6134
rect 3188 6102 3224 6134
rect 3256 6102 3292 6134
rect 3324 6102 3360 6134
rect 3392 6102 3428 6134
rect 3460 6102 3496 6134
rect 3528 6102 3564 6134
rect 3596 6102 3632 6134
rect 3664 6102 3700 6134
rect 3732 6102 3768 6134
rect 3800 6102 3836 6134
rect 3868 6102 3904 6134
rect 3936 6102 3972 6134
rect 4004 6102 4040 6134
rect 4072 6102 4108 6134
rect 4140 6102 4176 6134
rect 4208 6102 4244 6134
rect 4276 6102 4312 6134
rect 4344 6102 4380 6134
rect 4412 6102 4448 6134
rect 4480 6102 4516 6134
rect 4548 6102 4584 6134
rect 4616 6102 4652 6134
rect 4684 6102 4720 6134
rect 4752 6102 4788 6134
rect 4820 6102 4856 6134
rect 4888 6102 4924 6134
rect 4956 6102 4992 6134
rect 5024 6102 5060 6134
rect 5092 6102 5128 6134
rect 5160 6102 5196 6134
rect 5228 6102 5264 6134
rect 5296 6102 5332 6134
rect 5364 6102 5400 6134
rect 5432 6102 5468 6134
rect 5500 6102 5536 6134
rect 5568 6102 5604 6134
rect 5636 6102 5672 6134
rect 5704 6102 5740 6134
rect 5772 6102 5808 6134
rect 5840 6102 5876 6134
rect 5908 6102 5944 6134
rect 5976 6102 6012 6134
rect 6044 6102 6080 6134
rect 6112 6102 6148 6134
rect 6180 6102 6216 6134
rect 6248 6102 6284 6134
rect 6316 6102 6352 6134
rect 6384 6102 6420 6134
rect 6452 6102 6488 6134
rect 6520 6102 6556 6134
rect 6588 6102 6624 6134
rect 6656 6102 6692 6134
rect 6724 6102 6760 6134
rect 6792 6102 6828 6134
rect 6860 6102 6896 6134
rect 6928 6102 6964 6134
rect 6996 6102 7032 6134
rect 7064 6102 7100 6134
rect 7132 6102 7168 6134
rect 7200 6102 7236 6134
rect 7268 6102 7304 6134
rect 7336 6102 7372 6134
rect 7404 6102 7440 6134
rect 7472 6102 7508 6134
rect 7540 6102 7576 6134
rect 7608 6102 7644 6134
rect 7676 6102 7712 6134
rect 7744 6102 7780 6134
rect 7812 6102 7848 6134
rect 7880 6102 7916 6134
rect 7948 6102 7984 6134
rect 8016 6102 8052 6134
rect 8084 6102 8120 6134
rect 8152 6102 8188 6134
rect 8220 6102 8256 6134
rect 8288 6102 8324 6134
rect 8356 6102 8392 6134
rect 8424 6102 8460 6134
rect 8492 6102 8528 6134
rect 8560 6102 8596 6134
rect 8628 6102 8664 6134
rect 8696 6102 8732 6134
rect 8764 6102 8800 6134
rect 8832 6102 8868 6134
rect 8900 6102 8936 6134
rect 8968 6102 9004 6134
rect 9036 6102 9072 6134
rect 9104 6102 9140 6134
rect 9172 6102 9208 6134
rect 9240 6102 9276 6134
rect 9308 6102 9344 6134
rect 9376 6102 9412 6134
rect 9444 6102 9480 6134
rect 9512 6102 9548 6134
rect 9580 6102 9616 6134
rect 9648 6102 9684 6134
rect 9716 6102 9752 6134
rect 9784 6102 9820 6134
rect 9852 6102 9888 6134
rect 9920 6102 9956 6134
rect 9988 6102 10024 6134
rect 10056 6102 10092 6134
rect 10124 6102 10160 6134
rect 10192 6102 10228 6134
rect 10260 6102 10296 6134
rect 10328 6102 10364 6134
rect 10396 6102 10432 6134
rect 10464 6102 10500 6134
rect 10532 6102 10568 6134
rect 10600 6102 10636 6134
rect 10668 6102 10704 6134
rect 10736 6102 10772 6134
rect 10804 6102 10840 6134
rect 10872 6102 10908 6134
rect 10940 6102 10976 6134
rect 11008 6102 11044 6134
rect 11076 6102 11112 6134
rect 11144 6102 11180 6134
rect 11212 6102 11248 6134
rect 11280 6102 11316 6134
rect 11348 6102 11384 6134
rect 11416 6102 11452 6134
rect 11484 6102 11520 6134
rect 11552 6102 11588 6134
rect 11620 6102 11656 6134
rect 11688 6102 11724 6134
rect 11756 6102 11792 6134
rect 11824 6102 11860 6134
rect 11892 6102 11928 6134
rect 11960 6102 11996 6134
rect 12028 6102 12064 6134
rect 12096 6102 12132 6134
rect 12164 6102 12200 6134
rect 12232 6102 12268 6134
rect 12300 6102 12336 6134
rect 12368 6102 12404 6134
rect 12436 6102 12472 6134
rect 12504 6102 12540 6134
rect 12572 6102 12608 6134
rect 12640 6102 12676 6134
rect 12708 6102 12744 6134
rect 12776 6102 12812 6134
rect 12844 6102 12880 6134
rect 12912 6102 12948 6134
rect 12980 6102 13016 6134
rect 13048 6102 13084 6134
rect 13116 6102 13152 6134
rect 13184 6102 13220 6134
rect 13252 6102 13288 6134
rect 13320 6102 13356 6134
rect 13388 6102 13424 6134
rect 13456 6102 13492 6134
rect 13524 6102 13560 6134
rect 13592 6102 13628 6134
rect 13660 6102 13696 6134
rect 13728 6102 13764 6134
rect 13796 6102 13832 6134
rect 13864 6102 13900 6134
rect 13932 6102 13968 6134
rect 14000 6102 14036 6134
rect 14068 6102 14104 6134
rect 14136 6102 14172 6134
rect 14204 6102 14240 6134
rect 14272 6102 14308 6134
rect 14340 6102 14376 6134
rect 14408 6102 14444 6134
rect 14476 6102 14512 6134
rect 14544 6102 14580 6134
rect 14612 6102 14648 6134
rect 14680 6102 14716 6134
rect 14748 6102 14784 6134
rect 14816 6102 14852 6134
rect 14884 6102 14920 6134
rect 14952 6102 14988 6134
rect 15020 6102 15056 6134
rect 15088 6102 15124 6134
rect 15156 6102 15192 6134
rect 15224 6102 15260 6134
rect 15292 6102 15328 6134
rect 15360 6102 15396 6134
rect 15428 6102 15464 6134
rect 15496 6102 15532 6134
rect 15564 6102 15600 6134
rect 15632 6102 15668 6134
rect 15700 6102 15736 6134
rect 15768 6102 15804 6134
rect 15836 6102 15872 6134
rect 15904 6102 15940 6134
rect 15972 6102 16000 6134
rect 0 6084 16000 6102
rect 0 1200 30 6084
rect 15970 1200 16000 6084
<< psubdiffcont >>
rect 50 31384 82 31416
rect 64 27939 96 27971
rect 18 23089 50 23121
rect 15951 23078 15983 23110
<< nsubdiffcont >>
rect 50 33384 82 33416
rect 50 29684 82 29716
rect 28 12658 60 12690
rect 18 12542 50 12574
rect 15950 12542 15982 12574
rect 28 6102 60 6134
<< metal1 >>
rect 118 33384 150 33416
rect 186 33384 218 33416
rect 254 33384 286 33416
rect 322 33384 354 33416
rect 390 33384 422 33416
rect 458 33384 490 33416
rect 526 33384 558 33416
rect 594 33384 626 33416
rect 662 33384 694 33416
rect 730 33384 762 33416
rect 798 33384 830 33416
rect 866 33384 898 33416
rect 934 33384 966 33416
rect 1002 33384 1034 33416
rect 1070 33384 1102 33416
rect 1138 33384 1170 33416
rect 1206 33384 1238 33416
rect 1274 33384 1306 33416
rect 1342 33384 1374 33416
rect 1410 33384 1442 33416
rect 1478 33384 1510 33416
rect 1546 33384 1578 33416
rect 1614 33384 1646 33416
rect 1682 33384 1714 33416
rect 1750 33384 1782 33416
rect 1818 33384 1850 33416
rect 1886 33384 1918 33416
rect 1954 33384 1986 33416
rect 2022 33384 2054 33416
rect 2090 33384 2122 33416
rect 2158 33384 2190 33416
rect 2226 33384 2258 33416
rect 2294 33384 2326 33416
rect 2362 33384 2394 33416
rect 2430 33384 2462 33416
rect 2498 33384 2530 33416
rect 2566 33384 2598 33416
rect 2634 33384 2666 33416
rect 2702 33384 2734 33416
rect 2770 33384 2802 33416
rect 2838 33384 2870 33416
rect 2906 33384 2938 33416
rect 2974 33384 3006 33416
rect 3042 33384 3074 33416
rect 3110 33384 3142 33416
rect 3178 33384 3210 33416
rect 3246 33384 3278 33416
rect 3314 33384 3346 33416
rect 3382 33384 3414 33416
rect 3450 33384 3482 33416
rect 3518 33384 3550 33416
rect 3586 33384 3618 33416
rect 3654 33384 3686 33416
rect 3722 33384 3754 33416
rect 3790 33384 3822 33416
rect 3858 33384 3890 33416
rect 3926 33384 3958 33416
rect 3994 33384 4026 33416
rect 4062 33384 4094 33416
rect 4130 33384 4162 33416
rect 4198 33384 4230 33416
rect 4266 33384 4298 33416
rect 4334 33384 4366 33416
rect 4402 33384 4434 33416
rect 4470 33384 4502 33416
rect 4538 33384 4570 33416
rect 4606 33384 4638 33416
rect 4674 33384 4706 33416
rect 4742 33384 4774 33416
rect 4810 33384 4842 33416
rect 4878 33384 4910 33416
rect 4946 33384 4978 33416
rect 5014 33384 5046 33416
rect 5082 33384 5114 33416
rect 5150 33384 5182 33416
rect 5218 33384 5250 33416
rect 5286 33384 5318 33416
rect 5354 33384 5386 33416
rect 5422 33384 5454 33416
rect 5490 33384 5522 33416
rect 5558 33384 5590 33416
rect 5626 33384 5658 33416
rect 5694 33384 5726 33416
rect 5762 33384 5794 33416
rect 5830 33384 5862 33416
rect 5898 33384 5930 33416
rect 5966 33384 5998 33416
rect 6034 33384 6066 33416
rect 6102 33384 6134 33416
rect 6170 33384 6202 33416
rect 6238 33384 6270 33416
rect 6306 33384 6338 33416
rect 6374 33384 6406 33416
rect 6442 33384 6474 33416
rect 6510 33384 6542 33416
rect 6578 33384 6610 33416
rect 6646 33384 6678 33416
rect 6714 33384 6746 33416
rect 6782 33384 6814 33416
rect 6850 33384 6882 33416
rect 6918 33384 6950 33416
rect 6986 33384 7018 33416
rect 7054 33384 7086 33416
rect 7122 33384 7154 33416
rect 7190 33384 7222 33416
rect 7258 33384 7290 33416
rect 7326 33384 7358 33416
rect 7394 33384 7426 33416
rect 7462 33384 7494 33416
rect 7530 33384 7562 33416
rect 7598 33384 7630 33416
rect 7666 33384 7698 33416
rect 7734 33384 7766 33416
rect 7802 33384 7834 33416
rect 7870 33384 7902 33416
rect 7938 33384 7970 33416
rect 8006 33384 8038 33416
rect 8074 33384 8106 33416
rect 8142 33384 8174 33416
rect 8210 33384 8242 33416
rect 8278 33384 8310 33416
rect 8346 33384 8378 33416
rect 8414 33384 8446 33416
rect 8482 33384 8514 33416
rect 8550 33384 8582 33416
rect 8618 33384 8650 33416
rect 8686 33384 8718 33416
rect 8754 33384 8786 33416
rect 8822 33384 8854 33416
rect 8890 33384 8922 33416
rect 8958 33384 8990 33416
rect 9026 33384 9058 33416
rect 9094 33384 9126 33416
rect 9162 33384 9194 33416
rect 9230 33384 9262 33416
rect 9298 33384 9330 33416
rect 9366 33384 9398 33416
rect 9434 33384 9466 33416
rect 9502 33384 9534 33416
rect 9570 33384 9602 33416
rect 9638 33384 9670 33416
rect 9706 33384 9738 33416
rect 9774 33384 9806 33416
rect 9842 33384 9874 33416
rect 9910 33384 9942 33416
rect 9978 33384 10010 33416
rect 10046 33384 10078 33416
rect 10114 33384 10146 33416
rect 10182 33384 10214 33416
rect 10250 33384 10282 33416
rect 10318 33384 10350 33416
rect 10386 33384 10418 33416
rect 10454 33384 10486 33416
rect 10522 33384 10554 33416
rect 10590 33384 10622 33416
rect 10658 33384 10690 33416
rect 10726 33384 10758 33416
rect 10794 33384 10826 33416
rect 10862 33384 10894 33416
rect 10930 33384 10962 33416
rect 10998 33384 11030 33416
rect 11066 33384 11098 33416
rect 11134 33384 11166 33416
rect 11202 33384 11234 33416
rect 11270 33384 11302 33416
rect 11338 33384 11370 33416
rect 11406 33384 11438 33416
rect 11474 33384 11506 33416
rect 11542 33384 11574 33416
rect 11610 33384 11642 33416
rect 11678 33384 11710 33416
rect 11746 33384 11778 33416
rect 11814 33384 11846 33416
rect 11882 33384 11914 33416
rect 11950 33384 11982 33416
rect 12018 33384 12050 33416
rect 12086 33384 12118 33416
rect 12154 33384 12186 33416
rect 12222 33384 12254 33416
rect 12290 33384 12322 33416
rect 12358 33384 12390 33416
rect 12426 33384 12458 33416
rect 12494 33384 12526 33416
rect 12562 33384 12594 33416
rect 12630 33384 12662 33416
rect 12698 33384 12730 33416
rect 12766 33384 12798 33416
rect 12834 33384 12866 33416
rect 12902 33384 12934 33416
rect 12970 33384 13002 33416
rect 13038 33384 13070 33416
rect 13106 33384 13138 33416
rect 13174 33384 13206 33416
rect 13242 33384 13274 33416
rect 13310 33384 13342 33416
rect 13378 33384 13410 33416
rect 13446 33384 13478 33416
rect 13514 33384 13546 33416
rect 13582 33384 13614 33416
rect 13650 33384 13682 33416
rect 13718 33384 13750 33416
rect 13786 33384 13818 33416
rect 13854 33384 13886 33416
rect 13922 33384 13954 33416
rect 13990 33384 14022 33416
rect 14058 33384 14090 33416
rect 14126 33384 14158 33416
rect 14194 33384 14226 33416
rect 14262 33384 14294 33416
rect 14330 33384 14362 33416
rect 14398 33384 14430 33416
rect 14466 33384 14498 33416
rect 14534 33384 14566 33416
rect 14602 33384 14634 33416
rect 14670 33384 14702 33416
rect 14738 33384 14770 33416
rect 14806 33384 14838 33416
rect 14874 33384 14906 33416
rect 14942 33384 14974 33416
rect 15010 33384 15042 33416
rect 15078 33384 15110 33416
rect 15146 33384 15178 33416
rect 15214 33384 15246 33416
rect 15282 33384 15314 33416
rect 15350 33384 15382 33416
rect 15442 33384 15474 33416
rect 15510 33384 15542 33416
rect 15578 33384 15610 33416
rect 15646 33384 15678 33416
rect 15714 33384 15746 33416
rect 15782 33384 15814 33416
rect 15850 33384 15882 33416
rect 15918 33384 15950 33416
rect 118 29684 150 29716
rect 186 29684 218 29716
rect 254 29684 286 29716
rect 322 29684 354 29716
rect 390 29684 422 29716
rect 458 29684 490 29716
rect 526 29684 558 29716
rect 594 29684 626 29716
rect 662 29684 694 29716
rect 730 29684 762 29716
rect 798 29684 830 29716
rect 866 29684 898 29716
rect 934 29684 966 29716
rect 1002 29684 1034 29716
rect 1070 29684 1102 29716
rect 1138 29684 1170 29716
rect 1206 29684 1238 29716
rect 1274 29684 1306 29716
rect 1342 29684 1374 29716
rect 1410 29684 1442 29716
rect 1478 29684 1510 29716
rect 1546 29684 1578 29716
rect 1614 29684 1646 29716
rect 1682 29684 1714 29716
rect 1750 29684 1782 29716
rect 1818 29684 1850 29716
rect 1886 29684 1918 29716
rect 1954 29684 1986 29716
rect 2022 29684 2054 29716
rect 2090 29684 2122 29716
rect 2158 29684 2190 29716
rect 2226 29684 2258 29716
rect 2294 29684 2326 29716
rect 2362 29684 2394 29716
rect 2430 29684 2462 29716
rect 2498 29684 2530 29716
rect 2566 29684 2598 29716
rect 2634 29684 2666 29716
rect 2702 29684 2734 29716
rect 2770 29684 2802 29716
rect 2838 29684 2870 29716
rect 2906 29684 2938 29716
rect 2974 29684 3006 29716
rect 3042 29684 3074 29716
rect 3110 29684 3142 29716
rect 3178 29684 3210 29716
rect 3246 29684 3278 29716
rect 3314 29684 3346 29716
rect 3382 29684 3414 29716
rect 3450 29684 3482 29716
rect 3518 29684 3550 29716
rect 3586 29684 3618 29716
rect 3654 29684 3686 29716
rect 3722 29684 3754 29716
rect 3790 29684 3822 29716
rect 3858 29684 3890 29716
rect 3926 29684 3958 29716
rect 3994 29684 4026 29716
rect 4062 29684 4094 29716
rect 4130 29684 4162 29716
rect 4198 29684 4230 29716
rect 4266 29684 4298 29716
rect 4334 29684 4366 29716
rect 4402 29684 4434 29716
rect 4470 29684 4502 29716
rect 4538 29684 4570 29716
rect 4606 29684 4638 29716
rect 4674 29684 4706 29716
rect 4742 29684 4774 29716
rect 4810 29684 4842 29716
rect 4878 29684 4910 29716
rect 4946 29684 4978 29716
rect 5014 29684 5046 29716
rect 5082 29684 5114 29716
rect 5150 29684 5182 29716
rect 5218 29684 5250 29716
rect 5286 29684 5318 29716
rect 5354 29684 5386 29716
rect 5422 29684 5454 29716
rect 5490 29684 5522 29716
rect 5558 29684 5590 29716
rect 5626 29684 5658 29716
rect 5694 29684 5726 29716
rect 5762 29684 5794 29716
rect 5830 29684 5862 29716
rect 5898 29684 5930 29716
rect 5966 29684 5998 29716
rect 6034 29684 6066 29716
rect 6102 29684 6134 29716
rect 6170 29684 6202 29716
rect 6238 29684 6270 29716
rect 6306 29684 6338 29716
rect 6374 29684 6406 29716
rect 6442 29684 6474 29716
rect 6510 29684 6542 29716
rect 6578 29684 6610 29716
rect 6646 29684 6678 29716
rect 6714 29684 6746 29716
rect 6782 29684 6814 29716
rect 6850 29684 6882 29716
rect 6918 29684 6950 29716
rect 6986 29684 7018 29716
rect 7054 29684 7086 29716
rect 7122 29684 7154 29716
rect 7190 29684 7222 29716
rect 7258 29684 7290 29716
rect 7326 29684 7358 29716
rect 7394 29684 7426 29716
rect 7462 29684 7494 29716
rect 7530 29684 7562 29716
rect 7598 29684 7630 29716
rect 7666 29684 7698 29716
rect 7734 29684 7766 29716
rect 7802 29684 7834 29716
rect 7870 29684 7902 29716
rect 7938 29684 7970 29716
rect 8006 29684 8038 29716
rect 8074 29684 8106 29716
rect 8142 29684 8174 29716
rect 8210 29684 8242 29716
rect 8278 29684 8310 29716
rect 8346 29684 8378 29716
rect 8414 29684 8446 29716
rect 8482 29684 8514 29716
rect 8550 29684 8582 29716
rect 8618 29684 8650 29716
rect 8686 29684 8718 29716
rect 8754 29684 8786 29716
rect 8822 29684 8854 29716
rect 8890 29684 8922 29716
rect 8958 29684 8990 29716
rect 9026 29684 9058 29716
rect 9094 29684 9126 29716
rect 9162 29684 9194 29716
rect 9230 29684 9262 29716
rect 9298 29684 9330 29716
rect 9366 29684 9398 29716
rect 9434 29684 9466 29716
rect 9502 29684 9534 29716
rect 9570 29684 9602 29716
rect 9638 29684 9670 29716
rect 9706 29684 9738 29716
rect 9774 29684 9806 29716
rect 9842 29684 9874 29716
rect 9910 29684 9942 29716
rect 9978 29684 10010 29716
rect 10046 29684 10078 29716
rect 10114 29684 10146 29716
rect 10182 29684 10214 29716
rect 10250 29684 10282 29716
rect 10318 29684 10350 29716
rect 10386 29684 10418 29716
rect 10454 29684 10486 29716
rect 10522 29684 10554 29716
rect 10590 29684 10622 29716
rect 10658 29684 10690 29716
rect 10726 29684 10758 29716
rect 10794 29684 10826 29716
rect 10862 29684 10894 29716
rect 10930 29684 10962 29716
rect 10998 29684 11030 29716
rect 11066 29684 11098 29716
rect 11134 29684 11166 29716
rect 11202 29684 11234 29716
rect 11270 29684 11302 29716
rect 11338 29684 11370 29716
rect 11406 29684 11438 29716
rect 11474 29684 11506 29716
rect 11542 29684 11574 29716
rect 11610 29684 11642 29716
rect 11678 29684 11710 29716
rect 11746 29684 11778 29716
rect 11814 29684 11846 29716
rect 11882 29684 11914 29716
rect 11950 29684 11982 29716
rect 12018 29684 12050 29716
rect 12086 29684 12118 29716
rect 12154 29684 12186 29716
rect 12222 29684 12254 29716
rect 12290 29684 12322 29716
rect 12358 29684 12390 29716
rect 12426 29684 12458 29716
rect 12494 29684 12526 29716
rect 12562 29684 12594 29716
rect 12630 29684 12662 29716
rect 12698 29684 12730 29716
rect 12766 29684 12798 29716
rect 12834 29684 12866 29716
rect 12902 29684 12934 29716
rect 12970 29684 13002 29716
rect 13038 29684 13070 29716
rect 13106 29684 13138 29716
rect 13174 29684 13206 29716
rect 13242 29684 13274 29716
rect 13310 29684 13342 29716
rect 13378 29684 13410 29716
rect 13446 29684 13478 29716
rect 13514 29684 13546 29716
rect 13582 29684 13614 29716
rect 13650 29684 13682 29716
rect 13718 29684 13750 29716
rect 13786 29684 13818 29716
rect 13854 29684 13886 29716
rect 13922 29684 13954 29716
rect 13990 29684 14022 29716
rect 14058 29684 14090 29716
rect 14126 29684 14158 29716
rect 14194 29684 14226 29716
rect 14262 29684 14294 29716
rect 14330 29684 14362 29716
rect 14398 29684 14430 29716
rect 14466 29684 14498 29716
rect 14534 29684 14566 29716
rect 14602 29684 14634 29716
rect 14670 29684 14702 29716
rect 14738 29684 14770 29716
rect 14806 29684 14838 29716
rect 14874 29684 14906 29716
rect 14942 29684 14974 29716
rect 15010 29684 15042 29716
rect 15078 29684 15110 29716
rect 15146 29684 15178 29716
rect 15214 29684 15246 29716
rect 15282 29684 15314 29716
rect 15350 29684 15382 29716
rect 15442 29684 15474 29716
rect 15510 29684 15542 29716
rect 15578 29684 15610 29716
rect 15646 29684 15678 29716
rect 15714 29684 15746 29716
rect 15782 29684 15814 29716
rect 15850 29684 15882 29716
rect 15918 29684 15950 29716
rect 96 12658 128 12690
rect 164 12658 196 12690
rect 232 12658 264 12690
rect 300 12658 332 12690
rect 368 12658 400 12690
rect 436 12658 468 12690
rect 504 12658 536 12690
rect 572 12658 604 12690
rect 640 12658 672 12690
rect 708 12658 740 12690
rect 776 12658 808 12690
rect 844 12658 876 12690
rect 912 12658 944 12690
rect 980 12658 1012 12690
rect 1048 12658 1080 12690
rect 1116 12658 1148 12690
rect 1184 12658 1216 12690
rect 1252 12658 1284 12690
rect 1320 12658 1352 12690
rect 1388 12658 1420 12690
rect 1456 12658 1488 12690
rect 1524 12658 1556 12690
rect 1592 12658 1624 12690
rect 1660 12658 1692 12690
rect 1728 12658 1760 12690
rect 1796 12658 1828 12690
rect 1864 12658 1896 12690
rect 1932 12658 1964 12690
rect 2000 12658 2032 12690
rect 2068 12658 2100 12690
rect 2136 12658 2168 12690
rect 2204 12658 2236 12690
rect 2272 12658 2304 12690
rect 2340 12658 2372 12690
rect 2408 12658 2440 12690
rect 2476 12658 2508 12690
rect 2544 12658 2576 12690
rect 2612 12658 2644 12690
rect 2680 12658 2712 12690
rect 2748 12658 2780 12690
rect 2816 12658 2848 12690
rect 2884 12658 2916 12690
rect 2952 12658 2984 12690
rect 3020 12658 3052 12690
rect 3088 12658 3120 12690
rect 3156 12658 3188 12690
rect 3224 12658 3256 12690
rect 3292 12658 3324 12690
rect 3360 12658 3392 12690
rect 3428 12658 3460 12690
rect 3496 12658 3528 12690
rect 3564 12658 3596 12690
rect 3632 12658 3664 12690
rect 3700 12658 3732 12690
rect 3768 12658 3800 12690
rect 3836 12658 3868 12690
rect 3904 12658 3936 12690
rect 3972 12658 4004 12690
rect 4040 12658 4072 12690
rect 4108 12658 4140 12690
rect 4176 12658 4208 12690
rect 4244 12658 4276 12690
rect 4312 12658 4344 12690
rect 4380 12658 4412 12690
rect 4448 12658 4480 12690
rect 4516 12658 4548 12690
rect 4584 12658 4616 12690
rect 4652 12658 4684 12690
rect 4720 12658 4752 12690
rect 4788 12658 4820 12690
rect 4856 12658 4888 12690
rect 4924 12658 4956 12690
rect 4992 12658 5024 12690
rect 5060 12658 5092 12690
rect 5128 12658 5160 12690
rect 5196 12658 5228 12690
rect 5264 12658 5296 12690
rect 5332 12658 5364 12690
rect 5400 12658 5432 12690
rect 5468 12658 5500 12690
rect 5536 12658 5568 12690
rect 5604 12658 5636 12690
rect 5672 12658 5704 12690
rect 5740 12658 5772 12690
rect 5808 12658 5840 12690
rect 5876 12658 5908 12690
rect 5944 12658 5976 12690
rect 6012 12658 6044 12690
rect 6080 12658 6112 12690
rect 6148 12658 6180 12690
rect 6216 12658 6248 12690
rect 6284 12658 6316 12690
rect 6352 12658 6384 12690
rect 6420 12658 6452 12690
rect 6488 12658 6520 12690
rect 6556 12658 6588 12690
rect 6624 12658 6656 12690
rect 6692 12658 6724 12690
rect 6760 12658 6792 12690
rect 6828 12658 6860 12690
rect 6896 12658 6928 12690
rect 6964 12658 6996 12690
rect 7032 12658 7064 12690
rect 7100 12658 7132 12690
rect 7168 12658 7200 12690
rect 7236 12658 7268 12690
rect 7304 12658 7336 12690
rect 7372 12658 7404 12690
rect 7440 12658 7472 12690
rect 7508 12658 7540 12690
rect 7576 12658 7608 12690
rect 7644 12658 7676 12690
rect 7712 12658 7744 12690
rect 7780 12658 7812 12690
rect 7848 12658 7880 12690
rect 7916 12658 7948 12690
rect 7984 12658 8016 12690
rect 8052 12658 8084 12690
rect 8120 12658 8152 12690
rect 8188 12658 8220 12690
rect 8256 12658 8288 12690
rect 8324 12658 8356 12690
rect 8392 12658 8424 12690
rect 8460 12658 8492 12690
rect 8528 12658 8560 12690
rect 8596 12658 8628 12690
rect 8664 12658 8696 12690
rect 8732 12658 8764 12690
rect 8800 12658 8832 12690
rect 8868 12658 8900 12690
rect 8936 12658 8968 12690
rect 9004 12658 9036 12690
rect 9072 12658 9104 12690
rect 9140 12658 9172 12690
rect 9208 12658 9240 12690
rect 9276 12658 9308 12690
rect 9344 12658 9376 12690
rect 9412 12658 9444 12690
rect 9480 12658 9512 12690
rect 9548 12658 9580 12690
rect 9616 12658 9648 12690
rect 9684 12658 9716 12690
rect 9752 12658 9784 12690
rect 9820 12658 9852 12690
rect 9888 12658 9920 12690
rect 9956 12658 9988 12690
rect 10024 12658 10056 12690
rect 10092 12658 10124 12690
rect 10160 12658 10192 12690
rect 10228 12658 10260 12690
rect 10296 12658 10328 12690
rect 10364 12658 10396 12690
rect 10432 12658 10464 12690
rect 10500 12658 10532 12690
rect 10568 12658 10600 12690
rect 10636 12658 10668 12690
rect 10704 12658 10736 12690
rect 10772 12658 10804 12690
rect 10840 12658 10872 12690
rect 10908 12658 10940 12690
rect 10976 12658 11008 12690
rect 11044 12658 11076 12690
rect 11112 12658 11144 12690
rect 11180 12658 11212 12690
rect 11248 12658 11280 12690
rect 11316 12658 11348 12690
rect 11384 12658 11416 12690
rect 11452 12658 11484 12690
rect 11520 12658 11552 12690
rect 11588 12658 11620 12690
rect 11656 12658 11688 12690
rect 11724 12658 11756 12690
rect 11792 12658 11824 12690
rect 11860 12658 11892 12690
rect 11928 12658 11960 12690
rect 11996 12658 12028 12690
rect 12064 12658 12096 12690
rect 12132 12658 12164 12690
rect 12200 12658 12232 12690
rect 12268 12658 12300 12690
rect 12336 12658 12368 12690
rect 12404 12658 12436 12690
rect 12472 12658 12504 12690
rect 12540 12658 12572 12690
rect 12608 12658 12640 12690
rect 12676 12658 12708 12690
rect 12744 12658 12776 12690
rect 12812 12658 12844 12690
rect 12880 12658 12912 12690
rect 12948 12658 12980 12690
rect 13016 12658 13048 12690
rect 13084 12658 13116 12690
rect 13152 12658 13184 12690
rect 13220 12658 13252 12690
rect 13288 12658 13320 12690
rect 13356 12658 13388 12690
rect 13424 12658 13456 12690
rect 13492 12658 13524 12690
rect 13560 12658 13592 12690
rect 13628 12658 13660 12690
rect 13696 12658 13728 12690
rect 13764 12658 13796 12690
rect 13832 12658 13864 12690
rect 13900 12658 13932 12690
rect 13968 12658 14000 12690
rect 14036 12658 14068 12690
rect 14104 12658 14136 12690
rect 14172 12658 14204 12690
rect 14240 12658 14272 12690
rect 14308 12658 14340 12690
rect 14376 12658 14408 12690
rect 14444 12658 14476 12690
rect 14512 12658 14544 12690
rect 14580 12658 14612 12690
rect 14648 12658 14680 12690
rect 14716 12658 14748 12690
rect 14784 12658 14816 12690
rect 14852 12658 14884 12690
rect 14920 12658 14952 12690
rect 14988 12658 15020 12690
rect 15056 12658 15088 12690
rect 15124 12658 15156 12690
rect 15192 12658 15224 12690
rect 15260 12658 15292 12690
rect 15328 12658 15360 12690
rect 15396 12658 15428 12690
rect 15464 12658 15496 12690
rect 15532 12658 15564 12690
rect 15600 12658 15632 12690
rect 15668 12658 15700 12690
rect 15736 12658 15768 12690
rect 15804 12658 15836 12690
rect 15872 12658 15904 12690
rect 15940 12658 15972 12690
rect 18 12474 50 12506
rect 18 12406 50 12438
rect 18 12338 50 12370
rect 18 12270 50 12302
rect 18 12202 50 12234
rect 18 12134 50 12166
rect 18 12066 50 12098
rect 18 11998 50 12030
rect 18 11930 50 11962
rect 18 11862 50 11894
rect 18 11794 50 11826
rect 18 11726 50 11758
rect 18 11658 50 11690
rect 18 11590 50 11622
rect 18 11522 50 11554
rect 18 11454 50 11486
rect 18 11386 50 11418
rect 18 11318 50 11350
rect 18 11250 50 11282
rect 18 11182 50 11214
rect 18 11114 50 11146
rect 18 11046 50 11078
rect 18 10978 50 11010
rect 18 10910 50 10942
rect 18 10842 50 10874
rect 18 10774 50 10806
rect 18 10706 50 10738
rect 18 10638 50 10670
rect 18 10570 50 10602
rect 18 10502 50 10534
rect 18 10434 50 10466
rect 18 10366 50 10398
rect 18 10298 50 10330
rect 18 10230 50 10262
rect 18 10162 50 10194
rect 18 10094 50 10126
rect 18 10026 50 10058
rect 18 9958 50 9990
rect 18 9890 50 9922
rect 18 9822 50 9854
rect 18 9754 50 9786
rect 18 9686 50 9718
rect 18 9618 50 9650
rect 18 9550 50 9582
rect 18 9482 50 9514
rect 18 9414 50 9446
rect 18 9346 50 9378
rect 18 9278 50 9310
rect 18 9210 50 9242
rect 18 9142 50 9174
rect 18 9074 50 9106
rect 18 9006 50 9038
rect 18 8938 50 8970
rect 18 8870 50 8902
rect 18 8802 50 8834
rect 18 8734 50 8766
rect 18 8666 50 8698
rect 18 8598 50 8630
rect 18 8530 50 8562
rect 18 8462 50 8494
rect 18 8394 50 8426
rect 18 8326 50 8358
rect 18 8258 50 8290
rect 18 8190 50 8222
rect 18 8122 50 8154
rect 18 8054 50 8086
rect 18 7986 50 8018
rect 18 7918 50 7950
rect 18 7850 50 7882
rect 18 7782 50 7814
rect 18 7714 50 7746
rect 18 7646 50 7678
rect 18 7578 50 7610
rect 18 7510 50 7542
rect 18 7442 50 7474
rect 18 7374 50 7406
rect 18 7306 50 7338
rect 18 7238 50 7270
rect 18 7170 50 7202
rect 18 7102 50 7134
rect 18 7034 50 7066
rect 18 6966 50 6998
rect 18 6898 50 6930
rect 18 6830 50 6862
rect 18 6762 50 6794
rect 18 6694 50 6726
rect 18 6626 50 6658
rect 18 6558 50 6590
rect 18 6490 50 6522
rect 18 6422 50 6454
rect 18 6354 50 6386
rect 18 6286 50 6318
rect 18 6218 50 6250
rect 15950 12474 15982 12506
rect 15950 12406 15982 12438
rect 15950 12338 15982 12370
rect 15950 12270 15982 12302
rect 15950 12202 15982 12234
rect 15950 12134 15982 12166
rect 15950 12066 15982 12098
rect 15950 11998 15982 12030
rect 15950 11930 15982 11962
rect 15950 11862 15982 11894
rect 15950 11794 15982 11826
rect 15950 11726 15982 11758
rect 15950 11658 15982 11690
rect 15950 11590 15982 11622
rect 15950 11522 15982 11554
rect 15950 11454 15982 11486
rect 15950 11386 15982 11418
rect 15950 11318 15982 11350
rect 15950 11250 15982 11282
rect 15950 11182 15982 11214
rect 15950 11114 15982 11146
rect 15950 11046 15982 11078
rect 15950 10978 15982 11010
rect 15950 10910 15982 10942
rect 15950 10842 15982 10874
rect 15950 10774 15982 10806
rect 15950 10706 15982 10738
rect 15950 10638 15982 10670
rect 15950 10570 15982 10602
rect 15950 10502 15982 10534
rect 15950 10434 15982 10466
rect 15950 10366 15982 10398
rect 15950 10298 15982 10330
rect 15950 10230 15982 10262
rect 15950 10162 15982 10194
rect 15950 10094 15982 10126
rect 15950 10026 15982 10058
rect 15950 9958 15982 9990
rect 15950 9890 15982 9922
rect 15950 9822 15982 9854
rect 15950 9754 15982 9786
rect 15950 9686 15982 9718
rect 15950 9618 15982 9650
rect 15950 9550 15982 9582
rect 15950 9482 15982 9514
rect 15950 9414 15982 9446
rect 15950 9346 15982 9378
rect 15950 9278 15982 9310
rect 15950 9210 15982 9242
rect 15950 9142 15982 9174
rect 15950 9074 15982 9106
rect 15950 9006 15982 9038
rect 15950 8938 15982 8970
rect 15950 8870 15982 8902
rect 15950 8802 15982 8834
rect 15950 8734 15982 8766
rect 15950 8666 15982 8698
rect 15950 8598 15982 8630
rect 15950 8530 15982 8562
rect 15950 8462 15982 8494
rect 15950 8394 15982 8426
rect 15950 8326 15982 8358
rect 15950 8258 15982 8290
rect 15950 8190 15982 8222
rect 15950 8122 15982 8154
rect 15950 8054 15982 8086
rect 15950 7986 15982 8018
rect 15950 7918 15982 7950
rect 15950 7850 15982 7882
rect 15950 7782 15982 7814
rect 15950 7714 15982 7746
rect 15950 7646 15982 7678
rect 15950 7578 15982 7610
rect 15950 7510 15982 7542
rect 15950 7442 15982 7474
rect 15950 7374 15982 7406
rect 15950 7306 15982 7338
rect 15950 7238 15982 7270
rect 15950 7170 15982 7202
rect 15950 7102 15982 7134
rect 15950 7034 15982 7066
rect 15950 6966 15982 6998
rect 15950 6898 15982 6930
rect 15950 6830 15982 6862
rect 15950 6762 15982 6794
rect 15950 6694 15982 6726
rect 15950 6626 15982 6658
rect 15950 6558 15982 6590
rect 15950 6490 15982 6522
rect 15950 6422 15982 6454
rect 15950 6354 15982 6386
rect 15950 6286 15982 6318
rect 15950 6218 15982 6250
rect 96 6102 128 6134
rect 164 6102 196 6134
rect 232 6102 264 6134
rect 300 6102 332 6134
rect 368 6102 400 6134
rect 436 6102 468 6134
rect 504 6102 536 6134
rect 572 6102 604 6134
rect 640 6102 672 6134
rect 708 6102 740 6134
rect 776 6102 808 6134
rect 844 6102 876 6134
rect 912 6102 944 6134
rect 980 6102 1012 6134
rect 1048 6102 1080 6134
rect 1116 6102 1148 6134
rect 1184 6102 1216 6134
rect 1252 6102 1284 6134
rect 1320 6102 1352 6134
rect 1388 6102 1420 6134
rect 1456 6102 1488 6134
rect 1524 6102 1556 6134
rect 1592 6102 1624 6134
rect 1660 6102 1692 6134
rect 1728 6102 1760 6134
rect 1796 6102 1828 6134
rect 1864 6102 1896 6134
rect 1932 6102 1964 6134
rect 2000 6102 2032 6134
rect 2068 6102 2100 6134
rect 2136 6102 2168 6134
rect 2204 6102 2236 6134
rect 2272 6102 2304 6134
rect 2340 6102 2372 6134
rect 2408 6102 2440 6134
rect 2476 6102 2508 6134
rect 2544 6102 2576 6134
rect 2612 6102 2644 6134
rect 2680 6102 2712 6134
rect 2748 6102 2780 6134
rect 2816 6102 2848 6134
rect 2884 6102 2916 6134
rect 2952 6102 2984 6134
rect 3020 6102 3052 6134
rect 3088 6102 3120 6134
rect 3156 6102 3188 6134
rect 3224 6102 3256 6134
rect 3292 6102 3324 6134
rect 3360 6102 3392 6134
rect 3428 6102 3460 6134
rect 3496 6102 3528 6134
rect 3564 6102 3596 6134
rect 3632 6102 3664 6134
rect 3700 6102 3732 6134
rect 3768 6102 3800 6134
rect 3836 6102 3868 6134
rect 3904 6102 3936 6134
rect 3972 6102 4004 6134
rect 4040 6102 4072 6134
rect 4108 6102 4140 6134
rect 4176 6102 4208 6134
rect 4244 6102 4276 6134
rect 4312 6102 4344 6134
rect 4380 6102 4412 6134
rect 4448 6102 4480 6134
rect 4516 6102 4548 6134
rect 4584 6102 4616 6134
rect 4652 6102 4684 6134
rect 4720 6102 4752 6134
rect 4788 6102 4820 6134
rect 4856 6102 4888 6134
rect 4924 6102 4956 6134
rect 4992 6102 5024 6134
rect 5060 6102 5092 6134
rect 5128 6102 5160 6134
rect 5196 6102 5228 6134
rect 5264 6102 5296 6134
rect 5332 6102 5364 6134
rect 5400 6102 5432 6134
rect 5468 6102 5500 6134
rect 5536 6102 5568 6134
rect 5604 6102 5636 6134
rect 5672 6102 5704 6134
rect 5740 6102 5772 6134
rect 5808 6102 5840 6134
rect 5876 6102 5908 6134
rect 5944 6102 5976 6134
rect 6012 6102 6044 6134
rect 6080 6102 6112 6134
rect 6148 6102 6180 6134
rect 6216 6102 6248 6134
rect 6284 6102 6316 6134
rect 6352 6102 6384 6134
rect 6420 6102 6452 6134
rect 6488 6102 6520 6134
rect 6556 6102 6588 6134
rect 6624 6102 6656 6134
rect 6692 6102 6724 6134
rect 6760 6102 6792 6134
rect 6828 6102 6860 6134
rect 6896 6102 6928 6134
rect 6964 6102 6996 6134
rect 7032 6102 7064 6134
rect 7100 6102 7132 6134
rect 7168 6102 7200 6134
rect 7236 6102 7268 6134
rect 7304 6102 7336 6134
rect 7372 6102 7404 6134
rect 7440 6102 7472 6134
rect 7508 6102 7540 6134
rect 7576 6102 7608 6134
rect 7644 6102 7676 6134
rect 7712 6102 7744 6134
rect 7780 6102 7812 6134
rect 7848 6102 7880 6134
rect 7916 6102 7948 6134
rect 7984 6102 8016 6134
rect 8052 6102 8084 6134
rect 8120 6102 8152 6134
rect 8188 6102 8220 6134
rect 8256 6102 8288 6134
rect 8324 6102 8356 6134
rect 8392 6102 8424 6134
rect 8460 6102 8492 6134
rect 8528 6102 8560 6134
rect 8596 6102 8628 6134
rect 8664 6102 8696 6134
rect 8732 6102 8764 6134
rect 8800 6102 8832 6134
rect 8868 6102 8900 6134
rect 8936 6102 8968 6134
rect 9004 6102 9036 6134
rect 9072 6102 9104 6134
rect 9140 6102 9172 6134
rect 9208 6102 9240 6134
rect 9276 6102 9308 6134
rect 9344 6102 9376 6134
rect 9412 6102 9444 6134
rect 9480 6102 9512 6134
rect 9548 6102 9580 6134
rect 9616 6102 9648 6134
rect 9684 6102 9716 6134
rect 9752 6102 9784 6134
rect 9820 6102 9852 6134
rect 9888 6102 9920 6134
rect 9956 6102 9988 6134
rect 10024 6102 10056 6134
rect 10092 6102 10124 6134
rect 10160 6102 10192 6134
rect 10228 6102 10260 6134
rect 10296 6102 10328 6134
rect 10364 6102 10396 6134
rect 10432 6102 10464 6134
rect 10500 6102 10532 6134
rect 10568 6102 10600 6134
rect 10636 6102 10668 6134
rect 10704 6102 10736 6134
rect 10772 6102 10804 6134
rect 10840 6102 10872 6134
rect 10908 6102 10940 6134
rect 10976 6102 11008 6134
rect 11044 6102 11076 6134
rect 11112 6102 11144 6134
rect 11180 6102 11212 6134
rect 11248 6102 11280 6134
rect 11316 6102 11348 6134
rect 11384 6102 11416 6134
rect 11452 6102 11484 6134
rect 11520 6102 11552 6134
rect 11588 6102 11620 6134
rect 11656 6102 11688 6134
rect 11724 6102 11756 6134
rect 11792 6102 11824 6134
rect 11860 6102 11892 6134
rect 11928 6102 11960 6134
rect 11996 6102 12028 6134
rect 12064 6102 12096 6134
rect 12132 6102 12164 6134
rect 12200 6102 12232 6134
rect 12268 6102 12300 6134
rect 12336 6102 12368 6134
rect 12404 6102 12436 6134
rect 12472 6102 12504 6134
rect 12540 6102 12572 6134
rect 12608 6102 12640 6134
rect 12676 6102 12708 6134
rect 12744 6102 12776 6134
rect 12812 6102 12844 6134
rect 12880 6102 12912 6134
rect 12948 6102 12980 6134
rect 13016 6102 13048 6134
rect 13084 6102 13116 6134
rect 13152 6102 13184 6134
rect 13220 6102 13252 6134
rect 13288 6102 13320 6134
rect 13356 6102 13388 6134
rect 13424 6102 13456 6134
rect 13492 6102 13524 6134
rect 13560 6102 13592 6134
rect 13628 6102 13660 6134
rect 13696 6102 13728 6134
rect 13764 6102 13796 6134
rect 13832 6102 13864 6134
rect 13900 6102 13932 6134
rect 13968 6102 14000 6134
rect 14036 6102 14068 6134
rect 14104 6102 14136 6134
rect 14172 6102 14204 6134
rect 14240 6102 14272 6134
rect 14308 6102 14340 6134
rect 14376 6102 14408 6134
rect 14444 6102 14476 6134
rect 14512 6102 14544 6134
rect 14580 6102 14612 6134
rect 14648 6102 14680 6134
rect 14716 6102 14748 6134
rect 14784 6102 14816 6134
rect 14852 6102 14884 6134
rect 14920 6102 14952 6134
rect 14988 6102 15020 6134
rect 15056 6102 15088 6134
rect 15124 6102 15156 6134
rect 15192 6102 15224 6134
rect 15260 6102 15292 6134
rect 15328 6102 15360 6134
rect 15396 6102 15428 6134
rect 15464 6102 15496 6134
rect 15532 6102 15564 6134
rect 15600 6102 15632 6134
rect 15668 6102 15700 6134
rect 15736 6102 15768 6134
rect 15804 6102 15836 6134
rect 15872 6102 15904 6134
rect 15940 6102 15972 6134
rect 118 31384 150 31416
rect 186 31384 218 31416
rect 254 31384 286 31416
rect 322 31384 354 31416
rect 390 31384 422 31416
rect 458 31384 490 31416
rect 526 31384 558 31416
rect 594 31384 626 31416
rect 662 31384 694 31416
rect 730 31384 762 31416
rect 798 31384 830 31416
rect 866 31384 898 31416
rect 934 31384 966 31416
rect 1002 31384 1034 31416
rect 1070 31384 1102 31416
rect 1138 31384 1170 31416
rect 1206 31384 1238 31416
rect 1274 31384 1306 31416
rect 1342 31384 1374 31416
rect 1410 31384 1442 31416
rect 1478 31384 1510 31416
rect 1546 31384 1578 31416
rect 1614 31384 1646 31416
rect 1682 31384 1714 31416
rect 1750 31384 1782 31416
rect 1818 31384 1850 31416
rect 1886 31384 1918 31416
rect 1954 31384 1986 31416
rect 2022 31384 2054 31416
rect 2090 31384 2122 31416
rect 2158 31384 2190 31416
rect 2226 31384 2258 31416
rect 2294 31384 2326 31416
rect 2362 31384 2394 31416
rect 2430 31384 2462 31416
rect 2498 31384 2530 31416
rect 2566 31384 2598 31416
rect 2634 31384 2666 31416
rect 2702 31384 2734 31416
rect 2770 31384 2802 31416
rect 2838 31384 2870 31416
rect 2906 31384 2938 31416
rect 2974 31384 3006 31416
rect 3042 31384 3074 31416
rect 3110 31384 3142 31416
rect 3178 31384 3210 31416
rect 3246 31384 3278 31416
rect 3314 31384 3346 31416
rect 3382 31384 3414 31416
rect 3450 31384 3482 31416
rect 3518 31384 3550 31416
rect 3586 31384 3618 31416
rect 3654 31384 3686 31416
rect 3722 31384 3754 31416
rect 3790 31384 3822 31416
rect 3858 31384 3890 31416
rect 3926 31384 3958 31416
rect 3994 31384 4026 31416
rect 4062 31384 4094 31416
rect 4130 31384 4162 31416
rect 4198 31384 4230 31416
rect 4266 31384 4298 31416
rect 4334 31384 4366 31416
rect 4402 31384 4434 31416
rect 4470 31384 4502 31416
rect 4538 31384 4570 31416
rect 4606 31384 4638 31416
rect 4674 31384 4706 31416
rect 4742 31384 4774 31416
rect 4810 31384 4842 31416
rect 4878 31384 4910 31416
rect 4946 31384 4978 31416
rect 5014 31384 5046 31416
rect 5082 31384 5114 31416
rect 5150 31384 5182 31416
rect 5218 31384 5250 31416
rect 5286 31384 5318 31416
rect 5354 31384 5386 31416
rect 5422 31384 5454 31416
rect 5490 31384 5522 31416
rect 5558 31384 5590 31416
rect 5626 31384 5658 31416
rect 5694 31384 5726 31416
rect 5762 31384 5794 31416
rect 5830 31384 5862 31416
rect 5898 31384 5930 31416
rect 5966 31384 5998 31416
rect 6034 31384 6066 31416
rect 6102 31384 6134 31416
rect 6170 31384 6202 31416
rect 6238 31384 6270 31416
rect 6306 31384 6338 31416
rect 6374 31384 6406 31416
rect 6442 31384 6474 31416
rect 6510 31384 6542 31416
rect 6578 31384 6610 31416
rect 6646 31384 6678 31416
rect 6714 31384 6746 31416
rect 6782 31384 6814 31416
rect 6850 31384 6882 31416
rect 6918 31384 6950 31416
rect 6986 31384 7018 31416
rect 7054 31384 7086 31416
rect 7122 31384 7154 31416
rect 7190 31384 7222 31416
rect 7258 31384 7290 31416
rect 7326 31384 7358 31416
rect 7394 31384 7426 31416
rect 7462 31384 7494 31416
rect 7530 31384 7562 31416
rect 7598 31384 7630 31416
rect 7666 31384 7698 31416
rect 7734 31384 7766 31416
rect 7802 31384 7834 31416
rect 7870 31384 7902 31416
rect 7938 31384 7970 31416
rect 8006 31384 8038 31416
rect 8074 31384 8106 31416
rect 8142 31384 8174 31416
rect 8210 31384 8242 31416
rect 8278 31384 8310 31416
rect 8346 31384 8378 31416
rect 8414 31384 8446 31416
rect 8482 31384 8514 31416
rect 8550 31384 8582 31416
rect 8618 31384 8650 31416
rect 8686 31384 8718 31416
rect 8754 31384 8786 31416
rect 8822 31384 8854 31416
rect 8890 31384 8922 31416
rect 8958 31384 8990 31416
rect 9026 31384 9058 31416
rect 9094 31384 9126 31416
rect 9162 31384 9194 31416
rect 9230 31384 9262 31416
rect 9298 31384 9330 31416
rect 9366 31384 9398 31416
rect 9434 31384 9466 31416
rect 9502 31384 9534 31416
rect 9570 31384 9602 31416
rect 9638 31384 9670 31416
rect 9706 31384 9738 31416
rect 9774 31384 9806 31416
rect 9842 31384 9874 31416
rect 9910 31384 9942 31416
rect 9978 31384 10010 31416
rect 10046 31384 10078 31416
rect 10114 31384 10146 31416
rect 10182 31384 10214 31416
rect 10250 31384 10282 31416
rect 10318 31384 10350 31416
rect 10386 31384 10418 31416
rect 10454 31384 10486 31416
rect 10522 31384 10554 31416
rect 10590 31384 10622 31416
rect 10658 31384 10690 31416
rect 10726 31384 10758 31416
rect 10794 31384 10826 31416
rect 10862 31384 10894 31416
rect 10930 31384 10962 31416
rect 10998 31384 11030 31416
rect 11066 31384 11098 31416
rect 11134 31384 11166 31416
rect 11202 31384 11234 31416
rect 11270 31384 11302 31416
rect 11338 31384 11370 31416
rect 11406 31384 11438 31416
rect 11474 31384 11506 31416
rect 11542 31384 11574 31416
rect 11610 31384 11642 31416
rect 11678 31384 11710 31416
rect 11746 31384 11778 31416
rect 11814 31384 11846 31416
rect 11882 31384 11914 31416
rect 11950 31384 11982 31416
rect 12018 31384 12050 31416
rect 12086 31384 12118 31416
rect 12154 31384 12186 31416
rect 12222 31384 12254 31416
rect 12290 31384 12322 31416
rect 12358 31384 12390 31416
rect 12426 31384 12458 31416
rect 12494 31384 12526 31416
rect 12562 31384 12594 31416
rect 12630 31384 12662 31416
rect 12698 31384 12730 31416
rect 12766 31384 12798 31416
rect 12834 31384 12866 31416
rect 12902 31384 12934 31416
rect 12970 31384 13002 31416
rect 13038 31384 13070 31416
rect 13106 31384 13138 31416
rect 13174 31384 13206 31416
rect 13242 31384 13274 31416
rect 13310 31384 13342 31416
rect 13378 31384 13410 31416
rect 13446 31384 13478 31416
rect 13514 31384 13546 31416
rect 13582 31384 13614 31416
rect 13650 31384 13682 31416
rect 13718 31384 13750 31416
rect 13786 31384 13818 31416
rect 13854 31384 13886 31416
rect 13922 31384 13954 31416
rect 13990 31384 14022 31416
rect 14058 31384 14090 31416
rect 14126 31384 14158 31416
rect 14194 31384 14226 31416
rect 14262 31384 14294 31416
rect 14330 31384 14362 31416
rect 14398 31384 14430 31416
rect 14466 31384 14498 31416
rect 14534 31384 14566 31416
rect 14602 31384 14634 31416
rect 14670 31384 14702 31416
rect 14738 31384 14770 31416
rect 14806 31384 14838 31416
rect 14874 31384 14906 31416
rect 14942 31384 14974 31416
rect 15010 31384 15042 31416
rect 15078 31384 15110 31416
rect 15146 31384 15178 31416
rect 15214 31384 15246 31416
rect 15282 31384 15314 31416
rect 15350 31384 15382 31416
rect 15442 31384 15474 31416
rect 15510 31384 15542 31416
rect 15578 31384 15610 31416
rect 15646 31384 15678 31416
rect 15714 31384 15746 31416
rect 15782 31384 15814 31416
rect 15850 31384 15882 31416
rect 15918 31384 15950 31416
rect 136 27939 168 27971
rect 208 27939 240 27971
rect 280 27939 312 27971
rect 352 27939 384 27971
rect 424 27939 456 27971
rect 496 27939 528 27971
rect 568 27939 600 27971
rect 640 27939 672 27971
rect 712 27939 744 27971
rect 784 27939 816 27971
rect 856 27939 888 27971
rect 928 27939 960 27971
rect 1000 27939 1032 27971
rect 1072 27939 1104 27971
rect 1144 27939 1176 27971
rect 1216 27939 1248 27971
rect 1288 27939 1320 27971
rect 1360 27939 1392 27971
rect 1432 27939 1464 27971
rect 1504 27939 1536 27971
rect 1576 27939 1608 27971
rect 1648 27939 1680 27971
rect 1720 27939 1752 27971
rect 1792 27939 1824 27971
rect 1864 27939 1896 27971
rect 1936 27939 1968 27971
rect 2008 27939 2040 27971
rect 2080 27939 2112 27971
rect 2152 27939 2184 27971
rect 2224 27939 2256 27971
rect 2296 27939 2328 27971
rect 2368 27939 2400 27971
rect 2440 27939 2472 27971
rect 2512 27939 2544 27971
rect 2584 27939 2616 27971
rect 2656 27939 2688 27971
rect 2728 27939 2760 27971
rect 2800 27939 2832 27971
rect 2872 27939 2904 27971
rect 2944 27939 2976 27971
rect 3016 27939 3048 27971
rect 3088 27939 3120 27971
rect 3160 27939 3192 27971
rect 3232 27939 3264 27971
rect 3304 27939 3336 27971
rect 3376 27939 3408 27971
rect 3448 27939 3480 27971
rect 3520 27939 3552 27971
rect 3592 27939 3624 27971
rect 3664 27939 3696 27971
rect 3736 27939 3768 27971
rect 3808 27939 3840 27971
rect 3880 27939 3912 27971
rect 3952 27939 3984 27971
rect 4024 27939 4056 27971
rect 4096 27939 4128 27971
rect 4168 27939 4200 27971
rect 4240 27939 4272 27971
rect 4312 27939 4344 27971
rect 4384 27939 4416 27971
rect 4456 27939 4488 27971
rect 4528 27939 4560 27971
rect 4600 27939 4632 27971
rect 4672 27939 4704 27971
rect 4744 27939 4776 27971
rect 4816 27939 4848 27971
rect 4888 27939 4920 27971
rect 4960 27939 4992 27971
rect 5032 27939 5064 27971
rect 5104 27939 5136 27971
rect 5176 27939 5208 27971
rect 5248 27939 5280 27971
rect 5320 27939 5352 27971
rect 5392 27939 5424 27971
rect 5464 27939 5496 27971
rect 5536 27939 5568 27971
rect 5608 27939 5640 27971
rect 5680 27939 5712 27971
rect 5752 27939 5784 27971
rect 5824 27939 5856 27971
rect 5896 27939 5928 27971
rect 5968 27939 6000 27971
rect 6040 27939 6072 27971
rect 6112 27939 6144 27971
rect 6184 27939 6216 27971
rect 6256 27939 6288 27971
rect 6328 27939 6360 27971
rect 6400 27939 6432 27971
rect 6472 27939 6504 27971
rect 6544 27939 6576 27971
rect 6616 27939 6648 27971
rect 6688 27939 6720 27971
rect 6760 27939 6792 27971
rect 6832 27939 6864 27971
rect 6904 27939 6936 27971
rect 6976 27939 7008 27971
rect 7048 27939 7080 27971
rect 7120 27939 7152 27971
rect 7192 27939 7224 27971
rect 7264 27939 7296 27971
rect 7336 27939 7368 27971
rect 7408 27939 7440 27971
rect 7480 27939 7512 27971
rect 7552 27939 7584 27971
rect 7624 27939 7656 27971
rect 7696 27939 7728 27971
rect 7768 27939 7800 27971
rect 7840 27939 7872 27971
rect 7912 27939 7944 27971
rect 7984 27939 8016 27971
rect 8056 27939 8088 27971
rect 8128 27939 8160 27971
rect 8200 27939 8232 27971
rect 8272 27939 8304 27971
rect 8344 27939 8376 27971
rect 8416 27939 8448 27971
rect 8488 27939 8520 27971
rect 8560 27939 8592 27971
rect 8632 27939 8664 27971
rect 8704 27939 8736 27971
rect 8776 27939 8808 27971
rect 8848 27939 8880 27971
rect 8920 27939 8952 27971
rect 8992 27939 9024 27971
rect 9064 27939 9096 27971
rect 9136 27939 9168 27971
rect 9208 27939 9240 27971
rect 9280 27939 9312 27971
rect 9352 27939 9384 27971
rect 9424 27939 9456 27971
rect 9496 27939 9528 27971
rect 9568 27939 9600 27971
rect 9640 27939 9672 27971
rect 9712 27939 9744 27971
rect 9784 27939 9816 27971
rect 9856 27939 9888 27971
rect 9928 27939 9960 27971
rect 10000 27939 10032 27971
rect 10072 27939 10104 27971
rect 10144 27939 10176 27971
rect 10216 27939 10248 27971
rect 10288 27939 10320 27971
rect 10360 27939 10392 27971
rect 10432 27939 10464 27971
rect 10504 27939 10536 27971
rect 10576 27939 10608 27971
rect 10648 27939 10680 27971
rect 10720 27939 10752 27971
rect 10792 27939 10824 27971
rect 10864 27939 10896 27971
rect 10936 27939 10968 27971
rect 11008 27939 11040 27971
rect 11080 27939 11112 27971
rect 11152 27939 11184 27971
rect 11224 27939 11256 27971
rect 11296 27939 11328 27971
rect 11368 27939 11400 27971
rect 11440 27939 11472 27971
rect 11512 27939 11544 27971
rect 11584 27939 11616 27971
rect 11656 27939 11688 27971
rect 11728 27939 11760 27971
rect 11800 27939 11832 27971
rect 11872 27939 11904 27971
rect 11944 27939 11976 27971
rect 12016 27939 12048 27971
rect 12088 27939 12120 27971
rect 12160 27939 12192 27971
rect 12232 27939 12264 27971
rect 12304 27939 12336 27971
rect 12376 27939 12408 27971
rect 12448 27939 12480 27971
rect 12520 27939 12552 27971
rect 12592 27939 12624 27971
rect 12664 27939 12696 27971
rect 12736 27939 12768 27971
rect 12808 27939 12840 27971
rect 12880 27939 12912 27971
rect 12952 27939 12984 27971
rect 13024 27939 13056 27971
rect 13096 27939 13128 27971
rect 13168 27939 13200 27971
rect 13240 27939 13272 27971
rect 13312 27939 13344 27971
rect 13384 27939 13416 27971
rect 13456 27939 13488 27971
rect 13528 27939 13560 27971
rect 13600 27939 13632 27971
rect 13672 27939 13704 27971
rect 13744 27939 13776 27971
rect 13816 27939 13848 27971
rect 13888 27939 13920 27971
rect 13960 27939 13992 27971
rect 14032 27939 14064 27971
rect 14104 27939 14136 27971
rect 14176 27939 14208 27971
rect 14248 27939 14280 27971
rect 14320 27939 14352 27971
rect 14392 27939 14424 27971
rect 14464 27939 14496 27971
rect 14536 27939 14568 27971
rect 14608 27939 14640 27971
rect 14680 27939 14712 27971
rect 14752 27939 14784 27971
rect 14824 27939 14856 27971
rect 14896 27939 14928 27971
rect 14968 27939 15000 27971
rect 15040 27939 15072 27971
rect 15112 27939 15144 27971
rect 15184 27939 15216 27971
rect 15256 27939 15288 27971
rect 15328 27939 15360 27971
rect 15400 27939 15432 27971
rect 15472 27939 15504 27971
rect 15544 27939 15576 27971
rect 15616 27939 15648 27971
rect 15688 27939 15720 27971
rect 15760 27939 15792 27971
rect 15832 27939 15864 27971
rect 15904 27939 15936 27971
rect 64 27867 96 27899
rect 136 27867 168 27899
rect 208 27867 240 27899
rect 280 27867 312 27899
rect 352 27867 384 27899
rect 424 27867 456 27899
rect 496 27867 528 27899
rect 568 27867 600 27899
rect 640 27867 672 27899
rect 712 27867 744 27899
rect 784 27867 816 27899
rect 856 27867 888 27899
rect 928 27867 960 27899
rect 1000 27867 1032 27899
rect 1072 27867 1104 27899
rect 1144 27867 1176 27899
rect 1216 27867 1248 27899
rect 1288 27867 1320 27899
rect 1360 27867 1392 27899
rect 1432 27867 1464 27899
rect 1504 27867 1536 27899
rect 1576 27867 1608 27899
rect 1648 27867 1680 27899
rect 1720 27867 1752 27899
rect 1792 27867 1824 27899
rect 1864 27867 1896 27899
rect 1936 27867 1968 27899
rect 2008 27867 2040 27899
rect 2080 27867 2112 27899
rect 2152 27867 2184 27899
rect 2224 27867 2256 27899
rect 2296 27867 2328 27899
rect 2368 27867 2400 27899
rect 2440 27867 2472 27899
rect 2512 27867 2544 27899
rect 2584 27867 2616 27899
rect 2656 27867 2688 27899
rect 2728 27867 2760 27899
rect 2800 27867 2832 27899
rect 2872 27867 2904 27899
rect 2944 27867 2976 27899
rect 3016 27867 3048 27899
rect 3088 27867 3120 27899
rect 3160 27867 3192 27899
rect 3232 27867 3264 27899
rect 3304 27867 3336 27899
rect 3376 27867 3408 27899
rect 3448 27867 3480 27899
rect 3520 27867 3552 27899
rect 3592 27867 3624 27899
rect 3664 27867 3696 27899
rect 3736 27867 3768 27899
rect 3808 27867 3840 27899
rect 3880 27867 3912 27899
rect 3952 27867 3984 27899
rect 4024 27867 4056 27899
rect 4096 27867 4128 27899
rect 4168 27867 4200 27899
rect 4240 27867 4272 27899
rect 4312 27867 4344 27899
rect 4384 27867 4416 27899
rect 4456 27867 4488 27899
rect 4528 27867 4560 27899
rect 4600 27867 4632 27899
rect 4672 27867 4704 27899
rect 4744 27867 4776 27899
rect 4816 27867 4848 27899
rect 4888 27867 4920 27899
rect 4960 27867 4992 27899
rect 5032 27867 5064 27899
rect 5104 27867 5136 27899
rect 5176 27867 5208 27899
rect 5248 27867 5280 27899
rect 5320 27867 5352 27899
rect 5392 27867 5424 27899
rect 5464 27867 5496 27899
rect 5536 27867 5568 27899
rect 5608 27867 5640 27899
rect 5680 27867 5712 27899
rect 5752 27867 5784 27899
rect 5824 27867 5856 27899
rect 5896 27867 5928 27899
rect 5968 27867 6000 27899
rect 6040 27867 6072 27899
rect 6112 27867 6144 27899
rect 6184 27867 6216 27899
rect 6256 27867 6288 27899
rect 6328 27867 6360 27899
rect 6400 27867 6432 27899
rect 6472 27867 6504 27899
rect 6544 27867 6576 27899
rect 6616 27867 6648 27899
rect 6688 27867 6720 27899
rect 6760 27867 6792 27899
rect 6832 27867 6864 27899
rect 6904 27867 6936 27899
rect 6976 27867 7008 27899
rect 7048 27867 7080 27899
rect 7120 27867 7152 27899
rect 7192 27867 7224 27899
rect 7264 27867 7296 27899
rect 7336 27867 7368 27899
rect 7408 27867 7440 27899
rect 7480 27867 7512 27899
rect 7552 27867 7584 27899
rect 7624 27867 7656 27899
rect 7696 27867 7728 27899
rect 7768 27867 7800 27899
rect 7840 27867 7872 27899
rect 7912 27867 7944 27899
rect 7984 27867 8016 27899
rect 8056 27867 8088 27899
rect 8128 27867 8160 27899
rect 8200 27867 8232 27899
rect 8272 27867 8304 27899
rect 8344 27867 8376 27899
rect 8416 27867 8448 27899
rect 8488 27867 8520 27899
rect 8560 27867 8592 27899
rect 8632 27867 8664 27899
rect 8704 27867 8736 27899
rect 8776 27867 8808 27899
rect 8848 27867 8880 27899
rect 8920 27867 8952 27899
rect 8992 27867 9024 27899
rect 9064 27867 9096 27899
rect 9136 27867 9168 27899
rect 9208 27867 9240 27899
rect 9280 27867 9312 27899
rect 9352 27867 9384 27899
rect 9424 27867 9456 27899
rect 9496 27867 9528 27899
rect 9568 27867 9600 27899
rect 9640 27867 9672 27899
rect 9712 27867 9744 27899
rect 9784 27867 9816 27899
rect 9856 27867 9888 27899
rect 9928 27867 9960 27899
rect 10000 27867 10032 27899
rect 10072 27867 10104 27899
rect 10144 27867 10176 27899
rect 10216 27867 10248 27899
rect 10288 27867 10320 27899
rect 10360 27867 10392 27899
rect 10432 27867 10464 27899
rect 10504 27867 10536 27899
rect 10576 27867 10608 27899
rect 10648 27867 10680 27899
rect 10720 27867 10752 27899
rect 10792 27867 10824 27899
rect 10864 27867 10896 27899
rect 10936 27867 10968 27899
rect 11008 27867 11040 27899
rect 11080 27867 11112 27899
rect 11152 27867 11184 27899
rect 11224 27867 11256 27899
rect 11296 27867 11328 27899
rect 11368 27867 11400 27899
rect 11440 27867 11472 27899
rect 11512 27867 11544 27899
rect 11584 27867 11616 27899
rect 11656 27867 11688 27899
rect 11728 27867 11760 27899
rect 11800 27867 11832 27899
rect 11872 27867 11904 27899
rect 11944 27867 11976 27899
rect 12016 27867 12048 27899
rect 12088 27867 12120 27899
rect 12160 27867 12192 27899
rect 12232 27867 12264 27899
rect 12304 27867 12336 27899
rect 12376 27867 12408 27899
rect 12448 27867 12480 27899
rect 12520 27867 12552 27899
rect 12592 27867 12624 27899
rect 12664 27867 12696 27899
rect 12736 27867 12768 27899
rect 12808 27867 12840 27899
rect 12880 27867 12912 27899
rect 12952 27867 12984 27899
rect 13024 27867 13056 27899
rect 13096 27867 13128 27899
rect 13168 27867 13200 27899
rect 13240 27867 13272 27899
rect 13312 27867 13344 27899
rect 13384 27867 13416 27899
rect 13456 27867 13488 27899
rect 13528 27867 13560 27899
rect 13600 27867 13632 27899
rect 13672 27867 13704 27899
rect 13744 27867 13776 27899
rect 13816 27867 13848 27899
rect 13888 27867 13920 27899
rect 13960 27867 13992 27899
rect 14032 27867 14064 27899
rect 14104 27867 14136 27899
rect 14176 27867 14208 27899
rect 14248 27867 14280 27899
rect 14320 27867 14352 27899
rect 14392 27867 14424 27899
rect 14464 27867 14496 27899
rect 14536 27867 14568 27899
rect 14608 27867 14640 27899
rect 14680 27867 14712 27899
rect 14752 27867 14784 27899
rect 14824 27867 14856 27899
rect 14896 27867 14928 27899
rect 14968 27867 15000 27899
rect 15040 27867 15072 27899
rect 15112 27867 15144 27899
rect 15184 27867 15216 27899
rect 15256 27867 15288 27899
rect 15328 27867 15360 27899
rect 15400 27867 15432 27899
rect 15472 27867 15504 27899
rect 15544 27867 15576 27899
rect 15616 27867 15648 27899
rect 15688 27867 15720 27899
rect 15760 27867 15792 27899
rect 15832 27867 15864 27899
rect 15904 27867 15936 27899
rect 64 27795 96 27827
rect 136 27795 168 27827
rect 208 27795 240 27827
rect 280 27795 312 27827
rect 352 27795 384 27827
rect 424 27795 456 27827
rect 496 27795 528 27827
rect 568 27795 600 27827
rect 640 27795 672 27827
rect 712 27795 744 27827
rect 784 27795 816 27827
rect 856 27795 888 27827
rect 928 27795 960 27827
rect 1000 27795 1032 27827
rect 1072 27795 1104 27827
rect 1144 27795 1176 27827
rect 1216 27795 1248 27827
rect 1288 27795 1320 27827
rect 1360 27795 1392 27827
rect 1432 27795 1464 27827
rect 1504 27795 1536 27827
rect 1576 27795 1608 27827
rect 1648 27795 1680 27827
rect 1720 27795 1752 27827
rect 1792 27795 1824 27827
rect 1864 27795 1896 27827
rect 1936 27795 1968 27827
rect 2008 27795 2040 27827
rect 2080 27795 2112 27827
rect 2152 27795 2184 27827
rect 2224 27795 2256 27827
rect 2296 27795 2328 27827
rect 2368 27795 2400 27827
rect 2440 27795 2472 27827
rect 2512 27795 2544 27827
rect 2584 27795 2616 27827
rect 2656 27795 2688 27827
rect 2728 27795 2760 27827
rect 2800 27795 2832 27827
rect 2872 27795 2904 27827
rect 2944 27795 2976 27827
rect 3016 27795 3048 27827
rect 3088 27795 3120 27827
rect 3160 27795 3192 27827
rect 3232 27795 3264 27827
rect 3304 27795 3336 27827
rect 3376 27795 3408 27827
rect 3448 27795 3480 27827
rect 3520 27795 3552 27827
rect 3592 27795 3624 27827
rect 3664 27795 3696 27827
rect 3736 27795 3768 27827
rect 3808 27795 3840 27827
rect 3880 27795 3912 27827
rect 3952 27795 3984 27827
rect 4024 27795 4056 27827
rect 4096 27795 4128 27827
rect 4168 27795 4200 27827
rect 4240 27795 4272 27827
rect 4312 27795 4344 27827
rect 4384 27795 4416 27827
rect 4456 27795 4488 27827
rect 4528 27795 4560 27827
rect 4600 27795 4632 27827
rect 4672 27795 4704 27827
rect 4744 27795 4776 27827
rect 4816 27795 4848 27827
rect 4888 27795 4920 27827
rect 4960 27795 4992 27827
rect 5032 27795 5064 27827
rect 5104 27795 5136 27827
rect 5176 27795 5208 27827
rect 5248 27795 5280 27827
rect 5320 27795 5352 27827
rect 5392 27795 5424 27827
rect 5464 27795 5496 27827
rect 5536 27795 5568 27827
rect 5608 27795 5640 27827
rect 5680 27795 5712 27827
rect 5752 27795 5784 27827
rect 5824 27795 5856 27827
rect 5896 27795 5928 27827
rect 5968 27795 6000 27827
rect 6040 27795 6072 27827
rect 6112 27795 6144 27827
rect 6184 27795 6216 27827
rect 6256 27795 6288 27827
rect 6328 27795 6360 27827
rect 6400 27795 6432 27827
rect 6472 27795 6504 27827
rect 6544 27795 6576 27827
rect 6616 27795 6648 27827
rect 6688 27795 6720 27827
rect 6760 27795 6792 27827
rect 6832 27795 6864 27827
rect 6904 27795 6936 27827
rect 6976 27795 7008 27827
rect 7048 27795 7080 27827
rect 7120 27795 7152 27827
rect 7192 27795 7224 27827
rect 7264 27795 7296 27827
rect 7336 27795 7368 27827
rect 7408 27795 7440 27827
rect 7480 27795 7512 27827
rect 7552 27795 7584 27827
rect 7624 27795 7656 27827
rect 7696 27795 7728 27827
rect 7768 27795 7800 27827
rect 7840 27795 7872 27827
rect 7912 27795 7944 27827
rect 7984 27795 8016 27827
rect 8056 27795 8088 27827
rect 8128 27795 8160 27827
rect 8200 27795 8232 27827
rect 8272 27795 8304 27827
rect 8344 27795 8376 27827
rect 8416 27795 8448 27827
rect 8488 27795 8520 27827
rect 8560 27795 8592 27827
rect 8632 27795 8664 27827
rect 8704 27795 8736 27827
rect 8776 27795 8808 27827
rect 8848 27795 8880 27827
rect 8920 27795 8952 27827
rect 8992 27795 9024 27827
rect 9064 27795 9096 27827
rect 9136 27795 9168 27827
rect 9208 27795 9240 27827
rect 9280 27795 9312 27827
rect 9352 27795 9384 27827
rect 9424 27795 9456 27827
rect 9496 27795 9528 27827
rect 9568 27795 9600 27827
rect 9640 27795 9672 27827
rect 9712 27795 9744 27827
rect 9784 27795 9816 27827
rect 9856 27795 9888 27827
rect 9928 27795 9960 27827
rect 10000 27795 10032 27827
rect 10072 27795 10104 27827
rect 10144 27795 10176 27827
rect 10216 27795 10248 27827
rect 10288 27795 10320 27827
rect 10360 27795 10392 27827
rect 10432 27795 10464 27827
rect 10504 27795 10536 27827
rect 10576 27795 10608 27827
rect 10648 27795 10680 27827
rect 10720 27795 10752 27827
rect 10792 27795 10824 27827
rect 10864 27795 10896 27827
rect 10936 27795 10968 27827
rect 11008 27795 11040 27827
rect 11080 27795 11112 27827
rect 11152 27795 11184 27827
rect 11224 27795 11256 27827
rect 11296 27795 11328 27827
rect 11368 27795 11400 27827
rect 11440 27795 11472 27827
rect 11512 27795 11544 27827
rect 11584 27795 11616 27827
rect 11656 27795 11688 27827
rect 11728 27795 11760 27827
rect 11800 27795 11832 27827
rect 11872 27795 11904 27827
rect 11944 27795 11976 27827
rect 12016 27795 12048 27827
rect 12088 27795 12120 27827
rect 12160 27795 12192 27827
rect 12232 27795 12264 27827
rect 12304 27795 12336 27827
rect 12376 27795 12408 27827
rect 12448 27795 12480 27827
rect 12520 27795 12552 27827
rect 12592 27795 12624 27827
rect 12664 27795 12696 27827
rect 12736 27795 12768 27827
rect 12808 27795 12840 27827
rect 12880 27795 12912 27827
rect 12952 27795 12984 27827
rect 13024 27795 13056 27827
rect 13096 27795 13128 27827
rect 13168 27795 13200 27827
rect 13240 27795 13272 27827
rect 13312 27795 13344 27827
rect 13384 27795 13416 27827
rect 13456 27795 13488 27827
rect 13528 27795 13560 27827
rect 13600 27795 13632 27827
rect 13672 27795 13704 27827
rect 13744 27795 13776 27827
rect 13816 27795 13848 27827
rect 13888 27795 13920 27827
rect 13960 27795 13992 27827
rect 14032 27795 14064 27827
rect 14104 27795 14136 27827
rect 14176 27795 14208 27827
rect 14248 27795 14280 27827
rect 14320 27795 14352 27827
rect 14392 27795 14424 27827
rect 14464 27795 14496 27827
rect 14536 27795 14568 27827
rect 14608 27795 14640 27827
rect 14680 27795 14712 27827
rect 14752 27795 14784 27827
rect 14824 27795 14856 27827
rect 14896 27795 14928 27827
rect 14968 27795 15000 27827
rect 15040 27795 15072 27827
rect 15112 27795 15144 27827
rect 15184 27795 15216 27827
rect 15256 27795 15288 27827
rect 15328 27795 15360 27827
rect 15400 27795 15432 27827
rect 15472 27795 15504 27827
rect 15544 27795 15576 27827
rect 15616 27795 15648 27827
rect 15688 27795 15720 27827
rect 15760 27795 15792 27827
rect 15832 27795 15864 27827
rect 15904 27795 15936 27827
rect 64 27723 96 27755
rect 136 27723 168 27755
rect 208 27723 240 27755
rect 280 27723 312 27755
rect 352 27723 384 27755
rect 424 27723 456 27755
rect 496 27723 528 27755
rect 568 27723 600 27755
rect 640 27723 672 27755
rect 712 27723 744 27755
rect 784 27723 816 27755
rect 856 27723 888 27755
rect 928 27723 960 27755
rect 1000 27723 1032 27755
rect 1072 27723 1104 27755
rect 1144 27723 1176 27755
rect 1216 27723 1248 27755
rect 1288 27723 1320 27755
rect 1360 27723 1392 27755
rect 1432 27723 1464 27755
rect 1504 27723 1536 27755
rect 1576 27723 1608 27755
rect 1648 27723 1680 27755
rect 1720 27723 1752 27755
rect 1792 27723 1824 27755
rect 1864 27723 1896 27755
rect 1936 27723 1968 27755
rect 2008 27723 2040 27755
rect 2080 27723 2112 27755
rect 2152 27723 2184 27755
rect 2224 27723 2256 27755
rect 2296 27723 2328 27755
rect 2368 27723 2400 27755
rect 2440 27723 2472 27755
rect 2512 27723 2544 27755
rect 2584 27723 2616 27755
rect 2656 27723 2688 27755
rect 2728 27723 2760 27755
rect 2800 27723 2832 27755
rect 2872 27723 2904 27755
rect 2944 27723 2976 27755
rect 3016 27723 3048 27755
rect 3088 27723 3120 27755
rect 3160 27723 3192 27755
rect 3232 27723 3264 27755
rect 3304 27723 3336 27755
rect 3376 27723 3408 27755
rect 3448 27723 3480 27755
rect 3520 27723 3552 27755
rect 3592 27723 3624 27755
rect 3664 27723 3696 27755
rect 3736 27723 3768 27755
rect 3808 27723 3840 27755
rect 3880 27723 3912 27755
rect 3952 27723 3984 27755
rect 4024 27723 4056 27755
rect 4096 27723 4128 27755
rect 4168 27723 4200 27755
rect 4240 27723 4272 27755
rect 4312 27723 4344 27755
rect 4384 27723 4416 27755
rect 4456 27723 4488 27755
rect 4528 27723 4560 27755
rect 4600 27723 4632 27755
rect 4672 27723 4704 27755
rect 4744 27723 4776 27755
rect 4816 27723 4848 27755
rect 4888 27723 4920 27755
rect 4960 27723 4992 27755
rect 5032 27723 5064 27755
rect 5104 27723 5136 27755
rect 5176 27723 5208 27755
rect 5248 27723 5280 27755
rect 5320 27723 5352 27755
rect 5392 27723 5424 27755
rect 5464 27723 5496 27755
rect 5536 27723 5568 27755
rect 5608 27723 5640 27755
rect 5680 27723 5712 27755
rect 5752 27723 5784 27755
rect 5824 27723 5856 27755
rect 5896 27723 5928 27755
rect 5968 27723 6000 27755
rect 6040 27723 6072 27755
rect 6112 27723 6144 27755
rect 6184 27723 6216 27755
rect 6256 27723 6288 27755
rect 6328 27723 6360 27755
rect 6400 27723 6432 27755
rect 6472 27723 6504 27755
rect 6544 27723 6576 27755
rect 6616 27723 6648 27755
rect 6688 27723 6720 27755
rect 6760 27723 6792 27755
rect 6832 27723 6864 27755
rect 6904 27723 6936 27755
rect 6976 27723 7008 27755
rect 7048 27723 7080 27755
rect 7120 27723 7152 27755
rect 7192 27723 7224 27755
rect 7264 27723 7296 27755
rect 7336 27723 7368 27755
rect 7408 27723 7440 27755
rect 7480 27723 7512 27755
rect 7552 27723 7584 27755
rect 7624 27723 7656 27755
rect 7696 27723 7728 27755
rect 7768 27723 7800 27755
rect 7840 27723 7872 27755
rect 7912 27723 7944 27755
rect 7984 27723 8016 27755
rect 8056 27723 8088 27755
rect 8128 27723 8160 27755
rect 8200 27723 8232 27755
rect 8272 27723 8304 27755
rect 8344 27723 8376 27755
rect 8416 27723 8448 27755
rect 8488 27723 8520 27755
rect 8560 27723 8592 27755
rect 8632 27723 8664 27755
rect 8704 27723 8736 27755
rect 8776 27723 8808 27755
rect 8848 27723 8880 27755
rect 8920 27723 8952 27755
rect 8992 27723 9024 27755
rect 9064 27723 9096 27755
rect 9136 27723 9168 27755
rect 9208 27723 9240 27755
rect 9280 27723 9312 27755
rect 9352 27723 9384 27755
rect 9424 27723 9456 27755
rect 9496 27723 9528 27755
rect 9568 27723 9600 27755
rect 9640 27723 9672 27755
rect 9712 27723 9744 27755
rect 9784 27723 9816 27755
rect 9856 27723 9888 27755
rect 9928 27723 9960 27755
rect 10000 27723 10032 27755
rect 10072 27723 10104 27755
rect 10144 27723 10176 27755
rect 10216 27723 10248 27755
rect 10288 27723 10320 27755
rect 10360 27723 10392 27755
rect 10432 27723 10464 27755
rect 10504 27723 10536 27755
rect 10576 27723 10608 27755
rect 10648 27723 10680 27755
rect 10720 27723 10752 27755
rect 10792 27723 10824 27755
rect 10864 27723 10896 27755
rect 10936 27723 10968 27755
rect 11008 27723 11040 27755
rect 11080 27723 11112 27755
rect 11152 27723 11184 27755
rect 11224 27723 11256 27755
rect 11296 27723 11328 27755
rect 11368 27723 11400 27755
rect 11440 27723 11472 27755
rect 11512 27723 11544 27755
rect 11584 27723 11616 27755
rect 11656 27723 11688 27755
rect 11728 27723 11760 27755
rect 11800 27723 11832 27755
rect 11872 27723 11904 27755
rect 11944 27723 11976 27755
rect 12016 27723 12048 27755
rect 12088 27723 12120 27755
rect 12160 27723 12192 27755
rect 12232 27723 12264 27755
rect 12304 27723 12336 27755
rect 12376 27723 12408 27755
rect 12448 27723 12480 27755
rect 12520 27723 12552 27755
rect 12592 27723 12624 27755
rect 12664 27723 12696 27755
rect 12736 27723 12768 27755
rect 12808 27723 12840 27755
rect 12880 27723 12912 27755
rect 12952 27723 12984 27755
rect 13024 27723 13056 27755
rect 13096 27723 13128 27755
rect 13168 27723 13200 27755
rect 13240 27723 13272 27755
rect 13312 27723 13344 27755
rect 13384 27723 13416 27755
rect 13456 27723 13488 27755
rect 13528 27723 13560 27755
rect 13600 27723 13632 27755
rect 13672 27723 13704 27755
rect 13744 27723 13776 27755
rect 13816 27723 13848 27755
rect 13888 27723 13920 27755
rect 13960 27723 13992 27755
rect 14032 27723 14064 27755
rect 14104 27723 14136 27755
rect 14176 27723 14208 27755
rect 14248 27723 14280 27755
rect 14320 27723 14352 27755
rect 14392 27723 14424 27755
rect 14464 27723 14496 27755
rect 14536 27723 14568 27755
rect 14608 27723 14640 27755
rect 14680 27723 14712 27755
rect 14752 27723 14784 27755
rect 14824 27723 14856 27755
rect 14896 27723 14928 27755
rect 14968 27723 15000 27755
rect 15040 27723 15072 27755
rect 15112 27723 15144 27755
rect 15184 27723 15216 27755
rect 15256 27723 15288 27755
rect 15328 27723 15360 27755
rect 15400 27723 15432 27755
rect 15472 27723 15504 27755
rect 15544 27723 15576 27755
rect 15616 27723 15648 27755
rect 15688 27723 15720 27755
rect 15760 27723 15792 27755
rect 15832 27723 15864 27755
rect 15904 27723 15936 27755
rect 64 27651 96 27683
rect 136 27651 168 27683
rect 208 27651 240 27683
rect 280 27651 312 27683
rect 352 27651 384 27683
rect 424 27651 456 27683
rect 496 27651 528 27683
rect 568 27651 600 27683
rect 640 27651 672 27683
rect 712 27651 744 27683
rect 784 27651 816 27683
rect 856 27651 888 27683
rect 928 27651 960 27683
rect 1000 27651 1032 27683
rect 1072 27651 1104 27683
rect 1144 27651 1176 27683
rect 1216 27651 1248 27683
rect 1288 27651 1320 27683
rect 1360 27651 1392 27683
rect 1432 27651 1464 27683
rect 1504 27651 1536 27683
rect 1576 27651 1608 27683
rect 1648 27651 1680 27683
rect 1720 27651 1752 27683
rect 1792 27651 1824 27683
rect 1864 27651 1896 27683
rect 1936 27651 1968 27683
rect 2008 27651 2040 27683
rect 2080 27651 2112 27683
rect 2152 27651 2184 27683
rect 2224 27651 2256 27683
rect 2296 27651 2328 27683
rect 2368 27651 2400 27683
rect 2440 27651 2472 27683
rect 2512 27651 2544 27683
rect 2584 27651 2616 27683
rect 2656 27651 2688 27683
rect 2728 27651 2760 27683
rect 2800 27651 2832 27683
rect 2872 27651 2904 27683
rect 2944 27651 2976 27683
rect 3016 27651 3048 27683
rect 3088 27651 3120 27683
rect 3160 27651 3192 27683
rect 3232 27651 3264 27683
rect 3304 27651 3336 27683
rect 3376 27651 3408 27683
rect 3448 27651 3480 27683
rect 3520 27651 3552 27683
rect 3592 27651 3624 27683
rect 3664 27651 3696 27683
rect 3736 27651 3768 27683
rect 3808 27651 3840 27683
rect 3880 27651 3912 27683
rect 3952 27651 3984 27683
rect 4024 27651 4056 27683
rect 4096 27651 4128 27683
rect 4168 27651 4200 27683
rect 4240 27651 4272 27683
rect 4312 27651 4344 27683
rect 4384 27651 4416 27683
rect 4456 27651 4488 27683
rect 4528 27651 4560 27683
rect 4600 27651 4632 27683
rect 4672 27651 4704 27683
rect 4744 27651 4776 27683
rect 4816 27651 4848 27683
rect 4888 27651 4920 27683
rect 4960 27651 4992 27683
rect 5032 27651 5064 27683
rect 5104 27651 5136 27683
rect 5176 27651 5208 27683
rect 5248 27651 5280 27683
rect 5320 27651 5352 27683
rect 5392 27651 5424 27683
rect 5464 27651 5496 27683
rect 5536 27651 5568 27683
rect 5608 27651 5640 27683
rect 5680 27651 5712 27683
rect 5752 27651 5784 27683
rect 5824 27651 5856 27683
rect 5896 27651 5928 27683
rect 5968 27651 6000 27683
rect 6040 27651 6072 27683
rect 6112 27651 6144 27683
rect 6184 27651 6216 27683
rect 6256 27651 6288 27683
rect 6328 27651 6360 27683
rect 6400 27651 6432 27683
rect 6472 27651 6504 27683
rect 6544 27651 6576 27683
rect 6616 27651 6648 27683
rect 6688 27651 6720 27683
rect 6760 27651 6792 27683
rect 6832 27651 6864 27683
rect 6904 27651 6936 27683
rect 6976 27651 7008 27683
rect 7048 27651 7080 27683
rect 7120 27651 7152 27683
rect 7192 27651 7224 27683
rect 7264 27651 7296 27683
rect 7336 27651 7368 27683
rect 7408 27651 7440 27683
rect 7480 27651 7512 27683
rect 7552 27651 7584 27683
rect 7624 27651 7656 27683
rect 7696 27651 7728 27683
rect 7768 27651 7800 27683
rect 7840 27651 7872 27683
rect 7912 27651 7944 27683
rect 7984 27651 8016 27683
rect 8056 27651 8088 27683
rect 8128 27651 8160 27683
rect 8200 27651 8232 27683
rect 8272 27651 8304 27683
rect 8344 27651 8376 27683
rect 8416 27651 8448 27683
rect 8488 27651 8520 27683
rect 8560 27651 8592 27683
rect 8632 27651 8664 27683
rect 8704 27651 8736 27683
rect 8776 27651 8808 27683
rect 8848 27651 8880 27683
rect 8920 27651 8952 27683
rect 8992 27651 9024 27683
rect 9064 27651 9096 27683
rect 9136 27651 9168 27683
rect 9208 27651 9240 27683
rect 9280 27651 9312 27683
rect 9352 27651 9384 27683
rect 9424 27651 9456 27683
rect 9496 27651 9528 27683
rect 9568 27651 9600 27683
rect 9640 27651 9672 27683
rect 9712 27651 9744 27683
rect 9784 27651 9816 27683
rect 9856 27651 9888 27683
rect 9928 27651 9960 27683
rect 10000 27651 10032 27683
rect 10072 27651 10104 27683
rect 10144 27651 10176 27683
rect 10216 27651 10248 27683
rect 10288 27651 10320 27683
rect 10360 27651 10392 27683
rect 10432 27651 10464 27683
rect 10504 27651 10536 27683
rect 10576 27651 10608 27683
rect 10648 27651 10680 27683
rect 10720 27651 10752 27683
rect 10792 27651 10824 27683
rect 10864 27651 10896 27683
rect 10936 27651 10968 27683
rect 11008 27651 11040 27683
rect 11080 27651 11112 27683
rect 11152 27651 11184 27683
rect 11224 27651 11256 27683
rect 11296 27651 11328 27683
rect 11368 27651 11400 27683
rect 11440 27651 11472 27683
rect 11512 27651 11544 27683
rect 11584 27651 11616 27683
rect 11656 27651 11688 27683
rect 11728 27651 11760 27683
rect 11800 27651 11832 27683
rect 11872 27651 11904 27683
rect 11944 27651 11976 27683
rect 12016 27651 12048 27683
rect 12088 27651 12120 27683
rect 12160 27651 12192 27683
rect 12232 27651 12264 27683
rect 12304 27651 12336 27683
rect 12376 27651 12408 27683
rect 12448 27651 12480 27683
rect 12520 27651 12552 27683
rect 12592 27651 12624 27683
rect 12664 27651 12696 27683
rect 12736 27651 12768 27683
rect 12808 27651 12840 27683
rect 12880 27651 12912 27683
rect 12952 27651 12984 27683
rect 13024 27651 13056 27683
rect 13096 27651 13128 27683
rect 13168 27651 13200 27683
rect 13240 27651 13272 27683
rect 13312 27651 13344 27683
rect 13384 27651 13416 27683
rect 13456 27651 13488 27683
rect 13528 27651 13560 27683
rect 13600 27651 13632 27683
rect 13672 27651 13704 27683
rect 13744 27651 13776 27683
rect 13816 27651 13848 27683
rect 13888 27651 13920 27683
rect 13960 27651 13992 27683
rect 14032 27651 14064 27683
rect 14104 27651 14136 27683
rect 14176 27651 14208 27683
rect 14248 27651 14280 27683
rect 14320 27651 14352 27683
rect 14392 27651 14424 27683
rect 14464 27651 14496 27683
rect 14536 27651 14568 27683
rect 14608 27651 14640 27683
rect 14680 27651 14712 27683
rect 14752 27651 14784 27683
rect 14824 27651 14856 27683
rect 14896 27651 14928 27683
rect 14968 27651 15000 27683
rect 15040 27651 15072 27683
rect 15112 27651 15144 27683
rect 15184 27651 15216 27683
rect 15256 27651 15288 27683
rect 15328 27651 15360 27683
rect 15400 27651 15432 27683
rect 15472 27651 15504 27683
rect 15544 27651 15576 27683
rect 15616 27651 15648 27683
rect 15688 27651 15720 27683
rect 15760 27651 15792 27683
rect 15832 27651 15864 27683
rect 15904 27651 15936 27683
rect 64 27579 96 27611
rect 136 27579 168 27611
rect 208 27579 240 27611
rect 280 27579 312 27611
rect 352 27579 384 27611
rect 424 27579 456 27611
rect 496 27579 528 27611
rect 568 27579 600 27611
rect 640 27579 672 27611
rect 712 27579 744 27611
rect 784 27579 816 27611
rect 856 27579 888 27611
rect 928 27579 960 27611
rect 1000 27579 1032 27611
rect 1072 27579 1104 27611
rect 1144 27579 1176 27611
rect 1216 27579 1248 27611
rect 1288 27579 1320 27611
rect 1360 27579 1392 27611
rect 1432 27579 1464 27611
rect 1504 27579 1536 27611
rect 1576 27579 1608 27611
rect 1648 27579 1680 27611
rect 1720 27579 1752 27611
rect 1792 27579 1824 27611
rect 1864 27579 1896 27611
rect 1936 27579 1968 27611
rect 2008 27579 2040 27611
rect 2080 27579 2112 27611
rect 2152 27579 2184 27611
rect 2224 27579 2256 27611
rect 2296 27579 2328 27611
rect 2368 27579 2400 27611
rect 2440 27579 2472 27611
rect 2512 27579 2544 27611
rect 2584 27579 2616 27611
rect 2656 27579 2688 27611
rect 2728 27579 2760 27611
rect 2800 27579 2832 27611
rect 2872 27579 2904 27611
rect 2944 27579 2976 27611
rect 3016 27579 3048 27611
rect 3088 27579 3120 27611
rect 3160 27579 3192 27611
rect 3232 27579 3264 27611
rect 3304 27579 3336 27611
rect 3376 27579 3408 27611
rect 3448 27579 3480 27611
rect 3520 27579 3552 27611
rect 3592 27579 3624 27611
rect 3664 27579 3696 27611
rect 3736 27579 3768 27611
rect 3808 27579 3840 27611
rect 3880 27579 3912 27611
rect 3952 27579 3984 27611
rect 4024 27579 4056 27611
rect 4096 27579 4128 27611
rect 4168 27579 4200 27611
rect 4240 27579 4272 27611
rect 4312 27579 4344 27611
rect 4384 27579 4416 27611
rect 4456 27579 4488 27611
rect 4528 27579 4560 27611
rect 4600 27579 4632 27611
rect 4672 27579 4704 27611
rect 4744 27579 4776 27611
rect 4816 27579 4848 27611
rect 4888 27579 4920 27611
rect 4960 27579 4992 27611
rect 5032 27579 5064 27611
rect 5104 27579 5136 27611
rect 5176 27579 5208 27611
rect 5248 27579 5280 27611
rect 5320 27579 5352 27611
rect 5392 27579 5424 27611
rect 5464 27579 5496 27611
rect 5536 27579 5568 27611
rect 5608 27579 5640 27611
rect 5680 27579 5712 27611
rect 5752 27579 5784 27611
rect 5824 27579 5856 27611
rect 5896 27579 5928 27611
rect 5968 27579 6000 27611
rect 6040 27579 6072 27611
rect 6112 27579 6144 27611
rect 6184 27579 6216 27611
rect 6256 27579 6288 27611
rect 6328 27579 6360 27611
rect 6400 27579 6432 27611
rect 6472 27579 6504 27611
rect 6544 27579 6576 27611
rect 6616 27579 6648 27611
rect 6688 27579 6720 27611
rect 6760 27579 6792 27611
rect 6832 27579 6864 27611
rect 6904 27579 6936 27611
rect 6976 27579 7008 27611
rect 7048 27579 7080 27611
rect 7120 27579 7152 27611
rect 7192 27579 7224 27611
rect 7264 27579 7296 27611
rect 7336 27579 7368 27611
rect 7408 27579 7440 27611
rect 7480 27579 7512 27611
rect 7552 27579 7584 27611
rect 7624 27579 7656 27611
rect 7696 27579 7728 27611
rect 7768 27579 7800 27611
rect 7840 27579 7872 27611
rect 7912 27579 7944 27611
rect 7984 27579 8016 27611
rect 8056 27579 8088 27611
rect 8128 27579 8160 27611
rect 8200 27579 8232 27611
rect 8272 27579 8304 27611
rect 8344 27579 8376 27611
rect 8416 27579 8448 27611
rect 8488 27579 8520 27611
rect 8560 27579 8592 27611
rect 8632 27579 8664 27611
rect 8704 27579 8736 27611
rect 8776 27579 8808 27611
rect 8848 27579 8880 27611
rect 8920 27579 8952 27611
rect 8992 27579 9024 27611
rect 9064 27579 9096 27611
rect 9136 27579 9168 27611
rect 9208 27579 9240 27611
rect 9280 27579 9312 27611
rect 9352 27579 9384 27611
rect 9424 27579 9456 27611
rect 9496 27579 9528 27611
rect 9568 27579 9600 27611
rect 9640 27579 9672 27611
rect 9712 27579 9744 27611
rect 9784 27579 9816 27611
rect 9856 27579 9888 27611
rect 9928 27579 9960 27611
rect 10000 27579 10032 27611
rect 10072 27579 10104 27611
rect 10144 27579 10176 27611
rect 10216 27579 10248 27611
rect 10288 27579 10320 27611
rect 10360 27579 10392 27611
rect 10432 27579 10464 27611
rect 10504 27579 10536 27611
rect 10576 27579 10608 27611
rect 10648 27579 10680 27611
rect 10720 27579 10752 27611
rect 10792 27579 10824 27611
rect 10864 27579 10896 27611
rect 10936 27579 10968 27611
rect 11008 27579 11040 27611
rect 11080 27579 11112 27611
rect 11152 27579 11184 27611
rect 11224 27579 11256 27611
rect 11296 27579 11328 27611
rect 11368 27579 11400 27611
rect 11440 27579 11472 27611
rect 11512 27579 11544 27611
rect 11584 27579 11616 27611
rect 11656 27579 11688 27611
rect 11728 27579 11760 27611
rect 11800 27579 11832 27611
rect 11872 27579 11904 27611
rect 11944 27579 11976 27611
rect 12016 27579 12048 27611
rect 12088 27579 12120 27611
rect 12160 27579 12192 27611
rect 12232 27579 12264 27611
rect 12304 27579 12336 27611
rect 12376 27579 12408 27611
rect 12448 27579 12480 27611
rect 12520 27579 12552 27611
rect 12592 27579 12624 27611
rect 12664 27579 12696 27611
rect 12736 27579 12768 27611
rect 12808 27579 12840 27611
rect 12880 27579 12912 27611
rect 12952 27579 12984 27611
rect 13024 27579 13056 27611
rect 13096 27579 13128 27611
rect 13168 27579 13200 27611
rect 13240 27579 13272 27611
rect 13312 27579 13344 27611
rect 13384 27579 13416 27611
rect 13456 27579 13488 27611
rect 13528 27579 13560 27611
rect 13600 27579 13632 27611
rect 13672 27579 13704 27611
rect 13744 27579 13776 27611
rect 13816 27579 13848 27611
rect 13888 27579 13920 27611
rect 13960 27579 13992 27611
rect 14032 27579 14064 27611
rect 14104 27579 14136 27611
rect 14176 27579 14208 27611
rect 14248 27579 14280 27611
rect 14320 27579 14352 27611
rect 14392 27579 14424 27611
rect 14464 27579 14496 27611
rect 14536 27579 14568 27611
rect 14608 27579 14640 27611
rect 14680 27579 14712 27611
rect 14752 27579 14784 27611
rect 14824 27579 14856 27611
rect 14896 27579 14928 27611
rect 14968 27579 15000 27611
rect 15040 27579 15072 27611
rect 15112 27579 15144 27611
rect 15184 27579 15216 27611
rect 15256 27579 15288 27611
rect 15328 27579 15360 27611
rect 15400 27579 15432 27611
rect 15472 27579 15504 27611
rect 15544 27579 15576 27611
rect 15616 27579 15648 27611
rect 15688 27579 15720 27611
rect 15760 27579 15792 27611
rect 15832 27579 15864 27611
rect 15904 27579 15936 27611
rect 64 27507 96 27539
rect 136 27507 168 27539
rect 208 27507 240 27539
rect 280 27507 312 27539
rect 352 27507 384 27539
rect 424 27507 456 27539
rect 496 27507 528 27539
rect 568 27507 600 27539
rect 640 27507 672 27539
rect 712 27507 744 27539
rect 784 27507 816 27539
rect 856 27507 888 27539
rect 928 27507 960 27539
rect 1000 27507 1032 27539
rect 1072 27507 1104 27539
rect 1144 27507 1176 27539
rect 1216 27507 1248 27539
rect 1288 27507 1320 27539
rect 1360 27507 1392 27539
rect 1432 27507 1464 27539
rect 1504 27507 1536 27539
rect 1576 27507 1608 27539
rect 1648 27507 1680 27539
rect 1720 27507 1752 27539
rect 1792 27507 1824 27539
rect 1864 27507 1896 27539
rect 1936 27507 1968 27539
rect 2008 27507 2040 27539
rect 2080 27507 2112 27539
rect 2152 27507 2184 27539
rect 2224 27507 2256 27539
rect 2296 27507 2328 27539
rect 2368 27507 2400 27539
rect 2440 27507 2472 27539
rect 2512 27507 2544 27539
rect 2584 27507 2616 27539
rect 2656 27507 2688 27539
rect 2728 27507 2760 27539
rect 2800 27507 2832 27539
rect 2872 27507 2904 27539
rect 2944 27507 2976 27539
rect 3016 27507 3048 27539
rect 3088 27507 3120 27539
rect 3160 27507 3192 27539
rect 3232 27507 3264 27539
rect 3304 27507 3336 27539
rect 3376 27507 3408 27539
rect 3448 27507 3480 27539
rect 3520 27507 3552 27539
rect 3592 27507 3624 27539
rect 3664 27507 3696 27539
rect 3736 27507 3768 27539
rect 3808 27507 3840 27539
rect 3880 27507 3912 27539
rect 3952 27507 3984 27539
rect 4024 27507 4056 27539
rect 4096 27507 4128 27539
rect 4168 27507 4200 27539
rect 4240 27507 4272 27539
rect 4312 27507 4344 27539
rect 4384 27507 4416 27539
rect 4456 27507 4488 27539
rect 4528 27507 4560 27539
rect 4600 27507 4632 27539
rect 4672 27507 4704 27539
rect 4744 27507 4776 27539
rect 4816 27507 4848 27539
rect 4888 27507 4920 27539
rect 4960 27507 4992 27539
rect 5032 27507 5064 27539
rect 5104 27507 5136 27539
rect 5176 27507 5208 27539
rect 5248 27507 5280 27539
rect 5320 27507 5352 27539
rect 5392 27507 5424 27539
rect 5464 27507 5496 27539
rect 5536 27507 5568 27539
rect 5608 27507 5640 27539
rect 5680 27507 5712 27539
rect 5752 27507 5784 27539
rect 5824 27507 5856 27539
rect 5896 27507 5928 27539
rect 5968 27507 6000 27539
rect 6040 27507 6072 27539
rect 6112 27507 6144 27539
rect 6184 27507 6216 27539
rect 6256 27507 6288 27539
rect 6328 27507 6360 27539
rect 6400 27507 6432 27539
rect 6472 27507 6504 27539
rect 6544 27507 6576 27539
rect 6616 27507 6648 27539
rect 6688 27507 6720 27539
rect 6760 27507 6792 27539
rect 6832 27507 6864 27539
rect 6904 27507 6936 27539
rect 6976 27507 7008 27539
rect 7048 27507 7080 27539
rect 7120 27507 7152 27539
rect 7192 27507 7224 27539
rect 7264 27507 7296 27539
rect 7336 27507 7368 27539
rect 7408 27507 7440 27539
rect 7480 27507 7512 27539
rect 7552 27507 7584 27539
rect 7624 27507 7656 27539
rect 7696 27507 7728 27539
rect 7768 27507 7800 27539
rect 7840 27507 7872 27539
rect 7912 27507 7944 27539
rect 7984 27507 8016 27539
rect 8056 27507 8088 27539
rect 8128 27507 8160 27539
rect 8200 27507 8232 27539
rect 8272 27507 8304 27539
rect 8344 27507 8376 27539
rect 8416 27507 8448 27539
rect 8488 27507 8520 27539
rect 8560 27507 8592 27539
rect 8632 27507 8664 27539
rect 8704 27507 8736 27539
rect 8776 27507 8808 27539
rect 8848 27507 8880 27539
rect 8920 27507 8952 27539
rect 8992 27507 9024 27539
rect 9064 27507 9096 27539
rect 9136 27507 9168 27539
rect 9208 27507 9240 27539
rect 9280 27507 9312 27539
rect 9352 27507 9384 27539
rect 9424 27507 9456 27539
rect 9496 27507 9528 27539
rect 9568 27507 9600 27539
rect 9640 27507 9672 27539
rect 9712 27507 9744 27539
rect 9784 27507 9816 27539
rect 9856 27507 9888 27539
rect 9928 27507 9960 27539
rect 10000 27507 10032 27539
rect 10072 27507 10104 27539
rect 10144 27507 10176 27539
rect 10216 27507 10248 27539
rect 10288 27507 10320 27539
rect 10360 27507 10392 27539
rect 10432 27507 10464 27539
rect 10504 27507 10536 27539
rect 10576 27507 10608 27539
rect 10648 27507 10680 27539
rect 10720 27507 10752 27539
rect 10792 27507 10824 27539
rect 10864 27507 10896 27539
rect 10936 27507 10968 27539
rect 11008 27507 11040 27539
rect 11080 27507 11112 27539
rect 11152 27507 11184 27539
rect 11224 27507 11256 27539
rect 11296 27507 11328 27539
rect 11368 27507 11400 27539
rect 11440 27507 11472 27539
rect 11512 27507 11544 27539
rect 11584 27507 11616 27539
rect 11656 27507 11688 27539
rect 11728 27507 11760 27539
rect 11800 27507 11832 27539
rect 11872 27507 11904 27539
rect 11944 27507 11976 27539
rect 12016 27507 12048 27539
rect 12088 27507 12120 27539
rect 12160 27507 12192 27539
rect 12232 27507 12264 27539
rect 12304 27507 12336 27539
rect 12376 27507 12408 27539
rect 12448 27507 12480 27539
rect 12520 27507 12552 27539
rect 12592 27507 12624 27539
rect 12664 27507 12696 27539
rect 12736 27507 12768 27539
rect 12808 27507 12840 27539
rect 12880 27507 12912 27539
rect 12952 27507 12984 27539
rect 13024 27507 13056 27539
rect 13096 27507 13128 27539
rect 13168 27507 13200 27539
rect 13240 27507 13272 27539
rect 13312 27507 13344 27539
rect 13384 27507 13416 27539
rect 13456 27507 13488 27539
rect 13528 27507 13560 27539
rect 13600 27507 13632 27539
rect 13672 27507 13704 27539
rect 13744 27507 13776 27539
rect 13816 27507 13848 27539
rect 13888 27507 13920 27539
rect 13960 27507 13992 27539
rect 14032 27507 14064 27539
rect 14104 27507 14136 27539
rect 14176 27507 14208 27539
rect 14248 27507 14280 27539
rect 14320 27507 14352 27539
rect 14392 27507 14424 27539
rect 14464 27507 14496 27539
rect 14536 27507 14568 27539
rect 14608 27507 14640 27539
rect 14680 27507 14712 27539
rect 14752 27507 14784 27539
rect 14824 27507 14856 27539
rect 14896 27507 14928 27539
rect 14968 27507 15000 27539
rect 15040 27507 15072 27539
rect 15112 27507 15144 27539
rect 15184 27507 15216 27539
rect 15256 27507 15288 27539
rect 15328 27507 15360 27539
rect 15400 27507 15432 27539
rect 15472 27507 15504 27539
rect 15544 27507 15576 27539
rect 15616 27507 15648 27539
rect 15688 27507 15720 27539
rect 15760 27507 15792 27539
rect 15832 27507 15864 27539
rect 15904 27507 15936 27539
rect 64 27435 96 27467
rect 136 27435 168 27467
rect 208 27435 240 27467
rect 280 27435 312 27467
rect 352 27435 384 27467
rect 424 27435 456 27467
rect 496 27435 528 27467
rect 568 27435 600 27467
rect 640 27435 672 27467
rect 712 27435 744 27467
rect 784 27435 816 27467
rect 856 27435 888 27467
rect 928 27435 960 27467
rect 1000 27435 1032 27467
rect 1072 27435 1104 27467
rect 1144 27435 1176 27467
rect 1216 27435 1248 27467
rect 1288 27435 1320 27467
rect 1360 27435 1392 27467
rect 1432 27435 1464 27467
rect 1504 27435 1536 27467
rect 1576 27435 1608 27467
rect 1648 27435 1680 27467
rect 1720 27435 1752 27467
rect 1792 27435 1824 27467
rect 1864 27435 1896 27467
rect 1936 27435 1968 27467
rect 2008 27435 2040 27467
rect 2080 27435 2112 27467
rect 2152 27435 2184 27467
rect 2224 27435 2256 27467
rect 2296 27435 2328 27467
rect 2368 27435 2400 27467
rect 2440 27435 2472 27467
rect 2512 27435 2544 27467
rect 2584 27435 2616 27467
rect 2656 27435 2688 27467
rect 2728 27435 2760 27467
rect 2800 27435 2832 27467
rect 2872 27435 2904 27467
rect 2944 27435 2976 27467
rect 3016 27435 3048 27467
rect 3088 27435 3120 27467
rect 3160 27435 3192 27467
rect 3232 27435 3264 27467
rect 3304 27435 3336 27467
rect 3376 27435 3408 27467
rect 3448 27435 3480 27467
rect 3520 27435 3552 27467
rect 3592 27435 3624 27467
rect 3664 27435 3696 27467
rect 3736 27435 3768 27467
rect 3808 27435 3840 27467
rect 3880 27435 3912 27467
rect 3952 27435 3984 27467
rect 4024 27435 4056 27467
rect 4096 27435 4128 27467
rect 4168 27435 4200 27467
rect 4240 27435 4272 27467
rect 4312 27435 4344 27467
rect 4384 27435 4416 27467
rect 4456 27435 4488 27467
rect 4528 27435 4560 27467
rect 4600 27435 4632 27467
rect 4672 27435 4704 27467
rect 4744 27435 4776 27467
rect 4816 27435 4848 27467
rect 4888 27435 4920 27467
rect 4960 27435 4992 27467
rect 5032 27435 5064 27467
rect 5104 27435 5136 27467
rect 5176 27435 5208 27467
rect 5248 27435 5280 27467
rect 5320 27435 5352 27467
rect 5392 27435 5424 27467
rect 5464 27435 5496 27467
rect 5536 27435 5568 27467
rect 5608 27435 5640 27467
rect 5680 27435 5712 27467
rect 5752 27435 5784 27467
rect 5824 27435 5856 27467
rect 5896 27435 5928 27467
rect 5968 27435 6000 27467
rect 6040 27435 6072 27467
rect 6112 27435 6144 27467
rect 6184 27435 6216 27467
rect 6256 27435 6288 27467
rect 6328 27435 6360 27467
rect 6400 27435 6432 27467
rect 6472 27435 6504 27467
rect 6544 27435 6576 27467
rect 6616 27435 6648 27467
rect 6688 27435 6720 27467
rect 6760 27435 6792 27467
rect 6832 27435 6864 27467
rect 6904 27435 6936 27467
rect 6976 27435 7008 27467
rect 7048 27435 7080 27467
rect 7120 27435 7152 27467
rect 7192 27435 7224 27467
rect 7264 27435 7296 27467
rect 7336 27435 7368 27467
rect 7408 27435 7440 27467
rect 7480 27435 7512 27467
rect 7552 27435 7584 27467
rect 7624 27435 7656 27467
rect 7696 27435 7728 27467
rect 7768 27435 7800 27467
rect 7840 27435 7872 27467
rect 7912 27435 7944 27467
rect 7984 27435 8016 27467
rect 8056 27435 8088 27467
rect 8128 27435 8160 27467
rect 8200 27435 8232 27467
rect 8272 27435 8304 27467
rect 8344 27435 8376 27467
rect 8416 27435 8448 27467
rect 8488 27435 8520 27467
rect 8560 27435 8592 27467
rect 8632 27435 8664 27467
rect 8704 27435 8736 27467
rect 8776 27435 8808 27467
rect 8848 27435 8880 27467
rect 8920 27435 8952 27467
rect 8992 27435 9024 27467
rect 9064 27435 9096 27467
rect 9136 27435 9168 27467
rect 9208 27435 9240 27467
rect 9280 27435 9312 27467
rect 9352 27435 9384 27467
rect 9424 27435 9456 27467
rect 9496 27435 9528 27467
rect 9568 27435 9600 27467
rect 9640 27435 9672 27467
rect 9712 27435 9744 27467
rect 9784 27435 9816 27467
rect 9856 27435 9888 27467
rect 9928 27435 9960 27467
rect 10000 27435 10032 27467
rect 10072 27435 10104 27467
rect 10144 27435 10176 27467
rect 10216 27435 10248 27467
rect 10288 27435 10320 27467
rect 10360 27435 10392 27467
rect 10432 27435 10464 27467
rect 10504 27435 10536 27467
rect 10576 27435 10608 27467
rect 10648 27435 10680 27467
rect 10720 27435 10752 27467
rect 10792 27435 10824 27467
rect 10864 27435 10896 27467
rect 10936 27435 10968 27467
rect 11008 27435 11040 27467
rect 11080 27435 11112 27467
rect 11152 27435 11184 27467
rect 11224 27435 11256 27467
rect 11296 27435 11328 27467
rect 11368 27435 11400 27467
rect 11440 27435 11472 27467
rect 11512 27435 11544 27467
rect 11584 27435 11616 27467
rect 11656 27435 11688 27467
rect 11728 27435 11760 27467
rect 11800 27435 11832 27467
rect 11872 27435 11904 27467
rect 11944 27435 11976 27467
rect 12016 27435 12048 27467
rect 12088 27435 12120 27467
rect 12160 27435 12192 27467
rect 12232 27435 12264 27467
rect 12304 27435 12336 27467
rect 12376 27435 12408 27467
rect 12448 27435 12480 27467
rect 12520 27435 12552 27467
rect 12592 27435 12624 27467
rect 12664 27435 12696 27467
rect 12736 27435 12768 27467
rect 12808 27435 12840 27467
rect 12880 27435 12912 27467
rect 12952 27435 12984 27467
rect 13024 27435 13056 27467
rect 13096 27435 13128 27467
rect 13168 27435 13200 27467
rect 13240 27435 13272 27467
rect 13312 27435 13344 27467
rect 13384 27435 13416 27467
rect 13456 27435 13488 27467
rect 13528 27435 13560 27467
rect 13600 27435 13632 27467
rect 13672 27435 13704 27467
rect 13744 27435 13776 27467
rect 13816 27435 13848 27467
rect 13888 27435 13920 27467
rect 13960 27435 13992 27467
rect 14032 27435 14064 27467
rect 14104 27435 14136 27467
rect 14176 27435 14208 27467
rect 14248 27435 14280 27467
rect 14320 27435 14352 27467
rect 14392 27435 14424 27467
rect 14464 27435 14496 27467
rect 14536 27435 14568 27467
rect 14608 27435 14640 27467
rect 14680 27435 14712 27467
rect 14752 27435 14784 27467
rect 14824 27435 14856 27467
rect 14896 27435 14928 27467
rect 14968 27435 15000 27467
rect 15040 27435 15072 27467
rect 15112 27435 15144 27467
rect 15184 27435 15216 27467
rect 15256 27435 15288 27467
rect 15328 27435 15360 27467
rect 15400 27435 15432 27467
rect 15472 27435 15504 27467
rect 15544 27435 15576 27467
rect 15616 27435 15648 27467
rect 15688 27435 15720 27467
rect 15760 27435 15792 27467
rect 15832 27435 15864 27467
rect 15904 27435 15936 27467
rect 64 27363 96 27395
rect 136 27363 168 27395
rect 208 27363 240 27395
rect 280 27363 312 27395
rect 352 27363 384 27395
rect 424 27363 456 27395
rect 496 27363 528 27395
rect 568 27363 600 27395
rect 640 27363 672 27395
rect 712 27363 744 27395
rect 784 27363 816 27395
rect 856 27363 888 27395
rect 928 27363 960 27395
rect 1000 27363 1032 27395
rect 1072 27363 1104 27395
rect 1144 27363 1176 27395
rect 1216 27363 1248 27395
rect 1288 27363 1320 27395
rect 1360 27363 1392 27395
rect 1432 27363 1464 27395
rect 1504 27363 1536 27395
rect 1576 27363 1608 27395
rect 1648 27363 1680 27395
rect 1720 27363 1752 27395
rect 1792 27363 1824 27395
rect 1864 27363 1896 27395
rect 1936 27363 1968 27395
rect 2008 27363 2040 27395
rect 2080 27363 2112 27395
rect 2152 27363 2184 27395
rect 2224 27363 2256 27395
rect 2296 27363 2328 27395
rect 2368 27363 2400 27395
rect 2440 27363 2472 27395
rect 2512 27363 2544 27395
rect 2584 27363 2616 27395
rect 2656 27363 2688 27395
rect 2728 27363 2760 27395
rect 2800 27363 2832 27395
rect 2872 27363 2904 27395
rect 2944 27363 2976 27395
rect 3016 27363 3048 27395
rect 3088 27363 3120 27395
rect 3160 27363 3192 27395
rect 3232 27363 3264 27395
rect 3304 27363 3336 27395
rect 3376 27363 3408 27395
rect 3448 27363 3480 27395
rect 3520 27363 3552 27395
rect 3592 27363 3624 27395
rect 3664 27363 3696 27395
rect 3736 27363 3768 27395
rect 3808 27363 3840 27395
rect 3880 27363 3912 27395
rect 3952 27363 3984 27395
rect 4024 27363 4056 27395
rect 4096 27363 4128 27395
rect 4168 27363 4200 27395
rect 4240 27363 4272 27395
rect 4312 27363 4344 27395
rect 4384 27363 4416 27395
rect 4456 27363 4488 27395
rect 4528 27363 4560 27395
rect 4600 27363 4632 27395
rect 4672 27363 4704 27395
rect 4744 27363 4776 27395
rect 4816 27363 4848 27395
rect 4888 27363 4920 27395
rect 4960 27363 4992 27395
rect 5032 27363 5064 27395
rect 5104 27363 5136 27395
rect 5176 27363 5208 27395
rect 5248 27363 5280 27395
rect 5320 27363 5352 27395
rect 5392 27363 5424 27395
rect 5464 27363 5496 27395
rect 5536 27363 5568 27395
rect 5608 27363 5640 27395
rect 5680 27363 5712 27395
rect 5752 27363 5784 27395
rect 5824 27363 5856 27395
rect 5896 27363 5928 27395
rect 5968 27363 6000 27395
rect 6040 27363 6072 27395
rect 6112 27363 6144 27395
rect 6184 27363 6216 27395
rect 6256 27363 6288 27395
rect 6328 27363 6360 27395
rect 6400 27363 6432 27395
rect 6472 27363 6504 27395
rect 6544 27363 6576 27395
rect 6616 27363 6648 27395
rect 6688 27363 6720 27395
rect 6760 27363 6792 27395
rect 6832 27363 6864 27395
rect 6904 27363 6936 27395
rect 6976 27363 7008 27395
rect 7048 27363 7080 27395
rect 7120 27363 7152 27395
rect 7192 27363 7224 27395
rect 7264 27363 7296 27395
rect 7336 27363 7368 27395
rect 7408 27363 7440 27395
rect 7480 27363 7512 27395
rect 7552 27363 7584 27395
rect 7624 27363 7656 27395
rect 7696 27363 7728 27395
rect 7768 27363 7800 27395
rect 7840 27363 7872 27395
rect 7912 27363 7944 27395
rect 7984 27363 8016 27395
rect 8056 27363 8088 27395
rect 8128 27363 8160 27395
rect 8200 27363 8232 27395
rect 8272 27363 8304 27395
rect 8344 27363 8376 27395
rect 8416 27363 8448 27395
rect 8488 27363 8520 27395
rect 8560 27363 8592 27395
rect 8632 27363 8664 27395
rect 8704 27363 8736 27395
rect 8776 27363 8808 27395
rect 8848 27363 8880 27395
rect 8920 27363 8952 27395
rect 8992 27363 9024 27395
rect 9064 27363 9096 27395
rect 9136 27363 9168 27395
rect 9208 27363 9240 27395
rect 9280 27363 9312 27395
rect 9352 27363 9384 27395
rect 9424 27363 9456 27395
rect 9496 27363 9528 27395
rect 9568 27363 9600 27395
rect 9640 27363 9672 27395
rect 9712 27363 9744 27395
rect 9784 27363 9816 27395
rect 9856 27363 9888 27395
rect 9928 27363 9960 27395
rect 10000 27363 10032 27395
rect 10072 27363 10104 27395
rect 10144 27363 10176 27395
rect 10216 27363 10248 27395
rect 10288 27363 10320 27395
rect 10360 27363 10392 27395
rect 10432 27363 10464 27395
rect 10504 27363 10536 27395
rect 10576 27363 10608 27395
rect 10648 27363 10680 27395
rect 10720 27363 10752 27395
rect 10792 27363 10824 27395
rect 10864 27363 10896 27395
rect 10936 27363 10968 27395
rect 11008 27363 11040 27395
rect 11080 27363 11112 27395
rect 11152 27363 11184 27395
rect 11224 27363 11256 27395
rect 11296 27363 11328 27395
rect 11368 27363 11400 27395
rect 11440 27363 11472 27395
rect 11512 27363 11544 27395
rect 11584 27363 11616 27395
rect 11656 27363 11688 27395
rect 11728 27363 11760 27395
rect 11800 27363 11832 27395
rect 11872 27363 11904 27395
rect 11944 27363 11976 27395
rect 12016 27363 12048 27395
rect 12088 27363 12120 27395
rect 12160 27363 12192 27395
rect 12232 27363 12264 27395
rect 12304 27363 12336 27395
rect 12376 27363 12408 27395
rect 12448 27363 12480 27395
rect 12520 27363 12552 27395
rect 12592 27363 12624 27395
rect 12664 27363 12696 27395
rect 12736 27363 12768 27395
rect 12808 27363 12840 27395
rect 12880 27363 12912 27395
rect 12952 27363 12984 27395
rect 13024 27363 13056 27395
rect 13096 27363 13128 27395
rect 13168 27363 13200 27395
rect 13240 27363 13272 27395
rect 13312 27363 13344 27395
rect 13384 27363 13416 27395
rect 13456 27363 13488 27395
rect 13528 27363 13560 27395
rect 13600 27363 13632 27395
rect 13672 27363 13704 27395
rect 13744 27363 13776 27395
rect 13816 27363 13848 27395
rect 13888 27363 13920 27395
rect 13960 27363 13992 27395
rect 14032 27363 14064 27395
rect 14104 27363 14136 27395
rect 14176 27363 14208 27395
rect 14248 27363 14280 27395
rect 14320 27363 14352 27395
rect 14392 27363 14424 27395
rect 14464 27363 14496 27395
rect 14536 27363 14568 27395
rect 14608 27363 14640 27395
rect 14680 27363 14712 27395
rect 14752 27363 14784 27395
rect 14824 27363 14856 27395
rect 14896 27363 14928 27395
rect 14968 27363 15000 27395
rect 15040 27363 15072 27395
rect 15112 27363 15144 27395
rect 15184 27363 15216 27395
rect 15256 27363 15288 27395
rect 15328 27363 15360 27395
rect 15400 27363 15432 27395
rect 15472 27363 15504 27395
rect 15544 27363 15576 27395
rect 15616 27363 15648 27395
rect 15688 27363 15720 27395
rect 15760 27363 15792 27395
rect 15832 27363 15864 27395
rect 15904 27363 15936 27395
rect 64 27291 96 27323
rect 136 27291 168 27323
rect 208 27291 240 27323
rect 280 27291 312 27323
rect 352 27291 384 27323
rect 424 27291 456 27323
rect 496 27291 528 27323
rect 568 27291 600 27323
rect 640 27291 672 27323
rect 712 27291 744 27323
rect 784 27291 816 27323
rect 856 27291 888 27323
rect 928 27291 960 27323
rect 1000 27291 1032 27323
rect 1072 27291 1104 27323
rect 1144 27291 1176 27323
rect 1216 27291 1248 27323
rect 1288 27291 1320 27323
rect 1360 27291 1392 27323
rect 1432 27291 1464 27323
rect 1504 27291 1536 27323
rect 1576 27291 1608 27323
rect 1648 27291 1680 27323
rect 1720 27291 1752 27323
rect 1792 27291 1824 27323
rect 1864 27291 1896 27323
rect 1936 27291 1968 27323
rect 2008 27291 2040 27323
rect 2080 27291 2112 27323
rect 2152 27291 2184 27323
rect 2224 27291 2256 27323
rect 2296 27291 2328 27323
rect 2368 27291 2400 27323
rect 2440 27291 2472 27323
rect 2512 27291 2544 27323
rect 2584 27291 2616 27323
rect 2656 27291 2688 27323
rect 2728 27291 2760 27323
rect 2800 27291 2832 27323
rect 2872 27291 2904 27323
rect 2944 27291 2976 27323
rect 3016 27291 3048 27323
rect 3088 27291 3120 27323
rect 3160 27291 3192 27323
rect 3232 27291 3264 27323
rect 3304 27291 3336 27323
rect 3376 27291 3408 27323
rect 3448 27291 3480 27323
rect 3520 27291 3552 27323
rect 3592 27291 3624 27323
rect 3664 27291 3696 27323
rect 3736 27291 3768 27323
rect 3808 27291 3840 27323
rect 3880 27291 3912 27323
rect 3952 27291 3984 27323
rect 4024 27291 4056 27323
rect 4096 27291 4128 27323
rect 4168 27291 4200 27323
rect 4240 27291 4272 27323
rect 4312 27291 4344 27323
rect 4384 27291 4416 27323
rect 4456 27291 4488 27323
rect 4528 27291 4560 27323
rect 4600 27291 4632 27323
rect 4672 27291 4704 27323
rect 4744 27291 4776 27323
rect 4816 27291 4848 27323
rect 4888 27291 4920 27323
rect 4960 27291 4992 27323
rect 5032 27291 5064 27323
rect 5104 27291 5136 27323
rect 5176 27291 5208 27323
rect 5248 27291 5280 27323
rect 5320 27291 5352 27323
rect 5392 27291 5424 27323
rect 5464 27291 5496 27323
rect 5536 27291 5568 27323
rect 5608 27291 5640 27323
rect 5680 27291 5712 27323
rect 5752 27291 5784 27323
rect 5824 27291 5856 27323
rect 5896 27291 5928 27323
rect 5968 27291 6000 27323
rect 6040 27291 6072 27323
rect 6112 27291 6144 27323
rect 6184 27291 6216 27323
rect 6256 27291 6288 27323
rect 6328 27291 6360 27323
rect 6400 27291 6432 27323
rect 6472 27291 6504 27323
rect 6544 27291 6576 27323
rect 6616 27291 6648 27323
rect 6688 27291 6720 27323
rect 6760 27291 6792 27323
rect 6832 27291 6864 27323
rect 6904 27291 6936 27323
rect 6976 27291 7008 27323
rect 7048 27291 7080 27323
rect 7120 27291 7152 27323
rect 7192 27291 7224 27323
rect 7264 27291 7296 27323
rect 7336 27291 7368 27323
rect 7408 27291 7440 27323
rect 7480 27291 7512 27323
rect 7552 27291 7584 27323
rect 7624 27291 7656 27323
rect 7696 27291 7728 27323
rect 7768 27291 7800 27323
rect 7840 27291 7872 27323
rect 7912 27291 7944 27323
rect 7984 27291 8016 27323
rect 8056 27291 8088 27323
rect 8128 27291 8160 27323
rect 8200 27291 8232 27323
rect 8272 27291 8304 27323
rect 8344 27291 8376 27323
rect 8416 27291 8448 27323
rect 8488 27291 8520 27323
rect 8560 27291 8592 27323
rect 8632 27291 8664 27323
rect 8704 27291 8736 27323
rect 8776 27291 8808 27323
rect 8848 27291 8880 27323
rect 8920 27291 8952 27323
rect 8992 27291 9024 27323
rect 9064 27291 9096 27323
rect 9136 27291 9168 27323
rect 9208 27291 9240 27323
rect 9280 27291 9312 27323
rect 9352 27291 9384 27323
rect 9424 27291 9456 27323
rect 9496 27291 9528 27323
rect 9568 27291 9600 27323
rect 9640 27291 9672 27323
rect 9712 27291 9744 27323
rect 9784 27291 9816 27323
rect 9856 27291 9888 27323
rect 9928 27291 9960 27323
rect 10000 27291 10032 27323
rect 10072 27291 10104 27323
rect 10144 27291 10176 27323
rect 10216 27291 10248 27323
rect 10288 27291 10320 27323
rect 10360 27291 10392 27323
rect 10432 27291 10464 27323
rect 10504 27291 10536 27323
rect 10576 27291 10608 27323
rect 10648 27291 10680 27323
rect 10720 27291 10752 27323
rect 10792 27291 10824 27323
rect 10864 27291 10896 27323
rect 10936 27291 10968 27323
rect 11008 27291 11040 27323
rect 11080 27291 11112 27323
rect 11152 27291 11184 27323
rect 11224 27291 11256 27323
rect 11296 27291 11328 27323
rect 11368 27291 11400 27323
rect 11440 27291 11472 27323
rect 11512 27291 11544 27323
rect 11584 27291 11616 27323
rect 11656 27291 11688 27323
rect 11728 27291 11760 27323
rect 11800 27291 11832 27323
rect 11872 27291 11904 27323
rect 11944 27291 11976 27323
rect 12016 27291 12048 27323
rect 12088 27291 12120 27323
rect 12160 27291 12192 27323
rect 12232 27291 12264 27323
rect 12304 27291 12336 27323
rect 12376 27291 12408 27323
rect 12448 27291 12480 27323
rect 12520 27291 12552 27323
rect 12592 27291 12624 27323
rect 12664 27291 12696 27323
rect 12736 27291 12768 27323
rect 12808 27291 12840 27323
rect 12880 27291 12912 27323
rect 12952 27291 12984 27323
rect 13024 27291 13056 27323
rect 13096 27291 13128 27323
rect 13168 27291 13200 27323
rect 13240 27291 13272 27323
rect 13312 27291 13344 27323
rect 13384 27291 13416 27323
rect 13456 27291 13488 27323
rect 13528 27291 13560 27323
rect 13600 27291 13632 27323
rect 13672 27291 13704 27323
rect 13744 27291 13776 27323
rect 13816 27291 13848 27323
rect 13888 27291 13920 27323
rect 13960 27291 13992 27323
rect 14032 27291 14064 27323
rect 14104 27291 14136 27323
rect 14176 27291 14208 27323
rect 14248 27291 14280 27323
rect 14320 27291 14352 27323
rect 14392 27291 14424 27323
rect 14464 27291 14496 27323
rect 14536 27291 14568 27323
rect 14608 27291 14640 27323
rect 14680 27291 14712 27323
rect 14752 27291 14784 27323
rect 14824 27291 14856 27323
rect 14896 27291 14928 27323
rect 14968 27291 15000 27323
rect 15040 27291 15072 27323
rect 15112 27291 15144 27323
rect 15184 27291 15216 27323
rect 15256 27291 15288 27323
rect 15328 27291 15360 27323
rect 15400 27291 15432 27323
rect 15472 27291 15504 27323
rect 15544 27291 15576 27323
rect 15616 27291 15648 27323
rect 15688 27291 15720 27323
rect 15760 27291 15792 27323
rect 15832 27291 15864 27323
rect 15904 27291 15936 27323
rect 64 27219 96 27251
rect 136 27219 168 27251
rect 208 27219 240 27251
rect 280 27219 312 27251
rect 352 27219 384 27251
rect 424 27219 456 27251
rect 496 27219 528 27251
rect 568 27219 600 27251
rect 640 27219 672 27251
rect 712 27219 744 27251
rect 784 27219 816 27251
rect 856 27219 888 27251
rect 928 27219 960 27251
rect 1000 27219 1032 27251
rect 1072 27219 1104 27251
rect 1144 27219 1176 27251
rect 1216 27219 1248 27251
rect 1288 27219 1320 27251
rect 1360 27219 1392 27251
rect 1432 27219 1464 27251
rect 1504 27219 1536 27251
rect 1576 27219 1608 27251
rect 1648 27219 1680 27251
rect 1720 27219 1752 27251
rect 1792 27219 1824 27251
rect 1864 27219 1896 27251
rect 1936 27219 1968 27251
rect 2008 27219 2040 27251
rect 2080 27219 2112 27251
rect 2152 27219 2184 27251
rect 2224 27219 2256 27251
rect 2296 27219 2328 27251
rect 2368 27219 2400 27251
rect 2440 27219 2472 27251
rect 2512 27219 2544 27251
rect 2584 27219 2616 27251
rect 2656 27219 2688 27251
rect 2728 27219 2760 27251
rect 2800 27219 2832 27251
rect 2872 27219 2904 27251
rect 2944 27219 2976 27251
rect 3016 27219 3048 27251
rect 3088 27219 3120 27251
rect 3160 27219 3192 27251
rect 3232 27219 3264 27251
rect 3304 27219 3336 27251
rect 3376 27219 3408 27251
rect 3448 27219 3480 27251
rect 3520 27219 3552 27251
rect 3592 27219 3624 27251
rect 3664 27219 3696 27251
rect 3736 27219 3768 27251
rect 3808 27219 3840 27251
rect 3880 27219 3912 27251
rect 3952 27219 3984 27251
rect 4024 27219 4056 27251
rect 4096 27219 4128 27251
rect 4168 27219 4200 27251
rect 4240 27219 4272 27251
rect 4312 27219 4344 27251
rect 4384 27219 4416 27251
rect 4456 27219 4488 27251
rect 4528 27219 4560 27251
rect 4600 27219 4632 27251
rect 4672 27219 4704 27251
rect 4744 27219 4776 27251
rect 4816 27219 4848 27251
rect 4888 27219 4920 27251
rect 4960 27219 4992 27251
rect 5032 27219 5064 27251
rect 5104 27219 5136 27251
rect 5176 27219 5208 27251
rect 5248 27219 5280 27251
rect 5320 27219 5352 27251
rect 5392 27219 5424 27251
rect 5464 27219 5496 27251
rect 5536 27219 5568 27251
rect 5608 27219 5640 27251
rect 5680 27219 5712 27251
rect 5752 27219 5784 27251
rect 5824 27219 5856 27251
rect 5896 27219 5928 27251
rect 5968 27219 6000 27251
rect 6040 27219 6072 27251
rect 6112 27219 6144 27251
rect 6184 27219 6216 27251
rect 6256 27219 6288 27251
rect 6328 27219 6360 27251
rect 6400 27219 6432 27251
rect 6472 27219 6504 27251
rect 6544 27219 6576 27251
rect 6616 27219 6648 27251
rect 6688 27219 6720 27251
rect 6760 27219 6792 27251
rect 6832 27219 6864 27251
rect 6904 27219 6936 27251
rect 6976 27219 7008 27251
rect 7048 27219 7080 27251
rect 7120 27219 7152 27251
rect 7192 27219 7224 27251
rect 7264 27219 7296 27251
rect 7336 27219 7368 27251
rect 7408 27219 7440 27251
rect 7480 27219 7512 27251
rect 7552 27219 7584 27251
rect 7624 27219 7656 27251
rect 7696 27219 7728 27251
rect 7768 27219 7800 27251
rect 7840 27219 7872 27251
rect 7912 27219 7944 27251
rect 7984 27219 8016 27251
rect 8056 27219 8088 27251
rect 8128 27219 8160 27251
rect 8200 27219 8232 27251
rect 8272 27219 8304 27251
rect 8344 27219 8376 27251
rect 8416 27219 8448 27251
rect 8488 27219 8520 27251
rect 8560 27219 8592 27251
rect 8632 27219 8664 27251
rect 8704 27219 8736 27251
rect 8776 27219 8808 27251
rect 8848 27219 8880 27251
rect 8920 27219 8952 27251
rect 8992 27219 9024 27251
rect 9064 27219 9096 27251
rect 9136 27219 9168 27251
rect 9208 27219 9240 27251
rect 9280 27219 9312 27251
rect 9352 27219 9384 27251
rect 9424 27219 9456 27251
rect 9496 27219 9528 27251
rect 9568 27219 9600 27251
rect 9640 27219 9672 27251
rect 9712 27219 9744 27251
rect 9784 27219 9816 27251
rect 9856 27219 9888 27251
rect 9928 27219 9960 27251
rect 10000 27219 10032 27251
rect 10072 27219 10104 27251
rect 10144 27219 10176 27251
rect 10216 27219 10248 27251
rect 10288 27219 10320 27251
rect 10360 27219 10392 27251
rect 10432 27219 10464 27251
rect 10504 27219 10536 27251
rect 10576 27219 10608 27251
rect 10648 27219 10680 27251
rect 10720 27219 10752 27251
rect 10792 27219 10824 27251
rect 10864 27219 10896 27251
rect 10936 27219 10968 27251
rect 11008 27219 11040 27251
rect 11080 27219 11112 27251
rect 11152 27219 11184 27251
rect 11224 27219 11256 27251
rect 11296 27219 11328 27251
rect 11368 27219 11400 27251
rect 11440 27219 11472 27251
rect 11512 27219 11544 27251
rect 11584 27219 11616 27251
rect 11656 27219 11688 27251
rect 11728 27219 11760 27251
rect 11800 27219 11832 27251
rect 11872 27219 11904 27251
rect 11944 27219 11976 27251
rect 12016 27219 12048 27251
rect 12088 27219 12120 27251
rect 12160 27219 12192 27251
rect 12232 27219 12264 27251
rect 12304 27219 12336 27251
rect 12376 27219 12408 27251
rect 12448 27219 12480 27251
rect 12520 27219 12552 27251
rect 12592 27219 12624 27251
rect 12664 27219 12696 27251
rect 12736 27219 12768 27251
rect 12808 27219 12840 27251
rect 12880 27219 12912 27251
rect 12952 27219 12984 27251
rect 13024 27219 13056 27251
rect 13096 27219 13128 27251
rect 13168 27219 13200 27251
rect 13240 27219 13272 27251
rect 13312 27219 13344 27251
rect 13384 27219 13416 27251
rect 13456 27219 13488 27251
rect 13528 27219 13560 27251
rect 13600 27219 13632 27251
rect 13672 27219 13704 27251
rect 13744 27219 13776 27251
rect 13816 27219 13848 27251
rect 13888 27219 13920 27251
rect 13960 27219 13992 27251
rect 14032 27219 14064 27251
rect 14104 27219 14136 27251
rect 14176 27219 14208 27251
rect 14248 27219 14280 27251
rect 14320 27219 14352 27251
rect 14392 27219 14424 27251
rect 14464 27219 14496 27251
rect 14536 27219 14568 27251
rect 14608 27219 14640 27251
rect 14680 27219 14712 27251
rect 14752 27219 14784 27251
rect 14824 27219 14856 27251
rect 14896 27219 14928 27251
rect 14968 27219 15000 27251
rect 15040 27219 15072 27251
rect 15112 27219 15144 27251
rect 15184 27219 15216 27251
rect 15256 27219 15288 27251
rect 15328 27219 15360 27251
rect 15400 27219 15432 27251
rect 15472 27219 15504 27251
rect 15544 27219 15576 27251
rect 15616 27219 15648 27251
rect 15688 27219 15720 27251
rect 15760 27219 15792 27251
rect 15832 27219 15864 27251
rect 15904 27219 15936 27251
rect 64 27147 96 27179
rect 136 27147 168 27179
rect 208 27147 240 27179
rect 280 27147 312 27179
rect 352 27147 384 27179
rect 424 27147 456 27179
rect 496 27147 528 27179
rect 568 27147 600 27179
rect 640 27147 672 27179
rect 712 27147 744 27179
rect 784 27147 816 27179
rect 856 27147 888 27179
rect 928 27147 960 27179
rect 1000 27147 1032 27179
rect 1072 27147 1104 27179
rect 1144 27147 1176 27179
rect 1216 27147 1248 27179
rect 1288 27147 1320 27179
rect 1360 27147 1392 27179
rect 1432 27147 1464 27179
rect 1504 27147 1536 27179
rect 1576 27147 1608 27179
rect 1648 27147 1680 27179
rect 1720 27147 1752 27179
rect 1792 27147 1824 27179
rect 1864 27147 1896 27179
rect 1936 27147 1968 27179
rect 2008 27147 2040 27179
rect 2080 27147 2112 27179
rect 2152 27147 2184 27179
rect 2224 27147 2256 27179
rect 2296 27147 2328 27179
rect 2368 27147 2400 27179
rect 2440 27147 2472 27179
rect 2512 27147 2544 27179
rect 2584 27147 2616 27179
rect 2656 27147 2688 27179
rect 2728 27147 2760 27179
rect 2800 27147 2832 27179
rect 2872 27147 2904 27179
rect 2944 27147 2976 27179
rect 3016 27147 3048 27179
rect 3088 27147 3120 27179
rect 3160 27147 3192 27179
rect 3232 27147 3264 27179
rect 3304 27147 3336 27179
rect 3376 27147 3408 27179
rect 3448 27147 3480 27179
rect 3520 27147 3552 27179
rect 3592 27147 3624 27179
rect 3664 27147 3696 27179
rect 3736 27147 3768 27179
rect 3808 27147 3840 27179
rect 3880 27147 3912 27179
rect 3952 27147 3984 27179
rect 4024 27147 4056 27179
rect 4096 27147 4128 27179
rect 4168 27147 4200 27179
rect 4240 27147 4272 27179
rect 4312 27147 4344 27179
rect 4384 27147 4416 27179
rect 4456 27147 4488 27179
rect 4528 27147 4560 27179
rect 4600 27147 4632 27179
rect 4672 27147 4704 27179
rect 4744 27147 4776 27179
rect 4816 27147 4848 27179
rect 4888 27147 4920 27179
rect 4960 27147 4992 27179
rect 5032 27147 5064 27179
rect 5104 27147 5136 27179
rect 5176 27147 5208 27179
rect 5248 27147 5280 27179
rect 5320 27147 5352 27179
rect 5392 27147 5424 27179
rect 5464 27147 5496 27179
rect 5536 27147 5568 27179
rect 5608 27147 5640 27179
rect 5680 27147 5712 27179
rect 5752 27147 5784 27179
rect 5824 27147 5856 27179
rect 5896 27147 5928 27179
rect 5968 27147 6000 27179
rect 6040 27147 6072 27179
rect 6112 27147 6144 27179
rect 6184 27147 6216 27179
rect 6256 27147 6288 27179
rect 6328 27147 6360 27179
rect 6400 27147 6432 27179
rect 6472 27147 6504 27179
rect 6544 27147 6576 27179
rect 6616 27147 6648 27179
rect 6688 27147 6720 27179
rect 6760 27147 6792 27179
rect 6832 27147 6864 27179
rect 6904 27147 6936 27179
rect 6976 27147 7008 27179
rect 7048 27147 7080 27179
rect 7120 27147 7152 27179
rect 7192 27147 7224 27179
rect 7264 27147 7296 27179
rect 7336 27147 7368 27179
rect 7408 27147 7440 27179
rect 7480 27147 7512 27179
rect 7552 27147 7584 27179
rect 7624 27147 7656 27179
rect 7696 27147 7728 27179
rect 7768 27147 7800 27179
rect 7840 27147 7872 27179
rect 7912 27147 7944 27179
rect 7984 27147 8016 27179
rect 8056 27147 8088 27179
rect 8128 27147 8160 27179
rect 8200 27147 8232 27179
rect 8272 27147 8304 27179
rect 8344 27147 8376 27179
rect 8416 27147 8448 27179
rect 8488 27147 8520 27179
rect 8560 27147 8592 27179
rect 8632 27147 8664 27179
rect 8704 27147 8736 27179
rect 8776 27147 8808 27179
rect 8848 27147 8880 27179
rect 8920 27147 8952 27179
rect 8992 27147 9024 27179
rect 9064 27147 9096 27179
rect 9136 27147 9168 27179
rect 9208 27147 9240 27179
rect 9280 27147 9312 27179
rect 9352 27147 9384 27179
rect 9424 27147 9456 27179
rect 9496 27147 9528 27179
rect 9568 27147 9600 27179
rect 9640 27147 9672 27179
rect 9712 27147 9744 27179
rect 9784 27147 9816 27179
rect 9856 27147 9888 27179
rect 9928 27147 9960 27179
rect 10000 27147 10032 27179
rect 10072 27147 10104 27179
rect 10144 27147 10176 27179
rect 10216 27147 10248 27179
rect 10288 27147 10320 27179
rect 10360 27147 10392 27179
rect 10432 27147 10464 27179
rect 10504 27147 10536 27179
rect 10576 27147 10608 27179
rect 10648 27147 10680 27179
rect 10720 27147 10752 27179
rect 10792 27147 10824 27179
rect 10864 27147 10896 27179
rect 10936 27147 10968 27179
rect 11008 27147 11040 27179
rect 11080 27147 11112 27179
rect 11152 27147 11184 27179
rect 11224 27147 11256 27179
rect 11296 27147 11328 27179
rect 11368 27147 11400 27179
rect 11440 27147 11472 27179
rect 11512 27147 11544 27179
rect 11584 27147 11616 27179
rect 11656 27147 11688 27179
rect 11728 27147 11760 27179
rect 11800 27147 11832 27179
rect 11872 27147 11904 27179
rect 11944 27147 11976 27179
rect 12016 27147 12048 27179
rect 12088 27147 12120 27179
rect 12160 27147 12192 27179
rect 12232 27147 12264 27179
rect 12304 27147 12336 27179
rect 12376 27147 12408 27179
rect 12448 27147 12480 27179
rect 12520 27147 12552 27179
rect 12592 27147 12624 27179
rect 12664 27147 12696 27179
rect 12736 27147 12768 27179
rect 12808 27147 12840 27179
rect 12880 27147 12912 27179
rect 12952 27147 12984 27179
rect 13024 27147 13056 27179
rect 13096 27147 13128 27179
rect 13168 27147 13200 27179
rect 13240 27147 13272 27179
rect 13312 27147 13344 27179
rect 13384 27147 13416 27179
rect 13456 27147 13488 27179
rect 13528 27147 13560 27179
rect 13600 27147 13632 27179
rect 13672 27147 13704 27179
rect 13744 27147 13776 27179
rect 13816 27147 13848 27179
rect 13888 27147 13920 27179
rect 13960 27147 13992 27179
rect 14032 27147 14064 27179
rect 14104 27147 14136 27179
rect 14176 27147 14208 27179
rect 14248 27147 14280 27179
rect 14320 27147 14352 27179
rect 14392 27147 14424 27179
rect 14464 27147 14496 27179
rect 14536 27147 14568 27179
rect 14608 27147 14640 27179
rect 14680 27147 14712 27179
rect 14752 27147 14784 27179
rect 14824 27147 14856 27179
rect 14896 27147 14928 27179
rect 14968 27147 15000 27179
rect 15040 27147 15072 27179
rect 15112 27147 15144 27179
rect 15184 27147 15216 27179
rect 15256 27147 15288 27179
rect 15328 27147 15360 27179
rect 15400 27147 15432 27179
rect 15472 27147 15504 27179
rect 15544 27147 15576 27179
rect 15616 27147 15648 27179
rect 15688 27147 15720 27179
rect 15760 27147 15792 27179
rect 15832 27147 15864 27179
rect 15904 27147 15936 27179
rect 64 27075 96 27107
rect 136 27075 168 27107
rect 208 27075 240 27107
rect 280 27075 312 27107
rect 352 27075 384 27107
rect 424 27075 456 27107
rect 496 27075 528 27107
rect 568 27075 600 27107
rect 640 27075 672 27107
rect 712 27075 744 27107
rect 784 27075 816 27107
rect 856 27075 888 27107
rect 928 27075 960 27107
rect 1000 27075 1032 27107
rect 1072 27075 1104 27107
rect 1144 27075 1176 27107
rect 1216 27075 1248 27107
rect 1288 27075 1320 27107
rect 1360 27075 1392 27107
rect 1432 27075 1464 27107
rect 1504 27075 1536 27107
rect 1576 27075 1608 27107
rect 1648 27075 1680 27107
rect 1720 27075 1752 27107
rect 1792 27075 1824 27107
rect 1864 27075 1896 27107
rect 1936 27075 1968 27107
rect 2008 27075 2040 27107
rect 2080 27075 2112 27107
rect 2152 27075 2184 27107
rect 2224 27075 2256 27107
rect 2296 27075 2328 27107
rect 2368 27075 2400 27107
rect 2440 27075 2472 27107
rect 2512 27075 2544 27107
rect 2584 27075 2616 27107
rect 2656 27075 2688 27107
rect 2728 27075 2760 27107
rect 2800 27075 2832 27107
rect 2872 27075 2904 27107
rect 2944 27075 2976 27107
rect 3016 27075 3048 27107
rect 3088 27075 3120 27107
rect 3160 27075 3192 27107
rect 3232 27075 3264 27107
rect 3304 27075 3336 27107
rect 3376 27075 3408 27107
rect 3448 27075 3480 27107
rect 3520 27075 3552 27107
rect 3592 27075 3624 27107
rect 3664 27075 3696 27107
rect 3736 27075 3768 27107
rect 3808 27075 3840 27107
rect 3880 27075 3912 27107
rect 3952 27075 3984 27107
rect 4024 27075 4056 27107
rect 4096 27075 4128 27107
rect 4168 27075 4200 27107
rect 4240 27075 4272 27107
rect 4312 27075 4344 27107
rect 4384 27075 4416 27107
rect 4456 27075 4488 27107
rect 4528 27075 4560 27107
rect 4600 27075 4632 27107
rect 4672 27075 4704 27107
rect 4744 27075 4776 27107
rect 4816 27075 4848 27107
rect 4888 27075 4920 27107
rect 4960 27075 4992 27107
rect 5032 27075 5064 27107
rect 5104 27075 5136 27107
rect 5176 27075 5208 27107
rect 5248 27075 5280 27107
rect 5320 27075 5352 27107
rect 5392 27075 5424 27107
rect 5464 27075 5496 27107
rect 5536 27075 5568 27107
rect 5608 27075 5640 27107
rect 5680 27075 5712 27107
rect 5752 27075 5784 27107
rect 5824 27075 5856 27107
rect 5896 27075 5928 27107
rect 5968 27075 6000 27107
rect 6040 27075 6072 27107
rect 6112 27075 6144 27107
rect 6184 27075 6216 27107
rect 6256 27075 6288 27107
rect 6328 27075 6360 27107
rect 6400 27075 6432 27107
rect 6472 27075 6504 27107
rect 6544 27075 6576 27107
rect 6616 27075 6648 27107
rect 6688 27075 6720 27107
rect 6760 27075 6792 27107
rect 6832 27075 6864 27107
rect 6904 27075 6936 27107
rect 6976 27075 7008 27107
rect 7048 27075 7080 27107
rect 7120 27075 7152 27107
rect 7192 27075 7224 27107
rect 7264 27075 7296 27107
rect 7336 27075 7368 27107
rect 7408 27075 7440 27107
rect 7480 27075 7512 27107
rect 7552 27075 7584 27107
rect 7624 27075 7656 27107
rect 7696 27075 7728 27107
rect 7768 27075 7800 27107
rect 7840 27075 7872 27107
rect 7912 27075 7944 27107
rect 7984 27075 8016 27107
rect 8056 27075 8088 27107
rect 8128 27075 8160 27107
rect 8200 27075 8232 27107
rect 8272 27075 8304 27107
rect 8344 27075 8376 27107
rect 8416 27075 8448 27107
rect 8488 27075 8520 27107
rect 8560 27075 8592 27107
rect 8632 27075 8664 27107
rect 8704 27075 8736 27107
rect 8776 27075 8808 27107
rect 8848 27075 8880 27107
rect 8920 27075 8952 27107
rect 8992 27075 9024 27107
rect 9064 27075 9096 27107
rect 9136 27075 9168 27107
rect 9208 27075 9240 27107
rect 9280 27075 9312 27107
rect 9352 27075 9384 27107
rect 9424 27075 9456 27107
rect 9496 27075 9528 27107
rect 9568 27075 9600 27107
rect 9640 27075 9672 27107
rect 9712 27075 9744 27107
rect 9784 27075 9816 27107
rect 9856 27075 9888 27107
rect 9928 27075 9960 27107
rect 10000 27075 10032 27107
rect 10072 27075 10104 27107
rect 10144 27075 10176 27107
rect 10216 27075 10248 27107
rect 10288 27075 10320 27107
rect 10360 27075 10392 27107
rect 10432 27075 10464 27107
rect 10504 27075 10536 27107
rect 10576 27075 10608 27107
rect 10648 27075 10680 27107
rect 10720 27075 10752 27107
rect 10792 27075 10824 27107
rect 10864 27075 10896 27107
rect 10936 27075 10968 27107
rect 11008 27075 11040 27107
rect 11080 27075 11112 27107
rect 11152 27075 11184 27107
rect 11224 27075 11256 27107
rect 11296 27075 11328 27107
rect 11368 27075 11400 27107
rect 11440 27075 11472 27107
rect 11512 27075 11544 27107
rect 11584 27075 11616 27107
rect 11656 27075 11688 27107
rect 11728 27075 11760 27107
rect 11800 27075 11832 27107
rect 11872 27075 11904 27107
rect 11944 27075 11976 27107
rect 12016 27075 12048 27107
rect 12088 27075 12120 27107
rect 12160 27075 12192 27107
rect 12232 27075 12264 27107
rect 12304 27075 12336 27107
rect 12376 27075 12408 27107
rect 12448 27075 12480 27107
rect 12520 27075 12552 27107
rect 12592 27075 12624 27107
rect 12664 27075 12696 27107
rect 12736 27075 12768 27107
rect 12808 27075 12840 27107
rect 12880 27075 12912 27107
rect 12952 27075 12984 27107
rect 13024 27075 13056 27107
rect 13096 27075 13128 27107
rect 13168 27075 13200 27107
rect 13240 27075 13272 27107
rect 13312 27075 13344 27107
rect 13384 27075 13416 27107
rect 13456 27075 13488 27107
rect 13528 27075 13560 27107
rect 13600 27075 13632 27107
rect 13672 27075 13704 27107
rect 13744 27075 13776 27107
rect 13816 27075 13848 27107
rect 13888 27075 13920 27107
rect 13960 27075 13992 27107
rect 14032 27075 14064 27107
rect 14104 27075 14136 27107
rect 14176 27075 14208 27107
rect 14248 27075 14280 27107
rect 14320 27075 14352 27107
rect 14392 27075 14424 27107
rect 14464 27075 14496 27107
rect 14536 27075 14568 27107
rect 14608 27075 14640 27107
rect 14680 27075 14712 27107
rect 14752 27075 14784 27107
rect 14824 27075 14856 27107
rect 14896 27075 14928 27107
rect 14968 27075 15000 27107
rect 15040 27075 15072 27107
rect 15112 27075 15144 27107
rect 15184 27075 15216 27107
rect 15256 27075 15288 27107
rect 15328 27075 15360 27107
rect 15400 27075 15432 27107
rect 15472 27075 15504 27107
rect 15544 27075 15576 27107
rect 15616 27075 15648 27107
rect 15688 27075 15720 27107
rect 15760 27075 15792 27107
rect 15832 27075 15864 27107
rect 15904 27075 15936 27107
rect 64 27003 96 27035
rect 136 27003 168 27035
rect 208 27003 240 27035
rect 280 27003 312 27035
rect 352 27003 384 27035
rect 424 27003 456 27035
rect 496 27003 528 27035
rect 568 27003 600 27035
rect 640 27003 672 27035
rect 712 27003 744 27035
rect 784 27003 816 27035
rect 856 27003 888 27035
rect 928 27003 960 27035
rect 1000 27003 1032 27035
rect 1072 27003 1104 27035
rect 1144 27003 1176 27035
rect 1216 27003 1248 27035
rect 1288 27003 1320 27035
rect 1360 27003 1392 27035
rect 1432 27003 1464 27035
rect 1504 27003 1536 27035
rect 1576 27003 1608 27035
rect 1648 27003 1680 27035
rect 1720 27003 1752 27035
rect 1792 27003 1824 27035
rect 1864 27003 1896 27035
rect 1936 27003 1968 27035
rect 2008 27003 2040 27035
rect 2080 27003 2112 27035
rect 2152 27003 2184 27035
rect 2224 27003 2256 27035
rect 2296 27003 2328 27035
rect 2368 27003 2400 27035
rect 2440 27003 2472 27035
rect 2512 27003 2544 27035
rect 2584 27003 2616 27035
rect 2656 27003 2688 27035
rect 2728 27003 2760 27035
rect 2800 27003 2832 27035
rect 2872 27003 2904 27035
rect 2944 27003 2976 27035
rect 3016 27003 3048 27035
rect 3088 27003 3120 27035
rect 3160 27003 3192 27035
rect 3232 27003 3264 27035
rect 3304 27003 3336 27035
rect 3376 27003 3408 27035
rect 3448 27003 3480 27035
rect 3520 27003 3552 27035
rect 3592 27003 3624 27035
rect 3664 27003 3696 27035
rect 3736 27003 3768 27035
rect 3808 27003 3840 27035
rect 3880 27003 3912 27035
rect 3952 27003 3984 27035
rect 4024 27003 4056 27035
rect 4096 27003 4128 27035
rect 4168 27003 4200 27035
rect 4240 27003 4272 27035
rect 4312 27003 4344 27035
rect 4384 27003 4416 27035
rect 4456 27003 4488 27035
rect 4528 27003 4560 27035
rect 4600 27003 4632 27035
rect 4672 27003 4704 27035
rect 4744 27003 4776 27035
rect 4816 27003 4848 27035
rect 4888 27003 4920 27035
rect 4960 27003 4992 27035
rect 5032 27003 5064 27035
rect 5104 27003 5136 27035
rect 5176 27003 5208 27035
rect 5248 27003 5280 27035
rect 5320 27003 5352 27035
rect 5392 27003 5424 27035
rect 5464 27003 5496 27035
rect 5536 27003 5568 27035
rect 5608 27003 5640 27035
rect 5680 27003 5712 27035
rect 5752 27003 5784 27035
rect 5824 27003 5856 27035
rect 5896 27003 5928 27035
rect 5968 27003 6000 27035
rect 6040 27003 6072 27035
rect 6112 27003 6144 27035
rect 6184 27003 6216 27035
rect 6256 27003 6288 27035
rect 6328 27003 6360 27035
rect 6400 27003 6432 27035
rect 6472 27003 6504 27035
rect 6544 27003 6576 27035
rect 6616 27003 6648 27035
rect 6688 27003 6720 27035
rect 6760 27003 6792 27035
rect 6832 27003 6864 27035
rect 6904 27003 6936 27035
rect 6976 27003 7008 27035
rect 7048 27003 7080 27035
rect 7120 27003 7152 27035
rect 7192 27003 7224 27035
rect 7264 27003 7296 27035
rect 7336 27003 7368 27035
rect 7408 27003 7440 27035
rect 7480 27003 7512 27035
rect 7552 27003 7584 27035
rect 7624 27003 7656 27035
rect 7696 27003 7728 27035
rect 7768 27003 7800 27035
rect 7840 27003 7872 27035
rect 7912 27003 7944 27035
rect 7984 27003 8016 27035
rect 8056 27003 8088 27035
rect 8128 27003 8160 27035
rect 8200 27003 8232 27035
rect 8272 27003 8304 27035
rect 8344 27003 8376 27035
rect 8416 27003 8448 27035
rect 8488 27003 8520 27035
rect 8560 27003 8592 27035
rect 8632 27003 8664 27035
rect 8704 27003 8736 27035
rect 8776 27003 8808 27035
rect 8848 27003 8880 27035
rect 8920 27003 8952 27035
rect 8992 27003 9024 27035
rect 9064 27003 9096 27035
rect 9136 27003 9168 27035
rect 9208 27003 9240 27035
rect 9280 27003 9312 27035
rect 9352 27003 9384 27035
rect 9424 27003 9456 27035
rect 9496 27003 9528 27035
rect 9568 27003 9600 27035
rect 9640 27003 9672 27035
rect 9712 27003 9744 27035
rect 9784 27003 9816 27035
rect 9856 27003 9888 27035
rect 9928 27003 9960 27035
rect 10000 27003 10032 27035
rect 10072 27003 10104 27035
rect 10144 27003 10176 27035
rect 10216 27003 10248 27035
rect 10288 27003 10320 27035
rect 10360 27003 10392 27035
rect 10432 27003 10464 27035
rect 10504 27003 10536 27035
rect 10576 27003 10608 27035
rect 10648 27003 10680 27035
rect 10720 27003 10752 27035
rect 10792 27003 10824 27035
rect 10864 27003 10896 27035
rect 10936 27003 10968 27035
rect 11008 27003 11040 27035
rect 11080 27003 11112 27035
rect 11152 27003 11184 27035
rect 11224 27003 11256 27035
rect 11296 27003 11328 27035
rect 11368 27003 11400 27035
rect 11440 27003 11472 27035
rect 11512 27003 11544 27035
rect 11584 27003 11616 27035
rect 11656 27003 11688 27035
rect 11728 27003 11760 27035
rect 11800 27003 11832 27035
rect 11872 27003 11904 27035
rect 11944 27003 11976 27035
rect 12016 27003 12048 27035
rect 12088 27003 12120 27035
rect 12160 27003 12192 27035
rect 12232 27003 12264 27035
rect 12304 27003 12336 27035
rect 12376 27003 12408 27035
rect 12448 27003 12480 27035
rect 12520 27003 12552 27035
rect 12592 27003 12624 27035
rect 12664 27003 12696 27035
rect 12736 27003 12768 27035
rect 12808 27003 12840 27035
rect 12880 27003 12912 27035
rect 12952 27003 12984 27035
rect 13024 27003 13056 27035
rect 13096 27003 13128 27035
rect 13168 27003 13200 27035
rect 13240 27003 13272 27035
rect 13312 27003 13344 27035
rect 13384 27003 13416 27035
rect 13456 27003 13488 27035
rect 13528 27003 13560 27035
rect 13600 27003 13632 27035
rect 13672 27003 13704 27035
rect 13744 27003 13776 27035
rect 13816 27003 13848 27035
rect 13888 27003 13920 27035
rect 13960 27003 13992 27035
rect 14032 27003 14064 27035
rect 14104 27003 14136 27035
rect 14176 27003 14208 27035
rect 14248 27003 14280 27035
rect 14320 27003 14352 27035
rect 14392 27003 14424 27035
rect 14464 27003 14496 27035
rect 14536 27003 14568 27035
rect 14608 27003 14640 27035
rect 14680 27003 14712 27035
rect 14752 27003 14784 27035
rect 14824 27003 14856 27035
rect 14896 27003 14928 27035
rect 14968 27003 15000 27035
rect 15040 27003 15072 27035
rect 15112 27003 15144 27035
rect 15184 27003 15216 27035
rect 15256 27003 15288 27035
rect 15328 27003 15360 27035
rect 15400 27003 15432 27035
rect 15472 27003 15504 27035
rect 15544 27003 15576 27035
rect 15616 27003 15648 27035
rect 15688 27003 15720 27035
rect 15760 27003 15792 27035
rect 15832 27003 15864 27035
rect 15904 27003 15936 27035
rect 64 26931 96 26963
rect 136 26931 168 26963
rect 208 26931 240 26963
rect 280 26931 312 26963
rect 352 26931 384 26963
rect 424 26931 456 26963
rect 496 26931 528 26963
rect 568 26931 600 26963
rect 640 26931 672 26963
rect 712 26931 744 26963
rect 784 26931 816 26963
rect 856 26931 888 26963
rect 928 26931 960 26963
rect 1000 26931 1032 26963
rect 1072 26931 1104 26963
rect 1144 26931 1176 26963
rect 1216 26931 1248 26963
rect 1288 26931 1320 26963
rect 1360 26931 1392 26963
rect 1432 26931 1464 26963
rect 1504 26931 1536 26963
rect 1576 26931 1608 26963
rect 1648 26931 1680 26963
rect 1720 26931 1752 26963
rect 1792 26931 1824 26963
rect 1864 26931 1896 26963
rect 1936 26931 1968 26963
rect 2008 26931 2040 26963
rect 2080 26931 2112 26963
rect 2152 26931 2184 26963
rect 2224 26931 2256 26963
rect 2296 26931 2328 26963
rect 2368 26931 2400 26963
rect 2440 26931 2472 26963
rect 2512 26931 2544 26963
rect 2584 26931 2616 26963
rect 2656 26931 2688 26963
rect 2728 26931 2760 26963
rect 2800 26931 2832 26963
rect 2872 26931 2904 26963
rect 2944 26931 2976 26963
rect 3016 26931 3048 26963
rect 3088 26931 3120 26963
rect 3160 26931 3192 26963
rect 3232 26931 3264 26963
rect 3304 26931 3336 26963
rect 3376 26931 3408 26963
rect 3448 26931 3480 26963
rect 3520 26931 3552 26963
rect 3592 26931 3624 26963
rect 3664 26931 3696 26963
rect 3736 26931 3768 26963
rect 3808 26931 3840 26963
rect 3880 26931 3912 26963
rect 3952 26931 3984 26963
rect 4024 26931 4056 26963
rect 4096 26931 4128 26963
rect 4168 26931 4200 26963
rect 4240 26931 4272 26963
rect 4312 26931 4344 26963
rect 4384 26931 4416 26963
rect 4456 26931 4488 26963
rect 4528 26931 4560 26963
rect 4600 26931 4632 26963
rect 4672 26931 4704 26963
rect 4744 26931 4776 26963
rect 4816 26931 4848 26963
rect 4888 26931 4920 26963
rect 4960 26931 4992 26963
rect 5032 26931 5064 26963
rect 5104 26931 5136 26963
rect 5176 26931 5208 26963
rect 5248 26931 5280 26963
rect 5320 26931 5352 26963
rect 5392 26931 5424 26963
rect 5464 26931 5496 26963
rect 5536 26931 5568 26963
rect 5608 26931 5640 26963
rect 5680 26931 5712 26963
rect 5752 26931 5784 26963
rect 5824 26931 5856 26963
rect 5896 26931 5928 26963
rect 5968 26931 6000 26963
rect 6040 26931 6072 26963
rect 6112 26931 6144 26963
rect 6184 26931 6216 26963
rect 6256 26931 6288 26963
rect 6328 26931 6360 26963
rect 6400 26931 6432 26963
rect 6472 26931 6504 26963
rect 6544 26931 6576 26963
rect 6616 26931 6648 26963
rect 6688 26931 6720 26963
rect 6760 26931 6792 26963
rect 6832 26931 6864 26963
rect 6904 26931 6936 26963
rect 6976 26931 7008 26963
rect 7048 26931 7080 26963
rect 7120 26931 7152 26963
rect 7192 26931 7224 26963
rect 7264 26931 7296 26963
rect 7336 26931 7368 26963
rect 7408 26931 7440 26963
rect 7480 26931 7512 26963
rect 7552 26931 7584 26963
rect 7624 26931 7656 26963
rect 7696 26931 7728 26963
rect 7768 26931 7800 26963
rect 7840 26931 7872 26963
rect 7912 26931 7944 26963
rect 7984 26931 8016 26963
rect 8056 26931 8088 26963
rect 8128 26931 8160 26963
rect 8200 26931 8232 26963
rect 8272 26931 8304 26963
rect 8344 26931 8376 26963
rect 8416 26931 8448 26963
rect 8488 26931 8520 26963
rect 8560 26931 8592 26963
rect 8632 26931 8664 26963
rect 8704 26931 8736 26963
rect 8776 26931 8808 26963
rect 8848 26931 8880 26963
rect 8920 26931 8952 26963
rect 8992 26931 9024 26963
rect 9064 26931 9096 26963
rect 9136 26931 9168 26963
rect 9208 26931 9240 26963
rect 9280 26931 9312 26963
rect 9352 26931 9384 26963
rect 9424 26931 9456 26963
rect 9496 26931 9528 26963
rect 9568 26931 9600 26963
rect 9640 26931 9672 26963
rect 9712 26931 9744 26963
rect 9784 26931 9816 26963
rect 9856 26931 9888 26963
rect 9928 26931 9960 26963
rect 10000 26931 10032 26963
rect 10072 26931 10104 26963
rect 10144 26931 10176 26963
rect 10216 26931 10248 26963
rect 10288 26931 10320 26963
rect 10360 26931 10392 26963
rect 10432 26931 10464 26963
rect 10504 26931 10536 26963
rect 10576 26931 10608 26963
rect 10648 26931 10680 26963
rect 10720 26931 10752 26963
rect 10792 26931 10824 26963
rect 10864 26931 10896 26963
rect 10936 26931 10968 26963
rect 11008 26931 11040 26963
rect 11080 26931 11112 26963
rect 11152 26931 11184 26963
rect 11224 26931 11256 26963
rect 11296 26931 11328 26963
rect 11368 26931 11400 26963
rect 11440 26931 11472 26963
rect 11512 26931 11544 26963
rect 11584 26931 11616 26963
rect 11656 26931 11688 26963
rect 11728 26931 11760 26963
rect 11800 26931 11832 26963
rect 11872 26931 11904 26963
rect 11944 26931 11976 26963
rect 12016 26931 12048 26963
rect 12088 26931 12120 26963
rect 12160 26931 12192 26963
rect 12232 26931 12264 26963
rect 12304 26931 12336 26963
rect 12376 26931 12408 26963
rect 12448 26931 12480 26963
rect 12520 26931 12552 26963
rect 12592 26931 12624 26963
rect 12664 26931 12696 26963
rect 12736 26931 12768 26963
rect 12808 26931 12840 26963
rect 12880 26931 12912 26963
rect 12952 26931 12984 26963
rect 13024 26931 13056 26963
rect 13096 26931 13128 26963
rect 13168 26931 13200 26963
rect 13240 26931 13272 26963
rect 13312 26931 13344 26963
rect 13384 26931 13416 26963
rect 13456 26931 13488 26963
rect 13528 26931 13560 26963
rect 13600 26931 13632 26963
rect 13672 26931 13704 26963
rect 13744 26931 13776 26963
rect 13816 26931 13848 26963
rect 13888 26931 13920 26963
rect 13960 26931 13992 26963
rect 14032 26931 14064 26963
rect 14104 26931 14136 26963
rect 14176 26931 14208 26963
rect 14248 26931 14280 26963
rect 14320 26931 14352 26963
rect 14392 26931 14424 26963
rect 14464 26931 14496 26963
rect 14536 26931 14568 26963
rect 14608 26931 14640 26963
rect 14680 26931 14712 26963
rect 14752 26931 14784 26963
rect 14824 26931 14856 26963
rect 14896 26931 14928 26963
rect 14968 26931 15000 26963
rect 15040 26931 15072 26963
rect 15112 26931 15144 26963
rect 15184 26931 15216 26963
rect 15256 26931 15288 26963
rect 15328 26931 15360 26963
rect 15400 26931 15432 26963
rect 15472 26931 15504 26963
rect 15544 26931 15576 26963
rect 15616 26931 15648 26963
rect 15688 26931 15720 26963
rect 15760 26931 15792 26963
rect 15832 26931 15864 26963
rect 15904 26931 15936 26963
rect 64 26859 96 26891
rect 136 26859 168 26891
rect 208 26859 240 26891
rect 280 26859 312 26891
rect 352 26859 384 26891
rect 424 26859 456 26891
rect 496 26859 528 26891
rect 568 26859 600 26891
rect 640 26859 672 26891
rect 712 26859 744 26891
rect 784 26859 816 26891
rect 856 26859 888 26891
rect 928 26859 960 26891
rect 1000 26859 1032 26891
rect 1072 26859 1104 26891
rect 1144 26859 1176 26891
rect 1216 26859 1248 26891
rect 1288 26859 1320 26891
rect 1360 26859 1392 26891
rect 1432 26859 1464 26891
rect 1504 26859 1536 26891
rect 1576 26859 1608 26891
rect 1648 26859 1680 26891
rect 1720 26859 1752 26891
rect 1792 26859 1824 26891
rect 1864 26859 1896 26891
rect 1936 26859 1968 26891
rect 2008 26859 2040 26891
rect 2080 26859 2112 26891
rect 2152 26859 2184 26891
rect 2224 26859 2256 26891
rect 2296 26859 2328 26891
rect 2368 26859 2400 26891
rect 2440 26859 2472 26891
rect 2512 26859 2544 26891
rect 2584 26859 2616 26891
rect 2656 26859 2688 26891
rect 2728 26859 2760 26891
rect 2800 26859 2832 26891
rect 2872 26859 2904 26891
rect 2944 26859 2976 26891
rect 3016 26859 3048 26891
rect 3088 26859 3120 26891
rect 3160 26859 3192 26891
rect 3232 26859 3264 26891
rect 3304 26859 3336 26891
rect 3376 26859 3408 26891
rect 3448 26859 3480 26891
rect 3520 26859 3552 26891
rect 3592 26859 3624 26891
rect 3664 26859 3696 26891
rect 3736 26859 3768 26891
rect 3808 26859 3840 26891
rect 3880 26859 3912 26891
rect 3952 26859 3984 26891
rect 4024 26859 4056 26891
rect 4096 26859 4128 26891
rect 4168 26859 4200 26891
rect 4240 26859 4272 26891
rect 4312 26859 4344 26891
rect 4384 26859 4416 26891
rect 4456 26859 4488 26891
rect 4528 26859 4560 26891
rect 4600 26859 4632 26891
rect 4672 26859 4704 26891
rect 4744 26859 4776 26891
rect 4816 26859 4848 26891
rect 4888 26859 4920 26891
rect 4960 26859 4992 26891
rect 5032 26859 5064 26891
rect 5104 26859 5136 26891
rect 5176 26859 5208 26891
rect 5248 26859 5280 26891
rect 5320 26859 5352 26891
rect 5392 26859 5424 26891
rect 5464 26859 5496 26891
rect 5536 26859 5568 26891
rect 5608 26859 5640 26891
rect 5680 26859 5712 26891
rect 5752 26859 5784 26891
rect 5824 26859 5856 26891
rect 5896 26859 5928 26891
rect 5968 26859 6000 26891
rect 6040 26859 6072 26891
rect 6112 26859 6144 26891
rect 6184 26859 6216 26891
rect 6256 26859 6288 26891
rect 6328 26859 6360 26891
rect 6400 26859 6432 26891
rect 6472 26859 6504 26891
rect 6544 26859 6576 26891
rect 6616 26859 6648 26891
rect 6688 26859 6720 26891
rect 6760 26859 6792 26891
rect 6832 26859 6864 26891
rect 6904 26859 6936 26891
rect 6976 26859 7008 26891
rect 7048 26859 7080 26891
rect 7120 26859 7152 26891
rect 7192 26859 7224 26891
rect 7264 26859 7296 26891
rect 7336 26859 7368 26891
rect 7408 26859 7440 26891
rect 7480 26859 7512 26891
rect 7552 26859 7584 26891
rect 7624 26859 7656 26891
rect 7696 26859 7728 26891
rect 7768 26859 7800 26891
rect 7840 26859 7872 26891
rect 7912 26859 7944 26891
rect 7984 26859 8016 26891
rect 8056 26859 8088 26891
rect 8128 26859 8160 26891
rect 8200 26859 8232 26891
rect 8272 26859 8304 26891
rect 8344 26859 8376 26891
rect 8416 26859 8448 26891
rect 8488 26859 8520 26891
rect 8560 26859 8592 26891
rect 8632 26859 8664 26891
rect 8704 26859 8736 26891
rect 8776 26859 8808 26891
rect 8848 26859 8880 26891
rect 8920 26859 8952 26891
rect 8992 26859 9024 26891
rect 9064 26859 9096 26891
rect 9136 26859 9168 26891
rect 9208 26859 9240 26891
rect 9280 26859 9312 26891
rect 9352 26859 9384 26891
rect 9424 26859 9456 26891
rect 9496 26859 9528 26891
rect 9568 26859 9600 26891
rect 9640 26859 9672 26891
rect 9712 26859 9744 26891
rect 9784 26859 9816 26891
rect 9856 26859 9888 26891
rect 9928 26859 9960 26891
rect 10000 26859 10032 26891
rect 10072 26859 10104 26891
rect 10144 26859 10176 26891
rect 10216 26859 10248 26891
rect 10288 26859 10320 26891
rect 10360 26859 10392 26891
rect 10432 26859 10464 26891
rect 10504 26859 10536 26891
rect 10576 26859 10608 26891
rect 10648 26859 10680 26891
rect 10720 26859 10752 26891
rect 10792 26859 10824 26891
rect 10864 26859 10896 26891
rect 10936 26859 10968 26891
rect 11008 26859 11040 26891
rect 11080 26859 11112 26891
rect 11152 26859 11184 26891
rect 11224 26859 11256 26891
rect 11296 26859 11328 26891
rect 11368 26859 11400 26891
rect 11440 26859 11472 26891
rect 11512 26859 11544 26891
rect 11584 26859 11616 26891
rect 11656 26859 11688 26891
rect 11728 26859 11760 26891
rect 11800 26859 11832 26891
rect 11872 26859 11904 26891
rect 11944 26859 11976 26891
rect 12016 26859 12048 26891
rect 12088 26859 12120 26891
rect 12160 26859 12192 26891
rect 12232 26859 12264 26891
rect 12304 26859 12336 26891
rect 12376 26859 12408 26891
rect 12448 26859 12480 26891
rect 12520 26859 12552 26891
rect 12592 26859 12624 26891
rect 12664 26859 12696 26891
rect 12736 26859 12768 26891
rect 12808 26859 12840 26891
rect 12880 26859 12912 26891
rect 12952 26859 12984 26891
rect 13024 26859 13056 26891
rect 13096 26859 13128 26891
rect 13168 26859 13200 26891
rect 13240 26859 13272 26891
rect 13312 26859 13344 26891
rect 13384 26859 13416 26891
rect 13456 26859 13488 26891
rect 13528 26859 13560 26891
rect 13600 26859 13632 26891
rect 13672 26859 13704 26891
rect 13744 26859 13776 26891
rect 13816 26859 13848 26891
rect 13888 26859 13920 26891
rect 13960 26859 13992 26891
rect 14032 26859 14064 26891
rect 14104 26859 14136 26891
rect 14176 26859 14208 26891
rect 14248 26859 14280 26891
rect 14320 26859 14352 26891
rect 14392 26859 14424 26891
rect 14464 26859 14496 26891
rect 14536 26859 14568 26891
rect 14608 26859 14640 26891
rect 14680 26859 14712 26891
rect 14752 26859 14784 26891
rect 14824 26859 14856 26891
rect 14896 26859 14928 26891
rect 14968 26859 15000 26891
rect 15040 26859 15072 26891
rect 15112 26859 15144 26891
rect 15184 26859 15216 26891
rect 15256 26859 15288 26891
rect 15328 26859 15360 26891
rect 15400 26859 15432 26891
rect 15472 26859 15504 26891
rect 15544 26859 15576 26891
rect 15616 26859 15648 26891
rect 15688 26859 15720 26891
rect 15760 26859 15792 26891
rect 15832 26859 15864 26891
rect 15904 26859 15936 26891
rect 64 26787 96 26819
rect 136 26787 168 26819
rect 208 26787 240 26819
rect 280 26787 312 26819
rect 352 26787 384 26819
rect 424 26787 456 26819
rect 496 26787 528 26819
rect 568 26787 600 26819
rect 640 26787 672 26819
rect 712 26787 744 26819
rect 784 26787 816 26819
rect 856 26787 888 26819
rect 928 26787 960 26819
rect 1000 26787 1032 26819
rect 1072 26787 1104 26819
rect 1144 26787 1176 26819
rect 1216 26787 1248 26819
rect 1288 26787 1320 26819
rect 1360 26787 1392 26819
rect 1432 26787 1464 26819
rect 1504 26787 1536 26819
rect 1576 26787 1608 26819
rect 1648 26787 1680 26819
rect 1720 26787 1752 26819
rect 1792 26787 1824 26819
rect 1864 26787 1896 26819
rect 1936 26787 1968 26819
rect 2008 26787 2040 26819
rect 2080 26787 2112 26819
rect 2152 26787 2184 26819
rect 2224 26787 2256 26819
rect 2296 26787 2328 26819
rect 2368 26787 2400 26819
rect 2440 26787 2472 26819
rect 2512 26787 2544 26819
rect 2584 26787 2616 26819
rect 2656 26787 2688 26819
rect 2728 26787 2760 26819
rect 2800 26787 2832 26819
rect 2872 26787 2904 26819
rect 2944 26787 2976 26819
rect 3016 26787 3048 26819
rect 3088 26787 3120 26819
rect 3160 26787 3192 26819
rect 3232 26787 3264 26819
rect 3304 26787 3336 26819
rect 3376 26787 3408 26819
rect 3448 26787 3480 26819
rect 3520 26787 3552 26819
rect 3592 26787 3624 26819
rect 3664 26787 3696 26819
rect 3736 26787 3768 26819
rect 3808 26787 3840 26819
rect 3880 26787 3912 26819
rect 3952 26787 3984 26819
rect 4024 26787 4056 26819
rect 4096 26787 4128 26819
rect 4168 26787 4200 26819
rect 4240 26787 4272 26819
rect 4312 26787 4344 26819
rect 4384 26787 4416 26819
rect 4456 26787 4488 26819
rect 4528 26787 4560 26819
rect 4600 26787 4632 26819
rect 4672 26787 4704 26819
rect 4744 26787 4776 26819
rect 4816 26787 4848 26819
rect 4888 26787 4920 26819
rect 4960 26787 4992 26819
rect 5032 26787 5064 26819
rect 5104 26787 5136 26819
rect 5176 26787 5208 26819
rect 5248 26787 5280 26819
rect 5320 26787 5352 26819
rect 5392 26787 5424 26819
rect 5464 26787 5496 26819
rect 5536 26787 5568 26819
rect 5608 26787 5640 26819
rect 5680 26787 5712 26819
rect 5752 26787 5784 26819
rect 5824 26787 5856 26819
rect 5896 26787 5928 26819
rect 5968 26787 6000 26819
rect 6040 26787 6072 26819
rect 6112 26787 6144 26819
rect 6184 26787 6216 26819
rect 6256 26787 6288 26819
rect 6328 26787 6360 26819
rect 6400 26787 6432 26819
rect 6472 26787 6504 26819
rect 6544 26787 6576 26819
rect 6616 26787 6648 26819
rect 6688 26787 6720 26819
rect 6760 26787 6792 26819
rect 6832 26787 6864 26819
rect 6904 26787 6936 26819
rect 6976 26787 7008 26819
rect 7048 26787 7080 26819
rect 7120 26787 7152 26819
rect 7192 26787 7224 26819
rect 7264 26787 7296 26819
rect 7336 26787 7368 26819
rect 7408 26787 7440 26819
rect 7480 26787 7512 26819
rect 7552 26787 7584 26819
rect 7624 26787 7656 26819
rect 7696 26787 7728 26819
rect 7768 26787 7800 26819
rect 7840 26787 7872 26819
rect 7912 26787 7944 26819
rect 7984 26787 8016 26819
rect 8056 26787 8088 26819
rect 8128 26787 8160 26819
rect 8200 26787 8232 26819
rect 8272 26787 8304 26819
rect 8344 26787 8376 26819
rect 8416 26787 8448 26819
rect 8488 26787 8520 26819
rect 8560 26787 8592 26819
rect 8632 26787 8664 26819
rect 8704 26787 8736 26819
rect 8776 26787 8808 26819
rect 8848 26787 8880 26819
rect 8920 26787 8952 26819
rect 8992 26787 9024 26819
rect 9064 26787 9096 26819
rect 9136 26787 9168 26819
rect 9208 26787 9240 26819
rect 9280 26787 9312 26819
rect 9352 26787 9384 26819
rect 9424 26787 9456 26819
rect 9496 26787 9528 26819
rect 9568 26787 9600 26819
rect 9640 26787 9672 26819
rect 9712 26787 9744 26819
rect 9784 26787 9816 26819
rect 9856 26787 9888 26819
rect 9928 26787 9960 26819
rect 10000 26787 10032 26819
rect 10072 26787 10104 26819
rect 10144 26787 10176 26819
rect 10216 26787 10248 26819
rect 10288 26787 10320 26819
rect 10360 26787 10392 26819
rect 10432 26787 10464 26819
rect 10504 26787 10536 26819
rect 10576 26787 10608 26819
rect 10648 26787 10680 26819
rect 10720 26787 10752 26819
rect 10792 26787 10824 26819
rect 10864 26787 10896 26819
rect 10936 26787 10968 26819
rect 11008 26787 11040 26819
rect 11080 26787 11112 26819
rect 11152 26787 11184 26819
rect 11224 26787 11256 26819
rect 11296 26787 11328 26819
rect 11368 26787 11400 26819
rect 11440 26787 11472 26819
rect 11512 26787 11544 26819
rect 11584 26787 11616 26819
rect 11656 26787 11688 26819
rect 11728 26787 11760 26819
rect 11800 26787 11832 26819
rect 11872 26787 11904 26819
rect 11944 26787 11976 26819
rect 12016 26787 12048 26819
rect 12088 26787 12120 26819
rect 12160 26787 12192 26819
rect 12232 26787 12264 26819
rect 12304 26787 12336 26819
rect 12376 26787 12408 26819
rect 12448 26787 12480 26819
rect 12520 26787 12552 26819
rect 12592 26787 12624 26819
rect 12664 26787 12696 26819
rect 12736 26787 12768 26819
rect 12808 26787 12840 26819
rect 12880 26787 12912 26819
rect 12952 26787 12984 26819
rect 13024 26787 13056 26819
rect 13096 26787 13128 26819
rect 13168 26787 13200 26819
rect 13240 26787 13272 26819
rect 13312 26787 13344 26819
rect 13384 26787 13416 26819
rect 13456 26787 13488 26819
rect 13528 26787 13560 26819
rect 13600 26787 13632 26819
rect 13672 26787 13704 26819
rect 13744 26787 13776 26819
rect 13816 26787 13848 26819
rect 13888 26787 13920 26819
rect 13960 26787 13992 26819
rect 14032 26787 14064 26819
rect 14104 26787 14136 26819
rect 14176 26787 14208 26819
rect 14248 26787 14280 26819
rect 14320 26787 14352 26819
rect 14392 26787 14424 26819
rect 14464 26787 14496 26819
rect 14536 26787 14568 26819
rect 14608 26787 14640 26819
rect 14680 26787 14712 26819
rect 14752 26787 14784 26819
rect 14824 26787 14856 26819
rect 14896 26787 14928 26819
rect 14968 26787 15000 26819
rect 15040 26787 15072 26819
rect 15112 26787 15144 26819
rect 15184 26787 15216 26819
rect 15256 26787 15288 26819
rect 15328 26787 15360 26819
rect 15400 26787 15432 26819
rect 15472 26787 15504 26819
rect 15544 26787 15576 26819
rect 15616 26787 15648 26819
rect 15688 26787 15720 26819
rect 15760 26787 15792 26819
rect 15832 26787 15864 26819
rect 15904 26787 15936 26819
rect 64 26715 96 26747
rect 136 26715 168 26747
rect 208 26715 240 26747
rect 280 26715 312 26747
rect 352 26715 384 26747
rect 424 26715 456 26747
rect 496 26715 528 26747
rect 568 26715 600 26747
rect 640 26715 672 26747
rect 712 26715 744 26747
rect 784 26715 816 26747
rect 856 26715 888 26747
rect 928 26715 960 26747
rect 1000 26715 1032 26747
rect 1072 26715 1104 26747
rect 1144 26715 1176 26747
rect 1216 26715 1248 26747
rect 1288 26715 1320 26747
rect 1360 26715 1392 26747
rect 1432 26715 1464 26747
rect 1504 26715 1536 26747
rect 1576 26715 1608 26747
rect 1648 26715 1680 26747
rect 1720 26715 1752 26747
rect 1792 26715 1824 26747
rect 1864 26715 1896 26747
rect 1936 26715 1968 26747
rect 2008 26715 2040 26747
rect 2080 26715 2112 26747
rect 2152 26715 2184 26747
rect 2224 26715 2256 26747
rect 2296 26715 2328 26747
rect 2368 26715 2400 26747
rect 2440 26715 2472 26747
rect 2512 26715 2544 26747
rect 2584 26715 2616 26747
rect 2656 26715 2688 26747
rect 2728 26715 2760 26747
rect 2800 26715 2832 26747
rect 2872 26715 2904 26747
rect 2944 26715 2976 26747
rect 3016 26715 3048 26747
rect 3088 26715 3120 26747
rect 3160 26715 3192 26747
rect 3232 26715 3264 26747
rect 3304 26715 3336 26747
rect 3376 26715 3408 26747
rect 3448 26715 3480 26747
rect 3520 26715 3552 26747
rect 3592 26715 3624 26747
rect 3664 26715 3696 26747
rect 3736 26715 3768 26747
rect 3808 26715 3840 26747
rect 3880 26715 3912 26747
rect 3952 26715 3984 26747
rect 4024 26715 4056 26747
rect 4096 26715 4128 26747
rect 4168 26715 4200 26747
rect 4240 26715 4272 26747
rect 4312 26715 4344 26747
rect 4384 26715 4416 26747
rect 4456 26715 4488 26747
rect 4528 26715 4560 26747
rect 4600 26715 4632 26747
rect 4672 26715 4704 26747
rect 4744 26715 4776 26747
rect 4816 26715 4848 26747
rect 4888 26715 4920 26747
rect 4960 26715 4992 26747
rect 5032 26715 5064 26747
rect 5104 26715 5136 26747
rect 5176 26715 5208 26747
rect 5248 26715 5280 26747
rect 5320 26715 5352 26747
rect 5392 26715 5424 26747
rect 5464 26715 5496 26747
rect 5536 26715 5568 26747
rect 5608 26715 5640 26747
rect 5680 26715 5712 26747
rect 5752 26715 5784 26747
rect 5824 26715 5856 26747
rect 5896 26715 5928 26747
rect 5968 26715 6000 26747
rect 6040 26715 6072 26747
rect 6112 26715 6144 26747
rect 6184 26715 6216 26747
rect 6256 26715 6288 26747
rect 6328 26715 6360 26747
rect 6400 26715 6432 26747
rect 6472 26715 6504 26747
rect 6544 26715 6576 26747
rect 6616 26715 6648 26747
rect 6688 26715 6720 26747
rect 6760 26715 6792 26747
rect 6832 26715 6864 26747
rect 6904 26715 6936 26747
rect 6976 26715 7008 26747
rect 7048 26715 7080 26747
rect 7120 26715 7152 26747
rect 7192 26715 7224 26747
rect 7264 26715 7296 26747
rect 7336 26715 7368 26747
rect 7408 26715 7440 26747
rect 7480 26715 7512 26747
rect 7552 26715 7584 26747
rect 7624 26715 7656 26747
rect 7696 26715 7728 26747
rect 7768 26715 7800 26747
rect 7840 26715 7872 26747
rect 7912 26715 7944 26747
rect 7984 26715 8016 26747
rect 8056 26715 8088 26747
rect 8128 26715 8160 26747
rect 8200 26715 8232 26747
rect 8272 26715 8304 26747
rect 8344 26715 8376 26747
rect 8416 26715 8448 26747
rect 8488 26715 8520 26747
rect 8560 26715 8592 26747
rect 8632 26715 8664 26747
rect 8704 26715 8736 26747
rect 8776 26715 8808 26747
rect 8848 26715 8880 26747
rect 8920 26715 8952 26747
rect 8992 26715 9024 26747
rect 9064 26715 9096 26747
rect 9136 26715 9168 26747
rect 9208 26715 9240 26747
rect 9280 26715 9312 26747
rect 9352 26715 9384 26747
rect 9424 26715 9456 26747
rect 9496 26715 9528 26747
rect 9568 26715 9600 26747
rect 9640 26715 9672 26747
rect 9712 26715 9744 26747
rect 9784 26715 9816 26747
rect 9856 26715 9888 26747
rect 9928 26715 9960 26747
rect 10000 26715 10032 26747
rect 10072 26715 10104 26747
rect 10144 26715 10176 26747
rect 10216 26715 10248 26747
rect 10288 26715 10320 26747
rect 10360 26715 10392 26747
rect 10432 26715 10464 26747
rect 10504 26715 10536 26747
rect 10576 26715 10608 26747
rect 10648 26715 10680 26747
rect 10720 26715 10752 26747
rect 10792 26715 10824 26747
rect 10864 26715 10896 26747
rect 10936 26715 10968 26747
rect 11008 26715 11040 26747
rect 11080 26715 11112 26747
rect 11152 26715 11184 26747
rect 11224 26715 11256 26747
rect 11296 26715 11328 26747
rect 11368 26715 11400 26747
rect 11440 26715 11472 26747
rect 11512 26715 11544 26747
rect 11584 26715 11616 26747
rect 11656 26715 11688 26747
rect 11728 26715 11760 26747
rect 11800 26715 11832 26747
rect 11872 26715 11904 26747
rect 11944 26715 11976 26747
rect 12016 26715 12048 26747
rect 12088 26715 12120 26747
rect 12160 26715 12192 26747
rect 12232 26715 12264 26747
rect 12304 26715 12336 26747
rect 12376 26715 12408 26747
rect 12448 26715 12480 26747
rect 12520 26715 12552 26747
rect 12592 26715 12624 26747
rect 12664 26715 12696 26747
rect 12736 26715 12768 26747
rect 12808 26715 12840 26747
rect 12880 26715 12912 26747
rect 12952 26715 12984 26747
rect 13024 26715 13056 26747
rect 13096 26715 13128 26747
rect 13168 26715 13200 26747
rect 13240 26715 13272 26747
rect 13312 26715 13344 26747
rect 13384 26715 13416 26747
rect 13456 26715 13488 26747
rect 13528 26715 13560 26747
rect 13600 26715 13632 26747
rect 13672 26715 13704 26747
rect 13744 26715 13776 26747
rect 13816 26715 13848 26747
rect 13888 26715 13920 26747
rect 13960 26715 13992 26747
rect 14032 26715 14064 26747
rect 14104 26715 14136 26747
rect 14176 26715 14208 26747
rect 14248 26715 14280 26747
rect 14320 26715 14352 26747
rect 14392 26715 14424 26747
rect 14464 26715 14496 26747
rect 14536 26715 14568 26747
rect 14608 26715 14640 26747
rect 14680 26715 14712 26747
rect 14752 26715 14784 26747
rect 14824 26715 14856 26747
rect 14896 26715 14928 26747
rect 14968 26715 15000 26747
rect 15040 26715 15072 26747
rect 15112 26715 15144 26747
rect 15184 26715 15216 26747
rect 15256 26715 15288 26747
rect 15328 26715 15360 26747
rect 15400 26715 15432 26747
rect 15472 26715 15504 26747
rect 15544 26715 15576 26747
rect 15616 26715 15648 26747
rect 15688 26715 15720 26747
rect 15760 26715 15792 26747
rect 15832 26715 15864 26747
rect 15904 26715 15936 26747
rect 64 26643 96 26675
rect 136 26643 168 26675
rect 208 26643 240 26675
rect 280 26643 312 26675
rect 352 26643 384 26675
rect 424 26643 456 26675
rect 496 26643 528 26675
rect 568 26643 600 26675
rect 640 26643 672 26675
rect 712 26643 744 26675
rect 784 26643 816 26675
rect 856 26643 888 26675
rect 928 26643 960 26675
rect 1000 26643 1032 26675
rect 1072 26643 1104 26675
rect 1144 26643 1176 26675
rect 1216 26643 1248 26675
rect 1288 26643 1320 26675
rect 1360 26643 1392 26675
rect 1432 26643 1464 26675
rect 1504 26643 1536 26675
rect 1576 26643 1608 26675
rect 1648 26643 1680 26675
rect 1720 26643 1752 26675
rect 1792 26643 1824 26675
rect 1864 26643 1896 26675
rect 1936 26643 1968 26675
rect 2008 26643 2040 26675
rect 2080 26643 2112 26675
rect 2152 26643 2184 26675
rect 2224 26643 2256 26675
rect 2296 26643 2328 26675
rect 2368 26643 2400 26675
rect 2440 26643 2472 26675
rect 2512 26643 2544 26675
rect 2584 26643 2616 26675
rect 2656 26643 2688 26675
rect 2728 26643 2760 26675
rect 2800 26643 2832 26675
rect 2872 26643 2904 26675
rect 2944 26643 2976 26675
rect 3016 26643 3048 26675
rect 3088 26643 3120 26675
rect 3160 26643 3192 26675
rect 3232 26643 3264 26675
rect 3304 26643 3336 26675
rect 3376 26643 3408 26675
rect 3448 26643 3480 26675
rect 3520 26643 3552 26675
rect 3592 26643 3624 26675
rect 3664 26643 3696 26675
rect 3736 26643 3768 26675
rect 3808 26643 3840 26675
rect 3880 26643 3912 26675
rect 3952 26643 3984 26675
rect 4024 26643 4056 26675
rect 4096 26643 4128 26675
rect 4168 26643 4200 26675
rect 4240 26643 4272 26675
rect 4312 26643 4344 26675
rect 4384 26643 4416 26675
rect 4456 26643 4488 26675
rect 4528 26643 4560 26675
rect 4600 26643 4632 26675
rect 4672 26643 4704 26675
rect 4744 26643 4776 26675
rect 4816 26643 4848 26675
rect 4888 26643 4920 26675
rect 4960 26643 4992 26675
rect 5032 26643 5064 26675
rect 5104 26643 5136 26675
rect 5176 26643 5208 26675
rect 5248 26643 5280 26675
rect 5320 26643 5352 26675
rect 5392 26643 5424 26675
rect 5464 26643 5496 26675
rect 5536 26643 5568 26675
rect 5608 26643 5640 26675
rect 5680 26643 5712 26675
rect 5752 26643 5784 26675
rect 5824 26643 5856 26675
rect 5896 26643 5928 26675
rect 5968 26643 6000 26675
rect 6040 26643 6072 26675
rect 6112 26643 6144 26675
rect 6184 26643 6216 26675
rect 6256 26643 6288 26675
rect 6328 26643 6360 26675
rect 6400 26643 6432 26675
rect 6472 26643 6504 26675
rect 6544 26643 6576 26675
rect 6616 26643 6648 26675
rect 6688 26643 6720 26675
rect 6760 26643 6792 26675
rect 6832 26643 6864 26675
rect 6904 26643 6936 26675
rect 6976 26643 7008 26675
rect 7048 26643 7080 26675
rect 7120 26643 7152 26675
rect 7192 26643 7224 26675
rect 7264 26643 7296 26675
rect 7336 26643 7368 26675
rect 7408 26643 7440 26675
rect 7480 26643 7512 26675
rect 7552 26643 7584 26675
rect 7624 26643 7656 26675
rect 7696 26643 7728 26675
rect 7768 26643 7800 26675
rect 7840 26643 7872 26675
rect 7912 26643 7944 26675
rect 7984 26643 8016 26675
rect 8056 26643 8088 26675
rect 8128 26643 8160 26675
rect 8200 26643 8232 26675
rect 8272 26643 8304 26675
rect 8344 26643 8376 26675
rect 8416 26643 8448 26675
rect 8488 26643 8520 26675
rect 8560 26643 8592 26675
rect 8632 26643 8664 26675
rect 8704 26643 8736 26675
rect 8776 26643 8808 26675
rect 8848 26643 8880 26675
rect 8920 26643 8952 26675
rect 8992 26643 9024 26675
rect 9064 26643 9096 26675
rect 9136 26643 9168 26675
rect 9208 26643 9240 26675
rect 9280 26643 9312 26675
rect 9352 26643 9384 26675
rect 9424 26643 9456 26675
rect 9496 26643 9528 26675
rect 9568 26643 9600 26675
rect 9640 26643 9672 26675
rect 9712 26643 9744 26675
rect 9784 26643 9816 26675
rect 9856 26643 9888 26675
rect 9928 26643 9960 26675
rect 10000 26643 10032 26675
rect 10072 26643 10104 26675
rect 10144 26643 10176 26675
rect 10216 26643 10248 26675
rect 10288 26643 10320 26675
rect 10360 26643 10392 26675
rect 10432 26643 10464 26675
rect 10504 26643 10536 26675
rect 10576 26643 10608 26675
rect 10648 26643 10680 26675
rect 10720 26643 10752 26675
rect 10792 26643 10824 26675
rect 10864 26643 10896 26675
rect 10936 26643 10968 26675
rect 11008 26643 11040 26675
rect 11080 26643 11112 26675
rect 11152 26643 11184 26675
rect 11224 26643 11256 26675
rect 11296 26643 11328 26675
rect 11368 26643 11400 26675
rect 11440 26643 11472 26675
rect 11512 26643 11544 26675
rect 11584 26643 11616 26675
rect 11656 26643 11688 26675
rect 11728 26643 11760 26675
rect 11800 26643 11832 26675
rect 11872 26643 11904 26675
rect 11944 26643 11976 26675
rect 12016 26643 12048 26675
rect 12088 26643 12120 26675
rect 12160 26643 12192 26675
rect 12232 26643 12264 26675
rect 12304 26643 12336 26675
rect 12376 26643 12408 26675
rect 12448 26643 12480 26675
rect 12520 26643 12552 26675
rect 12592 26643 12624 26675
rect 12664 26643 12696 26675
rect 12736 26643 12768 26675
rect 12808 26643 12840 26675
rect 12880 26643 12912 26675
rect 12952 26643 12984 26675
rect 13024 26643 13056 26675
rect 13096 26643 13128 26675
rect 13168 26643 13200 26675
rect 13240 26643 13272 26675
rect 13312 26643 13344 26675
rect 13384 26643 13416 26675
rect 13456 26643 13488 26675
rect 13528 26643 13560 26675
rect 13600 26643 13632 26675
rect 13672 26643 13704 26675
rect 13744 26643 13776 26675
rect 13816 26643 13848 26675
rect 13888 26643 13920 26675
rect 13960 26643 13992 26675
rect 14032 26643 14064 26675
rect 14104 26643 14136 26675
rect 14176 26643 14208 26675
rect 14248 26643 14280 26675
rect 14320 26643 14352 26675
rect 14392 26643 14424 26675
rect 14464 26643 14496 26675
rect 14536 26643 14568 26675
rect 14608 26643 14640 26675
rect 14680 26643 14712 26675
rect 14752 26643 14784 26675
rect 14824 26643 14856 26675
rect 14896 26643 14928 26675
rect 14968 26643 15000 26675
rect 15040 26643 15072 26675
rect 15112 26643 15144 26675
rect 15184 26643 15216 26675
rect 15256 26643 15288 26675
rect 15328 26643 15360 26675
rect 15400 26643 15432 26675
rect 15472 26643 15504 26675
rect 15544 26643 15576 26675
rect 15616 26643 15648 26675
rect 15688 26643 15720 26675
rect 15760 26643 15792 26675
rect 15832 26643 15864 26675
rect 15904 26643 15936 26675
rect 64 26571 96 26603
rect 136 26571 168 26603
rect 208 26571 240 26603
rect 280 26571 312 26603
rect 352 26571 384 26603
rect 424 26571 456 26603
rect 496 26571 528 26603
rect 568 26571 600 26603
rect 640 26571 672 26603
rect 712 26571 744 26603
rect 784 26571 816 26603
rect 856 26571 888 26603
rect 928 26571 960 26603
rect 1000 26571 1032 26603
rect 1072 26571 1104 26603
rect 1144 26571 1176 26603
rect 1216 26571 1248 26603
rect 1288 26571 1320 26603
rect 1360 26571 1392 26603
rect 1432 26571 1464 26603
rect 1504 26571 1536 26603
rect 1576 26571 1608 26603
rect 1648 26571 1680 26603
rect 1720 26571 1752 26603
rect 1792 26571 1824 26603
rect 1864 26571 1896 26603
rect 1936 26571 1968 26603
rect 2008 26571 2040 26603
rect 2080 26571 2112 26603
rect 2152 26571 2184 26603
rect 2224 26571 2256 26603
rect 2296 26571 2328 26603
rect 2368 26571 2400 26603
rect 2440 26571 2472 26603
rect 2512 26571 2544 26603
rect 2584 26571 2616 26603
rect 2656 26571 2688 26603
rect 2728 26571 2760 26603
rect 2800 26571 2832 26603
rect 2872 26571 2904 26603
rect 2944 26571 2976 26603
rect 3016 26571 3048 26603
rect 3088 26571 3120 26603
rect 3160 26571 3192 26603
rect 3232 26571 3264 26603
rect 3304 26571 3336 26603
rect 3376 26571 3408 26603
rect 3448 26571 3480 26603
rect 3520 26571 3552 26603
rect 3592 26571 3624 26603
rect 3664 26571 3696 26603
rect 3736 26571 3768 26603
rect 3808 26571 3840 26603
rect 3880 26571 3912 26603
rect 3952 26571 3984 26603
rect 4024 26571 4056 26603
rect 4096 26571 4128 26603
rect 4168 26571 4200 26603
rect 4240 26571 4272 26603
rect 4312 26571 4344 26603
rect 4384 26571 4416 26603
rect 4456 26571 4488 26603
rect 4528 26571 4560 26603
rect 4600 26571 4632 26603
rect 4672 26571 4704 26603
rect 4744 26571 4776 26603
rect 4816 26571 4848 26603
rect 4888 26571 4920 26603
rect 4960 26571 4992 26603
rect 5032 26571 5064 26603
rect 5104 26571 5136 26603
rect 5176 26571 5208 26603
rect 5248 26571 5280 26603
rect 5320 26571 5352 26603
rect 5392 26571 5424 26603
rect 5464 26571 5496 26603
rect 5536 26571 5568 26603
rect 5608 26571 5640 26603
rect 5680 26571 5712 26603
rect 5752 26571 5784 26603
rect 5824 26571 5856 26603
rect 5896 26571 5928 26603
rect 5968 26571 6000 26603
rect 6040 26571 6072 26603
rect 6112 26571 6144 26603
rect 6184 26571 6216 26603
rect 6256 26571 6288 26603
rect 6328 26571 6360 26603
rect 6400 26571 6432 26603
rect 6472 26571 6504 26603
rect 6544 26571 6576 26603
rect 6616 26571 6648 26603
rect 6688 26571 6720 26603
rect 6760 26571 6792 26603
rect 6832 26571 6864 26603
rect 6904 26571 6936 26603
rect 6976 26571 7008 26603
rect 7048 26571 7080 26603
rect 7120 26571 7152 26603
rect 7192 26571 7224 26603
rect 7264 26571 7296 26603
rect 7336 26571 7368 26603
rect 7408 26571 7440 26603
rect 7480 26571 7512 26603
rect 7552 26571 7584 26603
rect 7624 26571 7656 26603
rect 7696 26571 7728 26603
rect 7768 26571 7800 26603
rect 7840 26571 7872 26603
rect 7912 26571 7944 26603
rect 7984 26571 8016 26603
rect 8056 26571 8088 26603
rect 8128 26571 8160 26603
rect 8200 26571 8232 26603
rect 8272 26571 8304 26603
rect 8344 26571 8376 26603
rect 8416 26571 8448 26603
rect 8488 26571 8520 26603
rect 8560 26571 8592 26603
rect 8632 26571 8664 26603
rect 8704 26571 8736 26603
rect 8776 26571 8808 26603
rect 8848 26571 8880 26603
rect 8920 26571 8952 26603
rect 8992 26571 9024 26603
rect 9064 26571 9096 26603
rect 9136 26571 9168 26603
rect 9208 26571 9240 26603
rect 9280 26571 9312 26603
rect 9352 26571 9384 26603
rect 9424 26571 9456 26603
rect 9496 26571 9528 26603
rect 9568 26571 9600 26603
rect 9640 26571 9672 26603
rect 9712 26571 9744 26603
rect 9784 26571 9816 26603
rect 9856 26571 9888 26603
rect 9928 26571 9960 26603
rect 10000 26571 10032 26603
rect 10072 26571 10104 26603
rect 10144 26571 10176 26603
rect 10216 26571 10248 26603
rect 10288 26571 10320 26603
rect 10360 26571 10392 26603
rect 10432 26571 10464 26603
rect 10504 26571 10536 26603
rect 10576 26571 10608 26603
rect 10648 26571 10680 26603
rect 10720 26571 10752 26603
rect 10792 26571 10824 26603
rect 10864 26571 10896 26603
rect 10936 26571 10968 26603
rect 11008 26571 11040 26603
rect 11080 26571 11112 26603
rect 11152 26571 11184 26603
rect 11224 26571 11256 26603
rect 11296 26571 11328 26603
rect 11368 26571 11400 26603
rect 11440 26571 11472 26603
rect 11512 26571 11544 26603
rect 11584 26571 11616 26603
rect 11656 26571 11688 26603
rect 11728 26571 11760 26603
rect 11800 26571 11832 26603
rect 11872 26571 11904 26603
rect 11944 26571 11976 26603
rect 12016 26571 12048 26603
rect 12088 26571 12120 26603
rect 12160 26571 12192 26603
rect 12232 26571 12264 26603
rect 12304 26571 12336 26603
rect 12376 26571 12408 26603
rect 12448 26571 12480 26603
rect 12520 26571 12552 26603
rect 12592 26571 12624 26603
rect 12664 26571 12696 26603
rect 12736 26571 12768 26603
rect 12808 26571 12840 26603
rect 12880 26571 12912 26603
rect 12952 26571 12984 26603
rect 13024 26571 13056 26603
rect 13096 26571 13128 26603
rect 13168 26571 13200 26603
rect 13240 26571 13272 26603
rect 13312 26571 13344 26603
rect 13384 26571 13416 26603
rect 13456 26571 13488 26603
rect 13528 26571 13560 26603
rect 13600 26571 13632 26603
rect 13672 26571 13704 26603
rect 13744 26571 13776 26603
rect 13816 26571 13848 26603
rect 13888 26571 13920 26603
rect 13960 26571 13992 26603
rect 14032 26571 14064 26603
rect 14104 26571 14136 26603
rect 14176 26571 14208 26603
rect 14248 26571 14280 26603
rect 14320 26571 14352 26603
rect 14392 26571 14424 26603
rect 14464 26571 14496 26603
rect 14536 26571 14568 26603
rect 14608 26571 14640 26603
rect 14680 26571 14712 26603
rect 14752 26571 14784 26603
rect 14824 26571 14856 26603
rect 14896 26571 14928 26603
rect 14968 26571 15000 26603
rect 15040 26571 15072 26603
rect 15112 26571 15144 26603
rect 15184 26571 15216 26603
rect 15256 26571 15288 26603
rect 15328 26571 15360 26603
rect 15400 26571 15432 26603
rect 15472 26571 15504 26603
rect 15544 26571 15576 26603
rect 15616 26571 15648 26603
rect 15688 26571 15720 26603
rect 15760 26571 15792 26603
rect 15832 26571 15864 26603
rect 15904 26571 15936 26603
rect 64 26499 96 26531
rect 136 26499 168 26531
rect 208 26499 240 26531
rect 280 26499 312 26531
rect 352 26499 384 26531
rect 424 26499 456 26531
rect 496 26499 528 26531
rect 568 26499 600 26531
rect 640 26499 672 26531
rect 712 26499 744 26531
rect 784 26499 816 26531
rect 856 26499 888 26531
rect 928 26499 960 26531
rect 1000 26499 1032 26531
rect 1072 26499 1104 26531
rect 1144 26499 1176 26531
rect 1216 26499 1248 26531
rect 1288 26499 1320 26531
rect 1360 26499 1392 26531
rect 1432 26499 1464 26531
rect 1504 26499 1536 26531
rect 1576 26499 1608 26531
rect 1648 26499 1680 26531
rect 1720 26499 1752 26531
rect 1792 26499 1824 26531
rect 1864 26499 1896 26531
rect 1936 26499 1968 26531
rect 2008 26499 2040 26531
rect 2080 26499 2112 26531
rect 2152 26499 2184 26531
rect 2224 26499 2256 26531
rect 2296 26499 2328 26531
rect 2368 26499 2400 26531
rect 2440 26499 2472 26531
rect 2512 26499 2544 26531
rect 2584 26499 2616 26531
rect 2656 26499 2688 26531
rect 2728 26499 2760 26531
rect 2800 26499 2832 26531
rect 2872 26499 2904 26531
rect 2944 26499 2976 26531
rect 3016 26499 3048 26531
rect 3088 26499 3120 26531
rect 3160 26499 3192 26531
rect 3232 26499 3264 26531
rect 3304 26499 3336 26531
rect 3376 26499 3408 26531
rect 3448 26499 3480 26531
rect 3520 26499 3552 26531
rect 3592 26499 3624 26531
rect 3664 26499 3696 26531
rect 3736 26499 3768 26531
rect 3808 26499 3840 26531
rect 3880 26499 3912 26531
rect 3952 26499 3984 26531
rect 4024 26499 4056 26531
rect 4096 26499 4128 26531
rect 4168 26499 4200 26531
rect 4240 26499 4272 26531
rect 4312 26499 4344 26531
rect 4384 26499 4416 26531
rect 4456 26499 4488 26531
rect 4528 26499 4560 26531
rect 4600 26499 4632 26531
rect 4672 26499 4704 26531
rect 4744 26499 4776 26531
rect 4816 26499 4848 26531
rect 4888 26499 4920 26531
rect 4960 26499 4992 26531
rect 5032 26499 5064 26531
rect 5104 26499 5136 26531
rect 5176 26499 5208 26531
rect 5248 26499 5280 26531
rect 5320 26499 5352 26531
rect 5392 26499 5424 26531
rect 5464 26499 5496 26531
rect 5536 26499 5568 26531
rect 5608 26499 5640 26531
rect 5680 26499 5712 26531
rect 5752 26499 5784 26531
rect 5824 26499 5856 26531
rect 5896 26499 5928 26531
rect 5968 26499 6000 26531
rect 6040 26499 6072 26531
rect 6112 26499 6144 26531
rect 6184 26499 6216 26531
rect 6256 26499 6288 26531
rect 6328 26499 6360 26531
rect 6400 26499 6432 26531
rect 6472 26499 6504 26531
rect 6544 26499 6576 26531
rect 6616 26499 6648 26531
rect 6688 26499 6720 26531
rect 6760 26499 6792 26531
rect 6832 26499 6864 26531
rect 6904 26499 6936 26531
rect 6976 26499 7008 26531
rect 7048 26499 7080 26531
rect 7120 26499 7152 26531
rect 7192 26499 7224 26531
rect 7264 26499 7296 26531
rect 7336 26499 7368 26531
rect 7408 26499 7440 26531
rect 7480 26499 7512 26531
rect 7552 26499 7584 26531
rect 7624 26499 7656 26531
rect 7696 26499 7728 26531
rect 7768 26499 7800 26531
rect 7840 26499 7872 26531
rect 7912 26499 7944 26531
rect 7984 26499 8016 26531
rect 8056 26499 8088 26531
rect 8128 26499 8160 26531
rect 8200 26499 8232 26531
rect 8272 26499 8304 26531
rect 8344 26499 8376 26531
rect 8416 26499 8448 26531
rect 8488 26499 8520 26531
rect 8560 26499 8592 26531
rect 8632 26499 8664 26531
rect 8704 26499 8736 26531
rect 8776 26499 8808 26531
rect 8848 26499 8880 26531
rect 8920 26499 8952 26531
rect 8992 26499 9024 26531
rect 9064 26499 9096 26531
rect 9136 26499 9168 26531
rect 9208 26499 9240 26531
rect 9280 26499 9312 26531
rect 9352 26499 9384 26531
rect 9424 26499 9456 26531
rect 9496 26499 9528 26531
rect 9568 26499 9600 26531
rect 9640 26499 9672 26531
rect 9712 26499 9744 26531
rect 9784 26499 9816 26531
rect 9856 26499 9888 26531
rect 9928 26499 9960 26531
rect 10000 26499 10032 26531
rect 10072 26499 10104 26531
rect 10144 26499 10176 26531
rect 10216 26499 10248 26531
rect 10288 26499 10320 26531
rect 10360 26499 10392 26531
rect 10432 26499 10464 26531
rect 10504 26499 10536 26531
rect 10576 26499 10608 26531
rect 10648 26499 10680 26531
rect 10720 26499 10752 26531
rect 10792 26499 10824 26531
rect 10864 26499 10896 26531
rect 10936 26499 10968 26531
rect 11008 26499 11040 26531
rect 11080 26499 11112 26531
rect 11152 26499 11184 26531
rect 11224 26499 11256 26531
rect 11296 26499 11328 26531
rect 11368 26499 11400 26531
rect 11440 26499 11472 26531
rect 11512 26499 11544 26531
rect 11584 26499 11616 26531
rect 11656 26499 11688 26531
rect 11728 26499 11760 26531
rect 11800 26499 11832 26531
rect 11872 26499 11904 26531
rect 11944 26499 11976 26531
rect 12016 26499 12048 26531
rect 12088 26499 12120 26531
rect 12160 26499 12192 26531
rect 12232 26499 12264 26531
rect 12304 26499 12336 26531
rect 12376 26499 12408 26531
rect 12448 26499 12480 26531
rect 12520 26499 12552 26531
rect 12592 26499 12624 26531
rect 12664 26499 12696 26531
rect 12736 26499 12768 26531
rect 12808 26499 12840 26531
rect 12880 26499 12912 26531
rect 12952 26499 12984 26531
rect 13024 26499 13056 26531
rect 13096 26499 13128 26531
rect 13168 26499 13200 26531
rect 13240 26499 13272 26531
rect 13312 26499 13344 26531
rect 13384 26499 13416 26531
rect 13456 26499 13488 26531
rect 13528 26499 13560 26531
rect 13600 26499 13632 26531
rect 13672 26499 13704 26531
rect 13744 26499 13776 26531
rect 13816 26499 13848 26531
rect 13888 26499 13920 26531
rect 13960 26499 13992 26531
rect 14032 26499 14064 26531
rect 14104 26499 14136 26531
rect 14176 26499 14208 26531
rect 14248 26499 14280 26531
rect 14320 26499 14352 26531
rect 14392 26499 14424 26531
rect 14464 26499 14496 26531
rect 14536 26499 14568 26531
rect 14608 26499 14640 26531
rect 14680 26499 14712 26531
rect 14752 26499 14784 26531
rect 14824 26499 14856 26531
rect 14896 26499 14928 26531
rect 14968 26499 15000 26531
rect 15040 26499 15072 26531
rect 15112 26499 15144 26531
rect 15184 26499 15216 26531
rect 15256 26499 15288 26531
rect 15328 26499 15360 26531
rect 15400 26499 15432 26531
rect 15472 26499 15504 26531
rect 15544 26499 15576 26531
rect 15616 26499 15648 26531
rect 15688 26499 15720 26531
rect 15760 26499 15792 26531
rect 15832 26499 15864 26531
rect 15904 26499 15936 26531
rect 64 26427 96 26459
rect 136 26427 168 26459
rect 208 26427 240 26459
rect 280 26427 312 26459
rect 352 26427 384 26459
rect 424 26427 456 26459
rect 496 26427 528 26459
rect 568 26427 600 26459
rect 640 26427 672 26459
rect 712 26427 744 26459
rect 784 26427 816 26459
rect 856 26427 888 26459
rect 928 26427 960 26459
rect 1000 26427 1032 26459
rect 1072 26427 1104 26459
rect 1144 26427 1176 26459
rect 1216 26427 1248 26459
rect 1288 26427 1320 26459
rect 1360 26427 1392 26459
rect 1432 26427 1464 26459
rect 1504 26427 1536 26459
rect 1576 26427 1608 26459
rect 1648 26427 1680 26459
rect 1720 26427 1752 26459
rect 1792 26427 1824 26459
rect 1864 26427 1896 26459
rect 1936 26427 1968 26459
rect 2008 26427 2040 26459
rect 2080 26427 2112 26459
rect 2152 26427 2184 26459
rect 2224 26427 2256 26459
rect 2296 26427 2328 26459
rect 2368 26427 2400 26459
rect 2440 26427 2472 26459
rect 2512 26427 2544 26459
rect 2584 26427 2616 26459
rect 2656 26427 2688 26459
rect 2728 26427 2760 26459
rect 2800 26427 2832 26459
rect 2872 26427 2904 26459
rect 2944 26427 2976 26459
rect 3016 26427 3048 26459
rect 3088 26427 3120 26459
rect 3160 26427 3192 26459
rect 3232 26427 3264 26459
rect 3304 26427 3336 26459
rect 3376 26427 3408 26459
rect 3448 26427 3480 26459
rect 3520 26427 3552 26459
rect 3592 26427 3624 26459
rect 3664 26427 3696 26459
rect 3736 26427 3768 26459
rect 3808 26427 3840 26459
rect 3880 26427 3912 26459
rect 3952 26427 3984 26459
rect 4024 26427 4056 26459
rect 4096 26427 4128 26459
rect 4168 26427 4200 26459
rect 4240 26427 4272 26459
rect 4312 26427 4344 26459
rect 4384 26427 4416 26459
rect 4456 26427 4488 26459
rect 4528 26427 4560 26459
rect 4600 26427 4632 26459
rect 4672 26427 4704 26459
rect 4744 26427 4776 26459
rect 4816 26427 4848 26459
rect 4888 26427 4920 26459
rect 4960 26427 4992 26459
rect 5032 26427 5064 26459
rect 5104 26427 5136 26459
rect 5176 26427 5208 26459
rect 5248 26427 5280 26459
rect 5320 26427 5352 26459
rect 5392 26427 5424 26459
rect 5464 26427 5496 26459
rect 5536 26427 5568 26459
rect 5608 26427 5640 26459
rect 5680 26427 5712 26459
rect 5752 26427 5784 26459
rect 5824 26427 5856 26459
rect 5896 26427 5928 26459
rect 5968 26427 6000 26459
rect 6040 26427 6072 26459
rect 6112 26427 6144 26459
rect 6184 26427 6216 26459
rect 6256 26427 6288 26459
rect 6328 26427 6360 26459
rect 6400 26427 6432 26459
rect 6472 26427 6504 26459
rect 6544 26427 6576 26459
rect 6616 26427 6648 26459
rect 6688 26427 6720 26459
rect 6760 26427 6792 26459
rect 6832 26427 6864 26459
rect 6904 26427 6936 26459
rect 6976 26427 7008 26459
rect 7048 26427 7080 26459
rect 7120 26427 7152 26459
rect 7192 26427 7224 26459
rect 7264 26427 7296 26459
rect 7336 26427 7368 26459
rect 7408 26427 7440 26459
rect 7480 26427 7512 26459
rect 7552 26427 7584 26459
rect 7624 26427 7656 26459
rect 7696 26427 7728 26459
rect 7768 26427 7800 26459
rect 7840 26427 7872 26459
rect 7912 26427 7944 26459
rect 7984 26427 8016 26459
rect 8056 26427 8088 26459
rect 8128 26427 8160 26459
rect 8200 26427 8232 26459
rect 8272 26427 8304 26459
rect 8344 26427 8376 26459
rect 8416 26427 8448 26459
rect 8488 26427 8520 26459
rect 8560 26427 8592 26459
rect 8632 26427 8664 26459
rect 8704 26427 8736 26459
rect 8776 26427 8808 26459
rect 8848 26427 8880 26459
rect 8920 26427 8952 26459
rect 8992 26427 9024 26459
rect 9064 26427 9096 26459
rect 9136 26427 9168 26459
rect 9208 26427 9240 26459
rect 9280 26427 9312 26459
rect 9352 26427 9384 26459
rect 9424 26427 9456 26459
rect 9496 26427 9528 26459
rect 9568 26427 9600 26459
rect 9640 26427 9672 26459
rect 9712 26427 9744 26459
rect 9784 26427 9816 26459
rect 9856 26427 9888 26459
rect 9928 26427 9960 26459
rect 10000 26427 10032 26459
rect 10072 26427 10104 26459
rect 10144 26427 10176 26459
rect 10216 26427 10248 26459
rect 10288 26427 10320 26459
rect 10360 26427 10392 26459
rect 10432 26427 10464 26459
rect 10504 26427 10536 26459
rect 10576 26427 10608 26459
rect 10648 26427 10680 26459
rect 10720 26427 10752 26459
rect 10792 26427 10824 26459
rect 10864 26427 10896 26459
rect 10936 26427 10968 26459
rect 11008 26427 11040 26459
rect 11080 26427 11112 26459
rect 11152 26427 11184 26459
rect 11224 26427 11256 26459
rect 11296 26427 11328 26459
rect 11368 26427 11400 26459
rect 11440 26427 11472 26459
rect 11512 26427 11544 26459
rect 11584 26427 11616 26459
rect 11656 26427 11688 26459
rect 11728 26427 11760 26459
rect 11800 26427 11832 26459
rect 11872 26427 11904 26459
rect 11944 26427 11976 26459
rect 12016 26427 12048 26459
rect 12088 26427 12120 26459
rect 12160 26427 12192 26459
rect 12232 26427 12264 26459
rect 12304 26427 12336 26459
rect 12376 26427 12408 26459
rect 12448 26427 12480 26459
rect 12520 26427 12552 26459
rect 12592 26427 12624 26459
rect 12664 26427 12696 26459
rect 12736 26427 12768 26459
rect 12808 26427 12840 26459
rect 12880 26427 12912 26459
rect 12952 26427 12984 26459
rect 13024 26427 13056 26459
rect 13096 26427 13128 26459
rect 13168 26427 13200 26459
rect 13240 26427 13272 26459
rect 13312 26427 13344 26459
rect 13384 26427 13416 26459
rect 13456 26427 13488 26459
rect 13528 26427 13560 26459
rect 13600 26427 13632 26459
rect 13672 26427 13704 26459
rect 13744 26427 13776 26459
rect 13816 26427 13848 26459
rect 13888 26427 13920 26459
rect 13960 26427 13992 26459
rect 14032 26427 14064 26459
rect 14104 26427 14136 26459
rect 14176 26427 14208 26459
rect 14248 26427 14280 26459
rect 14320 26427 14352 26459
rect 14392 26427 14424 26459
rect 14464 26427 14496 26459
rect 14536 26427 14568 26459
rect 14608 26427 14640 26459
rect 14680 26427 14712 26459
rect 14752 26427 14784 26459
rect 14824 26427 14856 26459
rect 14896 26427 14928 26459
rect 14968 26427 15000 26459
rect 15040 26427 15072 26459
rect 15112 26427 15144 26459
rect 15184 26427 15216 26459
rect 15256 26427 15288 26459
rect 15328 26427 15360 26459
rect 15400 26427 15432 26459
rect 15472 26427 15504 26459
rect 15544 26427 15576 26459
rect 15616 26427 15648 26459
rect 15688 26427 15720 26459
rect 15760 26427 15792 26459
rect 15832 26427 15864 26459
rect 15904 26427 15936 26459
rect 64 26355 96 26387
rect 136 26355 168 26387
rect 208 26355 240 26387
rect 280 26355 312 26387
rect 352 26355 384 26387
rect 424 26355 456 26387
rect 496 26355 528 26387
rect 568 26355 600 26387
rect 640 26355 672 26387
rect 712 26355 744 26387
rect 784 26355 816 26387
rect 856 26355 888 26387
rect 928 26355 960 26387
rect 1000 26355 1032 26387
rect 1072 26355 1104 26387
rect 1144 26355 1176 26387
rect 1216 26355 1248 26387
rect 1288 26355 1320 26387
rect 1360 26355 1392 26387
rect 1432 26355 1464 26387
rect 1504 26355 1536 26387
rect 1576 26355 1608 26387
rect 1648 26355 1680 26387
rect 1720 26355 1752 26387
rect 1792 26355 1824 26387
rect 1864 26355 1896 26387
rect 1936 26355 1968 26387
rect 2008 26355 2040 26387
rect 2080 26355 2112 26387
rect 2152 26355 2184 26387
rect 2224 26355 2256 26387
rect 2296 26355 2328 26387
rect 2368 26355 2400 26387
rect 2440 26355 2472 26387
rect 2512 26355 2544 26387
rect 2584 26355 2616 26387
rect 2656 26355 2688 26387
rect 2728 26355 2760 26387
rect 2800 26355 2832 26387
rect 2872 26355 2904 26387
rect 2944 26355 2976 26387
rect 3016 26355 3048 26387
rect 3088 26355 3120 26387
rect 3160 26355 3192 26387
rect 3232 26355 3264 26387
rect 3304 26355 3336 26387
rect 3376 26355 3408 26387
rect 3448 26355 3480 26387
rect 3520 26355 3552 26387
rect 3592 26355 3624 26387
rect 3664 26355 3696 26387
rect 3736 26355 3768 26387
rect 3808 26355 3840 26387
rect 3880 26355 3912 26387
rect 3952 26355 3984 26387
rect 4024 26355 4056 26387
rect 4096 26355 4128 26387
rect 4168 26355 4200 26387
rect 4240 26355 4272 26387
rect 4312 26355 4344 26387
rect 4384 26355 4416 26387
rect 4456 26355 4488 26387
rect 4528 26355 4560 26387
rect 4600 26355 4632 26387
rect 4672 26355 4704 26387
rect 4744 26355 4776 26387
rect 4816 26355 4848 26387
rect 4888 26355 4920 26387
rect 4960 26355 4992 26387
rect 5032 26355 5064 26387
rect 5104 26355 5136 26387
rect 5176 26355 5208 26387
rect 5248 26355 5280 26387
rect 5320 26355 5352 26387
rect 5392 26355 5424 26387
rect 5464 26355 5496 26387
rect 5536 26355 5568 26387
rect 5608 26355 5640 26387
rect 5680 26355 5712 26387
rect 5752 26355 5784 26387
rect 5824 26355 5856 26387
rect 5896 26355 5928 26387
rect 5968 26355 6000 26387
rect 6040 26355 6072 26387
rect 6112 26355 6144 26387
rect 6184 26355 6216 26387
rect 6256 26355 6288 26387
rect 6328 26355 6360 26387
rect 6400 26355 6432 26387
rect 6472 26355 6504 26387
rect 6544 26355 6576 26387
rect 6616 26355 6648 26387
rect 6688 26355 6720 26387
rect 6760 26355 6792 26387
rect 6832 26355 6864 26387
rect 6904 26355 6936 26387
rect 6976 26355 7008 26387
rect 7048 26355 7080 26387
rect 7120 26355 7152 26387
rect 7192 26355 7224 26387
rect 7264 26355 7296 26387
rect 7336 26355 7368 26387
rect 7408 26355 7440 26387
rect 7480 26355 7512 26387
rect 7552 26355 7584 26387
rect 7624 26355 7656 26387
rect 7696 26355 7728 26387
rect 7768 26355 7800 26387
rect 7840 26355 7872 26387
rect 7912 26355 7944 26387
rect 7984 26355 8016 26387
rect 8056 26355 8088 26387
rect 8128 26355 8160 26387
rect 8200 26355 8232 26387
rect 8272 26355 8304 26387
rect 8344 26355 8376 26387
rect 8416 26355 8448 26387
rect 8488 26355 8520 26387
rect 8560 26355 8592 26387
rect 8632 26355 8664 26387
rect 8704 26355 8736 26387
rect 8776 26355 8808 26387
rect 8848 26355 8880 26387
rect 8920 26355 8952 26387
rect 8992 26355 9024 26387
rect 9064 26355 9096 26387
rect 9136 26355 9168 26387
rect 9208 26355 9240 26387
rect 9280 26355 9312 26387
rect 9352 26355 9384 26387
rect 9424 26355 9456 26387
rect 9496 26355 9528 26387
rect 9568 26355 9600 26387
rect 9640 26355 9672 26387
rect 9712 26355 9744 26387
rect 9784 26355 9816 26387
rect 9856 26355 9888 26387
rect 9928 26355 9960 26387
rect 10000 26355 10032 26387
rect 10072 26355 10104 26387
rect 10144 26355 10176 26387
rect 10216 26355 10248 26387
rect 10288 26355 10320 26387
rect 10360 26355 10392 26387
rect 10432 26355 10464 26387
rect 10504 26355 10536 26387
rect 10576 26355 10608 26387
rect 10648 26355 10680 26387
rect 10720 26355 10752 26387
rect 10792 26355 10824 26387
rect 10864 26355 10896 26387
rect 10936 26355 10968 26387
rect 11008 26355 11040 26387
rect 11080 26355 11112 26387
rect 11152 26355 11184 26387
rect 11224 26355 11256 26387
rect 11296 26355 11328 26387
rect 11368 26355 11400 26387
rect 11440 26355 11472 26387
rect 11512 26355 11544 26387
rect 11584 26355 11616 26387
rect 11656 26355 11688 26387
rect 11728 26355 11760 26387
rect 11800 26355 11832 26387
rect 11872 26355 11904 26387
rect 11944 26355 11976 26387
rect 12016 26355 12048 26387
rect 12088 26355 12120 26387
rect 12160 26355 12192 26387
rect 12232 26355 12264 26387
rect 12304 26355 12336 26387
rect 12376 26355 12408 26387
rect 12448 26355 12480 26387
rect 12520 26355 12552 26387
rect 12592 26355 12624 26387
rect 12664 26355 12696 26387
rect 12736 26355 12768 26387
rect 12808 26355 12840 26387
rect 12880 26355 12912 26387
rect 12952 26355 12984 26387
rect 13024 26355 13056 26387
rect 13096 26355 13128 26387
rect 13168 26355 13200 26387
rect 13240 26355 13272 26387
rect 13312 26355 13344 26387
rect 13384 26355 13416 26387
rect 13456 26355 13488 26387
rect 13528 26355 13560 26387
rect 13600 26355 13632 26387
rect 13672 26355 13704 26387
rect 13744 26355 13776 26387
rect 13816 26355 13848 26387
rect 13888 26355 13920 26387
rect 13960 26355 13992 26387
rect 14032 26355 14064 26387
rect 14104 26355 14136 26387
rect 14176 26355 14208 26387
rect 14248 26355 14280 26387
rect 14320 26355 14352 26387
rect 14392 26355 14424 26387
rect 14464 26355 14496 26387
rect 14536 26355 14568 26387
rect 14608 26355 14640 26387
rect 14680 26355 14712 26387
rect 14752 26355 14784 26387
rect 14824 26355 14856 26387
rect 14896 26355 14928 26387
rect 14968 26355 15000 26387
rect 15040 26355 15072 26387
rect 15112 26355 15144 26387
rect 15184 26355 15216 26387
rect 15256 26355 15288 26387
rect 15328 26355 15360 26387
rect 15400 26355 15432 26387
rect 15472 26355 15504 26387
rect 15544 26355 15576 26387
rect 15616 26355 15648 26387
rect 15688 26355 15720 26387
rect 15760 26355 15792 26387
rect 15832 26355 15864 26387
rect 15904 26355 15936 26387
rect 64 26283 96 26315
rect 136 26283 168 26315
rect 208 26283 240 26315
rect 280 26283 312 26315
rect 352 26283 384 26315
rect 424 26283 456 26315
rect 496 26283 528 26315
rect 568 26283 600 26315
rect 640 26283 672 26315
rect 712 26283 744 26315
rect 784 26283 816 26315
rect 856 26283 888 26315
rect 928 26283 960 26315
rect 1000 26283 1032 26315
rect 1072 26283 1104 26315
rect 1144 26283 1176 26315
rect 1216 26283 1248 26315
rect 1288 26283 1320 26315
rect 1360 26283 1392 26315
rect 1432 26283 1464 26315
rect 1504 26283 1536 26315
rect 1576 26283 1608 26315
rect 1648 26283 1680 26315
rect 1720 26283 1752 26315
rect 1792 26283 1824 26315
rect 1864 26283 1896 26315
rect 1936 26283 1968 26315
rect 2008 26283 2040 26315
rect 2080 26283 2112 26315
rect 2152 26283 2184 26315
rect 2224 26283 2256 26315
rect 2296 26283 2328 26315
rect 2368 26283 2400 26315
rect 2440 26283 2472 26315
rect 2512 26283 2544 26315
rect 2584 26283 2616 26315
rect 2656 26283 2688 26315
rect 2728 26283 2760 26315
rect 2800 26283 2832 26315
rect 2872 26283 2904 26315
rect 2944 26283 2976 26315
rect 3016 26283 3048 26315
rect 3088 26283 3120 26315
rect 3160 26283 3192 26315
rect 3232 26283 3264 26315
rect 3304 26283 3336 26315
rect 3376 26283 3408 26315
rect 3448 26283 3480 26315
rect 3520 26283 3552 26315
rect 3592 26283 3624 26315
rect 3664 26283 3696 26315
rect 3736 26283 3768 26315
rect 3808 26283 3840 26315
rect 3880 26283 3912 26315
rect 3952 26283 3984 26315
rect 4024 26283 4056 26315
rect 4096 26283 4128 26315
rect 4168 26283 4200 26315
rect 4240 26283 4272 26315
rect 4312 26283 4344 26315
rect 4384 26283 4416 26315
rect 4456 26283 4488 26315
rect 4528 26283 4560 26315
rect 4600 26283 4632 26315
rect 4672 26283 4704 26315
rect 4744 26283 4776 26315
rect 4816 26283 4848 26315
rect 4888 26283 4920 26315
rect 4960 26283 4992 26315
rect 5032 26283 5064 26315
rect 5104 26283 5136 26315
rect 5176 26283 5208 26315
rect 5248 26283 5280 26315
rect 5320 26283 5352 26315
rect 5392 26283 5424 26315
rect 5464 26283 5496 26315
rect 5536 26283 5568 26315
rect 5608 26283 5640 26315
rect 5680 26283 5712 26315
rect 5752 26283 5784 26315
rect 5824 26283 5856 26315
rect 5896 26283 5928 26315
rect 5968 26283 6000 26315
rect 6040 26283 6072 26315
rect 6112 26283 6144 26315
rect 6184 26283 6216 26315
rect 6256 26283 6288 26315
rect 6328 26283 6360 26315
rect 6400 26283 6432 26315
rect 6472 26283 6504 26315
rect 6544 26283 6576 26315
rect 6616 26283 6648 26315
rect 6688 26283 6720 26315
rect 6760 26283 6792 26315
rect 6832 26283 6864 26315
rect 6904 26283 6936 26315
rect 6976 26283 7008 26315
rect 7048 26283 7080 26315
rect 7120 26283 7152 26315
rect 7192 26283 7224 26315
rect 7264 26283 7296 26315
rect 7336 26283 7368 26315
rect 7408 26283 7440 26315
rect 7480 26283 7512 26315
rect 7552 26283 7584 26315
rect 7624 26283 7656 26315
rect 7696 26283 7728 26315
rect 7768 26283 7800 26315
rect 7840 26283 7872 26315
rect 7912 26283 7944 26315
rect 7984 26283 8016 26315
rect 8056 26283 8088 26315
rect 8128 26283 8160 26315
rect 8200 26283 8232 26315
rect 8272 26283 8304 26315
rect 8344 26283 8376 26315
rect 8416 26283 8448 26315
rect 8488 26283 8520 26315
rect 8560 26283 8592 26315
rect 8632 26283 8664 26315
rect 8704 26283 8736 26315
rect 8776 26283 8808 26315
rect 8848 26283 8880 26315
rect 8920 26283 8952 26315
rect 8992 26283 9024 26315
rect 9064 26283 9096 26315
rect 9136 26283 9168 26315
rect 9208 26283 9240 26315
rect 9280 26283 9312 26315
rect 9352 26283 9384 26315
rect 9424 26283 9456 26315
rect 9496 26283 9528 26315
rect 9568 26283 9600 26315
rect 9640 26283 9672 26315
rect 9712 26283 9744 26315
rect 9784 26283 9816 26315
rect 9856 26283 9888 26315
rect 9928 26283 9960 26315
rect 10000 26283 10032 26315
rect 10072 26283 10104 26315
rect 10144 26283 10176 26315
rect 10216 26283 10248 26315
rect 10288 26283 10320 26315
rect 10360 26283 10392 26315
rect 10432 26283 10464 26315
rect 10504 26283 10536 26315
rect 10576 26283 10608 26315
rect 10648 26283 10680 26315
rect 10720 26283 10752 26315
rect 10792 26283 10824 26315
rect 10864 26283 10896 26315
rect 10936 26283 10968 26315
rect 11008 26283 11040 26315
rect 11080 26283 11112 26315
rect 11152 26283 11184 26315
rect 11224 26283 11256 26315
rect 11296 26283 11328 26315
rect 11368 26283 11400 26315
rect 11440 26283 11472 26315
rect 11512 26283 11544 26315
rect 11584 26283 11616 26315
rect 11656 26283 11688 26315
rect 11728 26283 11760 26315
rect 11800 26283 11832 26315
rect 11872 26283 11904 26315
rect 11944 26283 11976 26315
rect 12016 26283 12048 26315
rect 12088 26283 12120 26315
rect 12160 26283 12192 26315
rect 12232 26283 12264 26315
rect 12304 26283 12336 26315
rect 12376 26283 12408 26315
rect 12448 26283 12480 26315
rect 12520 26283 12552 26315
rect 12592 26283 12624 26315
rect 12664 26283 12696 26315
rect 12736 26283 12768 26315
rect 12808 26283 12840 26315
rect 12880 26283 12912 26315
rect 12952 26283 12984 26315
rect 13024 26283 13056 26315
rect 13096 26283 13128 26315
rect 13168 26283 13200 26315
rect 13240 26283 13272 26315
rect 13312 26283 13344 26315
rect 13384 26283 13416 26315
rect 13456 26283 13488 26315
rect 13528 26283 13560 26315
rect 13600 26283 13632 26315
rect 13672 26283 13704 26315
rect 13744 26283 13776 26315
rect 13816 26283 13848 26315
rect 13888 26283 13920 26315
rect 13960 26283 13992 26315
rect 14032 26283 14064 26315
rect 14104 26283 14136 26315
rect 14176 26283 14208 26315
rect 14248 26283 14280 26315
rect 14320 26283 14352 26315
rect 14392 26283 14424 26315
rect 14464 26283 14496 26315
rect 14536 26283 14568 26315
rect 14608 26283 14640 26315
rect 14680 26283 14712 26315
rect 14752 26283 14784 26315
rect 14824 26283 14856 26315
rect 14896 26283 14928 26315
rect 14968 26283 15000 26315
rect 15040 26283 15072 26315
rect 15112 26283 15144 26315
rect 15184 26283 15216 26315
rect 15256 26283 15288 26315
rect 15328 26283 15360 26315
rect 15400 26283 15432 26315
rect 15472 26283 15504 26315
rect 15544 26283 15576 26315
rect 15616 26283 15648 26315
rect 15688 26283 15720 26315
rect 15760 26283 15792 26315
rect 15832 26283 15864 26315
rect 15904 26283 15936 26315
rect 64 26211 96 26243
rect 136 26211 168 26243
rect 208 26211 240 26243
rect 280 26211 312 26243
rect 352 26211 384 26243
rect 424 26211 456 26243
rect 496 26211 528 26243
rect 568 26211 600 26243
rect 640 26211 672 26243
rect 712 26211 744 26243
rect 784 26211 816 26243
rect 856 26211 888 26243
rect 928 26211 960 26243
rect 1000 26211 1032 26243
rect 1072 26211 1104 26243
rect 1144 26211 1176 26243
rect 1216 26211 1248 26243
rect 1288 26211 1320 26243
rect 1360 26211 1392 26243
rect 1432 26211 1464 26243
rect 1504 26211 1536 26243
rect 1576 26211 1608 26243
rect 1648 26211 1680 26243
rect 1720 26211 1752 26243
rect 1792 26211 1824 26243
rect 1864 26211 1896 26243
rect 1936 26211 1968 26243
rect 2008 26211 2040 26243
rect 2080 26211 2112 26243
rect 2152 26211 2184 26243
rect 2224 26211 2256 26243
rect 2296 26211 2328 26243
rect 2368 26211 2400 26243
rect 2440 26211 2472 26243
rect 2512 26211 2544 26243
rect 2584 26211 2616 26243
rect 2656 26211 2688 26243
rect 2728 26211 2760 26243
rect 2800 26211 2832 26243
rect 2872 26211 2904 26243
rect 2944 26211 2976 26243
rect 3016 26211 3048 26243
rect 3088 26211 3120 26243
rect 3160 26211 3192 26243
rect 3232 26211 3264 26243
rect 3304 26211 3336 26243
rect 3376 26211 3408 26243
rect 3448 26211 3480 26243
rect 3520 26211 3552 26243
rect 3592 26211 3624 26243
rect 3664 26211 3696 26243
rect 3736 26211 3768 26243
rect 3808 26211 3840 26243
rect 3880 26211 3912 26243
rect 3952 26211 3984 26243
rect 4024 26211 4056 26243
rect 4096 26211 4128 26243
rect 4168 26211 4200 26243
rect 4240 26211 4272 26243
rect 4312 26211 4344 26243
rect 4384 26211 4416 26243
rect 4456 26211 4488 26243
rect 4528 26211 4560 26243
rect 4600 26211 4632 26243
rect 4672 26211 4704 26243
rect 4744 26211 4776 26243
rect 4816 26211 4848 26243
rect 4888 26211 4920 26243
rect 4960 26211 4992 26243
rect 5032 26211 5064 26243
rect 5104 26211 5136 26243
rect 5176 26211 5208 26243
rect 5248 26211 5280 26243
rect 5320 26211 5352 26243
rect 5392 26211 5424 26243
rect 5464 26211 5496 26243
rect 5536 26211 5568 26243
rect 5608 26211 5640 26243
rect 5680 26211 5712 26243
rect 5752 26211 5784 26243
rect 5824 26211 5856 26243
rect 5896 26211 5928 26243
rect 5968 26211 6000 26243
rect 6040 26211 6072 26243
rect 6112 26211 6144 26243
rect 6184 26211 6216 26243
rect 6256 26211 6288 26243
rect 6328 26211 6360 26243
rect 6400 26211 6432 26243
rect 6472 26211 6504 26243
rect 6544 26211 6576 26243
rect 6616 26211 6648 26243
rect 6688 26211 6720 26243
rect 6760 26211 6792 26243
rect 6832 26211 6864 26243
rect 6904 26211 6936 26243
rect 6976 26211 7008 26243
rect 7048 26211 7080 26243
rect 7120 26211 7152 26243
rect 7192 26211 7224 26243
rect 7264 26211 7296 26243
rect 7336 26211 7368 26243
rect 7408 26211 7440 26243
rect 7480 26211 7512 26243
rect 7552 26211 7584 26243
rect 7624 26211 7656 26243
rect 7696 26211 7728 26243
rect 7768 26211 7800 26243
rect 7840 26211 7872 26243
rect 7912 26211 7944 26243
rect 7984 26211 8016 26243
rect 8056 26211 8088 26243
rect 8128 26211 8160 26243
rect 8200 26211 8232 26243
rect 8272 26211 8304 26243
rect 8344 26211 8376 26243
rect 8416 26211 8448 26243
rect 8488 26211 8520 26243
rect 8560 26211 8592 26243
rect 8632 26211 8664 26243
rect 8704 26211 8736 26243
rect 8776 26211 8808 26243
rect 8848 26211 8880 26243
rect 8920 26211 8952 26243
rect 8992 26211 9024 26243
rect 9064 26211 9096 26243
rect 9136 26211 9168 26243
rect 9208 26211 9240 26243
rect 9280 26211 9312 26243
rect 9352 26211 9384 26243
rect 9424 26211 9456 26243
rect 9496 26211 9528 26243
rect 9568 26211 9600 26243
rect 9640 26211 9672 26243
rect 9712 26211 9744 26243
rect 9784 26211 9816 26243
rect 9856 26211 9888 26243
rect 9928 26211 9960 26243
rect 10000 26211 10032 26243
rect 10072 26211 10104 26243
rect 10144 26211 10176 26243
rect 10216 26211 10248 26243
rect 10288 26211 10320 26243
rect 10360 26211 10392 26243
rect 10432 26211 10464 26243
rect 10504 26211 10536 26243
rect 10576 26211 10608 26243
rect 10648 26211 10680 26243
rect 10720 26211 10752 26243
rect 10792 26211 10824 26243
rect 10864 26211 10896 26243
rect 10936 26211 10968 26243
rect 11008 26211 11040 26243
rect 11080 26211 11112 26243
rect 11152 26211 11184 26243
rect 11224 26211 11256 26243
rect 11296 26211 11328 26243
rect 11368 26211 11400 26243
rect 11440 26211 11472 26243
rect 11512 26211 11544 26243
rect 11584 26211 11616 26243
rect 11656 26211 11688 26243
rect 11728 26211 11760 26243
rect 11800 26211 11832 26243
rect 11872 26211 11904 26243
rect 11944 26211 11976 26243
rect 12016 26211 12048 26243
rect 12088 26211 12120 26243
rect 12160 26211 12192 26243
rect 12232 26211 12264 26243
rect 12304 26211 12336 26243
rect 12376 26211 12408 26243
rect 12448 26211 12480 26243
rect 12520 26211 12552 26243
rect 12592 26211 12624 26243
rect 12664 26211 12696 26243
rect 12736 26211 12768 26243
rect 12808 26211 12840 26243
rect 12880 26211 12912 26243
rect 12952 26211 12984 26243
rect 13024 26211 13056 26243
rect 13096 26211 13128 26243
rect 13168 26211 13200 26243
rect 13240 26211 13272 26243
rect 13312 26211 13344 26243
rect 13384 26211 13416 26243
rect 13456 26211 13488 26243
rect 13528 26211 13560 26243
rect 13600 26211 13632 26243
rect 13672 26211 13704 26243
rect 13744 26211 13776 26243
rect 13816 26211 13848 26243
rect 13888 26211 13920 26243
rect 13960 26211 13992 26243
rect 14032 26211 14064 26243
rect 14104 26211 14136 26243
rect 14176 26211 14208 26243
rect 14248 26211 14280 26243
rect 14320 26211 14352 26243
rect 14392 26211 14424 26243
rect 14464 26211 14496 26243
rect 14536 26211 14568 26243
rect 14608 26211 14640 26243
rect 14680 26211 14712 26243
rect 14752 26211 14784 26243
rect 14824 26211 14856 26243
rect 14896 26211 14928 26243
rect 14968 26211 15000 26243
rect 15040 26211 15072 26243
rect 15112 26211 15144 26243
rect 15184 26211 15216 26243
rect 15256 26211 15288 26243
rect 15328 26211 15360 26243
rect 15400 26211 15432 26243
rect 15472 26211 15504 26243
rect 15544 26211 15576 26243
rect 15616 26211 15648 26243
rect 15688 26211 15720 26243
rect 15760 26211 15792 26243
rect 15832 26211 15864 26243
rect 15904 26211 15936 26243
rect 64 26139 96 26171
rect 136 26139 168 26171
rect 208 26139 240 26171
rect 280 26139 312 26171
rect 352 26139 384 26171
rect 424 26139 456 26171
rect 496 26139 528 26171
rect 568 26139 600 26171
rect 640 26139 672 26171
rect 712 26139 744 26171
rect 784 26139 816 26171
rect 856 26139 888 26171
rect 928 26139 960 26171
rect 1000 26139 1032 26171
rect 1072 26139 1104 26171
rect 1144 26139 1176 26171
rect 1216 26139 1248 26171
rect 1288 26139 1320 26171
rect 1360 26139 1392 26171
rect 1432 26139 1464 26171
rect 1504 26139 1536 26171
rect 1576 26139 1608 26171
rect 1648 26139 1680 26171
rect 1720 26139 1752 26171
rect 1792 26139 1824 26171
rect 1864 26139 1896 26171
rect 1936 26139 1968 26171
rect 2008 26139 2040 26171
rect 2080 26139 2112 26171
rect 2152 26139 2184 26171
rect 2224 26139 2256 26171
rect 2296 26139 2328 26171
rect 2368 26139 2400 26171
rect 2440 26139 2472 26171
rect 2512 26139 2544 26171
rect 2584 26139 2616 26171
rect 2656 26139 2688 26171
rect 2728 26139 2760 26171
rect 2800 26139 2832 26171
rect 2872 26139 2904 26171
rect 2944 26139 2976 26171
rect 3016 26139 3048 26171
rect 3088 26139 3120 26171
rect 3160 26139 3192 26171
rect 3232 26139 3264 26171
rect 3304 26139 3336 26171
rect 3376 26139 3408 26171
rect 3448 26139 3480 26171
rect 3520 26139 3552 26171
rect 3592 26139 3624 26171
rect 3664 26139 3696 26171
rect 3736 26139 3768 26171
rect 3808 26139 3840 26171
rect 3880 26139 3912 26171
rect 3952 26139 3984 26171
rect 4024 26139 4056 26171
rect 4096 26139 4128 26171
rect 4168 26139 4200 26171
rect 4240 26139 4272 26171
rect 4312 26139 4344 26171
rect 4384 26139 4416 26171
rect 4456 26139 4488 26171
rect 4528 26139 4560 26171
rect 4600 26139 4632 26171
rect 4672 26139 4704 26171
rect 4744 26139 4776 26171
rect 4816 26139 4848 26171
rect 4888 26139 4920 26171
rect 4960 26139 4992 26171
rect 5032 26139 5064 26171
rect 5104 26139 5136 26171
rect 5176 26139 5208 26171
rect 5248 26139 5280 26171
rect 5320 26139 5352 26171
rect 5392 26139 5424 26171
rect 5464 26139 5496 26171
rect 5536 26139 5568 26171
rect 5608 26139 5640 26171
rect 5680 26139 5712 26171
rect 5752 26139 5784 26171
rect 5824 26139 5856 26171
rect 5896 26139 5928 26171
rect 5968 26139 6000 26171
rect 6040 26139 6072 26171
rect 6112 26139 6144 26171
rect 6184 26139 6216 26171
rect 6256 26139 6288 26171
rect 6328 26139 6360 26171
rect 6400 26139 6432 26171
rect 6472 26139 6504 26171
rect 6544 26139 6576 26171
rect 6616 26139 6648 26171
rect 6688 26139 6720 26171
rect 6760 26139 6792 26171
rect 6832 26139 6864 26171
rect 6904 26139 6936 26171
rect 6976 26139 7008 26171
rect 7048 26139 7080 26171
rect 7120 26139 7152 26171
rect 7192 26139 7224 26171
rect 7264 26139 7296 26171
rect 7336 26139 7368 26171
rect 7408 26139 7440 26171
rect 7480 26139 7512 26171
rect 7552 26139 7584 26171
rect 7624 26139 7656 26171
rect 7696 26139 7728 26171
rect 7768 26139 7800 26171
rect 7840 26139 7872 26171
rect 7912 26139 7944 26171
rect 7984 26139 8016 26171
rect 8056 26139 8088 26171
rect 8128 26139 8160 26171
rect 8200 26139 8232 26171
rect 8272 26139 8304 26171
rect 8344 26139 8376 26171
rect 8416 26139 8448 26171
rect 8488 26139 8520 26171
rect 8560 26139 8592 26171
rect 8632 26139 8664 26171
rect 8704 26139 8736 26171
rect 8776 26139 8808 26171
rect 8848 26139 8880 26171
rect 8920 26139 8952 26171
rect 8992 26139 9024 26171
rect 9064 26139 9096 26171
rect 9136 26139 9168 26171
rect 9208 26139 9240 26171
rect 9280 26139 9312 26171
rect 9352 26139 9384 26171
rect 9424 26139 9456 26171
rect 9496 26139 9528 26171
rect 9568 26139 9600 26171
rect 9640 26139 9672 26171
rect 9712 26139 9744 26171
rect 9784 26139 9816 26171
rect 9856 26139 9888 26171
rect 9928 26139 9960 26171
rect 10000 26139 10032 26171
rect 10072 26139 10104 26171
rect 10144 26139 10176 26171
rect 10216 26139 10248 26171
rect 10288 26139 10320 26171
rect 10360 26139 10392 26171
rect 10432 26139 10464 26171
rect 10504 26139 10536 26171
rect 10576 26139 10608 26171
rect 10648 26139 10680 26171
rect 10720 26139 10752 26171
rect 10792 26139 10824 26171
rect 10864 26139 10896 26171
rect 10936 26139 10968 26171
rect 11008 26139 11040 26171
rect 11080 26139 11112 26171
rect 11152 26139 11184 26171
rect 11224 26139 11256 26171
rect 11296 26139 11328 26171
rect 11368 26139 11400 26171
rect 11440 26139 11472 26171
rect 11512 26139 11544 26171
rect 11584 26139 11616 26171
rect 11656 26139 11688 26171
rect 11728 26139 11760 26171
rect 11800 26139 11832 26171
rect 11872 26139 11904 26171
rect 11944 26139 11976 26171
rect 12016 26139 12048 26171
rect 12088 26139 12120 26171
rect 12160 26139 12192 26171
rect 12232 26139 12264 26171
rect 12304 26139 12336 26171
rect 12376 26139 12408 26171
rect 12448 26139 12480 26171
rect 12520 26139 12552 26171
rect 12592 26139 12624 26171
rect 12664 26139 12696 26171
rect 12736 26139 12768 26171
rect 12808 26139 12840 26171
rect 12880 26139 12912 26171
rect 12952 26139 12984 26171
rect 13024 26139 13056 26171
rect 13096 26139 13128 26171
rect 13168 26139 13200 26171
rect 13240 26139 13272 26171
rect 13312 26139 13344 26171
rect 13384 26139 13416 26171
rect 13456 26139 13488 26171
rect 13528 26139 13560 26171
rect 13600 26139 13632 26171
rect 13672 26139 13704 26171
rect 13744 26139 13776 26171
rect 13816 26139 13848 26171
rect 13888 26139 13920 26171
rect 13960 26139 13992 26171
rect 14032 26139 14064 26171
rect 14104 26139 14136 26171
rect 14176 26139 14208 26171
rect 14248 26139 14280 26171
rect 14320 26139 14352 26171
rect 14392 26139 14424 26171
rect 14464 26139 14496 26171
rect 14536 26139 14568 26171
rect 14608 26139 14640 26171
rect 14680 26139 14712 26171
rect 14752 26139 14784 26171
rect 14824 26139 14856 26171
rect 14896 26139 14928 26171
rect 14968 26139 15000 26171
rect 15040 26139 15072 26171
rect 15112 26139 15144 26171
rect 15184 26139 15216 26171
rect 15256 26139 15288 26171
rect 15328 26139 15360 26171
rect 15400 26139 15432 26171
rect 15472 26139 15504 26171
rect 15544 26139 15576 26171
rect 15616 26139 15648 26171
rect 15688 26139 15720 26171
rect 15760 26139 15792 26171
rect 15832 26139 15864 26171
rect 15904 26139 15936 26171
rect 64 26067 96 26099
rect 136 26067 168 26099
rect 208 26067 240 26099
rect 280 26067 312 26099
rect 352 26067 384 26099
rect 424 26067 456 26099
rect 496 26067 528 26099
rect 568 26067 600 26099
rect 640 26067 672 26099
rect 712 26067 744 26099
rect 784 26067 816 26099
rect 856 26067 888 26099
rect 928 26067 960 26099
rect 1000 26067 1032 26099
rect 1072 26067 1104 26099
rect 1144 26067 1176 26099
rect 1216 26067 1248 26099
rect 1288 26067 1320 26099
rect 1360 26067 1392 26099
rect 1432 26067 1464 26099
rect 1504 26067 1536 26099
rect 1576 26067 1608 26099
rect 1648 26067 1680 26099
rect 1720 26067 1752 26099
rect 1792 26067 1824 26099
rect 1864 26067 1896 26099
rect 1936 26067 1968 26099
rect 2008 26067 2040 26099
rect 2080 26067 2112 26099
rect 2152 26067 2184 26099
rect 2224 26067 2256 26099
rect 2296 26067 2328 26099
rect 2368 26067 2400 26099
rect 2440 26067 2472 26099
rect 2512 26067 2544 26099
rect 2584 26067 2616 26099
rect 2656 26067 2688 26099
rect 2728 26067 2760 26099
rect 2800 26067 2832 26099
rect 2872 26067 2904 26099
rect 2944 26067 2976 26099
rect 3016 26067 3048 26099
rect 3088 26067 3120 26099
rect 3160 26067 3192 26099
rect 3232 26067 3264 26099
rect 3304 26067 3336 26099
rect 3376 26067 3408 26099
rect 3448 26067 3480 26099
rect 3520 26067 3552 26099
rect 3592 26067 3624 26099
rect 3664 26067 3696 26099
rect 3736 26067 3768 26099
rect 3808 26067 3840 26099
rect 3880 26067 3912 26099
rect 3952 26067 3984 26099
rect 4024 26067 4056 26099
rect 4096 26067 4128 26099
rect 4168 26067 4200 26099
rect 4240 26067 4272 26099
rect 4312 26067 4344 26099
rect 4384 26067 4416 26099
rect 4456 26067 4488 26099
rect 4528 26067 4560 26099
rect 4600 26067 4632 26099
rect 4672 26067 4704 26099
rect 4744 26067 4776 26099
rect 4816 26067 4848 26099
rect 4888 26067 4920 26099
rect 4960 26067 4992 26099
rect 5032 26067 5064 26099
rect 5104 26067 5136 26099
rect 5176 26067 5208 26099
rect 5248 26067 5280 26099
rect 5320 26067 5352 26099
rect 5392 26067 5424 26099
rect 5464 26067 5496 26099
rect 5536 26067 5568 26099
rect 5608 26067 5640 26099
rect 5680 26067 5712 26099
rect 5752 26067 5784 26099
rect 5824 26067 5856 26099
rect 5896 26067 5928 26099
rect 5968 26067 6000 26099
rect 6040 26067 6072 26099
rect 6112 26067 6144 26099
rect 6184 26067 6216 26099
rect 6256 26067 6288 26099
rect 6328 26067 6360 26099
rect 6400 26067 6432 26099
rect 6472 26067 6504 26099
rect 6544 26067 6576 26099
rect 6616 26067 6648 26099
rect 6688 26067 6720 26099
rect 6760 26067 6792 26099
rect 6832 26067 6864 26099
rect 6904 26067 6936 26099
rect 6976 26067 7008 26099
rect 7048 26067 7080 26099
rect 7120 26067 7152 26099
rect 7192 26067 7224 26099
rect 7264 26067 7296 26099
rect 7336 26067 7368 26099
rect 7408 26067 7440 26099
rect 7480 26067 7512 26099
rect 7552 26067 7584 26099
rect 7624 26067 7656 26099
rect 7696 26067 7728 26099
rect 7768 26067 7800 26099
rect 7840 26067 7872 26099
rect 7912 26067 7944 26099
rect 7984 26067 8016 26099
rect 8056 26067 8088 26099
rect 8128 26067 8160 26099
rect 8200 26067 8232 26099
rect 8272 26067 8304 26099
rect 8344 26067 8376 26099
rect 8416 26067 8448 26099
rect 8488 26067 8520 26099
rect 8560 26067 8592 26099
rect 8632 26067 8664 26099
rect 8704 26067 8736 26099
rect 8776 26067 8808 26099
rect 8848 26067 8880 26099
rect 8920 26067 8952 26099
rect 8992 26067 9024 26099
rect 9064 26067 9096 26099
rect 9136 26067 9168 26099
rect 9208 26067 9240 26099
rect 9280 26067 9312 26099
rect 9352 26067 9384 26099
rect 9424 26067 9456 26099
rect 9496 26067 9528 26099
rect 9568 26067 9600 26099
rect 9640 26067 9672 26099
rect 9712 26067 9744 26099
rect 9784 26067 9816 26099
rect 9856 26067 9888 26099
rect 9928 26067 9960 26099
rect 10000 26067 10032 26099
rect 10072 26067 10104 26099
rect 10144 26067 10176 26099
rect 10216 26067 10248 26099
rect 10288 26067 10320 26099
rect 10360 26067 10392 26099
rect 10432 26067 10464 26099
rect 10504 26067 10536 26099
rect 10576 26067 10608 26099
rect 10648 26067 10680 26099
rect 10720 26067 10752 26099
rect 10792 26067 10824 26099
rect 10864 26067 10896 26099
rect 10936 26067 10968 26099
rect 11008 26067 11040 26099
rect 11080 26067 11112 26099
rect 11152 26067 11184 26099
rect 11224 26067 11256 26099
rect 11296 26067 11328 26099
rect 11368 26067 11400 26099
rect 11440 26067 11472 26099
rect 11512 26067 11544 26099
rect 11584 26067 11616 26099
rect 11656 26067 11688 26099
rect 11728 26067 11760 26099
rect 11800 26067 11832 26099
rect 11872 26067 11904 26099
rect 11944 26067 11976 26099
rect 12016 26067 12048 26099
rect 12088 26067 12120 26099
rect 12160 26067 12192 26099
rect 12232 26067 12264 26099
rect 12304 26067 12336 26099
rect 12376 26067 12408 26099
rect 12448 26067 12480 26099
rect 12520 26067 12552 26099
rect 12592 26067 12624 26099
rect 12664 26067 12696 26099
rect 12736 26067 12768 26099
rect 12808 26067 12840 26099
rect 12880 26067 12912 26099
rect 12952 26067 12984 26099
rect 13024 26067 13056 26099
rect 13096 26067 13128 26099
rect 13168 26067 13200 26099
rect 13240 26067 13272 26099
rect 13312 26067 13344 26099
rect 13384 26067 13416 26099
rect 13456 26067 13488 26099
rect 13528 26067 13560 26099
rect 13600 26067 13632 26099
rect 13672 26067 13704 26099
rect 13744 26067 13776 26099
rect 13816 26067 13848 26099
rect 13888 26067 13920 26099
rect 13960 26067 13992 26099
rect 14032 26067 14064 26099
rect 14104 26067 14136 26099
rect 14176 26067 14208 26099
rect 14248 26067 14280 26099
rect 14320 26067 14352 26099
rect 14392 26067 14424 26099
rect 14464 26067 14496 26099
rect 14536 26067 14568 26099
rect 14608 26067 14640 26099
rect 14680 26067 14712 26099
rect 14752 26067 14784 26099
rect 14824 26067 14856 26099
rect 14896 26067 14928 26099
rect 14968 26067 15000 26099
rect 15040 26067 15072 26099
rect 15112 26067 15144 26099
rect 15184 26067 15216 26099
rect 15256 26067 15288 26099
rect 15328 26067 15360 26099
rect 15400 26067 15432 26099
rect 15472 26067 15504 26099
rect 15544 26067 15576 26099
rect 15616 26067 15648 26099
rect 15688 26067 15720 26099
rect 15760 26067 15792 26099
rect 15832 26067 15864 26099
rect 15904 26067 15936 26099
rect 64 25995 96 26027
rect 136 25995 168 26027
rect 208 25995 240 26027
rect 280 25995 312 26027
rect 352 25995 384 26027
rect 424 25995 456 26027
rect 496 25995 528 26027
rect 568 25995 600 26027
rect 640 25995 672 26027
rect 712 25995 744 26027
rect 784 25995 816 26027
rect 856 25995 888 26027
rect 928 25995 960 26027
rect 1000 25995 1032 26027
rect 1072 25995 1104 26027
rect 1144 25995 1176 26027
rect 1216 25995 1248 26027
rect 1288 25995 1320 26027
rect 1360 25995 1392 26027
rect 1432 25995 1464 26027
rect 1504 25995 1536 26027
rect 1576 25995 1608 26027
rect 1648 25995 1680 26027
rect 1720 25995 1752 26027
rect 1792 25995 1824 26027
rect 1864 25995 1896 26027
rect 1936 25995 1968 26027
rect 2008 25995 2040 26027
rect 2080 25995 2112 26027
rect 2152 25995 2184 26027
rect 2224 25995 2256 26027
rect 2296 25995 2328 26027
rect 2368 25995 2400 26027
rect 2440 25995 2472 26027
rect 2512 25995 2544 26027
rect 2584 25995 2616 26027
rect 2656 25995 2688 26027
rect 2728 25995 2760 26027
rect 2800 25995 2832 26027
rect 2872 25995 2904 26027
rect 2944 25995 2976 26027
rect 3016 25995 3048 26027
rect 3088 25995 3120 26027
rect 3160 25995 3192 26027
rect 3232 25995 3264 26027
rect 3304 25995 3336 26027
rect 3376 25995 3408 26027
rect 3448 25995 3480 26027
rect 3520 25995 3552 26027
rect 3592 25995 3624 26027
rect 3664 25995 3696 26027
rect 3736 25995 3768 26027
rect 3808 25995 3840 26027
rect 3880 25995 3912 26027
rect 3952 25995 3984 26027
rect 4024 25995 4056 26027
rect 4096 25995 4128 26027
rect 4168 25995 4200 26027
rect 4240 25995 4272 26027
rect 4312 25995 4344 26027
rect 4384 25995 4416 26027
rect 4456 25995 4488 26027
rect 4528 25995 4560 26027
rect 4600 25995 4632 26027
rect 4672 25995 4704 26027
rect 4744 25995 4776 26027
rect 4816 25995 4848 26027
rect 4888 25995 4920 26027
rect 4960 25995 4992 26027
rect 5032 25995 5064 26027
rect 5104 25995 5136 26027
rect 5176 25995 5208 26027
rect 5248 25995 5280 26027
rect 5320 25995 5352 26027
rect 5392 25995 5424 26027
rect 5464 25995 5496 26027
rect 5536 25995 5568 26027
rect 5608 25995 5640 26027
rect 5680 25995 5712 26027
rect 5752 25995 5784 26027
rect 5824 25995 5856 26027
rect 5896 25995 5928 26027
rect 5968 25995 6000 26027
rect 6040 25995 6072 26027
rect 6112 25995 6144 26027
rect 6184 25995 6216 26027
rect 6256 25995 6288 26027
rect 6328 25995 6360 26027
rect 6400 25995 6432 26027
rect 6472 25995 6504 26027
rect 6544 25995 6576 26027
rect 6616 25995 6648 26027
rect 6688 25995 6720 26027
rect 6760 25995 6792 26027
rect 6832 25995 6864 26027
rect 6904 25995 6936 26027
rect 6976 25995 7008 26027
rect 7048 25995 7080 26027
rect 7120 25995 7152 26027
rect 7192 25995 7224 26027
rect 7264 25995 7296 26027
rect 7336 25995 7368 26027
rect 7408 25995 7440 26027
rect 7480 25995 7512 26027
rect 7552 25995 7584 26027
rect 7624 25995 7656 26027
rect 7696 25995 7728 26027
rect 7768 25995 7800 26027
rect 7840 25995 7872 26027
rect 7912 25995 7944 26027
rect 7984 25995 8016 26027
rect 8056 25995 8088 26027
rect 8128 25995 8160 26027
rect 8200 25995 8232 26027
rect 8272 25995 8304 26027
rect 8344 25995 8376 26027
rect 8416 25995 8448 26027
rect 8488 25995 8520 26027
rect 8560 25995 8592 26027
rect 8632 25995 8664 26027
rect 8704 25995 8736 26027
rect 8776 25995 8808 26027
rect 8848 25995 8880 26027
rect 8920 25995 8952 26027
rect 8992 25995 9024 26027
rect 9064 25995 9096 26027
rect 9136 25995 9168 26027
rect 9208 25995 9240 26027
rect 9280 25995 9312 26027
rect 9352 25995 9384 26027
rect 9424 25995 9456 26027
rect 9496 25995 9528 26027
rect 9568 25995 9600 26027
rect 9640 25995 9672 26027
rect 9712 25995 9744 26027
rect 9784 25995 9816 26027
rect 9856 25995 9888 26027
rect 9928 25995 9960 26027
rect 10000 25995 10032 26027
rect 10072 25995 10104 26027
rect 10144 25995 10176 26027
rect 10216 25995 10248 26027
rect 10288 25995 10320 26027
rect 10360 25995 10392 26027
rect 10432 25995 10464 26027
rect 10504 25995 10536 26027
rect 10576 25995 10608 26027
rect 10648 25995 10680 26027
rect 10720 25995 10752 26027
rect 10792 25995 10824 26027
rect 10864 25995 10896 26027
rect 10936 25995 10968 26027
rect 11008 25995 11040 26027
rect 11080 25995 11112 26027
rect 11152 25995 11184 26027
rect 11224 25995 11256 26027
rect 11296 25995 11328 26027
rect 11368 25995 11400 26027
rect 11440 25995 11472 26027
rect 11512 25995 11544 26027
rect 11584 25995 11616 26027
rect 11656 25995 11688 26027
rect 11728 25995 11760 26027
rect 11800 25995 11832 26027
rect 11872 25995 11904 26027
rect 11944 25995 11976 26027
rect 12016 25995 12048 26027
rect 12088 25995 12120 26027
rect 12160 25995 12192 26027
rect 12232 25995 12264 26027
rect 12304 25995 12336 26027
rect 12376 25995 12408 26027
rect 12448 25995 12480 26027
rect 12520 25995 12552 26027
rect 12592 25995 12624 26027
rect 12664 25995 12696 26027
rect 12736 25995 12768 26027
rect 12808 25995 12840 26027
rect 12880 25995 12912 26027
rect 12952 25995 12984 26027
rect 13024 25995 13056 26027
rect 13096 25995 13128 26027
rect 13168 25995 13200 26027
rect 13240 25995 13272 26027
rect 13312 25995 13344 26027
rect 13384 25995 13416 26027
rect 13456 25995 13488 26027
rect 13528 25995 13560 26027
rect 13600 25995 13632 26027
rect 13672 25995 13704 26027
rect 13744 25995 13776 26027
rect 13816 25995 13848 26027
rect 13888 25995 13920 26027
rect 13960 25995 13992 26027
rect 14032 25995 14064 26027
rect 14104 25995 14136 26027
rect 14176 25995 14208 26027
rect 14248 25995 14280 26027
rect 14320 25995 14352 26027
rect 14392 25995 14424 26027
rect 14464 25995 14496 26027
rect 14536 25995 14568 26027
rect 14608 25995 14640 26027
rect 14680 25995 14712 26027
rect 14752 25995 14784 26027
rect 14824 25995 14856 26027
rect 14896 25995 14928 26027
rect 14968 25995 15000 26027
rect 15040 25995 15072 26027
rect 15112 25995 15144 26027
rect 15184 25995 15216 26027
rect 15256 25995 15288 26027
rect 15328 25995 15360 26027
rect 15400 25995 15432 26027
rect 15472 25995 15504 26027
rect 15544 25995 15576 26027
rect 15616 25995 15648 26027
rect 15688 25995 15720 26027
rect 15760 25995 15792 26027
rect 15832 25995 15864 26027
rect 15904 25995 15936 26027
rect 64 25923 96 25955
rect 136 25923 168 25955
rect 208 25923 240 25955
rect 280 25923 312 25955
rect 352 25923 384 25955
rect 424 25923 456 25955
rect 496 25923 528 25955
rect 568 25923 600 25955
rect 640 25923 672 25955
rect 712 25923 744 25955
rect 784 25923 816 25955
rect 856 25923 888 25955
rect 928 25923 960 25955
rect 1000 25923 1032 25955
rect 1072 25923 1104 25955
rect 1144 25923 1176 25955
rect 1216 25923 1248 25955
rect 1288 25923 1320 25955
rect 1360 25923 1392 25955
rect 1432 25923 1464 25955
rect 1504 25923 1536 25955
rect 1576 25923 1608 25955
rect 1648 25923 1680 25955
rect 1720 25923 1752 25955
rect 1792 25923 1824 25955
rect 1864 25923 1896 25955
rect 1936 25923 1968 25955
rect 2008 25923 2040 25955
rect 2080 25923 2112 25955
rect 2152 25923 2184 25955
rect 2224 25923 2256 25955
rect 2296 25923 2328 25955
rect 2368 25923 2400 25955
rect 2440 25923 2472 25955
rect 2512 25923 2544 25955
rect 2584 25923 2616 25955
rect 2656 25923 2688 25955
rect 2728 25923 2760 25955
rect 2800 25923 2832 25955
rect 2872 25923 2904 25955
rect 2944 25923 2976 25955
rect 3016 25923 3048 25955
rect 3088 25923 3120 25955
rect 3160 25923 3192 25955
rect 3232 25923 3264 25955
rect 3304 25923 3336 25955
rect 3376 25923 3408 25955
rect 3448 25923 3480 25955
rect 3520 25923 3552 25955
rect 3592 25923 3624 25955
rect 3664 25923 3696 25955
rect 3736 25923 3768 25955
rect 3808 25923 3840 25955
rect 3880 25923 3912 25955
rect 3952 25923 3984 25955
rect 4024 25923 4056 25955
rect 4096 25923 4128 25955
rect 4168 25923 4200 25955
rect 4240 25923 4272 25955
rect 4312 25923 4344 25955
rect 4384 25923 4416 25955
rect 4456 25923 4488 25955
rect 4528 25923 4560 25955
rect 4600 25923 4632 25955
rect 4672 25923 4704 25955
rect 4744 25923 4776 25955
rect 4816 25923 4848 25955
rect 4888 25923 4920 25955
rect 4960 25923 4992 25955
rect 5032 25923 5064 25955
rect 5104 25923 5136 25955
rect 5176 25923 5208 25955
rect 5248 25923 5280 25955
rect 5320 25923 5352 25955
rect 5392 25923 5424 25955
rect 5464 25923 5496 25955
rect 5536 25923 5568 25955
rect 5608 25923 5640 25955
rect 5680 25923 5712 25955
rect 5752 25923 5784 25955
rect 5824 25923 5856 25955
rect 5896 25923 5928 25955
rect 5968 25923 6000 25955
rect 6040 25923 6072 25955
rect 6112 25923 6144 25955
rect 6184 25923 6216 25955
rect 6256 25923 6288 25955
rect 6328 25923 6360 25955
rect 6400 25923 6432 25955
rect 6472 25923 6504 25955
rect 6544 25923 6576 25955
rect 6616 25923 6648 25955
rect 6688 25923 6720 25955
rect 6760 25923 6792 25955
rect 6832 25923 6864 25955
rect 6904 25923 6936 25955
rect 6976 25923 7008 25955
rect 7048 25923 7080 25955
rect 7120 25923 7152 25955
rect 7192 25923 7224 25955
rect 7264 25923 7296 25955
rect 7336 25923 7368 25955
rect 7408 25923 7440 25955
rect 7480 25923 7512 25955
rect 7552 25923 7584 25955
rect 7624 25923 7656 25955
rect 7696 25923 7728 25955
rect 7768 25923 7800 25955
rect 7840 25923 7872 25955
rect 7912 25923 7944 25955
rect 7984 25923 8016 25955
rect 8056 25923 8088 25955
rect 8128 25923 8160 25955
rect 8200 25923 8232 25955
rect 8272 25923 8304 25955
rect 8344 25923 8376 25955
rect 8416 25923 8448 25955
rect 8488 25923 8520 25955
rect 8560 25923 8592 25955
rect 8632 25923 8664 25955
rect 8704 25923 8736 25955
rect 8776 25923 8808 25955
rect 8848 25923 8880 25955
rect 8920 25923 8952 25955
rect 8992 25923 9024 25955
rect 9064 25923 9096 25955
rect 9136 25923 9168 25955
rect 9208 25923 9240 25955
rect 9280 25923 9312 25955
rect 9352 25923 9384 25955
rect 9424 25923 9456 25955
rect 9496 25923 9528 25955
rect 9568 25923 9600 25955
rect 9640 25923 9672 25955
rect 9712 25923 9744 25955
rect 9784 25923 9816 25955
rect 9856 25923 9888 25955
rect 9928 25923 9960 25955
rect 10000 25923 10032 25955
rect 10072 25923 10104 25955
rect 10144 25923 10176 25955
rect 10216 25923 10248 25955
rect 10288 25923 10320 25955
rect 10360 25923 10392 25955
rect 10432 25923 10464 25955
rect 10504 25923 10536 25955
rect 10576 25923 10608 25955
rect 10648 25923 10680 25955
rect 10720 25923 10752 25955
rect 10792 25923 10824 25955
rect 10864 25923 10896 25955
rect 10936 25923 10968 25955
rect 11008 25923 11040 25955
rect 11080 25923 11112 25955
rect 11152 25923 11184 25955
rect 11224 25923 11256 25955
rect 11296 25923 11328 25955
rect 11368 25923 11400 25955
rect 11440 25923 11472 25955
rect 11512 25923 11544 25955
rect 11584 25923 11616 25955
rect 11656 25923 11688 25955
rect 11728 25923 11760 25955
rect 11800 25923 11832 25955
rect 11872 25923 11904 25955
rect 11944 25923 11976 25955
rect 12016 25923 12048 25955
rect 12088 25923 12120 25955
rect 12160 25923 12192 25955
rect 12232 25923 12264 25955
rect 12304 25923 12336 25955
rect 12376 25923 12408 25955
rect 12448 25923 12480 25955
rect 12520 25923 12552 25955
rect 12592 25923 12624 25955
rect 12664 25923 12696 25955
rect 12736 25923 12768 25955
rect 12808 25923 12840 25955
rect 12880 25923 12912 25955
rect 12952 25923 12984 25955
rect 13024 25923 13056 25955
rect 13096 25923 13128 25955
rect 13168 25923 13200 25955
rect 13240 25923 13272 25955
rect 13312 25923 13344 25955
rect 13384 25923 13416 25955
rect 13456 25923 13488 25955
rect 13528 25923 13560 25955
rect 13600 25923 13632 25955
rect 13672 25923 13704 25955
rect 13744 25923 13776 25955
rect 13816 25923 13848 25955
rect 13888 25923 13920 25955
rect 13960 25923 13992 25955
rect 14032 25923 14064 25955
rect 14104 25923 14136 25955
rect 14176 25923 14208 25955
rect 14248 25923 14280 25955
rect 14320 25923 14352 25955
rect 14392 25923 14424 25955
rect 14464 25923 14496 25955
rect 14536 25923 14568 25955
rect 14608 25923 14640 25955
rect 14680 25923 14712 25955
rect 14752 25923 14784 25955
rect 14824 25923 14856 25955
rect 14896 25923 14928 25955
rect 14968 25923 15000 25955
rect 15040 25923 15072 25955
rect 15112 25923 15144 25955
rect 15184 25923 15216 25955
rect 15256 25923 15288 25955
rect 15328 25923 15360 25955
rect 15400 25923 15432 25955
rect 15472 25923 15504 25955
rect 15544 25923 15576 25955
rect 15616 25923 15648 25955
rect 15688 25923 15720 25955
rect 15760 25923 15792 25955
rect 15832 25923 15864 25955
rect 15904 25923 15936 25955
rect 64 25851 96 25883
rect 136 25851 168 25883
rect 208 25851 240 25883
rect 280 25851 312 25883
rect 352 25851 384 25883
rect 424 25851 456 25883
rect 496 25851 528 25883
rect 568 25851 600 25883
rect 640 25851 672 25883
rect 712 25851 744 25883
rect 784 25851 816 25883
rect 856 25851 888 25883
rect 928 25851 960 25883
rect 1000 25851 1032 25883
rect 1072 25851 1104 25883
rect 1144 25851 1176 25883
rect 1216 25851 1248 25883
rect 1288 25851 1320 25883
rect 1360 25851 1392 25883
rect 1432 25851 1464 25883
rect 1504 25851 1536 25883
rect 1576 25851 1608 25883
rect 1648 25851 1680 25883
rect 1720 25851 1752 25883
rect 1792 25851 1824 25883
rect 1864 25851 1896 25883
rect 1936 25851 1968 25883
rect 2008 25851 2040 25883
rect 2080 25851 2112 25883
rect 2152 25851 2184 25883
rect 2224 25851 2256 25883
rect 2296 25851 2328 25883
rect 2368 25851 2400 25883
rect 2440 25851 2472 25883
rect 2512 25851 2544 25883
rect 2584 25851 2616 25883
rect 2656 25851 2688 25883
rect 2728 25851 2760 25883
rect 2800 25851 2832 25883
rect 2872 25851 2904 25883
rect 2944 25851 2976 25883
rect 3016 25851 3048 25883
rect 3088 25851 3120 25883
rect 3160 25851 3192 25883
rect 3232 25851 3264 25883
rect 3304 25851 3336 25883
rect 3376 25851 3408 25883
rect 3448 25851 3480 25883
rect 3520 25851 3552 25883
rect 3592 25851 3624 25883
rect 3664 25851 3696 25883
rect 3736 25851 3768 25883
rect 3808 25851 3840 25883
rect 3880 25851 3912 25883
rect 3952 25851 3984 25883
rect 4024 25851 4056 25883
rect 4096 25851 4128 25883
rect 4168 25851 4200 25883
rect 4240 25851 4272 25883
rect 4312 25851 4344 25883
rect 4384 25851 4416 25883
rect 4456 25851 4488 25883
rect 4528 25851 4560 25883
rect 4600 25851 4632 25883
rect 4672 25851 4704 25883
rect 4744 25851 4776 25883
rect 4816 25851 4848 25883
rect 4888 25851 4920 25883
rect 4960 25851 4992 25883
rect 5032 25851 5064 25883
rect 5104 25851 5136 25883
rect 5176 25851 5208 25883
rect 5248 25851 5280 25883
rect 5320 25851 5352 25883
rect 5392 25851 5424 25883
rect 5464 25851 5496 25883
rect 5536 25851 5568 25883
rect 5608 25851 5640 25883
rect 5680 25851 5712 25883
rect 5752 25851 5784 25883
rect 5824 25851 5856 25883
rect 5896 25851 5928 25883
rect 5968 25851 6000 25883
rect 6040 25851 6072 25883
rect 6112 25851 6144 25883
rect 6184 25851 6216 25883
rect 6256 25851 6288 25883
rect 6328 25851 6360 25883
rect 6400 25851 6432 25883
rect 6472 25851 6504 25883
rect 6544 25851 6576 25883
rect 6616 25851 6648 25883
rect 6688 25851 6720 25883
rect 6760 25851 6792 25883
rect 6832 25851 6864 25883
rect 6904 25851 6936 25883
rect 6976 25851 7008 25883
rect 7048 25851 7080 25883
rect 7120 25851 7152 25883
rect 7192 25851 7224 25883
rect 7264 25851 7296 25883
rect 7336 25851 7368 25883
rect 7408 25851 7440 25883
rect 7480 25851 7512 25883
rect 7552 25851 7584 25883
rect 7624 25851 7656 25883
rect 7696 25851 7728 25883
rect 7768 25851 7800 25883
rect 7840 25851 7872 25883
rect 7912 25851 7944 25883
rect 7984 25851 8016 25883
rect 8056 25851 8088 25883
rect 8128 25851 8160 25883
rect 8200 25851 8232 25883
rect 8272 25851 8304 25883
rect 8344 25851 8376 25883
rect 8416 25851 8448 25883
rect 8488 25851 8520 25883
rect 8560 25851 8592 25883
rect 8632 25851 8664 25883
rect 8704 25851 8736 25883
rect 8776 25851 8808 25883
rect 8848 25851 8880 25883
rect 8920 25851 8952 25883
rect 8992 25851 9024 25883
rect 9064 25851 9096 25883
rect 9136 25851 9168 25883
rect 9208 25851 9240 25883
rect 9280 25851 9312 25883
rect 9352 25851 9384 25883
rect 9424 25851 9456 25883
rect 9496 25851 9528 25883
rect 9568 25851 9600 25883
rect 9640 25851 9672 25883
rect 9712 25851 9744 25883
rect 9784 25851 9816 25883
rect 9856 25851 9888 25883
rect 9928 25851 9960 25883
rect 10000 25851 10032 25883
rect 10072 25851 10104 25883
rect 10144 25851 10176 25883
rect 10216 25851 10248 25883
rect 10288 25851 10320 25883
rect 10360 25851 10392 25883
rect 10432 25851 10464 25883
rect 10504 25851 10536 25883
rect 10576 25851 10608 25883
rect 10648 25851 10680 25883
rect 10720 25851 10752 25883
rect 10792 25851 10824 25883
rect 10864 25851 10896 25883
rect 10936 25851 10968 25883
rect 11008 25851 11040 25883
rect 11080 25851 11112 25883
rect 11152 25851 11184 25883
rect 11224 25851 11256 25883
rect 11296 25851 11328 25883
rect 11368 25851 11400 25883
rect 11440 25851 11472 25883
rect 11512 25851 11544 25883
rect 11584 25851 11616 25883
rect 11656 25851 11688 25883
rect 11728 25851 11760 25883
rect 11800 25851 11832 25883
rect 11872 25851 11904 25883
rect 11944 25851 11976 25883
rect 12016 25851 12048 25883
rect 12088 25851 12120 25883
rect 12160 25851 12192 25883
rect 12232 25851 12264 25883
rect 12304 25851 12336 25883
rect 12376 25851 12408 25883
rect 12448 25851 12480 25883
rect 12520 25851 12552 25883
rect 12592 25851 12624 25883
rect 12664 25851 12696 25883
rect 12736 25851 12768 25883
rect 12808 25851 12840 25883
rect 12880 25851 12912 25883
rect 12952 25851 12984 25883
rect 13024 25851 13056 25883
rect 13096 25851 13128 25883
rect 13168 25851 13200 25883
rect 13240 25851 13272 25883
rect 13312 25851 13344 25883
rect 13384 25851 13416 25883
rect 13456 25851 13488 25883
rect 13528 25851 13560 25883
rect 13600 25851 13632 25883
rect 13672 25851 13704 25883
rect 13744 25851 13776 25883
rect 13816 25851 13848 25883
rect 13888 25851 13920 25883
rect 13960 25851 13992 25883
rect 14032 25851 14064 25883
rect 14104 25851 14136 25883
rect 14176 25851 14208 25883
rect 14248 25851 14280 25883
rect 14320 25851 14352 25883
rect 14392 25851 14424 25883
rect 14464 25851 14496 25883
rect 14536 25851 14568 25883
rect 14608 25851 14640 25883
rect 14680 25851 14712 25883
rect 14752 25851 14784 25883
rect 14824 25851 14856 25883
rect 14896 25851 14928 25883
rect 14968 25851 15000 25883
rect 15040 25851 15072 25883
rect 15112 25851 15144 25883
rect 15184 25851 15216 25883
rect 15256 25851 15288 25883
rect 15328 25851 15360 25883
rect 15400 25851 15432 25883
rect 15472 25851 15504 25883
rect 15544 25851 15576 25883
rect 15616 25851 15648 25883
rect 15688 25851 15720 25883
rect 15760 25851 15792 25883
rect 15832 25851 15864 25883
rect 15904 25851 15936 25883
rect 64 25779 96 25811
rect 136 25779 168 25811
rect 208 25779 240 25811
rect 280 25779 312 25811
rect 352 25779 384 25811
rect 424 25779 456 25811
rect 496 25779 528 25811
rect 568 25779 600 25811
rect 640 25779 672 25811
rect 712 25779 744 25811
rect 784 25779 816 25811
rect 856 25779 888 25811
rect 928 25779 960 25811
rect 1000 25779 1032 25811
rect 1072 25779 1104 25811
rect 1144 25779 1176 25811
rect 1216 25779 1248 25811
rect 1288 25779 1320 25811
rect 1360 25779 1392 25811
rect 1432 25779 1464 25811
rect 1504 25779 1536 25811
rect 1576 25779 1608 25811
rect 1648 25779 1680 25811
rect 1720 25779 1752 25811
rect 1792 25779 1824 25811
rect 1864 25779 1896 25811
rect 1936 25779 1968 25811
rect 2008 25779 2040 25811
rect 2080 25779 2112 25811
rect 2152 25779 2184 25811
rect 2224 25779 2256 25811
rect 2296 25779 2328 25811
rect 2368 25779 2400 25811
rect 2440 25779 2472 25811
rect 2512 25779 2544 25811
rect 2584 25779 2616 25811
rect 2656 25779 2688 25811
rect 2728 25779 2760 25811
rect 2800 25779 2832 25811
rect 2872 25779 2904 25811
rect 2944 25779 2976 25811
rect 3016 25779 3048 25811
rect 3088 25779 3120 25811
rect 3160 25779 3192 25811
rect 3232 25779 3264 25811
rect 3304 25779 3336 25811
rect 3376 25779 3408 25811
rect 3448 25779 3480 25811
rect 3520 25779 3552 25811
rect 3592 25779 3624 25811
rect 3664 25779 3696 25811
rect 3736 25779 3768 25811
rect 3808 25779 3840 25811
rect 3880 25779 3912 25811
rect 3952 25779 3984 25811
rect 4024 25779 4056 25811
rect 4096 25779 4128 25811
rect 4168 25779 4200 25811
rect 4240 25779 4272 25811
rect 4312 25779 4344 25811
rect 4384 25779 4416 25811
rect 4456 25779 4488 25811
rect 4528 25779 4560 25811
rect 4600 25779 4632 25811
rect 4672 25779 4704 25811
rect 4744 25779 4776 25811
rect 4816 25779 4848 25811
rect 4888 25779 4920 25811
rect 4960 25779 4992 25811
rect 5032 25779 5064 25811
rect 5104 25779 5136 25811
rect 5176 25779 5208 25811
rect 5248 25779 5280 25811
rect 5320 25779 5352 25811
rect 5392 25779 5424 25811
rect 5464 25779 5496 25811
rect 5536 25779 5568 25811
rect 5608 25779 5640 25811
rect 5680 25779 5712 25811
rect 5752 25779 5784 25811
rect 5824 25779 5856 25811
rect 5896 25779 5928 25811
rect 5968 25779 6000 25811
rect 6040 25779 6072 25811
rect 6112 25779 6144 25811
rect 6184 25779 6216 25811
rect 6256 25779 6288 25811
rect 6328 25779 6360 25811
rect 6400 25779 6432 25811
rect 6472 25779 6504 25811
rect 6544 25779 6576 25811
rect 6616 25779 6648 25811
rect 6688 25779 6720 25811
rect 6760 25779 6792 25811
rect 6832 25779 6864 25811
rect 6904 25779 6936 25811
rect 6976 25779 7008 25811
rect 7048 25779 7080 25811
rect 7120 25779 7152 25811
rect 7192 25779 7224 25811
rect 7264 25779 7296 25811
rect 7336 25779 7368 25811
rect 7408 25779 7440 25811
rect 7480 25779 7512 25811
rect 7552 25779 7584 25811
rect 7624 25779 7656 25811
rect 7696 25779 7728 25811
rect 7768 25779 7800 25811
rect 7840 25779 7872 25811
rect 7912 25779 7944 25811
rect 7984 25779 8016 25811
rect 8056 25779 8088 25811
rect 8128 25779 8160 25811
rect 8200 25779 8232 25811
rect 8272 25779 8304 25811
rect 8344 25779 8376 25811
rect 8416 25779 8448 25811
rect 8488 25779 8520 25811
rect 8560 25779 8592 25811
rect 8632 25779 8664 25811
rect 8704 25779 8736 25811
rect 8776 25779 8808 25811
rect 8848 25779 8880 25811
rect 8920 25779 8952 25811
rect 8992 25779 9024 25811
rect 9064 25779 9096 25811
rect 9136 25779 9168 25811
rect 9208 25779 9240 25811
rect 9280 25779 9312 25811
rect 9352 25779 9384 25811
rect 9424 25779 9456 25811
rect 9496 25779 9528 25811
rect 9568 25779 9600 25811
rect 9640 25779 9672 25811
rect 9712 25779 9744 25811
rect 9784 25779 9816 25811
rect 9856 25779 9888 25811
rect 9928 25779 9960 25811
rect 10000 25779 10032 25811
rect 10072 25779 10104 25811
rect 10144 25779 10176 25811
rect 10216 25779 10248 25811
rect 10288 25779 10320 25811
rect 10360 25779 10392 25811
rect 10432 25779 10464 25811
rect 10504 25779 10536 25811
rect 10576 25779 10608 25811
rect 10648 25779 10680 25811
rect 10720 25779 10752 25811
rect 10792 25779 10824 25811
rect 10864 25779 10896 25811
rect 10936 25779 10968 25811
rect 11008 25779 11040 25811
rect 11080 25779 11112 25811
rect 11152 25779 11184 25811
rect 11224 25779 11256 25811
rect 11296 25779 11328 25811
rect 11368 25779 11400 25811
rect 11440 25779 11472 25811
rect 11512 25779 11544 25811
rect 11584 25779 11616 25811
rect 11656 25779 11688 25811
rect 11728 25779 11760 25811
rect 11800 25779 11832 25811
rect 11872 25779 11904 25811
rect 11944 25779 11976 25811
rect 12016 25779 12048 25811
rect 12088 25779 12120 25811
rect 12160 25779 12192 25811
rect 12232 25779 12264 25811
rect 12304 25779 12336 25811
rect 12376 25779 12408 25811
rect 12448 25779 12480 25811
rect 12520 25779 12552 25811
rect 12592 25779 12624 25811
rect 12664 25779 12696 25811
rect 12736 25779 12768 25811
rect 12808 25779 12840 25811
rect 12880 25779 12912 25811
rect 12952 25779 12984 25811
rect 13024 25779 13056 25811
rect 13096 25779 13128 25811
rect 13168 25779 13200 25811
rect 13240 25779 13272 25811
rect 13312 25779 13344 25811
rect 13384 25779 13416 25811
rect 13456 25779 13488 25811
rect 13528 25779 13560 25811
rect 13600 25779 13632 25811
rect 13672 25779 13704 25811
rect 13744 25779 13776 25811
rect 13816 25779 13848 25811
rect 13888 25779 13920 25811
rect 13960 25779 13992 25811
rect 14032 25779 14064 25811
rect 14104 25779 14136 25811
rect 14176 25779 14208 25811
rect 14248 25779 14280 25811
rect 14320 25779 14352 25811
rect 14392 25779 14424 25811
rect 14464 25779 14496 25811
rect 14536 25779 14568 25811
rect 14608 25779 14640 25811
rect 14680 25779 14712 25811
rect 14752 25779 14784 25811
rect 14824 25779 14856 25811
rect 14896 25779 14928 25811
rect 14968 25779 15000 25811
rect 15040 25779 15072 25811
rect 15112 25779 15144 25811
rect 15184 25779 15216 25811
rect 15256 25779 15288 25811
rect 15328 25779 15360 25811
rect 15400 25779 15432 25811
rect 15472 25779 15504 25811
rect 15544 25779 15576 25811
rect 15616 25779 15648 25811
rect 15688 25779 15720 25811
rect 15760 25779 15792 25811
rect 15832 25779 15864 25811
rect 15904 25779 15936 25811
rect 64 25707 96 25739
rect 136 25707 168 25739
rect 208 25707 240 25739
rect 280 25707 312 25739
rect 352 25707 384 25739
rect 424 25707 456 25739
rect 496 25707 528 25739
rect 568 25707 600 25739
rect 640 25707 672 25739
rect 712 25707 744 25739
rect 784 25707 816 25739
rect 856 25707 888 25739
rect 928 25707 960 25739
rect 1000 25707 1032 25739
rect 1072 25707 1104 25739
rect 1144 25707 1176 25739
rect 1216 25707 1248 25739
rect 1288 25707 1320 25739
rect 1360 25707 1392 25739
rect 1432 25707 1464 25739
rect 1504 25707 1536 25739
rect 1576 25707 1608 25739
rect 1648 25707 1680 25739
rect 1720 25707 1752 25739
rect 1792 25707 1824 25739
rect 1864 25707 1896 25739
rect 1936 25707 1968 25739
rect 2008 25707 2040 25739
rect 2080 25707 2112 25739
rect 2152 25707 2184 25739
rect 2224 25707 2256 25739
rect 2296 25707 2328 25739
rect 2368 25707 2400 25739
rect 2440 25707 2472 25739
rect 2512 25707 2544 25739
rect 2584 25707 2616 25739
rect 2656 25707 2688 25739
rect 2728 25707 2760 25739
rect 2800 25707 2832 25739
rect 2872 25707 2904 25739
rect 2944 25707 2976 25739
rect 3016 25707 3048 25739
rect 3088 25707 3120 25739
rect 3160 25707 3192 25739
rect 3232 25707 3264 25739
rect 3304 25707 3336 25739
rect 3376 25707 3408 25739
rect 3448 25707 3480 25739
rect 3520 25707 3552 25739
rect 3592 25707 3624 25739
rect 3664 25707 3696 25739
rect 3736 25707 3768 25739
rect 3808 25707 3840 25739
rect 3880 25707 3912 25739
rect 3952 25707 3984 25739
rect 4024 25707 4056 25739
rect 4096 25707 4128 25739
rect 4168 25707 4200 25739
rect 4240 25707 4272 25739
rect 4312 25707 4344 25739
rect 4384 25707 4416 25739
rect 4456 25707 4488 25739
rect 4528 25707 4560 25739
rect 4600 25707 4632 25739
rect 4672 25707 4704 25739
rect 4744 25707 4776 25739
rect 4816 25707 4848 25739
rect 4888 25707 4920 25739
rect 4960 25707 4992 25739
rect 5032 25707 5064 25739
rect 5104 25707 5136 25739
rect 5176 25707 5208 25739
rect 5248 25707 5280 25739
rect 5320 25707 5352 25739
rect 5392 25707 5424 25739
rect 5464 25707 5496 25739
rect 5536 25707 5568 25739
rect 5608 25707 5640 25739
rect 5680 25707 5712 25739
rect 5752 25707 5784 25739
rect 5824 25707 5856 25739
rect 5896 25707 5928 25739
rect 5968 25707 6000 25739
rect 6040 25707 6072 25739
rect 6112 25707 6144 25739
rect 6184 25707 6216 25739
rect 6256 25707 6288 25739
rect 6328 25707 6360 25739
rect 6400 25707 6432 25739
rect 6472 25707 6504 25739
rect 6544 25707 6576 25739
rect 6616 25707 6648 25739
rect 6688 25707 6720 25739
rect 6760 25707 6792 25739
rect 6832 25707 6864 25739
rect 6904 25707 6936 25739
rect 6976 25707 7008 25739
rect 7048 25707 7080 25739
rect 7120 25707 7152 25739
rect 7192 25707 7224 25739
rect 7264 25707 7296 25739
rect 7336 25707 7368 25739
rect 7408 25707 7440 25739
rect 7480 25707 7512 25739
rect 7552 25707 7584 25739
rect 7624 25707 7656 25739
rect 7696 25707 7728 25739
rect 7768 25707 7800 25739
rect 7840 25707 7872 25739
rect 7912 25707 7944 25739
rect 7984 25707 8016 25739
rect 8056 25707 8088 25739
rect 8128 25707 8160 25739
rect 8200 25707 8232 25739
rect 8272 25707 8304 25739
rect 8344 25707 8376 25739
rect 8416 25707 8448 25739
rect 8488 25707 8520 25739
rect 8560 25707 8592 25739
rect 8632 25707 8664 25739
rect 8704 25707 8736 25739
rect 8776 25707 8808 25739
rect 8848 25707 8880 25739
rect 8920 25707 8952 25739
rect 8992 25707 9024 25739
rect 9064 25707 9096 25739
rect 9136 25707 9168 25739
rect 9208 25707 9240 25739
rect 9280 25707 9312 25739
rect 9352 25707 9384 25739
rect 9424 25707 9456 25739
rect 9496 25707 9528 25739
rect 9568 25707 9600 25739
rect 9640 25707 9672 25739
rect 9712 25707 9744 25739
rect 9784 25707 9816 25739
rect 9856 25707 9888 25739
rect 9928 25707 9960 25739
rect 10000 25707 10032 25739
rect 10072 25707 10104 25739
rect 10144 25707 10176 25739
rect 10216 25707 10248 25739
rect 10288 25707 10320 25739
rect 10360 25707 10392 25739
rect 10432 25707 10464 25739
rect 10504 25707 10536 25739
rect 10576 25707 10608 25739
rect 10648 25707 10680 25739
rect 10720 25707 10752 25739
rect 10792 25707 10824 25739
rect 10864 25707 10896 25739
rect 10936 25707 10968 25739
rect 11008 25707 11040 25739
rect 11080 25707 11112 25739
rect 11152 25707 11184 25739
rect 11224 25707 11256 25739
rect 11296 25707 11328 25739
rect 11368 25707 11400 25739
rect 11440 25707 11472 25739
rect 11512 25707 11544 25739
rect 11584 25707 11616 25739
rect 11656 25707 11688 25739
rect 11728 25707 11760 25739
rect 11800 25707 11832 25739
rect 11872 25707 11904 25739
rect 11944 25707 11976 25739
rect 12016 25707 12048 25739
rect 12088 25707 12120 25739
rect 12160 25707 12192 25739
rect 12232 25707 12264 25739
rect 12304 25707 12336 25739
rect 12376 25707 12408 25739
rect 12448 25707 12480 25739
rect 12520 25707 12552 25739
rect 12592 25707 12624 25739
rect 12664 25707 12696 25739
rect 12736 25707 12768 25739
rect 12808 25707 12840 25739
rect 12880 25707 12912 25739
rect 12952 25707 12984 25739
rect 13024 25707 13056 25739
rect 13096 25707 13128 25739
rect 13168 25707 13200 25739
rect 13240 25707 13272 25739
rect 13312 25707 13344 25739
rect 13384 25707 13416 25739
rect 13456 25707 13488 25739
rect 13528 25707 13560 25739
rect 13600 25707 13632 25739
rect 13672 25707 13704 25739
rect 13744 25707 13776 25739
rect 13816 25707 13848 25739
rect 13888 25707 13920 25739
rect 13960 25707 13992 25739
rect 14032 25707 14064 25739
rect 14104 25707 14136 25739
rect 14176 25707 14208 25739
rect 14248 25707 14280 25739
rect 14320 25707 14352 25739
rect 14392 25707 14424 25739
rect 14464 25707 14496 25739
rect 14536 25707 14568 25739
rect 14608 25707 14640 25739
rect 14680 25707 14712 25739
rect 14752 25707 14784 25739
rect 14824 25707 14856 25739
rect 14896 25707 14928 25739
rect 14968 25707 15000 25739
rect 15040 25707 15072 25739
rect 15112 25707 15144 25739
rect 15184 25707 15216 25739
rect 15256 25707 15288 25739
rect 15328 25707 15360 25739
rect 15400 25707 15432 25739
rect 15472 25707 15504 25739
rect 15544 25707 15576 25739
rect 15616 25707 15648 25739
rect 15688 25707 15720 25739
rect 15760 25707 15792 25739
rect 15832 25707 15864 25739
rect 15904 25707 15936 25739
rect 64 25635 96 25667
rect 136 25635 168 25667
rect 208 25635 240 25667
rect 280 25635 312 25667
rect 352 25635 384 25667
rect 424 25635 456 25667
rect 496 25635 528 25667
rect 568 25635 600 25667
rect 640 25635 672 25667
rect 712 25635 744 25667
rect 784 25635 816 25667
rect 856 25635 888 25667
rect 928 25635 960 25667
rect 1000 25635 1032 25667
rect 1072 25635 1104 25667
rect 1144 25635 1176 25667
rect 1216 25635 1248 25667
rect 1288 25635 1320 25667
rect 1360 25635 1392 25667
rect 1432 25635 1464 25667
rect 1504 25635 1536 25667
rect 1576 25635 1608 25667
rect 1648 25635 1680 25667
rect 1720 25635 1752 25667
rect 1792 25635 1824 25667
rect 1864 25635 1896 25667
rect 1936 25635 1968 25667
rect 2008 25635 2040 25667
rect 2080 25635 2112 25667
rect 2152 25635 2184 25667
rect 2224 25635 2256 25667
rect 2296 25635 2328 25667
rect 2368 25635 2400 25667
rect 2440 25635 2472 25667
rect 2512 25635 2544 25667
rect 2584 25635 2616 25667
rect 2656 25635 2688 25667
rect 2728 25635 2760 25667
rect 2800 25635 2832 25667
rect 2872 25635 2904 25667
rect 2944 25635 2976 25667
rect 3016 25635 3048 25667
rect 3088 25635 3120 25667
rect 3160 25635 3192 25667
rect 3232 25635 3264 25667
rect 3304 25635 3336 25667
rect 3376 25635 3408 25667
rect 3448 25635 3480 25667
rect 3520 25635 3552 25667
rect 3592 25635 3624 25667
rect 3664 25635 3696 25667
rect 3736 25635 3768 25667
rect 3808 25635 3840 25667
rect 3880 25635 3912 25667
rect 3952 25635 3984 25667
rect 4024 25635 4056 25667
rect 4096 25635 4128 25667
rect 4168 25635 4200 25667
rect 4240 25635 4272 25667
rect 4312 25635 4344 25667
rect 4384 25635 4416 25667
rect 4456 25635 4488 25667
rect 4528 25635 4560 25667
rect 4600 25635 4632 25667
rect 4672 25635 4704 25667
rect 4744 25635 4776 25667
rect 4816 25635 4848 25667
rect 4888 25635 4920 25667
rect 4960 25635 4992 25667
rect 5032 25635 5064 25667
rect 5104 25635 5136 25667
rect 5176 25635 5208 25667
rect 5248 25635 5280 25667
rect 5320 25635 5352 25667
rect 5392 25635 5424 25667
rect 5464 25635 5496 25667
rect 5536 25635 5568 25667
rect 5608 25635 5640 25667
rect 5680 25635 5712 25667
rect 5752 25635 5784 25667
rect 5824 25635 5856 25667
rect 5896 25635 5928 25667
rect 5968 25635 6000 25667
rect 6040 25635 6072 25667
rect 6112 25635 6144 25667
rect 6184 25635 6216 25667
rect 6256 25635 6288 25667
rect 6328 25635 6360 25667
rect 6400 25635 6432 25667
rect 6472 25635 6504 25667
rect 6544 25635 6576 25667
rect 6616 25635 6648 25667
rect 6688 25635 6720 25667
rect 6760 25635 6792 25667
rect 6832 25635 6864 25667
rect 6904 25635 6936 25667
rect 6976 25635 7008 25667
rect 7048 25635 7080 25667
rect 7120 25635 7152 25667
rect 7192 25635 7224 25667
rect 7264 25635 7296 25667
rect 7336 25635 7368 25667
rect 7408 25635 7440 25667
rect 7480 25635 7512 25667
rect 7552 25635 7584 25667
rect 7624 25635 7656 25667
rect 7696 25635 7728 25667
rect 7768 25635 7800 25667
rect 7840 25635 7872 25667
rect 7912 25635 7944 25667
rect 7984 25635 8016 25667
rect 8056 25635 8088 25667
rect 8128 25635 8160 25667
rect 8200 25635 8232 25667
rect 8272 25635 8304 25667
rect 8344 25635 8376 25667
rect 8416 25635 8448 25667
rect 8488 25635 8520 25667
rect 8560 25635 8592 25667
rect 8632 25635 8664 25667
rect 8704 25635 8736 25667
rect 8776 25635 8808 25667
rect 8848 25635 8880 25667
rect 8920 25635 8952 25667
rect 8992 25635 9024 25667
rect 9064 25635 9096 25667
rect 9136 25635 9168 25667
rect 9208 25635 9240 25667
rect 9280 25635 9312 25667
rect 9352 25635 9384 25667
rect 9424 25635 9456 25667
rect 9496 25635 9528 25667
rect 9568 25635 9600 25667
rect 9640 25635 9672 25667
rect 9712 25635 9744 25667
rect 9784 25635 9816 25667
rect 9856 25635 9888 25667
rect 9928 25635 9960 25667
rect 10000 25635 10032 25667
rect 10072 25635 10104 25667
rect 10144 25635 10176 25667
rect 10216 25635 10248 25667
rect 10288 25635 10320 25667
rect 10360 25635 10392 25667
rect 10432 25635 10464 25667
rect 10504 25635 10536 25667
rect 10576 25635 10608 25667
rect 10648 25635 10680 25667
rect 10720 25635 10752 25667
rect 10792 25635 10824 25667
rect 10864 25635 10896 25667
rect 10936 25635 10968 25667
rect 11008 25635 11040 25667
rect 11080 25635 11112 25667
rect 11152 25635 11184 25667
rect 11224 25635 11256 25667
rect 11296 25635 11328 25667
rect 11368 25635 11400 25667
rect 11440 25635 11472 25667
rect 11512 25635 11544 25667
rect 11584 25635 11616 25667
rect 11656 25635 11688 25667
rect 11728 25635 11760 25667
rect 11800 25635 11832 25667
rect 11872 25635 11904 25667
rect 11944 25635 11976 25667
rect 12016 25635 12048 25667
rect 12088 25635 12120 25667
rect 12160 25635 12192 25667
rect 12232 25635 12264 25667
rect 12304 25635 12336 25667
rect 12376 25635 12408 25667
rect 12448 25635 12480 25667
rect 12520 25635 12552 25667
rect 12592 25635 12624 25667
rect 12664 25635 12696 25667
rect 12736 25635 12768 25667
rect 12808 25635 12840 25667
rect 12880 25635 12912 25667
rect 12952 25635 12984 25667
rect 13024 25635 13056 25667
rect 13096 25635 13128 25667
rect 13168 25635 13200 25667
rect 13240 25635 13272 25667
rect 13312 25635 13344 25667
rect 13384 25635 13416 25667
rect 13456 25635 13488 25667
rect 13528 25635 13560 25667
rect 13600 25635 13632 25667
rect 13672 25635 13704 25667
rect 13744 25635 13776 25667
rect 13816 25635 13848 25667
rect 13888 25635 13920 25667
rect 13960 25635 13992 25667
rect 14032 25635 14064 25667
rect 14104 25635 14136 25667
rect 14176 25635 14208 25667
rect 14248 25635 14280 25667
rect 14320 25635 14352 25667
rect 14392 25635 14424 25667
rect 14464 25635 14496 25667
rect 14536 25635 14568 25667
rect 14608 25635 14640 25667
rect 14680 25635 14712 25667
rect 14752 25635 14784 25667
rect 14824 25635 14856 25667
rect 14896 25635 14928 25667
rect 14968 25635 15000 25667
rect 15040 25635 15072 25667
rect 15112 25635 15144 25667
rect 15184 25635 15216 25667
rect 15256 25635 15288 25667
rect 15328 25635 15360 25667
rect 15400 25635 15432 25667
rect 15472 25635 15504 25667
rect 15544 25635 15576 25667
rect 15616 25635 15648 25667
rect 15688 25635 15720 25667
rect 15760 25635 15792 25667
rect 15832 25635 15864 25667
rect 15904 25635 15936 25667
rect 64 25563 96 25595
rect 136 25563 168 25595
rect 208 25563 240 25595
rect 280 25563 312 25595
rect 352 25563 384 25595
rect 424 25563 456 25595
rect 496 25563 528 25595
rect 568 25563 600 25595
rect 640 25563 672 25595
rect 712 25563 744 25595
rect 784 25563 816 25595
rect 856 25563 888 25595
rect 928 25563 960 25595
rect 1000 25563 1032 25595
rect 1072 25563 1104 25595
rect 1144 25563 1176 25595
rect 1216 25563 1248 25595
rect 1288 25563 1320 25595
rect 1360 25563 1392 25595
rect 1432 25563 1464 25595
rect 1504 25563 1536 25595
rect 1576 25563 1608 25595
rect 1648 25563 1680 25595
rect 1720 25563 1752 25595
rect 1792 25563 1824 25595
rect 1864 25563 1896 25595
rect 1936 25563 1968 25595
rect 2008 25563 2040 25595
rect 2080 25563 2112 25595
rect 2152 25563 2184 25595
rect 2224 25563 2256 25595
rect 2296 25563 2328 25595
rect 2368 25563 2400 25595
rect 2440 25563 2472 25595
rect 2512 25563 2544 25595
rect 2584 25563 2616 25595
rect 2656 25563 2688 25595
rect 2728 25563 2760 25595
rect 2800 25563 2832 25595
rect 2872 25563 2904 25595
rect 2944 25563 2976 25595
rect 3016 25563 3048 25595
rect 3088 25563 3120 25595
rect 3160 25563 3192 25595
rect 3232 25563 3264 25595
rect 3304 25563 3336 25595
rect 3376 25563 3408 25595
rect 3448 25563 3480 25595
rect 3520 25563 3552 25595
rect 3592 25563 3624 25595
rect 3664 25563 3696 25595
rect 3736 25563 3768 25595
rect 3808 25563 3840 25595
rect 3880 25563 3912 25595
rect 3952 25563 3984 25595
rect 4024 25563 4056 25595
rect 4096 25563 4128 25595
rect 4168 25563 4200 25595
rect 4240 25563 4272 25595
rect 4312 25563 4344 25595
rect 4384 25563 4416 25595
rect 4456 25563 4488 25595
rect 4528 25563 4560 25595
rect 4600 25563 4632 25595
rect 4672 25563 4704 25595
rect 4744 25563 4776 25595
rect 4816 25563 4848 25595
rect 4888 25563 4920 25595
rect 4960 25563 4992 25595
rect 5032 25563 5064 25595
rect 5104 25563 5136 25595
rect 5176 25563 5208 25595
rect 5248 25563 5280 25595
rect 5320 25563 5352 25595
rect 5392 25563 5424 25595
rect 5464 25563 5496 25595
rect 5536 25563 5568 25595
rect 5608 25563 5640 25595
rect 5680 25563 5712 25595
rect 5752 25563 5784 25595
rect 5824 25563 5856 25595
rect 5896 25563 5928 25595
rect 5968 25563 6000 25595
rect 6040 25563 6072 25595
rect 6112 25563 6144 25595
rect 6184 25563 6216 25595
rect 6256 25563 6288 25595
rect 6328 25563 6360 25595
rect 6400 25563 6432 25595
rect 6472 25563 6504 25595
rect 6544 25563 6576 25595
rect 6616 25563 6648 25595
rect 6688 25563 6720 25595
rect 6760 25563 6792 25595
rect 6832 25563 6864 25595
rect 6904 25563 6936 25595
rect 6976 25563 7008 25595
rect 7048 25563 7080 25595
rect 7120 25563 7152 25595
rect 7192 25563 7224 25595
rect 7264 25563 7296 25595
rect 7336 25563 7368 25595
rect 7408 25563 7440 25595
rect 7480 25563 7512 25595
rect 7552 25563 7584 25595
rect 7624 25563 7656 25595
rect 7696 25563 7728 25595
rect 7768 25563 7800 25595
rect 7840 25563 7872 25595
rect 7912 25563 7944 25595
rect 7984 25563 8016 25595
rect 8056 25563 8088 25595
rect 8128 25563 8160 25595
rect 8200 25563 8232 25595
rect 8272 25563 8304 25595
rect 8344 25563 8376 25595
rect 8416 25563 8448 25595
rect 8488 25563 8520 25595
rect 8560 25563 8592 25595
rect 8632 25563 8664 25595
rect 8704 25563 8736 25595
rect 8776 25563 8808 25595
rect 8848 25563 8880 25595
rect 8920 25563 8952 25595
rect 8992 25563 9024 25595
rect 9064 25563 9096 25595
rect 9136 25563 9168 25595
rect 9208 25563 9240 25595
rect 9280 25563 9312 25595
rect 9352 25563 9384 25595
rect 9424 25563 9456 25595
rect 9496 25563 9528 25595
rect 9568 25563 9600 25595
rect 9640 25563 9672 25595
rect 9712 25563 9744 25595
rect 9784 25563 9816 25595
rect 9856 25563 9888 25595
rect 9928 25563 9960 25595
rect 10000 25563 10032 25595
rect 10072 25563 10104 25595
rect 10144 25563 10176 25595
rect 10216 25563 10248 25595
rect 10288 25563 10320 25595
rect 10360 25563 10392 25595
rect 10432 25563 10464 25595
rect 10504 25563 10536 25595
rect 10576 25563 10608 25595
rect 10648 25563 10680 25595
rect 10720 25563 10752 25595
rect 10792 25563 10824 25595
rect 10864 25563 10896 25595
rect 10936 25563 10968 25595
rect 11008 25563 11040 25595
rect 11080 25563 11112 25595
rect 11152 25563 11184 25595
rect 11224 25563 11256 25595
rect 11296 25563 11328 25595
rect 11368 25563 11400 25595
rect 11440 25563 11472 25595
rect 11512 25563 11544 25595
rect 11584 25563 11616 25595
rect 11656 25563 11688 25595
rect 11728 25563 11760 25595
rect 11800 25563 11832 25595
rect 11872 25563 11904 25595
rect 11944 25563 11976 25595
rect 12016 25563 12048 25595
rect 12088 25563 12120 25595
rect 12160 25563 12192 25595
rect 12232 25563 12264 25595
rect 12304 25563 12336 25595
rect 12376 25563 12408 25595
rect 12448 25563 12480 25595
rect 12520 25563 12552 25595
rect 12592 25563 12624 25595
rect 12664 25563 12696 25595
rect 12736 25563 12768 25595
rect 12808 25563 12840 25595
rect 12880 25563 12912 25595
rect 12952 25563 12984 25595
rect 13024 25563 13056 25595
rect 13096 25563 13128 25595
rect 13168 25563 13200 25595
rect 13240 25563 13272 25595
rect 13312 25563 13344 25595
rect 13384 25563 13416 25595
rect 13456 25563 13488 25595
rect 13528 25563 13560 25595
rect 13600 25563 13632 25595
rect 13672 25563 13704 25595
rect 13744 25563 13776 25595
rect 13816 25563 13848 25595
rect 13888 25563 13920 25595
rect 13960 25563 13992 25595
rect 14032 25563 14064 25595
rect 14104 25563 14136 25595
rect 14176 25563 14208 25595
rect 14248 25563 14280 25595
rect 14320 25563 14352 25595
rect 14392 25563 14424 25595
rect 14464 25563 14496 25595
rect 14536 25563 14568 25595
rect 14608 25563 14640 25595
rect 14680 25563 14712 25595
rect 14752 25563 14784 25595
rect 14824 25563 14856 25595
rect 14896 25563 14928 25595
rect 14968 25563 15000 25595
rect 15040 25563 15072 25595
rect 15112 25563 15144 25595
rect 15184 25563 15216 25595
rect 15256 25563 15288 25595
rect 15328 25563 15360 25595
rect 15400 25563 15432 25595
rect 15472 25563 15504 25595
rect 15544 25563 15576 25595
rect 15616 25563 15648 25595
rect 15688 25563 15720 25595
rect 15760 25563 15792 25595
rect 15832 25563 15864 25595
rect 15904 25563 15936 25595
rect 64 25491 96 25523
rect 136 25491 168 25523
rect 208 25491 240 25523
rect 280 25491 312 25523
rect 352 25491 384 25523
rect 424 25491 456 25523
rect 496 25491 528 25523
rect 568 25491 600 25523
rect 640 25491 672 25523
rect 712 25491 744 25523
rect 784 25491 816 25523
rect 856 25491 888 25523
rect 928 25491 960 25523
rect 1000 25491 1032 25523
rect 1072 25491 1104 25523
rect 1144 25491 1176 25523
rect 1216 25491 1248 25523
rect 1288 25491 1320 25523
rect 1360 25491 1392 25523
rect 1432 25491 1464 25523
rect 1504 25491 1536 25523
rect 1576 25491 1608 25523
rect 1648 25491 1680 25523
rect 1720 25491 1752 25523
rect 1792 25491 1824 25523
rect 1864 25491 1896 25523
rect 1936 25491 1968 25523
rect 2008 25491 2040 25523
rect 2080 25491 2112 25523
rect 2152 25491 2184 25523
rect 2224 25491 2256 25523
rect 2296 25491 2328 25523
rect 2368 25491 2400 25523
rect 2440 25491 2472 25523
rect 2512 25491 2544 25523
rect 2584 25491 2616 25523
rect 2656 25491 2688 25523
rect 2728 25491 2760 25523
rect 2800 25491 2832 25523
rect 2872 25491 2904 25523
rect 2944 25491 2976 25523
rect 3016 25491 3048 25523
rect 3088 25491 3120 25523
rect 3160 25491 3192 25523
rect 3232 25491 3264 25523
rect 3304 25491 3336 25523
rect 3376 25491 3408 25523
rect 3448 25491 3480 25523
rect 3520 25491 3552 25523
rect 3592 25491 3624 25523
rect 3664 25491 3696 25523
rect 3736 25491 3768 25523
rect 3808 25491 3840 25523
rect 3880 25491 3912 25523
rect 3952 25491 3984 25523
rect 4024 25491 4056 25523
rect 4096 25491 4128 25523
rect 4168 25491 4200 25523
rect 4240 25491 4272 25523
rect 4312 25491 4344 25523
rect 4384 25491 4416 25523
rect 4456 25491 4488 25523
rect 4528 25491 4560 25523
rect 4600 25491 4632 25523
rect 4672 25491 4704 25523
rect 4744 25491 4776 25523
rect 4816 25491 4848 25523
rect 4888 25491 4920 25523
rect 4960 25491 4992 25523
rect 5032 25491 5064 25523
rect 5104 25491 5136 25523
rect 5176 25491 5208 25523
rect 5248 25491 5280 25523
rect 5320 25491 5352 25523
rect 5392 25491 5424 25523
rect 5464 25491 5496 25523
rect 5536 25491 5568 25523
rect 5608 25491 5640 25523
rect 5680 25491 5712 25523
rect 5752 25491 5784 25523
rect 5824 25491 5856 25523
rect 5896 25491 5928 25523
rect 5968 25491 6000 25523
rect 6040 25491 6072 25523
rect 6112 25491 6144 25523
rect 6184 25491 6216 25523
rect 6256 25491 6288 25523
rect 6328 25491 6360 25523
rect 6400 25491 6432 25523
rect 6472 25491 6504 25523
rect 6544 25491 6576 25523
rect 6616 25491 6648 25523
rect 6688 25491 6720 25523
rect 6760 25491 6792 25523
rect 6832 25491 6864 25523
rect 6904 25491 6936 25523
rect 6976 25491 7008 25523
rect 7048 25491 7080 25523
rect 7120 25491 7152 25523
rect 7192 25491 7224 25523
rect 7264 25491 7296 25523
rect 7336 25491 7368 25523
rect 7408 25491 7440 25523
rect 7480 25491 7512 25523
rect 7552 25491 7584 25523
rect 7624 25491 7656 25523
rect 7696 25491 7728 25523
rect 7768 25491 7800 25523
rect 7840 25491 7872 25523
rect 7912 25491 7944 25523
rect 7984 25491 8016 25523
rect 8056 25491 8088 25523
rect 8128 25491 8160 25523
rect 8200 25491 8232 25523
rect 8272 25491 8304 25523
rect 8344 25491 8376 25523
rect 8416 25491 8448 25523
rect 8488 25491 8520 25523
rect 8560 25491 8592 25523
rect 8632 25491 8664 25523
rect 8704 25491 8736 25523
rect 8776 25491 8808 25523
rect 8848 25491 8880 25523
rect 8920 25491 8952 25523
rect 8992 25491 9024 25523
rect 9064 25491 9096 25523
rect 9136 25491 9168 25523
rect 9208 25491 9240 25523
rect 9280 25491 9312 25523
rect 9352 25491 9384 25523
rect 9424 25491 9456 25523
rect 9496 25491 9528 25523
rect 9568 25491 9600 25523
rect 9640 25491 9672 25523
rect 9712 25491 9744 25523
rect 9784 25491 9816 25523
rect 9856 25491 9888 25523
rect 9928 25491 9960 25523
rect 10000 25491 10032 25523
rect 10072 25491 10104 25523
rect 10144 25491 10176 25523
rect 10216 25491 10248 25523
rect 10288 25491 10320 25523
rect 10360 25491 10392 25523
rect 10432 25491 10464 25523
rect 10504 25491 10536 25523
rect 10576 25491 10608 25523
rect 10648 25491 10680 25523
rect 10720 25491 10752 25523
rect 10792 25491 10824 25523
rect 10864 25491 10896 25523
rect 10936 25491 10968 25523
rect 11008 25491 11040 25523
rect 11080 25491 11112 25523
rect 11152 25491 11184 25523
rect 11224 25491 11256 25523
rect 11296 25491 11328 25523
rect 11368 25491 11400 25523
rect 11440 25491 11472 25523
rect 11512 25491 11544 25523
rect 11584 25491 11616 25523
rect 11656 25491 11688 25523
rect 11728 25491 11760 25523
rect 11800 25491 11832 25523
rect 11872 25491 11904 25523
rect 11944 25491 11976 25523
rect 12016 25491 12048 25523
rect 12088 25491 12120 25523
rect 12160 25491 12192 25523
rect 12232 25491 12264 25523
rect 12304 25491 12336 25523
rect 12376 25491 12408 25523
rect 12448 25491 12480 25523
rect 12520 25491 12552 25523
rect 12592 25491 12624 25523
rect 12664 25491 12696 25523
rect 12736 25491 12768 25523
rect 12808 25491 12840 25523
rect 12880 25491 12912 25523
rect 12952 25491 12984 25523
rect 13024 25491 13056 25523
rect 13096 25491 13128 25523
rect 13168 25491 13200 25523
rect 13240 25491 13272 25523
rect 13312 25491 13344 25523
rect 13384 25491 13416 25523
rect 13456 25491 13488 25523
rect 13528 25491 13560 25523
rect 13600 25491 13632 25523
rect 13672 25491 13704 25523
rect 13744 25491 13776 25523
rect 13816 25491 13848 25523
rect 13888 25491 13920 25523
rect 13960 25491 13992 25523
rect 14032 25491 14064 25523
rect 14104 25491 14136 25523
rect 14176 25491 14208 25523
rect 14248 25491 14280 25523
rect 14320 25491 14352 25523
rect 14392 25491 14424 25523
rect 14464 25491 14496 25523
rect 14536 25491 14568 25523
rect 14608 25491 14640 25523
rect 14680 25491 14712 25523
rect 14752 25491 14784 25523
rect 14824 25491 14856 25523
rect 14896 25491 14928 25523
rect 14968 25491 15000 25523
rect 15040 25491 15072 25523
rect 15112 25491 15144 25523
rect 15184 25491 15216 25523
rect 15256 25491 15288 25523
rect 15328 25491 15360 25523
rect 15400 25491 15432 25523
rect 15472 25491 15504 25523
rect 15544 25491 15576 25523
rect 15616 25491 15648 25523
rect 15688 25491 15720 25523
rect 15760 25491 15792 25523
rect 15832 25491 15864 25523
rect 15904 25491 15936 25523
rect 64 25419 96 25451
rect 136 25419 168 25451
rect 208 25419 240 25451
rect 280 25419 312 25451
rect 352 25419 384 25451
rect 424 25419 456 25451
rect 496 25419 528 25451
rect 568 25419 600 25451
rect 640 25419 672 25451
rect 712 25419 744 25451
rect 784 25419 816 25451
rect 856 25419 888 25451
rect 928 25419 960 25451
rect 1000 25419 1032 25451
rect 1072 25419 1104 25451
rect 1144 25419 1176 25451
rect 1216 25419 1248 25451
rect 1288 25419 1320 25451
rect 1360 25419 1392 25451
rect 1432 25419 1464 25451
rect 1504 25419 1536 25451
rect 1576 25419 1608 25451
rect 1648 25419 1680 25451
rect 1720 25419 1752 25451
rect 1792 25419 1824 25451
rect 1864 25419 1896 25451
rect 1936 25419 1968 25451
rect 2008 25419 2040 25451
rect 2080 25419 2112 25451
rect 2152 25419 2184 25451
rect 2224 25419 2256 25451
rect 2296 25419 2328 25451
rect 2368 25419 2400 25451
rect 2440 25419 2472 25451
rect 2512 25419 2544 25451
rect 2584 25419 2616 25451
rect 2656 25419 2688 25451
rect 2728 25419 2760 25451
rect 2800 25419 2832 25451
rect 2872 25419 2904 25451
rect 2944 25419 2976 25451
rect 3016 25419 3048 25451
rect 3088 25419 3120 25451
rect 3160 25419 3192 25451
rect 3232 25419 3264 25451
rect 3304 25419 3336 25451
rect 3376 25419 3408 25451
rect 3448 25419 3480 25451
rect 3520 25419 3552 25451
rect 3592 25419 3624 25451
rect 3664 25419 3696 25451
rect 3736 25419 3768 25451
rect 3808 25419 3840 25451
rect 3880 25419 3912 25451
rect 3952 25419 3984 25451
rect 4024 25419 4056 25451
rect 4096 25419 4128 25451
rect 4168 25419 4200 25451
rect 4240 25419 4272 25451
rect 4312 25419 4344 25451
rect 4384 25419 4416 25451
rect 4456 25419 4488 25451
rect 4528 25419 4560 25451
rect 4600 25419 4632 25451
rect 4672 25419 4704 25451
rect 4744 25419 4776 25451
rect 4816 25419 4848 25451
rect 4888 25419 4920 25451
rect 4960 25419 4992 25451
rect 5032 25419 5064 25451
rect 5104 25419 5136 25451
rect 5176 25419 5208 25451
rect 5248 25419 5280 25451
rect 5320 25419 5352 25451
rect 5392 25419 5424 25451
rect 5464 25419 5496 25451
rect 5536 25419 5568 25451
rect 5608 25419 5640 25451
rect 5680 25419 5712 25451
rect 5752 25419 5784 25451
rect 5824 25419 5856 25451
rect 5896 25419 5928 25451
rect 5968 25419 6000 25451
rect 6040 25419 6072 25451
rect 6112 25419 6144 25451
rect 6184 25419 6216 25451
rect 6256 25419 6288 25451
rect 6328 25419 6360 25451
rect 6400 25419 6432 25451
rect 6472 25419 6504 25451
rect 6544 25419 6576 25451
rect 6616 25419 6648 25451
rect 6688 25419 6720 25451
rect 6760 25419 6792 25451
rect 6832 25419 6864 25451
rect 6904 25419 6936 25451
rect 6976 25419 7008 25451
rect 7048 25419 7080 25451
rect 7120 25419 7152 25451
rect 7192 25419 7224 25451
rect 7264 25419 7296 25451
rect 7336 25419 7368 25451
rect 7408 25419 7440 25451
rect 7480 25419 7512 25451
rect 7552 25419 7584 25451
rect 7624 25419 7656 25451
rect 7696 25419 7728 25451
rect 7768 25419 7800 25451
rect 7840 25419 7872 25451
rect 7912 25419 7944 25451
rect 7984 25419 8016 25451
rect 8056 25419 8088 25451
rect 8128 25419 8160 25451
rect 8200 25419 8232 25451
rect 8272 25419 8304 25451
rect 8344 25419 8376 25451
rect 8416 25419 8448 25451
rect 8488 25419 8520 25451
rect 8560 25419 8592 25451
rect 8632 25419 8664 25451
rect 8704 25419 8736 25451
rect 8776 25419 8808 25451
rect 8848 25419 8880 25451
rect 8920 25419 8952 25451
rect 8992 25419 9024 25451
rect 9064 25419 9096 25451
rect 9136 25419 9168 25451
rect 9208 25419 9240 25451
rect 9280 25419 9312 25451
rect 9352 25419 9384 25451
rect 9424 25419 9456 25451
rect 9496 25419 9528 25451
rect 9568 25419 9600 25451
rect 9640 25419 9672 25451
rect 9712 25419 9744 25451
rect 9784 25419 9816 25451
rect 9856 25419 9888 25451
rect 9928 25419 9960 25451
rect 10000 25419 10032 25451
rect 10072 25419 10104 25451
rect 10144 25419 10176 25451
rect 10216 25419 10248 25451
rect 10288 25419 10320 25451
rect 10360 25419 10392 25451
rect 10432 25419 10464 25451
rect 10504 25419 10536 25451
rect 10576 25419 10608 25451
rect 10648 25419 10680 25451
rect 10720 25419 10752 25451
rect 10792 25419 10824 25451
rect 10864 25419 10896 25451
rect 10936 25419 10968 25451
rect 11008 25419 11040 25451
rect 11080 25419 11112 25451
rect 11152 25419 11184 25451
rect 11224 25419 11256 25451
rect 11296 25419 11328 25451
rect 11368 25419 11400 25451
rect 11440 25419 11472 25451
rect 11512 25419 11544 25451
rect 11584 25419 11616 25451
rect 11656 25419 11688 25451
rect 11728 25419 11760 25451
rect 11800 25419 11832 25451
rect 11872 25419 11904 25451
rect 11944 25419 11976 25451
rect 12016 25419 12048 25451
rect 12088 25419 12120 25451
rect 12160 25419 12192 25451
rect 12232 25419 12264 25451
rect 12304 25419 12336 25451
rect 12376 25419 12408 25451
rect 12448 25419 12480 25451
rect 12520 25419 12552 25451
rect 12592 25419 12624 25451
rect 12664 25419 12696 25451
rect 12736 25419 12768 25451
rect 12808 25419 12840 25451
rect 12880 25419 12912 25451
rect 12952 25419 12984 25451
rect 13024 25419 13056 25451
rect 13096 25419 13128 25451
rect 13168 25419 13200 25451
rect 13240 25419 13272 25451
rect 13312 25419 13344 25451
rect 13384 25419 13416 25451
rect 13456 25419 13488 25451
rect 13528 25419 13560 25451
rect 13600 25419 13632 25451
rect 13672 25419 13704 25451
rect 13744 25419 13776 25451
rect 13816 25419 13848 25451
rect 13888 25419 13920 25451
rect 13960 25419 13992 25451
rect 14032 25419 14064 25451
rect 14104 25419 14136 25451
rect 14176 25419 14208 25451
rect 14248 25419 14280 25451
rect 14320 25419 14352 25451
rect 14392 25419 14424 25451
rect 14464 25419 14496 25451
rect 14536 25419 14568 25451
rect 14608 25419 14640 25451
rect 14680 25419 14712 25451
rect 14752 25419 14784 25451
rect 14824 25419 14856 25451
rect 14896 25419 14928 25451
rect 14968 25419 15000 25451
rect 15040 25419 15072 25451
rect 15112 25419 15144 25451
rect 15184 25419 15216 25451
rect 15256 25419 15288 25451
rect 15328 25419 15360 25451
rect 15400 25419 15432 25451
rect 15472 25419 15504 25451
rect 15544 25419 15576 25451
rect 15616 25419 15648 25451
rect 15688 25419 15720 25451
rect 15760 25419 15792 25451
rect 15832 25419 15864 25451
rect 15904 25419 15936 25451
rect 64 25347 96 25379
rect 136 25347 168 25379
rect 208 25347 240 25379
rect 280 25347 312 25379
rect 352 25347 384 25379
rect 424 25347 456 25379
rect 496 25347 528 25379
rect 568 25347 600 25379
rect 640 25347 672 25379
rect 712 25347 744 25379
rect 784 25347 816 25379
rect 856 25347 888 25379
rect 928 25347 960 25379
rect 1000 25347 1032 25379
rect 1072 25347 1104 25379
rect 1144 25347 1176 25379
rect 1216 25347 1248 25379
rect 1288 25347 1320 25379
rect 1360 25347 1392 25379
rect 1432 25347 1464 25379
rect 1504 25347 1536 25379
rect 1576 25347 1608 25379
rect 1648 25347 1680 25379
rect 1720 25347 1752 25379
rect 1792 25347 1824 25379
rect 1864 25347 1896 25379
rect 1936 25347 1968 25379
rect 2008 25347 2040 25379
rect 2080 25347 2112 25379
rect 2152 25347 2184 25379
rect 2224 25347 2256 25379
rect 2296 25347 2328 25379
rect 2368 25347 2400 25379
rect 2440 25347 2472 25379
rect 2512 25347 2544 25379
rect 2584 25347 2616 25379
rect 2656 25347 2688 25379
rect 2728 25347 2760 25379
rect 2800 25347 2832 25379
rect 2872 25347 2904 25379
rect 2944 25347 2976 25379
rect 3016 25347 3048 25379
rect 3088 25347 3120 25379
rect 3160 25347 3192 25379
rect 3232 25347 3264 25379
rect 3304 25347 3336 25379
rect 3376 25347 3408 25379
rect 3448 25347 3480 25379
rect 3520 25347 3552 25379
rect 3592 25347 3624 25379
rect 3664 25347 3696 25379
rect 3736 25347 3768 25379
rect 3808 25347 3840 25379
rect 3880 25347 3912 25379
rect 3952 25347 3984 25379
rect 4024 25347 4056 25379
rect 4096 25347 4128 25379
rect 4168 25347 4200 25379
rect 4240 25347 4272 25379
rect 4312 25347 4344 25379
rect 4384 25347 4416 25379
rect 4456 25347 4488 25379
rect 4528 25347 4560 25379
rect 4600 25347 4632 25379
rect 4672 25347 4704 25379
rect 4744 25347 4776 25379
rect 4816 25347 4848 25379
rect 4888 25347 4920 25379
rect 4960 25347 4992 25379
rect 5032 25347 5064 25379
rect 5104 25347 5136 25379
rect 5176 25347 5208 25379
rect 5248 25347 5280 25379
rect 5320 25347 5352 25379
rect 5392 25347 5424 25379
rect 5464 25347 5496 25379
rect 5536 25347 5568 25379
rect 5608 25347 5640 25379
rect 5680 25347 5712 25379
rect 5752 25347 5784 25379
rect 5824 25347 5856 25379
rect 5896 25347 5928 25379
rect 5968 25347 6000 25379
rect 6040 25347 6072 25379
rect 6112 25347 6144 25379
rect 6184 25347 6216 25379
rect 6256 25347 6288 25379
rect 6328 25347 6360 25379
rect 6400 25347 6432 25379
rect 6472 25347 6504 25379
rect 6544 25347 6576 25379
rect 6616 25347 6648 25379
rect 6688 25347 6720 25379
rect 6760 25347 6792 25379
rect 6832 25347 6864 25379
rect 6904 25347 6936 25379
rect 6976 25347 7008 25379
rect 7048 25347 7080 25379
rect 7120 25347 7152 25379
rect 7192 25347 7224 25379
rect 7264 25347 7296 25379
rect 7336 25347 7368 25379
rect 7408 25347 7440 25379
rect 7480 25347 7512 25379
rect 7552 25347 7584 25379
rect 7624 25347 7656 25379
rect 7696 25347 7728 25379
rect 7768 25347 7800 25379
rect 7840 25347 7872 25379
rect 7912 25347 7944 25379
rect 7984 25347 8016 25379
rect 8056 25347 8088 25379
rect 8128 25347 8160 25379
rect 8200 25347 8232 25379
rect 8272 25347 8304 25379
rect 8344 25347 8376 25379
rect 8416 25347 8448 25379
rect 8488 25347 8520 25379
rect 8560 25347 8592 25379
rect 8632 25347 8664 25379
rect 8704 25347 8736 25379
rect 8776 25347 8808 25379
rect 8848 25347 8880 25379
rect 8920 25347 8952 25379
rect 8992 25347 9024 25379
rect 9064 25347 9096 25379
rect 9136 25347 9168 25379
rect 9208 25347 9240 25379
rect 9280 25347 9312 25379
rect 9352 25347 9384 25379
rect 9424 25347 9456 25379
rect 9496 25347 9528 25379
rect 9568 25347 9600 25379
rect 9640 25347 9672 25379
rect 9712 25347 9744 25379
rect 9784 25347 9816 25379
rect 9856 25347 9888 25379
rect 9928 25347 9960 25379
rect 10000 25347 10032 25379
rect 10072 25347 10104 25379
rect 10144 25347 10176 25379
rect 10216 25347 10248 25379
rect 10288 25347 10320 25379
rect 10360 25347 10392 25379
rect 10432 25347 10464 25379
rect 10504 25347 10536 25379
rect 10576 25347 10608 25379
rect 10648 25347 10680 25379
rect 10720 25347 10752 25379
rect 10792 25347 10824 25379
rect 10864 25347 10896 25379
rect 10936 25347 10968 25379
rect 11008 25347 11040 25379
rect 11080 25347 11112 25379
rect 11152 25347 11184 25379
rect 11224 25347 11256 25379
rect 11296 25347 11328 25379
rect 11368 25347 11400 25379
rect 11440 25347 11472 25379
rect 11512 25347 11544 25379
rect 11584 25347 11616 25379
rect 11656 25347 11688 25379
rect 11728 25347 11760 25379
rect 11800 25347 11832 25379
rect 11872 25347 11904 25379
rect 11944 25347 11976 25379
rect 12016 25347 12048 25379
rect 12088 25347 12120 25379
rect 12160 25347 12192 25379
rect 12232 25347 12264 25379
rect 12304 25347 12336 25379
rect 12376 25347 12408 25379
rect 12448 25347 12480 25379
rect 12520 25347 12552 25379
rect 12592 25347 12624 25379
rect 12664 25347 12696 25379
rect 12736 25347 12768 25379
rect 12808 25347 12840 25379
rect 12880 25347 12912 25379
rect 12952 25347 12984 25379
rect 13024 25347 13056 25379
rect 13096 25347 13128 25379
rect 13168 25347 13200 25379
rect 13240 25347 13272 25379
rect 13312 25347 13344 25379
rect 13384 25347 13416 25379
rect 13456 25347 13488 25379
rect 13528 25347 13560 25379
rect 13600 25347 13632 25379
rect 13672 25347 13704 25379
rect 13744 25347 13776 25379
rect 13816 25347 13848 25379
rect 13888 25347 13920 25379
rect 13960 25347 13992 25379
rect 14032 25347 14064 25379
rect 14104 25347 14136 25379
rect 14176 25347 14208 25379
rect 14248 25347 14280 25379
rect 14320 25347 14352 25379
rect 14392 25347 14424 25379
rect 14464 25347 14496 25379
rect 14536 25347 14568 25379
rect 14608 25347 14640 25379
rect 14680 25347 14712 25379
rect 14752 25347 14784 25379
rect 14824 25347 14856 25379
rect 14896 25347 14928 25379
rect 14968 25347 15000 25379
rect 15040 25347 15072 25379
rect 15112 25347 15144 25379
rect 15184 25347 15216 25379
rect 15256 25347 15288 25379
rect 15328 25347 15360 25379
rect 15400 25347 15432 25379
rect 15472 25347 15504 25379
rect 15544 25347 15576 25379
rect 15616 25347 15648 25379
rect 15688 25347 15720 25379
rect 15760 25347 15792 25379
rect 15832 25347 15864 25379
rect 15904 25347 15936 25379
rect 64 25275 96 25307
rect 136 25275 168 25307
rect 208 25275 240 25307
rect 280 25275 312 25307
rect 352 25275 384 25307
rect 424 25275 456 25307
rect 496 25275 528 25307
rect 568 25275 600 25307
rect 640 25275 672 25307
rect 712 25275 744 25307
rect 784 25275 816 25307
rect 856 25275 888 25307
rect 928 25275 960 25307
rect 1000 25275 1032 25307
rect 1072 25275 1104 25307
rect 1144 25275 1176 25307
rect 1216 25275 1248 25307
rect 1288 25275 1320 25307
rect 1360 25275 1392 25307
rect 1432 25275 1464 25307
rect 1504 25275 1536 25307
rect 1576 25275 1608 25307
rect 1648 25275 1680 25307
rect 1720 25275 1752 25307
rect 1792 25275 1824 25307
rect 1864 25275 1896 25307
rect 1936 25275 1968 25307
rect 2008 25275 2040 25307
rect 2080 25275 2112 25307
rect 2152 25275 2184 25307
rect 2224 25275 2256 25307
rect 2296 25275 2328 25307
rect 2368 25275 2400 25307
rect 2440 25275 2472 25307
rect 2512 25275 2544 25307
rect 2584 25275 2616 25307
rect 2656 25275 2688 25307
rect 2728 25275 2760 25307
rect 2800 25275 2832 25307
rect 2872 25275 2904 25307
rect 2944 25275 2976 25307
rect 3016 25275 3048 25307
rect 3088 25275 3120 25307
rect 3160 25275 3192 25307
rect 3232 25275 3264 25307
rect 3304 25275 3336 25307
rect 3376 25275 3408 25307
rect 3448 25275 3480 25307
rect 3520 25275 3552 25307
rect 3592 25275 3624 25307
rect 3664 25275 3696 25307
rect 3736 25275 3768 25307
rect 3808 25275 3840 25307
rect 3880 25275 3912 25307
rect 3952 25275 3984 25307
rect 4024 25275 4056 25307
rect 4096 25275 4128 25307
rect 4168 25275 4200 25307
rect 4240 25275 4272 25307
rect 4312 25275 4344 25307
rect 4384 25275 4416 25307
rect 4456 25275 4488 25307
rect 4528 25275 4560 25307
rect 4600 25275 4632 25307
rect 4672 25275 4704 25307
rect 4744 25275 4776 25307
rect 4816 25275 4848 25307
rect 4888 25275 4920 25307
rect 4960 25275 4992 25307
rect 5032 25275 5064 25307
rect 5104 25275 5136 25307
rect 5176 25275 5208 25307
rect 5248 25275 5280 25307
rect 5320 25275 5352 25307
rect 5392 25275 5424 25307
rect 5464 25275 5496 25307
rect 5536 25275 5568 25307
rect 5608 25275 5640 25307
rect 5680 25275 5712 25307
rect 5752 25275 5784 25307
rect 5824 25275 5856 25307
rect 5896 25275 5928 25307
rect 5968 25275 6000 25307
rect 6040 25275 6072 25307
rect 6112 25275 6144 25307
rect 6184 25275 6216 25307
rect 6256 25275 6288 25307
rect 6328 25275 6360 25307
rect 6400 25275 6432 25307
rect 6472 25275 6504 25307
rect 6544 25275 6576 25307
rect 6616 25275 6648 25307
rect 6688 25275 6720 25307
rect 6760 25275 6792 25307
rect 6832 25275 6864 25307
rect 6904 25275 6936 25307
rect 6976 25275 7008 25307
rect 7048 25275 7080 25307
rect 7120 25275 7152 25307
rect 7192 25275 7224 25307
rect 7264 25275 7296 25307
rect 7336 25275 7368 25307
rect 7408 25275 7440 25307
rect 7480 25275 7512 25307
rect 7552 25275 7584 25307
rect 7624 25275 7656 25307
rect 7696 25275 7728 25307
rect 7768 25275 7800 25307
rect 7840 25275 7872 25307
rect 7912 25275 7944 25307
rect 7984 25275 8016 25307
rect 8056 25275 8088 25307
rect 8128 25275 8160 25307
rect 8200 25275 8232 25307
rect 8272 25275 8304 25307
rect 8344 25275 8376 25307
rect 8416 25275 8448 25307
rect 8488 25275 8520 25307
rect 8560 25275 8592 25307
rect 8632 25275 8664 25307
rect 8704 25275 8736 25307
rect 8776 25275 8808 25307
rect 8848 25275 8880 25307
rect 8920 25275 8952 25307
rect 8992 25275 9024 25307
rect 9064 25275 9096 25307
rect 9136 25275 9168 25307
rect 9208 25275 9240 25307
rect 9280 25275 9312 25307
rect 9352 25275 9384 25307
rect 9424 25275 9456 25307
rect 9496 25275 9528 25307
rect 9568 25275 9600 25307
rect 9640 25275 9672 25307
rect 9712 25275 9744 25307
rect 9784 25275 9816 25307
rect 9856 25275 9888 25307
rect 9928 25275 9960 25307
rect 10000 25275 10032 25307
rect 10072 25275 10104 25307
rect 10144 25275 10176 25307
rect 10216 25275 10248 25307
rect 10288 25275 10320 25307
rect 10360 25275 10392 25307
rect 10432 25275 10464 25307
rect 10504 25275 10536 25307
rect 10576 25275 10608 25307
rect 10648 25275 10680 25307
rect 10720 25275 10752 25307
rect 10792 25275 10824 25307
rect 10864 25275 10896 25307
rect 10936 25275 10968 25307
rect 11008 25275 11040 25307
rect 11080 25275 11112 25307
rect 11152 25275 11184 25307
rect 11224 25275 11256 25307
rect 11296 25275 11328 25307
rect 11368 25275 11400 25307
rect 11440 25275 11472 25307
rect 11512 25275 11544 25307
rect 11584 25275 11616 25307
rect 11656 25275 11688 25307
rect 11728 25275 11760 25307
rect 11800 25275 11832 25307
rect 11872 25275 11904 25307
rect 11944 25275 11976 25307
rect 12016 25275 12048 25307
rect 12088 25275 12120 25307
rect 12160 25275 12192 25307
rect 12232 25275 12264 25307
rect 12304 25275 12336 25307
rect 12376 25275 12408 25307
rect 12448 25275 12480 25307
rect 12520 25275 12552 25307
rect 12592 25275 12624 25307
rect 12664 25275 12696 25307
rect 12736 25275 12768 25307
rect 12808 25275 12840 25307
rect 12880 25275 12912 25307
rect 12952 25275 12984 25307
rect 13024 25275 13056 25307
rect 13096 25275 13128 25307
rect 13168 25275 13200 25307
rect 13240 25275 13272 25307
rect 13312 25275 13344 25307
rect 13384 25275 13416 25307
rect 13456 25275 13488 25307
rect 13528 25275 13560 25307
rect 13600 25275 13632 25307
rect 13672 25275 13704 25307
rect 13744 25275 13776 25307
rect 13816 25275 13848 25307
rect 13888 25275 13920 25307
rect 13960 25275 13992 25307
rect 14032 25275 14064 25307
rect 14104 25275 14136 25307
rect 14176 25275 14208 25307
rect 14248 25275 14280 25307
rect 14320 25275 14352 25307
rect 14392 25275 14424 25307
rect 14464 25275 14496 25307
rect 14536 25275 14568 25307
rect 14608 25275 14640 25307
rect 14680 25275 14712 25307
rect 14752 25275 14784 25307
rect 14824 25275 14856 25307
rect 14896 25275 14928 25307
rect 14968 25275 15000 25307
rect 15040 25275 15072 25307
rect 15112 25275 15144 25307
rect 15184 25275 15216 25307
rect 15256 25275 15288 25307
rect 15328 25275 15360 25307
rect 15400 25275 15432 25307
rect 15472 25275 15504 25307
rect 15544 25275 15576 25307
rect 15616 25275 15648 25307
rect 15688 25275 15720 25307
rect 15760 25275 15792 25307
rect 15832 25275 15864 25307
rect 15904 25275 15936 25307
rect 64 25203 96 25235
rect 136 25203 168 25235
rect 208 25203 240 25235
rect 280 25203 312 25235
rect 352 25203 384 25235
rect 424 25203 456 25235
rect 496 25203 528 25235
rect 568 25203 600 25235
rect 640 25203 672 25235
rect 712 25203 744 25235
rect 784 25203 816 25235
rect 856 25203 888 25235
rect 928 25203 960 25235
rect 1000 25203 1032 25235
rect 1072 25203 1104 25235
rect 1144 25203 1176 25235
rect 1216 25203 1248 25235
rect 1288 25203 1320 25235
rect 1360 25203 1392 25235
rect 1432 25203 1464 25235
rect 1504 25203 1536 25235
rect 1576 25203 1608 25235
rect 1648 25203 1680 25235
rect 1720 25203 1752 25235
rect 1792 25203 1824 25235
rect 1864 25203 1896 25235
rect 1936 25203 1968 25235
rect 2008 25203 2040 25235
rect 2080 25203 2112 25235
rect 2152 25203 2184 25235
rect 2224 25203 2256 25235
rect 2296 25203 2328 25235
rect 2368 25203 2400 25235
rect 2440 25203 2472 25235
rect 2512 25203 2544 25235
rect 2584 25203 2616 25235
rect 2656 25203 2688 25235
rect 2728 25203 2760 25235
rect 2800 25203 2832 25235
rect 2872 25203 2904 25235
rect 2944 25203 2976 25235
rect 3016 25203 3048 25235
rect 3088 25203 3120 25235
rect 3160 25203 3192 25235
rect 3232 25203 3264 25235
rect 3304 25203 3336 25235
rect 3376 25203 3408 25235
rect 3448 25203 3480 25235
rect 3520 25203 3552 25235
rect 3592 25203 3624 25235
rect 3664 25203 3696 25235
rect 3736 25203 3768 25235
rect 3808 25203 3840 25235
rect 3880 25203 3912 25235
rect 3952 25203 3984 25235
rect 4024 25203 4056 25235
rect 4096 25203 4128 25235
rect 4168 25203 4200 25235
rect 4240 25203 4272 25235
rect 4312 25203 4344 25235
rect 4384 25203 4416 25235
rect 4456 25203 4488 25235
rect 4528 25203 4560 25235
rect 4600 25203 4632 25235
rect 4672 25203 4704 25235
rect 4744 25203 4776 25235
rect 4816 25203 4848 25235
rect 4888 25203 4920 25235
rect 4960 25203 4992 25235
rect 5032 25203 5064 25235
rect 5104 25203 5136 25235
rect 5176 25203 5208 25235
rect 5248 25203 5280 25235
rect 5320 25203 5352 25235
rect 5392 25203 5424 25235
rect 5464 25203 5496 25235
rect 5536 25203 5568 25235
rect 5608 25203 5640 25235
rect 5680 25203 5712 25235
rect 5752 25203 5784 25235
rect 5824 25203 5856 25235
rect 5896 25203 5928 25235
rect 5968 25203 6000 25235
rect 6040 25203 6072 25235
rect 6112 25203 6144 25235
rect 6184 25203 6216 25235
rect 6256 25203 6288 25235
rect 6328 25203 6360 25235
rect 6400 25203 6432 25235
rect 6472 25203 6504 25235
rect 6544 25203 6576 25235
rect 6616 25203 6648 25235
rect 6688 25203 6720 25235
rect 6760 25203 6792 25235
rect 6832 25203 6864 25235
rect 6904 25203 6936 25235
rect 6976 25203 7008 25235
rect 7048 25203 7080 25235
rect 7120 25203 7152 25235
rect 7192 25203 7224 25235
rect 7264 25203 7296 25235
rect 7336 25203 7368 25235
rect 7408 25203 7440 25235
rect 7480 25203 7512 25235
rect 7552 25203 7584 25235
rect 7624 25203 7656 25235
rect 7696 25203 7728 25235
rect 7768 25203 7800 25235
rect 7840 25203 7872 25235
rect 7912 25203 7944 25235
rect 7984 25203 8016 25235
rect 8056 25203 8088 25235
rect 8128 25203 8160 25235
rect 8200 25203 8232 25235
rect 8272 25203 8304 25235
rect 8344 25203 8376 25235
rect 8416 25203 8448 25235
rect 8488 25203 8520 25235
rect 8560 25203 8592 25235
rect 8632 25203 8664 25235
rect 8704 25203 8736 25235
rect 8776 25203 8808 25235
rect 8848 25203 8880 25235
rect 8920 25203 8952 25235
rect 8992 25203 9024 25235
rect 9064 25203 9096 25235
rect 9136 25203 9168 25235
rect 9208 25203 9240 25235
rect 9280 25203 9312 25235
rect 9352 25203 9384 25235
rect 9424 25203 9456 25235
rect 9496 25203 9528 25235
rect 9568 25203 9600 25235
rect 9640 25203 9672 25235
rect 9712 25203 9744 25235
rect 9784 25203 9816 25235
rect 9856 25203 9888 25235
rect 9928 25203 9960 25235
rect 10000 25203 10032 25235
rect 10072 25203 10104 25235
rect 10144 25203 10176 25235
rect 10216 25203 10248 25235
rect 10288 25203 10320 25235
rect 10360 25203 10392 25235
rect 10432 25203 10464 25235
rect 10504 25203 10536 25235
rect 10576 25203 10608 25235
rect 10648 25203 10680 25235
rect 10720 25203 10752 25235
rect 10792 25203 10824 25235
rect 10864 25203 10896 25235
rect 10936 25203 10968 25235
rect 11008 25203 11040 25235
rect 11080 25203 11112 25235
rect 11152 25203 11184 25235
rect 11224 25203 11256 25235
rect 11296 25203 11328 25235
rect 11368 25203 11400 25235
rect 11440 25203 11472 25235
rect 11512 25203 11544 25235
rect 11584 25203 11616 25235
rect 11656 25203 11688 25235
rect 11728 25203 11760 25235
rect 11800 25203 11832 25235
rect 11872 25203 11904 25235
rect 11944 25203 11976 25235
rect 12016 25203 12048 25235
rect 12088 25203 12120 25235
rect 12160 25203 12192 25235
rect 12232 25203 12264 25235
rect 12304 25203 12336 25235
rect 12376 25203 12408 25235
rect 12448 25203 12480 25235
rect 12520 25203 12552 25235
rect 12592 25203 12624 25235
rect 12664 25203 12696 25235
rect 12736 25203 12768 25235
rect 12808 25203 12840 25235
rect 12880 25203 12912 25235
rect 12952 25203 12984 25235
rect 13024 25203 13056 25235
rect 13096 25203 13128 25235
rect 13168 25203 13200 25235
rect 13240 25203 13272 25235
rect 13312 25203 13344 25235
rect 13384 25203 13416 25235
rect 13456 25203 13488 25235
rect 13528 25203 13560 25235
rect 13600 25203 13632 25235
rect 13672 25203 13704 25235
rect 13744 25203 13776 25235
rect 13816 25203 13848 25235
rect 13888 25203 13920 25235
rect 13960 25203 13992 25235
rect 14032 25203 14064 25235
rect 14104 25203 14136 25235
rect 14176 25203 14208 25235
rect 14248 25203 14280 25235
rect 14320 25203 14352 25235
rect 14392 25203 14424 25235
rect 14464 25203 14496 25235
rect 14536 25203 14568 25235
rect 14608 25203 14640 25235
rect 14680 25203 14712 25235
rect 14752 25203 14784 25235
rect 14824 25203 14856 25235
rect 14896 25203 14928 25235
rect 14968 25203 15000 25235
rect 15040 25203 15072 25235
rect 15112 25203 15144 25235
rect 15184 25203 15216 25235
rect 15256 25203 15288 25235
rect 15328 25203 15360 25235
rect 15400 25203 15432 25235
rect 15472 25203 15504 25235
rect 15544 25203 15576 25235
rect 15616 25203 15648 25235
rect 15688 25203 15720 25235
rect 15760 25203 15792 25235
rect 15832 25203 15864 25235
rect 15904 25203 15936 25235
rect 64 25131 96 25163
rect 136 25131 168 25163
rect 208 25131 240 25163
rect 280 25131 312 25163
rect 352 25131 384 25163
rect 424 25131 456 25163
rect 496 25131 528 25163
rect 568 25131 600 25163
rect 640 25131 672 25163
rect 712 25131 744 25163
rect 784 25131 816 25163
rect 856 25131 888 25163
rect 928 25131 960 25163
rect 1000 25131 1032 25163
rect 1072 25131 1104 25163
rect 1144 25131 1176 25163
rect 1216 25131 1248 25163
rect 1288 25131 1320 25163
rect 1360 25131 1392 25163
rect 1432 25131 1464 25163
rect 1504 25131 1536 25163
rect 1576 25131 1608 25163
rect 1648 25131 1680 25163
rect 1720 25131 1752 25163
rect 1792 25131 1824 25163
rect 1864 25131 1896 25163
rect 1936 25131 1968 25163
rect 2008 25131 2040 25163
rect 2080 25131 2112 25163
rect 2152 25131 2184 25163
rect 2224 25131 2256 25163
rect 2296 25131 2328 25163
rect 2368 25131 2400 25163
rect 2440 25131 2472 25163
rect 2512 25131 2544 25163
rect 2584 25131 2616 25163
rect 2656 25131 2688 25163
rect 2728 25131 2760 25163
rect 2800 25131 2832 25163
rect 2872 25131 2904 25163
rect 2944 25131 2976 25163
rect 3016 25131 3048 25163
rect 3088 25131 3120 25163
rect 3160 25131 3192 25163
rect 3232 25131 3264 25163
rect 3304 25131 3336 25163
rect 3376 25131 3408 25163
rect 3448 25131 3480 25163
rect 3520 25131 3552 25163
rect 3592 25131 3624 25163
rect 3664 25131 3696 25163
rect 3736 25131 3768 25163
rect 3808 25131 3840 25163
rect 3880 25131 3912 25163
rect 3952 25131 3984 25163
rect 4024 25131 4056 25163
rect 4096 25131 4128 25163
rect 4168 25131 4200 25163
rect 4240 25131 4272 25163
rect 4312 25131 4344 25163
rect 4384 25131 4416 25163
rect 4456 25131 4488 25163
rect 4528 25131 4560 25163
rect 4600 25131 4632 25163
rect 4672 25131 4704 25163
rect 4744 25131 4776 25163
rect 4816 25131 4848 25163
rect 4888 25131 4920 25163
rect 4960 25131 4992 25163
rect 5032 25131 5064 25163
rect 5104 25131 5136 25163
rect 5176 25131 5208 25163
rect 5248 25131 5280 25163
rect 5320 25131 5352 25163
rect 5392 25131 5424 25163
rect 5464 25131 5496 25163
rect 5536 25131 5568 25163
rect 5608 25131 5640 25163
rect 5680 25131 5712 25163
rect 5752 25131 5784 25163
rect 5824 25131 5856 25163
rect 5896 25131 5928 25163
rect 5968 25131 6000 25163
rect 6040 25131 6072 25163
rect 6112 25131 6144 25163
rect 6184 25131 6216 25163
rect 6256 25131 6288 25163
rect 6328 25131 6360 25163
rect 6400 25131 6432 25163
rect 6472 25131 6504 25163
rect 6544 25131 6576 25163
rect 6616 25131 6648 25163
rect 6688 25131 6720 25163
rect 6760 25131 6792 25163
rect 6832 25131 6864 25163
rect 6904 25131 6936 25163
rect 6976 25131 7008 25163
rect 7048 25131 7080 25163
rect 7120 25131 7152 25163
rect 7192 25131 7224 25163
rect 7264 25131 7296 25163
rect 7336 25131 7368 25163
rect 7408 25131 7440 25163
rect 7480 25131 7512 25163
rect 7552 25131 7584 25163
rect 7624 25131 7656 25163
rect 7696 25131 7728 25163
rect 7768 25131 7800 25163
rect 7840 25131 7872 25163
rect 7912 25131 7944 25163
rect 7984 25131 8016 25163
rect 8056 25131 8088 25163
rect 8128 25131 8160 25163
rect 8200 25131 8232 25163
rect 8272 25131 8304 25163
rect 8344 25131 8376 25163
rect 8416 25131 8448 25163
rect 8488 25131 8520 25163
rect 8560 25131 8592 25163
rect 8632 25131 8664 25163
rect 8704 25131 8736 25163
rect 8776 25131 8808 25163
rect 8848 25131 8880 25163
rect 8920 25131 8952 25163
rect 8992 25131 9024 25163
rect 9064 25131 9096 25163
rect 9136 25131 9168 25163
rect 9208 25131 9240 25163
rect 9280 25131 9312 25163
rect 9352 25131 9384 25163
rect 9424 25131 9456 25163
rect 9496 25131 9528 25163
rect 9568 25131 9600 25163
rect 9640 25131 9672 25163
rect 9712 25131 9744 25163
rect 9784 25131 9816 25163
rect 9856 25131 9888 25163
rect 9928 25131 9960 25163
rect 10000 25131 10032 25163
rect 10072 25131 10104 25163
rect 10144 25131 10176 25163
rect 10216 25131 10248 25163
rect 10288 25131 10320 25163
rect 10360 25131 10392 25163
rect 10432 25131 10464 25163
rect 10504 25131 10536 25163
rect 10576 25131 10608 25163
rect 10648 25131 10680 25163
rect 10720 25131 10752 25163
rect 10792 25131 10824 25163
rect 10864 25131 10896 25163
rect 10936 25131 10968 25163
rect 11008 25131 11040 25163
rect 11080 25131 11112 25163
rect 11152 25131 11184 25163
rect 11224 25131 11256 25163
rect 11296 25131 11328 25163
rect 11368 25131 11400 25163
rect 11440 25131 11472 25163
rect 11512 25131 11544 25163
rect 11584 25131 11616 25163
rect 11656 25131 11688 25163
rect 11728 25131 11760 25163
rect 11800 25131 11832 25163
rect 11872 25131 11904 25163
rect 11944 25131 11976 25163
rect 12016 25131 12048 25163
rect 12088 25131 12120 25163
rect 12160 25131 12192 25163
rect 12232 25131 12264 25163
rect 12304 25131 12336 25163
rect 12376 25131 12408 25163
rect 12448 25131 12480 25163
rect 12520 25131 12552 25163
rect 12592 25131 12624 25163
rect 12664 25131 12696 25163
rect 12736 25131 12768 25163
rect 12808 25131 12840 25163
rect 12880 25131 12912 25163
rect 12952 25131 12984 25163
rect 13024 25131 13056 25163
rect 13096 25131 13128 25163
rect 13168 25131 13200 25163
rect 13240 25131 13272 25163
rect 13312 25131 13344 25163
rect 13384 25131 13416 25163
rect 13456 25131 13488 25163
rect 13528 25131 13560 25163
rect 13600 25131 13632 25163
rect 13672 25131 13704 25163
rect 13744 25131 13776 25163
rect 13816 25131 13848 25163
rect 13888 25131 13920 25163
rect 13960 25131 13992 25163
rect 14032 25131 14064 25163
rect 14104 25131 14136 25163
rect 14176 25131 14208 25163
rect 14248 25131 14280 25163
rect 14320 25131 14352 25163
rect 14392 25131 14424 25163
rect 14464 25131 14496 25163
rect 14536 25131 14568 25163
rect 14608 25131 14640 25163
rect 14680 25131 14712 25163
rect 14752 25131 14784 25163
rect 14824 25131 14856 25163
rect 14896 25131 14928 25163
rect 14968 25131 15000 25163
rect 15040 25131 15072 25163
rect 15112 25131 15144 25163
rect 15184 25131 15216 25163
rect 15256 25131 15288 25163
rect 15328 25131 15360 25163
rect 15400 25131 15432 25163
rect 15472 25131 15504 25163
rect 15544 25131 15576 25163
rect 15616 25131 15648 25163
rect 15688 25131 15720 25163
rect 15760 25131 15792 25163
rect 15832 25131 15864 25163
rect 15904 25131 15936 25163
rect 64 25059 96 25091
rect 136 25059 168 25091
rect 208 25059 240 25091
rect 280 25059 312 25091
rect 352 25059 384 25091
rect 424 25059 456 25091
rect 496 25059 528 25091
rect 568 25059 600 25091
rect 640 25059 672 25091
rect 712 25059 744 25091
rect 784 25059 816 25091
rect 856 25059 888 25091
rect 928 25059 960 25091
rect 1000 25059 1032 25091
rect 1072 25059 1104 25091
rect 1144 25059 1176 25091
rect 1216 25059 1248 25091
rect 1288 25059 1320 25091
rect 1360 25059 1392 25091
rect 1432 25059 1464 25091
rect 1504 25059 1536 25091
rect 1576 25059 1608 25091
rect 1648 25059 1680 25091
rect 1720 25059 1752 25091
rect 1792 25059 1824 25091
rect 1864 25059 1896 25091
rect 1936 25059 1968 25091
rect 2008 25059 2040 25091
rect 2080 25059 2112 25091
rect 2152 25059 2184 25091
rect 2224 25059 2256 25091
rect 2296 25059 2328 25091
rect 2368 25059 2400 25091
rect 2440 25059 2472 25091
rect 2512 25059 2544 25091
rect 2584 25059 2616 25091
rect 2656 25059 2688 25091
rect 2728 25059 2760 25091
rect 2800 25059 2832 25091
rect 2872 25059 2904 25091
rect 2944 25059 2976 25091
rect 3016 25059 3048 25091
rect 3088 25059 3120 25091
rect 3160 25059 3192 25091
rect 3232 25059 3264 25091
rect 3304 25059 3336 25091
rect 3376 25059 3408 25091
rect 3448 25059 3480 25091
rect 3520 25059 3552 25091
rect 3592 25059 3624 25091
rect 3664 25059 3696 25091
rect 3736 25059 3768 25091
rect 3808 25059 3840 25091
rect 3880 25059 3912 25091
rect 3952 25059 3984 25091
rect 4024 25059 4056 25091
rect 4096 25059 4128 25091
rect 4168 25059 4200 25091
rect 4240 25059 4272 25091
rect 4312 25059 4344 25091
rect 4384 25059 4416 25091
rect 4456 25059 4488 25091
rect 4528 25059 4560 25091
rect 4600 25059 4632 25091
rect 4672 25059 4704 25091
rect 4744 25059 4776 25091
rect 4816 25059 4848 25091
rect 4888 25059 4920 25091
rect 4960 25059 4992 25091
rect 5032 25059 5064 25091
rect 5104 25059 5136 25091
rect 5176 25059 5208 25091
rect 5248 25059 5280 25091
rect 5320 25059 5352 25091
rect 5392 25059 5424 25091
rect 5464 25059 5496 25091
rect 5536 25059 5568 25091
rect 5608 25059 5640 25091
rect 5680 25059 5712 25091
rect 5752 25059 5784 25091
rect 5824 25059 5856 25091
rect 5896 25059 5928 25091
rect 5968 25059 6000 25091
rect 6040 25059 6072 25091
rect 6112 25059 6144 25091
rect 6184 25059 6216 25091
rect 6256 25059 6288 25091
rect 6328 25059 6360 25091
rect 6400 25059 6432 25091
rect 6472 25059 6504 25091
rect 6544 25059 6576 25091
rect 6616 25059 6648 25091
rect 6688 25059 6720 25091
rect 6760 25059 6792 25091
rect 6832 25059 6864 25091
rect 6904 25059 6936 25091
rect 6976 25059 7008 25091
rect 7048 25059 7080 25091
rect 7120 25059 7152 25091
rect 7192 25059 7224 25091
rect 7264 25059 7296 25091
rect 7336 25059 7368 25091
rect 7408 25059 7440 25091
rect 7480 25059 7512 25091
rect 7552 25059 7584 25091
rect 7624 25059 7656 25091
rect 7696 25059 7728 25091
rect 7768 25059 7800 25091
rect 7840 25059 7872 25091
rect 7912 25059 7944 25091
rect 7984 25059 8016 25091
rect 8056 25059 8088 25091
rect 8128 25059 8160 25091
rect 8200 25059 8232 25091
rect 8272 25059 8304 25091
rect 8344 25059 8376 25091
rect 8416 25059 8448 25091
rect 8488 25059 8520 25091
rect 8560 25059 8592 25091
rect 8632 25059 8664 25091
rect 8704 25059 8736 25091
rect 8776 25059 8808 25091
rect 8848 25059 8880 25091
rect 8920 25059 8952 25091
rect 8992 25059 9024 25091
rect 9064 25059 9096 25091
rect 9136 25059 9168 25091
rect 9208 25059 9240 25091
rect 9280 25059 9312 25091
rect 9352 25059 9384 25091
rect 9424 25059 9456 25091
rect 9496 25059 9528 25091
rect 9568 25059 9600 25091
rect 9640 25059 9672 25091
rect 9712 25059 9744 25091
rect 9784 25059 9816 25091
rect 9856 25059 9888 25091
rect 9928 25059 9960 25091
rect 10000 25059 10032 25091
rect 10072 25059 10104 25091
rect 10144 25059 10176 25091
rect 10216 25059 10248 25091
rect 10288 25059 10320 25091
rect 10360 25059 10392 25091
rect 10432 25059 10464 25091
rect 10504 25059 10536 25091
rect 10576 25059 10608 25091
rect 10648 25059 10680 25091
rect 10720 25059 10752 25091
rect 10792 25059 10824 25091
rect 10864 25059 10896 25091
rect 10936 25059 10968 25091
rect 11008 25059 11040 25091
rect 11080 25059 11112 25091
rect 11152 25059 11184 25091
rect 11224 25059 11256 25091
rect 11296 25059 11328 25091
rect 11368 25059 11400 25091
rect 11440 25059 11472 25091
rect 11512 25059 11544 25091
rect 11584 25059 11616 25091
rect 11656 25059 11688 25091
rect 11728 25059 11760 25091
rect 11800 25059 11832 25091
rect 11872 25059 11904 25091
rect 11944 25059 11976 25091
rect 12016 25059 12048 25091
rect 12088 25059 12120 25091
rect 12160 25059 12192 25091
rect 12232 25059 12264 25091
rect 12304 25059 12336 25091
rect 12376 25059 12408 25091
rect 12448 25059 12480 25091
rect 12520 25059 12552 25091
rect 12592 25059 12624 25091
rect 12664 25059 12696 25091
rect 12736 25059 12768 25091
rect 12808 25059 12840 25091
rect 12880 25059 12912 25091
rect 12952 25059 12984 25091
rect 13024 25059 13056 25091
rect 13096 25059 13128 25091
rect 13168 25059 13200 25091
rect 13240 25059 13272 25091
rect 13312 25059 13344 25091
rect 13384 25059 13416 25091
rect 13456 25059 13488 25091
rect 13528 25059 13560 25091
rect 13600 25059 13632 25091
rect 13672 25059 13704 25091
rect 13744 25059 13776 25091
rect 13816 25059 13848 25091
rect 13888 25059 13920 25091
rect 13960 25059 13992 25091
rect 14032 25059 14064 25091
rect 14104 25059 14136 25091
rect 14176 25059 14208 25091
rect 14248 25059 14280 25091
rect 14320 25059 14352 25091
rect 14392 25059 14424 25091
rect 14464 25059 14496 25091
rect 14536 25059 14568 25091
rect 14608 25059 14640 25091
rect 14680 25059 14712 25091
rect 14752 25059 14784 25091
rect 14824 25059 14856 25091
rect 14896 25059 14928 25091
rect 14968 25059 15000 25091
rect 15040 25059 15072 25091
rect 15112 25059 15144 25091
rect 15184 25059 15216 25091
rect 15256 25059 15288 25091
rect 15328 25059 15360 25091
rect 15400 25059 15432 25091
rect 15472 25059 15504 25091
rect 15544 25059 15576 25091
rect 15616 25059 15648 25091
rect 15688 25059 15720 25091
rect 15760 25059 15792 25091
rect 15832 25059 15864 25091
rect 15904 25059 15936 25091
rect 64 24987 96 25019
rect 136 24987 168 25019
rect 208 24987 240 25019
rect 280 24987 312 25019
rect 352 24987 384 25019
rect 424 24987 456 25019
rect 496 24987 528 25019
rect 568 24987 600 25019
rect 640 24987 672 25019
rect 712 24987 744 25019
rect 784 24987 816 25019
rect 856 24987 888 25019
rect 928 24987 960 25019
rect 1000 24987 1032 25019
rect 1072 24987 1104 25019
rect 1144 24987 1176 25019
rect 1216 24987 1248 25019
rect 1288 24987 1320 25019
rect 1360 24987 1392 25019
rect 1432 24987 1464 25019
rect 1504 24987 1536 25019
rect 1576 24987 1608 25019
rect 1648 24987 1680 25019
rect 1720 24987 1752 25019
rect 1792 24987 1824 25019
rect 1864 24987 1896 25019
rect 1936 24987 1968 25019
rect 2008 24987 2040 25019
rect 2080 24987 2112 25019
rect 2152 24987 2184 25019
rect 2224 24987 2256 25019
rect 2296 24987 2328 25019
rect 2368 24987 2400 25019
rect 2440 24987 2472 25019
rect 2512 24987 2544 25019
rect 2584 24987 2616 25019
rect 2656 24987 2688 25019
rect 2728 24987 2760 25019
rect 2800 24987 2832 25019
rect 2872 24987 2904 25019
rect 2944 24987 2976 25019
rect 3016 24987 3048 25019
rect 3088 24987 3120 25019
rect 3160 24987 3192 25019
rect 3232 24987 3264 25019
rect 3304 24987 3336 25019
rect 3376 24987 3408 25019
rect 3448 24987 3480 25019
rect 3520 24987 3552 25019
rect 3592 24987 3624 25019
rect 3664 24987 3696 25019
rect 3736 24987 3768 25019
rect 3808 24987 3840 25019
rect 3880 24987 3912 25019
rect 3952 24987 3984 25019
rect 4024 24987 4056 25019
rect 4096 24987 4128 25019
rect 4168 24987 4200 25019
rect 4240 24987 4272 25019
rect 4312 24987 4344 25019
rect 4384 24987 4416 25019
rect 4456 24987 4488 25019
rect 4528 24987 4560 25019
rect 4600 24987 4632 25019
rect 4672 24987 4704 25019
rect 4744 24987 4776 25019
rect 4816 24987 4848 25019
rect 4888 24987 4920 25019
rect 4960 24987 4992 25019
rect 5032 24987 5064 25019
rect 5104 24987 5136 25019
rect 5176 24987 5208 25019
rect 5248 24987 5280 25019
rect 5320 24987 5352 25019
rect 5392 24987 5424 25019
rect 5464 24987 5496 25019
rect 5536 24987 5568 25019
rect 5608 24987 5640 25019
rect 5680 24987 5712 25019
rect 5752 24987 5784 25019
rect 5824 24987 5856 25019
rect 5896 24987 5928 25019
rect 5968 24987 6000 25019
rect 6040 24987 6072 25019
rect 6112 24987 6144 25019
rect 6184 24987 6216 25019
rect 6256 24987 6288 25019
rect 6328 24987 6360 25019
rect 6400 24987 6432 25019
rect 6472 24987 6504 25019
rect 6544 24987 6576 25019
rect 6616 24987 6648 25019
rect 6688 24987 6720 25019
rect 6760 24987 6792 25019
rect 6832 24987 6864 25019
rect 6904 24987 6936 25019
rect 6976 24987 7008 25019
rect 7048 24987 7080 25019
rect 7120 24987 7152 25019
rect 7192 24987 7224 25019
rect 7264 24987 7296 25019
rect 7336 24987 7368 25019
rect 7408 24987 7440 25019
rect 7480 24987 7512 25019
rect 7552 24987 7584 25019
rect 7624 24987 7656 25019
rect 7696 24987 7728 25019
rect 7768 24987 7800 25019
rect 7840 24987 7872 25019
rect 7912 24987 7944 25019
rect 7984 24987 8016 25019
rect 8056 24987 8088 25019
rect 8128 24987 8160 25019
rect 8200 24987 8232 25019
rect 8272 24987 8304 25019
rect 8344 24987 8376 25019
rect 8416 24987 8448 25019
rect 8488 24987 8520 25019
rect 8560 24987 8592 25019
rect 8632 24987 8664 25019
rect 8704 24987 8736 25019
rect 8776 24987 8808 25019
rect 8848 24987 8880 25019
rect 8920 24987 8952 25019
rect 8992 24987 9024 25019
rect 9064 24987 9096 25019
rect 9136 24987 9168 25019
rect 9208 24987 9240 25019
rect 9280 24987 9312 25019
rect 9352 24987 9384 25019
rect 9424 24987 9456 25019
rect 9496 24987 9528 25019
rect 9568 24987 9600 25019
rect 9640 24987 9672 25019
rect 9712 24987 9744 25019
rect 9784 24987 9816 25019
rect 9856 24987 9888 25019
rect 9928 24987 9960 25019
rect 10000 24987 10032 25019
rect 10072 24987 10104 25019
rect 10144 24987 10176 25019
rect 10216 24987 10248 25019
rect 10288 24987 10320 25019
rect 10360 24987 10392 25019
rect 10432 24987 10464 25019
rect 10504 24987 10536 25019
rect 10576 24987 10608 25019
rect 10648 24987 10680 25019
rect 10720 24987 10752 25019
rect 10792 24987 10824 25019
rect 10864 24987 10896 25019
rect 10936 24987 10968 25019
rect 11008 24987 11040 25019
rect 11080 24987 11112 25019
rect 11152 24987 11184 25019
rect 11224 24987 11256 25019
rect 11296 24987 11328 25019
rect 11368 24987 11400 25019
rect 11440 24987 11472 25019
rect 11512 24987 11544 25019
rect 11584 24987 11616 25019
rect 11656 24987 11688 25019
rect 11728 24987 11760 25019
rect 11800 24987 11832 25019
rect 11872 24987 11904 25019
rect 11944 24987 11976 25019
rect 12016 24987 12048 25019
rect 12088 24987 12120 25019
rect 12160 24987 12192 25019
rect 12232 24987 12264 25019
rect 12304 24987 12336 25019
rect 12376 24987 12408 25019
rect 12448 24987 12480 25019
rect 12520 24987 12552 25019
rect 12592 24987 12624 25019
rect 12664 24987 12696 25019
rect 12736 24987 12768 25019
rect 12808 24987 12840 25019
rect 12880 24987 12912 25019
rect 12952 24987 12984 25019
rect 13024 24987 13056 25019
rect 13096 24987 13128 25019
rect 13168 24987 13200 25019
rect 13240 24987 13272 25019
rect 13312 24987 13344 25019
rect 13384 24987 13416 25019
rect 13456 24987 13488 25019
rect 13528 24987 13560 25019
rect 13600 24987 13632 25019
rect 13672 24987 13704 25019
rect 13744 24987 13776 25019
rect 13816 24987 13848 25019
rect 13888 24987 13920 25019
rect 13960 24987 13992 25019
rect 14032 24987 14064 25019
rect 14104 24987 14136 25019
rect 14176 24987 14208 25019
rect 14248 24987 14280 25019
rect 14320 24987 14352 25019
rect 14392 24987 14424 25019
rect 14464 24987 14496 25019
rect 14536 24987 14568 25019
rect 14608 24987 14640 25019
rect 14680 24987 14712 25019
rect 14752 24987 14784 25019
rect 14824 24987 14856 25019
rect 14896 24987 14928 25019
rect 14968 24987 15000 25019
rect 15040 24987 15072 25019
rect 15112 24987 15144 25019
rect 15184 24987 15216 25019
rect 15256 24987 15288 25019
rect 15328 24987 15360 25019
rect 15400 24987 15432 25019
rect 15472 24987 15504 25019
rect 15544 24987 15576 25019
rect 15616 24987 15648 25019
rect 15688 24987 15720 25019
rect 15760 24987 15792 25019
rect 15832 24987 15864 25019
rect 15904 24987 15936 25019
rect 64 24915 96 24947
rect 136 24915 168 24947
rect 208 24915 240 24947
rect 280 24915 312 24947
rect 352 24915 384 24947
rect 424 24915 456 24947
rect 496 24915 528 24947
rect 568 24915 600 24947
rect 640 24915 672 24947
rect 712 24915 744 24947
rect 784 24915 816 24947
rect 856 24915 888 24947
rect 928 24915 960 24947
rect 1000 24915 1032 24947
rect 1072 24915 1104 24947
rect 1144 24915 1176 24947
rect 1216 24915 1248 24947
rect 1288 24915 1320 24947
rect 1360 24915 1392 24947
rect 1432 24915 1464 24947
rect 1504 24915 1536 24947
rect 1576 24915 1608 24947
rect 1648 24915 1680 24947
rect 1720 24915 1752 24947
rect 1792 24915 1824 24947
rect 1864 24915 1896 24947
rect 1936 24915 1968 24947
rect 2008 24915 2040 24947
rect 2080 24915 2112 24947
rect 2152 24915 2184 24947
rect 2224 24915 2256 24947
rect 2296 24915 2328 24947
rect 2368 24915 2400 24947
rect 2440 24915 2472 24947
rect 2512 24915 2544 24947
rect 2584 24915 2616 24947
rect 2656 24915 2688 24947
rect 2728 24915 2760 24947
rect 2800 24915 2832 24947
rect 2872 24915 2904 24947
rect 2944 24915 2976 24947
rect 3016 24915 3048 24947
rect 3088 24915 3120 24947
rect 3160 24915 3192 24947
rect 3232 24915 3264 24947
rect 3304 24915 3336 24947
rect 3376 24915 3408 24947
rect 3448 24915 3480 24947
rect 3520 24915 3552 24947
rect 3592 24915 3624 24947
rect 3664 24915 3696 24947
rect 3736 24915 3768 24947
rect 3808 24915 3840 24947
rect 3880 24915 3912 24947
rect 3952 24915 3984 24947
rect 4024 24915 4056 24947
rect 4096 24915 4128 24947
rect 4168 24915 4200 24947
rect 4240 24915 4272 24947
rect 4312 24915 4344 24947
rect 4384 24915 4416 24947
rect 4456 24915 4488 24947
rect 4528 24915 4560 24947
rect 4600 24915 4632 24947
rect 4672 24915 4704 24947
rect 4744 24915 4776 24947
rect 4816 24915 4848 24947
rect 4888 24915 4920 24947
rect 4960 24915 4992 24947
rect 5032 24915 5064 24947
rect 5104 24915 5136 24947
rect 5176 24915 5208 24947
rect 5248 24915 5280 24947
rect 5320 24915 5352 24947
rect 5392 24915 5424 24947
rect 5464 24915 5496 24947
rect 5536 24915 5568 24947
rect 5608 24915 5640 24947
rect 5680 24915 5712 24947
rect 5752 24915 5784 24947
rect 5824 24915 5856 24947
rect 5896 24915 5928 24947
rect 5968 24915 6000 24947
rect 6040 24915 6072 24947
rect 6112 24915 6144 24947
rect 6184 24915 6216 24947
rect 6256 24915 6288 24947
rect 6328 24915 6360 24947
rect 6400 24915 6432 24947
rect 6472 24915 6504 24947
rect 6544 24915 6576 24947
rect 6616 24915 6648 24947
rect 6688 24915 6720 24947
rect 6760 24915 6792 24947
rect 6832 24915 6864 24947
rect 6904 24915 6936 24947
rect 6976 24915 7008 24947
rect 7048 24915 7080 24947
rect 7120 24915 7152 24947
rect 7192 24915 7224 24947
rect 7264 24915 7296 24947
rect 7336 24915 7368 24947
rect 7408 24915 7440 24947
rect 7480 24915 7512 24947
rect 7552 24915 7584 24947
rect 7624 24915 7656 24947
rect 7696 24915 7728 24947
rect 7768 24915 7800 24947
rect 7840 24915 7872 24947
rect 7912 24915 7944 24947
rect 7984 24915 8016 24947
rect 8056 24915 8088 24947
rect 8128 24915 8160 24947
rect 8200 24915 8232 24947
rect 8272 24915 8304 24947
rect 8344 24915 8376 24947
rect 8416 24915 8448 24947
rect 8488 24915 8520 24947
rect 8560 24915 8592 24947
rect 8632 24915 8664 24947
rect 8704 24915 8736 24947
rect 8776 24915 8808 24947
rect 8848 24915 8880 24947
rect 8920 24915 8952 24947
rect 8992 24915 9024 24947
rect 9064 24915 9096 24947
rect 9136 24915 9168 24947
rect 9208 24915 9240 24947
rect 9280 24915 9312 24947
rect 9352 24915 9384 24947
rect 9424 24915 9456 24947
rect 9496 24915 9528 24947
rect 9568 24915 9600 24947
rect 9640 24915 9672 24947
rect 9712 24915 9744 24947
rect 9784 24915 9816 24947
rect 9856 24915 9888 24947
rect 9928 24915 9960 24947
rect 10000 24915 10032 24947
rect 10072 24915 10104 24947
rect 10144 24915 10176 24947
rect 10216 24915 10248 24947
rect 10288 24915 10320 24947
rect 10360 24915 10392 24947
rect 10432 24915 10464 24947
rect 10504 24915 10536 24947
rect 10576 24915 10608 24947
rect 10648 24915 10680 24947
rect 10720 24915 10752 24947
rect 10792 24915 10824 24947
rect 10864 24915 10896 24947
rect 10936 24915 10968 24947
rect 11008 24915 11040 24947
rect 11080 24915 11112 24947
rect 11152 24915 11184 24947
rect 11224 24915 11256 24947
rect 11296 24915 11328 24947
rect 11368 24915 11400 24947
rect 11440 24915 11472 24947
rect 11512 24915 11544 24947
rect 11584 24915 11616 24947
rect 11656 24915 11688 24947
rect 11728 24915 11760 24947
rect 11800 24915 11832 24947
rect 11872 24915 11904 24947
rect 11944 24915 11976 24947
rect 12016 24915 12048 24947
rect 12088 24915 12120 24947
rect 12160 24915 12192 24947
rect 12232 24915 12264 24947
rect 12304 24915 12336 24947
rect 12376 24915 12408 24947
rect 12448 24915 12480 24947
rect 12520 24915 12552 24947
rect 12592 24915 12624 24947
rect 12664 24915 12696 24947
rect 12736 24915 12768 24947
rect 12808 24915 12840 24947
rect 12880 24915 12912 24947
rect 12952 24915 12984 24947
rect 13024 24915 13056 24947
rect 13096 24915 13128 24947
rect 13168 24915 13200 24947
rect 13240 24915 13272 24947
rect 13312 24915 13344 24947
rect 13384 24915 13416 24947
rect 13456 24915 13488 24947
rect 13528 24915 13560 24947
rect 13600 24915 13632 24947
rect 13672 24915 13704 24947
rect 13744 24915 13776 24947
rect 13816 24915 13848 24947
rect 13888 24915 13920 24947
rect 13960 24915 13992 24947
rect 14032 24915 14064 24947
rect 14104 24915 14136 24947
rect 14176 24915 14208 24947
rect 14248 24915 14280 24947
rect 14320 24915 14352 24947
rect 14392 24915 14424 24947
rect 14464 24915 14496 24947
rect 14536 24915 14568 24947
rect 14608 24915 14640 24947
rect 14680 24915 14712 24947
rect 14752 24915 14784 24947
rect 14824 24915 14856 24947
rect 14896 24915 14928 24947
rect 14968 24915 15000 24947
rect 15040 24915 15072 24947
rect 15112 24915 15144 24947
rect 15184 24915 15216 24947
rect 15256 24915 15288 24947
rect 15328 24915 15360 24947
rect 15400 24915 15432 24947
rect 15472 24915 15504 24947
rect 15544 24915 15576 24947
rect 15616 24915 15648 24947
rect 15688 24915 15720 24947
rect 15760 24915 15792 24947
rect 15832 24915 15864 24947
rect 15904 24915 15936 24947
rect 64 24843 96 24875
rect 136 24843 168 24875
rect 208 24843 240 24875
rect 280 24843 312 24875
rect 352 24843 384 24875
rect 424 24843 456 24875
rect 496 24843 528 24875
rect 568 24843 600 24875
rect 640 24843 672 24875
rect 712 24843 744 24875
rect 784 24843 816 24875
rect 856 24843 888 24875
rect 928 24843 960 24875
rect 1000 24843 1032 24875
rect 1072 24843 1104 24875
rect 1144 24843 1176 24875
rect 1216 24843 1248 24875
rect 1288 24843 1320 24875
rect 1360 24843 1392 24875
rect 1432 24843 1464 24875
rect 1504 24843 1536 24875
rect 1576 24843 1608 24875
rect 1648 24843 1680 24875
rect 1720 24843 1752 24875
rect 1792 24843 1824 24875
rect 1864 24843 1896 24875
rect 1936 24843 1968 24875
rect 2008 24843 2040 24875
rect 2080 24843 2112 24875
rect 2152 24843 2184 24875
rect 2224 24843 2256 24875
rect 2296 24843 2328 24875
rect 2368 24843 2400 24875
rect 2440 24843 2472 24875
rect 2512 24843 2544 24875
rect 2584 24843 2616 24875
rect 2656 24843 2688 24875
rect 2728 24843 2760 24875
rect 2800 24843 2832 24875
rect 2872 24843 2904 24875
rect 2944 24843 2976 24875
rect 3016 24843 3048 24875
rect 3088 24843 3120 24875
rect 3160 24843 3192 24875
rect 3232 24843 3264 24875
rect 3304 24843 3336 24875
rect 3376 24843 3408 24875
rect 3448 24843 3480 24875
rect 3520 24843 3552 24875
rect 3592 24843 3624 24875
rect 3664 24843 3696 24875
rect 3736 24843 3768 24875
rect 3808 24843 3840 24875
rect 3880 24843 3912 24875
rect 3952 24843 3984 24875
rect 4024 24843 4056 24875
rect 4096 24843 4128 24875
rect 4168 24843 4200 24875
rect 4240 24843 4272 24875
rect 4312 24843 4344 24875
rect 4384 24843 4416 24875
rect 4456 24843 4488 24875
rect 4528 24843 4560 24875
rect 4600 24843 4632 24875
rect 4672 24843 4704 24875
rect 4744 24843 4776 24875
rect 4816 24843 4848 24875
rect 4888 24843 4920 24875
rect 4960 24843 4992 24875
rect 5032 24843 5064 24875
rect 5104 24843 5136 24875
rect 5176 24843 5208 24875
rect 5248 24843 5280 24875
rect 5320 24843 5352 24875
rect 5392 24843 5424 24875
rect 5464 24843 5496 24875
rect 5536 24843 5568 24875
rect 5608 24843 5640 24875
rect 5680 24843 5712 24875
rect 5752 24843 5784 24875
rect 5824 24843 5856 24875
rect 5896 24843 5928 24875
rect 5968 24843 6000 24875
rect 6040 24843 6072 24875
rect 6112 24843 6144 24875
rect 6184 24843 6216 24875
rect 6256 24843 6288 24875
rect 6328 24843 6360 24875
rect 6400 24843 6432 24875
rect 6472 24843 6504 24875
rect 6544 24843 6576 24875
rect 6616 24843 6648 24875
rect 6688 24843 6720 24875
rect 6760 24843 6792 24875
rect 6832 24843 6864 24875
rect 6904 24843 6936 24875
rect 6976 24843 7008 24875
rect 7048 24843 7080 24875
rect 7120 24843 7152 24875
rect 7192 24843 7224 24875
rect 7264 24843 7296 24875
rect 7336 24843 7368 24875
rect 7408 24843 7440 24875
rect 7480 24843 7512 24875
rect 7552 24843 7584 24875
rect 7624 24843 7656 24875
rect 7696 24843 7728 24875
rect 7768 24843 7800 24875
rect 7840 24843 7872 24875
rect 7912 24843 7944 24875
rect 7984 24843 8016 24875
rect 8056 24843 8088 24875
rect 8128 24843 8160 24875
rect 8200 24843 8232 24875
rect 8272 24843 8304 24875
rect 8344 24843 8376 24875
rect 8416 24843 8448 24875
rect 8488 24843 8520 24875
rect 8560 24843 8592 24875
rect 8632 24843 8664 24875
rect 8704 24843 8736 24875
rect 8776 24843 8808 24875
rect 8848 24843 8880 24875
rect 8920 24843 8952 24875
rect 8992 24843 9024 24875
rect 9064 24843 9096 24875
rect 9136 24843 9168 24875
rect 9208 24843 9240 24875
rect 9280 24843 9312 24875
rect 9352 24843 9384 24875
rect 9424 24843 9456 24875
rect 9496 24843 9528 24875
rect 9568 24843 9600 24875
rect 9640 24843 9672 24875
rect 9712 24843 9744 24875
rect 9784 24843 9816 24875
rect 9856 24843 9888 24875
rect 9928 24843 9960 24875
rect 10000 24843 10032 24875
rect 10072 24843 10104 24875
rect 10144 24843 10176 24875
rect 10216 24843 10248 24875
rect 10288 24843 10320 24875
rect 10360 24843 10392 24875
rect 10432 24843 10464 24875
rect 10504 24843 10536 24875
rect 10576 24843 10608 24875
rect 10648 24843 10680 24875
rect 10720 24843 10752 24875
rect 10792 24843 10824 24875
rect 10864 24843 10896 24875
rect 10936 24843 10968 24875
rect 11008 24843 11040 24875
rect 11080 24843 11112 24875
rect 11152 24843 11184 24875
rect 11224 24843 11256 24875
rect 11296 24843 11328 24875
rect 11368 24843 11400 24875
rect 11440 24843 11472 24875
rect 11512 24843 11544 24875
rect 11584 24843 11616 24875
rect 11656 24843 11688 24875
rect 11728 24843 11760 24875
rect 11800 24843 11832 24875
rect 11872 24843 11904 24875
rect 11944 24843 11976 24875
rect 12016 24843 12048 24875
rect 12088 24843 12120 24875
rect 12160 24843 12192 24875
rect 12232 24843 12264 24875
rect 12304 24843 12336 24875
rect 12376 24843 12408 24875
rect 12448 24843 12480 24875
rect 12520 24843 12552 24875
rect 12592 24843 12624 24875
rect 12664 24843 12696 24875
rect 12736 24843 12768 24875
rect 12808 24843 12840 24875
rect 12880 24843 12912 24875
rect 12952 24843 12984 24875
rect 13024 24843 13056 24875
rect 13096 24843 13128 24875
rect 13168 24843 13200 24875
rect 13240 24843 13272 24875
rect 13312 24843 13344 24875
rect 13384 24843 13416 24875
rect 13456 24843 13488 24875
rect 13528 24843 13560 24875
rect 13600 24843 13632 24875
rect 13672 24843 13704 24875
rect 13744 24843 13776 24875
rect 13816 24843 13848 24875
rect 13888 24843 13920 24875
rect 13960 24843 13992 24875
rect 14032 24843 14064 24875
rect 14104 24843 14136 24875
rect 14176 24843 14208 24875
rect 14248 24843 14280 24875
rect 14320 24843 14352 24875
rect 14392 24843 14424 24875
rect 14464 24843 14496 24875
rect 14536 24843 14568 24875
rect 14608 24843 14640 24875
rect 14680 24843 14712 24875
rect 14752 24843 14784 24875
rect 14824 24843 14856 24875
rect 14896 24843 14928 24875
rect 14968 24843 15000 24875
rect 15040 24843 15072 24875
rect 15112 24843 15144 24875
rect 15184 24843 15216 24875
rect 15256 24843 15288 24875
rect 15328 24843 15360 24875
rect 15400 24843 15432 24875
rect 15472 24843 15504 24875
rect 15544 24843 15576 24875
rect 15616 24843 15648 24875
rect 15688 24843 15720 24875
rect 15760 24843 15792 24875
rect 15832 24843 15864 24875
rect 15904 24843 15936 24875
rect 64 24771 96 24803
rect 136 24771 168 24803
rect 208 24771 240 24803
rect 280 24771 312 24803
rect 352 24771 384 24803
rect 424 24771 456 24803
rect 496 24771 528 24803
rect 568 24771 600 24803
rect 640 24771 672 24803
rect 712 24771 744 24803
rect 784 24771 816 24803
rect 856 24771 888 24803
rect 928 24771 960 24803
rect 1000 24771 1032 24803
rect 1072 24771 1104 24803
rect 1144 24771 1176 24803
rect 1216 24771 1248 24803
rect 1288 24771 1320 24803
rect 1360 24771 1392 24803
rect 1432 24771 1464 24803
rect 1504 24771 1536 24803
rect 1576 24771 1608 24803
rect 1648 24771 1680 24803
rect 1720 24771 1752 24803
rect 1792 24771 1824 24803
rect 1864 24771 1896 24803
rect 1936 24771 1968 24803
rect 2008 24771 2040 24803
rect 2080 24771 2112 24803
rect 2152 24771 2184 24803
rect 2224 24771 2256 24803
rect 2296 24771 2328 24803
rect 2368 24771 2400 24803
rect 2440 24771 2472 24803
rect 2512 24771 2544 24803
rect 2584 24771 2616 24803
rect 2656 24771 2688 24803
rect 2728 24771 2760 24803
rect 2800 24771 2832 24803
rect 2872 24771 2904 24803
rect 2944 24771 2976 24803
rect 3016 24771 3048 24803
rect 3088 24771 3120 24803
rect 3160 24771 3192 24803
rect 3232 24771 3264 24803
rect 3304 24771 3336 24803
rect 3376 24771 3408 24803
rect 3448 24771 3480 24803
rect 3520 24771 3552 24803
rect 3592 24771 3624 24803
rect 3664 24771 3696 24803
rect 3736 24771 3768 24803
rect 3808 24771 3840 24803
rect 3880 24771 3912 24803
rect 3952 24771 3984 24803
rect 4024 24771 4056 24803
rect 4096 24771 4128 24803
rect 4168 24771 4200 24803
rect 4240 24771 4272 24803
rect 4312 24771 4344 24803
rect 4384 24771 4416 24803
rect 4456 24771 4488 24803
rect 4528 24771 4560 24803
rect 4600 24771 4632 24803
rect 4672 24771 4704 24803
rect 4744 24771 4776 24803
rect 4816 24771 4848 24803
rect 4888 24771 4920 24803
rect 4960 24771 4992 24803
rect 5032 24771 5064 24803
rect 5104 24771 5136 24803
rect 5176 24771 5208 24803
rect 5248 24771 5280 24803
rect 5320 24771 5352 24803
rect 5392 24771 5424 24803
rect 5464 24771 5496 24803
rect 5536 24771 5568 24803
rect 5608 24771 5640 24803
rect 5680 24771 5712 24803
rect 5752 24771 5784 24803
rect 5824 24771 5856 24803
rect 5896 24771 5928 24803
rect 5968 24771 6000 24803
rect 6040 24771 6072 24803
rect 6112 24771 6144 24803
rect 6184 24771 6216 24803
rect 6256 24771 6288 24803
rect 6328 24771 6360 24803
rect 6400 24771 6432 24803
rect 6472 24771 6504 24803
rect 6544 24771 6576 24803
rect 6616 24771 6648 24803
rect 6688 24771 6720 24803
rect 6760 24771 6792 24803
rect 6832 24771 6864 24803
rect 6904 24771 6936 24803
rect 6976 24771 7008 24803
rect 7048 24771 7080 24803
rect 7120 24771 7152 24803
rect 7192 24771 7224 24803
rect 7264 24771 7296 24803
rect 7336 24771 7368 24803
rect 7408 24771 7440 24803
rect 7480 24771 7512 24803
rect 7552 24771 7584 24803
rect 7624 24771 7656 24803
rect 7696 24771 7728 24803
rect 7768 24771 7800 24803
rect 7840 24771 7872 24803
rect 7912 24771 7944 24803
rect 7984 24771 8016 24803
rect 8056 24771 8088 24803
rect 8128 24771 8160 24803
rect 8200 24771 8232 24803
rect 8272 24771 8304 24803
rect 8344 24771 8376 24803
rect 8416 24771 8448 24803
rect 8488 24771 8520 24803
rect 8560 24771 8592 24803
rect 8632 24771 8664 24803
rect 8704 24771 8736 24803
rect 8776 24771 8808 24803
rect 8848 24771 8880 24803
rect 8920 24771 8952 24803
rect 8992 24771 9024 24803
rect 9064 24771 9096 24803
rect 9136 24771 9168 24803
rect 9208 24771 9240 24803
rect 9280 24771 9312 24803
rect 9352 24771 9384 24803
rect 9424 24771 9456 24803
rect 9496 24771 9528 24803
rect 9568 24771 9600 24803
rect 9640 24771 9672 24803
rect 9712 24771 9744 24803
rect 9784 24771 9816 24803
rect 9856 24771 9888 24803
rect 9928 24771 9960 24803
rect 10000 24771 10032 24803
rect 10072 24771 10104 24803
rect 10144 24771 10176 24803
rect 10216 24771 10248 24803
rect 10288 24771 10320 24803
rect 10360 24771 10392 24803
rect 10432 24771 10464 24803
rect 10504 24771 10536 24803
rect 10576 24771 10608 24803
rect 10648 24771 10680 24803
rect 10720 24771 10752 24803
rect 10792 24771 10824 24803
rect 10864 24771 10896 24803
rect 10936 24771 10968 24803
rect 11008 24771 11040 24803
rect 11080 24771 11112 24803
rect 11152 24771 11184 24803
rect 11224 24771 11256 24803
rect 11296 24771 11328 24803
rect 11368 24771 11400 24803
rect 11440 24771 11472 24803
rect 11512 24771 11544 24803
rect 11584 24771 11616 24803
rect 11656 24771 11688 24803
rect 11728 24771 11760 24803
rect 11800 24771 11832 24803
rect 11872 24771 11904 24803
rect 11944 24771 11976 24803
rect 12016 24771 12048 24803
rect 12088 24771 12120 24803
rect 12160 24771 12192 24803
rect 12232 24771 12264 24803
rect 12304 24771 12336 24803
rect 12376 24771 12408 24803
rect 12448 24771 12480 24803
rect 12520 24771 12552 24803
rect 12592 24771 12624 24803
rect 12664 24771 12696 24803
rect 12736 24771 12768 24803
rect 12808 24771 12840 24803
rect 12880 24771 12912 24803
rect 12952 24771 12984 24803
rect 13024 24771 13056 24803
rect 13096 24771 13128 24803
rect 13168 24771 13200 24803
rect 13240 24771 13272 24803
rect 13312 24771 13344 24803
rect 13384 24771 13416 24803
rect 13456 24771 13488 24803
rect 13528 24771 13560 24803
rect 13600 24771 13632 24803
rect 13672 24771 13704 24803
rect 13744 24771 13776 24803
rect 13816 24771 13848 24803
rect 13888 24771 13920 24803
rect 13960 24771 13992 24803
rect 14032 24771 14064 24803
rect 14104 24771 14136 24803
rect 14176 24771 14208 24803
rect 14248 24771 14280 24803
rect 14320 24771 14352 24803
rect 14392 24771 14424 24803
rect 14464 24771 14496 24803
rect 14536 24771 14568 24803
rect 14608 24771 14640 24803
rect 14680 24771 14712 24803
rect 14752 24771 14784 24803
rect 14824 24771 14856 24803
rect 14896 24771 14928 24803
rect 14968 24771 15000 24803
rect 15040 24771 15072 24803
rect 15112 24771 15144 24803
rect 15184 24771 15216 24803
rect 15256 24771 15288 24803
rect 15328 24771 15360 24803
rect 15400 24771 15432 24803
rect 15472 24771 15504 24803
rect 15544 24771 15576 24803
rect 15616 24771 15648 24803
rect 15688 24771 15720 24803
rect 15760 24771 15792 24803
rect 15832 24771 15864 24803
rect 15904 24771 15936 24803
rect 64 24699 96 24731
rect 136 24699 168 24731
rect 208 24699 240 24731
rect 280 24699 312 24731
rect 352 24699 384 24731
rect 424 24699 456 24731
rect 496 24699 528 24731
rect 568 24699 600 24731
rect 640 24699 672 24731
rect 712 24699 744 24731
rect 784 24699 816 24731
rect 856 24699 888 24731
rect 928 24699 960 24731
rect 1000 24699 1032 24731
rect 1072 24699 1104 24731
rect 1144 24699 1176 24731
rect 1216 24699 1248 24731
rect 1288 24699 1320 24731
rect 1360 24699 1392 24731
rect 1432 24699 1464 24731
rect 1504 24699 1536 24731
rect 1576 24699 1608 24731
rect 1648 24699 1680 24731
rect 1720 24699 1752 24731
rect 1792 24699 1824 24731
rect 1864 24699 1896 24731
rect 1936 24699 1968 24731
rect 2008 24699 2040 24731
rect 2080 24699 2112 24731
rect 2152 24699 2184 24731
rect 2224 24699 2256 24731
rect 2296 24699 2328 24731
rect 2368 24699 2400 24731
rect 2440 24699 2472 24731
rect 2512 24699 2544 24731
rect 2584 24699 2616 24731
rect 2656 24699 2688 24731
rect 2728 24699 2760 24731
rect 2800 24699 2832 24731
rect 2872 24699 2904 24731
rect 2944 24699 2976 24731
rect 3016 24699 3048 24731
rect 3088 24699 3120 24731
rect 3160 24699 3192 24731
rect 3232 24699 3264 24731
rect 3304 24699 3336 24731
rect 3376 24699 3408 24731
rect 3448 24699 3480 24731
rect 3520 24699 3552 24731
rect 3592 24699 3624 24731
rect 3664 24699 3696 24731
rect 3736 24699 3768 24731
rect 3808 24699 3840 24731
rect 3880 24699 3912 24731
rect 3952 24699 3984 24731
rect 4024 24699 4056 24731
rect 4096 24699 4128 24731
rect 4168 24699 4200 24731
rect 4240 24699 4272 24731
rect 4312 24699 4344 24731
rect 4384 24699 4416 24731
rect 4456 24699 4488 24731
rect 4528 24699 4560 24731
rect 4600 24699 4632 24731
rect 4672 24699 4704 24731
rect 4744 24699 4776 24731
rect 4816 24699 4848 24731
rect 4888 24699 4920 24731
rect 4960 24699 4992 24731
rect 5032 24699 5064 24731
rect 5104 24699 5136 24731
rect 5176 24699 5208 24731
rect 5248 24699 5280 24731
rect 5320 24699 5352 24731
rect 5392 24699 5424 24731
rect 5464 24699 5496 24731
rect 5536 24699 5568 24731
rect 5608 24699 5640 24731
rect 5680 24699 5712 24731
rect 5752 24699 5784 24731
rect 5824 24699 5856 24731
rect 5896 24699 5928 24731
rect 5968 24699 6000 24731
rect 6040 24699 6072 24731
rect 6112 24699 6144 24731
rect 6184 24699 6216 24731
rect 6256 24699 6288 24731
rect 6328 24699 6360 24731
rect 6400 24699 6432 24731
rect 6472 24699 6504 24731
rect 6544 24699 6576 24731
rect 6616 24699 6648 24731
rect 6688 24699 6720 24731
rect 6760 24699 6792 24731
rect 6832 24699 6864 24731
rect 6904 24699 6936 24731
rect 6976 24699 7008 24731
rect 7048 24699 7080 24731
rect 7120 24699 7152 24731
rect 7192 24699 7224 24731
rect 7264 24699 7296 24731
rect 7336 24699 7368 24731
rect 7408 24699 7440 24731
rect 7480 24699 7512 24731
rect 7552 24699 7584 24731
rect 7624 24699 7656 24731
rect 7696 24699 7728 24731
rect 7768 24699 7800 24731
rect 7840 24699 7872 24731
rect 7912 24699 7944 24731
rect 7984 24699 8016 24731
rect 8056 24699 8088 24731
rect 8128 24699 8160 24731
rect 8200 24699 8232 24731
rect 8272 24699 8304 24731
rect 8344 24699 8376 24731
rect 8416 24699 8448 24731
rect 8488 24699 8520 24731
rect 8560 24699 8592 24731
rect 8632 24699 8664 24731
rect 8704 24699 8736 24731
rect 8776 24699 8808 24731
rect 8848 24699 8880 24731
rect 8920 24699 8952 24731
rect 8992 24699 9024 24731
rect 9064 24699 9096 24731
rect 9136 24699 9168 24731
rect 9208 24699 9240 24731
rect 9280 24699 9312 24731
rect 9352 24699 9384 24731
rect 9424 24699 9456 24731
rect 9496 24699 9528 24731
rect 9568 24699 9600 24731
rect 9640 24699 9672 24731
rect 9712 24699 9744 24731
rect 9784 24699 9816 24731
rect 9856 24699 9888 24731
rect 9928 24699 9960 24731
rect 10000 24699 10032 24731
rect 10072 24699 10104 24731
rect 10144 24699 10176 24731
rect 10216 24699 10248 24731
rect 10288 24699 10320 24731
rect 10360 24699 10392 24731
rect 10432 24699 10464 24731
rect 10504 24699 10536 24731
rect 10576 24699 10608 24731
rect 10648 24699 10680 24731
rect 10720 24699 10752 24731
rect 10792 24699 10824 24731
rect 10864 24699 10896 24731
rect 10936 24699 10968 24731
rect 11008 24699 11040 24731
rect 11080 24699 11112 24731
rect 11152 24699 11184 24731
rect 11224 24699 11256 24731
rect 11296 24699 11328 24731
rect 11368 24699 11400 24731
rect 11440 24699 11472 24731
rect 11512 24699 11544 24731
rect 11584 24699 11616 24731
rect 11656 24699 11688 24731
rect 11728 24699 11760 24731
rect 11800 24699 11832 24731
rect 11872 24699 11904 24731
rect 11944 24699 11976 24731
rect 12016 24699 12048 24731
rect 12088 24699 12120 24731
rect 12160 24699 12192 24731
rect 12232 24699 12264 24731
rect 12304 24699 12336 24731
rect 12376 24699 12408 24731
rect 12448 24699 12480 24731
rect 12520 24699 12552 24731
rect 12592 24699 12624 24731
rect 12664 24699 12696 24731
rect 12736 24699 12768 24731
rect 12808 24699 12840 24731
rect 12880 24699 12912 24731
rect 12952 24699 12984 24731
rect 13024 24699 13056 24731
rect 13096 24699 13128 24731
rect 13168 24699 13200 24731
rect 13240 24699 13272 24731
rect 13312 24699 13344 24731
rect 13384 24699 13416 24731
rect 13456 24699 13488 24731
rect 13528 24699 13560 24731
rect 13600 24699 13632 24731
rect 13672 24699 13704 24731
rect 13744 24699 13776 24731
rect 13816 24699 13848 24731
rect 13888 24699 13920 24731
rect 13960 24699 13992 24731
rect 14032 24699 14064 24731
rect 14104 24699 14136 24731
rect 14176 24699 14208 24731
rect 14248 24699 14280 24731
rect 14320 24699 14352 24731
rect 14392 24699 14424 24731
rect 14464 24699 14496 24731
rect 14536 24699 14568 24731
rect 14608 24699 14640 24731
rect 14680 24699 14712 24731
rect 14752 24699 14784 24731
rect 14824 24699 14856 24731
rect 14896 24699 14928 24731
rect 14968 24699 15000 24731
rect 15040 24699 15072 24731
rect 15112 24699 15144 24731
rect 15184 24699 15216 24731
rect 15256 24699 15288 24731
rect 15328 24699 15360 24731
rect 15400 24699 15432 24731
rect 15472 24699 15504 24731
rect 15544 24699 15576 24731
rect 15616 24699 15648 24731
rect 15688 24699 15720 24731
rect 15760 24699 15792 24731
rect 15832 24699 15864 24731
rect 15904 24699 15936 24731
rect 64 24627 96 24659
rect 136 24627 168 24659
rect 208 24627 240 24659
rect 280 24627 312 24659
rect 352 24627 384 24659
rect 424 24627 456 24659
rect 496 24627 528 24659
rect 568 24627 600 24659
rect 640 24627 672 24659
rect 712 24627 744 24659
rect 784 24627 816 24659
rect 856 24627 888 24659
rect 928 24627 960 24659
rect 1000 24627 1032 24659
rect 1072 24627 1104 24659
rect 1144 24627 1176 24659
rect 1216 24627 1248 24659
rect 1288 24627 1320 24659
rect 1360 24627 1392 24659
rect 1432 24627 1464 24659
rect 1504 24627 1536 24659
rect 1576 24627 1608 24659
rect 1648 24627 1680 24659
rect 1720 24627 1752 24659
rect 1792 24627 1824 24659
rect 1864 24627 1896 24659
rect 1936 24627 1968 24659
rect 2008 24627 2040 24659
rect 2080 24627 2112 24659
rect 2152 24627 2184 24659
rect 2224 24627 2256 24659
rect 2296 24627 2328 24659
rect 2368 24627 2400 24659
rect 2440 24627 2472 24659
rect 2512 24627 2544 24659
rect 2584 24627 2616 24659
rect 2656 24627 2688 24659
rect 2728 24627 2760 24659
rect 2800 24627 2832 24659
rect 2872 24627 2904 24659
rect 2944 24627 2976 24659
rect 3016 24627 3048 24659
rect 3088 24627 3120 24659
rect 3160 24627 3192 24659
rect 3232 24627 3264 24659
rect 3304 24627 3336 24659
rect 3376 24627 3408 24659
rect 3448 24627 3480 24659
rect 3520 24627 3552 24659
rect 3592 24627 3624 24659
rect 3664 24627 3696 24659
rect 3736 24627 3768 24659
rect 3808 24627 3840 24659
rect 3880 24627 3912 24659
rect 3952 24627 3984 24659
rect 4024 24627 4056 24659
rect 4096 24627 4128 24659
rect 4168 24627 4200 24659
rect 4240 24627 4272 24659
rect 4312 24627 4344 24659
rect 4384 24627 4416 24659
rect 4456 24627 4488 24659
rect 4528 24627 4560 24659
rect 4600 24627 4632 24659
rect 4672 24627 4704 24659
rect 4744 24627 4776 24659
rect 4816 24627 4848 24659
rect 4888 24627 4920 24659
rect 4960 24627 4992 24659
rect 5032 24627 5064 24659
rect 5104 24627 5136 24659
rect 5176 24627 5208 24659
rect 5248 24627 5280 24659
rect 5320 24627 5352 24659
rect 5392 24627 5424 24659
rect 5464 24627 5496 24659
rect 5536 24627 5568 24659
rect 5608 24627 5640 24659
rect 5680 24627 5712 24659
rect 5752 24627 5784 24659
rect 5824 24627 5856 24659
rect 5896 24627 5928 24659
rect 5968 24627 6000 24659
rect 6040 24627 6072 24659
rect 6112 24627 6144 24659
rect 6184 24627 6216 24659
rect 6256 24627 6288 24659
rect 6328 24627 6360 24659
rect 6400 24627 6432 24659
rect 6472 24627 6504 24659
rect 6544 24627 6576 24659
rect 6616 24627 6648 24659
rect 6688 24627 6720 24659
rect 6760 24627 6792 24659
rect 6832 24627 6864 24659
rect 6904 24627 6936 24659
rect 6976 24627 7008 24659
rect 7048 24627 7080 24659
rect 7120 24627 7152 24659
rect 7192 24627 7224 24659
rect 7264 24627 7296 24659
rect 7336 24627 7368 24659
rect 7408 24627 7440 24659
rect 7480 24627 7512 24659
rect 7552 24627 7584 24659
rect 7624 24627 7656 24659
rect 7696 24627 7728 24659
rect 7768 24627 7800 24659
rect 7840 24627 7872 24659
rect 7912 24627 7944 24659
rect 7984 24627 8016 24659
rect 8056 24627 8088 24659
rect 8128 24627 8160 24659
rect 8200 24627 8232 24659
rect 8272 24627 8304 24659
rect 8344 24627 8376 24659
rect 8416 24627 8448 24659
rect 8488 24627 8520 24659
rect 8560 24627 8592 24659
rect 8632 24627 8664 24659
rect 8704 24627 8736 24659
rect 8776 24627 8808 24659
rect 8848 24627 8880 24659
rect 8920 24627 8952 24659
rect 8992 24627 9024 24659
rect 9064 24627 9096 24659
rect 9136 24627 9168 24659
rect 9208 24627 9240 24659
rect 9280 24627 9312 24659
rect 9352 24627 9384 24659
rect 9424 24627 9456 24659
rect 9496 24627 9528 24659
rect 9568 24627 9600 24659
rect 9640 24627 9672 24659
rect 9712 24627 9744 24659
rect 9784 24627 9816 24659
rect 9856 24627 9888 24659
rect 9928 24627 9960 24659
rect 10000 24627 10032 24659
rect 10072 24627 10104 24659
rect 10144 24627 10176 24659
rect 10216 24627 10248 24659
rect 10288 24627 10320 24659
rect 10360 24627 10392 24659
rect 10432 24627 10464 24659
rect 10504 24627 10536 24659
rect 10576 24627 10608 24659
rect 10648 24627 10680 24659
rect 10720 24627 10752 24659
rect 10792 24627 10824 24659
rect 10864 24627 10896 24659
rect 10936 24627 10968 24659
rect 11008 24627 11040 24659
rect 11080 24627 11112 24659
rect 11152 24627 11184 24659
rect 11224 24627 11256 24659
rect 11296 24627 11328 24659
rect 11368 24627 11400 24659
rect 11440 24627 11472 24659
rect 11512 24627 11544 24659
rect 11584 24627 11616 24659
rect 11656 24627 11688 24659
rect 11728 24627 11760 24659
rect 11800 24627 11832 24659
rect 11872 24627 11904 24659
rect 11944 24627 11976 24659
rect 12016 24627 12048 24659
rect 12088 24627 12120 24659
rect 12160 24627 12192 24659
rect 12232 24627 12264 24659
rect 12304 24627 12336 24659
rect 12376 24627 12408 24659
rect 12448 24627 12480 24659
rect 12520 24627 12552 24659
rect 12592 24627 12624 24659
rect 12664 24627 12696 24659
rect 12736 24627 12768 24659
rect 12808 24627 12840 24659
rect 12880 24627 12912 24659
rect 12952 24627 12984 24659
rect 13024 24627 13056 24659
rect 13096 24627 13128 24659
rect 13168 24627 13200 24659
rect 13240 24627 13272 24659
rect 13312 24627 13344 24659
rect 13384 24627 13416 24659
rect 13456 24627 13488 24659
rect 13528 24627 13560 24659
rect 13600 24627 13632 24659
rect 13672 24627 13704 24659
rect 13744 24627 13776 24659
rect 13816 24627 13848 24659
rect 13888 24627 13920 24659
rect 13960 24627 13992 24659
rect 14032 24627 14064 24659
rect 14104 24627 14136 24659
rect 14176 24627 14208 24659
rect 14248 24627 14280 24659
rect 14320 24627 14352 24659
rect 14392 24627 14424 24659
rect 14464 24627 14496 24659
rect 14536 24627 14568 24659
rect 14608 24627 14640 24659
rect 14680 24627 14712 24659
rect 14752 24627 14784 24659
rect 14824 24627 14856 24659
rect 14896 24627 14928 24659
rect 14968 24627 15000 24659
rect 15040 24627 15072 24659
rect 15112 24627 15144 24659
rect 15184 24627 15216 24659
rect 15256 24627 15288 24659
rect 15328 24627 15360 24659
rect 15400 24627 15432 24659
rect 15472 24627 15504 24659
rect 15544 24627 15576 24659
rect 15616 24627 15648 24659
rect 15688 24627 15720 24659
rect 15760 24627 15792 24659
rect 15832 24627 15864 24659
rect 15904 24627 15936 24659
rect 64 24555 96 24587
rect 136 24555 168 24587
rect 208 24555 240 24587
rect 280 24555 312 24587
rect 352 24555 384 24587
rect 424 24555 456 24587
rect 496 24555 528 24587
rect 568 24555 600 24587
rect 640 24555 672 24587
rect 712 24555 744 24587
rect 784 24555 816 24587
rect 856 24555 888 24587
rect 928 24555 960 24587
rect 1000 24555 1032 24587
rect 1072 24555 1104 24587
rect 1144 24555 1176 24587
rect 1216 24555 1248 24587
rect 1288 24555 1320 24587
rect 1360 24555 1392 24587
rect 1432 24555 1464 24587
rect 1504 24555 1536 24587
rect 1576 24555 1608 24587
rect 1648 24555 1680 24587
rect 1720 24555 1752 24587
rect 1792 24555 1824 24587
rect 1864 24555 1896 24587
rect 1936 24555 1968 24587
rect 2008 24555 2040 24587
rect 2080 24555 2112 24587
rect 2152 24555 2184 24587
rect 2224 24555 2256 24587
rect 2296 24555 2328 24587
rect 2368 24555 2400 24587
rect 2440 24555 2472 24587
rect 2512 24555 2544 24587
rect 2584 24555 2616 24587
rect 2656 24555 2688 24587
rect 2728 24555 2760 24587
rect 2800 24555 2832 24587
rect 2872 24555 2904 24587
rect 2944 24555 2976 24587
rect 3016 24555 3048 24587
rect 3088 24555 3120 24587
rect 3160 24555 3192 24587
rect 3232 24555 3264 24587
rect 3304 24555 3336 24587
rect 3376 24555 3408 24587
rect 3448 24555 3480 24587
rect 3520 24555 3552 24587
rect 3592 24555 3624 24587
rect 3664 24555 3696 24587
rect 3736 24555 3768 24587
rect 3808 24555 3840 24587
rect 3880 24555 3912 24587
rect 3952 24555 3984 24587
rect 4024 24555 4056 24587
rect 4096 24555 4128 24587
rect 4168 24555 4200 24587
rect 4240 24555 4272 24587
rect 4312 24555 4344 24587
rect 4384 24555 4416 24587
rect 4456 24555 4488 24587
rect 4528 24555 4560 24587
rect 4600 24555 4632 24587
rect 4672 24555 4704 24587
rect 4744 24555 4776 24587
rect 4816 24555 4848 24587
rect 4888 24555 4920 24587
rect 4960 24555 4992 24587
rect 5032 24555 5064 24587
rect 5104 24555 5136 24587
rect 5176 24555 5208 24587
rect 5248 24555 5280 24587
rect 5320 24555 5352 24587
rect 5392 24555 5424 24587
rect 5464 24555 5496 24587
rect 5536 24555 5568 24587
rect 5608 24555 5640 24587
rect 5680 24555 5712 24587
rect 5752 24555 5784 24587
rect 5824 24555 5856 24587
rect 5896 24555 5928 24587
rect 5968 24555 6000 24587
rect 6040 24555 6072 24587
rect 6112 24555 6144 24587
rect 6184 24555 6216 24587
rect 6256 24555 6288 24587
rect 6328 24555 6360 24587
rect 6400 24555 6432 24587
rect 6472 24555 6504 24587
rect 6544 24555 6576 24587
rect 6616 24555 6648 24587
rect 6688 24555 6720 24587
rect 6760 24555 6792 24587
rect 6832 24555 6864 24587
rect 6904 24555 6936 24587
rect 6976 24555 7008 24587
rect 7048 24555 7080 24587
rect 7120 24555 7152 24587
rect 7192 24555 7224 24587
rect 7264 24555 7296 24587
rect 7336 24555 7368 24587
rect 7408 24555 7440 24587
rect 7480 24555 7512 24587
rect 7552 24555 7584 24587
rect 7624 24555 7656 24587
rect 7696 24555 7728 24587
rect 7768 24555 7800 24587
rect 7840 24555 7872 24587
rect 7912 24555 7944 24587
rect 7984 24555 8016 24587
rect 8056 24555 8088 24587
rect 8128 24555 8160 24587
rect 8200 24555 8232 24587
rect 8272 24555 8304 24587
rect 8344 24555 8376 24587
rect 8416 24555 8448 24587
rect 8488 24555 8520 24587
rect 8560 24555 8592 24587
rect 8632 24555 8664 24587
rect 8704 24555 8736 24587
rect 8776 24555 8808 24587
rect 8848 24555 8880 24587
rect 8920 24555 8952 24587
rect 8992 24555 9024 24587
rect 9064 24555 9096 24587
rect 9136 24555 9168 24587
rect 9208 24555 9240 24587
rect 9280 24555 9312 24587
rect 9352 24555 9384 24587
rect 9424 24555 9456 24587
rect 9496 24555 9528 24587
rect 9568 24555 9600 24587
rect 9640 24555 9672 24587
rect 9712 24555 9744 24587
rect 9784 24555 9816 24587
rect 9856 24555 9888 24587
rect 9928 24555 9960 24587
rect 10000 24555 10032 24587
rect 10072 24555 10104 24587
rect 10144 24555 10176 24587
rect 10216 24555 10248 24587
rect 10288 24555 10320 24587
rect 10360 24555 10392 24587
rect 10432 24555 10464 24587
rect 10504 24555 10536 24587
rect 10576 24555 10608 24587
rect 10648 24555 10680 24587
rect 10720 24555 10752 24587
rect 10792 24555 10824 24587
rect 10864 24555 10896 24587
rect 10936 24555 10968 24587
rect 11008 24555 11040 24587
rect 11080 24555 11112 24587
rect 11152 24555 11184 24587
rect 11224 24555 11256 24587
rect 11296 24555 11328 24587
rect 11368 24555 11400 24587
rect 11440 24555 11472 24587
rect 11512 24555 11544 24587
rect 11584 24555 11616 24587
rect 11656 24555 11688 24587
rect 11728 24555 11760 24587
rect 11800 24555 11832 24587
rect 11872 24555 11904 24587
rect 11944 24555 11976 24587
rect 12016 24555 12048 24587
rect 12088 24555 12120 24587
rect 12160 24555 12192 24587
rect 12232 24555 12264 24587
rect 12304 24555 12336 24587
rect 12376 24555 12408 24587
rect 12448 24555 12480 24587
rect 12520 24555 12552 24587
rect 12592 24555 12624 24587
rect 12664 24555 12696 24587
rect 12736 24555 12768 24587
rect 12808 24555 12840 24587
rect 12880 24555 12912 24587
rect 12952 24555 12984 24587
rect 13024 24555 13056 24587
rect 13096 24555 13128 24587
rect 13168 24555 13200 24587
rect 13240 24555 13272 24587
rect 13312 24555 13344 24587
rect 13384 24555 13416 24587
rect 13456 24555 13488 24587
rect 13528 24555 13560 24587
rect 13600 24555 13632 24587
rect 13672 24555 13704 24587
rect 13744 24555 13776 24587
rect 13816 24555 13848 24587
rect 13888 24555 13920 24587
rect 13960 24555 13992 24587
rect 14032 24555 14064 24587
rect 14104 24555 14136 24587
rect 14176 24555 14208 24587
rect 14248 24555 14280 24587
rect 14320 24555 14352 24587
rect 14392 24555 14424 24587
rect 14464 24555 14496 24587
rect 14536 24555 14568 24587
rect 14608 24555 14640 24587
rect 14680 24555 14712 24587
rect 14752 24555 14784 24587
rect 14824 24555 14856 24587
rect 14896 24555 14928 24587
rect 14968 24555 15000 24587
rect 15040 24555 15072 24587
rect 15112 24555 15144 24587
rect 15184 24555 15216 24587
rect 15256 24555 15288 24587
rect 15328 24555 15360 24587
rect 15400 24555 15432 24587
rect 15472 24555 15504 24587
rect 15544 24555 15576 24587
rect 15616 24555 15648 24587
rect 15688 24555 15720 24587
rect 15760 24555 15792 24587
rect 15832 24555 15864 24587
rect 15904 24555 15936 24587
rect 64 24483 96 24515
rect 136 24483 168 24515
rect 208 24483 240 24515
rect 280 24483 312 24515
rect 352 24483 384 24515
rect 424 24483 456 24515
rect 496 24483 528 24515
rect 568 24483 600 24515
rect 640 24483 672 24515
rect 712 24483 744 24515
rect 784 24483 816 24515
rect 856 24483 888 24515
rect 928 24483 960 24515
rect 1000 24483 1032 24515
rect 1072 24483 1104 24515
rect 1144 24483 1176 24515
rect 1216 24483 1248 24515
rect 1288 24483 1320 24515
rect 1360 24483 1392 24515
rect 1432 24483 1464 24515
rect 1504 24483 1536 24515
rect 1576 24483 1608 24515
rect 1648 24483 1680 24515
rect 1720 24483 1752 24515
rect 1792 24483 1824 24515
rect 1864 24483 1896 24515
rect 1936 24483 1968 24515
rect 2008 24483 2040 24515
rect 2080 24483 2112 24515
rect 2152 24483 2184 24515
rect 2224 24483 2256 24515
rect 2296 24483 2328 24515
rect 2368 24483 2400 24515
rect 2440 24483 2472 24515
rect 2512 24483 2544 24515
rect 2584 24483 2616 24515
rect 2656 24483 2688 24515
rect 2728 24483 2760 24515
rect 2800 24483 2832 24515
rect 2872 24483 2904 24515
rect 2944 24483 2976 24515
rect 3016 24483 3048 24515
rect 3088 24483 3120 24515
rect 3160 24483 3192 24515
rect 3232 24483 3264 24515
rect 3304 24483 3336 24515
rect 3376 24483 3408 24515
rect 3448 24483 3480 24515
rect 3520 24483 3552 24515
rect 3592 24483 3624 24515
rect 3664 24483 3696 24515
rect 3736 24483 3768 24515
rect 3808 24483 3840 24515
rect 3880 24483 3912 24515
rect 3952 24483 3984 24515
rect 4024 24483 4056 24515
rect 4096 24483 4128 24515
rect 4168 24483 4200 24515
rect 4240 24483 4272 24515
rect 4312 24483 4344 24515
rect 4384 24483 4416 24515
rect 4456 24483 4488 24515
rect 4528 24483 4560 24515
rect 4600 24483 4632 24515
rect 4672 24483 4704 24515
rect 4744 24483 4776 24515
rect 4816 24483 4848 24515
rect 4888 24483 4920 24515
rect 4960 24483 4992 24515
rect 5032 24483 5064 24515
rect 5104 24483 5136 24515
rect 5176 24483 5208 24515
rect 5248 24483 5280 24515
rect 5320 24483 5352 24515
rect 5392 24483 5424 24515
rect 5464 24483 5496 24515
rect 5536 24483 5568 24515
rect 5608 24483 5640 24515
rect 5680 24483 5712 24515
rect 5752 24483 5784 24515
rect 5824 24483 5856 24515
rect 5896 24483 5928 24515
rect 5968 24483 6000 24515
rect 6040 24483 6072 24515
rect 6112 24483 6144 24515
rect 6184 24483 6216 24515
rect 6256 24483 6288 24515
rect 6328 24483 6360 24515
rect 6400 24483 6432 24515
rect 6472 24483 6504 24515
rect 6544 24483 6576 24515
rect 6616 24483 6648 24515
rect 6688 24483 6720 24515
rect 6760 24483 6792 24515
rect 6832 24483 6864 24515
rect 6904 24483 6936 24515
rect 6976 24483 7008 24515
rect 7048 24483 7080 24515
rect 7120 24483 7152 24515
rect 7192 24483 7224 24515
rect 7264 24483 7296 24515
rect 7336 24483 7368 24515
rect 7408 24483 7440 24515
rect 7480 24483 7512 24515
rect 7552 24483 7584 24515
rect 7624 24483 7656 24515
rect 7696 24483 7728 24515
rect 7768 24483 7800 24515
rect 7840 24483 7872 24515
rect 7912 24483 7944 24515
rect 7984 24483 8016 24515
rect 8056 24483 8088 24515
rect 8128 24483 8160 24515
rect 8200 24483 8232 24515
rect 8272 24483 8304 24515
rect 8344 24483 8376 24515
rect 8416 24483 8448 24515
rect 8488 24483 8520 24515
rect 8560 24483 8592 24515
rect 8632 24483 8664 24515
rect 8704 24483 8736 24515
rect 8776 24483 8808 24515
rect 8848 24483 8880 24515
rect 8920 24483 8952 24515
rect 8992 24483 9024 24515
rect 9064 24483 9096 24515
rect 9136 24483 9168 24515
rect 9208 24483 9240 24515
rect 9280 24483 9312 24515
rect 9352 24483 9384 24515
rect 9424 24483 9456 24515
rect 9496 24483 9528 24515
rect 9568 24483 9600 24515
rect 9640 24483 9672 24515
rect 9712 24483 9744 24515
rect 9784 24483 9816 24515
rect 9856 24483 9888 24515
rect 9928 24483 9960 24515
rect 10000 24483 10032 24515
rect 10072 24483 10104 24515
rect 10144 24483 10176 24515
rect 10216 24483 10248 24515
rect 10288 24483 10320 24515
rect 10360 24483 10392 24515
rect 10432 24483 10464 24515
rect 10504 24483 10536 24515
rect 10576 24483 10608 24515
rect 10648 24483 10680 24515
rect 10720 24483 10752 24515
rect 10792 24483 10824 24515
rect 10864 24483 10896 24515
rect 10936 24483 10968 24515
rect 11008 24483 11040 24515
rect 11080 24483 11112 24515
rect 11152 24483 11184 24515
rect 11224 24483 11256 24515
rect 11296 24483 11328 24515
rect 11368 24483 11400 24515
rect 11440 24483 11472 24515
rect 11512 24483 11544 24515
rect 11584 24483 11616 24515
rect 11656 24483 11688 24515
rect 11728 24483 11760 24515
rect 11800 24483 11832 24515
rect 11872 24483 11904 24515
rect 11944 24483 11976 24515
rect 12016 24483 12048 24515
rect 12088 24483 12120 24515
rect 12160 24483 12192 24515
rect 12232 24483 12264 24515
rect 12304 24483 12336 24515
rect 12376 24483 12408 24515
rect 12448 24483 12480 24515
rect 12520 24483 12552 24515
rect 12592 24483 12624 24515
rect 12664 24483 12696 24515
rect 12736 24483 12768 24515
rect 12808 24483 12840 24515
rect 12880 24483 12912 24515
rect 12952 24483 12984 24515
rect 13024 24483 13056 24515
rect 13096 24483 13128 24515
rect 13168 24483 13200 24515
rect 13240 24483 13272 24515
rect 13312 24483 13344 24515
rect 13384 24483 13416 24515
rect 13456 24483 13488 24515
rect 13528 24483 13560 24515
rect 13600 24483 13632 24515
rect 13672 24483 13704 24515
rect 13744 24483 13776 24515
rect 13816 24483 13848 24515
rect 13888 24483 13920 24515
rect 13960 24483 13992 24515
rect 14032 24483 14064 24515
rect 14104 24483 14136 24515
rect 14176 24483 14208 24515
rect 14248 24483 14280 24515
rect 14320 24483 14352 24515
rect 14392 24483 14424 24515
rect 14464 24483 14496 24515
rect 14536 24483 14568 24515
rect 14608 24483 14640 24515
rect 14680 24483 14712 24515
rect 14752 24483 14784 24515
rect 14824 24483 14856 24515
rect 14896 24483 14928 24515
rect 14968 24483 15000 24515
rect 15040 24483 15072 24515
rect 15112 24483 15144 24515
rect 15184 24483 15216 24515
rect 15256 24483 15288 24515
rect 15328 24483 15360 24515
rect 15400 24483 15432 24515
rect 15472 24483 15504 24515
rect 15544 24483 15576 24515
rect 15616 24483 15648 24515
rect 15688 24483 15720 24515
rect 15760 24483 15792 24515
rect 15832 24483 15864 24515
rect 15904 24483 15936 24515
rect 64 24411 96 24443
rect 136 24411 168 24443
rect 208 24411 240 24443
rect 280 24411 312 24443
rect 352 24411 384 24443
rect 424 24411 456 24443
rect 496 24411 528 24443
rect 568 24411 600 24443
rect 640 24411 672 24443
rect 712 24411 744 24443
rect 784 24411 816 24443
rect 856 24411 888 24443
rect 928 24411 960 24443
rect 1000 24411 1032 24443
rect 1072 24411 1104 24443
rect 1144 24411 1176 24443
rect 1216 24411 1248 24443
rect 1288 24411 1320 24443
rect 1360 24411 1392 24443
rect 1432 24411 1464 24443
rect 1504 24411 1536 24443
rect 1576 24411 1608 24443
rect 1648 24411 1680 24443
rect 1720 24411 1752 24443
rect 1792 24411 1824 24443
rect 1864 24411 1896 24443
rect 1936 24411 1968 24443
rect 2008 24411 2040 24443
rect 2080 24411 2112 24443
rect 2152 24411 2184 24443
rect 2224 24411 2256 24443
rect 2296 24411 2328 24443
rect 2368 24411 2400 24443
rect 2440 24411 2472 24443
rect 2512 24411 2544 24443
rect 2584 24411 2616 24443
rect 2656 24411 2688 24443
rect 2728 24411 2760 24443
rect 2800 24411 2832 24443
rect 2872 24411 2904 24443
rect 2944 24411 2976 24443
rect 3016 24411 3048 24443
rect 3088 24411 3120 24443
rect 3160 24411 3192 24443
rect 3232 24411 3264 24443
rect 3304 24411 3336 24443
rect 3376 24411 3408 24443
rect 3448 24411 3480 24443
rect 3520 24411 3552 24443
rect 3592 24411 3624 24443
rect 3664 24411 3696 24443
rect 3736 24411 3768 24443
rect 3808 24411 3840 24443
rect 3880 24411 3912 24443
rect 3952 24411 3984 24443
rect 4024 24411 4056 24443
rect 4096 24411 4128 24443
rect 4168 24411 4200 24443
rect 4240 24411 4272 24443
rect 4312 24411 4344 24443
rect 4384 24411 4416 24443
rect 4456 24411 4488 24443
rect 4528 24411 4560 24443
rect 4600 24411 4632 24443
rect 4672 24411 4704 24443
rect 4744 24411 4776 24443
rect 4816 24411 4848 24443
rect 4888 24411 4920 24443
rect 4960 24411 4992 24443
rect 5032 24411 5064 24443
rect 5104 24411 5136 24443
rect 5176 24411 5208 24443
rect 5248 24411 5280 24443
rect 5320 24411 5352 24443
rect 5392 24411 5424 24443
rect 5464 24411 5496 24443
rect 5536 24411 5568 24443
rect 5608 24411 5640 24443
rect 5680 24411 5712 24443
rect 5752 24411 5784 24443
rect 5824 24411 5856 24443
rect 5896 24411 5928 24443
rect 5968 24411 6000 24443
rect 6040 24411 6072 24443
rect 6112 24411 6144 24443
rect 6184 24411 6216 24443
rect 6256 24411 6288 24443
rect 6328 24411 6360 24443
rect 6400 24411 6432 24443
rect 6472 24411 6504 24443
rect 6544 24411 6576 24443
rect 6616 24411 6648 24443
rect 6688 24411 6720 24443
rect 6760 24411 6792 24443
rect 6832 24411 6864 24443
rect 6904 24411 6936 24443
rect 6976 24411 7008 24443
rect 7048 24411 7080 24443
rect 7120 24411 7152 24443
rect 7192 24411 7224 24443
rect 7264 24411 7296 24443
rect 7336 24411 7368 24443
rect 7408 24411 7440 24443
rect 7480 24411 7512 24443
rect 7552 24411 7584 24443
rect 7624 24411 7656 24443
rect 7696 24411 7728 24443
rect 7768 24411 7800 24443
rect 7840 24411 7872 24443
rect 7912 24411 7944 24443
rect 7984 24411 8016 24443
rect 8056 24411 8088 24443
rect 8128 24411 8160 24443
rect 8200 24411 8232 24443
rect 8272 24411 8304 24443
rect 8344 24411 8376 24443
rect 8416 24411 8448 24443
rect 8488 24411 8520 24443
rect 8560 24411 8592 24443
rect 8632 24411 8664 24443
rect 8704 24411 8736 24443
rect 8776 24411 8808 24443
rect 8848 24411 8880 24443
rect 8920 24411 8952 24443
rect 8992 24411 9024 24443
rect 9064 24411 9096 24443
rect 9136 24411 9168 24443
rect 9208 24411 9240 24443
rect 9280 24411 9312 24443
rect 9352 24411 9384 24443
rect 9424 24411 9456 24443
rect 9496 24411 9528 24443
rect 9568 24411 9600 24443
rect 9640 24411 9672 24443
rect 9712 24411 9744 24443
rect 9784 24411 9816 24443
rect 9856 24411 9888 24443
rect 9928 24411 9960 24443
rect 10000 24411 10032 24443
rect 10072 24411 10104 24443
rect 10144 24411 10176 24443
rect 10216 24411 10248 24443
rect 10288 24411 10320 24443
rect 10360 24411 10392 24443
rect 10432 24411 10464 24443
rect 10504 24411 10536 24443
rect 10576 24411 10608 24443
rect 10648 24411 10680 24443
rect 10720 24411 10752 24443
rect 10792 24411 10824 24443
rect 10864 24411 10896 24443
rect 10936 24411 10968 24443
rect 11008 24411 11040 24443
rect 11080 24411 11112 24443
rect 11152 24411 11184 24443
rect 11224 24411 11256 24443
rect 11296 24411 11328 24443
rect 11368 24411 11400 24443
rect 11440 24411 11472 24443
rect 11512 24411 11544 24443
rect 11584 24411 11616 24443
rect 11656 24411 11688 24443
rect 11728 24411 11760 24443
rect 11800 24411 11832 24443
rect 11872 24411 11904 24443
rect 11944 24411 11976 24443
rect 12016 24411 12048 24443
rect 12088 24411 12120 24443
rect 12160 24411 12192 24443
rect 12232 24411 12264 24443
rect 12304 24411 12336 24443
rect 12376 24411 12408 24443
rect 12448 24411 12480 24443
rect 12520 24411 12552 24443
rect 12592 24411 12624 24443
rect 12664 24411 12696 24443
rect 12736 24411 12768 24443
rect 12808 24411 12840 24443
rect 12880 24411 12912 24443
rect 12952 24411 12984 24443
rect 13024 24411 13056 24443
rect 13096 24411 13128 24443
rect 13168 24411 13200 24443
rect 13240 24411 13272 24443
rect 13312 24411 13344 24443
rect 13384 24411 13416 24443
rect 13456 24411 13488 24443
rect 13528 24411 13560 24443
rect 13600 24411 13632 24443
rect 13672 24411 13704 24443
rect 13744 24411 13776 24443
rect 13816 24411 13848 24443
rect 13888 24411 13920 24443
rect 13960 24411 13992 24443
rect 14032 24411 14064 24443
rect 14104 24411 14136 24443
rect 14176 24411 14208 24443
rect 14248 24411 14280 24443
rect 14320 24411 14352 24443
rect 14392 24411 14424 24443
rect 14464 24411 14496 24443
rect 14536 24411 14568 24443
rect 14608 24411 14640 24443
rect 14680 24411 14712 24443
rect 14752 24411 14784 24443
rect 14824 24411 14856 24443
rect 14896 24411 14928 24443
rect 14968 24411 15000 24443
rect 15040 24411 15072 24443
rect 15112 24411 15144 24443
rect 15184 24411 15216 24443
rect 15256 24411 15288 24443
rect 15328 24411 15360 24443
rect 15400 24411 15432 24443
rect 15472 24411 15504 24443
rect 15544 24411 15576 24443
rect 15616 24411 15648 24443
rect 15688 24411 15720 24443
rect 15760 24411 15792 24443
rect 15832 24411 15864 24443
rect 15904 24411 15936 24443
rect 64 24339 96 24371
rect 136 24339 168 24371
rect 208 24339 240 24371
rect 280 24339 312 24371
rect 352 24339 384 24371
rect 424 24339 456 24371
rect 496 24339 528 24371
rect 568 24339 600 24371
rect 640 24339 672 24371
rect 712 24339 744 24371
rect 784 24339 816 24371
rect 856 24339 888 24371
rect 928 24339 960 24371
rect 1000 24339 1032 24371
rect 1072 24339 1104 24371
rect 1144 24339 1176 24371
rect 1216 24339 1248 24371
rect 1288 24339 1320 24371
rect 1360 24339 1392 24371
rect 1432 24339 1464 24371
rect 1504 24339 1536 24371
rect 1576 24339 1608 24371
rect 1648 24339 1680 24371
rect 1720 24339 1752 24371
rect 1792 24339 1824 24371
rect 1864 24339 1896 24371
rect 1936 24339 1968 24371
rect 2008 24339 2040 24371
rect 2080 24339 2112 24371
rect 2152 24339 2184 24371
rect 2224 24339 2256 24371
rect 2296 24339 2328 24371
rect 2368 24339 2400 24371
rect 2440 24339 2472 24371
rect 2512 24339 2544 24371
rect 2584 24339 2616 24371
rect 2656 24339 2688 24371
rect 2728 24339 2760 24371
rect 2800 24339 2832 24371
rect 2872 24339 2904 24371
rect 2944 24339 2976 24371
rect 3016 24339 3048 24371
rect 3088 24339 3120 24371
rect 3160 24339 3192 24371
rect 3232 24339 3264 24371
rect 3304 24339 3336 24371
rect 3376 24339 3408 24371
rect 3448 24339 3480 24371
rect 3520 24339 3552 24371
rect 3592 24339 3624 24371
rect 3664 24339 3696 24371
rect 3736 24339 3768 24371
rect 3808 24339 3840 24371
rect 3880 24339 3912 24371
rect 3952 24339 3984 24371
rect 4024 24339 4056 24371
rect 4096 24339 4128 24371
rect 4168 24339 4200 24371
rect 4240 24339 4272 24371
rect 4312 24339 4344 24371
rect 4384 24339 4416 24371
rect 4456 24339 4488 24371
rect 4528 24339 4560 24371
rect 4600 24339 4632 24371
rect 4672 24339 4704 24371
rect 4744 24339 4776 24371
rect 4816 24339 4848 24371
rect 4888 24339 4920 24371
rect 4960 24339 4992 24371
rect 5032 24339 5064 24371
rect 5104 24339 5136 24371
rect 5176 24339 5208 24371
rect 5248 24339 5280 24371
rect 5320 24339 5352 24371
rect 5392 24339 5424 24371
rect 5464 24339 5496 24371
rect 5536 24339 5568 24371
rect 5608 24339 5640 24371
rect 5680 24339 5712 24371
rect 5752 24339 5784 24371
rect 5824 24339 5856 24371
rect 5896 24339 5928 24371
rect 5968 24339 6000 24371
rect 6040 24339 6072 24371
rect 6112 24339 6144 24371
rect 6184 24339 6216 24371
rect 6256 24339 6288 24371
rect 6328 24339 6360 24371
rect 6400 24339 6432 24371
rect 6472 24339 6504 24371
rect 6544 24339 6576 24371
rect 6616 24339 6648 24371
rect 6688 24339 6720 24371
rect 6760 24339 6792 24371
rect 6832 24339 6864 24371
rect 6904 24339 6936 24371
rect 6976 24339 7008 24371
rect 7048 24339 7080 24371
rect 7120 24339 7152 24371
rect 7192 24339 7224 24371
rect 7264 24339 7296 24371
rect 7336 24339 7368 24371
rect 7408 24339 7440 24371
rect 7480 24339 7512 24371
rect 7552 24339 7584 24371
rect 7624 24339 7656 24371
rect 7696 24339 7728 24371
rect 7768 24339 7800 24371
rect 7840 24339 7872 24371
rect 7912 24339 7944 24371
rect 7984 24339 8016 24371
rect 8056 24339 8088 24371
rect 8128 24339 8160 24371
rect 8200 24339 8232 24371
rect 8272 24339 8304 24371
rect 8344 24339 8376 24371
rect 8416 24339 8448 24371
rect 8488 24339 8520 24371
rect 8560 24339 8592 24371
rect 8632 24339 8664 24371
rect 8704 24339 8736 24371
rect 8776 24339 8808 24371
rect 8848 24339 8880 24371
rect 8920 24339 8952 24371
rect 8992 24339 9024 24371
rect 9064 24339 9096 24371
rect 9136 24339 9168 24371
rect 9208 24339 9240 24371
rect 9280 24339 9312 24371
rect 9352 24339 9384 24371
rect 9424 24339 9456 24371
rect 9496 24339 9528 24371
rect 9568 24339 9600 24371
rect 9640 24339 9672 24371
rect 9712 24339 9744 24371
rect 9784 24339 9816 24371
rect 9856 24339 9888 24371
rect 9928 24339 9960 24371
rect 10000 24339 10032 24371
rect 10072 24339 10104 24371
rect 10144 24339 10176 24371
rect 10216 24339 10248 24371
rect 10288 24339 10320 24371
rect 10360 24339 10392 24371
rect 10432 24339 10464 24371
rect 10504 24339 10536 24371
rect 10576 24339 10608 24371
rect 10648 24339 10680 24371
rect 10720 24339 10752 24371
rect 10792 24339 10824 24371
rect 10864 24339 10896 24371
rect 10936 24339 10968 24371
rect 11008 24339 11040 24371
rect 11080 24339 11112 24371
rect 11152 24339 11184 24371
rect 11224 24339 11256 24371
rect 11296 24339 11328 24371
rect 11368 24339 11400 24371
rect 11440 24339 11472 24371
rect 11512 24339 11544 24371
rect 11584 24339 11616 24371
rect 11656 24339 11688 24371
rect 11728 24339 11760 24371
rect 11800 24339 11832 24371
rect 11872 24339 11904 24371
rect 11944 24339 11976 24371
rect 12016 24339 12048 24371
rect 12088 24339 12120 24371
rect 12160 24339 12192 24371
rect 12232 24339 12264 24371
rect 12304 24339 12336 24371
rect 12376 24339 12408 24371
rect 12448 24339 12480 24371
rect 12520 24339 12552 24371
rect 12592 24339 12624 24371
rect 12664 24339 12696 24371
rect 12736 24339 12768 24371
rect 12808 24339 12840 24371
rect 12880 24339 12912 24371
rect 12952 24339 12984 24371
rect 13024 24339 13056 24371
rect 13096 24339 13128 24371
rect 13168 24339 13200 24371
rect 13240 24339 13272 24371
rect 13312 24339 13344 24371
rect 13384 24339 13416 24371
rect 13456 24339 13488 24371
rect 13528 24339 13560 24371
rect 13600 24339 13632 24371
rect 13672 24339 13704 24371
rect 13744 24339 13776 24371
rect 13816 24339 13848 24371
rect 13888 24339 13920 24371
rect 13960 24339 13992 24371
rect 14032 24339 14064 24371
rect 14104 24339 14136 24371
rect 14176 24339 14208 24371
rect 14248 24339 14280 24371
rect 14320 24339 14352 24371
rect 14392 24339 14424 24371
rect 14464 24339 14496 24371
rect 14536 24339 14568 24371
rect 14608 24339 14640 24371
rect 14680 24339 14712 24371
rect 14752 24339 14784 24371
rect 14824 24339 14856 24371
rect 14896 24339 14928 24371
rect 14968 24339 15000 24371
rect 15040 24339 15072 24371
rect 15112 24339 15144 24371
rect 15184 24339 15216 24371
rect 15256 24339 15288 24371
rect 15328 24339 15360 24371
rect 15400 24339 15432 24371
rect 15472 24339 15504 24371
rect 15544 24339 15576 24371
rect 15616 24339 15648 24371
rect 15688 24339 15720 24371
rect 15760 24339 15792 24371
rect 15832 24339 15864 24371
rect 15904 24339 15936 24371
rect 64 24267 96 24299
rect 136 24267 168 24299
rect 208 24267 240 24299
rect 280 24267 312 24299
rect 352 24267 384 24299
rect 424 24267 456 24299
rect 496 24267 528 24299
rect 568 24267 600 24299
rect 640 24267 672 24299
rect 712 24267 744 24299
rect 784 24267 816 24299
rect 856 24267 888 24299
rect 928 24267 960 24299
rect 1000 24267 1032 24299
rect 1072 24267 1104 24299
rect 1144 24267 1176 24299
rect 1216 24267 1248 24299
rect 1288 24267 1320 24299
rect 1360 24267 1392 24299
rect 1432 24267 1464 24299
rect 1504 24267 1536 24299
rect 1576 24267 1608 24299
rect 1648 24267 1680 24299
rect 1720 24267 1752 24299
rect 1792 24267 1824 24299
rect 1864 24267 1896 24299
rect 1936 24267 1968 24299
rect 2008 24267 2040 24299
rect 2080 24267 2112 24299
rect 2152 24267 2184 24299
rect 2224 24267 2256 24299
rect 2296 24267 2328 24299
rect 2368 24267 2400 24299
rect 2440 24267 2472 24299
rect 2512 24267 2544 24299
rect 2584 24267 2616 24299
rect 2656 24267 2688 24299
rect 2728 24267 2760 24299
rect 2800 24267 2832 24299
rect 2872 24267 2904 24299
rect 2944 24267 2976 24299
rect 3016 24267 3048 24299
rect 3088 24267 3120 24299
rect 3160 24267 3192 24299
rect 3232 24267 3264 24299
rect 3304 24267 3336 24299
rect 3376 24267 3408 24299
rect 3448 24267 3480 24299
rect 3520 24267 3552 24299
rect 3592 24267 3624 24299
rect 3664 24267 3696 24299
rect 3736 24267 3768 24299
rect 3808 24267 3840 24299
rect 3880 24267 3912 24299
rect 3952 24267 3984 24299
rect 4024 24267 4056 24299
rect 4096 24267 4128 24299
rect 4168 24267 4200 24299
rect 4240 24267 4272 24299
rect 4312 24267 4344 24299
rect 4384 24267 4416 24299
rect 4456 24267 4488 24299
rect 4528 24267 4560 24299
rect 4600 24267 4632 24299
rect 4672 24267 4704 24299
rect 4744 24267 4776 24299
rect 4816 24267 4848 24299
rect 4888 24267 4920 24299
rect 4960 24267 4992 24299
rect 5032 24267 5064 24299
rect 5104 24267 5136 24299
rect 5176 24267 5208 24299
rect 5248 24267 5280 24299
rect 5320 24267 5352 24299
rect 5392 24267 5424 24299
rect 5464 24267 5496 24299
rect 5536 24267 5568 24299
rect 5608 24267 5640 24299
rect 5680 24267 5712 24299
rect 5752 24267 5784 24299
rect 5824 24267 5856 24299
rect 5896 24267 5928 24299
rect 5968 24267 6000 24299
rect 6040 24267 6072 24299
rect 6112 24267 6144 24299
rect 6184 24267 6216 24299
rect 6256 24267 6288 24299
rect 6328 24267 6360 24299
rect 6400 24267 6432 24299
rect 6472 24267 6504 24299
rect 6544 24267 6576 24299
rect 6616 24267 6648 24299
rect 6688 24267 6720 24299
rect 6760 24267 6792 24299
rect 6832 24267 6864 24299
rect 6904 24267 6936 24299
rect 6976 24267 7008 24299
rect 7048 24267 7080 24299
rect 7120 24267 7152 24299
rect 7192 24267 7224 24299
rect 7264 24267 7296 24299
rect 7336 24267 7368 24299
rect 7408 24267 7440 24299
rect 7480 24267 7512 24299
rect 7552 24267 7584 24299
rect 7624 24267 7656 24299
rect 7696 24267 7728 24299
rect 7768 24267 7800 24299
rect 7840 24267 7872 24299
rect 7912 24267 7944 24299
rect 7984 24267 8016 24299
rect 8056 24267 8088 24299
rect 8128 24267 8160 24299
rect 8200 24267 8232 24299
rect 8272 24267 8304 24299
rect 8344 24267 8376 24299
rect 8416 24267 8448 24299
rect 8488 24267 8520 24299
rect 8560 24267 8592 24299
rect 8632 24267 8664 24299
rect 8704 24267 8736 24299
rect 8776 24267 8808 24299
rect 8848 24267 8880 24299
rect 8920 24267 8952 24299
rect 8992 24267 9024 24299
rect 9064 24267 9096 24299
rect 9136 24267 9168 24299
rect 9208 24267 9240 24299
rect 9280 24267 9312 24299
rect 9352 24267 9384 24299
rect 9424 24267 9456 24299
rect 9496 24267 9528 24299
rect 9568 24267 9600 24299
rect 9640 24267 9672 24299
rect 9712 24267 9744 24299
rect 9784 24267 9816 24299
rect 9856 24267 9888 24299
rect 9928 24267 9960 24299
rect 10000 24267 10032 24299
rect 10072 24267 10104 24299
rect 10144 24267 10176 24299
rect 10216 24267 10248 24299
rect 10288 24267 10320 24299
rect 10360 24267 10392 24299
rect 10432 24267 10464 24299
rect 10504 24267 10536 24299
rect 10576 24267 10608 24299
rect 10648 24267 10680 24299
rect 10720 24267 10752 24299
rect 10792 24267 10824 24299
rect 10864 24267 10896 24299
rect 10936 24267 10968 24299
rect 11008 24267 11040 24299
rect 11080 24267 11112 24299
rect 11152 24267 11184 24299
rect 11224 24267 11256 24299
rect 11296 24267 11328 24299
rect 11368 24267 11400 24299
rect 11440 24267 11472 24299
rect 11512 24267 11544 24299
rect 11584 24267 11616 24299
rect 11656 24267 11688 24299
rect 11728 24267 11760 24299
rect 11800 24267 11832 24299
rect 11872 24267 11904 24299
rect 11944 24267 11976 24299
rect 12016 24267 12048 24299
rect 12088 24267 12120 24299
rect 12160 24267 12192 24299
rect 12232 24267 12264 24299
rect 12304 24267 12336 24299
rect 12376 24267 12408 24299
rect 12448 24267 12480 24299
rect 12520 24267 12552 24299
rect 12592 24267 12624 24299
rect 12664 24267 12696 24299
rect 12736 24267 12768 24299
rect 12808 24267 12840 24299
rect 12880 24267 12912 24299
rect 12952 24267 12984 24299
rect 13024 24267 13056 24299
rect 13096 24267 13128 24299
rect 13168 24267 13200 24299
rect 13240 24267 13272 24299
rect 13312 24267 13344 24299
rect 13384 24267 13416 24299
rect 13456 24267 13488 24299
rect 13528 24267 13560 24299
rect 13600 24267 13632 24299
rect 13672 24267 13704 24299
rect 13744 24267 13776 24299
rect 13816 24267 13848 24299
rect 13888 24267 13920 24299
rect 13960 24267 13992 24299
rect 14032 24267 14064 24299
rect 14104 24267 14136 24299
rect 14176 24267 14208 24299
rect 14248 24267 14280 24299
rect 14320 24267 14352 24299
rect 14392 24267 14424 24299
rect 14464 24267 14496 24299
rect 14536 24267 14568 24299
rect 14608 24267 14640 24299
rect 14680 24267 14712 24299
rect 14752 24267 14784 24299
rect 14824 24267 14856 24299
rect 14896 24267 14928 24299
rect 14968 24267 15000 24299
rect 15040 24267 15072 24299
rect 15112 24267 15144 24299
rect 15184 24267 15216 24299
rect 15256 24267 15288 24299
rect 15328 24267 15360 24299
rect 15400 24267 15432 24299
rect 15472 24267 15504 24299
rect 15544 24267 15576 24299
rect 15616 24267 15648 24299
rect 15688 24267 15720 24299
rect 15760 24267 15792 24299
rect 15832 24267 15864 24299
rect 15904 24267 15936 24299
rect 64 24195 96 24227
rect 136 24195 168 24227
rect 208 24195 240 24227
rect 280 24195 312 24227
rect 352 24195 384 24227
rect 424 24195 456 24227
rect 496 24195 528 24227
rect 568 24195 600 24227
rect 640 24195 672 24227
rect 712 24195 744 24227
rect 784 24195 816 24227
rect 856 24195 888 24227
rect 928 24195 960 24227
rect 1000 24195 1032 24227
rect 1072 24195 1104 24227
rect 1144 24195 1176 24227
rect 1216 24195 1248 24227
rect 1288 24195 1320 24227
rect 1360 24195 1392 24227
rect 1432 24195 1464 24227
rect 1504 24195 1536 24227
rect 1576 24195 1608 24227
rect 1648 24195 1680 24227
rect 1720 24195 1752 24227
rect 1792 24195 1824 24227
rect 1864 24195 1896 24227
rect 1936 24195 1968 24227
rect 2008 24195 2040 24227
rect 2080 24195 2112 24227
rect 2152 24195 2184 24227
rect 2224 24195 2256 24227
rect 2296 24195 2328 24227
rect 2368 24195 2400 24227
rect 2440 24195 2472 24227
rect 2512 24195 2544 24227
rect 2584 24195 2616 24227
rect 2656 24195 2688 24227
rect 2728 24195 2760 24227
rect 2800 24195 2832 24227
rect 2872 24195 2904 24227
rect 2944 24195 2976 24227
rect 3016 24195 3048 24227
rect 3088 24195 3120 24227
rect 3160 24195 3192 24227
rect 3232 24195 3264 24227
rect 3304 24195 3336 24227
rect 3376 24195 3408 24227
rect 3448 24195 3480 24227
rect 3520 24195 3552 24227
rect 3592 24195 3624 24227
rect 3664 24195 3696 24227
rect 3736 24195 3768 24227
rect 3808 24195 3840 24227
rect 3880 24195 3912 24227
rect 3952 24195 3984 24227
rect 4024 24195 4056 24227
rect 4096 24195 4128 24227
rect 4168 24195 4200 24227
rect 4240 24195 4272 24227
rect 4312 24195 4344 24227
rect 4384 24195 4416 24227
rect 4456 24195 4488 24227
rect 4528 24195 4560 24227
rect 4600 24195 4632 24227
rect 4672 24195 4704 24227
rect 4744 24195 4776 24227
rect 4816 24195 4848 24227
rect 4888 24195 4920 24227
rect 4960 24195 4992 24227
rect 5032 24195 5064 24227
rect 5104 24195 5136 24227
rect 5176 24195 5208 24227
rect 5248 24195 5280 24227
rect 5320 24195 5352 24227
rect 5392 24195 5424 24227
rect 5464 24195 5496 24227
rect 5536 24195 5568 24227
rect 5608 24195 5640 24227
rect 5680 24195 5712 24227
rect 5752 24195 5784 24227
rect 5824 24195 5856 24227
rect 5896 24195 5928 24227
rect 5968 24195 6000 24227
rect 6040 24195 6072 24227
rect 6112 24195 6144 24227
rect 6184 24195 6216 24227
rect 6256 24195 6288 24227
rect 6328 24195 6360 24227
rect 6400 24195 6432 24227
rect 6472 24195 6504 24227
rect 6544 24195 6576 24227
rect 6616 24195 6648 24227
rect 6688 24195 6720 24227
rect 6760 24195 6792 24227
rect 6832 24195 6864 24227
rect 6904 24195 6936 24227
rect 6976 24195 7008 24227
rect 7048 24195 7080 24227
rect 7120 24195 7152 24227
rect 7192 24195 7224 24227
rect 7264 24195 7296 24227
rect 7336 24195 7368 24227
rect 7408 24195 7440 24227
rect 7480 24195 7512 24227
rect 7552 24195 7584 24227
rect 7624 24195 7656 24227
rect 7696 24195 7728 24227
rect 7768 24195 7800 24227
rect 7840 24195 7872 24227
rect 7912 24195 7944 24227
rect 7984 24195 8016 24227
rect 8056 24195 8088 24227
rect 8128 24195 8160 24227
rect 8200 24195 8232 24227
rect 8272 24195 8304 24227
rect 8344 24195 8376 24227
rect 8416 24195 8448 24227
rect 8488 24195 8520 24227
rect 8560 24195 8592 24227
rect 8632 24195 8664 24227
rect 8704 24195 8736 24227
rect 8776 24195 8808 24227
rect 8848 24195 8880 24227
rect 8920 24195 8952 24227
rect 8992 24195 9024 24227
rect 9064 24195 9096 24227
rect 9136 24195 9168 24227
rect 9208 24195 9240 24227
rect 9280 24195 9312 24227
rect 9352 24195 9384 24227
rect 9424 24195 9456 24227
rect 9496 24195 9528 24227
rect 9568 24195 9600 24227
rect 9640 24195 9672 24227
rect 9712 24195 9744 24227
rect 9784 24195 9816 24227
rect 9856 24195 9888 24227
rect 9928 24195 9960 24227
rect 10000 24195 10032 24227
rect 10072 24195 10104 24227
rect 10144 24195 10176 24227
rect 10216 24195 10248 24227
rect 10288 24195 10320 24227
rect 10360 24195 10392 24227
rect 10432 24195 10464 24227
rect 10504 24195 10536 24227
rect 10576 24195 10608 24227
rect 10648 24195 10680 24227
rect 10720 24195 10752 24227
rect 10792 24195 10824 24227
rect 10864 24195 10896 24227
rect 10936 24195 10968 24227
rect 11008 24195 11040 24227
rect 11080 24195 11112 24227
rect 11152 24195 11184 24227
rect 11224 24195 11256 24227
rect 11296 24195 11328 24227
rect 11368 24195 11400 24227
rect 11440 24195 11472 24227
rect 11512 24195 11544 24227
rect 11584 24195 11616 24227
rect 11656 24195 11688 24227
rect 11728 24195 11760 24227
rect 11800 24195 11832 24227
rect 11872 24195 11904 24227
rect 11944 24195 11976 24227
rect 12016 24195 12048 24227
rect 12088 24195 12120 24227
rect 12160 24195 12192 24227
rect 12232 24195 12264 24227
rect 12304 24195 12336 24227
rect 12376 24195 12408 24227
rect 12448 24195 12480 24227
rect 12520 24195 12552 24227
rect 12592 24195 12624 24227
rect 12664 24195 12696 24227
rect 12736 24195 12768 24227
rect 12808 24195 12840 24227
rect 12880 24195 12912 24227
rect 12952 24195 12984 24227
rect 13024 24195 13056 24227
rect 13096 24195 13128 24227
rect 13168 24195 13200 24227
rect 13240 24195 13272 24227
rect 13312 24195 13344 24227
rect 13384 24195 13416 24227
rect 13456 24195 13488 24227
rect 13528 24195 13560 24227
rect 13600 24195 13632 24227
rect 13672 24195 13704 24227
rect 13744 24195 13776 24227
rect 13816 24195 13848 24227
rect 13888 24195 13920 24227
rect 13960 24195 13992 24227
rect 14032 24195 14064 24227
rect 14104 24195 14136 24227
rect 14176 24195 14208 24227
rect 14248 24195 14280 24227
rect 14320 24195 14352 24227
rect 14392 24195 14424 24227
rect 14464 24195 14496 24227
rect 14536 24195 14568 24227
rect 14608 24195 14640 24227
rect 14680 24195 14712 24227
rect 14752 24195 14784 24227
rect 14824 24195 14856 24227
rect 14896 24195 14928 24227
rect 14968 24195 15000 24227
rect 15040 24195 15072 24227
rect 15112 24195 15144 24227
rect 15184 24195 15216 24227
rect 15256 24195 15288 24227
rect 15328 24195 15360 24227
rect 15400 24195 15432 24227
rect 15472 24195 15504 24227
rect 15544 24195 15576 24227
rect 15616 24195 15648 24227
rect 15688 24195 15720 24227
rect 15760 24195 15792 24227
rect 15832 24195 15864 24227
rect 15904 24195 15936 24227
rect 64 24123 96 24155
rect 136 24123 168 24155
rect 208 24123 240 24155
rect 280 24123 312 24155
rect 352 24123 384 24155
rect 424 24123 456 24155
rect 496 24123 528 24155
rect 568 24123 600 24155
rect 640 24123 672 24155
rect 712 24123 744 24155
rect 784 24123 816 24155
rect 856 24123 888 24155
rect 928 24123 960 24155
rect 1000 24123 1032 24155
rect 1072 24123 1104 24155
rect 1144 24123 1176 24155
rect 1216 24123 1248 24155
rect 1288 24123 1320 24155
rect 1360 24123 1392 24155
rect 1432 24123 1464 24155
rect 1504 24123 1536 24155
rect 1576 24123 1608 24155
rect 1648 24123 1680 24155
rect 1720 24123 1752 24155
rect 1792 24123 1824 24155
rect 1864 24123 1896 24155
rect 1936 24123 1968 24155
rect 2008 24123 2040 24155
rect 2080 24123 2112 24155
rect 2152 24123 2184 24155
rect 2224 24123 2256 24155
rect 2296 24123 2328 24155
rect 2368 24123 2400 24155
rect 2440 24123 2472 24155
rect 2512 24123 2544 24155
rect 2584 24123 2616 24155
rect 2656 24123 2688 24155
rect 2728 24123 2760 24155
rect 2800 24123 2832 24155
rect 2872 24123 2904 24155
rect 2944 24123 2976 24155
rect 3016 24123 3048 24155
rect 3088 24123 3120 24155
rect 3160 24123 3192 24155
rect 3232 24123 3264 24155
rect 3304 24123 3336 24155
rect 3376 24123 3408 24155
rect 3448 24123 3480 24155
rect 3520 24123 3552 24155
rect 3592 24123 3624 24155
rect 3664 24123 3696 24155
rect 3736 24123 3768 24155
rect 3808 24123 3840 24155
rect 3880 24123 3912 24155
rect 3952 24123 3984 24155
rect 4024 24123 4056 24155
rect 4096 24123 4128 24155
rect 4168 24123 4200 24155
rect 4240 24123 4272 24155
rect 4312 24123 4344 24155
rect 4384 24123 4416 24155
rect 4456 24123 4488 24155
rect 4528 24123 4560 24155
rect 4600 24123 4632 24155
rect 4672 24123 4704 24155
rect 4744 24123 4776 24155
rect 4816 24123 4848 24155
rect 4888 24123 4920 24155
rect 4960 24123 4992 24155
rect 5032 24123 5064 24155
rect 5104 24123 5136 24155
rect 5176 24123 5208 24155
rect 5248 24123 5280 24155
rect 5320 24123 5352 24155
rect 5392 24123 5424 24155
rect 5464 24123 5496 24155
rect 5536 24123 5568 24155
rect 5608 24123 5640 24155
rect 5680 24123 5712 24155
rect 5752 24123 5784 24155
rect 5824 24123 5856 24155
rect 5896 24123 5928 24155
rect 5968 24123 6000 24155
rect 6040 24123 6072 24155
rect 6112 24123 6144 24155
rect 6184 24123 6216 24155
rect 6256 24123 6288 24155
rect 6328 24123 6360 24155
rect 6400 24123 6432 24155
rect 6472 24123 6504 24155
rect 6544 24123 6576 24155
rect 6616 24123 6648 24155
rect 6688 24123 6720 24155
rect 6760 24123 6792 24155
rect 6832 24123 6864 24155
rect 6904 24123 6936 24155
rect 6976 24123 7008 24155
rect 7048 24123 7080 24155
rect 7120 24123 7152 24155
rect 7192 24123 7224 24155
rect 7264 24123 7296 24155
rect 7336 24123 7368 24155
rect 7408 24123 7440 24155
rect 7480 24123 7512 24155
rect 7552 24123 7584 24155
rect 7624 24123 7656 24155
rect 7696 24123 7728 24155
rect 7768 24123 7800 24155
rect 7840 24123 7872 24155
rect 7912 24123 7944 24155
rect 7984 24123 8016 24155
rect 8056 24123 8088 24155
rect 8128 24123 8160 24155
rect 8200 24123 8232 24155
rect 8272 24123 8304 24155
rect 8344 24123 8376 24155
rect 8416 24123 8448 24155
rect 8488 24123 8520 24155
rect 8560 24123 8592 24155
rect 8632 24123 8664 24155
rect 8704 24123 8736 24155
rect 8776 24123 8808 24155
rect 8848 24123 8880 24155
rect 8920 24123 8952 24155
rect 8992 24123 9024 24155
rect 9064 24123 9096 24155
rect 9136 24123 9168 24155
rect 9208 24123 9240 24155
rect 9280 24123 9312 24155
rect 9352 24123 9384 24155
rect 9424 24123 9456 24155
rect 9496 24123 9528 24155
rect 9568 24123 9600 24155
rect 9640 24123 9672 24155
rect 9712 24123 9744 24155
rect 9784 24123 9816 24155
rect 9856 24123 9888 24155
rect 9928 24123 9960 24155
rect 10000 24123 10032 24155
rect 10072 24123 10104 24155
rect 10144 24123 10176 24155
rect 10216 24123 10248 24155
rect 10288 24123 10320 24155
rect 10360 24123 10392 24155
rect 10432 24123 10464 24155
rect 10504 24123 10536 24155
rect 10576 24123 10608 24155
rect 10648 24123 10680 24155
rect 10720 24123 10752 24155
rect 10792 24123 10824 24155
rect 10864 24123 10896 24155
rect 10936 24123 10968 24155
rect 11008 24123 11040 24155
rect 11080 24123 11112 24155
rect 11152 24123 11184 24155
rect 11224 24123 11256 24155
rect 11296 24123 11328 24155
rect 11368 24123 11400 24155
rect 11440 24123 11472 24155
rect 11512 24123 11544 24155
rect 11584 24123 11616 24155
rect 11656 24123 11688 24155
rect 11728 24123 11760 24155
rect 11800 24123 11832 24155
rect 11872 24123 11904 24155
rect 11944 24123 11976 24155
rect 12016 24123 12048 24155
rect 12088 24123 12120 24155
rect 12160 24123 12192 24155
rect 12232 24123 12264 24155
rect 12304 24123 12336 24155
rect 12376 24123 12408 24155
rect 12448 24123 12480 24155
rect 12520 24123 12552 24155
rect 12592 24123 12624 24155
rect 12664 24123 12696 24155
rect 12736 24123 12768 24155
rect 12808 24123 12840 24155
rect 12880 24123 12912 24155
rect 12952 24123 12984 24155
rect 13024 24123 13056 24155
rect 13096 24123 13128 24155
rect 13168 24123 13200 24155
rect 13240 24123 13272 24155
rect 13312 24123 13344 24155
rect 13384 24123 13416 24155
rect 13456 24123 13488 24155
rect 13528 24123 13560 24155
rect 13600 24123 13632 24155
rect 13672 24123 13704 24155
rect 13744 24123 13776 24155
rect 13816 24123 13848 24155
rect 13888 24123 13920 24155
rect 13960 24123 13992 24155
rect 14032 24123 14064 24155
rect 14104 24123 14136 24155
rect 14176 24123 14208 24155
rect 14248 24123 14280 24155
rect 14320 24123 14352 24155
rect 14392 24123 14424 24155
rect 14464 24123 14496 24155
rect 14536 24123 14568 24155
rect 14608 24123 14640 24155
rect 14680 24123 14712 24155
rect 14752 24123 14784 24155
rect 14824 24123 14856 24155
rect 14896 24123 14928 24155
rect 14968 24123 15000 24155
rect 15040 24123 15072 24155
rect 15112 24123 15144 24155
rect 15184 24123 15216 24155
rect 15256 24123 15288 24155
rect 15328 24123 15360 24155
rect 15400 24123 15432 24155
rect 15472 24123 15504 24155
rect 15544 24123 15576 24155
rect 15616 24123 15648 24155
rect 15688 24123 15720 24155
rect 15760 24123 15792 24155
rect 15832 24123 15864 24155
rect 15904 24123 15936 24155
rect 64 24051 96 24083
rect 136 24051 168 24083
rect 208 24051 240 24083
rect 280 24051 312 24083
rect 352 24051 384 24083
rect 424 24051 456 24083
rect 496 24051 528 24083
rect 568 24051 600 24083
rect 640 24051 672 24083
rect 712 24051 744 24083
rect 784 24051 816 24083
rect 856 24051 888 24083
rect 928 24051 960 24083
rect 1000 24051 1032 24083
rect 1072 24051 1104 24083
rect 1144 24051 1176 24083
rect 1216 24051 1248 24083
rect 1288 24051 1320 24083
rect 1360 24051 1392 24083
rect 1432 24051 1464 24083
rect 1504 24051 1536 24083
rect 1576 24051 1608 24083
rect 1648 24051 1680 24083
rect 1720 24051 1752 24083
rect 1792 24051 1824 24083
rect 1864 24051 1896 24083
rect 1936 24051 1968 24083
rect 2008 24051 2040 24083
rect 2080 24051 2112 24083
rect 2152 24051 2184 24083
rect 2224 24051 2256 24083
rect 2296 24051 2328 24083
rect 2368 24051 2400 24083
rect 2440 24051 2472 24083
rect 2512 24051 2544 24083
rect 2584 24051 2616 24083
rect 2656 24051 2688 24083
rect 2728 24051 2760 24083
rect 2800 24051 2832 24083
rect 2872 24051 2904 24083
rect 2944 24051 2976 24083
rect 3016 24051 3048 24083
rect 3088 24051 3120 24083
rect 3160 24051 3192 24083
rect 3232 24051 3264 24083
rect 3304 24051 3336 24083
rect 3376 24051 3408 24083
rect 3448 24051 3480 24083
rect 3520 24051 3552 24083
rect 3592 24051 3624 24083
rect 3664 24051 3696 24083
rect 3736 24051 3768 24083
rect 3808 24051 3840 24083
rect 3880 24051 3912 24083
rect 3952 24051 3984 24083
rect 4024 24051 4056 24083
rect 4096 24051 4128 24083
rect 4168 24051 4200 24083
rect 4240 24051 4272 24083
rect 4312 24051 4344 24083
rect 4384 24051 4416 24083
rect 4456 24051 4488 24083
rect 4528 24051 4560 24083
rect 4600 24051 4632 24083
rect 4672 24051 4704 24083
rect 4744 24051 4776 24083
rect 4816 24051 4848 24083
rect 4888 24051 4920 24083
rect 4960 24051 4992 24083
rect 5032 24051 5064 24083
rect 5104 24051 5136 24083
rect 5176 24051 5208 24083
rect 5248 24051 5280 24083
rect 5320 24051 5352 24083
rect 5392 24051 5424 24083
rect 5464 24051 5496 24083
rect 5536 24051 5568 24083
rect 5608 24051 5640 24083
rect 5680 24051 5712 24083
rect 5752 24051 5784 24083
rect 5824 24051 5856 24083
rect 5896 24051 5928 24083
rect 5968 24051 6000 24083
rect 6040 24051 6072 24083
rect 6112 24051 6144 24083
rect 6184 24051 6216 24083
rect 6256 24051 6288 24083
rect 6328 24051 6360 24083
rect 6400 24051 6432 24083
rect 6472 24051 6504 24083
rect 6544 24051 6576 24083
rect 6616 24051 6648 24083
rect 6688 24051 6720 24083
rect 6760 24051 6792 24083
rect 6832 24051 6864 24083
rect 6904 24051 6936 24083
rect 6976 24051 7008 24083
rect 7048 24051 7080 24083
rect 7120 24051 7152 24083
rect 7192 24051 7224 24083
rect 7264 24051 7296 24083
rect 7336 24051 7368 24083
rect 7408 24051 7440 24083
rect 7480 24051 7512 24083
rect 7552 24051 7584 24083
rect 7624 24051 7656 24083
rect 7696 24051 7728 24083
rect 7768 24051 7800 24083
rect 7840 24051 7872 24083
rect 7912 24051 7944 24083
rect 7984 24051 8016 24083
rect 8056 24051 8088 24083
rect 8128 24051 8160 24083
rect 8200 24051 8232 24083
rect 8272 24051 8304 24083
rect 8344 24051 8376 24083
rect 8416 24051 8448 24083
rect 8488 24051 8520 24083
rect 8560 24051 8592 24083
rect 8632 24051 8664 24083
rect 8704 24051 8736 24083
rect 8776 24051 8808 24083
rect 8848 24051 8880 24083
rect 8920 24051 8952 24083
rect 8992 24051 9024 24083
rect 9064 24051 9096 24083
rect 9136 24051 9168 24083
rect 9208 24051 9240 24083
rect 9280 24051 9312 24083
rect 9352 24051 9384 24083
rect 9424 24051 9456 24083
rect 9496 24051 9528 24083
rect 9568 24051 9600 24083
rect 9640 24051 9672 24083
rect 9712 24051 9744 24083
rect 9784 24051 9816 24083
rect 9856 24051 9888 24083
rect 9928 24051 9960 24083
rect 10000 24051 10032 24083
rect 10072 24051 10104 24083
rect 10144 24051 10176 24083
rect 10216 24051 10248 24083
rect 10288 24051 10320 24083
rect 10360 24051 10392 24083
rect 10432 24051 10464 24083
rect 10504 24051 10536 24083
rect 10576 24051 10608 24083
rect 10648 24051 10680 24083
rect 10720 24051 10752 24083
rect 10792 24051 10824 24083
rect 10864 24051 10896 24083
rect 10936 24051 10968 24083
rect 11008 24051 11040 24083
rect 11080 24051 11112 24083
rect 11152 24051 11184 24083
rect 11224 24051 11256 24083
rect 11296 24051 11328 24083
rect 11368 24051 11400 24083
rect 11440 24051 11472 24083
rect 11512 24051 11544 24083
rect 11584 24051 11616 24083
rect 11656 24051 11688 24083
rect 11728 24051 11760 24083
rect 11800 24051 11832 24083
rect 11872 24051 11904 24083
rect 11944 24051 11976 24083
rect 12016 24051 12048 24083
rect 12088 24051 12120 24083
rect 12160 24051 12192 24083
rect 12232 24051 12264 24083
rect 12304 24051 12336 24083
rect 12376 24051 12408 24083
rect 12448 24051 12480 24083
rect 12520 24051 12552 24083
rect 12592 24051 12624 24083
rect 12664 24051 12696 24083
rect 12736 24051 12768 24083
rect 12808 24051 12840 24083
rect 12880 24051 12912 24083
rect 12952 24051 12984 24083
rect 13024 24051 13056 24083
rect 13096 24051 13128 24083
rect 13168 24051 13200 24083
rect 13240 24051 13272 24083
rect 13312 24051 13344 24083
rect 13384 24051 13416 24083
rect 13456 24051 13488 24083
rect 13528 24051 13560 24083
rect 13600 24051 13632 24083
rect 13672 24051 13704 24083
rect 13744 24051 13776 24083
rect 13816 24051 13848 24083
rect 13888 24051 13920 24083
rect 13960 24051 13992 24083
rect 14032 24051 14064 24083
rect 14104 24051 14136 24083
rect 14176 24051 14208 24083
rect 14248 24051 14280 24083
rect 14320 24051 14352 24083
rect 14392 24051 14424 24083
rect 14464 24051 14496 24083
rect 14536 24051 14568 24083
rect 14608 24051 14640 24083
rect 14680 24051 14712 24083
rect 14752 24051 14784 24083
rect 14824 24051 14856 24083
rect 14896 24051 14928 24083
rect 14968 24051 15000 24083
rect 15040 24051 15072 24083
rect 15112 24051 15144 24083
rect 15184 24051 15216 24083
rect 15256 24051 15288 24083
rect 15328 24051 15360 24083
rect 15400 24051 15432 24083
rect 15472 24051 15504 24083
rect 15544 24051 15576 24083
rect 15616 24051 15648 24083
rect 15688 24051 15720 24083
rect 15760 24051 15792 24083
rect 15832 24051 15864 24083
rect 15904 24051 15936 24083
rect 64 23979 96 24011
rect 136 23979 168 24011
rect 208 23979 240 24011
rect 280 23979 312 24011
rect 352 23979 384 24011
rect 424 23979 456 24011
rect 496 23979 528 24011
rect 568 23979 600 24011
rect 640 23979 672 24011
rect 712 23979 744 24011
rect 784 23979 816 24011
rect 856 23979 888 24011
rect 928 23979 960 24011
rect 1000 23979 1032 24011
rect 1072 23979 1104 24011
rect 1144 23979 1176 24011
rect 1216 23979 1248 24011
rect 1288 23979 1320 24011
rect 1360 23979 1392 24011
rect 1432 23979 1464 24011
rect 1504 23979 1536 24011
rect 1576 23979 1608 24011
rect 1648 23979 1680 24011
rect 1720 23979 1752 24011
rect 1792 23979 1824 24011
rect 1864 23979 1896 24011
rect 1936 23979 1968 24011
rect 2008 23979 2040 24011
rect 2080 23979 2112 24011
rect 2152 23979 2184 24011
rect 2224 23979 2256 24011
rect 2296 23979 2328 24011
rect 2368 23979 2400 24011
rect 2440 23979 2472 24011
rect 2512 23979 2544 24011
rect 2584 23979 2616 24011
rect 2656 23979 2688 24011
rect 2728 23979 2760 24011
rect 2800 23979 2832 24011
rect 2872 23979 2904 24011
rect 2944 23979 2976 24011
rect 3016 23979 3048 24011
rect 3088 23979 3120 24011
rect 3160 23979 3192 24011
rect 3232 23979 3264 24011
rect 3304 23979 3336 24011
rect 3376 23979 3408 24011
rect 3448 23979 3480 24011
rect 3520 23979 3552 24011
rect 3592 23979 3624 24011
rect 3664 23979 3696 24011
rect 3736 23979 3768 24011
rect 3808 23979 3840 24011
rect 3880 23979 3912 24011
rect 3952 23979 3984 24011
rect 4024 23979 4056 24011
rect 4096 23979 4128 24011
rect 4168 23979 4200 24011
rect 4240 23979 4272 24011
rect 4312 23979 4344 24011
rect 4384 23979 4416 24011
rect 4456 23979 4488 24011
rect 4528 23979 4560 24011
rect 4600 23979 4632 24011
rect 4672 23979 4704 24011
rect 4744 23979 4776 24011
rect 4816 23979 4848 24011
rect 4888 23979 4920 24011
rect 4960 23979 4992 24011
rect 5032 23979 5064 24011
rect 5104 23979 5136 24011
rect 5176 23979 5208 24011
rect 5248 23979 5280 24011
rect 5320 23979 5352 24011
rect 5392 23979 5424 24011
rect 5464 23979 5496 24011
rect 5536 23979 5568 24011
rect 5608 23979 5640 24011
rect 5680 23979 5712 24011
rect 5752 23979 5784 24011
rect 5824 23979 5856 24011
rect 5896 23979 5928 24011
rect 5968 23979 6000 24011
rect 6040 23979 6072 24011
rect 6112 23979 6144 24011
rect 6184 23979 6216 24011
rect 6256 23979 6288 24011
rect 6328 23979 6360 24011
rect 6400 23979 6432 24011
rect 6472 23979 6504 24011
rect 6544 23979 6576 24011
rect 6616 23979 6648 24011
rect 6688 23979 6720 24011
rect 6760 23979 6792 24011
rect 6832 23979 6864 24011
rect 6904 23979 6936 24011
rect 6976 23979 7008 24011
rect 7048 23979 7080 24011
rect 7120 23979 7152 24011
rect 7192 23979 7224 24011
rect 7264 23979 7296 24011
rect 7336 23979 7368 24011
rect 7408 23979 7440 24011
rect 7480 23979 7512 24011
rect 7552 23979 7584 24011
rect 7624 23979 7656 24011
rect 7696 23979 7728 24011
rect 7768 23979 7800 24011
rect 7840 23979 7872 24011
rect 7912 23979 7944 24011
rect 7984 23979 8016 24011
rect 8056 23979 8088 24011
rect 8128 23979 8160 24011
rect 8200 23979 8232 24011
rect 8272 23979 8304 24011
rect 8344 23979 8376 24011
rect 8416 23979 8448 24011
rect 8488 23979 8520 24011
rect 8560 23979 8592 24011
rect 8632 23979 8664 24011
rect 8704 23979 8736 24011
rect 8776 23979 8808 24011
rect 8848 23979 8880 24011
rect 8920 23979 8952 24011
rect 8992 23979 9024 24011
rect 9064 23979 9096 24011
rect 9136 23979 9168 24011
rect 9208 23979 9240 24011
rect 9280 23979 9312 24011
rect 9352 23979 9384 24011
rect 9424 23979 9456 24011
rect 9496 23979 9528 24011
rect 9568 23979 9600 24011
rect 9640 23979 9672 24011
rect 9712 23979 9744 24011
rect 9784 23979 9816 24011
rect 9856 23979 9888 24011
rect 9928 23979 9960 24011
rect 10000 23979 10032 24011
rect 10072 23979 10104 24011
rect 10144 23979 10176 24011
rect 10216 23979 10248 24011
rect 10288 23979 10320 24011
rect 10360 23979 10392 24011
rect 10432 23979 10464 24011
rect 10504 23979 10536 24011
rect 10576 23979 10608 24011
rect 10648 23979 10680 24011
rect 10720 23979 10752 24011
rect 10792 23979 10824 24011
rect 10864 23979 10896 24011
rect 10936 23979 10968 24011
rect 11008 23979 11040 24011
rect 11080 23979 11112 24011
rect 11152 23979 11184 24011
rect 11224 23979 11256 24011
rect 11296 23979 11328 24011
rect 11368 23979 11400 24011
rect 11440 23979 11472 24011
rect 11512 23979 11544 24011
rect 11584 23979 11616 24011
rect 11656 23979 11688 24011
rect 11728 23979 11760 24011
rect 11800 23979 11832 24011
rect 11872 23979 11904 24011
rect 11944 23979 11976 24011
rect 12016 23979 12048 24011
rect 12088 23979 12120 24011
rect 12160 23979 12192 24011
rect 12232 23979 12264 24011
rect 12304 23979 12336 24011
rect 12376 23979 12408 24011
rect 12448 23979 12480 24011
rect 12520 23979 12552 24011
rect 12592 23979 12624 24011
rect 12664 23979 12696 24011
rect 12736 23979 12768 24011
rect 12808 23979 12840 24011
rect 12880 23979 12912 24011
rect 12952 23979 12984 24011
rect 13024 23979 13056 24011
rect 13096 23979 13128 24011
rect 13168 23979 13200 24011
rect 13240 23979 13272 24011
rect 13312 23979 13344 24011
rect 13384 23979 13416 24011
rect 13456 23979 13488 24011
rect 13528 23979 13560 24011
rect 13600 23979 13632 24011
rect 13672 23979 13704 24011
rect 13744 23979 13776 24011
rect 13816 23979 13848 24011
rect 13888 23979 13920 24011
rect 13960 23979 13992 24011
rect 14032 23979 14064 24011
rect 14104 23979 14136 24011
rect 14176 23979 14208 24011
rect 14248 23979 14280 24011
rect 14320 23979 14352 24011
rect 14392 23979 14424 24011
rect 14464 23979 14496 24011
rect 14536 23979 14568 24011
rect 14608 23979 14640 24011
rect 14680 23979 14712 24011
rect 14752 23979 14784 24011
rect 14824 23979 14856 24011
rect 14896 23979 14928 24011
rect 14968 23979 15000 24011
rect 15040 23979 15072 24011
rect 15112 23979 15144 24011
rect 15184 23979 15216 24011
rect 15256 23979 15288 24011
rect 15328 23979 15360 24011
rect 15400 23979 15432 24011
rect 15472 23979 15504 24011
rect 15544 23979 15576 24011
rect 15616 23979 15648 24011
rect 15688 23979 15720 24011
rect 15760 23979 15792 24011
rect 15832 23979 15864 24011
rect 15904 23979 15936 24011
rect 64 23907 96 23939
rect 136 23907 168 23939
rect 208 23907 240 23939
rect 280 23907 312 23939
rect 352 23907 384 23939
rect 424 23907 456 23939
rect 496 23907 528 23939
rect 568 23907 600 23939
rect 640 23907 672 23939
rect 712 23907 744 23939
rect 784 23907 816 23939
rect 856 23907 888 23939
rect 928 23907 960 23939
rect 1000 23907 1032 23939
rect 1072 23907 1104 23939
rect 1144 23907 1176 23939
rect 1216 23907 1248 23939
rect 1288 23907 1320 23939
rect 1360 23907 1392 23939
rect 1432 23907 1464 23939
rect 1504 23907 1536 23939
rect 1576 23907 1608 23939
rect 1648 23907 1680 23939
rect 1720 23907 1752 23939
rect 1792 23907 1824 23939
rect 1864 23907 1896 23939
rect 1936 23907 1968 23939
rect 2008 23907 2040 23939
rect 2080 23907 2112 23939
rect 2152 23907 2184 23939
rect 2224 23907 2256 23939
rect 2296 23907 2328 23939
rect 2368 23907 2400 23939
rect 2440 23907 2472 23939
rect 2512 23907 2544 23939
rect 2584 23907 2616 23939
rect 2656 23907 2688 23939
rect 2728 23907 2760 23939
rect 2800 23907 2832 23939
rect 2872 23907 2904 23939
rect 2944 23907 2976 23939
rect 3016 23907 3048 23939
rect 3088 23907 3120 23939
rect 3160 23907 3192 23939
rect 3232 23907 3264 23939
rect 3304 23907 3336 23939
rect 3376 23907 3408 23939
rect 3448 23907 3480 23939
rect 3520 23907 3552 23939
rect 3592 23907 3624 23939
rect 3664 23907 3696 23939
rect 3736 23907 3768 23939
rect 3808 23907 3840 23939
rect 3880 23907 3912 23939
rect 3952 23907 3984 23939
rect 4024 23907 4056 23939
rect 4096 23907 4128 23939
rect 4168 23907 4200 23939
rect 4240 23907 4272 23939
rect 4312 23907 4344 23939
rect 4384 23907 4416 23939
rect 4456 23907 4488 23939
rect 4528 23907 4560 23939
rect 4600 23907 4632 23939
rect 4672 23907 4704 23939
rect 4744 23907 4776 23939
rect 4816 23907 4848 23939
rect 4888 23907 4920 23939
rect 4960 23907 4992 23939
rect 5032 23907 5064 23939
rect 5104 23907 5136 23939
rect 5176 23907 5208 23939
rect 5248 23907 5280 23939
rect 5320 23907 5352 23939
rect 5392 23907 5424 23939
rect 5464 23907 5496 23939
rect 5536 23907 5568 23939
rect 5608 23907 5640 23939
rect 5680 23907 5712 23939
rect 5752 23907 5784 23939
rect 5824 23907 5856 23939
rect 5896 23907 5928 23939
rect 5968 23907 6000 23939
rect 6040 23907 6072 23939
rect 6112 23907 6144 23939
rect 6184 23907 6216 23939
rect 6256 23907 6288 23939
rect 6328 23907 6360 23939
rect 6400 23907 6432 23939
rect 6472 23907 6504 23939
rect 6544 23907 6576 23939
rect 6616 23907 6648 23939
rect 6688 23907 6720 23939
rect 6760 23907 6792 23939
rect 6832 23907 6864 23939
rect 6904 23907 6936 23939
rect 6976 23907 7008 23939
rect 7048 23907 7080 23939
rect 7120 23907 7152 23939
rect 7192 23907 7224 23939
rect 7264 23907 7296 23939
rect 7336 23907 7368 23939
rect 7408 23907 7440 23939
rect 7480 23907 7512 23939
rect 7552 23907 7584 23939
rect 7624 23907 7656 23939
rect 7696 23907 7728 23939
rect 7768 23907 7800 23939
rect 7840 23907 7872 23939
rect 7912 23907 7944 23939
rect 7984 23907 8016 23939
rect 8056 23907 8088 23939
rect 8128 23907 8160 23939
rect 8200 23907 8232 23939
rect 8272 23907 8304 23939
rect 8344 23907 8376 23939
rect 8416 23907 8448 23939
rect 8488 23907 8520 23939
rect 8560 23907 8592 23939
rect 8632 23907 8664 23939
rect 8704 23907 8736 23939
rect 8776 23907 8808 23939
rect 8848 23907 8880 23939
rect 8920 23907 8952 23939
rect 8992 23907 9024 23939
rect 9064 23907 9096 23939
rect 9136 23907 9168 23939
rect 9208 23907 9240 23939
rect 9280 23907 9312 23939
rect 9352 23907 9384 23939
rect 9424 23907 9456 23939
rect 9496 23907 9528 23939
rect 9568 23907 9600 23939
rect 9640 23907 9672 23939
rect 9712 23907 9744 23939
rect 9784 23907 9816 23939
rect 9856 23907 9888 23939
rect 9928 23907 9960 23939
rect 10000 23907 10032 23939
rect 10072 23907 10104 23939
rect 10144 23907 10176 23939
rect 10216 23907 10248 23939
rect 10288 23907 10320 23939
rect 10360 23907 10392 23939
rect 10432 23907 10464 23939
rect 10504 23907 10536 23939
rect 10576 23907 10608 23939
rect 10648 23907 10680 23939
rect 10720 23907 10752 23939
rect 10792 23907 10824 23939
rect 10864 23907 10896 23939
rect 10936 23907 10968 23939
rect 11008 23907 11040 23939
rect 11080 23907 11112 23939
rect 11152 23907 11184 23939
rect 11224 23907 11256 23939
rect 11296 23907 11328 23939
rect 11368 23907 11400 23939
rect 11440 23907 11472 23939
rect 11512 23907 11544 23939
rect 11584 23907 11616 23939
rect 11656 23907 11688 23939
rect 11728 23907 11760 23939
rect 11800 23907 11832 23939
rect 11872 23907 11904 23939
rect 11944 23907 11976 23939
rect 12016 23907 12048 23939
rect 12088 23907 12120 23939
rect 12160 23907 12192 23939
rect 12232 23907 12264 23939
rect 12304 23907 12336 23939
rect 12376 23907 12408 23939
rect 12448 23907 12480 23939
rect 12520 23907 12552 23939
rect 12592 23907 12624 23939
rect 12664 23907 12696 23939
rect 12736 23907 12768 23939
rect 12808 23907 12840 23939
rect 12880 23907 12912 23939
rect 12952 23907 12984 23939
rect 13024 23907 13056 23939
rect 13096 23907 13128 23939
rect 13168 23907 13200 23939
rect 13240 23907 13272 23939
rect 13312 23907 13344 23939
rect 13384 23907 13416 23939
rect 13456 23907 13488 23939
rect 13528 23907 13560 23939
rect 13600 23907 13632 23939
rect 13672 23907 13704 23939
rect 13744 23907 13776 23939
rect 13816 23907 13848 23939
rect 13888 23907 13920 23939
rect 13960 23907 13992 23939
rect 14032 23907 14064 23939
rect 14104 23907 14136 23939
rect 14176 23907 14208 23939
rect 14248 23907 14280 23939
rect 14320 23907 14352 23939
rect 14392 23907 14424 23939
rect 14464 23907 14496 23939
rect 14536 23907 14568 23939
rect 14608 23907 14640 23939
rect 14680 23907 14712 23939
rect 14752 23907 14784 23939
rect 14824 23907 14856 23939
rect 14896 23907 14928 23939
rect 14968 23907 15000 23939
rect 15040 23907 15072 23939
rect 15112 23907 15144 23939
rect 15184 23907 15216 23939
rect 15256 23907 15288 23939
rect 15328 23907 15360 23939
rect 15400 23907 15432 23939
rect 15472 23907 15504 23939
rect 15544 23907 15576 23939
rect 15616 23907 15648 23939
rect 15688 23907 15720 23939
rect 15760 23907 15792 23939
rect 15832 23907 15864 23939
rect 15904 23907 15936 23939
rect 64 23835 96 23867
rect 136 23835 168 23867
rect 208 23835 240 23867
rect 280 23835 312 23867
rect 352 23835 384 23867
rect 424 23835 456 23867
rect 496 23835 528 23867
rect 568 23835 600 23867
rect 640 23835 672 23867
rect 712 23835 744 23867
rect 784 23835 816 23867
rect 856 23835 888 23867
rect 928 23835 960 23867
rect 1000 23835 1032 23867
rect 1072 23835 1104 23867
rect 1144 23835 1176 23867
rect 1216 23835 1248 23867
rect 1288 23835 1320 23867
rect 1360 23835 1392 23867
rect 1432 23835 1464 23867
rect 1504 23835 1536 23867
rect 1576 23835 1608 23867
rect 1648 23835 1680 23867
rect 1720 23835 1752 23867
rect 1792 23835 1824 23867
rect 1864 23835 1896 23867
rect 1936 23835 1968 23867
rect 2008 23835 2040 23867
rect 2080 23835 2112 23867
rect 2152 23835 2184 23867
rect 2224 23835 2256 23867
rect 2296 23835 2328 23867
rect 2368 23835 2400 23867
rect 2440 23835 2472 23867
rect 2512 23835 2544 23867
rect 2584 23835 2616 23867
rect 2656 23835 2688 23867
rect 2728 23835 2760 23867
rect 2800 23835 2832 23867
rect 2872 23835 2904 23867
rect 2944 23835 2976 23867
rect 3016 23835 3048 23867
rect 3088 23835 3120 23867
rect 3160 23835 3192 23867
rect 3232 23835 3264 23867
rect 3304 23835 3336 23867
rect 3376 23835 3408 23867
rect 3448 23835 3480 23867
rect 3520 23835 3552 23867
rect 3592 23835 3624 23867
rect 3664 23835 3696 23867
rect 3736 23835 3768 23867
rect 3808 23835 3840 23867
rect 3880 23835 3912 23867
rect 3952 23835 3984 23867
rect 4024 23835 4056 23867
rect 4096 23835 4128 23867
rect 4168 23835 4200 23867
rect 4240 23835 4272 23867
rect 4312 23835 4344 23867
rect 4384 23835 4416 23867
rect 4456 23835 4488 23867
rect 4528 23835 4560 23867
rect 4600 23835 4632 23867
rect 4672 23835 4704 23867
rect 4744 23835 4776 23867
rect 4816 23835 4848 23867
rect 4888 23835 4920 23867
rect 4960 23835 4992 23867
rect 5032 23835 5064 23867
rect 5104 23835 5136 23867
rect 5176 23835 5208 23867
rect 5248 23835 5280 23867
rect 5320 23835 5352 23867
rect 5392 23835 5424 23867
rect 5464 23835 5496 23867
rect 5536 23835 5568 23867
rect 5608 23835 5640 23867
rect 5680 23835 5712 23867
rect 5752 23835 5784 23867
rect 5824 23835 5856 23867
rect 5896 23835 5928 23867
rect 5968 23835 6000 23867
rect 6040 23835 6072 23867
rect 6112 23835 6144 23867
rect 6184 23835 6216 23867
rect 6256 23835 6288 23867
rect 6328 23835 6360 23867
rect 6400 23835 6432 23867
rect 6472 23835 6504 23867
rect 6544 23835 6576 23867
rect 6616 23835 6648 23867
rect 6688 23835 6720 23867
rect 6760 23835 6792 23867
rect 6832 23835 6864 23867
rect 6904 23835 6936 23867
rect 6976 23835 7008 23867
rect 7048 23835 7080 23867
rect 7120 23835 7152 23867
rect 7192 23835 7224 23867
rect 7264 23835 7296 23867
rect 7336 23835 7368 23867
rect 7408 23835 7440 23867
rect 7480 23835 7512 23867
rect 7552 23835 7584 23867
rect 7624 23835 7656 23867
rect 7696 23835 7728 23867
rect 7768 23835 7800 23867
rect 7840 23835 7872 23867
rect 7912 23835 7944 23867
rect 7984 23835 8016 23867
rect 8056 23835 8088 23867
rect 8128 23835 8160 23867
rect 8200 23835 8232 23867
rect 8272 23835 8304 23867
rect 8344 23835 8376 23867
rect 8416 23835 8448 23867
rect 8488 23835 8520 23867
rect 8560 23835 8592 23867
rect 8632 23835 8664 23867
rect 8704 23835 8736 23867
rect 8776 23835 8808 23867
rect 8848 23835 8880 23867
rect 8920 23835 8952 23867
rect 8992 23835 9024 23867
rect 9064 23835 9096 23867
rect 9136 23835 9168 23867
rect 9208 23835 9240 23867
rect 9280 23835 9312 23867
rect 9352 23835 9384 23867
rect 9424 23835 9456 23867
rect 9496 23835 9528 23867
rect 9568 23835 9600 23867
rect 9640 23835 9672 23867
rect 9712 23835 9744 23867
rect 9784 23835 9816 23867
rect 9856 23835 9888 23867
rect 9928 23835 9960 23867
rect 10000 23835 10032 23867
rect 10072 23835 10104 23867
rect 10144 23835 10176 23867
rect 10216 23835 10248 23867
rect 10288 23835 10320 23867
rect 10360 23835 10392 23867
rect 10432 23835 10464 23867
rect 10504 23835 10536 23867
rect 10576 23835 10608 23867
rect 10648 23835 10680 23867
rect 10720 23835 10752 23867
rect 10792 23835 10824 23867
rect 10864 23835 10896 23867
rect 10936 23835 10968 23867
rect 11008 23835 11040 23867
rect 11080 23835 11112 23867
rect 11152 23835 11184 23867
rect 11224 23835 11256 23867
rect 11296 23835 11328 23867
rect 11368 23835 11400 23867
rect 11440 23835 11472 23867
rect 11512 23835 11544 23867
rect 11584 23835 11616 23867
rect 11656 23835 11688 23867
rect 11728 23835 11760 23867
rect 11800 23835 11832 23867
rect 11872 23835 11904 23867
rect 11944 23835 11976 23867
rect 12016 23835 12048 23867
rect 12088 23835 12120 23867
rect 12160 23835 12192 23867
rect 12232 23835 12264 23867
rect 12304 23835 12336 23867
rect 12376 23835 12408 23867
rect 12448 23835 12480 23867
rect 12520 23835 12552 23867
rect 12592 23835 12624 23867
rect 12664 23835 12696 23867
rect 12736 23835 12768 23867
rect 12808 23835 12840 23867
rect 12880 23835 12912 23867
rect 12952 23835 12984 23867
rect 13024 23835 13056 23867
rect 13096 23835 13128 23867
rect 13168 23835 13200 23867
rect 13240 23835 13272 23867
rect 13312 23835 13344 23867
rect 13384 23835 13416 23867
rect 13456 23835 13488 23867
rect 13528 23835 13560 23867
rect 13600 23835 13632 23867
rect 13672 23835 13704 23867
rect 13744 23835 13776 23867
rect 13816 23835 13848 23867
rect 13888 23835 13920 23867
rect 13960 23835 13992 23867
rect 14032 23835 14064 23867
rect 14104 23835 14136 23867
rect 14176 23835 14208 23867
rect 14248 23835 14280 23867
rect 14320 23835 14352 23867
rect 14392 23835 14424 23867
rect 14464 23835 14496 23867
rect 14536 23835 14568 23867
rect 14608 23835 14640 23867
rect 14680 23835 14712 23867
rect 14752 23835 14784 23867
rect 14824 23835 14856 23867
rect 14896 23835 14928 23867
rect 14968 23835 15000 23867
rect 15040 23835 15072 23867
rect 15112 23835 15144 23867
rect 15184 23835 15216 23867
rect 15256 23835 15288 23867
rect 15328 23835 15360 23867
rect 15400 23835 15432 23867
rect 15472 23835 15504 23867
rect 15544 23835 15576 23867
rect 15616 23835 15648 23867
rect 15688 23835 15720 23867
rect 15760 23835 15792 23867
rect 15832 23835 15864 23867
rect 15904 23835 15936 23867
rect 64 23763 96 23795
rect 136 23763 168 23795
rect 208 23763 240 23795
rect 280 23763 312 23795
rect 352 23763 384 23795
rect 424 23763 456 23795
rect 496 23763 528 23795
rect 568 23763 600 23795
rect 640 23763 672 23795
rect 712 23763 744 23795
rect 784 23763 816 23795
rect 856 23763 888 23795
rect 928 23763 960 23795
rect 1000 23763 1032 23795
rect 1072 23763 1104 23795
rect 1144 23763 1176 23795
rect 1216 23763 1248 23795
rect 1288 23763 1320 23795
rect 1360 23763 1392 23795
rect 1432 23763 1464 23795
rect 1504 23763 1536 23795
rect 1576 23763 1608 23795
rect 1648 23763 1680 23795
rect 1720 23763 1752 23795
rect 1792 23763 1824 23795
rect 1864 23763 1896 23795
rect 1936 23763 1968 23795
rect 2008 23763 2040 23795
rect 2080 23763 2112 23795
rect 2152 23763 2184 23795
rect 2224 23763 2256 23795
rect 2296 23763 2328 23795
rect 2368 23763 2400 23795
rect 2440 23763 2472 23795
rect 2512 23763 2544 23795
rect 2584 23763 2616 23795
rect 2656 23763 2688 23795
rect 2728 23763 2760 23795
rect 2800 23763 2832 23795
rect 2872 23763 2904 23795
rect 2944 23763 2976 23795
rect 3016 23763 3048 23795
rect 3088 23763 3120 23795
rect 3160 23763 3192 23795
rect 3232 23763 3264 23795
rect 3304 23763 3336 23795
rect 3376 23763 3408 23795
rect 3448 23763 3480 23795
rect 3520 23763 3552 23795
rect 3592 23763 3624 23795
rect 3664 23763 3696 23795
rect 3736 23763 3768 23795
rect 3808 23763 3840 23795
rect 3880 23763 3912 23795
rect 3952 23763 3984 23795
rect 4024 23763 4056 23795
rect 4096 23763 4128 23795
rect 4168 23763 4200 23795
rect 4240 23763 4272 23795
rect 4312 23763 4344 23795
rect 4384 23763 4416 23795
rect 4456 23763 4488 23795
rect 4528 23763 4560 23795
rect 4600 23763 4632 23795
rect 4672 23763 4704 23795
rect 4744 23763 4776 23795
rect 4816 23763 4848 23795
rect 4888 23763 4920 23795
rect 4960 23763 4992 23795
rect 5032 23763 5064 23795
rect 5104 23763 5136 23795
rect 5176 23763 5208 23795
rect 5248 23763 5280 23795
rect 5320 23763 5352 23795
rect 5392 23763 5424 23795
rect 5464 23763 5496 23795
rect 5536 23763 5568 23795
rect 5608 23763 5640 23795
rect 5680 23763 5712 23795
rect 5752 23763 5784 23795
rect 5824 23763 5856 23795
rect 5896 23763 5928 23795
rect 5968 23763 6000 23795
rect 6040 23763 6072 23795
rect 6112 23763 6144 23795
rect 6184 23763 6216 23795
rect 6256 23763 6288 23795
rect 6328 23763 6360 23795
rect 6400 23763 6432 23795
rect 6472 23763 6504 23795
rect 6544 23763 6576 23795
rect 6616 23763 6648 23795
rect 6688 23763 6720 23795
rect 6760 23763 6792 23795
rect 6832 23763 6864 23795
rect 6904 23763 6936 23795
rect 6976 23763 7008 23795
rect 7048 23763 7080 23795
rect 7120 23763 7152 23795
rect 7192 23763 7224 23795
rect 7264 23763 7296 23795
rect 7336 23763 7368 23795
rect 7408 23763 7440 23795
rect 7480 23763 7512 23795
rect 7552 23763 7584 23795
rect 7624 23763 7656 23795
rect 7696 23763 7728 23795
rect 7768 23763 7800 23795
rect 7840 23763 7872 23795
rect 7912 23763 7944 23795
rect 7984 23763 8016 23795
rect 8056 23763 8088 23795
rect 8128 23763 8160 23795
rect 8200 23763 8232 23795
rect 8272 23763 8304 23795
rect 8344 23763 8376 23795
rect 8416 23763 8448 23795
rect 8488 23763 8520 23795
rect 8560 23763 8592 23795
rect 8632 23763 8664 23795
rect 8704 23763 8736 23795
rect 8776 23763 8808 23795
rect 8848 23763 8880 23795
rect 8920 23763 8952 23795
rect 8992 23763 9024 23795
rect 9064 23763 9096 23795
rect 9136 23763 9168 23795
rect 9208 23763 9240 23795
rect 9280 23763 9312 23795
rect 9352 23763 9384 23795
rect 9424 23763 9456 23795
rect 9496 23763 9528 23795
rect 9568 23763 9600 23795
rect 9640 23763 9672 23795
rect 9712 23763 9744 23795
rect 9784 23763 9816 23795
rect 9856 23763 9888 23795
rect 9928 23763 9960 23795
rect 10000 23763 10032 23795
rect 10072 23763 10104 23795
rect 10144 23763 10176 23795
rect 10216 23763 10248 23795
rect 10288 23763 10320 23795
rect 10360 23763 10392 23795
rect 10432 23763 10464 23795
rect 10504 23763 10536 23795
rect 10576 23763 10608 23795
rect 10648 23763 10680 23795
rect 10720 23763 10752 23795
rect 10792 23763 10824 23795
rect 10864 23763 10896 23795
rect 10936 23763 10968 23795
rect 11008 23763 11040 23795
rect 11080 23763 11112 23795
rect 11152 23763 11184 23795
rect 11224 23763 11256 23795
rect 11296 23763 11328 23795
rect 11368 23763 11400 23795
rect 11440 23763 11472 23795
rect 11512 23763 11544 23795
rect 11584 23763 11616 23795
rect 11656 23763 11688 23795
rect 11728 23763 11760 23795
rect 11800 23763 11832 23795
rect 11872 23763 11904 23795
rect 11944 23763 11976 23795
rect 12016 23763 12048 23795
rect 12088 23763 12120 23795
rect 12160 23763 12192 23795
rect 12232 23763 12264 23795
rect 12304 23763 12336 23795
rect 12376 23763 12408 23795
rect 12448 23763 12480 23795
rect 12520 23763 12552 23795
rect 12592 23763 12624 23795
rect 12664 23763 12696 23795
rect 12736 23763 12768 23795
rect 12808 23763 12840 23795
rect 12880 23763 12912 23795
rect 12952 23763 12984 23795
rect 13024 23763 13056 23795
rect 13096 23763 13128 23795
rect 13168 23763 13200 23795
rect 13240 23763 13272 23795
rect 13312 23763 13344 23795
rect 13384 23763 13416 23795
rect 13456 23763 13488 23795
rect 13528 23763 13560 23795
rect 13600 23763 13632 23795
rect 13672 23763 13704 23795
rect 13744 23763 13776 23795
rect 13816 23763 13848 23795
rect 13888 23763 13920 23795
rect 13960 23763 13992 23795
rect 14032 23763 14064 23795
rect 14104 23763 14136 23795
rect 14176 23763 14208 23795
rect 14248 23763 14280 23795
rect 14320 23763 14352 23795
rect 14392 23763 14424 23795
rect 14464 23763 14496 23795
rect 14536 23763 14568 23795
rect 14608 23763 14640 23795
rect 14680 23763 14712 23795
rect 14752 23763 14784 23795
rect 14824 23763 14856 23795
rect 14896 23763 14928 23795
rect 14968 23763 15000 23795
rect 15040 23763 15072 23795
rect 15112 23763 15144 23795
rect 15184 23763 15216 23795
rect 15256 23763 15288 23795
rect 15328 23763 15360 23795
rect 15400 23763 15432 23795
rect 15472 23763 15504 23795
rect 15544 23763 15576 23795
rect 15616 23763 15648 23795
rect 15688 23763 15720 23795
rect 15760 23763 15792 23795
rect 15832 23763 15864 23795
rect 15904 23763 15936 23795
rect 64 23691 96 23723
rect 136 23691 168 23723
rect 208 23691 240 23723
rect 280 23691 312 23723
rect 352 23691 384 23723
rect 424 23691 456 23723
rect 496 23691 528 23723
rect 568 23691 600 23723
rect 640 23691 672 23723
rect 712 23691 744 23723
rect 784 23691 816 23723
rect 856 23691 888 23723
rect 928 23691 960 23723
rect 1000 23691 1032 23723
rect 1072 23691 1104 23723
rect 1144 23691 1176 23723
rect 1216 23691 1248 23723
rect 1288 23691 1320 23723
rect 1360 23691 1392 23723
rect 1432 23691 1464 23723
rect 1504 23691 1536 23723
rect 1576 23691 1608 23723
rect 1648 23691 1680 23723
rect 1720 23691 1752 23723
rect 1792 23691 1824 23723
rect 1864 23691 1896 23723
rect 1936 23691 1968 23723
rect 2008 23691 2040 23723
rect 2080 23691 2112 23723
rect 2152 23691 2184 23723
rect 2224 23691 2256 23723
rect 2296 23691 2328 23723
rect 2368 23691 2400 23723
rect 2440 23691 2472 23723
rect 2512 23691 2544 23723
rect 2584 23691 2616 23723
rect 2656 23691 2688 23723
rect 2728 23691 2760 23723
rect 2800 23691 2832 23723
rect 2872 23691 2904 23723
rect 2944 23691 2976 23723
rect 3016 23691 3048 23723
rect 3088 23691 3120 23723
rect 3160 23691 3192 23723
rect 3232 23691 3264 23723
rect 3304 23691 3336 23723
rect 3376 23691 3408 23723
rect 3448 23691 3480 23723
rect 3520 23691 3552 23723
rect 3592 23691 3624 23723
rect 3664 23691 3696 23723
rect 3736 23691 3768 23723
rect 3808 23691 3840 23723
rect 3880 23691 3912 23723
rect 3952 23691 3984 23723
rect 4024 23691 4056 23723
rect 4096 23691 4128 23723
rect 4168 23691 4200 23723
rect 4240 23691 4272 23723
rect 4312 23691 4344 23723
rect 4384 23691 4416 23723
rect 4456 23691 4488 23723
rect 4528 23691 4560 23723
rect 4600 23691 4632 23723
rect 4672 23691 4704 23723
rect 4744 23691 4776 23723
rect 4816 23691 4848 23723
rect 4888 23691 4920 23723
rect 4960 23691 4992 23723
rect 5032 23691 5064 23723
rect 5104 23691 5136 23723
rect 5176 23691 5208 23723
rect 5248 23691 5280 23723
rect 5320 23691 5352 23723
rect 5392 23691 5424 23723
rect 5464 23691 5496 23723
rect 5536 23691 5568 23723
rect 5608 23691 5640 23723
rect 5680 23691 5712 23723
rect 5752 23691 5784 23723
rect 5824 23691 5856 23723
rect 5896 23691 5928 23723
rect 5968 23691 6000 23723
rect 6040 23691 6072 23723
rect 6112 23691 6144 23723
rect 6184 23691 6216 23723
rect 6256 23691 6288 23723
rect 6328 23691 6360 23723
rect 6400 23691 6432 23723
rect 6472 23691 6504 23723
rect 6544 23691 6576 23723
rect 6616 23691 6648 23723
rect 6688 23691 6720 23723
rect 6760 23691 6792 23723
rect 6832 23691 6864 23723
rect 6904 23691 6936 23723
rect 6976 23691 7008 23723
rect 7048 23691 7080 23723
rect 7120 23691 7152 23723
rect 7192 23691 7224 23723
rect 7264 23691 7296 23723
rect 7336 23691 7368 23723
rect 7408 23691 7440 23723
rect 7480 23691 7512 23723
rect 7552 23691 7584 23723
rect 7624 23691 7656 23723
rect 7696 23691 7728 23723
rect 7768 23691 7800 23723
rect 7840 23691 7872 23723
rect 7912 23691 7944 23723
rect 7984 23691 8016 23723
rect 8056 23691 8088 23723
rect 8128 23691 8160 23723
rect 8200 23691 8232 23723
rect 8272 23691 8304 23723
rect 8344 23691 8376 23723
rect 8416 23691 8448 23723
rect 8488 23691 8520 23723
rect 8560 23691 8592 23723
rect 8632 23691 8664 23723
rect 8704 23691 8736 23723
rect 8776 23691 8808 23723
rect 8848 23691 8880 23723
rect 8920 23691 8952 23723
rect 8992 23691 9024 23723
rect 9064 23691 9096 23723
rect 9136 23691 9168 23723
rect 9208 23691 9240 23723
rect 9280 23691 9312 23723
rect 9352 23691 9384 23723
rect 9424 23691 9456 23723
rect 9496 23691 9528 23723
rect 9568 23691 9600 23723
rect 9640 23691 9672 23723
rect 9712 23691 9744 23723
rect 9784 23691 9816 23723
rect 9856 23691 9888 23723
rect 9928 23691 9960 23723
rect 10000 23691 10032 23723
rect 10072 23691 10104 23723
rect 10144 23691 10176 23723
rect 10216 23691 10248 23723
rect 10288 23691 10320 23723
rect 10360 23691 10392 23723
rect 10432 23691 10464 23723
rect 10504 23691 10536 23723
rect 10576 23691 10608 23723
rect 10648 23691 10680 23723
rect 10720 23691 10752 23723
rect 10792 23691 10824 23723
rect 10864 23691 10896 23723
rect 10936 23691 10968 23723
rect 11008 23691 11040 23723
rect 11080 23691 11112 23723
rect 11152 23691 11184 23723
rect 11224 23691 11256 23723
rect 11296 23691 11328 23723
rect 11368 23691 11400 23723
rect 11440 23691 11472 23723
rect 11512 23691 11544 23723
rect 11584 23691 11616 23723
rect 11656 23691 11688 23723
rect 11728 23691 11760 23723
rect 11800 23691 11832 23723
rect 11872 23691 11904 23723
rect 11944 23691 11976 23723
rect 12016 23691 12048 23723
rect 12088 23691 12120 23723
rect 12160 23691 12192 23723
rect 12232 23691 12264 23723
rect 12304 23691 12336 23723
rect 12376 23691 12408 23723
rect 12448 23691 12480 23723
rect 12520 23691 12552 23723
rect 12592 23691 12624 23723
rect 12664 23691 12696 23723
rect 12736 23691 12768 23723
rect 12808 23691 12840 23723
rect 12880 23691 12912 23723
rect 12952 23691 12984 23723
rect 13024 23691 13056 23723
rect 13096 23691 13128 23723
rect 13168 23691 13200 23723
rect 13240 23691 13272 23723
rect 13312 23691 13344 23723
rect 13384 23691 13416 23723
rect 13456 23691 13488 23723
rect 13528 23691 13560 23723
rect 13600 23691 13632 23723
rect 13672 23691 13704 23723
rect 13744 23691 13776 23723
rect 13816 23691 13848 23723
rect 13888 23691 13920 23723
rect 13960 23691 13992 23723
rect 14032 23691 14064 23723
rect 14104 23691 14136 23723
rect 14176 23691 14208 23723
rect 14248 23691 14280 23723
rect 14320 23691 14352 23723
rect 14392 23691 14424 23723
rect 14464 23691 14496 23723
rect 14536 23691 14568 23723
rect 14608 23691 14640 23723
rect 14680 23691 14712 23723
rect 14752 23691 14784 23723
rect 14824 23691 14856 23723
rect 14896 23691 14928 23723
rect 14968 23691 15000 23723
rect 15040 23691 15072 23723
rect 15112 23691 15144 23723
rect 15184 23691 15216 23723
rect 15256 23691 15288 23723
rect 15328 23691 15360 23723
rect 15400 23691 15432 23723
rect 15472 23691 15504 23723
rect 15544 23691 15576 23723
rect 15616 23691 15648 23723
rect 15688 23691 15720 23723
rect 15760 23691 15792 23723
rect 15832 23691 15864 23723
rect 15904 23691 15936 23723
rect 64 23619 96 23651
rect 136 23619 168 23651
rect 208 23619 240 23651
rect 280 23619 312 23651
rect 352 23619 384 23651
rect 424 23619 456 23651
rect 496 23619 528 23651
rect 568 23619 600 23651
rect 640 23619 672 23651
rect 712 23619 744 23651
rect 784 23619 816 23651
rect 856 23619 888 23651
rect 928 23619 960 23651
rect 1000 23619 1032 23651
rect 1072 23619 1104 23651
rect 1144 23619 1176 23651
rect 1216 23619 1248 23651
rect 1288 23619 1320 23651
rect 1360 23619 1392 23651
rect 1432 23619 1464 23651
rect 1504 23619 1536 23651
rect 1576 23619 1608 23651
rect 1648 23619 1680 23651
rect 1720 23619 1752 23651
rect 1792 23619 1824 23651
rect 1864 23619 1896 23651
rect 1936 23619 1968 23651
rect 2008 23619 2040 23651
rect 2080 23619 2112 23651
rect 2152 23619 2184 23651
rect 2224 23619 2256 23651
rect 2296 23619 2328 23651
rect 2368 23619 2400 23651
rect 2440 23619 2472 23651
rect 2512 23619 2544 23651
rect 2584 23619 2616 23651
rect 2656 23619 2688 23651
rect 2728 23619 2760 23651
rect 2800 23619 2832 23651
rect 2872 23619 2904 23651
rect 2944 23619 2976 23651
rect 3016 23619 3048 23651
rect 3088 23619 3120 23651
rect 3160 23619 3192 23651
rect 3232 23619 3264 23651
rect 3304 23619 3336 23651
rect 3376 23619 3408 23651
rect 3448 23619 3480 23651
rect 3520 23619 3552 23651
rect 3592 23619 3624 23651
rect 3664 23619 3696 23651
rect 3736 23619 3768 23651
rect 3808 23619 3840 23651
rect 3880 23619 3912 23651
rect 3952 23619 3984 23651
rect 4024 23619 4056 23651
rect 4096 23619 4128 23651
rect 4168 23619 4200 23651
rect 4240 23619 4272 23651
rect 4312 23619 4344 23651
rect 4384 23619 4416 23651
rect 4456 23619 4488 23651
rect 4528 23619 4560 23651
rect 4600 23619 4632 23651
rect 4672 23619 4704 23651
rect 4744 23619 4776 23651
rect 4816 23619 4848 23651
rect 4888 23619 4920 23651
rect 4960 23619 4992 23651
rect 5032 23619 5064 23651
rect 5104 23619 5136 23651
rect 5176 23619 5208 23651
rect 5248 23619 5280 23651
rect 5320 23619 5352 23651
rect 5392 23619 5424 23651
rect 5464 23619 5496 23651
rect 5536 23619 5568 23651
rect 5608 23619 5640 23651
rect 5680 23619 5712 23651
rect 5752 23619 5784 23651
rect 5824 23619 5856 23651
rect 5896 23619 5928 23651
rect 5968 23619 6000 23651
rect 6040 23619 6072 23651
rect 6112 23619 6144 23651
rect 6184 23619 6216 23651
rect 6256 23619 6288 23651
rect 6328 23619 6360 23651
rect 6400 23619 6432 23651
rect 6472 23619 6504 23651
rect 6544 23619 6576 23651
rect 6616 23619 6648 23651
rect 6688 23619 6720 23651
rect 6760 23619 6792 23651
rect 6832 23619 6864 23651
rect 6904 23619 6936 23651
rect 6976 23619 7008 23651
rect 7048 23619 7080 23651
rect 7120 23619 7152 23651
rect 7192 23619 7224 23651
rect 7264 23619 7296 23651
rect 7336 23619 7368 23651
rect 7408 23619 7440 23651
rect 7480 23619 7512 23651
rect 7552 23619 7584 23651
rect 7624 23619 7656 23651
rect 7696 23619 7728 23651
rect 7768 23619 7800 23651
rect 7840 23619 7872 23651
rect 7912 23619 7944 23651
rect 7984 23619 8016 23651
rect 8056 23619 8088 23651
rect 8128 23619 8160 23651
rect 8200 23619 8232 23651
rect 8272 23619 8304 23651
rect 8344 23619 8376 23651
rect 8416 23619 8448 23651
rect 8488 23619 8520 23651
rect 8560 23619 8592 23651
rect 8632 23619 8664 23651
rect 8704 23619 8736 23651
rect 8776 23619 8808 23651
rect 8848 23619 8880 23651
rect 8920 23619 8952 23651
rect 8992 23619 9024 23651
rect 9064 23619 9096 23651
rect 9136 23619 9168 23651
rect 9208 23619 9240 23651
rect 9280 23619 9312 23651
rect 9352 23619 9384 23651
rect 9424 23619 9456 23651
rect 9496 23619 9528 23651
rect 9568 23619 9600 23651
rect 9640 23619 9672 23651
rect 9712 23619 9744 23651
rect 9784 23619 9816 23651
rect 9856 23619 9888 23651
rect 9928 23619 9960 23651
rect 10000 23619 10032 23651
rect 10072 23619 10104 23651
rect 10144 23619 10176 23651
rect 10216 23619 10248 23651
rect 10288 23619 10320 23651
rect 10360 23619 10392 23651
rect 10432 23619 10464 23651
rect 10504 23619 10536 23651
rect 10576 23619 10608 23651
rect 10648 23619 10680 23651
rect 10720 23619 10752 23651
rect 10792 23619 10824 23651
rect 10864 23619 10896 23651
rect 10936 23619 10968 23651
rect 11008 23619 11040 23651
rect 11080 23619 11112 23651
rect 11152 23619 11184 23651
rect 11224 23619 11256 23651
rect 11296 23619 11328 23651
rect 11368 23619 11400 23651
rect 11440 23619 11472 23651
rect 11512 23619 11544 23651
rect 11584 23619 11616 23651
rect 11656 23619 11688 23651
rect 11728 23619 11760 23651
rect 11800 23619 11832 23651
rect 11872 23619 11904 23651
rect 11944 23619 11976 23651
rect 12016 23619 12048 23651
rect 12088 23619 12120 23651
rect 12160 23619 12192 23651
rect 12232 23619 12264 23651
rect 12304 23619 12336 23651
rect 12376 23619 12408 23651
rect 12448 23619 12480 23651
rect 12520 23619 12552 23651
rect 12592 23619 12624 23651
rect 12664 23619 12696 23651
rect 12736 23619 12768 23651
rect 12808 23619 12840 23651
rect 12880 23619 12912 23651
rect 12952 23619 12984 23651
rect 13024 23619 13056 23651
rect 13096 23619 13128 23651
rect 13168 23619 13200 23651
rect 13240 23619 13272 23651
rect 13312 23619 13344 23651
rect 13384 23619 13416 23651
rect 13456 23619 13488 23651
rect 13528 23619 13560 23651
rect 13600 23619 13632 23651
rect 13672 23619 13704 23651
rect 13744 23619 13776 23651
rect 13816 23619 13848 23651
rect 13888 23619 13920 23651
rect 13960 23619 13992 23651
rect 14032 23619 14064 23651
rect 14104 23619 14136 23651
rect 14176 23619 14208 23651
rect 14248 23619 14280 23651
rect 14320 23619 14352 23651
rect 14392 23619 14424 23651
rect 14464 23619 14496 23651
rect 14536 23619 14568 23651
rect 14608 23619 14640 23651
rect 14680 23619 14712 23651
rect 14752 23619 14784 23651
rect 14824 23619 14856 23651
rect 14896 23619 14928 23651
rect 14968 23619 15000 23651
rect 15040 23619 15072 23651
rect 15112 23619 15144 23651
rect 15184 23619 15216 23651
rect 15256 23619 15288 23651
rect 15328 23619 15360 23651
rect 15400 23619 15432 23651
rect 15472 23619 15504 23651
rect 15544 23619 15576 23651
rect 15616 23619 15648 23651
rect 15688 23619 15720 23651
rect 15760 23619 15792 23651
rect 15832 23619 15864 23651
rect 15904 23619 15936 23651
rect 64 23547 96 23579
rect 136 23547 168 23579
rect 208 23547 240 23579
rect 280 23547 312 23579
rect 352 23547 384 23579
rect 424 23547 456 23579
rect 496 23547 528 23579
rect 568 23547 600 23579
rect 640 23547 672 23579
rect 712 23547 744 23579
rect 784 23547 816 23579
rect 856 23547 888 23579
rect 928 23547 960 23579
rect 1000 23547 1032 23579
rect 1072 23547 1104 23579
rect 1144 23547 1176 23579
rect 1216 23547 1248 23579
rect 1288 23547 1320 23579
rect 1360 23547 1392 23579
rect 1432 23547 1464 23579
rect 1504 23547 1536 23579
rect 1576 23547 1608 23579
rect 1648 23547 1680 23579
rect 1720 23547 1752 23579
rect 1792 23547 1824 23579
rect 1864 23547 1896 23579
rect 1936 23547 1968 23579
rect 2008 23547 2040 23579
rect 2080 23547 2112 23579
rect 2152 23547 2184 23579
rect 2224 23547 2256 23579
rect 2296 23547 2328 23579
rect 2368 23547 2400 23579
rect 2440 23547 2472 23579
rect 2512 23547 2544 23579
rect 2584 23547 2616 23579
rect 2656 23547 2688 23579
rect 2728 23547 2760 23579
rect 2800 23547 2832 23579
rect 2872 23547 2904 23579
rect 2944 23547 2976 23579
rect 3016 23547 3048 23579
rect 3088 23547 3120 23579
rect 3160 23547 3192 23579
rect 3232 23547 3264 23579
rect 3304 23547 3336 23579
rect 3376 23547 3408 23579
rect 3448 23547 3480 23579
rect 3520 23547 3552 23579
rect 3592 23547 3624 23579
rect 3664 23547 3696 23579
rect 3736 23547 3768 23579
rect 3808 23547 3840 23579
rect 3880 23547 3912 23579
rect 3952 23547 3984 23579
rect 4024 23547 4056 23579
rect 4096 23547 4128 23579
rect 4168 23547 4200 23579
rect 4240 23547 4272 23579
rect 4312 23547 4344 23579
rect 4384 23547 4416 23579
rect 4456 23547 4488 23579
rect 4528 23547 4560 23579
rect 4600 23547 4632 23579
rect 4672 23547 4704 23579
rect 4744 23547 4776 23579
rect 4816 23547 4848 23579
rect 4888 23547 4920 23579
rect 4960 23547 4992 23579
rect 5032 23547 5064 23579
rect 5104 23547 5136 23579
rect 5176 23547 5208 23579
rect 5248 23547 5280 23579
rect 5320 23547 5352 23579
rect 5392 23547 5424 23579
rect 5464 23547 5496 23579
rect 5536 23547 5568 23579
rect 5608 23547 5640 23579
rect 5680 23547 5712 23579
rect 5752 23547 5784 23579
rect 5824 23547 5856 23579
rect 5896 23547 5928 23579
rect 5968 23547 6000 23579
rect 6040 23547 6072 23579
rect 6112 23547 6144 23579
rect 6184 23547 6216 23579
rect 6256 23547 6288 23579
rect 6328 23547 6360 23579
rect 6400 23547 6432 23579
rect 6472 23547 6504 23579
rect 6544 23547 6576 23579
rect 6616 23547 6648 23579
rect 6688 23547 6720 23579
rect 6760 23547 6792 23579
rect 6832 23547 6864 23579
rect 6904 23547 6936 23579
rect 6976 23547 7008 23579
rect 7048 23547 7080 23579
rect 7120 23547 7152 23579
rect 7192 23547 7224 23579
rect 7264 23547 7296 23579
rect 7336 23547 7368 23579
rect 7408 23547 7440 23579
rect 7480 23547 7512 23579
rect 7552 23547 7584 23579
rect 7624 23547 7656 23579
rect 7696 23547 7728 23579
rect 7768 23547 7800 23579
rect 7840 23547 7872 23579
rect 7912 23547 7944 23579
rect 7984 23547 8016 23579
rect 8056 23547 8088 23579
rect 8128 23547 8160 23579
rect 8200 23547 8232 23579
rect 8272 23547 8304 23579
rect 8344 23547 8376 23579
rect 8416 23547 8448 23579
rect 8488 23547 8520 23579
rect 8560 23547 8592 23579
rect 8632 23547 8664 23579
rect 8704 23547 8736 23579
rect 8776 23547 8808 23579
rect 8848 23547 8880 23579
rect 8920 23547 8952 23579
rect 8992 23547 9024 23579
rect 9064 23547 9096 23579
rect 9136 23547 9168 23579
rect 9208 23547 9240 23579
rect 9280 23547 9312 23579
rect 9352 23547 9384 23579
rect 9424 23547 9456 23579
rect 9496 23547 9528 23579
rect 9568 23547 9600 23579
rect 9640 23547 9672 23579
rect 9712 23547 9744 23579
rect 9784 23547 9816 23579
rect 9856 23547 9888 23579
rect 9928 23547 9960 23579
rect 10000 23547 10032 23579
rect 10072 23547 10104 23579
rect 10144 23547 10176 23579
rect 10216 23547 10248 23579
rect 10288 23547 10320 23579
rect 10360 23547 10392 23579
rect 10432 23547 10464 23579
rect 10504 23547 10536 23579
rect 10576 23547 10608 23579
rect 10648 23547 10680 23579
rect 10720 23547 10752 23579
rect 10792 23547 10824 23579
rect 10864 23547 10896 23579
rect 10936 23547 10968 23579
rect 11008 23547 11040 23579
rect 11080 23547 11112 23579
rect 11152 23547 11184 23579
rect 11224 23547 11256 23579
rect 11296 23547 11328 23579
rect 11368 23547 11400 23579
rect 11440 23547 11472 23579
rect 11512 23547 11544 23579
rect 11584 23547 11616 23579
rect 11656 23547 11688 23579
rect 11728 23547 11760 23579
rect 11800 23547 11832 23579
rect 11872 23547 11904 23579
rect 11944 23547 11976 23579
rect 12016 23547 12048 23579
rect 12088 23547 12120 23579
rect 12160 23547 12192 23579
rect 12232 23547 12264 23579
rect 12304 23547 12336 23579
rect 12376 23547 12408 23579
rect 12448 23547 12480 23579
rect 12520 23547 12552 23579
rect 12592 23547 12624 23579
rect 12664 23547 12696 23579
rect 12736 23547 12768 23579
rect 12808 23547 12840 23579
rect 12880 23547 12912 23579
rect 12952 23547 12984 23579
rect 13024 23547 13056 23579
rect 13096 23547 13128 23579
rect 13168 23547 13200 23579
rect 13240 23547 13272 23579
rect 13312 23547 13344 23579
rect 13384 23547 13416 23579
rect 13456 23547 13488 23579
rect 13528 23547 13560 23579
rect 13600 23547 13632 23579
rect 13672 23547 13704 23579
rect 13744 23547 13776 23579
rect 13816 23547 13848 23579
rect 13888 23547 13920 23579
rect 13960 23547 13992 23579
rect 14032 23547 14064 23579
rect 14104 23547 14136 23579
rect 14176 23547 14208 23579
rect 14248 23547 14280 23579
rect 14320 23547 14352 23579
rect 14392 23547 14424 23579
rect 14464 23547 14496 23579
rect 14536 23547 14568 23579
rect 14608 23547 14640 23579
rect 14680 23547 14712 23579
rect 14752 23547 14784 23579
rect 14824 23547 14856 23579
rect 14896 23547 14928 23579
rect 14968 23547 15000 23579
rect 15040 23547 15072 23579
rect 15112 23547 15144 23579
rect 15184 23547 15216 23579
rect 15256 23547 15288 23579
rect 15328 23547 15360 23579
rect 15400 23547 15432 23579
rect 15472 23547 15504 23579
rect 15544 23547 15576 23579
rect 15616 23547 15648 23579
rect 15688 23547 15720 23579
rect 15760 23547 15792 23579
rect 15832 23547 15864 23579
rect 15904 23547 15936 23579
rect 64 23475 96 23507
rect 136 23475 168 23507
rect 208 23475 240 23507
rect 280 23475 312 23507
rect 352 23475 384 23507
rect 424 23475 456 23507
rect 496 23475 528 23507
rect 568 23475 600 23507
rect 640 23475 672 23507
rect 712 23475 744 23507
rect 784 23475 816 23507
rect 856 23475 888 23507
rect 928 23475 960 23507
rect 1000 23475 1032 23507
rect 1072 23475 1104 23507
rect 1144 23475 1176 23507
rect 1216 23475 1248 23507
rect 1288 23475 1320 23507
rect 1360 23475 1392 23507
rect 1432 23475 1464 23507
rect 1504 23475 1536 23507
rect 1576 23475 1608 23507
rect 1648 23475 1680 23507
rect 1720 23475 1752 23507
rect 1792 23475 1824 23507
rect 1864 23475 1896 23507
rect 1936 23475 1968 23507
rect 2008 23475 2040 23507
rect 2080 23475 2112 23507
rect 2152 23475 2184 23507
rect 2224 23475 2256 23507
rect 2296 23475 2328 23507
rect 2368 23475 2400 23507
rect 2440 23475 2472 23507
rect 2512 23475 2544 23507
rect 2584 23475 2616 23507
rect 2656 23475 2688 23507
rect 2728 23475 2760 23507
rect 2800 23475 2832 23507
rect 2872 23475 2904 23507
rect 2944 23475 2976 23507
rect 3016 23475 3048 23507
rect 3088 23475 3120 23507
rect 3160 23475 3192 23507
rect 3232 23475 3264 23507
rect 3304 23475 3336 23507
rect 3376 23475 3408 23507
rect 3448 23475 3480 23507
rect 3520 23475 3552 23507
rect 3592 23475 3624 23507
rect 3664 23475 3696 23507
rect 3736 23475 3768 23507
rect 3808 23475 3840 23507
rect 3880 23475 3912 23507
rect 3952 23475 3984 23507
rect 4024 23475 4056 23507
rect 4096 23475 4128 23507
rect 4168 23475 4200 23507
rect 4240 23475 4272 23507
rect 4312 23475 4344 23507
rect 4384 23475 4416 23507
rect 4456 23475 4488 23507
rect 4528 23475 4560 23507
rect 4600 23475 4632 23507
rect 4672 23475 4704 23507
rect 4744 23475 4776 23507
rect 4816 23475 4848 23507
rect 4888 23475 4920 23507
rect 4960 23475 4992 23507
rect 5032 23475 5064 23507
rect 5104 23475 5136 23507
rect 5176 23475 5208 23507
rect 5248 23475 5280 23507
rect 5320 23475 5352 23507
rect 5392 23475 5424 23507
rect 5464 23475 5496 23507
rect 5536 23475 5568 23507
rect 5608 23475 5640 23507
rect 5680 23475 5712 23507
rect 5752 23475 5784 23507
rect 5824 23475 5856 23507
rect 5896 23475 5928 23507
rect 5968 23475 6000 23507
rect 6040 23475 6072 23507
rect 6112 23475 6144 23507
rect 6184 23475 6216 23507
rect 6256 23475 6288 23507
rect 6328 23475 6360 23507
rect 6400 23475 6432 23507
rect 6472 23475 6504 23507
rect 6544 23475 6576 23507
rect 6616 23475 6648 23507
rect 6688 23475 6720 23507
rect 6760 23475 6792 23507
rect 6832 23475 6864 23507
rect 6904 23475 6936 23507
rect 6976 23475 7008 23507
rect 7048 23475 7080 23507
rect 7120 23475 7152 23507
rect 7192 23475 7224 23507
rect 7264 23475 7296 23507
rect 7336 23475 7368 23507
rect 7408 23475 7440 23507
rect 7480 23475 7512 23507
rect 7552 23475 7584 23507
rect 7624 23475 7656 23507
rect 7696 23475 7728 23507
rect 7768 23475 7800 23507
rect 7840 23475 7872 23507
rect 7912 23475 7944 23507
rect 7984 23475 8016 23507
rect 8056 23475 8088 23507
rect 8128 23475 8160 23507
rect 8200 23475 8232 23507
rect 8272 23475 8304 23507
rect 8344 23475 8376 23507
rect 8416 23475 8448 23507
rect 8488 23475 8520 23507
rect 8560 23475 8592 23507
rect 8632 23475 8664 23507
rect 8704 23475 8736 23507
rect 8776 23475 8808 23507
rect 8848 23475 8880 23507
rect 8920 23475 8952 23507
rect 8992 23475 9024 23507
rect 9064 23475 9096 23507
rect 9136 23475 9168 23507
rect 9208 23475 9240 23507
rect 9280 23475 9312 23507
rect 9352 23475 9384 23507
rect 9424 23475 9456 23507
rect 9496 23475 9528 23507
rect 9568 23475 9600 23507
rect 9640 23475 9672 23507
rect 9712 23475 9744 23507
rect 9784 23475 9816 23507
rect 9856 23475 9888 23507
rect 9928 23475 9960 23507
rect 10000 23475 10032 23507
rect 10072 23475 10104 23507
rect 10144 23475 10176 23507
rect 10216 23475 10248 23507
rect 10288 23475 10320 23507
rect 10360 23475 10392 23507
rect 10432 23475 10464 23507
rect 10504 23475 10536 23507
rect 10576 23475 10608 23507
rect 10648 23475 10680 23507
rect 10720 23475 10752 23507
rect 10792 23475 10824 23507
rect 10864 23475 10896 23507
rect 10936 23475 10968 23507
rect 11008 23475 11040 23507
rect 11080 23475 11112 23507
rect 11152 23475 11184 23507
rect 11224 23475 11256 23507
rect 11296 23475 11328 23507
rect 11368 23475 11400 23507
rect 11440 23475 11472 23507
rect 11512 23475 11544 23507
rect 11584 23475 11616 23507
rect 11656 23475 11688 23507
rect 11728 23475 11760 23507
rect 11800 23475 11832 23507
rect 11872 23475 11904 23507
rect 11944 23475 11976 23507
rect 12016 23475 12048 23507
rect 12088 23475 12120 23507
rect 12160 23475 12192 23507
rect 12232 23475 12264 23507
rect 12304 23475 12336 23507
rect 12376 23475 12408 23507
rect 12448 23475 12480 23507
rect 12520 23475 12552 23507
rect 12592 23475 12624 23507
rect 12664 23475 12696 23507
rect 12736 23475 12768 23507
rect 12808 23475 12840 23507
rect 12880 23475 12912 23507
rect 12952 23475 12984 23507
rect 13024 23475 13056 23507
rect 13096 23475 13128 23507
rect 13168 23475 13200 23507
rect 13240 23475 13272 23507
rect 13312 23475 13344 23507
rect 13384 23475 13416 23507
rect 13456 23475 13488 23507
rect 13528 23475 13560 23507
rect 13600 23475 13632 23507
rect 13672 23475 13704 23507
rect 13744 23475 13776 23507
rect 13816 23475 13848 23507
rect 13888 23475 13920 23507
rect 13960 23475 13992 23507
rect 14032 23475 14064 23507
rect 14104 23475 14136 23507
rect 14176 23475 14208 23507
rect 14248 23475 14280 23507
rect 14320 23475 14352 23507
rect 14392 23475 14424 23507
rect 14464 23475 14496 23507
rect 14536 23475 14568 23507
rect 14608 23475 14640 23507
rect 14680 23475 14712 23507
rect 14752 23475 14784 23507
rect 14824 23475 14856 23507
rect 14896 23475 14928 23507
rect 14968 23475 15000 23507
rect 15040 23475 15072 23507
rect 15112 23475 15144 23507
rect 15184 23475 15216 23507
rect 15256 23475 15288 23507
rect 15328 23475 15360 23507
rect 15400 23475 15432 23507
rect 15472 23475 15504 23507
rect 15544 23475 15576 23507
rect 15616 23475 15648 23507
rect 15688 23475 15720 23507
rect 15760 23475 15792 23507
rect 15832 23475 15864 23507
rect 15904 23475 15936 23507
rect 64 23403 96 23435
rect 136 23403 168 23435
rect 208 23403 240 23435
rect 280 23403 312 23435
rect 352 23403 384 23435
rect 424 23403 456 23435
rect 496 23403 528 23435
rect 568 23403 600 23435
rect 640 23403 672 23435
rect 712 23403 744 23435
rect 784 23403 816 23435
rect 856 23403 888 23435
rect 928 23403 960 23435
rect 1000 23403 1032 23435
rect 1072 23403 1104 23435
rect 1144 23403 1176 23435
rect 1216 23403 1248 23435
rect 1288 23403 1320 23435
rect 1360 23403 1392 23435
rect 1432 23403 1464 23435
rect 1504 23403 1536 23435
rect 1576 23403 1608 23435
rect 1648 23403 1680 23435
rect 1720 23403 1752 23435
rect 1792 23403 1824 23435
rect 1864 23403 1896 23435
rect 1936 23403 1968 23435
rect 2008 23403 2040 23435
rect 2080 23403 2112 23435
rect 2152 23403 2184 23435
rect 2224 23403 2256 23435
rect 2296 23403 2328 23435
rect 2368 23403 2400 23435
rect 2440 23403 2472 23435
rect 2512 23403 2544 23435
rect 2584 23403 2616 23435
rect 2656 23403 2688 23435
rect 2728 23403 2760 23435
rect 2800 23403 2832 23435
rect 2872 23403 2904 23435
rect 2944 23403 2976 23435
rect 3016 23403 3048 23435
rect 3088 23403 3120 23435
rect 3160 23403 3192 23435
rect 3232 23403 3264 23435
rect 3304 23403 3336 23435
rect 3376 23403 3408 23435
rect 3448 23403 3480 23435
rect 3520 23403 3552 23435
rect 3592 23403 3624 23435
rect 3664 23403 3696 23435
rect 3736 23403 3768 23435
rect 3808 23403 3840 23435
rect 3880 23403 3912 23435
rect 3952 23403 3984 23435
rect 4024 23403 4056 23435
rect 4096 23403 4128 23435
rect 4168 23403 4200 23435
rect 4240 23403 4272 23435
rect 4312 23403 4344 23435
rect 4384 23403 4416 23435
rect 4456 23403 4488 23435
rect 4528 23403 4560 23435
rect 4600 23403 4632 23435
rect 4672 23403 4704 23435
rect 4744 23403 4776 23435
rect 4816 23403 4848 23435
rect 4888 23403 4920 23435
rect 4960 23403 4992 23435
rect 5032 23403 5064 23435
rect 5104 23403 5136 23435
rect 5176 23403 5208 23435
rect 5248 23403 5280 23435
rect 5320 23403 5352 23435
rect 5392 23403 5424 23435
rect 5464 23403 5496 23435
rect 5536 23403 5568 23435
rect 5608 23403 5640 23435
rect 5680 23403 5712 23435
rect 5752 23403 5784 23435
rect 5824 23403 5856 23435
rect 5896 23403 5928 23435
rect 5968 23403 6000 23435
rect 6040 23403 6072 23435
rect 6112 23403 6144 23435
rect 6184 23403 6216 23435
rect 6256 23403 6288 23435
rect 6328 23403 6360 23435
rect 6400 23403 6432 23435
rect 6472 23403 6504 23435
rect 6544 23403 6576 23435
rect 6616 23403 6648 23435
rect 6688 23403 6720 23435
rect 6760 23403 6792 23435
rect 6832 23403 6864 23435
rect 6904 23403 6936 23435
rect 6976 23403 7008 23435
rect 7048 23403 7080 23435
rect 7120 23403 7152 23435
rect 7192 23403 7224 23435
rect 7264 23403 7296 23435
rect 7336 23403 7368 23435
rect 7408 23403 7440 23435
rect 7480 23403 7512 23435
rect 7552 23403 7584 23435
rect 7624 23403 7656 23435
rect 7696 23403 7728 23435
rect 7768 23403 7800 23435
rect 7840 23403 7872 23435
rect 7912 23403 7944 23435
rect 7984 23403 8016 23435
rect 8056 23403 8088 23435
rect 8128 23403 8160 23435
rect 8200 23403 8232 23435
rect 8272 23403 8304 23435
rect 8344 23403 8376 23435
rect 8416 23403 8448 23435
rect 8488 23403 8520 23435
rect 8560 23403 8592 23435
rect 8632 23403 8664 23435
rect 8704 23403 8736 23435
rect 8776 23403 8808 23435
rect 8848 23403 8880 23435
rect 8920 23403 8952 23435
rect 8992 23403 9024 23435
rect 9064 23403 9096 23435
rect 9136 23403 9168 23435
rect 9208 23403 9240 23435
rect 9280 23403 9312 23435
rect 9352 23403 9384 23435
rect 9424 23403 9456 23435
rect 9496 23403 9528 23435
rect 9568 23403 9600 23435
rect 9640 23403 9672 23435
rect 9712 23403 9744 23435
rect 9784 23403 9816 23435
rect 9856 23403 9888 23435
rect 9928 23403 9960 23435
rect 10000 23403 10032 23435
rect 10072 23403 10104 23435
rect 10144 23403 10176 23435
rect 10216 23403 10248 23435
rect 10288 23403 10320 23435
rect 10360 23403 10392 23435
rect 10432 23403 10464 23435
rect 10504 23403 10536 23435
rect 10576 23403 10608 23435
rect 10648 23403 10680 23435
rect 10720 23403 10752 23435
rect 10792 23403 10824 23435
rect 10864 23403 10896 23435
rect 10936 23403 10968 23435
rect 11008 23403 11040 23435
rect 11080 23403 11112 23435
rect 11152 23403 11184 23435
rect 11224 23403 11256 23435
rect 11296 23403 11328 23435
rect 11368 23403 11400 23435
rect 11440 23403 11472 23435
rect 11512 23403 11544 23435
rect 11584 23403 11616 23435
rect 11656 23403 11688 23435
rect 11728 23403 11760 23435
rect 11800 23403 11832 23435
rect 11872 23403 11904 23435
rect 11944 23403 11976 23435
rect 12016 23403 12048 23435
rect 12088 23403 12120 23435
rect 12160 23403 12192 23435
rect 12232 23403 12264 23435
rect 12304 23403 12336 23435
rect 12376 23403 12408 23435
rect 12448 23403 12480 23435
rect 12520 23403 12552 23435
rect 12592 23403 12624 23435
rect 12664 23403 12696 23435
rect 12736 23403 12768 23435
rect 12808 23403 12840 23435
rect 12880 23403 12912 23435
rect 12952 23403 12984 23435
rect 13024 23403 13056 23435
rect 13096 23403 13128 23435
rect 13168 23403 13200 23435
rect 13240 23403 13272 23435
rect 13312 23403 13344 23435
rect 13384 23403 13416 23435
rect 13456 23403 13488 23435
rect 13528 23403 13560 23435
rect 13600 23403 13632 23435
rect 13672 23403 13704 23435
rect 13744 23403 13776 23435
rect 13816 23403 13848 23435
rect 13888 23403 13920 23435
rect 13960 23403 13992 23435
rect 14032 23403 14064 23435
rect 14104 23403 14136 23435
rect 14176 23403 14208 23435
rect 14248 23403 14280 23435
rect 14320 23403 14352 23435
rect 14392 23403 14424 23435
rect 14464 23403 14496 23435
rect 14536 23403 14568 23435
rect 14608 23403 14640 23435
rect 14680 23403 14712 23435
rect 14752 23403 14784 23435
rect 14824 23403 14856 23435
rect 14896 23403 14928 23435
rect 14968 23403 15000 23435
rect 15040 23403 15072 23435
rect 15112 23403 15144 23435
rect 15184 23403 15216 23435
rect 15256 23403 15288 23435
rect 15328 23403 15360 23435
rect 15400 23403 15432 23435
rect 15472 23403 15504 23435
rect 15544 23403 15576 23435
rect 15616 23403 15648 23435
rect 15688 23403 15720 23435
rect 15760 23403 15792 23435
rect 15832 23403 15864 23435
rect 15904 23403 15936 23435
rect 64 23331 96 23363
rect 136 23331 168 23363
rect 208 23331 240 23363
rect 280 23331 312 23363
rect 352 23331 384 23363
rect 424 23331 456 23363
rect 496 23331 528 23363
rect 568 23331 600 23363
rect 640 23331 672 23363
rect 712 23331 744 23363
rect 784 23331 816 23363
rect 856 23331 888 23363
rect 928 23331 960 23363
rect 1000 23331 1032 23363
rect 1072 23331 1104 23363
rect 1144 23331 1176 23363
rect 1216 23331 1248 23363
rect 1288 23331 1320 23363
rect 1360 23331 1392 23363
rect 1432 23331 1464 23363
rect 1504 23331 1536 23363
rect 1576 23331 1608 23363
rect 1648 23331 1680 23363
rect 1720 23331 1752 23363
rect 1792 23331 1824 23363
rect 1864 23331 1896 23363
rect 1936 23331 1968 23363
rect 2008 23331 2040 23363
rect 2080 23331 2112 23363
rect 2152 23331 2184 23363
rect 2224 23331 2256 23363
rect 2296 23331 2328 23363
rect 2368 23331 2400 23363
rect 2440 23331 2472 23363
rect 2512 23331 2544 23363
rect 2584 23331 2616 23363
rect 2656 23331 2688 23363
rect 2728 23331 2760 23363
rect 2800 23331 2832 23363
rect 2872 23331 2904 23363
rect 2944 23331 2976 23363
rect 3016 23331 3048 23363
rect 3088 23331 3120 23363
rect 3160 23331 3192 23363
rect 3232 23331 3264 23363
rect 3304 23331 3336 23363
rect 3376 23331 3408 23363
rect 3448 23331 3480 23363
rect 3520 23331 3552 23363
rect 3592 23331 3624 23363
rect 3664 23331 3696 23363
rect 3736 23331 3768 23363
rect 3808 23331 3840 23363
rect 3880 23331 3912 23363
rect 3952 23331 3984 23363
rect 4024 23331 4056 23363
rect 4096 23331 4128 23363
rect 4168 23331 4200 23363
rect 4240 23331 4272 23363
rect 4312 23331 4344 23363
rect 4384 23331 4416 23363
rect 4456 23331 4488 23363
rect 4528 23331 4560 23363
rect 4600 23331 4632 23363
rect 4672 23331 4704 23363
rect 4744 23331 4776 23363
rect 4816 23331 4848 23363
rect 4888 23331 4920 23363
rect 4960 23331 4992 23363
rect 5032 23331 5064 23363
rect 5104 23331 5136 23363
rect 5176 23331 5208 23363
rect 5248 23331 5280 23363
rect 5320 23331 5352 23363
rect 5392 23331 5424 23363
rect 5464 23331 5496 23363
rect 5536 23331 5568 23363
rect 5608 23331 5640 23363
rect 5680 23331 5712 23363
rect 5752 23331 5784 23363
rect 5824 23331 5856 23363
rect 5896 23331 5928 23363
rect 5968 23331 6000 23363
rect 6040 23331 6072 23363
rect 6112 23331 6144 23363
rect 6184 23331 6216 23363
rect 6256 23331 6288 23363
rect 6328 23331 6360 23363
rect 6400 23331 6432 23363
rect 6472 23331 6504 23363
rect 6544 23331 6576 23363
rect 6616 23331 6648 23363
rect 6688 23331 6720 23363
rect 6760 23331 6792 23363
rect 6832 23331 6864 23363
rect 6904 23331 6936 23363
rect 6976 23331 7008 23363
rect 7048 23331 7080 23363
rect 7120 23331 7152 23363
rect 7192 23331 7224 23363
rect 7264 23331 7296 23363
rect 7336 23331 7368 23363
rect 7408 23331 7440 23363
rect 7480 23331 7512 23363
rect 7552 23331 7584 23363
rect 7624 23331 7656 23363
rect 7696 23331 7728 23363
rect 7768 23331 7800 23363
rect 7840 23331 7872 23363
rect 7912 23331 7944 23363
rect 7984 23331 8016 23363
rect 8056 23331 8088 23363
rect 8128 23331 8160 23363
rect 8200 23331 8232 23363
rect 8272 23331 8304 23363
rect 8344 23331 8376 23363
rect 8416 23331 8448 23363
rect 8488 23331 8520 23363
rect 8560 23331 8592 23363
rect 8632 23331 8664 23363
rect 8704 23331 8736 23363
rect 8776 23331 8808 23363
rect 8848 23331 8880 23363
rect 8920 23331 8952 23363
rect 8992 23331 9024 23363
rect 9064 23331 9096 23363
rect 9136 23331 9168 23363
rect 9208 23331 9240 23363
rect 9280 23331 9312 23363
rect 9352 23331 9384 23363
rect 9424 23331 9456 23363
rect 9496 23331 9528 23363
rect 9568 23331 9600 23363
rect 9640 23331 9672 23363
rect 9712 23331 9744 23363
rect 9784 23331 9816 23363
rect 9856 23331 9888 23363
rect 9928 23331 9960 23363
rect 10000 23331 10032 23363
rect 10072 23331 10104 23363
rect 10144 23331 10176 23363
rect 10216 23331 10248 23363
rect 10288 23331 10320 23363
rect 10360 23331 10392 23363
rect 10432 23331 10464 23363
rect 10504 23331 10536 23363
rect 10576 23331 10608 23363
rect 10648 23331 10680 23363
rect 10720 23331 10752 23363
rect 10792 23331 10824 23363
rect 10864 23331 10896 23363
rect 10936 23331 10968 23363
rect 11008 23331 11040 23363
rect 11080 23331 11112 23363
rect 11152 23331 11184 23363
rect 11224 23331 11256 23363
rect 11296 23331 11328 23363
rect 11368 23331 11400 23363
rect 11440 23331 11472 23363
rect 11512 23331 11544 23363
rect 11584 23331 11616 23363
rect 11656 23331 11688 23363
rect 11728 23331 11760 23363
rect 11800 23331 11832 23363
rect 11872 23331 11904 23363
rect 11944 23331 11976 23363
rect 12016 23331 12048 23363
rect 12088 23331 12120 23363
rect 12160 23331 12192 23363
rect 12232 23331 12264 23363
rect 12304 23331 12336 23363
rect 12376 23331 12408 23363
rect 12448 23331 12480 23363
rect 12520 23331 12552 23363
rect 12592 23331 12624 23363
rect 12664 23331 12696 23363
rect 12736 23331 12768 23363
rect 12808 23331 12840 23363
rect 12880 23331 12912 23363
rect 12952 23331 12984 23363
rect 13024 23331 13056 23363
rect 13096 23331 13128 23363
rect 13168 23331 13200 23363
rect 13240 23331 13272 23363
rect 13312 23331 13344 23363
rect 13384 23331 13416 23363
rect 13456 23331 13488 23363
rect 13528 23331 13560 23363
rect 13600 23331 13632 23363
rect 13672 23331 13704 23363
rect 13744 23331 13776 23363
rect 13816 23331 13848 23363
rect 13888 23331 13920 23363
rect 13960 23331 13992 23363
rect 14032 23331 14064 23363
rect 14104 23331 14136 23363
rect 14176 23331 14208 23363
rect 14248 23331 14280 23363
rect 14320 23331 14352 23363
rect 14392 23331 14424 23363
rect 14464 23331 14496 23363
rect 14536 23331 14568 23363
rect 14608 23331 14640 23363
rect 14680 23331 14712 23363
rect 14752 23331 14784 23363
rect 14824 23331 14856 23363
rect 14896 23331 14928 23363
rect 14968 23331 15000 23363
rect 15040 23331 15072 23363
rect 15112 23331 15144 23363
rect 15184 23331 15216 23363
rect 15256 23331 15288 23363
rect 15328 23331 15360 23363
rect 15400 23331 15432 23363
rect 15472 23331 15504 23363
rect 15544 23331 15576 23363
rect 15616 23331 15648 23363
rect 15688 23331 15720 23363
rect 15760 23331 15792 23363
rect 15832 23331 15864 23363
rect 15904 23331 15936 23363
rect 64 23259 96 23291
rect 136 23259 168 23291
rect 208 23259 240 23291
rect 280 23259 312 23291
rect 352 23259 384 23291
rect 424 23259 456 23291
rect 496 23259 528 23291
rect 568 23259 600 23291
rect 640 23259 672 23291
rect 712 23259 744 23291
rect 784 23259 816 23291
rect 856 23259 888 23291
rect 928 23259 960 23291
rect 1000 23259 1032 23291
rect 1072 23259 1104 23291
rect 1144 23259 1176 23291
rect 1216 23259 1248 23291
rect 1288 23259 1320 23291
rect 1360 23259 1392 23291
rect 1432 23259 1464 23291
rect 1504 23259 1536 23291
rect 1576 23259 1608 23291
rect 1648 23259 1680 23291
rect 1720 23259 1752 23291
rect 1792 23259 1824 23291
rect 1864 23259 1896 23291
rect 1936 23259 1968 23291
rect 2008 23259 2040 23291
rect 2080 23259 2112 23291
rect 2152 23259 2184 23291
rect 2224 23259 2256 23291
rect 2296 23259 2328 23291
rect 2368 23259 2400 23291
rect 2440 23259 2472 23291
rect 2512 23259 2544 23291
rect 2584 23259 2616 23291
rect 2656 23259 2688 23291
rect 2728 23259 2760 23291
rect 2800 23259 2832 23291
rect 2872 23259 2904 23291
rect 2944 23259 2976 23291
rect 3016 23259 3048 23291
rect 3088 23259 3120 23291
rect 3160 23259 3192 23291
rect 3232 23259 3264 23291
rect 3304 23259 3336 23291
rect 3376 23259 3408 23291
rect 3448 23259 3480 23291
rect 3520 23259 3552 23291
rect 3592 23259 3624 23291
rect 3664 23259 3696 23291
rect 3736 23259 3768 23291
rect 3808 23259 3840 23291
rect 3880 23259 3912 23291
rect 3952 23259 3984 23291
rect 4024 23259 4056 23291
rect 4096 23259 4128 23291
rect 4168 23259 4200 23291
rect 4240 23259 4272 23291
rect 4312 23259 4344 23291
rect 4384 23259 4416 23291
rect 4456 23259 4488 23291
rect 4528 23259 4560 23291
rect 4600 23259 4632 23291
rect 4672 23259 4704 23291
rect 4744 23259 4776 23291
rect 4816 23259 4848 23291
rect 4888 23259 4920 23291
rect 4960 23259 4992 23291
rect 5032 23259 5064 23291
rect 5104 23259 5136 23291
rect 5176 23259 5208 23291
rect 5248 23259 5280 23291
rect 5320 23259 5352 23291
rect 5392 23259 5424 23291
rect 5464 23259 5496 23291
rect 5536 23259 5568 23291
rect 5608 23259 5640 23291
rect 5680 23259 5712 23291
rect 5752 23259 5784 23291
rect 5824 23259 5856 23291
rect 5896 23259 5928 23291
rect 5968 23259 6000 23291
rect 6040 23259 6072 23291
rect 6112 23259 6144 23291
rect 6184 23259 6216 23291
rect 6256 23259 6288 23291
rect 6328 23259 6360 23291
rect 6400 23259 6432 23291
rect 6472 23259 6504 23291
rect 6544 23259 6576 23291
rect 6616 23259 6648 23291
rect 6688 23259 6720 23291
rect 6760 23259 6792 23291
rect 6832 23259 6864 23291
rect 6904 23259 6936 23291
rect 6976 23259 7008 23291
rect 7048 23259 7080 23291
rect 7120 23259 7152 23291
rect 7192 23259 7224 23291
rect 7264 23259 7296 23291
rect 7336 23259 7368 23291
rect 7408 23259 7440 23291
rect 7480 23259 7512 23291
rect 7552 23259 7584 23291
rect 7624 23259 7656 23291
rect 7696 23259 7728 23291
rect 7768 23259 7800 23291
rect 7840 23259 7872 23291
rect 7912 23259 7944 23291
rect 7984 23259 8016 23291
rect 8056 23259 8088 23291
rect 8128 23259 8160 23291
rect 8200 23259 8232 23291
rect 8272 23259 8304 23291
rect 8344 23259 8376 23291
rect 8416 23259 8448 23291
rect 8488 23259 8520 23291
rect 8560 23259 8592 23291
rect 8632 23259 8664 23291
rect 8704 23259 8736 23291
rect 8776 23259 8808 23291
rect 8848 23259 8880 23291
rect 8920 23259 8952 23291
rect 8992 23259 9024 23291
rect 9064 23259 9096 23291
rect 9136 23259 9168 23291
rect 9208 23259 9240 23291
rect 9280 23259 9312 23291
rect 9352 23259 9384 23291
rect 9424 23259 9456 23291
rect 9496 23259 9528 23291
rect 9568 23259 9600 23291
rect 9640 23259 9672 23291
rect 9712 23259 9744 23291
rect 9784 23259 9816 23291
rect 9856 23259 9888 23291
rect 9928 23259 9960 23291
rect 10000 23259 10032 23291
rect 10072 23259 10104 23291
rect 10144 23259 10176 23291
rect 10216 23259 10248 23291
rect 10288 23259 10320 23291
rect 10360 23259 10392 23291
rect 10432 23259 10464 23291
rect 10504 23259 10536 23291
rect 10576 23259 10608 23291
rect 10648 23259 10680 23291
rect 10720 23259 10752 23291
rect 10792 23259 10824 23291
rect 10864 23259 10896 23291
rect 10936 23259 10968 23291
rect 11008 23259 11040 23291
rect 11080 23259 11112 23291
rect 11152 23259 11184 23291
rect 11224 23259 11256 23291
rect 11296 23259 11328 23291
rect 11368 23259 11400 23291
rect 11440 23259 11472 23291
rect 11512 23259 11544 23291
rect 11584 23259 11616 23291
rect 11656 23259 11688 23291
rect 11728 23259 11760 23291
rect 11800 23259 11832 23291
rect 11872 23259 11904 23291
rect 11944 23259 11976 23291
rect 12016 23259 12048 23291
rect 12088 23259 12120 23291
rect 12160 23259 12192 23291
rect 12232 23259 12264 23291
rect 12304 23259 12336 23291
rect 12376 23259 12408 23291
rect 12448 23259 12480 23291
rect 12520 23259 12552 23291
rect 12592 23259 12624 23291
rect 12664 23259 12696 23291
rect 12736 23259 12768 23291
rect 12808 23259 12840 23291
rect 12880 23259 12912 23291
rect 12952 23259 12984 23291
rect 13024 23259 13056 23291
rect 13096 23259 13128 23291
rect 13168 23259 13200 23291
rect 13240 23259 13272 23291
rect 13312 23259 13344 23291
rect 13384 23259 13416 23291
rect 13456 23259 13488 23291
rect 13528 23259 13560 23291
rect 13600 23259 13632 23291
rect 13672 23259 13704 23291
rect 13744 23259 13776 23291
rect 13816 23259 13848 23291
rect 13888 23259 13920 23291
rect 13960 23259 13992 23291
rect 14032 23259 14064 23291
rect 14104 23259 14136 23291
rect 14176 23259 14208 23291
rect 14248 23259 14280 23291
rect 14320 23259 14352 23291
rect 14392 23259 14424 23291
rect 14464 23259 14496 23291
rect 14536 23259 14568 23291
rect 14608 23259 14640 23291
rect 14680 23259 14712 23291
rect 14752 23259 14784 23291
rect 14824 23259 14856 23291
rect 14896 23259 14928 23291
rect 14968 23259 15000 23291
rect 15040 23259 15072 23291
rect 15112 23259 15144 23291
rect 15184 23259 15216 23291
rect 15256 23259 15288 23291
rect 15328 23259 15360 23291
rect 15400 23259 15432 23291
rect 15472 23259 15504 23291
rect 15544 23259 15576 23291
rect 15616 23259 15648 23291
rect 15688 23259 15720 23291
rect 15760 23259 15792 23291
rect 15832 23259 15864 23291
rect 15904 23259 15936 23291
rect 64 23187 96 23219
rect 136 23187 168 23219
rect 208 23187 240 23219
rect 280 23187 312 23219
rect 352 23187 384 23219
rect 424 23187 456 23219
rect 496 23187 528 23219
rect 568 23187 600 23219
rect 640 23187 672 23219
rect 712 23187 744 23219
rect 784 23187 816 23219
rect 856 23187 888 23219
rect 928 23187 960 23219
rect 1000 23187 1032 23219
rect 1072 23187 1104 23219
rect 1144 23187 1176 23219
rect 1216 23187 1248 23219
rect 1288 23187 1320 23219
rect 1360 23187 1392 23219
rect 1432 23187 1464 23219
rect 1504 23187 1536 23219
rect 1576 23187 1608 23219
rect 1648 23187 1680 23219
rect 1720 23187 1752 23219
rect 1792 23187 1824 23219
rect 1864 23187 1896 23219
rect 1936 23187 1968 23219
rect 2008 23187 2040 23219
rect 2080 23187 2112 23219
rect 2152 23187 2184 23219
rect 2224 23187 2256 23219
rect 2296 23187 2328 23219
rect 2368 23187 2400 23219
rect 2440 23187 2472 23219
rect 2512 23187 2544 23219
rect 2584 23187 2616 23219
rect 2656 23187 2688 23219
rect 2728 23187 2760 23219
rect 2800 23187 2832 23219
rect 2872 23187 2904 23219
rect 2944 23187 2976 23219
rect 3016 23187 3048 23219
rect 3088 23187 3120 23219
rect 3160 23187 3192 23219
rect 3232 23187 3264 23219
rect 3304 23187 3336 23219
rect 3376 23187 3408 23219
rect 3448 23187 3480 23219
rect 3520 23187 3552 23219
rect 3592 23187 3624 23219
rect 3664 23187 3696 23219
rect 3736 23187 3768 23219
rect 3808 23187 3840 23219
rect 3880 23187 3912 23219
rect 3952 23187 3984 23219
rect 4024 23187 4056 23219
rect 4096 23187 4128 23219
rect 4168 23187 4200 23219
rect 4240 23187 4272 23219
rect 4312 23187 4344 23219
rect 4384 23187 4416 23219
rect 4456 23187 4488 23219
rect 4528 23187 4560 23219
rect 4600 23187 4632 23219
rect 4672 23187 4704 23219
rect 4744 23187 4776 23219
rect 4816 23187 4848 23219
rect 4888 23187 4920 23219
rect 4960 23187 4992 23219
rect 5032 23187 5064 23219
rect 5104 23187 5136 23219
rect 5176 23187 5208 23219
rect 5248 23187 5280 23219
rect 5320 23187 5352 23219
rect 5392 23187 5424 23219
rect 5464 23187 5496 23219
rect 5536 23187 5568 23219
rect 5608 23187 5640 23219
rect 5680 23187 5712 23219
rect 5752 23187 5784 23219
rect 5824 23187 5856 23219
rect 5896 23187 5928 23219
rect 5968 23187 6000 23219
rect 6040 23187 6072 23219
rect 6112 23187 6144 23219
rect 6184 23187 6216 23219
rect 6256 23187 6288 23219
rect 6328 23187 6360 23219
rect 6400 23187 6432 23219
rect 6472 23187 6504 23219
rect 6544 23187 6576 23219
rect 6616 23187 6648 23219
rect 6688 23187 6720 23219
rect 6760 23187 6792 23219
rect 6832 23187 6864 23219
rect 6904 23187 6936 23219
rect 6976 23187 7008 23219
rect 7048 23187 7080 23219
rect 7120 23187 7152 23219
rect 7192 23187 7224 23219
rect 7264 23187 7296 23219
rect 7336 23187 7368 23219
rect 7408 23187 7440 23219
rect 7480 23187 7512 23219
rect 7552 23187 7584 23219
rect 7624 23187 7656 23219
rect 7696 23187 7728 23219
rect 7768 23187 7800 23219
rect 7840 23187 7872 23219
rect 7912 23187 7944 23219
rect 7984 23187 8016 23219
rect 8056 23187 8088 23219
rect 8128 23187 8160 23219
rect 8200 23187 8232 23219
rect 8272 23187 8304 23219
rect 8344 23187 8376 23219
rect 8416 23187 8448 23219
rect 8488 23187 8520 23219
rect 8560 23187 8592 23219
rect 8632 23187 8664 23219
rect 8704 23187 8736 23219
rect 8776 23187 8808 23219
rect 8848 23187 8880 23219
rect 8920 23187 8952 23219
rect 8992 23187 9024 23219
rect 9064 23187 9096 23219
rect 9136 23187 9168 23219
rect 9208 23187 9240 23219
rect 9280 23187 9312 23219
rect 9352 23187 9384 23219
rect 9424 23187 9456 23219
rect 9496 23187 9528 23219
rect 9568 23187 9600 23219
rect 9640 23187 9672 23219
rect 9712 23187 9744 23219
rect 9784 23187 9816 23219
rect 9856 23187 9888 23219
rect 9928 23187 9960 23219
rect 10000 23187 10032 23219
rect 10072 23187 10104 23219
rect 10144 23187 10176 23219
rect 10216 23187 10248 23219
rect 10288 23187 10320 23219
rect 10360 23187 10392 23219
rect 10432 23187 10464 23219
rect 10504 23187 10536 23219
rect 10576 23187 10608 23219
rect 10648 23187 10680 23219
rect 10720 23187 10752 23219
rect 10792 23187 10824 23219
rect 10864 23187 10896 23219
rect 10936 23187 10968 23219
rect 11008 23187 11040 23219
rect 11080 23187 11112 23219
rect 11152 23187 11184 23219
rect 11224 23187 11256 23219
rect 11296 23187 11328 23219
rect 11368 23187 11400 23219
rect 11440 23187 11472 23219
rect 11512 23187 11544 23219
rect 11584 23187 11616 23219
rect 11656 23187 11688 23219
rect 11728 23187 11760 23219
rect 11800 23187 11832 23219
rect 11872 23187 11904 23219
rect 11944 23187 11976 23219
rect 12016 23187 12048 23219
rect 12088 23187 12120 23219
rect 12160 23187 12192 23219
rect 12232 23187 12264 23219
rect 12304 23187 12336 23219
rect 12376 23187 12408 23219
rect 12448 23187 12480 23219
rect 12520 23187 12552 23219
rect 12592 23187 12624 23219
rect 12664 23187 12696 23219
rect 12736 23187 12768 23219
rect 12808 23187 12840 23219
rect 12880 23187 12912 23219
rect 12952 23187 12984 23219
rect 13024 23187 13056 23219
rect 13096 23187 13128 23219
rect 13168 23187 13200 23219
rect 13240 23187 13272 23219
rect 13312 23187 13344 23219
rect 13384 23187 13416 23219
rect 13456 23187 13488 23219
rect 13528 23187 13560 23219
rect 13600 23187 13632 23219
rect 13672 23187 13704 23219
rect 13744 23187 13776 23219
rect 13816 23187 13848 23219
rect 13888 23187 13920 23219
rect 13960 23187 13992 23219
rect 14032 23187 14064 23219
rect 14104 23187 14136 23219
rect 14176 23187 14208 23219
rect 14248 23187 14280 23219
rect 14320 23187 14352 23219
rect 14392 23187 14424 23219
rect 14464 23187 14496 23219
rect 14536 23187 14568 23219
rect 14608 23187 14640 23219
rect 14680 23187 14712 23219
rect 14752 23187 14784 23219
rect 14824 23187 14856 23219
rect 14896 23187 14928 23219
rect 14968 23187 15000 23219
rect 15040 23187 15072 23219
rect 15112 23187 15144 23219
rect 15184 23187 15216 23219
rect 15256 23187 15288 23219
rect 15328 23187 15360 23219
rect 15400 23187 15432 23219
rect 15472 23187 15504 23219
rect 15544 23187 15576 23219
rect 15616 23187 15648 23219
rect 15688 23187 15720 23219
rect 15760 23187 15792 23219
rect 15832 23187 15864 23219
rect 15904 23187 15936 23219
rect 18 23021 50 23053
rect 18 22952 50 22984
rect 18 22883 50 22915
rect 18 22814 50 22846
rect 18 22745 50 22777
rect 18 22676 50 22708
rect 18 22607 50 22639
rect 18 22538 50 22570
rect 18 22469 50 22501
rect 18 22400 50 22432
rect 18 22331 50 22363
rect 18 22262 50 22294
rect 18 22193 50 22225
rect 18 22124 50 22156
rect 18 22055 50 22087
rect 18 21986 50 22018
rect 18 21917 50 21949
rect 18 21848 50 21880
rect 18 21779 50 21811
rect 18 21710 50 21742
rect 18 21641 50 21673
rect 18 21572 50 21604
rect 18 21503 50 21535
rect 18 21434 50 21466
rect 18 21365 50 21397
rect 18 21296 50 21328
rect 18 21227 50 21259
rect 18 21158 50 21190
rect 18 21089 50 21121
rect 18 21020 50 21052
rect 18 20951 50 20983
rect 18 20882 50 20914
rect 18 20813 50 20845
rect 18 20744 50 20776
rect 18 20675 50 20707
rect 18 20606 50 20638
rect 18 20537 50 20569
rect 18 20468 50 20500
rect 18 20399 50 20431
rect 18 20330 50 20362
rect 18 20261 50 20293
rect 18 20192 50 20224
rect 18 20123 50 20155
rect 18 20054 50 20086
rect 18 19985 50 20017
rect 18 19916 50 19948
rect 18 19847 50 19879
rect 18 19778 50 19810
rect 18 19709 50 19741
rect 18 19640 50 19672
rect 18 19571 50 19603
rect 18 19502 50 19534
rect 18 19433 50 19465
rect 18 19364 50 19396
rect 18 19295 50 19327
rect 18 19226 50 19258
rect 18 19157 50 19189
rect 18 19088 50 19120
rect 18 19019 50 19051
rect 18 18950 50 18982
rect 18 18881 50 18913
rect 18 18812 50 18844
rect 18 18743 50 18775
rect 18 18674 50 18706
rect 18 18605 50 18637
rect 18 18536 50 18568
rect 18 18467 50 18499
rect 18 18398 50 18430
rect 18 18329 50 18361
rect 18 18260 50 18292
rect 18 18191 50 18223
rect 18 18122 50 18154
rect 18 18053 50 18085
rect 18 17984 50 18016
rect 18 17915 50 17947
rect 18 17846 50 17878
rect 18 17777 50 17809
rect 18 17708 50 17740
rect 18 17639 50 17671
rect 18 17570 50 17602
rect 18 17502 50 17534
rect 15951 23010 15983 23042
rect 15951 22942 15983 22974
rect 15951 22874 15983 22906
rect 15951 22806 15983 22838
rect 15951 22738 15983 22770
rect 15951 22670 15983 22702
rect 15951 22602 15983 22634
rect 15951 22534 15983 22566
rect 15951 22466 15983 22498
rect 15951 22398 15983 22430
rect 15951 22330 15983 22362
rect 15951 22262 15983 22294
rect 15951 22194 15983 22226
rect 15951 22126 15983 22158
rect 15951 22058 15983 22090
rect 15951 21990 15983 22022
rect 15951 21922 15983 21954
rect 15951 21854 15983 21886
rect 15951 21786 15983 21818
rect 15951 21718 15983 21750
rect 15951 21650 15983 21682
rect 15951 21582 15983 21614
rect 15951 21514 15983 21546
rect 15951 21446 15983 21478
rect 15951 21378 15983 21410
rect 15951 21310 15983 21342
rect 15951 21242 15983 21274
rect 15951 21174 15983 21206
rect 15951 21106 15983 21138
rect 15951 21038 15983 21070
rect 15951 20970 15983 21002
rect 15951 20902 15983 20934
rect 15951 20834 15983 20866
rect 15951 20766 15983 20798
rect 15951 20698 15983 20730
rect 15951 20630 15983 20662
rect 15951 20562 15983 20594
rect 15951 20494 15983 20526
rect 15951 20426 15983 20458
rect 15951 20358 15983 20390
rect 15951 20290 15983 20322
rect 15951 20222 15983 20254
rect 15951 20154 15983 20186
rect 15951 20086 15983 20118
rect 15951 20018 15983 20050
rect 15951 19950 15983 19982
rect 15951 19882 15983 19914
rect 15951 19814 15983 19846
rect 15951 19746 15983 19778
rect 15951 19678 15983 19710
rect 15951 19610 15983 19642
rect 15951 19542 15983 19574
rect 15951 19474 15983 19506
rect 15951 19406 15983 19438
rect 15951 19338 15983 19370
rect 15951 19270 15983 19302
rect 15951 19202 15983 19234
rect 15951 19134 15983 19166
rect 15951 19066 15983 19098
rect 15951 18998 15983 19030
rect 15951 18930 15983 18962
rect 15951 18862 15983 18894
rect 15951 18794 15983 18826
rect 15951 18726 15983 18758
rect 15951 18658 15983 18690
rect 15951 18590 15983 18622
rect 15951 18522 15983 18554
rect 15951 18454 15983 18486
rect 15951 18386 15983 18418
rect 15951 18318 15983 18350
rect 15951 18250 15983 18282
rect 15951 18182 15983 18214
rect 15951 18114 15983 18146
rect 15951 18046 15983 18078
rect 15951 17978 15983 18010
rect 15951 17910 15983 17942
rect 15951 17842 15983 17874
rect 15951 17774 15983 17806
rect 15951 17706 15983 17738
rect 15951 17638 15983 17670
rect 15951 17570 15983 17602
rect 15951 17502 15983 17534
rect 41 33420 657 33429
rect 41 33416 42 33420
rect 656 33416 657 33420
rect 15343 33420 15959 33429
rect 15343 33416 15344 33420
rect 15958 33416 15959 33420
rect 0 33384 42 33416
rect 656 33384 662 33416
rect 694 33384 730 33416
rect 762 33384 798 33416
rect 830 33384 866 33416
rect 898 33384 934 33416
rect 966 33384 1002 33416
rect 1034 33384 1070 33416
rect 1102 33384 1138 33416
rect 1170 33384 1206 33416
rect 1238 33384 1274 33416
rect 1306 33384 1342 33416
rect 1374 33384 1410 33416
rect 1442 33384 1478 33416
rect 1510 33384 1546 33416
rect 1578 33384 1614 33416
rect 1646 33384 1682 33416
rect 1714 33384 1750 33416
rect 1782 33384 1818 33416
rect 1850 33384 1886 33416
rect 1918 33384 1954 33416
rect 1986 33384 2022 33416
rect 2054 33384 2090 33416
rect 2122 33384 2158 33416
rect 2190 33384 2226 33416
rect 2258 33384 2294 33416
rect 2326 33384 2362 33416
rect 2394 33384 2430 33416
rect 2462 33384 2498 33416
rect 2530 33384 2566 33416
rect 2598 33384 2634 33416
rect 2666 33384 2702 33416
rect 2734 33384 2770 33416
rect 2802 33384 2838 33416
rect 2870 33384 2906 33416
rect 2938 33384 2974 33416
rect 3006 33384 3042 33416
rect 3074 33384 3110 33416
rect 3142 33384 3178 33416
rect 3210 33384 3246 33416
rect 3278 33384 3314 33416
rect 3346 33384 3382 33416
rect 3414 33384 3450 33416
rect 3482 33384 3518 33416
rect 3550 33384 3586 33416
rect 3618 33384 3654 33416
rect 3686 33384 3722 33416
rect 3754 33384 3790 33416
rect 3822 33384 3858 33416
rect 3890 33384 3926 33416
rect 3958 33384 3994 33416
rect 4026 33384 4062 33416
rect 4094 33384 4130 33416
rect 4162 33384 4198 33416
rect 4230 33384 4266 33416
rect 4298 33384 4334 33416
rect 4366 33384 4402 33416
rect 4434 33384 4470 33416
rect 4502 33384 4538 33416
rect 4570 33384 4606 33416
rect 4638 33384 4674 33416
rect 4706 33384 4742 33416
rect 4774 33384 4810 33416
rect 4842 33384 4878 33416
rect 4910 33384 4946 33416
rect 4978 33384 5014 33416
rect 5046 33384 5082 33416
rect 5114 33384 5150 33416
rect 5182 33384 5218 33416
rect 5250 33384 5286 33416
rect 5318 33384 5354 33416
rect 5386 33384 5422 33416
rect 5454 33384 5490 33416
rect 5522 33384 5558 33416
rect 5590 33384 5626 33416
rect 5658 33384 5694 33416
rect 5726 33384 5762 33416
rect 5794 33384 5830 33416
rect 5862 33384 5898 33416
rect 5930 33384 5966 33416
rect 5998 33384 6034 33416
rect 6066 33384 6102 33416
rect 6134 33384 6170 33416
rect 6202 33384 6238 33416
rect 6270 33384 6306 33416
rect 6338 33384 6374 33416
rect 6406 33384 6442 33416
rect 6474 33384 6510 33416
rect 6542 33384 6578 33416
rect 6610 33384 6646 33416
rect 6678 33384 6714 33416
rect 6746 33384 6782 33416
rect 6814 33384 6850 33416
rect 6882 33384 6918 33416
rect 6950 33384 6986 33416
rect 7018 33384 7054 33416
rect 7086 33384 7122 33416
rect 7154 33384 7190 33416
rect 7222 33384 7258 33416
rect 7290 33384 7326 33416
rect 7358 33384 7394 33416
rect 7426 33384 7462 33416
rect 7494 33384 7530 33416
rect 7562 33384 7598 33416
rect 7630 33384 7666 33416
rect 7698 33384 7734 33416
rect 7766 33384 7802 33416
rect 7834 33384 7870 33416
rect 7902 33384 7938 33416
rect 7970 33384 8006 33416
rect 8038 33384 8074 33416
rect 8106 33384 8142 33416
rect 8174 33384 8210 33416
rect 8242 33384 8278 33416
rect 8310 33384 8346 33416
rect 8378 33384 8414 33416
rect 8446 33384 8482 33416
rect 8514 33384 8550 33416
rect 8582 33384 8618 33416
rect 8650 33384 8686 33416
rect 8718 33384 8754 33416
rect 8786 33384 8822 33416
rect 8854 33384 8890 33416
rect 8922 33384 8958 33416
rect 8990 33384 9026 33416
rect 9058 33384 9094 33416
rect 9126 33384 9162 33416
rect 9194 33384 9230 33416
rect 9262 33384 9298 33416
rect 9330 33384 9366 33416
rect 9398 33384 9434 33416
rect 9466 33384 9502 33416
rect 9534 33384 9570 33416
rect 9602 33384 9638 33416
rect 9670 33384 9706 33416
rect 9738 33384 9774 33416
rect 9806 33384 9842 33416
rect 9874 33384 9910 33416
rect 9942 33384 9978 33416
rect 10010 33384 10046 33416
rect 10078 33384 10114 33416
rect 10146 33384 10182 33416
rect 10214 33384 10250 33416
rect 10282 33384 10318 33416
rect 10350 33384 10386 33416
rect 10418 33384 10454 33416
rect 10486 33384 10522 33416
rect 10554 33384 10590 33416
rect 10622 33384 10658 33416
rect 10690 33384 10726 33416
rect 10758 33384 10794 33416
rect 10826 33384 10862 33416
rect 10894 33384 10930 33416
rect 10962 33384 10998 33416
rect 11030 33384 11066 33416
rect 11098 33384 11134 33416
rect 11166 33384 11202 33416
rect 11234 33384 11270 33416
rect 11302 33384 11338 33416
rect 11370 33384 11406 33416
rect 11438 33384 11474 33416
rect 11506 33384 11542 33416
rect 11574 33384 11610 33416
rect 11642 33384 11678 33416
rect 11710 33384 11746 33416
rect 11778 33384 11814 33416
rect 11846 33384 11882 33416
rect 11914 33384 11950 33416
rect 11982 33384 12018 33416
rect 12050 33384 12086 33416
rect 12118 33384 12154 33416
rect 12186 33384 12222 33416
rect 12254 33384 12290 33416
rect 12322 33384 12358 33416
rect 12390 33384 12426 33416
rect 12458 33384 12494 33416
rect 12526 33384 12562 33416
rect 12594 33384 12630 33416
rect 12662 33384 12698 33416
rect 12730 33384 12766 33416
rect 12798 33384 12834 33416
rect 12866 33384 12902 33416
rect 12934 33384 12970 33416
rect 13002 33384 13038 33416
rect 13070 33384 13106 33416
rect 13138 33384 13174 33416
rect 13206 33384 13242 33416
rect 13274 33384 13310 33416
rect 13342 33384 13378 33416
rect 13410 33384 13446 33416
rect 13478 33384 13514 33416
rect 13546 33384 13582 33416
rect 13614 33384 13650 33416
rect 13682 33384 13718 33416
rect 13750 33384 13786 33416
rect 13818 33384 13854 33416
rect 13886 33384 13922 33416
rect 13954 33384 13990 33416
rect 14022 33384 14058 33416
rect 14090 33384 14126 33416
rect 14158 33384 14194 33416
rect 14226 33384 14262 33416
rect 14294 33384 14330 33416
rect 14362 33384 14398 33416
rect 14430 33384 14466 33416
rect 14498 33384 14534 33416
rect 14566 33384 14602 33416
rect 14634 33384 14670 33416
rect 14702 33384 14738 33416
rect 14770 33384 14806 33416
rect 14838 33384 14874 33416
rect 14906 33384 14942 33416
rect 14974 33384 15010 33416
rect 15042 33384 15078 33416
rect 15110 33384 15146 33416
rect 15178 33384 15214 33416
rect 15246 33384 15282 33416
rect 15314 33384 15344 33416
rect 15958 33384 16000 33416
rect 41 33380 42 33384
rect 656 33380 657 33384
rect 41 33371 657 33380
rect 15343 33380 15344 33384
rect 15958 33380 15959 33384
rect 15343 33371 15959 33380
rect 41 31420 657 31429
rect 41 31416 42 31420
rect 656 31416 657 31420
rect 15343 31420 15959 31429
rect 15343 31416 15344 31420
rect 15958 31416 15959 31420
rect 0 31384 42 31416
rect 656 31384 662 31416
rect 694 31384 730 31416
rect 762 31384 798 31416
rect 830 31384 866 31416
rect 898 31384 934 31416
rect 966 31384 1002 31416
rect 1034 31384 1070 31416
rect 1102 31384 1138 31416
rect 1170 31384 1206 31416
rect 1238 31384 1274 31416
rect 1306 31384 1342 31416
rect 1374 31384 1410 31416
rect 1442 31384 1478 31416
rect 1510 31384 1546 31416
rect 1578 31384 1614 31416
rect 1646 31384 1682 31416
rect 1714 31384 1750 31416
rect 1782 31384 1818 31416
rect 1850 31384 1886 31416
rect 1918 31384 1954 31416
rect 1986 31384 2022 31416
rect 2054 31384 2090 31416
rect 2122 31384 2158 31416
rect 2190 31384 2226 31416
rect 2258 31384 2294 31416
rect 2326 31384 2362 31416
rect 2394 31384 2430 31416
rect 2462 31384 2498 31416
rect 2530 31384 2566 31416
rect 2598 31384 2634 31416
rect 2666 31384 2702 31416
rect 2734 31384 2770 31416
rect 2802 31384 2838 31416
rect 2870 31384 2906 31416
rect 2938 31384 2974 31416
rect 3006 31384 3042 31416
rect 3074 31384 3110 31416
rect 3142 31384 3178 31416
rect 3210 31384 3246 31416
rect 3278 31384 3314 31416
rect 3346 31384 3382 31416
rect 3414 31384 3450 31416
rect 3482 31384 3518 31416
rect 3550 31384 3586 31416
rect 3618 31384 3654 31416
rect 3686 31384 3722 31416
rect 3754 31384 3790 31416
rect 3822 31384 3858 31416
rect 3890 31384 3926 31416
rect 3958 31384 3994 31416
rect 4026 31384 4062 31416
rect 4094 31384 4130 31416
rect 4162 31384 4198 31416
rect 4230 31384 4266 31416
rect 4298 31384 4334 31416
rect 4366 31384 4402 31416
rect 4434 31384 4470 31416
rect 4502 31384 4538 31416
rect 4570 31384 4606 31416
rect 4638 31384 4674 31416
rect 4706 31384 4742 31416
rect 4774 31384 4810 31416
rect 4842 31384 4878 31416
rect 4910 31384 4946 31416
rect 4978 31384 5014 31416
rect 5046 31384 5082 31416
rect 5114 31384 5150 31416
rect 5182 31384 5218 31416
rect 5250 31384 5286 31416
rect 5318 31384 5354 31416
rect 5386 31384 5422 31416
rect 5454 31384 5490 31416
rect 5522 31384 5558 31416
rect 5590 31384 5626 31416
rect 5658 31384 5694 31416
rect 5726 31384 5762 31416
rect 5794 31384 5830 31416
rect 5862 31384 5898 31416
rect 5930 31384 5966 31416
rect 5998 31384 6034 31416
rect 6066 31384 6102 31416
rect 6134 31384 6170 31416
rect 6202 31384 6238 31416
rect 6270 31384 6306 31416
rect 6338 31384 6374 31416
rect 6406 31384 6442 31416
rect 6474 31384 6510 31416
rect 6542 31384 6578 31416
rect 6610 31384 6646 31416
rect 6678 31384 6714 31416
rect 6746 31384 6782 31416
rect 6814 31384 6850 31416
rect 6882 31384 6918 31416
rect 6950 31384 6986 31416
rect 7018 31384 7054 31416
rect 7086 31384 7122 31416
rect 7154 31384 7190 31416
rect 7222 31384 7258 31416
rect 7290 31384 7326 31416
rect 7358 31384 7394 31416
rect 7426 31384 7462 31416
rect 7494 31384 7530 31416
rect 7562 31384 7598 31416
rect 7630 31384 7666 31416
rect 7698 31384 7734 31416
rect 7766 31384 7802 31416
rect 7834 31384 7870 31416
rect 7902 31384 7938 31416
rect 7970 31384 8006 31416
rect 8038 31384 8074 31416
rect 8106 31384 8142 31416
rect 8174 31384 8210 31416
rect 8242 31384 8278 31416
rect 8310 31384 8346 31416
rect 8378 31384 8414 31416
rect 8446 31384 8482 31416
rect 8514 31384 8550 31416
rect 8582 31384 8618 31416
rect 8650 31384 8686 31416
rect 8718 31384 8754 31416
rect 8786 31384 8822 31416
rect 8854 31384 8890 31416
rect 8922 31384 8958 31416
rect 8990 31384 9026 31416
rect 9058 31384 9094 31416
rect 9126 31384 9162 31416
rect 9194 31384 9230 31416
rect 9262 31384 9298 31416
rect 9330 31384 9366 31416
rect 9398 31384 9434 31416
rect 9466 31384 9502 31416
rect 9534 31384 9570 31416
rect 9602 31384 9638 31416
rect 9670 31384 9706 31416
rect 9738 31384 9774 31416
rect 9806 31384 9842 31416
rect 9874 31384 9910 31416
rect 9942 31384 9978 31416
rect 10010 31384 10046 31416
rect 10078 31384 10114 31416
rect 10146 31384 10182 31416
rect 10214 31384 10250 31416
rect 10282 31384 10318 31416
rect 10350 31384 10386 31416
rect 10418 31384 10454 31416
rect 10486 31384 10522 31416
rect 10554 31384 10590 31416
rect 10622 31384 10658 31416
rect 10690 31384 10726 31416
rect 10758 31384 10794 31416
rect 10826 31384 10862 31416
rect 10894 31384 10930 31416
rect 10962 31384 10998 31416
rect 11030 31384 11066 31416
rect 11098 31384 11134 31416
rect 11166 31384 11202 31416
rect 11234 31384 11270 31416
rect 11302 31384 11338 31416
rect 11370 31384 11406 31416
rect 11438 31384 11474 31416
rect 11506 31384 11542 31416
rect 11574 31384 11610 31416
rect 11642 31384 11678 31416
rect 11710 31384 11746 31416
rect 11778 31384 11814 31416
rect 11846 31384 11882 31416
rect 11914 31384 11950 31416
rect 11982 31384 12018 31416
rect 12050 31384 12086 31416
rect 12118 31384 12154 31416
rect 12186 31384 12222 31416
rect 12254 31384 12290 31416
rect 12322 31384 12358 31416
rect 12390 31384 12426 31416
rect 12458 31384 12494 31416
rect 12526 31384 12562 31416
rect 12594 31384 12630 31416
rect 12662 31384 12698 31416
rect 12730 31384 12766 31416
rect 12798 31384 12834 31416
rect 12866 31384 12902 31416
rect 12934 31384 12970 31416
rect 13002 31384 13038 31416
rect 13070 31384 13106 31416
rect 13138 31384 13174 31416
rect 13206 31384 13242 31416
rect 13274 31384 13310 31416
rect 13342 31384 13378 31416
rect 13410 31384 13446 31416
rect 13478 31384 13514 31416
rect 13546 31384 13582 31416
rect 13614 31384 13650 31416
rect 13682 31384 13718 31416
rect 13750 31384 13786 31416
rect 13818 31384 13854 31416
rect 13886 31384 13922 31416
rect 13954 31384 13990 31416
rect 14022 31384 14058 31416
rect 14090 31384 14126 31416
rect 14158 31384 14194 31416
rect 14226 31384 14262 31416
rect 14294 31384 14330 31416
rect 14362 31384 14398 31416
rect 14430 31384 14466 31416
rect 14498 31384 14534 31416
rect 14566 31384 14602 31416
rect 14634 31384 14670 31416
rect 14702 31384 14738 31416
rect 14770 31384 14806 31416
rect 14838 31384 14874 31416
rect 14906 31384 14942 31416
rect 14974 31384 15010 31416
rect 15042 31384 15078 31416
rect 15110 31384 15146 31416
rect 15178 31384 15214 31416
rect 15246 31384 15282 31416
rect 15314 31384 15344 31416
rect 15958 31384 16000 31416
rect 41 31380 42 31384
rect 656 31380 657 31384
rect 41 31371 657 31380
rect 15343 31380 15344 31384
rect 15958 31380 15959 31384
rect 15343 31371 15959 31380
rect 15835 29720 15959 29729
rect 15835 29716 15836 29720
rect 15958 29716 15959 29720
rect 0 29684 50 29716
rect 82 29684 118 29716
rect 150 29684 186 29716
rect 218 29684 254 29716
rect 286 29684 322 29716
rect 354 29684 390 29716
rect 422 29684 458 29716
rect 490 29684 526 29716
rect 558 29684 594 29716
rect 626 29684 662 29716
rect 694 29684 730 29716
rect 762 29684 798 29716
rect 830 29684 866 29716
rect 898 29684 934 29716
rect 966 29684 1002 29716
rect 1034 29684 1070 29716
rect 1102 29684 1138 29716
rect 1170 29684 1206 29716
rect 1238 29684 1274 29716
rect 1306 29684 1342 29716
rect 1374 29684 1410 29716
rect 1442 29684 1478 29716
rect 1510 29684 1546 29716
rect 1578 29684 1614 29716
rect 1646 29684 1682 29716
rect 1714 29684 1750 29716
rect 1782 29684 1818 29716
rect 1850 29684 1886 29716
rect 1918 29684 1954 29716
rect 1986 29684 2022 29716
rect 2054 29684 2090 29716
rect 2122 29684 2158 29716
rect 2190 29684 2226 29716
rect 2258 29684 2294 29716
rect 2326 29684 2362 29716
rect 2394 29684 2430 29716
rect 2462 29684 2498 29716
rect 2530 29684 2566 29716
rect 2598 29684 2634 29716
rect 2666 29684 2702 29716
rect 2734 29684 2770 29716
rect 2802 29684 2838 29716
rect 2870 29684 2906 29716
rect 2938 29684 2974 29716
rect 3006 29684 3042 29716
rect 3074 29684 3110 29716
rect 3142 29684 3178 29716
rect 3210 29684 3246 29716
rect 3278 29684 3314 29716
rect 3346 29684 3382 29716
rect 3414 29684 3450 29716
rect 3482 29684 3518 29716
rect 3550 29684 3586 29716
rect 3618 29684 3654 29716
rect 3686 29684 3722 29716
rect 3754 29684 3790 29716
rect 3822 29684 3858 29716
rect 3890 29684 3926 29716
rect 3958 29684 3994 29716
rect 4026 29684 4062 29716
rect 4094 29684 4130 29716
rect 4162 29684 4198 29716
rect 4230 29684 4266 29716
rect 4298 29684 4334 29716
rect 4366 29684 4402 29716
rect 4434 29684 4470 29716
rect 4502 29684 4538 29716
rect 4570 29684 4606 29716
rect 4638 29684 4674 29716
rect 4706 29684 4742 29716
rect 4774 29684 4810 29716
rect 4842 29684 4878 29716
rect 4910 29684 4946 29716
rect 4978 29684 5014 29716
rect 5046 29684 5082 29716
rect 5114 29684 5150 29716
rect 5182 29684 5218 29716
rect 5250 29684 5286 29716
rect 5318 29684 5354 29716
rect 5386 29684 5422 29716
rect 5454 29684 5490 29716
rect 5522 29684 5558 29716
rect 5590 29684 5626 29716
rect 5658 29684 5694 29716
rect 5726 29684 5762 29716
rect 5794 29684 5830 29716
rect 5862 29684 5898 29716
rect 5930 29684 5966 29716
rect 5998 29684 6034 29716
rect 6066 29684 6102 29716
rect 6134 29684 6170 29716
rect 6202 29684 6238 29716
rect 6270 29684 6306 29716
rect 6338 29684 6374 29716
rect 6406 29684 6442 29716
rect 6474 29684 6510 29716
rect 6542 29684 6578 29716
rect 6610 29684 6646 29716
rect 6678 29684 6714 29716
rect 6746 29684 6782 29716
rect 6814 29684 6850 29716
rect 6882 29684 6918 29716
rect 6950 29684 6986 29716
rect 7018 29684 7054 29716
rect 7086 29684 7122 29716
rect 7154 29684 7190 29716
rect 7222 29684 7258 29716
rect 7290 29684 7326 29716
rect 7358 29684 7394 29716
rect 7426 29684 7462 29716
rect 7494 29684 7530 29716
rect 7562 29684 7598 29716
rect 7630 29684 7666 29716
rect 7698 29684 7734 29716
rect 7766 29684 7802 29716
rect 7834 29684 7870 29716
rect 7902 29684 7938 29716
rect 7970 29684 8006 29716
rect 8038 29684 8074 29716
rect 8106 29684 8142 29716
rect 8174 29684 8210 29716
rect 8242 29684 8278 29716
rect 8310 29684 8346 29716
rect 8378 29684 8414 29716
rect 8446 29684 8482 29716
rect 8514 29684 8550 29716
rect 8582 29684 8618 29716
rect 8650 29684 8686 29716
rect 8718 29684 8754 29716
rect 8786 29684 8822 29716
rect 8854 29684 8890 29716
rect 8922 29684 8958 29716
rect 8990 29684 9026 29716
rect 9058 29684 9094 29716
rect 9126 29684 9162 29716
rect 9194 29684 9230 29716
rect 9262 29684 9298 29716
rect 9330 29684 9366 29716
rect 9398 29684 9434 29716
rect 9466 29684 9502 29716
rect 9534 29684 9570 29716
rect 9602 29684 9638 29716
rect 9670 29684 9706 29716
rect 9738 29684 9774 29716
rect 9806 29684 9842 29716
rect 9874 29684 9910 29716
rect 9942 29684 9978 29716
rect 10010 29684 10046 29716
rect 10078 29684 10114 29716
rect 10146 29684 10182 29716
rect 10214 29684 10250 29716
rect 10282 29684 10318 29716
rect 10350 29684 10386 29716
rect 10418 29684 10454 29716
rect 10486 29684 10522 29716
rect 10554 29684 10590 29716
rect 10622 29684 10658 29716
rect 10690 29684 10726 29716
rect 10758 29684 10794 29716
rect 10826 29684 10862 29716
rect 10894 29684 10930 29716
rect 10962 29684 10998 29716
rect 11030 29684 11066 29716
rect 11098 29684 11134 29716
rect 11166 29684 11202 29716
rect 11234 29684 11270 29716
rect 11302 29684 11338 29716
rect 11370 29684 11406 29716
rect 11438 29684 11474 29716
rect 11506 29684 11542 29716
rect 11574 29684 11610 29716
rect 11642 29684 11678 29716
rect 11710 29684 11746 29716
rect 11778 29684 11814 29716
rect 11846 29684 11882 29716
rect 11914 29684 11950 29716
rect 11982 29684 12018 29716
rect 12050 29684 12086 29716
rect 12118 29684 12154 29716
rect 12186 29684 12222 29716
rect 12254 29684 12290 29716
rect 12322 29684 12358 29716
rect 12390 29684 12426 29716
rect 12458 29684 12494 29716
rect 12526 29684 12562 29716
rect 12594 29684 12630 29716
rect 12662 29684 12698 29716
rect 12730 29684 12766 29716
rect 12798 29684 12834 29716
rect 12866 29684 12902 29716
rect 12934 29684 12970 29716
rect 13002 29684 13038 29716
rect 13070 29684 13106 29716
rect 13138 29684 13174 29716
rect 13206 29684 13242 29716
rect 13274 29684 13310 29716
rect 13342 29684 13378 29716
rect 13410 29684 13446 29716
rect 13478 29684 13514 29716
rect 13546 29684 13582 29716
rect 13614 29684 13650 29716
rect 13682 29684 13718 29716
rect 13750 29684 13786 29716
rect 13818 29684 13854 29716
rect 13886 29684 13922 29716
rect 13954 29684 13990 29716
rect 14022 29684 14058 29716
rect 14090 29684 14126 29716
rect 14158 29684 14194 29716
rect 14226 29684 14262 29716
rect 14294 29684 14330 29716
rect 14362 29684 14398 29716
rect 14430 29684 14466 29716
rect 14498 29684 14534 29716
rect 14566 29684 14602 29716
rect 14634 29684 14670 29716
rect 14702 29684 14738 29716
rect 14770 29684 14806 29716
rect 14838 29684 14874 29716
rect 14906 29684 14942 29716
rect 14974 29684 15010 29716
rect 15042 29684 15078 29716
rect 15110 29684 15146 29716
rect 15178 29684 15214 29716
rect 15246 29684 15282 29716
rect 15314 29684 15350 29716
rect 15382 29684 15442 29716
rect 15474 29684 15510 29716
rect 15542 29684 15578 29716
rect 15610 29684 15646 29716
rect 15678 29684 15714 29716
rect 15746 29684 15782 29716
rect 15814 29684 15836 29716
rect 15958 29684 16000 29716
rect 15835 29680 15836 29684
rect 15958 29680 15959 29684
rect 15835 29671 15959 29680
rect 0 27971 16000 28034
rect 0 27939 64 27971
rect 96 27939 136 27971
rect 168 27939 208 27971
rect 240 27939 280 27971
rect 312 27939 352 27971
rect 384 27939 424 27971
rect 456 27939 496 27971
rect 528 27939 568 27971
rect 600 27939 640 27971
rect 672 27939 712 27971
rect 744 27939 784 27971
rect 816 27939 856 27971
rect 888 27939 928 27971
rect 960 27939 1000 27971
rect 1032 27939 1072 27971
rect 1104 27939 1144 27971
rect 1176 27939 1216 27971
rect 1248 27939 1288 27971
rect 1320 27939 1360 27971
rect 1392 27939 1432 27971
rect 1464 27939 1504 27971
rect 1536 27939 1576 27971
rect 1608 27939 1648 27971
rect 1680 27939 1720 27971
rect 1752 27939 1792 27971
rect 1824 27939 1864 27971
rect 1896 27939 1936 27971
rect 1968 27939 2008 27971
rect 2040 27939 2080 27971
rect 2112 27939 2152 27971
rect 2184 27939 2224 27971
rect 2256 27939 2296 27971
rect 2328 27939 2368 27971
rect 2400 27939 2440 27971
rect 2472 27939 2512 27971
rect 2544 27939 2584 27971
rect 2616 27939 2656 27971
rect 2688 27939 2728 27971
rect 2760 27939 2800 27971
rect 2832 27939 2872 27971
rect 2904 27939 2944 27971
rect 2976 27939 3016 27971
rect 3048 27939 3088 27971
rect 3120 27939 3160 27971
rect 3192 27939 3232 27971
rect 3264 27939 3304 27971
rect 3336 27939 3376 27971
rect 3408 27939 3448 27971
rect 3480 27939 3520 27971
rect 3552 27939 3592 27971
rect 3624 27939 3664 27971
rect 3696 27939 3736 27971
rect 3768 27939 3808 27971
rect 3840 27939 3880 27971
rect 3912 27939 3952 27971
rect 3984 27939 4024 27971
rect 4056 27939 4096 27971
rect 4128 27939 4168 27971
rect 4200 27939 4240 27971
rect 4272 27939 4312 27971
rect 4344 27939 4384 27971
rect 4416 27939 4456 27971
rect 4488 27939 4528 27971
rect 4560 27939 4600 27971
rect 4632 27939 4672 27971
rect 4704 27939 4744 27971
rect 4776 27939 4816 27971
rect 4848 27939 4888 27971
rect 4920 27939 4960 27971
rect 4992 27939 5032 27971
rect 5064 27939 5104 27971
rect 5136 27939 5176 27971
rect 5208 27939 5248 27971
rect 5280 27939 5320 27971
rect 5352 27939 5392 27971
rect 5424 27939 5464 27971
rect 5496 27939 5536 27971
rect 5568 27939 5608 27971
rect 5640 27939 5680 27971
rect 5712 27939 5752 27971
rect 5784 27939 5824 27971
rect 5856 27939 5896 27971
rect 5928 27939 5968 27971
rect 6000 27939 6040 27971
rect 6072 27939 6112 27971
rect 6144 27939 6184 27971
rect 6216 27939 6256 27971
rect 6288 27939 6328 27971
rect 6360 27939 6400 27971
rect 6432 27939 6472 27971
rect 6504 27939 6544 27971
rect 6576 27939 6616 27971
rect 6648 27939 6688 27971
rect 6720 27939 6760 27971
rect 6792 27939 6832 27971
rect 6864 27939 6904 27971
rect 6936 27939 6976 27971
rect 7008 27939 7048 27971
rect 7080 27939 7120 27971
rect 7152 27939 7192 27971
rect 7224 27939 7264 27971
rect 7296 27939 7336 27971
rect 7368 27939 7408 27971
rect 7440 27939 7480 27971
rect 7512 27939 7552 27971
rect 7584 27939 7624 27971
rect 7656 27939 7696 27971
rect 7728 27939 7768 27971
rect 7800 27939 7840 27971
rect 7872 27939 7912 27971
rect 7944 27939 7984 27971
rect 8016 27939 8056 27971
rect 8088 27939 8128 27971
rect 8160 27939 8200 27971
rect 8232 27939 8272 27971
rect 8304 27939 8344 27971
rect 8376 27939 8416 27971
rect 8448 27939 8488 27971
rect 8520 27939 8560 27971
rect 8592 27939 8632 27971
rect 8664 27939 8704 27971
rect 8736 27939 8776 27971
rect 8808 27939 8848 27971
rect 8880 27939 8920 27971
rect 8952 27939 8992 27971
rect 9024 27939 9064 27971
rect 9096 27939 9136 27971
rect 9168 27939 9208 27971
rect 9240 27939 9280 27971
rect 9312 27939 9352 27971
rect 9384 27939 9424 27971
rect 9456 27939 9496 27971
rect 9528 27939 9568 27971
rect 9600 27939 9640 27971
rect 9672 27939 9712 27971
rect 9744 27939 9784 27971
rect 9816 27939 9856 27971
rect 9888 27939 9928 27971
rect 9960 27939 10000 27971
rect 10032 27939 10072 27971
rect 10104 27939 10144 27971
rect 10176 27939 10216 27971
rect 10248 27939 10288 27971
rect 10320 27939 10360 27971
rect 10392 27939 10432 27971
rect 10464 27939 10504 27971
rect 10536 27939 10576 27971
rect 10608 27939 10648 27971
rect 10680 27939 10720 27971
rect 10752 27939 10792 27971
rect 10824 27939 10864 27971
rect 10896 27939 10936 27971
rect 10968 27939 11008 27971
rect 11040 27939 11080 27971
rect 11112 27939 11152 27971
rect 11184 27939 11224 27971
rect 11256 27939 11296 27971
rect 11328 27939 11368 27971
rect 11400 27939 11440 27971
rect 11472 27939 11512 27971
rect 11544 27939 11584 27971
rect 11616 27939 11656 27971
rect 11688 27939 11728 27971
rect 11760 27939 11800 27971
rect 11832 27939 11872 27971
rect 11904 27939 11944 27971
rect 11976 27939 12016 27971
rect 12048 27939 12088 27971
rect 12120 27939 12160 27971
rect 12192 27939 12232 27971
rect 12264 27939 12304 27971
rect 12336 27939 12376 27971
rect 12408 27939 12448 27971
rect 12480 27939 12520 27971
rect 12552 27939 12592 27971
rect 12624 27939 12664 27971
rect 12696 27939 12736 27971
rect 12768 27939 12808 27971
rect 12840 27939 12880 27971
rect 12912 27939 12952 27971
rect 12984 27939 13024 27971
rect 13056 27939 13096 27971
rect 13128 27939 13168 27971
rect 13200 27939 13240 27971
rect 13272 27939 13312 27971
rect 13344 27939 13384 27971
rect 13416 27939 13456 27971
rect 13488 27939 13528 27971
rect 13560 27939 13600 27971
rect 13632 27939 13672 27971
rect 13704 27939 13744 27971
rect 13776 27939 13816 27971
rect 13848 27939 13888 27971
rect 13920 27939 13960 27971
rect 13992 27939 14032 27971
rect 14064 27939 14104 27971
rect 14136 27939 14176 27971
rect 14208 27939 14248 27971
rect 14280 27939 14320 27971
rect 14352 27939 14392 27971
rect 14424 27939 14464 27971
rect 14496 27939 14536 27971
rect 14568 27939 14608 27971
rect 14640 27939 14680 27971
rect 14712 27939 14752 27971
rect 14784 27939 14824 27971
rect 14856 27939 14896 27971
rect 14928 27939 14968 27971
rect 15000 27939 15040 27971
rect 15072 27939 15112 27971
rect 15144 27939 15184 27971
rect 15216 27939 15256 27971
rect 15288 27939 15328 27971
rect 15360 27939 15400 27971
rect 15432 27939 15472 27971
rect 15504 27939 15544 27971
rect 15576 27939 15616 27971
rect 15648 27939 15688 27971
rect 15720 27939 15760 27971
rect 15792 27939 15832 27971
rect 15864 27939 15904 27971
rect 15936 27939 16000 27971
rect 0 27899 16000 27939
rect 0 27867 64 27899
rect 96 27867 136 27899
rect 168 27867 208 27899
rect 240 27867 280 27899
rect 312 27867 352 27899
rect 384 27867 424 27899
rect 456 27867 496 27899
rect 528 27867 568 27899
rect 600 27867 640 27899
rect 672 27867 712 27899
rect 744 27867 784 27899
rect 816 27867 856 27899
rect 888 27867 928 27899
rect 960 27867 1000 27899
rect 1032 27867 1072 27899
rect 1104 27867 1144 27899
rect 1176 27867 1216 27899
rect 1248 27867 1288 27899
rect 1320 27867 1360 27899
rect 1392 27867 1432 27899
rect 1464 27867 1504 27899
rect 1536 27867 1576 27899
rect 1608 27867 1648 27899
rect 1680 27867 1720 27899
rect 1752 27867 1792 27899
rect 1824 27867 1864 27899
rect 1896 27867 1936 27899
rect 1968 27867 2008 27899
rect 2040 27867 2080 27899
rect 2112 27867 2152 27899
rect 2184 27867 2224 27899
rect 2256 27867 2296 27899
rect 2328 27867 2368 27899
rect 2400 27867 2440 27899
rect 2472 27867 2512 27899
rect 2544 27867 2584 27899
rect 2616 27867 2656 27899
rect 2688 27867 2728 27899
rect 2760 27867 2800 27899
rect 2832 27867 2872 27899
rect 2904 27867 2944 27899
rect 2976 27867 3016 27899
rect 3048 27867 3088 27899
rect 3120 27867 3160 27899
rect 3192 27867 3232 27899
rect 3264 27867 3304 27899
rect 3336 27867 3376 27899
rect 3408 27867 3448 27899
rect 3480 27867 3520 27899
rect 3552 27867 3592 27899
rect 3624 27867 3664 27899
rect 3696 27867 3736 27899
rect 3768 27867 3808 27899
rect 3840 27867 3880 27899
rect 3912 27867 3952 27899
rect 3984 27867 4024 27899
rect 4056 27867 4096 27899
rect 4128 27867 4168 27899
rect 4200 27867 4240 27899
rect 4272 27867 4312 27899
rect 4344 27867 4384 27899
rect 4416 27867 4456 27899
rect 4488 27867 4528 27899
rect 4560 27867 4600 27899
rect 4632 27867 4672 27899
rect 4704 27867 4744 27899
rect 4776 27867 4816 27899
rect 4848 27867 4888 27899
rect 4920 27867 4960 27899
rect 4992 27867 5032 27899
rect 5064 27867 5104 27899
rect 5136 27867 5176 27899
rect 5208 27867 5248 27899
rect 5280 27867 5320 27899
rect 5352 27867 5392 27899
rect 5424 27867 5464 27899
rect 5496 27867 5536 27899
rect 5568 27867 5608 27899
rect 5640 27867 5680 27899
rect 5712 27867 5752 27899
rect 5784 27867 5824 27899
rect 5856 27867 5896 27899
rect 5928 27867 5968 27899
rect 6000 27867 6040 27899
rect 6072 27867 6112 27899
rect 6144 27867 6184 27899
rect 6216 27867 6256 27899
rect 6288 27867 6328 27899
rect 6360 27867 6400 27899
rect 6432 27867 6472 27899
rect 6504 27867 6544 27899
rect 6576 27867 6616 27899
rect 6648 27867 6688 27899
rect 6720 27867 6760 27899
rect 6792 27867 6832 27899
rect 6864 27867 6904 27899
rect 6936 27867 6976 27899
rect 7008 27867 7048 27899
rect 7080 27867 7120 27899
rect 7152 27867 7192 27899
rect 7224 27867 7264 27899
rect 7296 27867 7336 27899
rect 7368 27867 7408 27899
rect 7440 27867 7480 27899
rect 7512 27867 7552 27899
rect 7584 27867 7624 27899
rect 7656 27867 7696 27899
rect 7728 27867 7768 27899
rect 7800 27867 7840 27899
rect 7872 27867 7912 27899
rect 7944 27867 7984 27899
rect 8016 27867 8056 27899
rect 8088 27867 8128 27899
rect 8160 27867 8200 27899
rect 8232 27867 8272 27899
rect 8304 27867 8344 27899
rect 8376 27867 8416 27899
rect 8448 27867 8488 27899
rect 8520 27867 8560 27899
rect 8592 27867 8632 27899
rect 8664 27867 8704 27899
rect 8736 27867 8776 27899
rect 8808 27867 8848 27899
rect 8880 27867 8920 27899
rect 8952 27867 8992 27899
rect 9024 27867 9064 27899
rect 9096 27867 9136 27899
rect 9168 27867 9208 27899
rect 9240 27867 9280 27899
rect 9312 27867 9352 27899
rect 9384 27867 9424 27899
rect 9456 27867 9496 27899
rect 9528 27867 9568 27899
rect 9600 27867 9640 27899
rect 9672 27867 9712 27899
rect 9744 27867 9784 27899
rect 9816 27867 9856 27899
rect 9888 27867 9928 27899
rect 9960 27867 10000 27899
rect 10032 27867 10072 27899
rect 10104 27867 10144 27899
rect 10176 27867 10216 27899
rect 10248 27867 10288 27899
rect 10320 27867 10360 27899
rect 10392 27867 10432 27899
rect 10464 27867 10504 27899
rect 10536 27867 10576 27899
rect 10608 27867 10648 27899
rect 10680 27867 10720 27899
rect 10752 27867 10792 27899
rect 10824 27867 10864 27899
rect 10896 27867 10936 27899
rect 10968 27867 11008 27899
rect 11040 27867 11080 27899
rect 11112 27867 11152 27899
rect 11184 27867 11224 27899
rect 11256 27867 11296 27899
rect 11328 27867 11368 27899
rect 11400 27867 11440 27899
rect 11472 27867 11512 27899
rect 11544 27867 11584 27899
rect 11616 27867 11656 27899
rect 11688 27867 11728 27899
rect 11760 27867 11800 27899
rect 11832 27867 11872 27899
rect 11904 27867 11944 27899
rect 11976 27867 12016 27899
rect 12048 27867 12088 27899
rect 12120 27867 12160 27899
rect 12192 27867 12232 27899
rect 12264 27867 12304 27899
rect 12336 27867 12376 27899
rect 12408 27867 12448 27899
rect 12480 27867 12520 27899
rect 12552 27867 12592 27899
rect 12624 27867 12664 27899
rect 12696 27867 12736 27899
rect 12768 27867 12808 27899
rect 12840 27867 12880 27899
rect 12912 27867 12952 27899
rect 12984 27867 13024 27899
rect 13056 27867 13096 27899
rect 13128 27867 13168 27899
rect 13200 27867 13240 27899
rect 13272 27867 13312 27899
rect 13344 27867 13384 27899
rect 13416 27867 13456 27899
rect 13488 27867 13528 27899
rect 13560 27867 13600 27899
rect 13632 27867 13672 27899
rect 13704 27867 13744 27899
rect 13776 27867 13816 27899
rect 13848 27867 13888 27899
rect 13920 27867 13960 27899
rect 13992 27867 14032 27899
rect 14064 27867 14104 27899
rect 14136 27867 14176 27899
rect 14208 27867 14248 27899
rect 14280 27867 14320 27899
rect 14352 27867 14392 27899
rect 14424 27867 14464 27899
rect 14496 27867 14536 27899
rect 14568 27867 14608 27899
rect 14640 27867 14680 27899
rect 14712 27867 14752 27899
rect 14784 27867 14824 27899
rect 14856 27867 14896 27899
rect 14928 27867 14968 27899
rect 15000 27867 15040 27899
rect 15072 27867 15112 27899
rect 15144 27867 15184 27899
rect 15216 27867 15256 27899
rect 15288 27867 15328 27899
rect 15360 27867 15400 27899
rect 15432 27867 15472 27899
rect 15504 27867 15544 27899
rect 15576 27867 15616 27899
rect 15648 27867 15688 27899
rect 15720 27867 15760 27899
rect 15792 27867 15832 27899
rect 15864 27867 15904 27899
rect 15936 27867 16000 27899
rect 0 27827 16000 27867
rect 0 27795 64 27827
rect 96 27795 136 27827
rect 168 27795 208 27827
rect 240 27795 280 27827
rect 312 27795 352 27827
rect 384 27795 424 27827
rect 456 27795 496 27827
rect 528 27795 568 27827
rect 600 27795 640 27827
rect 672 27795 712 27827
rect 744 27795 784 27827
rect 816 27795 856 27827
rect 888 27795 928 27827
rect 960 27795 1000 27827
rect 1032 27795 1072 27827
rect 1104 27795 1144 27827
rect 1176 27795 1216 27827
rect 1248 27795 1288 27827
rect 1320 27795 1360 27827
rect 1392 27795 1432 27827
rect 1464 27795 1504 27827
rect 1536 27795 1576 27827
rect 1608 27795 1648 27827
rect 1680 27795 1720 27827
rect 1752 27795 1792 27827
rect 1824 27795 1864 27827
rect 1896 27795 1936 27827
rect 1968 27795 2008 27827
rect 2040 27795 2080 27827
rect 2112 27795 2152 27827
rect 2184 27795 2224 27827
rect 2256 27795 2296 27827
rect 2328 27795 2368 27827
rect 2400 27795 2440 27827
rect 2472 27795 2512 27827
rect 2544 27795 2584 27827
rect 2616 27795 2656 27827
rect 2688 27795 2728 27827
rect 2760 27795 2800 27827
rect 2832 27795 2872 27827
rect 2904 27795 2944 27827
rect 2976 27795 3016 27827
rect 3048 27795 3088 27827
rect 3120 27795 3160 27827
rect 3192 27795 3232 27827
rect 3264 27795 3304 27827
rect 3336 27795 3376 27827
rect 3408 27795 3448 27827
rect 3480 27795 3520 27827
rect 3552 27795 3592 27827
rect 3624 27795 3664 27827
rect 3696 27795 3736 27827
rect 3768 27795 3808 27827
rect 3840 27795 3880 27827
rect 3912 27795 3952 27827
rect 3984 27795 4024 27827
rect 4056 27795 4096 27827
rect 4128 27795 4168 27827
rect 4200 27795 4240 27827
rect 4272 27795 4312 27827
rect 4344 27795 4384 27827
rect 4416 27795 4456 27827
rect 4488 27795 4528 27827
rect 4560 27795 4600 27827
rect 4632 27795 4672 27827
rect 4704 27795 4744 27827
rect 4776 27795 4816 27827
rect 4848 27795 4888 27827
rect 4920 27795 4960 27827
rect 4992 27795 5032 27827
rect 5064 27795 5104 27827
rect 5136 27795 5176 27827
rect 5208 27795 5248 27827
rect 5280 27795 5320 27827
rect 5352 27795 5392 27827
rect 5424 27795 5464 27827
rect 5496 27795 5536 27827
rect 5568 27795 5608 27827
rect 5640 27795 5680 27827
rect 5712 27795 5752 27827
rect 5784 27795 5824 27827
rect 5856 27795 5896 27827
rect 5928 27795 5968 27827
rect 6000 27795 6040 27827
rect 6072 27795 6112 27827
rect 6144 27795 6184 27827
rect 6216 27795 6256 27827
rect 6288 27795 6328 27827
rect 6360 27795 6400 27827
rect 6432 27795 6472 27827
rect 6504 27795 6544 27827
rect 6576 27795 6616 27827
rect 6648 27795 6688 27827
rect 6720 27795 6760 27827
rect 6792 27795 6832 27827
rect 6864 27795 6904 27827
rect 6936 27795 6976 27827
rect 7008 27795 7048 27827
rect 7080 27795 7120 27827
rect 7152 27795 7192 27827
rect 7224 27795 7264 27827
rect 7296 27795 7336 27827
rect 7368 27795 7408 27827
rect 7440 27795 7480 27827
rect 7512 27795 7552 27827
rect 7584 27795 7624 27827
rect 7656 27795 7696 27827
rect 7728 27795 7768 27827
rect 7800 27795 7840 27827
rect 7872 27795 7912 27827
rect 7944 27795 7984 27827
rect 8016 27795 8056 27827
rect 8088 27795 8128 27827
rect 8160 27795 8200 27827
rect 8232 27795 8272 27827
rect 8304 27795 8344 27827
rect 8376 27795 8416 27827
rect 8448 27795 8488 27827
rect 8520 27795 8560 27827
rect 8592 27795 8632 27827
rect 8664 27795 8704 27827
rect 8736 27795 8776 27827
rect 8808 27795 8848 27827
rect 8880 27795 8920 27827
rect 8952 27795 8992 27827
rect 9024 27795 9064 27827
rect 9096 27795 9136 27827
rect 9168 27795 9208 27827
rect 9240 27795 9280 27827
rect 9312 27795 9352 27827
rect 9384 27795 9424 27827
rect 9456 27795 9496 27827
rect 9528 27795 9568 27827
rect 9600 27795 9640 27827
rect 9672 27795 9712 27827
rect 9744 27795 9784 27827
rect 9816 27795 9856 27827
rect 9888 27795 9928 27827
rect 9960 27795 10000 27827
rect 10032 27795 10072 27827
rect 10104 27795 10144 27827
rect 10176 27795 10216 27827
rect 10248 27795 10288 27827
rect 10320 27795 10360 27827
rect 10392 27795 10432 27827
rect 10464 27795 10504 27827
rect 10536 27795 10576 27827
rect 10608 27795 10648 27827
rect 10680 27795 10720 27827
rect 10752 27795 10792 27827
rect 10824 27795 10864 27827
rect 10896 27795 10936 27827
rect 10968 27795 11008 27827
rect 11040 27795 11080 27827
rect 11112 27795 11152 27827
rect 11184 27795 11224 27827
rect 11256 27795 11296 27827
rect 11328 27795 11368 27827
rect 11400 27795 11440 27827
rect 11472 27795 11512 27827
rect 11544 27795 11584 27827
rect 11616 27795 11656 27827
rect 11688 27795 11728 27827
rect 11760 27795 11800 27827
rect 11832 27795 11872 27827
rect 11904 27795 11944 27827
rect 11976 27795 12016 27827
rect 12048 27795 12088 27827
rect 12120 27795 12160 27827
rect 12192 27795 12232 27827
rect 12264 27795 12304 27827
rect 12336 27795 12376 27827
rect 12408 27795 12448 27827
rect 12480 27795 12520 27827
rect 12552 27795 12592 27827
rect 12624 27795 12664 27827
rect 12696 27795 12736 27827
rect 12768 27795 12808 27827
rect 12840 27795 12880 27827
rect 12912 27795 12952 27827
rect 12984 27795 13024 27827
rect 13056 27795 13096 27827
rect 13128 27795 13168 27827
rect 13200 27795 13240 27827
rect 13272 27795 13312 27827
rect 13344 27795 13384 27827
rect 13416 27795 13456 27827
rect 13488 27795 13528 27827
rect 13560 27795 13600 27827
rect 13632 27795 13672 27827
rect 13704 27795 13744 27827
rect 13776 27795 13816 27827
rect 13848 27795 13888 27827
rect 13920 27795 13960 27827
rect 13992 27795 14032 27827
rect 14064 27795 14104 27827
rect 14136 27795 14176 27827
rect 14208 27795 14248 27827
rect 14280 27795 14320 27827
rect 14352 27795 14392 27827
rect 14424 27795 14464 27827
rect 14496 27795 14536 27827
rect 14568 27795 14608 27827
rect 14640 27795 14680 27827
rect 14712 27795 14752 27827
rect 14784 27795 14824 27827
rect 14856 27795 14896 27827
rect 14928 27795 14968 27827
rect 15000 27795 15040 27827
rect 15072 27795 15112 27827
rect 15144 27795 15184 27827
rect 15216 27795 15256 27827
rect 15288 27795 15328 27827
rect 15360 27795 15400 27827
rect 15432 27795 15472 27827
rect 15504 27795 15544 27827
rect 15576 27795 15616 27827
rect 15648 27795 15688 27827
rect 15720 27795 15760 27827
rect 15792 27795 15832 27827
rect 15864 27795 15904 27827
rect 15936 27795 16000 27827
rect 0 27755 16000 27795
rect 0 27723 64 27755
rect 96 27723 136 27755
rect 168 27723 208 27755
rect 240 27723 280 27755
rect 312 27723 352 27755
rect 384 27723 424 27755
rect 456 27723 496 27755
rect 528 27723 568 27755
rect 600 27723 640 27755
rect 672 27723 712 27755
rect 744 27723 784 27755
rect 816 27723 856 27755
rect 888 27723 928 27755
rect 960 27723 1000 27755
rect 1032 27723 1072 27755
rect 1104 27723 1144 27755
rect 1176 27723 1216 27755
rect 1248 27723 1288 27755
rect 1320 27723 1360 27755
rect 1392 27723 1432 27755
rect 1464 27723 1504 27755
rect 1536 27723 1576 27755
rect 1608 27723 1648 27755
rect 1680 27723 1720 27755
rect 1752 27723 1792 27755
rect 1824 27723 1864 27755
rect 1896 27723 1936 27755
rect 1968 27723 2008 27755
rect 2040 27723 2080 27755
rect 2112 27723 2152 27755
rect 2184 27723 2224 27755
rect 2256 27723 2296 27755
rect 2328 27723 2368 27755
rect 2400 27723 2440 27755
rect 2472 27723 2512 27755
rect 2544 27723 2584 27755
rect 2616 27723 2656 27755
rect 2688 27723 2728 27755
rect 2760 27723 2800 27755
rect 2832 27723 2872 27755
rect 2904 27723 2944 27755
rect 2976 27723 3016 27755
rect 3048 27723 3088 27755
rect 3120 27723 3160 27755
rect 3192 27723 3232 27755
rect 3264 27723 3304 27755
rect 3336 27723 3376 27755
rect 3408 27723 3448 27755
rect 3480 27723 3520 27755
rect 3552 27723 3592 27755
rect 3624 27723 3664 27755
rect 3696 27723 3736 27755
rect 3768 27723 3808 27755
rect 3840 27723 3880 27755
rect 3912 27723 3952 27755
rect 3984 27723 4024 27755
rect 4056 27723 4096 27755
rect 4128 27723 4168 27755
rect 4200 27723 4240 27755
rect 4272 27723 4312 27755
rect 4344 27723 4384 27755
rect 4416 27723 4456 27755
rect 4488 27723 4528 27755
rect 4560 27723 4600 27755
rect 4632 27723 4672 27755
rect 4704 27723 4744 27755
rect 4776 27723 4816 27755
rect 4848 27723 4888 27755
rect 4920 27723 4960 27755
rect 4992 27723 5032 27755
rect 5064 27723 5104 27755
rect 5136 27723 5176 27755
rect 5208 27723 5248 27755
rect 5280 27723 5320 27755
rect 5352 27723 5392 27755
rect 5424 27723 5464 27755
rect 5496 27723 5536 27755
rect 5568 27723 5608 27755
rect 5640 27723 5680 27755
rect 5712 27723 5752 27755
rect 5784 27723 5824 27755
rect 5856 27723 5896 27755
rect 5928 27723 5968 27755
rect 6000 27723 6040 27755
rect 6072 27723 6112 27755
rect 6144 27723 6184 27755
rect 6216 27723 6256 27755
rect 6288 27723 6328 27755
rect 6360 27723 6400 27755
rect 6432 27723 6472 27755
rect 6504 27723 6544 27755
rect 6576 27723 6616 27755
rect 6648 27723 6688 27755
rect 6720 27723 6760 27755
rect 6792 27723 6832 27755
rect 6864 27723 6904 27755
rect 6936 27723 6976 27755
rect 7008 27723 7048 27755
rect 7080 27723 7120 27755
rect 7152 27723 7192 27755
rect 7224 27723 7264 27755
rect 7296 27723 7336 27755
rect 7368 27723 7408 27755
rect 7440 27723 7480 27755
rect 7512 27723 7552 27755
rect 7584 27723 7624 27755
rect 7656 27723 7696 27755
rect 7728 27723 7768 27755
rect 7800 27723 7840 27755
rect 7872 27723 7912 27755
rect 7944 27723 7984 27755
rect 8016 27723 8056 27755
rect 8088 27723 8128 27755
rect 8160 27723 8200 27755
rect 8232 27723 8272 27755
rect 8304 27723 8344 27755
rect 8376 27723 8416 27755
rect 8448 27723 8488 27755
rect 8520 27723 8560 27755
rect 8592 27723 8632 27755
rect 8664 27723 8704 27755
rect 8736 27723 8776 27755
rect 8808 27723 8848 27755
rect 8880 27723 8920 27755
rect 8952 27723 8992 27755
rect 9024 27723 9064 27755
rect 9096 27723 9136 27755
rect 9168 27723 9208 27755
rect 9240 27723 9280 27755
rect 9312 27723 9352 27755
rect 9384 27723 9424 27755
rect 9456 27723 9496 27755
rect 9528 27723 9568 27755
rect 9600 27723 9640 27755
rect 9672 27723 9712 27755
rect 9744 27723 9784 27755
rect 9816 27723 9856 27755
rect 9888 27723 9928 27755
rect 9960 27723 10000 27755
rect 10032 27723 10072 27755
rect 10104 27723 10144 27755
rect 10176 27723 10216 27755
rect 10248 27723 10288 27755
rect 10320 27723 10360 27755
rect 10392 27723 10432 27755
rect 10464 27723 10504 27755
rect 10536 27723 10576 27755
rect 10608 27723 10648 27755
rect 10680 27723 10720 27755
rect 10752 27723 10792 27755
rect 10824 27723 10864 27755
rect 10896 27723 10936 27755
rect 10968 27723 11008 27755
rect 11040 27723 11080 27755
rect 11112 27723 11152 27755
rect 11184 27723 11224 27755
rect 11256 27723 11296 27755
rect 11328 27723 11368 27755
rect 11400 27723 11440 27755
rect 11472 27723 11512 27755
rect 11544 27723 11584 27755
rect 11616 27723 11656 27755
rect 11688 27723 11728 27755
rect 11760 27723 11800 27755
rect 11832 27723 11872 27755
rect 11904 27723 11944 27755
rect 11976 27723 12016 27755
rect 12048 27723 12088 27755
rect 12120 27723 12160 27755
rect 12192 27723 12232 27755
rect 12264 27723 12304 27755
rect 12336 27723 12376 27755
rect 12408 27723 12448 27755
rect 12480 27723 12520 27755
rect 12552 27723 12592 27755
rect 12624 27723 12664 27755
rect 12696 27723 12736 27755
rect 12768 27723 12808 27755
rect 12840 27723 12880 27755
rect 12912 27723 12952 27755
rect 12984 27723 13024 27755
rect 13056 27723 13096 27755
rect 13128 27723 13168 27755
rect 13200 27723 13240 27755
rect 13272 27723 13312 27755
rect 13344 27723 13384 27755
rect 13416 27723 13456 27755
rect 13488 27723 13528 27755
rect 13560 27723 13600 27755
rect 13632 27723 13672 27755
rect 13704 27723 13744 27755
rect 13776 27723 13816 27755
rect 13848 27723 13888 27755
rect 13920 27723 13960 27755
rect 13992 27723 14032 27755
rect 14064 27723 14104 27755
rect 14136 27723 14176 27755
rect 14208 27723 14248 27755
rect 14280 27723 14320 27755
rect 14352 27723 14392 27755
rect 14424 27723 14464 27755
rect 14496 27723 14536 27755
rect 14568 27723 14608 27755
rect 14640 27723 14680 27755
rect 14712 27723 14752 27755
rect 14784 27723 14824 27755
rect 14856 27723 14896 27755
rect 14928 27723 14968 27755
rect 15000 27723 15040 27755
rect 15072 27723 15112 27755
rect 15144 27723 15184 27755
rect 15216 27723 15256 27755
rect 15288 27723 15328 27755
rect 15360 27723 15400 27755
rect 15432 27723 15472 27755
rect 15504 27723 15544 27755
rect 15576 27723 15616 27755
rect 15648 27723 15688 27755
rect 15720 27723 15760 27755
rect 15792 27723 15832 27755
rect 15864 27723 15904 27755
rect 15936 27723 16000 27755
rect 0 27683 16000 27723
rect 0 27651 64 27683
rect 96 27651 136 27683
rect 168 27651 208 27683
rect 240 27651 280 27683
rect 312 27651 352 27683
rect 384 27651 424 27683
rect 456 27651 496 27683
rect 528 27651 568 27683
rect 600 27651 640 27683
rect 672 27651 712 27683
rect 744 27651 784 27683
rect 816 27651 856 27683
rect 888 27651 928 27683
rect 960 27651 1000 27683
rect 1032 27651 1072 27683
rect 1104 27651 1144 27683
rect 1176 27651 1216 27683
rect 1248 27651 1288 27683
rect 1320 27651 1360 27683
rect 1392 27651 1432 27683
rect 1464 27651 1504 27683
rect 1536 27651 1576 27683
rect 1608 27651 1648 27683
rect 1680 27651 1720 27683
rect 1752 27651 1792 27683
rect 1824 27651 1864 27683
rect 1896 27651 1936 27683
rect 1968 27651 2008 27683
rect 2040 27651 2080 27683
rect 2112 27651 2152 27683
rect 2184 27651 2224 27683
rect 2256 27651 2296 27683
rect 2328 27651 2368 27683
rect 2400 27651 2440 27683
rect 2472 27651 2512 27683
rect 2544 27651 2584 27683
rect 2616 27651 2656 27683
rect 2688 27651 2728 27683
rect 2760 27651 2800 27683
rect 2832 27651 2872 27683
rect 2904 27651 2944 27683
rect 2976 27651 3016 27683
rect 3048 27651 3088 27683
rect 3120 27651 3160 27683
rect 3192 27651 3232 27683
rect 3264 27651 3304 27683
rect 3336 27651 3376 27683
rect 3408 27651 3448 27683
rect 3480 27651 3520 27683
rect 3552 27651 3592 27683
rect 3624 27651 3664 27683
rect 3696 27651 3736 27683
rect 3768 27651 3808 27683
rect 3840 27651 3880 27683
rect 3912 27651 3952 27683
rect 3984 27651 4024 27683
rect 4056 27651 4096 27683
rect 4128 27651 4168 27683
rect 4200 27651 4240 27683
rect 4272 27651 4312 27683
rect 4344 27651 4384 27683
rect 4416 27651 4456 27683
rect 4488 27651 4528 27683
rect 4560 27651 4600 27683
rect 4632 27651 4672 27683
rect 4704 27651 4744 27683
rect 4776 27651 4816 27683
rect 4848 27651 4888 27683
rect 4920 27651 4960 27683
rect 4992 27651 5032 27683
rect 5064 27651 5104 27683
rect 5136 27651 5176 27683
rect 5208 27651 5248 27683
rect 5280 27651 5320 27683
rect 5352 27651 5392 27683
rect 5424 27651 5464 27683
rect 5496 27651 5536 27683
rect 5568 27651 5608 27683
rect 5640 27651 5680 27683
rect 5712 27651 5752 27683
rect 5784 27651 5824 27683
rect 5856 27651 5896 27683
rect 5928 27651 5968 27683
rect 6000 27651 6040 27683
rect 6072 27651 6112 27683
rect 6144 27651 6184 27683
rect 6216 27651 6256 27683
rect 6288 27651 6328 27683
rect 6360 27651 6400 27683
rect 6432 27651 6472 27683
rect 6504 27651 6544 27683
rect 6576 27651 6616 27683
rect 6648 27651 6688 27683
rect 6720 27651 6760 27683
rect 6792 27651 6832 27683
rect 6864 27651 6904 27683
rect 6936 27651 6976 27683
rect 7008 27651 7048 27683
rect 7080 27651 7120 27683
rect 7152 27651 7192 27683
rect 7224 27651 7264 27683
rect 7296 27651 7336 27683
rect 7368 27651 7408 27683
rect 7440 27651 7480 27683
rect 7512 27651 7552 27683
rect 7584 27651 7624 27683
rect 7656 27651 7696 27683
rect 7728 27651 7768 27683
rect 7800 27651 7840 27683
rect 7872 27651 7912 27683
rect 7944 27651 7984 27683
rect 8016 27651 8056 27683
rect 8088 27651 8128 27683
rect 8160 27651 8200 27683
rect 8232 27651 8272 27683
rect 8304 27651 8344 27683
rect 8376 27651 8416 27683
rect 8448 27651 8488 27683
rect 8520 27651 8560 27683
rect 8592 27651 8632 27683
rect 8664 27651 8704 27683
rect 8736 27651 8776 27683
rect 8808 27651 8848 27683
rect 8880 27651 8920 27683
rect 8952 27651 8992 27683
rect 9024 27651 9064 27683
rect 9096 27651 9136 27683
rect 9168 27651 9208 27683
rect 9240 27651 9280 27683
rect 9312 27651 9352 27683
rect 9384 27651 9424 27683
rect 9456 27651 9496 27683
rect 9528 27651 9568 27683
rect 9600 27651 9640 27683
rect 9672 27651 9712 27683
rect 9744 27651 9784 27683
rect 9816 27651 9856 27683
rect 9888 27651 9928 27683
rect 9960 27651 10000 27683
rect 10032 27651 10072 27683
rect 10104 27651 10144 27683
rect 10176 27651 10216 27683
rect 10248 27651 10288 27683
rect 10320 27651 10360 27683
rect 10392 27651 10432 27683
rect 10464 27651 10504 27683
rect 10536 27651 10576 27683
rect 10608 27651 10648 27683
rect 10680 27651 10720 27683
rect 10752 27651 10792 27683
rect 10824 27651 10864 27683
rect 10896 27651 10936 27683
rect 10968 27651 11008 27683
rect 11040 27651 11080 27683
rect 11112 27651 11152 27683
rect 11184 27651 11224 27683
rect 11256 27651 11296 27683
rect 11328 27651 11368 27683
rect 11400 27651 11440 27683
rect 11472 27651 11512 27683
rect 11544 27651 11584 27683
rect 11616 27651 11656 27683
rect 11688 27651 11728 27683
rect 11760 27651 11800 27683
rect 11832 27651 11872 27683
rect 11904 27651 11944 27683
rect 11976 27651 12016 27683
rect 12048 27651 12088 27683
rect 12120 27651 12160 27683
rect 12192 27651 12232 27683
rect 12264 27651 12304 27683
rect 12336 27651 12376 27683
rect 12408 27651 12448 27683
rect 12480 27651 12520 27683
rect 12552 27651 12592 27683
rect 12624 27651 12664 27683
rect 12696 27651 12736 27683
rect 12768 27651 12808 27683
rect 12840 27651 12880 27683
rect 12912 27651 12952 27683
rect 12984 27651 13024 27683
rect 13056 27651 13096 27683
rect 13128 27651 13168 27683
rect 13200 27651 13240 27683
rect 13272 27651 13312 27683
rect 13344 27651 13384 27683
rect 13416 27651 13456 27683
rect 13488 27651 13528 27683
rect 13560 27651 13600 27683
rect 13632 27651 13672 27683
rect 13704 27651 13744 27683
rect 13776 27651 13816 27683
rect 13848 27651 13888 27683
rect 13920 27651 13960 27683
rect 13992 27651 14032 27683
rect 14064 27651 14104 27683
rect 14136 27651 14176 27683
rect 14208 27651 14248 27683
rect 14280 27651 14320 27683
rect 14352 27651 14392 27683
rect 14424 27651 14464 27683
rect 14496 27651 14536 27683
rect 14568 27651 14608 27683
rect 14640 27651 14680 27683
rect 14712 27651 14752 27683
rect 14784 27651 14824 27683
rect 14856 27651 14896 27683
rect 14928 27651 14968 27683
rect 15000 27651 15040 27683
rect 15072 27651 15112 27683
rect 15144 27651 15184 27683
rect 15216 27651 15256 27683
rect 15288 27651 15328 27683
rect 15360 27651 15400 27683
rect 15432 27651 15472 27683
rect 15504 27651 15544 27683
rect 15576 27651 15616 27683
rect 15648 27651 15688 27683
rect 15720 27651 15760 27683
rect 15792 27651 15832 27683
rect 15864 27651 15904 27683
rect 15936 27651 16000 27683
rect 0 27611 16000 27651
rect 0 27579 64 27611
rect 96 27579 136 27611
rect 168 27579 208 27611
rect 240 27579 280 27611
rect 312 27579 352 27611
rect 384 27579 424 27611
rect 456 27579 496 27611
rect 528 27579 568 27611
rect 600 27579 640 27611
rect 672 27579 712 27611
rect 744 27579 784 27611
rect 816 27579 856 27611
rect 888 27579 928 27611
rect 960 27579 1000 27611
rect 1032 27579 1072 27611
rect 1104 27579 1144 27611
rect 1176 27579 1216 27611
rect 1248 27579 1288 27611
rect 1320 27579 1360 27611
rect 1392 27579 1432 27611
rect 1464 27579 1504 27611
rect 1536 27579 1576 27611
rect 1608 27579 1648 27611
rect 1680 27579 1720 27611
rect 1752 27579 1792 27611
rect 1824 27579 1864 27611
rect 1896 27579 1936 27611
rect 1968 27579 2008 27611
rect 2040 27579 2080 27611
rect 2112 27579 2152 27611
rect 2184 27579 2224 27611
rect 2256 27579 2296 27611
rect 2328 27579 2368 27611
rect 2400 27579 2440 27611
rect 2472 27579 2512 27611
rect 2544 27579 2584 27611
rect 2616 27579 2656 27611
rect 2688 27579 2728 27611
rect 2760 27579 2800 27611
rect 2832 27579 2872 27611
rect 2904 27579 2944 27611
rect 2976 27579 3016 27611
rect 3048 27579 3088 27611
rect 3120 27579 3160 27611
rect 3192 27579 3232 27611
rect 3264 27579 3304 27611
rect 3336 27579 3376 27611
rect 3408 27579 3448 27611
rect 3480 27579 3520 27611
rect 3552 27579 3592 27611
rect 3624 27579 3664 27611
rect 3696 27579 3736 27611
rect 3768 27579 3808 27611
rect 3840 27579 3880 27611
rect 3912 27579 3952 27611
rect 3984 27579 4024 27611
rect 4056 27579 4096 27611
rect 4128 27579 4168 27611
rect 4200 27579 4240 27611
rect 4272 27579 4312 27611
rect 4344 27579 4384 27611
rect 4416 27579 4456 27611
rect 4488 27579 4528 27611
rect 4560 27579 4600 27611
rect 4632 27579 4672 27611
rect 4704 27579 4744 27611
rect 4776 27579 4816 27611
rect 4848 27579 4888 27611
rect 4920 27579 4960 27611
rect 4992 27579 5032 27611
rect 5064 27579 5104 27611
rect 5136 27579 5176 27611
rect 5208 27579 5248 27611
rect 5280 27579 5320 27611
rect 5352 27579 5392 27611
rect 5424 27579 5464 27611
rect 5496 27579 5536 27611
rect 5568 27579 5608 27611
rect 5640 27579 5680 27611
rect 5712 27579 5752 27611
rect 5784 27579 5824 27611
rect 5856 27579 5896 27611
rect 5928 27579 5968 27611
rect 6000 27579 6040 27611
rect 6072 27579 6112 27611
rect 6144 27579 6184 27611
rect 6216 27579 6256 27611
rect 6288 27579 6328 27611
rect 6360 27579 6400 27611
rect 6432 27579 6472 27611
rect 6504 27579 6544 27611
rect 6576 27579 6616 27611
rect 6648 27579 6688 27611
rect 6720 27579 6760 27611
rect 6792 27579 6832 27611
rect 6864 27579 6904 27611
rect 6936 27579 6976 27611
rect 7008 27579 7048 27611
rect 7080 27579 7120 27611
rect 7152 27579 7192 27611
rect 7224 27579 7264 27611
rect 7296 27579 7336 27611
rect 7368 27579 7408 27611
rect 7440 27579 7480 27611
rect 7512 27579 7552 27611
rect 7584 27579 7624 27611
rect 7656 27579 7696 27611
rect 7728 27579 7768 27611
rect 7800 27579 7840 27611
rect 7872 27579 7912 27611
rect 7944 27579 7984 27611
rect 8016 27579 8056 27611
rect 8088 27579 8128 27611
rect 8160 27579 8200 27611
rect 8232 27579 8272 27611
rect 8304 27579 8344 27611
rect 8376 27579 8416 27611
rect 8448 27579 8488 27611
rect 8520 27579 8560 27611
rect 8592 27579 8632 27611
rect 8664 27579 8704 27611
rect 8736 27579 8776 27611
rect 8808 27579 8848 27611
rect 8880 27579 8920 27611
rect 8952 27579 8992 27611
rect 9024 27579 9064 27611
rect 9096 27579 9136 27611
rect 9168 27579 9208 27611
rect 9240 27579 9280 27611
rect 9312 27579 9352 27611
rect 9384 27579 9424 27611
rect 9456 27579 9496 27611
rect 9528 27579 9568 27611
rect 9600 27579 9640 27611
rect 9672 27579 9712 27611
rect 9744 27579 9784 27611
rect 9816 27579 9856 27611
rect 9888 27579 9928 27611
rect 9960 27579 10000 27611
rect 10032 27579 10072 27611
rect 10104 27579 10144 27611
rect 10176 27579 10216 27611
rect 10248 27579 10288 27611
rect 10320 27579 10360 27611
rect 10392 27579 10432 27611
rect 10464 27579 10504 27611
rect 10536 27579 10576 27611
rect 10608 27579 10648 27611
rect 10680 27579 10720 27611
rect 10752 27579 10792 27611
rect 10824 27579 10864 27611
rect 10896 27579 10936 27611
rect 10968 27579 11008 27611
rect 11040 27579 11080 27611
rect 11112 27579 11152 27611
rect 11184 27579 11224 27611
rect 11256 27579 11296 27611
rect 11328 27579 11368 27611
rect 11400 27579 11440 27611
rect 11472 27579 11512 27611
rect 11544 27579 11584 27611
rect 11616 27579 11656 27611
rect 11688 27579 11728 27611
rect 11760 27579 11800 27611
rect 11832 27579 11872 27611
rect 11904 27579 11944 27611
rect 11976 27579 12016 27611
rect 12048 27579 12088 27611
rect 12120 27579 12160 27611
rect 12192 27579 12232 27611
rect 12264 27579 12304 27611
rect 12336 27579 12376 27611
rect 12408 27579 12448 27611
rect 12480 27579 12520 27611
rect 12552 27579 12592 27611
rect 12624 27579 12664 27611
rect 12696 27579 12736 27611
rect 12768 27579 12808 27611
rect 12840 27579 12880 27611
rect 12912 27579 12952 27611
rect 12984 27579 13024 27611
rect 13056 27579 13096 27611
rect 13128 27579 13168 27611
rect 13200 27579 13240 27611
rect 13272 27579 13312 27611
rect 13344 27579 13384 27611
rect 13416 27579 13456 27611
rect 13488 27579 13528 27611
rect 13560 27579 13600 27611
rect 13632 27579 13672 27611
rect 13704 27579 13744 27611
rect 13776 27579 13816 27611
rect 13848 27579 13888 27611
rect 13920 27579 13960 27611
rect 13992 27579 14032 27611
rect 14064 27579 14104 27611
rect 14136 27579 14176 27611
rect 14208 27579 14248 27611
rect 14280 27579 14320 27611
rect 14352 27579 14392 27611
rect 14424 27579 14464 27611
rect 14496 27579 14536 27611
rect 14568 27579 14608 27611
rect 14640 27579 14680 27611
rect 14712 27579 14752 27611
rect 14784 27579 14824 27611
rect 14856 27579 14896 27611
rect 14928 27579 14968 27611
rect 15000 27579 15040 27611
rect 15072 27579 15112 27611
rect 15144 27579 15184 27611
rect 15216 27579 15256 27611
rect 15288 27579 15328 27611
rect 15360 27579 15400 27611
rect 15432 27579 15472 27611
rect 15504 27579 15544 27611
rect 15576 27579 15616 27611
rect 15648 27579 15688 27611
rect 15720 27579 15760 27611
rect 15792 27579 15832 27611
rect 15864 27579 15904 27611
rect 15936 27579 16000 27611
rect 0 27539 16000 27579
rect 0 27507 64 27539
rect 96 27507 136 27539
rect 168 27507 208 27539
rect 240 27507 280 27539
rect 312 27507 352 27539
rect 384 27507 424 27539
rect 456 27507 496 27539
rect 528 27507 568 27539
rect 600 27507 640 27539
rect 672 27507 712 27539
rect 744 27507 784 27539
rect 816 27507 856 27539
rect 888 27507 928 27539
rect 960 27507 1000 27539
rect 1032 27507 1072 27539
rect 1104 27507 1144 27539
rect 1176 27507 1216 27539
rect 1248 27507 1288 27539
rect 1320 27507 1360 27539
rect 1392 27507 1432 27539
rect 1464 27507 1504 27539
rect 1536 27507 1576 27539
rect 1608 27507 1648 27539
rect 1680 27507 1720 27539
rect 1752 27507 1792 27539
rect 1824 27507 1864 27539
rect 1896 27507 1936 27539
rect 1968 27507 2008 27539
rect 2040 27507 2080 27539
rect 2112 27507 2152 27539
rect 2184 27507 2224 27539
rect 2256 27507 2296 27539
rect 2328 27507 2368 27539
rect 2400 27507 2440 27539
rect 2472 27507 2512 27539
rect 2544 27507 2584 27539
rect 2616 27507 2656 27539
rect 2688 27507 2728 27539
rect 2760 27507 2800 27539
rect 2832 27507 2872 27539
rect 2904 27507 2944 27539
rect 2976 27507 3016 27539
rect 3048 27507 3088 27539
rect 3120 27507 3160 27539
rect 3192 27507 3232 27539
rect 3264 27507 3304 27539
rect 3336 27507 3376 27539
rect 3408 27507 3448 27539
rect 3480 27507 3520 27539
rect 3552 27507 3592 27539
rect 3624 27507 3664 27539
rect 3696 27507 3736 27539
rect 3768 27507 3808 27539
rect 3840 27507 3880 27539
rect 3912 27507 3952 27539
rect 3984 27507 4024 27539
rect 4056 27507 4096 27539
rect 4128 27507 4168 27539
rect 4200 27507 4240 27539
rect 4272 27507 4312 27539
rect 4344 27507 4384 27539
rect 4416 27507 4456 27539
rect 4488 27507 4528 27539
rect 4560 27507 4600 27539
rect 4632 27507 4672 27539
rect 4704 27507 4744 27539
rect 4776 27507 4816 27539
rect 4848 27507 4888 27539
rect 4920 27507 4960 27539
rect 4992 27507 5032 27539
rect 5064 27507 5104 27539
rect 5136 27507 5176 27539
rect 5208 27507 5248 27539
rect 5280 27507 5320 27539
rect 5352 27507 5392 27539
rect 5424 27507 5464 27539
rect 5496 27507 5536 27539
rect 5568 27507 5608 27539
rect 5640 27507 5680 27539
rect 5712 27507 5752 27539
rect 5784 27507 5824 27539
rect 5856 27507 5896 27539
rect 5928 27507 5968 27539
rect 6000 27507 6040 27539
rect 6072 27507 6112 27539
rect 6144 27507 6184 27539
rect 6216 27507 6256 27539
rect 6288 27507 6328 27539
rect 6360 27507 6400 27539
rect 6432 27507 6472 27539
rect 6504 27507 6544 27539
rect 6576 27507 6616 27539
rect 6648 27507 6688 27539
rect 6720 27507 6760 27539
rect 6792 27507 6832 27539
rect 6864 27507 6904 27539
rect 6936 27507 6976 27539
rect 7008 27507 7048 27539
rect 7080 27507 7120 27539
rect 7152 27507 7192 27539
rect 7224 27507 7264 27539
rect 7296 27507 7336 27539
rect 7368 27507 7408 27539
rect 7440 27507 7480 27539
rect 7512 27507 7552 27539
rect 7584 27507 7624 27539
rect 7656 27507 7696 27539
rect 7728 27507 7768 27539
rect 7800 27507 7840 27539
rect 7872 27507 7912 27539
rect 7944 27507 7984 27539
rect 8016 27507 8056 27539
rect 8088 27507 8128 27539
rect 8160 27507 8200 27539
rect 8232 27507 8272 27539
rect 8304 27507 8344 27539
rect 8376 27507 8416 27539
rect 8448 27507 8488 27539
rect 8520 27507 8560 27539
rect 8592 27507 8632 27539
rect 8664 27507 8704 27539
rect 8736 27507 8776 27539
rect 8808 27507 8848 27539
rect 8880 27507 8920 27539
rect 8952 27507 8992 27539
rect 9024 27507 9064 27539
rect 9096 27507 9136 27539
rect 9168 27507 9208 27539
rect 9240 27507 9280 27539
rect 9312 27507 9352 27539
rect 9384 27507 9424 27539
rect 9456 27507 9496 27539
rect 9528 27507 9568 27539
rect 9600 27507 9640 27539
rect 9672 27507 9712 27539
rect 9744 27507 9784 27539
rect 9816 27507 9856 27539
rect 9888 27507 9928 27539
rect 9960 27507 10000 27539
rect 10032 27507 10072 27539
rect 10104 27507 10144 27539
rect 10176 27507 10216 27539
rect 10248 27507 10288 27539
rect 10320 27507 10360 27539
rect 10392 27507 10432 27539
rect 10464 27507 10504 27539
rect 10536 27507 10576 27539
rect 10608 27507 10648 27539
rect 10680 27507 10720 27539
rect 10752 27507 10792 27539
rect 10824 27507 10864 27539
rect 10896 27507 10936 27539
rect 10968 27507 11008 27539
rect 11040 27507 11080 27539
rect 11112 27507 11152 27539
rect 11184 27507 11224 27539
rect 11256 27507 11296 27539
rect 11328 27507 11368 27539
rect 11400 27507 11440 27539
rect 11472 27507 11512 27539
rect 11544 27507 11584 27539
rect 11616 27507 11656 27539
rect 11688 27507 11728 27539
rect 11760 27507 11800 27539
rect 11832 27507 11872 27539
rect 11904 27507 11944 27539
rect 11976 27507 12016 27539
rect 12048 27507 12088 27539
rect 12120 27507 12160 27539
rect 12192 27507 12232 27539
rect 12264 27507 12304 27539
rect 12336 27507 12376 27539
rect 12408 27507 12448 27539
rect 12480 27507 12520 27539
rect 12552 27507 12592 27539
rect 12624 27507 12664 27539
rect 12696 27507 12736 27539
rect 12768 27507 12808 27539
rect 12840 27507 12880 27539
rect 12912 27507 12952 27539
rect 12984 27507 13024 27539
rect 13056 27507 13096 27539
rect 13128 27507 13168 27539
rect 13200 27507 13240 27539
rect 13272 27507 13312 27539
rect 13344 27507 13384 27539
rect 13416 27507 13456 27539
rect 13488 27507 13528 27539
rect 13560 27507 13600 27539
rect 13632 27507 13672 27539
rect 13704 27507 13744 27539
rect 13776 27507 13816 27539
rect 13848 27507 13888 27539
rect 13920 27507 13960 27539
rect 13992 27507 14032 27539
rect 14064 27507 14104 27539
rect 14136 27507 14176 27539
rect 14208 27507 14248 27539
rect 14280 27507 14320 27539
rect 14352 27507 14392 27539
rect 14424 27507 14464 27539
rect 14496 27507 14536 27539
rect 14568 27507 14608 27539
rect 14640 27507 14680 27539
rect 14712 27507 14752 27539
rect 14784 27507 14824 27539
rect 14856 27507 14896 27539
rect 14928 27507 14968 27539
rect 15000 27507 15040 27539
rect 15072 27507 15112 27539
rect 15144 27507 15184 27539
rect 15216 27507 15256 27539
rect 15288 27507 15328 27539
rect 15360 27507 15400 27539
rect 15432 27507 15472 27539
rect 15504 27507 15544 27539
rect 15576 27507 15616 27539
rect 15648 27507 15688 27539
rect 15720 27507 15760 27539
rect 15792 27507 15832 27539
rect 15864 27507 15904 27539
rect 15936 27507 16000 27539
rect 0 27467 16000 27507
rect 0 27435 64 27467
rect 96 27435 136 27467
rect 168 27435 208 27467
rect 240 27435 280 27467
rect 312 27435 352 27467
rect 384 27435 424 27467
rect 456 27435 496 27467
rect 528 27435 568 27467
rect 600 27435 640 27467
rect 672 27435 712 27467
rect 744 27435 784 27467
rect 816 27435 856 27467
rect 888 27435 928 27467
rect 960 27435 1000 27467
rect 1032 27435 1072 27467
rect 1104 27435 1144 27467
rect 1176 27435 1216 27467
rect 1248 27435 1288 27467
rect 1320 27435 1360 27467
rect 1392 27435 1432 27467
rect 1464 27435 1504 27467
rect 1536 27435 1576 27467
rect 1608 27435 1648 27467
rect 1680 27435 1720 27467
rect 1752 27435 1792 27467
rect 1824 27435 1864 27467
rect 1896 27435 1936 27467
rect 1968 27435 2008 27467
rect 2040 27435 2080 27467
rect 2112 27435 2152 27467
rect 2184 27435 2224 27467
rect 2256 27435 2296 27467
rect 2328 27435 2368 27467
rect 2400 27435 2440 27467
rect 2472 27435 2512 27467
rect 2544 27435 2584 27467
rect 2616 27435 2656 27467
rect 2688 27435 2728 27467
rect 2760 27435 2800 27467
rect 2832 27435 2872 27467
rect 2904 27435 2944 27467
rect 2976 27435 3016 27467
rect 3048 27435 3088 27467
rect 3120 27435 3160 27467
rect 3192 27435 3232 27467
rect 3264 27435 3304 27467
rect 3336 27435 3376 27467
rect 3408 27435 3448 27467
rect 3480 27435 3520 27467
rect 3552 27435 3592 27467
rect 3624 27435 3664 27467
rect 3696 27435 3736 27467
rect 3768 27435 3808 27467
rect 3840 27435 3880 27467
rect 3912 27435 3952 27467
rect 3984 27435 4024 27467
rect 4056 27435 4096 27467
rect 4128 27435 4168 27467
rect 4200 27435 4240 27467
rect 4272 27435 4312 27467
rect 4344 27435 4384 27467
rect 4416 27435 4456 27467
rect 4488 27435 4528 27467
rect 4560 27435 4600 27467
rect 4632 27435 4672 27467
rect 4704 27435 4744 27467
rect 4776 27435 4816 27467
rect 4848 27435 4888 27467
rect 4920 27435 4960 27467
rect 4992 27435 5032 27467
rect 5064 27435 5104 27467
rect 5136 27435 5176 27467
rect 5208 27435 5248 27467
rect 5280 27435 5320 27467
rect 5352 27435 5392 27467
rect 5424 27435 5464 27467
rect 5496 27435 5536 27467
rect 5568 27435 5608 27467
rect 5640 27435 5680 27467
rect 5712 27435 5752 27467
rect 5784 27435 5824 27467
rect 5856 27435 5896 27467
rect 5928 27435 5968 27467
rect 6000 27435 6040 27467
rect 6072 27435 6112 27467
rect 6144 27435 6184 27467
rect 6216 27435 6256 27467
rect 6288 27435 6328 27467
rect 6360 27435 6400 27467
rect 6432 27435 6472 27467
rect 6504 27435 6544 27467
rect 6576 27435 6616 27467
rect 6648 27435 6688 27467
rect 6720 27435 6760 27467
rect 6792 27435 6832 27467
rect 6864 27435 6904 27467
rect 6936 27435 6976 27467
rect 7008 27435 7048 27467
rect 7080 27435 7120 27467
rect 7152 27435 7192 27467
rect 7224 27435 7264 27467
rect 7296 27435 7336 27467
rect 7368 27435 7408 27467
rect 7440 27435 7480 27467
rect 7512 27435 7552 27467
rect 7584 27435 7624 27467
rect 7656 27435 7696 27467
rect 7728 27435 7768 27467
rect 7800 27435 7840 27467
rect 7872 27435 7912 27467
rect 7944 27435 7984 27467
rect 8016 27435 8056 27467
rect 8088 27435 8128 27467
rect 8160 27435 8200 27467
rect 8232 27435 8272 27467
rect 8304 27435 8344 27467
rect 8376 27435 8416 27467
rect 8448 27435 8488 27467
rect 8520 27435 8560 27467
rect 8592 27435 8632 27467
rect 8664 27435 8704 27467
rect 8736 27435 8776 27467
rect 8808 27435 8848 27467
rect 8880 27435 8920 27467
rect 8952 27435 8992 27467
rect 9024 27435 9064 27467
rect 9096 27435 9136 27467
rect 9168 27435 9208 27467
rect 9240 27435 9280 27467
rect 9312 27435 9352 27467
rect 9384 27435 9424 27467
rect 9456 27435 9496 27467
rect 9528 27435 9568 27467
rect 9600 27435 9640 27467
rect 9672 27435 9712 27467
rect 9744 27435 9784 27467
rect 9816 27435 9856 27467
rect 9888 27435 9928 27467
rect 9960 27435 10000 27467
rect 10032 27435 10072 27467
rect 10104 27435 10144 27467
rect 10176 27435 10216 27467
rect 10248 27435 10288 27467
rect 10320 27435 10360 27467
rect 10392 27435 10432 27467
rect 10464 27435 10504 27467
rect 10536 27435 10576 27467
rect 10608 27435 10648 27467
rect 10680 27435 10720 27467
rect 10752 27435 10792 27467
rect 10824 27435 10864 27467
rect 10896 27435 10936 27467
rect 10968 27435 11008 27467
rect 11040 27435 11080 27467
rect 11112 27435 11152 27467
rect 11184 27435 11224 27467
rect 11256 27435 11296 27467
rect 11328 27435 11368 27467
rect 11400 27435 11440 27467
rect 11472 27435 11512 27467
rect 11544 27435 11584 27467
rect 11616 27435 11656 27467
rect 11688 27435 11728 27467
rect 11760 27435 11800 27467
rect 11832 27435 11872 27467
rect 11904 27435 11944 27467
rect 11976 27435 12016 27467
rect 12048 27435 12088 27467
rect 12120 27435 12160 27467
rect 12192 27435 12232 27467
rect 12264 27435 12304 27467
rect 12336 27435 12376 27467
rect 12408 27435 12448 27467
rect 12480 27435 12520 27467
rect 12552 27435 12592 27467
rect 12624 27435 12664 27467
rect 12696 27435 12736 27467
rect 12768 27435 12808 27467
rect 12840 27435 12880 27467
rect 12912 27435 12952 27467
rect 12984 27435 13024 27467
rect 13056 27435 13096 27467
rect 13128 27435 13168 27467
rect 13200 27435 13240 27467
rect 13272 27435 13312 27467
rect 13344 27435 13384 27467
rect 13416 27435 13456 27467
rect 13488 27435 13528 27467
rect 13560 27435 13600 27467
rect 13632 27435 13672 27467
rect 13704 27435 13744 27467
rect 13776 27435 13816 27467
rect 13848 27435 13888 27467
rect 13920 27435 13960 27467
rect 13992 27435 14032 27467
rect 14064 27435 14104 27467
rect 14136 27435 14176 27467
rect 14208 27435 14248 27467
rect 14280 27435 14320 27467
rect 14352 27435 14392 27467
rect 14424 27435 14464 27467
rect 14496 27435 14536 27467
rect 14568 27435 14608 27467
rect 14640 27435 14680 27467
rect 14712 27435 14752 27467
rect 14784 27435 14824 27467
rect 14856 27435 14896 27467
rect 14928 27435 14968 27467
rect 15000 27435 15040 27467
rect 15072 27435 15112 27467
rect 15144 27435 15184 27467
rect 15216 27435 15256 27467
rect 15288 27435 15328 27467
rect 15360 27435 15400 27467
rect 15432 27435 15472 27467
rect 15504 27435 15544 27467
rect 15576 27435 15616 27467
rect 15648 27435 15688 27467
rect 15720 27435 15760 27467
rect 15792 27435 15832 27467
rect 15864 27435 15904 27467
rect 15936 27435 16000 27467
rect 0 27395 16000 27435
rect 0 27363 64 27395
rect 96 27363 136 27395
rect 168 27363 208 27395
rect 240 27363 280 27395
rect 312 27363 352 27395
rect 384 27363 424 27395
rect 456 27363 496 27395
rect 528 27363 568 27395
rect 600 27363 640 27395
rect 672 27363 712 27395
rect 744 27363 784 27395
rect 816 27363 856 27395
rect 888 27363 928 27395
rect 960 27363 1000 27395
rect 1032 27363 1072 27395
rect 1104 27363 1144 27395
rect 1176 27363 1216 27395
rect 1248 27363 1288 27395
rect 1320 27363 1360 27395
rect 1392 27363 1432 27395
rect 1464 27363 1504 27395
rect 1536 27363 1576 27395
rect 1608 27363 1648 27395
rect 1680 27363 1720 27395
rect 1752 27363 1792 27395
rect 1824 27363 1864 27395
rect 1896 27363 1936 27395
rect 1968 27363 2008 27395
rect 2040 27363 2080 27395
rect 2112 27363 2152 27395
rect 2184 27363 2224 27395
rect 2256 27363 2296 27395
rect 2328 27363 2368 27395
rect 2400 27363 2440 27395
rect 2472 27363 2512 27395
rect 2544 27363 2584 27395
rect 2616 27363 2656 27395
rect 2688 27363 2728 27395
rect 2760 27363 2800 27395
rect 2832 27363 2872 27395
rect 2904 27363 2944 27395
rect 2976 27363 3016 27395
rect 3048 27363 3088 27395
rect 3120 27363 3160 27395
rect 3192 27363 3232 27395
rect 3264 27363 3304 27395
rect 3336 27363 3376 27395
rect 3408 27363 3448 27395
rect 3480 27363 3520 27395
rect 3552 27363 3592 27395
rect 3624 27363 3664 27395
rect 3696 27363 3736 27395
rect 3768 27363 3808 27395
rect 3840 27363 3880 27395
rect 3912 27363 3952 27395
rect 3984 27363 4024 27395
rect 4056 27363 4096 27395
rect 4128 27363 4168 27395
rect 4200 27363 4240 27395
rect 4272 27363 4312 27395
rect 4344 27363 4384 27395
rect 4416 27363 4456 27395
rect 4488 27363 4528 27395
rect 4560 27363 4600 27395
rect 4632 27363 4672 27395
rect 4704 27363 4744 27395
rect 4776 27363 4816 27395
rect 4848 27363 4888 27395
rect 4920 27363 4960 27395
rect 4992 27363 5032 27395
rect 5064 27363 5104 27395
rect 5136 27363 5176 27395
rect 5208 27363 5248 27395
rect 5280 27363 5320 27395
rect 5352 27363 5392 27395
rect 5424 27363 5464 27395
rect 5496 27363 5536 27395
rect 5568 27363 5608 27395
rect 5640 27363 5680 27395
rect 5712 27363 5752 27395
rect 5784 27363 5824 27395
rect 5856 27363 5896 27395
rect 5928 27363 5968 27395
rect 6000 27363 6040 27395
rect 6072 27363 6112 27395
rect 6144 27363 6184 27395
rect 6216 27363 6256 27395
rect 6288 27363 6328 27395
rect 6360 27363 6400 27395
rect 6432 27363 6472 27395
rect 6504 27363 6544 27395
rect 6576 27363 6616 27395
rect 6648 27363 6688 27395
rect 6720 27363 6760 27395
rect 6792 27363 6832 27395
rect 6864 27363 6904 27395
rect 6936 27363 6976 27395
rect 7008 27363 7048 27395
rect 7080 27363 7120 27395
rect 7152 27363 7192 27395
rect 7224 27363 7264 27395
rect 7296 27363 7336 27395
rect 7368 27363 7408 27395
rect 7440 27363 7480 27395
rect 7512 27363 7552 27395
rect 7584 27363 7624 27395
rect 7656 27363 7696 27395
rect 7728 27363 7768 27395
rect 7800 27363 7840 27395
rect 7872 27363 7912 27395
rect 7944 27363 7984 27395
rect 8016 27363 8056 27395
rect 8088 27363 8128 27395
rect 8160 27363 8200 27395
rect 8232 27363 8272 27395
rect 8304 27363 8344 27395
rect 8376 27363 8416 27395
rect 8448 27363 8488 27395
rect 8520 27363 8560 27395
rect 8592 27363 8632 27395
rect 8664 27363 8704 27395
rect 8736 27363 8776 27395
rect 8808 27363 8848 27395
rect 8880 27363 8920 27395
rect 8952 27363 8992 27395
rect 9024 27363 9064 27395
rect 9096 27363 9136 27395
rect 9168 27363 9208 27395
rect 9240 27363 9280 27395
rect 9312 27363 9352 27395
rect 9384 27363 9424 27395
rect 9456 27363 9496 27395
rect 9528 27363 9568 27395
rect 9600 27363 9640 27395
rect 9672 27363 9712 27395
rect 9744 27363 9784 27395
rect 9816 27363 9856 27395
rect 9888 27363 9928 27395
rect 9960 27363 10000 27395
rect 10032 27363 10072 27395
rect 10104 27363 10144 27395
rect 10176 27363 10216 27395
rect 10248 27363 10288 27395
rect 10320 27363 10360 27395
rect 10392 27363 10432 27395
rect 10464 27363 10504 27395
rect 10536 27363 10576 27395
rect 10608 27363 10648 27395
rect 10680 27363 10720 27395
rect 10752 27363 10792 27395
rect 10824 27363 10864 27395
rect 10896 27363 10936 27395
rect 10968 27363 11008 27395
rect 11040 27363 11080 27395
rect 11112 27363 11152 27395
rect 11184 27363 11224 27395
rect 11256 27363 11296 27395
rect 11328 27363 11368 27395
rect 11400 27363 11440 27395
rect 11472 27363 11512 27395
rect 11544 27363 11584 27395
rect 11616 27363 11656 27395
rect 11688 27363 11728 27395
rect 11760 27363 11800 27395
rect 11832 27363 11872 27395
rect 11904 27363 11944 27395
rect 11976 27363 12016 27395
rect 12048 27363 12088 27395
rect 12120 27363 12160 27395
rect 12192 27363 12232 27395
rect 12264 27363 12304 27395
rect 12336 27363 12376 27395
rect 12408 27363 12448 27395
rect 12480 27363 12520 27395
rect 12552 27363 12592 27395
rect 12624 27363 12664 27395
rect 12696 27363 12736 27395
rect 12768 27363 12808 27395
rect 12840 27363 12880 27395
rect 12912 27363 12952 27395
rect 12984 27363 13024 27395
rect 13056 27363 13096 27395
rect 13128 27363 13168 27395
rect 13200 27363 13240 27395
rect 13272 27363 13312 27395
rect 13344 27363 13384 27395
rect 13416 27363 13456 27395
rect 13488 27363 13528 27395
rect 13560 27363 13600 27395
rect 13632 27363 13672 27395
rect 13704 27363 13744 27395
rect 13776 27363 13816 27395
rect 13848 27363 13888 27395
rect 13920 27363 13960 27395
rect 13992 27363 14032 27395
rect 14064 27363 14104 27395
rect 14136 27363 14176 27395
rect 14208 27363 14248 27395
rect 14280 27363 14320 27395
rect 14352 27363 14392 27395
rect 14424 27363 14464 27395
rect 14496 27363 14536 27395
rect 14568 27363 14608 27395
rect 14640 27363 14680 27395
rect 14712 27363 14752 27395
rect 14784 27363 14824 27395
rect 14856 27363 14896 27395
rect 14928 27363 14968 27395
rect 15000 27363 15040 27395
rect 15072 27363 15112 27395
rect 15144 27363 15184 27395
rect 15216 27363 15256 27395
rect 15288 27363 15328 27395
rect 15360 27363 15400 27395
rect 15432 27363 15472 27395
rect 15504 27363 15544 27395
rect 15576 27363 15616 27395
rect 15648 27363 15688 27395
rect 15720 27363 15760 27395
rect 15792 27363 15832 27395
rect 15864 27363 15904 27395
rect 15936 27363 16000 27395
rect 0 27323 16000 27363
rect 0 27291 64 27323
rect 96 27291 136 27323
rect 168 27291 208 27323
rect 240 27291 280 27323
rect 312 27291 352 27323
rect 384 27291 424 27323
rect 456 27291 496 27323
rect 528 27291 568 27323
rect 600 27291 640 27323
rect 672 27291 712 27323
rect 744 27291 784 27323
rect 816 27291 856 27323
rect 888 27291 928 27323
rect 960 27291 1000 27323
rect 1032 27291 1072 27323
rect 1104 27291 1144 27323
rect 1176 27291 1216 27323
rect 1248 27291 1288 27323
rect 1320 27291 1360 27323
rect 1392 27291 1432 27323
rect 1464 27291 1504 27323
rect 1536 27291 1576 27323
rect 1608 27291 1648 27323
rect 1680 27291 1720 27323
rect 1752 27291 1792 27323
rect 1824 27291 1864 27323
rect 1896 27291 1936 27323
rect 1968 27291 2008 27323
rect 2040 27291 2080 27323
rect 2112 27291 2152 27323
rect 2184 27291 2224 27323
rect 2256 27291 2296 27323
rect 2328 27291 2368 27323
rect 2400 27291 2440 27323
rect 2472 27291 2512 27323
rect 2544 27291 2584 27323
rect 2616 27291 2656 27323
rect 2688 27291 2728 27323
rect 2760 27291 2800 27323
rect 2832 27291 2872 27323
rect 2904 27291 2944 27323
rect 2976 27291 3016 27323
rect 3048 27291 3088 27323
rect 3120 27291 3160 27323
rect 3192 27291 3232 27323
rect 3264 27291 3304 27323
rect 3336 27291 3376 27323
rect 3408 27291 3448 27323
rect 3480 27291 3520 27323
rect 3552 27291 3592 27323
rect 3624 27291 3664 27323
rect 3696 27291 3736 27323
rect 3768 27291 3808 27323
rect 3840 27291 3880 27323
rect 3912 27291 3952 27323
rect 3984 27291 4024 27323
rect 4056 27291 4096 27323
rect 4128 27291 4168 27323
rect 4200 27291 4240 27323
rect 4272 27291 4312 27323
rect 4344 27291 4384 27323
rect 4416 27291 4456 27323
rect 4488 27291 4528 27323
rect 4560 27291 4600 27323
rect 4632 27291 4672 27323
rect 4704 27291 4744 27323
rect 4776 27291 4816 27323
rect 4848 27291 4888 27323
rect 4920 27291 4960 27323
rect 4992 27291 5032 27323
rect 5064 27291 5104 27323
rect 5136 27291 5176 27323
rect 5208 27291 5248 27323
rect 5280 27291 5320 27323
rect 5352 27291 5392 27323
rect 5424 27291 5464 27323
rect 5496 27291 5536 27323
rect 5568 27291 5608 27323
rect 5640 27291 5680 27323
rect 5712 27291 5752 27323
rect 5784 27291 5824 27323
rect 5856 27291 5896 27323
rect 5928 27291 5968 27323
rect 6000 27291 6040 27323
rect 6072 27291 6112 27323
rect 6144 27291 6184 27323
rect 6216 27291 6256 27323
rect 6288 27291 6328 27323
rect 6360 27291 6400 27323
rect 6432 27291 6472 27323
rect 6504 27291 6544 27323
rect 6576 27291 6616 27323
rect 6648 27291 6688 27323
rect 6720 27291 6760 27323
rect 6792 27291 6832 27323
rect 6864 27291 6904 27323
rect 6936 27291 6976 27323
rect 7008 27291 7048 27323
rect 7080 27291 7120 27323
rect 7152 27291 7192 27323
rect 7224 27291 7264 27323
rect 7296 27291 7336 27323
rect 7368 27291 7408 27323
rect 7440 27291 7480 27323
rect 7512 27291 7552 27323
rect 7584 27291 7624 27323
rect 7656 27291 7696 27323
rect 7728 27291 7768 27323
rect 7800 27291 7840 27323
rect 7872 27291 7912 27323
rect 7944 27291 7984 27323
rect 8016 27291 8056 27323
rect 8088 27291 8128 27323
rect 8160 27291 8200 27323
rect 8232 27291 8272 27323
rect 8304 27291 8344 27323
rect 8376 27291 8416 27323
rect 8448 27291 8488 27323
rect 8520 27291 8560 27323
rect 8592 27291 8632 27323
rect 8664 27291 8704 27323
rect 8736 27291 8776 27323
rect 8808 27291 8848 27323
rect 8880 27291 8920 27323
rect 8952 27291 8992 27323
rect 9024 27291 9064 27323
rect 9096 27291 9136 27323
rect 9168 27291 9208 27323
rect 9240 27291 9280 27323
rect 9312 27291 9352 27323
rect 9384 27291 9424 27323
rect 9456 27291 9496 27323
rect 9528 27291 9568 27323
rect 9600 27291 9640 27323
rect 9672 27291 9712 27323
rect 9744 27291 9784 27323
rect 9816 27291 9856 27323
rect 9888 27291 9928 27323
rect 9960 27291 10000 27323
rect 10032 27291 10072 27323
rect 10104 27291 10144 27323
rect 10176 27291 10216 27323
rect 10248 27291 10288 27323
rect 10320 27291 10360 27323
rect 10392 27291 10432 27323
rect 10464 27291 10504 27323
rect 10536 27291 10576 27323
rect 10608 27291 10648 27323
rect 10680 27291 10720 27323
rect 10752 27291 10792 27323
rect 10824 27291 10864 27323
rect 10896 27291 10936 27323
rect 10968 27291 11008 27323
rect 11040 27291 11080 27323
rect 11112 27291 11152 27323
rect 11184 27291 11224 27323
rect 11256 27291 11296 27323
rect 11328 27291 11368 27323
rect 11400 27291 11440 27323
rect 11472 27291 11512 27323
rect 11544 27291 11584 27323
rect 11616 27291 11656 27323
rect 11688 27291 11728 27323
rect 11760 27291 11800 27323
rect 11832 27291 11872 27323
rect 11904 27291 11944 27323
rect 11976 27291 12016 27323
rect 12048 27291 12088 27323
rect 12120 27291 12160 27323
rect 12192 27291 12232 27323
rect 12264 27291 12304 27323
rect 12336 27291 12376 27323
rect 12408 27291 12448 27323
rect 12480 27291 12520 27323
rect 12552 27291 12592 27323
rect 12624 27291 12664 27323
rect 12696 27291 12736 27323
rect 12768 27291 12808 27323
rect 12840 27291 12880 27323
rect 12912 27291 12952 27323
rect 12984 27291 13024 27323
rect 13056 27291 13096 27323
rect 13128 27291 13168 27323
rect 13200 27291 13240 27323
rect 13272 27291 13312 27323
rect 13344 27291 13384 27323
rect 13416 27291 13456 27323
rect 13488 27291 13528 27323
rect 13560 27291 13600 27323
rect 13632 27291 13672 27323
rect 13704 27291 13744 27323
rect 13776 27291 13816 27323
rect 13848 27291 13888 27323
rect 13920 27291 13960 27323
rect 13992 27291 14032 27323
rect 14064 27291 14104 27323
rect 14136 27291 14176 27323
rect 14208 27291 14248 27323
rect 14280 27291 14320 27323
rect 14352 27291 14392 27323
rect 14424 27291 14464 27323
rect 14496 27291 14536 27323
rect 14568 27291 14608 27323
rect 14640 27291 14680 27323
rect 14712 27291 14752 27323
rect 14784 27291 14824 27323
rect 14856 27291 14896 27323
rect 14928 27291 14968 27323
rect 15000 27291 15040 27323
rect 15072 27291 15112 27323
rect 15144 27291 15184 27323
rect 15216 27291 15256 27323
rect 15288 27291 15328 27323
rect 15360 27291 15400 27323
rect 15432 27291 15472 27323
rect 15504 27291 15544 27323
rect 15576 27291 15616 27323
rect 15648 27291 15688 27323
rect 15720 27291 15760 27323
rect 15792 27291 15832 27323
rect 15864 27291 15904 27323
rect 15936 27291 16000 27323
rect 0 27251 16000 27291
rect 0 27219 64 27251
rect 96 27219 136 27251
rect 168 27219 208 27251
rect 240 27219 280 27251
rect 312 27219 352 27251
rect 384 27219 424 27251
rect 456 27219 496 27251
rect 528 27219 568 27251
rect 600 27219 640 27251
rect 672 27219 712 27251
rect 744 27219 784 27251
rect 816 27219 856 27251
rect 888 27219 928 27251
rect 960 27219 1000 27251
rect 1032 27219 1072 27251
rect 1104 27219 1144 27251
rect 1176 27219 1216 27251
rect 1248 27219 1288 27251
rect 1320 27219 1360 27251
rect 1392 27219 1432 27251
rect 1464 27219 1504 27251
rect 1536 27219 1576 27251
rect 1608 27219 1648 27251
rect 1680 27219 1720 27251
rect 1752 27219 1792 27251
rect 1824 27219 1864 27251
rect 1896 27219 1936 27251
rect 1968 27219 2008 27251
rect 2040 27219 2080 27251
rect 2112 27219 2152 27251
rect 2184 27219 2224 27251
rect 2256 27219 2296 27251
rect 2328 27219 2368 27251
rect 2400 27219 2440 27251
rect 2472 27219 2512 27251
rect 2544 27219 2584 27251
rect 2616 27219 2656 27251
rect 2688 27219 2728 27251
rect 2760 27219 2800 27251
rect 2832 27219 2872 27251
rect 2904 27219 2944 27251
rect 2976 27219 3016 27251
rect 3048 27219 3088 27251
rect 3120 27219 3160 27251
rect 3192 27219 3232 27251
rect 3264 27219 3304 27251
rect 3336 27219 3376 27251
rect 3408 27219 3448 27251
rect 3480 27219 3520 27251
rect 3552 27219 3592 27251
rect 3624 27219 3664 27251
rect 3696 27219 3736 27251
rect 3768 27219 3808 27251
rect 3840 27219 3880 27251
rect 3912 27219 3952 27251
rect 3984 27219 4024 27251
rect 4056 27219 4096 27251
rect 4128 27219 4168 27251
rect 4200 27219 4240 27251
rect 4272 27219 4312 27251
rect 4344 27219 4384 27251
rect 4416 27219 4456 27251
rect 4488 27219 4528 27251
rect 4560 27219 4600 27251
rect 4632 27219 4672 27251
rect 4704 27219 4744 27251
rect 4776 27219 4816 27251
rect 4848 27219 4888 27251
rect 4920 27219 4960 27251
rect 4992 27219 5032 27251
rect 5064 27219 5104 27251
rect 5136 27219 5176 27251
rect 5208 27219 5248 27251
rect 5280 27219 5320 27251
rect 5352 27219 5392 27251
rect 5424 27219 5464 27251
rect 5496 27219 5536 27251
rect 5568 27219 5608 27251
rect 5640 27219 5680 27251
rect 5712 27219 5752 27251
rect 5784 27219 5824 27251
rect 5856 27219 5896 27251
rect 5928 27219 5968 27251
rect 6000 27219 6040 27251
rect 6072 27219 6112 27251
rect 6144 27219 6184 27251
rect 6216 27219 6256 27251
rect 6288 27219 6328 27251
rect 6360 27219 6400 27251
rect 6432 27219 6472 27251
rect 6504 27219 6544 27251
rect 6576 27219 6616 27251
rect 6648 27219 6688 27251
rect 6720 27219 6760 27251
rect 6792 27219 6832 27251
rect 6864 27219 6904 27251
rect 6936 27219 6976 27251
rect 7008 27219 7048 27251
rect 7080 27219 7120 27251
rect 7152 27219 7192 27251
rect 7224 27219 7264 27251
rect 7296 27219 7336 27251
rect 7368 27219 7408 27251
rect 7440 27219 7480 27251
rect 7512 27219 7552 27251
rect 7584 27219 7624 27251
rect 7656 27219 7696 27251
rect 7728 27219 7768 27251
rect 7800 27219 7840 27251
rect 7872 27219 7912 27251
rect 7944 27219 7984 27251
rect 8016 27219 8056 27251
rect 8088 27219 8128 27251
rect 8160 27219 8200 27251
rect 8232 27219 8272 27251
rect 8304 27219 8344 27251
rect 8376 27219 8416 27251
rect 8448 27219 8488 27251
rect 8520 27219 8560 27251
rect 8592 27219 8632 27251
rect 8664 27219 8704 27251
rect 8736 27219 8776 27251
rect 8808 27219 8848 27251
rect 8880 27219 8920 27251
rect 8952 27219 8992 27251
rect 9024 27219 9064 27251
rect 9096 27219 9136 27251
rect 9168 27219 9208 27251
rect 9240 27219 9280 27251
rect 9312 27219 9352 27251
rect 9384 27219 9424 27251
rect 9456 27219 9496 27251
rect 9528 27219 9568 27251
rect 9600 27219 9640 27251
rect 9672 27219 9712 27251
rect 9744 27219 9784 27251
rect 9816 27219 9856 27251
rect 9888 27219 9928 27251
rect 9960 27219 10000 27251
rect 10032 27219 10072 27251
rect 10104 27219 10144 27251
rect 10176 27219 10216 27251
rect 10248 27219 10288 27251
rect 10320 27219 10360 27251
rect 10392 27219 10432 27251
rect 10464 27219 10504 27251
rect 10536 27219 10576 27251
rect 10608 27219 10648 27251
rect 10680 27219 10720 27251
rect 10752 27219 10792 27251
rect 10824 27219 10864 27251
rect 10896 27219 10936 27251
rect 10968 27219 11008 27251
rect 11040 27219 11080 27251
rect 11112 27219 11152 27251
rect 11184 27219 11224 27251
rect 11256 27219 11296 27251
rect 11328 27219 11368 27251
rect 11400 27219 11440 27251
rect 11472 27219 11512 27251
rect 11544 27219 11584 27251
rect 11616 27219 11656 27251
rect 11688 27219 11728 27251
rect 11760 27219 11800 27251
rect 11832 27219 11872 27251
rect 11904 27219 11944 27251
rect 11976 27219 12016 27251
rect 12048 27219 12088 27251
rect 12120 27219 12160 27251
rect 12192 27219 12232 27251
rect 12264 27219 12304 27251
rect 12336 27219 12376 27251
rect 12408 27219 12448 27251
rect 12480 27219 12520 27251
rect 12552 27219 12592 27251
rect 12624 27219 12664 27251
rect 12696 27219 12736 27251
rect 12768 27219 12808 27251
rect 12840 27219 12880 27251
rect 12912 27219 12952 27251
rect 12984 27219 13024 27251
rect 13056 27219 13096 27251
rect 13128 27219 13168 27251
rect 13200 27219 13240 27251
rect 13272 27219 13312 27251
rect 13344 27219 13384 27251
rect 13416 27219 13456 27251
rect 13488 27219 13528 27251
rect 13560 27219 13600 27251
rect 13632 27219 13672 27251
rect 13704 27219 13744 27251
rect 13776 27219 13816 27251
rect 13848 27219 13888 27251
rect 13920 27219 13960 27251
rect 13992 27219 14032 27251
rect 14064 27219 14104 27251
rect 14136 27219 14176 27251
rect 14208 27219 14248 27251
rect 14280 27219 14320 27251
rect 14352 27219 14392 27251
rect 14424 27219 14464 27251
rect 14496 27219 14536 27251
rect 14568 27219 14608 27251
rect 14640 27219 14680 27251
rect 14712 27219 14752 27251
rect 14784 27219 14824 27251
rect 14856 27219 14896 27251
rect 14928 27219 14968 27251
rect 15000 27219 15040 27251
rect 15072 27219 15112 27251
rect 15144 27219 15184 27251
rect 15216 27219 15256 27251
rect 15288 27219 15328 27251
rect 15360 27219 15400 27251
rect 15432 27219 15472 27251
rect 15504 27219 15544 27251
rect 15576 27219 15616 27251
rect 15648 27219 15688 27251
rect 15720 27219 15760 27251
rect 15792 27219 15832 27251
rect 15864 27219 15904 27251
rect 15936 27219 16000 27251
rect 0 27179 16000 27219
rect 0 27147 64 27179
rect 96 27147 136 27179
rect 168 27147 208 27179
rect 240 27147 280 27179
rect 312 27147 352 27179
rect 384 27147 424 27179
rect 456 27147 496 27179
rect 528 27147 568 27179
rect 600 27147 640 27179
rect 672 27147 712 27179
rect 744 27147 784 27179
rect 816 27147 856 27179
rect 888 27147 928 27179
rect 960 27147 1000 27179
rect 1032 27147 1072 27179
rect 1104 27147 1144 27179
rect 1176 27147 1216 27179
rect 1248 27147 1288 27179
rect 1320 27147 1360 27179
rect 1392 27147 1432 27179
rect 1464 27147 1504 27179
rect 1536 27147 1576 27179
rect 1608 27147 1648 27179
rect 1680 27147 1720 27179
rect 1752 27147 1792 27179
rect 1824 27147 1864 27179
rect 1896 27147 1936 27179
rect 1968 27147 2008 27179
rect 2040 27147 2080 27179
rect 2112 27147 2152 27179
rect 2184 27147 2224 27179
rect 2256 27147 2296 27179
rect 2328 27147 2368 27179
rect 2400 27147 2440 27179
rect 2472 27147 2512 27179
rect 2544 27147 2584 27179
rect 2616 27147 2656 27179
rect 2688 27147 2728 27179
rect 2760 27147 2800 27179
rect 2832 27147 2872 27179
rect 2904 27147 2944 27179
rect 2976 27147 3016 27179
rect 3048 27147 3088 27179
rect 3120 27147 3160 27179
rect 3192 27147 3232 27179
rect 3264 27147 3304 27179
rect 3336 27147 3376 27179
rect 3408 27147 3448 27179
rect 3480 27147 3520 27179
rect 3552 27147 3592 27179
rect 3624 27147 3664 27179
rect 3696 27147 3736 27179
rect 3768 27147 3808 27179
rect 3840 27147 3880 27179
rect 3912 27147 3952 27179
rect 3984 27147 4024 27179
rect 4056 27147 4096 27179
rect 4128 27147 4168 27179
rect 4200 27147 4240 27179
rect 4272 27147 4312 27179
rect 4344 27147 4384 27179
rect 4416 27147 4456 27179
rect 4488 27147 4528 27179
rect 4560 27147 4600 27179
rect 4632 27147 4672 27179
rect 4704 27147 4744 27179
rect 4776 27147 4816 27179
rect 4848 27147 4888 27179
rect 4920 27147 4960 27179
rect 4992 27147 5032 27179
rect 5064 27147 5104 27179
rect 5136 27147 5176 27179
rect 5208 27147 5248 27179
rect 5280 27147 5320 27179
rect 5352 27147 5392 27179
rect 5424 27147 5464 27179
rect 5496 27147 5536 27179
rect 5568 27147 5608 27179
rect 5640 27147 5680 27179
rect 5712 27147 5752 27179
rect 5784 27147 5824 27179
rect 5856 27147 5896 27179
rect 5928 27147 5968 27179
rect 6000 27147 6040 27179
rect 6072 27147 6112 27179
rect 6144 27147 6184 27179
rect 6216 27147 6256 27179
rect 6288 27147 6328 27179
rect 6360 27147 6400 27179
rect 6432 27147 6472 27179
rect 6504 27147 6544 27179
rect 6576 27147 6616 27179
rect 6648 27147 6688 27179
rect 6720 27147 6760 27179
rect 6792 27147 6832 27179
rect 6864 27147 6904 27179
rect 6936 27147 6976 27179
rect 7008 27147 7048 27179
rect 7080 27147 7120 27179
rect 7152 27147 7192 27179
rect 7224 27147 7264 27179
rect 7296 27147 7336 27179
rect 7368 27147 7408 27179
rect 7440 27147 7480 27179
rect 7512 27147 7552 27179
rect 7584 27147 7624 27179
rect 7656 27147 7696 27179
rect 7728 27147 7768 27179
rect 7800 27147 7840 27179
rect 7872 27147 7912 27179
rect 7944 27147 7984 27179
rect 8016 27147 8056 27179
rect 8088 27147 8128 27179
rect 8160 27147 8200 27179
rect 8232 27147 8272 27179
rect 8304 27147 8344 27179
rect 8376 27147 8416 27179
rect 8448 27147 8488 27179
rect 8520 27147 8560 27179
rect 8592 27147 8632 27179
rect 8664 27147 8704 27179
rect 8736 27147 8776 27179
rect 8808 27147 8848 27179
rect 8880 27147 8920 27179
rect 8952 27147 8992 27179
rect 9024 27147 9064 27179
rect 9096 27147 9136 27179
rect 9168 27147 9208 27179
rect 9240 27147 9280 27179
rect 9312 27147 9352 27179
rect 9384 27147 9424 27179
rect 9456 27147 9496 27179
rect 9528 27147 9568 27179
rect 9600 27147 9640 27179
rect 9672 27147 9712 27179
rect 9744 27147 9784 27179
rect 9816 27147 9856 27179
rect 9888 27147 9928 27179
rect 9960 27147 10000 27179
rect 10032 27147 10072 27179
rect 10104 27147 10144 27179
rect 10176 27147 10216 27179
rect 10248 27147 10288 27179
rect 10320 27147 10360 27179
rect 10392 27147 10432 27179
rect 10464 27147 10504 27179
rect 10536 27147 10576 27179
rect 10608 27147 10648 27179
rect 10680 27147 10720 27179
rect 10752 27147 10792 27179
rect 10824 27147 10864 27179
rect 10896 27147 10936 27179
rect 10968 27147 11008 27179
rect 11040 27147 11080 27179
rect 11112 27147 11152 27179
rect 11184 27147 11224 27179
rect 11256 27147 11296 27179
rect 11328 27147 11368 27179
rect 11400 27147 11440 27179
rect 11472 27147 11512 27179
rect 11544 27147 11584 27179
rect 11616 27147 11656 27179
rect 11688 27147 11728 27179
rect 11760 27147 11800 27179
rect 11832 27147 11872 27179
rect 11904 27147 11944 27179
rect 11976 27147 12016 27179
rect 12048 27147 12088 27179
rect 12120 27147 12160 27179
rect 12192 27147 12232 27179
rect 12264 27147 12304 27179
rect 12336 27147 12376 27179
rect 12408 27147 12448 27179
rect 12480 27147 12520 27179
rect 12552 27147 12592 27179
rect 12624 27147 12664 27179
rect 12696 27147 12736 27179
rect 12768 27147 12808 27179
rect 12840 27147 12880 27179
rect 12912 27147 12952 27179
rect 12984 27147 13024 27179
rect 13056 27147 13096 27179
rect 13128 27147 13168 27179
rect 13200 27147 13240 27179
rect 13272 27147 13312 27179
rect 13344 27147 13384 27179
rect 13416 27147 13456 27179
rect 13488 27147 13528 27179
rect 13560 27147 13600 27179
rect 13632 27147 13672 27179
rect 13704 27147 13744 27179
rect 13776 27147 13816 27179
rect 13848 27147 13888 27179
rect 13920 27147 13960 27179
rect 13992 27147 14032 27179
rect 14064 27147 14104 27179
rect 14136 27147 14176 27179
rect 14208 27147 14248 27179
rect 14280 27147 14320 27179
rect 14352 27147 14392 27179
rect 14424 27147 14464 27179
rect 14496 27147 14536 27179
rect 14568 27147 14608 27179
rect 14640 27147 14680 27179
rect 14712 27147 14752 27179
rect 14784 27147 14824 27179
rect 14856 27147 14896 27179
rect 14928 27147 14968 27179
rect 15000 27147 15040 27179
rect 15072 27147 15112 27179
rect 15144 27147 15184 27179
rect 15216 27147 15256 27179
rect 15288 27147 15328 27179
rect 15360 27147 15400 27179
rect 15432 27147 15472 27179
rect 15504 27147 15544 27179
rect 15576 27147 15616 27179
rect 15648 27147 15688 27179
rect 15720 27147 15760 27179
rect 15792 27147 15832 27179
rect 15864 27147 15904 27179
rect 15936 27147 16000 27179
rect 0 27107 16000 27147
rect 0 27075 64 27107
rect 96 27075 136 27107
rect 168 27075 208 27107
rect 240 27075 280 27107
rect 312 27075 352 27107
rect 384 27075 424 27107
rect 456 27075 496 27107
rect 528 27075 568 27107
rect 600 27075 640 27107
rect 672 27075 712 27107
rect 744 27075 784 27107
rect 816 27075 856 27107
rect 888 27075 928 27107
rect 960 27075 1000 27107
rect 1032 27075 1072 27107
rect 1104 27075 1144 27107
rect 1176 27075 1216 27107
rect 1248 27075 1288 27107
rect 1320 27075 1360 27107
rect 1392 27075 1432 27107
rect 1464 27075 1504 27107
rect 1536 27075 1576 27107
rect 1608 27075 1648 27107
rect 1680 27075 1720 27107
rect 1752 27075 1792 27107
rect 1824 27075 1864 27107
rect 1896 27075 1936 27107
rect 1968 27075 2008 27107
rect 2040 27075 2080 27107
rect 2112 27075 2152 27107
rect 2184 27075 2224 27107
rect 2256 27075 2296 27107
rect 2328 27075 2368 27107
rect 2400 27075 2440 27107
rect 2472 27075 2512 27107
rect 2544 27075 2584 27107
rect 2616 27075 2656 27107
rect 2688 27075 2728 27107
rect 2760 27075 2800 27107
rect 2832 27075 2872 27107
rect 2904 27075 2944 27107
rect 2976 27075 3016 27107
rect 3048 27075 3088 27107
rect 3120 27075 3160 27107
rect 3192 27075 3232 27107
rect 3264 27075 3304 27107
rect 3336 27075 3376 27107
rect 3408 27075 3448 27107
rect 3480 27075 3520 27107
rect 3552 27075 3592 27107
rect 3624 27075 3664 27107
rect 3696 27075 3736 27107
rect 3768 27075 3808 27107
rect 3840 27075 3880 27107
rect 3912 27075 3952 27107
rect 3984 27075 4024 27107
rect 4056 27075 4096 27107
rect 4128 27075 4168 27107
rect 4200 27075 4240 27107
rect 4272 27075 4312 27107
rect 4344 27075 4384 27107
rect 4416 27075 4456 27107
rect 4488 27075 4528 27107
rect 4560 27075 4600 27107
rect 4632 27075 4672 27107
rect 4704 27075 4744 27107
rect 4776 27075 4816 27107
rect 4848 27075 4888 27107
rect 4920 27075 4960 27107
rect 4992 27075 5032 27107
rect 5064 27075 5104 27107
rect 5136 27075 5176 27107
rect 5208 27075 5248 27107
rect 5280 27075 5320 27107
rect 5352 27075 5392 27107
rect 5424 27075 5464 27107
rect 5496 27075 5536 27107
rect 5568 27075 5608 27107
rect 5640 27075 5680 27107
rect 5712 27075 5752 27107
rect 5784 27075 5824 27107
rect 5856 27075 5896 27107
rect 5928 27075 5968 27107
rect 6000 27075 6040 27107
rect 6072 27075 6112 27107
rect 6144 27075 6184 27107
rect 6216 27075 6256 27107
rect 6288 27075 6328 27107
rect 6360 27075 6400 27107
rect 6432 27075 6472 27107
rect 6504 27075 6544 27107
rect 6576 27075 6616 27107
rect 6648 27075 6688 27107
rect 6720 27075 6760 27107
rect 6792 27075 6832 27107
rect 6864 27075 6904 27107
rect 6936 27075 6976 27107
rect 7008 27075 7048 27107
rect 7080 27075 7120 27107
rect 7152 27075 7192 27107
rect 7224 27075 7264 27107
rect 7296 27075 7336 27107
rect 7368 27075 7408 27107
rect 7440 27075 7480 27107
rect 7512 27075 7552 27107
rect 7584 27075 7624 27107
rect 7656 27075 7696 27107
rect 7728 27075 7768 27107
rect 7800 27075 7840 27107
rect 7872 27075 7912 27107
rect 7944 27075 7984 27107
rect 8016 27075 8056 27107
rect 8088 27075 8128 27107
rect 8160 27075 8200 27107
rect 8232 27075 8272 27107
rect 8304 27075 8344 27107
rect 8376 27075 8416 27107
rect 8448 27075 8488 27107
rect 8520 27075 8560 27107
rect 8592 27075 8632 27107
rect 8664 27075 8704 27107
rect 8736 27075 8776 27107
rect 8808 27075 8848 27107
rect 8880 27075 8920 27107
rect 8952 27075 8992 27107
rect 9024 27075 9064 27107
rect 9096 27075 9136 27107
rect 9168 27075 9208 27107
rect 9240 27075 9280 27107
rect 9312 27075 9352 27107
rect 9384 27075 9424 27107
rect 9456 27075 9496 27107
rect 9528 27075 9568 27107
rect 9600 27075 9640 27107
rect 9672 27075 9712 27107
rect 9744 27075 9784 27107
rect 9816 27075 9856 27107
rect 9888 27075 9928 27107
rect 9960 27075 10000 27107
rect 10032 27075 10072 27107
rect 10104 27075 10144 27107
rect 10176 27075 10216 27107
rect 10248 27075 10288 27107
rect 10320 27075 10360 27107
rect 10392 27075 10432 27107
rect 10464 27075 10504 27107
rect 10536 27075 10576 27107
rect 10608 27075 10648 27107
rect 10680 27075 10720 27107
rect 10752 27075 10792 27107
rect 10824 27075 10864 27107
rect 10896 27075 10936 27107
rect 10968 27075 11008 27107
rect 11040 27075 11080 27107
rect 11112 27075 11152 27107
rect 11184 27075 11224 27107
rect 11256 27075 11296 27107
rect 11328 27075 11368 27107
rect 11400 27075 11440 27107
rect 11472 27075 11512 27107
rect 11544 27075 11584 27107
rect 11616 27075 11656 27107
rect 11688 27075 11728 27107
rect 11760 27075 11800 27107
rect 11832 27075 11872 27107
rect 11904 27075 11944 27107
rect 11976 27075 12016 27107
rect 12048 27075 12088 27107
rect 12120 27075 12160 27107
rect 12192 27075 12232 27107
rect 12264 27075 12304 27107
rect 12336 27075 12376 27107
rect 12408 27075 12448 27107
rect 12480 27075 12520 27107
rect 12552 27075 12592 27107
rect 12624 27075 12664 27107
rect 12696 27075 12736 27107
rect 12768 27075 12808 27107
rect 12840 27075 12880 27107
rect 12912 27075 12952 27107
rect 12984 27075 13024 27107
rect 13056 27075 13096 27107
rect 13128 27075 13168 27107
rect 13200 27075 13240 27107
rect 13272 27075 13312 27107
rect 13344 27075 13384 27107
rect 13416 27075 13456 27107
rect 13488 27075 13528 27107
rect 13560 27075 13600 27107
rect 13632 27075 13672 27107
rect 13704 27075 13744 27107
rect 13776 27075 13816 27107
rect 13848 27075 13888 27107
rect 13920 27075 13960 27107
rect 13992 27075 14032 27107
rect 14064 27075 14104 27107
rect 14136 27075 14176 27107
rect 14208 27075 14248 27107
rect 14280 27075 14320 27107
rect 14352 27075 14392 27107
rect 14424 27075 14464 27107
rect 14496 27075 14536 27107
rect 14568 27075 14608 27107
rect 14640 27075 14680 27107
rect 14712 27075 14752 27107
rect 14784 27075 14824 27107
rect 14856 27075 14896 27107
rect 14928 27075 14968 27107
rect 15000 27075 15040 27107
rect 15072 27075 15112 27107
rect 15144 27075 15184 27107
rect 15216 27075 15256 27107
rect 15288 27075 15328 27107
rect 15360 27075 15400 27107
rect 15432 27075 15472 27107
rect 15504 27075 15544 27107
rect 15576 27075 15616 27107
rect 15648 27075 15688 27107
rect 15720 27075 15760 27107
rect 15792 27075 15832 27107
rect 15864 27075 15904 27107
rect 15936 27075 16000 27107
rect 0 27035 16000 27075
rect 0 27003 64 27035
rect 96 27003 136 27035
rect 168 27003 208 27035
rect 240 27003 280 27035
rect 312 27003 352 27035
rect 384 27003 424 27035
rect 456 27003 496 27035
rect 528 27003 568 27035
rect 600 27003 640 27035
rect 672 27003 712 27035
rect 744 27003 784 27035
rect 816 27003 856 27035
rect 888 27003 928 27035
rect 960 27003 1000 27035
rect 1032 27003 1072 27035
rect 1104 27003 1144 27035
rect 1176 27003 1216 27035
rect 1248 27003 1288 27035
rect 1320 27003 1360 27035
rect 1392 27003 1432 27035
rect 1464 27003 1504 27035
rect 1536 27003 1576 27035
rect 1608 27003 1648 27035
rect 1680 27003 1720 27035
rect 1752 27003 1792 27035
rect 1824 27003 1864 27035
rect 1896 27003 1936 27035
rect 1968 27003 2008 27035
rect 2040 27003 2080 27035
rect 2112 27003 2152 27035
rect 2184 27003 2224 27035
rect 2256 27003 2296 27035
rect 2328 27003 2368 27035
rect 2400 27003 2440 27035
rect 2472 27003 2512 27035
rect 2544 27003 2584 27035
rect 2616 27003 2656 27035
rect 2688 27003 2728 27035
rect 2760 27003 2800 27035
rect 2832 27003 2872 27035
rect 2904 27003 2944 27035
rect 2976 27003 3016 27035
rect 3048 27003 3088 27035
rect 3120 27003 3160 27035
rect 3192 27003 3232 27035
rect 3264 27003 3304 27035
rect 3336 27003 3376 27035
rect 3408 27003 3448 27035
rect 3480 27003 3520 27035
rect 3552 27003 3592 27035
rect 3624 27003 3664 27035
rect 3696 27003 3736 27035
rect 3768 27003 3808 27035
rect 3840 27003 3880 27035
rect 3912 27003 3952 27035
rect 3984 27003 4024 27035
rect 4056 27003 4096 27035
rect 4128 27003 4168 27035
rect 4200 27003 4240 27035
rect 4272 27003 4312 27035
rect 4344 27003 4384 27035
rect 4416 27003 4456 27035
rect 4488 27003 4528 27035
rect 4560 27003 4600 27035
rect 4632 27003 4672 27035
rect 4704 27003 4744 27035
rect 4776 27003 4816 27035
rect 4848 27003 4888 27035
rect 4920 27003 4960 27035
rect 4992 27003 5032 27035
rect 5064 27003 5104 27035
rect 5136 27003 5176 27035
rect 5208 27003 5248 27035
rect 5280 27003 5320 27035
rect 5352 27003 5392 27035
rect 5424 27003 5464 27035
rect 5496 27003 5536 27035
rect 5568 27003 5608 27035
rect 5640 27003 5680 27035
rect 5712 27003 5752 27035
rect 5784 27003 5824 27035
rect 5856 27003 5896 27035
rect 5928 27003 5968 27035
rect 6000 27003 6040 27035
rect 6072 27003 6112 27035
rect 6144 27003 6184 27035
rect 6216 27003 6256 27035
rect 6288 27003 6328 27035
rect 6360 27003 6400 27035
rect 6432 27003 6472 27035
rect 6504 27003 6544 27035
rect 6576 27003 6616 27035
rect 6648 27003 6688 27035
rect 6720 27003 6760 27035
rect 6792 27003 6832 27035
rect 6864 27003 6904 27035
rect 6936 27003 6976 27035
rect 7008 27003 7048 27035
rect 7080 27003 7120 27035
rect 7152 27003 7192 27035
rect 7224 27003 7264 27035
rect 7296 27003 7336 27035
rect 7368 27003 7408 27035
rect 7440 27003 7480 27035
rect 7512 27003 7552 27035
rect 7584 27003 7624 27035
rect 7656 27003 7696 27035
rect 7728 27003 7768 27035
rect 7800 27003 7840 27035
rect 7872 27003 7912 27035
rect 7944 27003 7984 27035
rect 8016 27003 8056 27035
rect 8088 27003 8128 27035
rect 8160 27003 8200 27035
rect 8232 27003 8272 27035
rect 8304 27003 8344 27035
rect 8376 27003 8416 27035
rect 8448 27003 8488 27035
rect 8520 27003 8560 27035
rect 8592 27003 8632 27035
rect 8664 27003 8704 27035
rect 8736 27003 8776 27035
rect 8808 27003 8848 27035
rect 8880 27003 8920 27035
rect 8952 27003 8992 27035
rect 9024 27003 9064 27035
rect 9096 27003 9136 27035
rect 9168 27003 9208 27035
rect 9240 27003 9280 27035
rect 9312 27003 9352 27035
rect 9384 27003 9424 27035
rect 9456 27003 9496 27035
rect 9528 27003 9568 27035
rect 9600 27003 9640 27035
rect 9672 27003 9712 27035
rect 9744 27003 9784 27035
rect 9816 27003 9856 27035
rect 9888 27003 9928 27035
rect 9960 27003 10000 27035
rect 10032 27003 10072 27035
rect 10104 27003 10144 27035
rect 10176 27003 10216 27035
rect 10248 27003 10288 27035
rect 10320 27003 10360 27035
rect 10392 27003 10432 27035
rect 10464 27003 10504 27035
rect 10536 27003 10576 27035
rect 10608 27003 10648 27035
rect 10680 27003 10720 27035
rect 10752 27003 10792 27035
rect 10824 27003 10864 27035
rect 10896 27003 10936 27035
rect 10968 27003 11008 27035
rect 11040 27003 11080 27035
rect 11112 27003 11152 27035
rect 11184 27003 11224 27035
rect 11256 27003 11296 27035
rect 11328 27003 11368 27035
rect 11400 27003 11440 27035
rect 11472 27003 11512 27035
rect 11544 27003 11584 27035
rect 11616 27003 11656 27035
rect 11688 27003 11728 27035
rect 11760 27003 11800 27035
rect 11832 27003 11872 27035
rect 11904 27003 11944 27035
rect 11976 27003 12016 27035
rect 12048 27003 12088 27035
rect 12120 27003 12160 27035
rect 12192 27003 12232 27035
rect 12264 27003 12304 27035
rect 12336 27003 12376 27035
rect 12408 27003 12448 27035
rect 12480 27003 12520 27035
rect 12552 27003 12592 27035
rect 12624 27003 12664 27035
rect 12696 27003 12736 27035
rect 12768 27003 12808 27035
rect 12840 27003 12880 27035
rect 12912 27003 12952 27035
rect 12984 27003 13024 27035
rect 13056 27003 13096 27035
rect 13128 27003 13168 27035
rect 13200 27003 13240 27035
rect 13272 27003 13312 27035
rect 13344 27003 13384 27035
rect 13416 27003 13456 27035
rect 13488 27003 13528 27035
rect 13560 27003 13600 27035
rect 13632 27003 13672 27035
rect 13704 27003 13744 27035
rect 13776 27003 13816 27035
rect 13848 27003 13888 27035
rect 13920 27003 13960 27035
rect 13992 27003 14032 27035
rect 14064 27003 14104 27035
rect 14136 27003 14176 27035
rect 14208 27003 14248 27035
rect 14280 27003 14320 27035
rect 14352 27003 14392 27035
rect 14424 27003 14464 27035
rect 14496 27003 14536 27035
rect 14568 27003 14608 27035
rect 14640 27003 14680 27035
rect 14712 27003 14752 27035
rect 14784 27003 14824 27035
rect 14856 27003 14896 27035
rect 14928 27003 14968 27035
rect 15000 27003 15040 27035
rect 15072 27003 15112 27035
rect 15144 27003 15184 27035
rect 15216 27003 15256 27035
rect 15288 27003 15328 27035
rect 15360 27003 15400 27035
rect 15432 27003 15472 27035
rect 15504 27003 15544 27035
rect 15576 27003 15616 27035
rect 15648 27003 15688 27035
rect 15720 27003 15760 27035
rect 15792 27003 15832 27035
rect 15864 27003 15904 27035
rect 15936 27003 16000 27035
rect 0 26963 16000 27003
rect 0 26931 64 26963
rect 96 26931 136 26963
rect 168 26931 208 26963
rect 240 26931 280 26963
rect 312 26931 352 26963
rect 384 26931 424 26963
rect 456 26931 496 26963
rect 528 26931 568 26963
rect 600 26931 640 26963
rect 672 26931 712 26963
rect 744 26931 784 26963
rect 816 26931 856 26963
rect 888 26931 928 26963
rect 960 26931 1000 26963
rect 1032 26931 1072 26963
rect 1104 26931 1144 26963
rect 1176 26931 1216 26963
rect 1248 26931 1288 26963
rect 1320 26931 1360 26963
rect 1392 26931 1432 26963
rect 1464 26931 1504 26963
rect 1536 26931 1576 26963
rect 1608 26931 1648 26963
rect 1680 26931 1720 26963
rect 1752 26931 1792 26963
rect 1824 26931 1864 26963
rect 1896 26931 1936 26963
rect 1968 26931 2008 26963
rect 2040 26931 2080 26963
rect 2112 26931 2152 26963
rect 2184 26931 2224 26963
rect 2256 26931 2296 26963
rect 2328 26931 2368 26963
rect 2400 26931 2440 26963
rect 2472 26931 2512 26963
rect 2544 26931 2584 26963
rect 2616 26931 2656 26963
rect 2688 26931 2728 26963
rect 2760 26931 2800 26963
rect 2832 26931 2872 26963
rect 2904 26931 2944 26963
rect 2976 26931 3016 26963
rect 3048 26931 3088 26963
rect 3120 26931 3160 26963
rect 3192 26931 3232 26963
rect 3264 26931 3304 26963
rect 3336 26931 3376 26963
rect 3408 26931 3448 26963
rect 3480 26931 3520 26963
rect 3552 26931 3592 26963
rect 3624 26931 3664 26963
rect 3696 26931 3736 26963
rect 3768 26931 3808 26963
rect 3840 26931 3880 26963
rect 3912 26931 3952 26963
rect 3984 26931 4024 26963
rect 4056 26931 4096 26963
rect 4128 26931 4168 26963
rect 4200 26931 4240 26963
rect 4272 26931 4312 26963
rect 4344 26931 4384 26963
rect 4416 26931 4456 26963
rect 4488 26931 4528 26963
rect 4560 26931 4600 26963
rect 4632 26931 4672 26963
rect 4704 26931 4744 26963
rect 4776 26931 4816 26963
rect 4848 26931 4888 26963
rect 4920 26931 4960 26963
rect 4992 26931 5032 26963
rect 5064 26931 5104 26963
rect 5136 26931 5176 26963
rect 5208 26931 5248 26963
rect 5280 26931 5320 26963
rect 5352 26931 5392 26963
rect 5424 26931 5464 26963
rect 5496 26931 5536 26963
rect 5568 26931 5608 26963
rect 5640 26931 5680 26963
rect 5712 26931 5752 26963
rect 5784 26931 5824 26963
rect 5856 26931 5896 26963
rect 5928 26931 5968 26963
rect 6000 26931 6040 26963
rect 6072 26931 6112 26963
rect 6144 26931 6184 26963
rect 6216 26931 6256 26963
rect 6288 26931 6328 26963
rect 6360 26931 6400 26963
rect 6432 26931 6472 26963
rect 6504 26931 6544 26963
rect 6576 26931 6616 26963
rect 6648 26931 6688 26963
rect 6720 26931 6760 26963
rect 6792 26931 6832 26963
rect 6864 26931 6904 26963
rect 6936 26931 6976 26963
rect 7008 26931 7048 26963
rect 7080 26931 7120 26963
rect 7152 26931 7192 26963
rect 7224 26931 7264 26963
rect 7296 26931 7336 26963
rect 7368 26931 7408 26963
rect 7440 26931 7480 26963
rect 7512 26931 7552 26963
rect 7584 26931 7624 26963
rect 7656 26931 7696 26963
rect 7728 26931 7768 26963
rect 7800 26931 7840 26963
rect 7872 26931 7912 26963
rect 7944 26931 7984 26963
rect 8016 26931 8056 26963
rect 8088 26931 8128 26963
rect 8160 26931 8200 26963
rect 8232 26931 8272 26963
rect 8304 26931 8344 26963
rect 8376 26931 8416 26963
rect 8448 26931 8488 26963
rect 8520 26931 8560 26963
rect 8592 26931 8632 26963
rect 8664 26931 8704 26963
rect 8736 26931 8776 26963
rect 8808 26931 8848 26963
rect 8880 26931 8920 26963
rect 8952 26931 8992 26963
rect 9024 26931 9064 26963
rect 9096 26931 9136 26963
rect 9168 26931 9208 26963
rect 9240 26931 9280 26963
rect 9312 26931 9352 26963
rect 9384 26931 9424 26963
rect 9456 26931 9496 26963
rect 9528 26931 9568 26963
rect 9600 26931 9640 26963
rect 9672 26931 9712 26963
rect 9744 26931 9784 26963
rect 9816 26931 9856 26963
rect 9888 26931 9928 26963
rect 9960 26931 10000 26963
rect 10032 26931 10072 26963
rect 10104 26931 10144 26963
rect 10176 26931 10216 26963
rect 10248 26931 10288 26963
rect 10320 26931 10360 26963
rect 10392 26931 10432 26963
rect 10464 26931 10504 26963
rect 10536 26931 10576 26963
rect 10608 26931 10648 26963
rect 10680 26931 10720 26963
rect 10752 26931 10792 26963
rect 10824 26931 10864 26963
rect 10896 26931 10936 26963
rect 10968 26931 11008 26963
rect 11040 26931 11080 26963
rect 11112 26931 11152 26963
rect 11184 26931 11224 26963
rect 11256 26931 11296 26963
rect 11328 26931 11368 26963
rect 11400 26931 11440 26963
rect 11472 26931 11512 26963
rect 11544 26931 11584 26963
rect 11616 26931 11656 26963
rect 11688 26931 11728 26963
rect 11760 26931 11800 26963
rect 11832 26931 11872 26963
rect 11904 26931 11944 26963
rect 11976 26931 12016 26963
rect 12048 26931 12088 26963
rect 12120 26931 12160 26963
rect 12192 26931 12232 26963
rect 12264 26931 12304 26963
rect 12336 26931 12376 26963
rect 12408 26931 12448 26963
rect 12480 26931 12520 26963
rect 12552 26931 12592 26963
rect 12624 26931 12664 26963
rect 12696 26931 12736 26963
rect 12768 26931 12808 26963
rect 12840 26931 12880 26963
rect 12912 26931 12952 26963
rect 12984 26931 13024 26963
rect 13056 26931 13096 26963
rect 13128 26931 13168 26963
rect 13200 26931 13240 26963
rect 13272 26931 13312 26963
rect 13344 26931 13384 26963
rect 13416 26931 13456 26963
rect 13488 26931 13528 26963
rect 13560 26931 13600 26963
rect 13632 26931 13672 26963
rect 13704 26931 13744 26963
rect 13776 26931 13816 26963
rect 13848 26931 13888 26963
rect 13920 26931 13960 26963
rect 13992 26931 14032 26963
rect 14064 26931 14104 26963
rect 14136 26931 14176 26963
rect 14208 26931 14248 26963
rect 14280 26931 14320 26963
rect 14352 26931 14392 26963
rect 14424 26931 14464 26963
rect 14496 26931 14536 26963
rect 14568 26931 14608 26963
rect 14640 26931 14680 26963
rect 14712 26931 14752 26963
rect 14784 26931 14824 26963
rect 14856 26931 14896 26963
rect 14928 26931 14968 26963
rect 15000 26931 15040 26963
rect 15072 26931 15112 26963
rect 15144 26931 15184 26963
rect 15216 26931 15256 26963
rect 15288 26931 15328 26963
rect 15360 26931 15400 26963
rect 15432 26931 15472 26963
rect 15504 26931 15544 26963
rect 15576 26931 15616 26963
rect 15648 26931 15688 26963
rect 15720 26931 15760 26963
rect 15792 26931 15832 26963
rect 15864 26931 15904 26963
rect 15936 26931 16000 26963
rect 0 26891 16000 26931
rect 0 26859 64 26891
rect 96 26859 136 26891
rect 168 26859 208 26891
rect 240 26859 280 26891
rect 312 26859 352 26891
rect 384 26859 424 26891
rect 456 26859 496 26891
rect 528 26859 568 26891
rect 600 26859 640 26891
rect 672 26859 712 26891
rect 744 26859 784 26891
rect 816 26859 856 26891
rect 888 26859 928 26891
rect 960 26859 1000 26891
rect 1032 26859 1072 26891
rect 1104 26859 1144 26891
rect 1176 26859 1216 26891
rect 1248 26859 1288 26891
rect 1320 26859 1360 26891
rect 1392 26859 1432 26891
rect 1464 26859 1504 26891
rect 1536 26859 1576 26891
rect 1608 26859 1648 26891
rect 1680 26859 1720 26891
rect 1752 26859 1792 26891
rect 1824 26859 1864 26891
rect 1896 26859 1936 26891
rect 1968 26859 2008 26891
rect 2040 26859 2080 26891
rect 2112 26859 2152 26891
rect 2184 26859 2224 26891
rect 2256 26859 2296 26891
rect 2328 26859 2368 26891
rect 2400 26859 2440 26891
rect 2472 26859 2512 26891
rect 2544 26859 2584 26891
rect 2616 26859 2656 26891
rect 2688 26859 2728 26891
rect 2760 26859 2800 26891
rect 2832 26859 2872 26891
rect 2904 26859 2944 26891
rect 2976 26859 3016 26891
rect 3048 26859 3088 26891
rect 3120 26859 3160 26891
rect 3192 26859 3232 26891
rect 3264 26859 3304 26891
rect 3336 26859 3376 26891
rect 3408 26859 3448 26891
rect 3480 26859 3520 26891
rect 3552 26859 3592 26891
rect 3624 26859 3664 26891
rect 3696 26859 3736 26891
rect 3768 26859 3808 26891
rect 3840 26859 3880 26891
rect 3912 26859 3952 26891
rect 3984 26859 4024 26891
rect 4056 26859 4096 26891
rect 4128 26859 4168 26891
rect 4200 26859 4240 26891
rect 4272 26859 4312 26891
rect 4344 26859 4384 26891
rect 4416 26859 4456 26891
rect 4488 26859 4528 26891
rect 4560 26859 4600 26891
rect 4632 26859 4672 26891
rect 4704 26859 4744 26891
rect 4776 26859 4816 26891
rect 4848 26859 4888 26891
rect 4920 26859 4960 26891
rect 4992 26859 5032 26891
rect 5064 26859 5104 26891
rect 5136 26859 5176 26891
rect 5208 26859 5248 26891
rect 5280 26859 5320 26891
rect 5352 26859 5392 26891
rect 5424 26859 5464 26891
rect 5496 26859 5536 26891
rect 5568 26859 5608 26891
rect 5640 26859 5680 26891
rect 5712 26859 5752 26891
rect 5784 26859 5824 26891
rect 5856 26859 5896 26891
rect 5928 26859 5968 26891
rect 6000 26859 6040 26891
rect 6072 26859 6112 26891
rect 6144 26859 6184 26891
rect 6216 26859 6256 26891
rect 6288 26859 6328 26891
rect 6360 26859 6400 26891
rect 6432 26859 6472 26891
rect 6504 26859 6544 26891
rect 6576 26859 6616 26891
rect 6648 26859 6688 26891
rect 6720 26859 6760 26891
rect 6792 26859 6832 26891
rect 6864 26859 6904 26891
rect 6936 26859 6976 26891
rect 7008 26859 7048 26891
rect 7080 26859 7120 26891
rect 7152 26859 7192 26891
rect 7224 26859 7264 26891
rect 7296 26859 7336 26891
rect 7368 26859 7408 26891
rect 7440 26859 7480 26891
rect 7512 26859 7552 26891
rect 7584 26859 7624 26891
rect 7656 26859 7696 26891
rect 7728 26859 7768 26891
rect 7800 26859 7840 26891
rect 7872 26859 7912 26891
rect 7944 26859 7984 26891
rect 8016 26859 8056 26891
rect 8088 26859 8128 26891
rect 8160 26859 8200 26891
rect 8232 26859 8272 26891
rect 8304 26859 8344 26891
rect 8376 26859 8416 26891
rect 8448 26859 8488 26891
rect 8520 26859 8560 26891
rect 8592 26859 8632 26891
rect 8664 26859 8704 26891
rect 8736 26859 8776 26891
rect 8808 26859 8848 26891
rect 8880 26859 8920 26891
rect 8952 26859 8992 26891
rect 9024 26859 9064 26891
rect 9096 26859 9136 26891
rect 9168 26859 9208 26891
rect 9240 26859 9280 26891
rect 9312 26859 9352 26891
rect 9384 26859 9424 26891
rect 9456 26859 9496 26891
rect 9528 26859 9568 26891
rect 9600 26859 9640 26891
rect 9672 26859 9712 26891
rect 9744 26859 9784 26891
rect 9816 26859 9856 26891
rect 9888 26859 9928 26891
rect 9960 26859 10000 26891
rect 10032 26859 10072 26891
rect 10104 26859 10144 26891
rect 10176 26859 10216 26891
rect 10248 26859 10288 26891
rect 10320 26859 10360 26891
rect 10392 26859 10432 26891
rect 10464 26859 10504 26891
rect 10536 26859 10576 26891
rect 10608 26859 10648 26891
rect 10680 26859 10720 26891
rect 10752 26859 10792 26891
rect 10824 26859 10864 26891
rect 10896 26859 10936 26891
rect 10968 26859 11008 26891
rect 11040 26859 11080 26891
rect 11112 26859 11152 26891
rect 11184 26859 11224 26891
rect 11256 26859 11296 26891
rect 11328 26859 11368 26891
rect 11400 26859 11440 26891
rect 11472 26859 11512 26891
rect 11544 26859 11584 26891
rect 11616 26859 11656 26891
rect 11688 26859 11728 26891
rect 11760 26859 11800 26891
rect 11832 26859 11872 26891
rect 11904 26859 11944 26891
rect 11976 26859 12016 26891
rect 12048 26859 12088 26891
rect 12120 26859 12160 26891
rect 12192 26859 12232 26891
rect 12264 26859 12304 26891
rect 12336 26859 12376 26891
rect 12408 26859 12448 26891
rect 12480 26859 12520 26891
rect 12552 26859 12592 26891
rect 12624 26859 12664 26891
rect 12696 26859 12736 26891
rect 12768 26859 12808 26891
rect 12840 26859 12880 26891
rect 12912 26859 12952 26891
rect 12984 26859 13024 26891
rect 13056 26859 13096 26891
rect 13128 26859 13168 26891
rect 13200 26859 13240 26891
rect 13272 26859 13312 26891
rect 13344 26859 13384 26891
rect 13416 26859 13456 26891
rect 13488 26859 13528 26891
rect 13560 26859 13600 26891
rect 13632 26859 13672 26891
rect 13704 26859 13744 26891
rect 13776 26859 13816 26891
rect 13848 26859 13888 26891
rect 13920 26859 13960 26891
rect 13992 26859 14032 26891
rect 14064 26859 14104 26891
rect 14136 26859 14176 26891
rect 14208 26859 14248 26891
rect 14280 26859 14320 26891
rect 14352 26859 14392 26891
rect 14424 26859 14464 26891
rect 14496 26859 14536 26891
rect 14568 26859 14608 26891
rect 14640 26859 14680 26891
rect 14712 26859 14752 26891
rect 14784 26859 14824 26891
rect 14856 26859 14896 26891
rect 14928 26859 14968 26891
rect 15000 26859 15040 26891
rect 15072 26859 15112 26891
rect 15144 26859 15184 26891
rect 15216 26859 15256 26891
rect 15288 26859 15328 26891
rect 15360 26859 15400 26891
rect 15432 26859 15472 26891
rect 15504 26859 15544 26891
rect 15576 26859 15616 26891
rect 15648 26859 15688 26891
rect 15720 26859 15760 26891
rect 15792 26859 15832 26891
rect 15864 26859 15904 26891
rect 15936 26859 16000 26891
rect 0 26819 16000 26859
rect 0 26787 64 26819
rect 96 26787 136 26819
rect 168 26787 208 26819
rect 240 26787 280 26819
rect 312 26787 352 26819
rect 384 26787 424 26819
rect 456 26787 496 26819
rect 528 26787 568 26819
rect 600 26787 640 26819
rect 672 26787 712 26819
rect 744 26787 784 26819
rect 816 26787 856 26819
rect 888 26787 928 26819
rect 960 26787 1000 26819
rect 1032 26787 1072 26819
rect 1104 26787 1144 26819
rect 1176 26787 1216 26819
rect 1248 26787 1288 26819
rect 1320 26787 1360 26819
rect 1392 26787 1432 26819
rect 1464 26787 1504 26819
rect 1536 26787 1576 26819
rect 1608 26787 1648 26819
rect 1680 26787 1720 26819
rect 1752 26787 1792 26819
rect 1824 26787 1864 26819
rect 1896 26787 1936 26819
rect 1968 26787 2008 26819
rect 2040 26787 2080 26819
rect 2112 26787 2152 26819
rect 2184 26787 2224 26819
rect 2256 26787 2296 26819
rect 2328 26787 2368 26819
rect 2400 26787 2440 26819
rect 2472 26787 2512 26819
rect 2544 26787 2584 26819
rect 2616 26787 2656 26819
rect 2688 26787 2728 26819
rect 2760 26787 2800 26819
rect 2832 26787 2872 26819
rect 2904 26787 2944 26819
rect 2976 26787 3016 26819
rect 3048 26787 3088 26819
rect 3120 26787 3160 26819
rect 3192 26787 3232 26819
rect 3264 26787 3304 26819
rect 3336 26787 3376 26819
rect 3408 26787 3448 26819
rect 3480 26787 3520 26819
rect 3552 26787 3592 26819
rect 3624 26787 3664 26819
rect 3696 26787 3736 26819
rect 3768 26787 3808 26819
rect 3840 26787 3880 26819
rect 3912 26787 3952 26819
rect 3984 26787 4024 26819
rect 4056 26787 4096 26819
rect 4128 26787 4168 26819
rect 4200 26787 4240 26819
rect 4272 26787 4312 26819
rect 4344 26787 4384 26819
rect 4416 26787 4456 26819
rect 4488 26787 4528 26819
rect 4560 26787 4600 26819
rect 4632 26787 4672 26819
rect 4704 26787 4744 26819
rect 4776 26787 4816 26819
rect 4848 26787 4888 26819
rect 4920 26787 4960 26819
rect 4992 26787 5032 26819
rect 5064 26787 5104 26819
rect 5136 26787 5176 26819
rect 5208 26787 5248 26819
rect 5280 26787 5320 26819
rect 5352 26787 5392 26819
rect 5424 26787 5464 26819
rect 5496 26787 5536 26819
rect 5568 26787 5608 26819
rect 5640 26787 5680 26819
rect 5712 26787 5752 26819
rect 5784 26787 5824 26819
rect 5856 26787 5896 26819
rect 5928 26787 5968 26819
rect 6000 26787 6040 26819
rect 6072 26787 6112 26819
rect 6144 26787 6184 26819
rect 6216 26787 6256 26819
rect 6288 26787 6328 26819
rect 6360 26787 6400 26819
rect 6432 26787 6472 26819
rect 6504 26787 6544 26819
rect 6576 26787 6616 26819
rect 6648 26787 6688 26819
rect 6720 26787 6760 26819
rect 6792 26787 6832 26819
rect 6864 26787 6904 26819
rect 6936 26787 6976 26819
rect 7008 26787 7048 26819
rect 7080 26787 7120 26819
rect 7152 26787 7192 26819
rect 7224 26787 7264 26819
rect 7296 26787 7336 26819
rect 7368 26787 7408 26819
rect 7440 26787 7480 26819
rect 7512 26787 7552 26819
rect 7584 26787 7624 26819
rect 7656 26787 7696 26819
rect 7728 26787 7768 26819
rect 7800 26787 7840 26819
rect 7872 26787 7912 26819
rect 7944 26787 7984 26819
rect 8016 26787 8056 26819
rect 8088 26787 8128 26819
rect 8160 26787 8200 26819
rect 8232 26787 8272 26819
rect 8304 26787 8344 26819
rect 8376 26787 8416 26819
rect 8448 26787 8488 26819
rect 8520 26787 8560 26819
rect 8592 26787 8632 26819
rect 8664 26787 8704 26819
rect 8736 26787 8776 26819
rect 8808 26787 8848 26819
rect 8880 26787 8920 26819
rect 8952 26787 8992 26819
rect 9024 26787 9064 26819
rect 9096 26787 9136 26819
rect 9168 26787 9208 26819
rect 9240 26787 9280 26819
rect 9312 26787 9352 26819
rect 9384 26787 9424 26819
rect 9456 26787 9496 26819
rect 9528 26787 9568 26819
rect 9600 26787 9640 26819
rect 9672 26787 9712 26819
rect 9744 26787 9784 26819
rect 9816 26787 9856 26819
rect 9888 26787 9928 26819
rect 9960 26787 10000 26819
rect 10032 26787 10072 26819
rect 10104 26787 10144 26819
rect 10176 26787 10216 26819
rect 10248 26787 10288 26819
rect 10320 26787 10360 26819
rect 10392 26787 10432 26819
rect 10464 26787 10504 26819
rect 10536 26787 10576 26819
rect 10608 26787 10648 26819
rect 10680 26787 10720 26819
rect 10752 26787 10792 26819
rect 10824 26787 10864 26819
rect 10896 26787 10936 26819
rect 10968 26787 11008 26819
rect 11040 26787 11080 26819
rect 11112 26787 11152 26819
rect 11184 26787 11224 26819
rect 11256 26787 11296 26819
rect 11328 26787 11368 26819
rect 11400 26787 11440 26819
rect 11472 26787 11512 26819
rect 11544 26787 11584 26819
rect 11616 26787 11656 26819
rect 11688 26787 11728 26819
rect 11760 26787 11800 26819
rect 11832 26787 11872 26819
rect 11904 26787 11944 26819
rect 11976 26787 12016 26819
rect 12048 26787 12088 26819
rect 12120 26787 12160 26819
rect 12192 26787 12232 26819
rect 12264 26787 12304 26819
rect 12336 26787 12376 26819
rect 12408 26787 12448 26819
rect 12480 26787 12520 26819
rect 12552 26787 12592 26819
rect 12624 26787 12664 26819
rect 12696 26787 12736 26819
rect 12768 26787 12808 26819
rect 12840 26787 12880 26819
rect 12912 26787 12952 26819
rect 12984 26787 13024 26819
rect 13056 26787 13096 26819
rect 13128 26787 13168 26819
rect 13200 26787 13240 26819
rect 13272 26787 13312 26819
rect 13344 26787 13384 26819
rect 13416 26787 13456 26819
rect 13488 26787 13528 26819
rect 13560 26787 13600 26819
rect 13632 26787 13672 26819
rect 13704 26787 13744 26819
rect 13776 26787 13816 26819
rect 13848 26787 13888 26819
rect 13920 26787 13960 26819
rect 13992 26787 14032 26819
rect 14064 26787 14104 26819
rect 14136 26787 14176 26819
rect 14208 26787 14248 26819
rect 14280 26787 14320 26819
rect 14352 26787 14392 26819
rect 14424 26787 14464 26819
rect 14496 26787 14536 26819
rect 14568 26787 14608 26819
rect 14640 26787 14680 26819
rect 14712 26787 14752 26819
rect 14784 26787 14824 26819
rect 14856 26787 14896 26819
rect 14928 26787 14968 26819
rect 15000 26787 15040 26819
rect 15072 26787 15112 26819
rect 15144 26787 15184 26819
rect 15216 26787 15256 26819
rect 15288 26787 15328 26819
rect 15360 26787 15400 26819
rect 15432 26787 15472 26819
rect 15504 26787 15544 26819
rect 15576 26787 15616 26819
rect 15648 26787 15688 26819
rect 15720 26787 15760 26819
rect 15792 26787 15832 26819
rect 15864 26787 15904 26819
rect 15936 26787 16000 26819
rect 0 26755 16000 26787
rect 0 26715 51 26755
rect 91 26747 149 26755
rect 189 26747 247 26755
rect 287 26747 345 26755
rect 385 26747 443 26755
rect 483 26747 541 26755
rect 581 26747 639 26755
rect 679 26747 737 26755
rect 777 26747 835 26755
rect 875 26747 933 26755
rect 973 26747 1031 26755
rect 1071 26747 1129 26755
rect 1169 26747 16000 26755
rect 96 26715 136 26747
rect 189 26715 208 26747
rect 240 26715 247 26747
rect 312 26715 345 26747
rect 385 26715 424 26747
rect 483 26715 496 26747
rect 528 26715 541 26747
rect 600 26715 639 26747
rect 679 26715 712 26747
rect 777 26715 784 26747
rect 816 26715 835 26747
rect 888 26715 928 26747
rect 973 26715 1000 26747
rect 1071 26715 1072 26747
rect 1104 26715 1129 26747
rect 1176 26715 1216 26747
rect 1248 26715 1288 26747
rect 1320 26715 1360 26747
rect 1392 26715 1432 26747
rect 1464 26715 1504 26747
rect 1536 26715 1576 26747
rect 1608 26715 1648 26747
rect 1680 26715 1720 26747
rect 1752 26715 1792 26747
rect 1824 26715 1864 26747
rect 1896 26715 1936 26747
rect 1968 26715 2008 26747
rect 2040 26715 2080 26747
rect 2112 26715 2152 26747
rect 2184 26715 2224 26747
rect 2256 26715 2296 26747
rect 2328 26715 2368 26747
rect 2400 26715 2440 26747
rect 2472 26715 2512 26747
rect 2544 26715 2584 26747
rect 2616 26715 2656 26747
rect 2688 26715 2728 26747
rect 2760 26715 2800 26747
rect 2832 26715 2872 26747
rect 2904 26715 2944 26747
rect 2976 26715 3016 26747
rect 3048 26715 3088 26747
rect 3120 26715 3160 26747
rect 3192 26715 3232 26747
rect 3264 26715 3304 26747
rect 3336 26715 3376 26747
rect 3408 26715 3448 26747
rect 3480 26715 3520 26747
rect 3552 26715 3592 26747
rect 3624 26715 3664 26747
rect 3696 26715 3736 26747
rect 3768 26715 3808 26747
rect 3840 26715 3880 26747
rect 3912 26715 3952 26747
rect 3984 26715 4024 26747
rect 4056 26715 4096 26747
rect 4128 26715 4168 26747
rect 4200 26715 4240 26747
rect 4272 26715 4312 26747
rect 4344 26715 4384 26747
rect 4416 26715 4456 26747
rect 4488 26715 4528 26747
rect 4560 26715 4600 26747
rect 4632 26715 4672 26747
rect 4704 26715 4744 26747
rect 4776 26715 4816 26747
rect 4848 26715 4888 26747
rect 4920 26715 4960 26747
rect 4992 26715 5032 26747
rect 5064 26715 5104 26747
rect 5136 26715 5176 26747
rect 5208 26715 5248 26747
rect 5280 26715 5320 26747
rect 5352 26715 5392 26747
rect 5424 26715 5464 26747
rect 5496 26715 5536 26747
rect 5568 26715 5608 26747
rect 5640 26715 5680 26747
rect 5712 26715 5752 26747
rect 5784 26715 5824 26747
rect 5856 26715 5896 26747
rect 5928 26715 5968 26747
rect 6000 26715 6040 26747
rect 6072 26715 6112 26747
rect 6144 26715 6184 26747
rect 6216 26715 6256 26747
rect 6288 26715 6328 26747
rect 6360 26715 6400 26747
rect 6432 26715 6472 26747
rect 6504 26715 6544 26747
rect 6576 26715 6616 26747
rect 6648 26715 6688 26747
rect 6720 26715 6760 26747
rect 6792 26715 6832 26747
rect 6864 26715 6904 26747
rect 6936 26715 6976 26747
rect 7008 26715 7048 26747
rect 7080 26715 7120 26747
rect 7152 26715 7192 26747
rect 7224 26715 7264 26747
rect 7296 26715 7336 26747
rect 7368 26715 7408 26747
rect 7440 26715 7480 26747
rect 7512 26715 7552 26747
rect 7584 26715 7624 26747
rect 7656 26715 7696 26747
rect 7728 26715 7768 26747
rect 7800 26715 7840 26747
rect 7872 26715 7912 26747
rect 7944 26715 7984 26747
rect 8016 26715 8056 26747
rect 8088 26715 8128 26747
rect 8160 26715 8200 26747
rect 8232 26715 8272 26747
rect 8304 26715 8344 26747
rect 8376 26715 8416 26747
rect 8448 26715 8488 26747
rect 8520 26715 8560 26747
rect 8592 26715 8632 26747
rect 8664 26715 8704 26747
rect 8736 26715 8776 26747
rect 8808 26715 8848 26747
rect 8880 26715 8920 26747
rect 8952 26715 8992 26747
rect 9024 26715 9064 26747
rect 9096 26715 9136 26747
rect 9168 26715 9208 26747
rect 9240 26715 9280 26747
rect 9312 26715 9352 26747
rect 9384 26715 9424 26747
rect 9456 26715 9496 26747
rect 9528 26715 9568 26747
rect 9600 26715 9640 26747
rect 9672 26715 9712 26747
rect 9744 26715 9784 26747
rect 9816 26715 9856 26747
rect 9888 26715 9928 26747
rect 9960 26715 10000 26747
rect 10032 26715 10072 26747
rect 10104 26715 10144 26747
rect 10176 26715 10216 26747
rect 10248 26715 10288 26747
rect 10320 26715 10360 26747
rect 10392 26715 10432 26747
rect 10464 26715 10504 26747
rect 10536 26715 10576 26747
rect 10608 26715 10648 26747
rect 10680 26715 10720 26747
rect 10752 26715 10792 26747
rect 10824 26715 10864 26747
rect 10896 26715 10936 26747
rect 10968 26715 11008 26747
rect 11040 26715 11080 26747
rect 11112 26715 11152 26747
rect 11184 26715 11224 26747
rect 11256 26715 11296 26747
rect 11328 26715 11368 26747
rect 11400 26715 11440 26747
rect 11472 26715 11512 26747
rect 11544 26715 11584 26747
rect 11616 26715 11656 26747
rect 11688 26715 11728 26747
rect 11760 26715 11800 26747
rect 11832 26715 11872 26747
rect 11904 26715 11944 26747
rect 11976 26715 12016 26747
rect 12048 26715 12088 26747
rect 12120 26715 12160 26747
rect 12192 26715 12232 26747
rect 12264 26715 12304 26747
rect 12336 26715 12376 26747
rect 12408 26715 12448 26747
rect 12480 26715 12520 26747
rect 12552 26715 12592 26747
rect 12624 26715 12664 26747
rect 12696 26715 12736 26747
rect 12768 26715 12808 26747
rect 12840 26715 12880 26747
rect 12912 26715 12952 26747
rect 12984 26715 13024 26747
rect 13056 26715 13096 26747
rect 13128 26715 13168 26747
rect 13200 26715 13240 26747
rect 13272 26715 13312 26747
rect 13344 26715 13384 26747
rect 13416 26715 13456 26747
rect 13488 26715 13528 26747
rect 13560 26715 13600 26747
rect 13632 26715 13672 26747
rect 13704 26715 13744 26747
rect 13776 26715 13816 26747
rect 13848 26715 13888 26747
rect 13920 26715 13960 26747
rect 13992 26715 14032 26747
rect 14064 26715 14104 26747
rect 14136 26715 14176 26747
rect 14208 26715 14248 26747
rect 14280 26715 14320 26747
rect 14352 26715 14392 26747
rect 14424 26715 14464 26747
rect 14496 26715 14536 26747
rect 14568 26715 14608 26747
rect 14640 26715 14680 26747
rect 14712 26715 14752 26747
rect 14784 26715 14824 26747
rect 14856 26715 14896 26747
rect 14928 26715 14968 26747
rect 15000 26715 15040 26747
rect 15072 26715 15112 26747
rect 15144 26715 15184 26747
rect 15216 26715 15256 26747
rect 15288 26715 15328 26747
rect 15360 26715 15400 26747
rect 15432 26715 15472 26747
rect 15504 26715 15544 26747
rect 15576 26715 15616 26747
rect 15648 26715 15688 26747
rect 15720 26715 15760 26747
rect 15792 26715 15832 26747
rect 15864 26715 15904 26747
rect 15936 26715 16000 26747
rect 0 26675 16000 26715
rect 0 26657 64 26675
rect 0 26617 51 26657
rect 96 26643 136 26675
rect 168 26657 208 26675
rect 189 26643 208 26657
rect 240 26657 280 26675
rect 312 26657 352 26675
rect 384 26657 424 26675
rect 456 26657 496 26675
rect 240 26643 247 26657
rect 312 26643 345 26657
rect 385 26643 424 26657
rect 483 26643 496 26657
rect 528 26657 568 26675
rect 600 26657 640 26675
rect 672 26657 712 26675
rect 744 26657 784 26675
rect 528 26643 541 26657
rect 600 26643 639 26657
rect 679 26643 712 26657
rect 777 26643 784 26657
rect 816 26657 856 26675
rect 816 26643 835 26657
rect 888 26643 928 26675
rect 960 26657 1000 26675
rect 1032 26657 1072 26675
rect 973 26643 1000 26657
rect 1071 26643 1072 26657
rect 1104 26657 1144 26675
rect 1104 26643 1129 26657
rect 1176 26643 1216 26675
rect 1248 26643 1288 26675
rect 1320 26643 1360 26675
rect 1392 26643 1432 26675
rect 1464 26643 1504 26675
rect 1536 26643 1576 26675
rect 1608 26643 1648 26675
rect 1680 26643 1720 26675
rect 1752 26643 1792 26675
rect 1824 26643 1864 26675
rect 1896 26643 1936 26675
rect 1968 26643 2008 26675
rect 2040 26643 2080 26675
rect 2112 26643 2152 26675
rect 2184 26643 2224 26675
rect 2256 26643 2296 26675
rect 2328 26643 2368 26675
rect 2400 26643 2440 26675
rect 2472 26643 2512 26675
rect 2544 26643 2584 26675
rect 2616 26643 2656 26675
rect 2688 26643 2728 26675
rect 2760 26643 2800 26675
rect 2832 26643 2872 26675
rect 2904 26643 2944 26675
rect 2976 26643 3016 26675
rect 3048 26643 3088 26675
rect 3120 26643 3160 26675
rect 3192 26643 3232 26675
rect 3264 26643 3304 26675
rect 3336 26643 3376 26675
rect 3408 26643 3448 26675
rect 3480 26643 3520 26675
rect 3552 26643 3592 26675
rect 3624 26643 3664 26675
rect 3696 26643 3736 26675
rect 3768 26643 3808 26675
rect 3840 26643 3880 26675
rect 3912 26643 3952 26675
rect 3984 26643 4024 26675
rect 4056 26643 4096 26675
rect 4128 26643 4168 26675
rect 4200 26643 4240 26675
rect 4272 26643 4312 26675
rect 4344 26643 4384 26675
rect 4416 26643 4456 26675
rect 4488 26643 4528 26675
rect 4560 26643 4600 26675
rect 4632 26643 4672 26675
rect 4704 26643 4744 26675
rect 4776 26643 4816 26675
rect 4848 26643 4888 26675
rect 4920 26643 4960 26675
rect 4992 26643 5032 26675
rect 5064 26643 5104 26675
rect 5136 26643 5176 26675
rect 5208 26643 5248 26675
rect 5280 26643 5320 26675
rect 5352 26643 5392 26675
rect 5424 26643 5464 26675
rect 5496 26643 5536 26675
rect 5568 26643 5608 26675
rect 5640 26643 5680 26675
rect 5712 26643 5752 26675
rect 5784 26643 5824 26675
rect 5856 26643 5896 26675
rect 5928 26643 5968 26675
rect 6000 26643 6040 26675
rect 6072 26643 6112 26675
rect 6144 26643 6184 26675
rect 6216 26643 6256 26675
rect 6288 26643 6328 26675
rect 6360 26643 6400 26675
rect 6432 26643 6472 26675
rect 6504 26643 6544 26675
rect 6576 26643 6616 26675
rect 6648 26643 6688 26675
rect 6720 26643 6760 26675
rect 6792 26643 6832 26675
rect 6864 26643 6904 26675
rect 6936 26643 6976 26675
rect 7008 26643 7048 26675
rect 7080 26643 7120 26675
rect 7152 26643 7192 26675
rect 7224 26643 7264 26675
rect 7296 26643 7336 26675
rect 7368 26643 7408 26675
rect 7440 26643 7480 26675
rect 7512 26643 7552 26675
rect 7584 26643 7624 26675
rect 7656 26643 7696 26675
rect 7728 26643 7768 26675
rect 7800 26643 7840 26675
rect 7872 26643 7912 26675
rect 7944 26643 7984 26675
rect 8016 26643 8056 26675
rect 8088 26643 8128 26675
rect 8160 26643 8200 26675
rect 8232 26643 8272 26675
rect 8304 26643 8344 26675
rect 8376 26643 8416 26675
rect 8448 26643 8488 26675
rect 8520 26643 8560 26675
rect 8592 26643 8632 26675
rect 8664 26643 8704 26675
rect 8736 26643 8776 26675
rect 8808 26643 8848 26675
rect 8880 26643 8920 26675
rect 8952 26643 8992 26675
rect 9024 26643 9064 26675
rect 9096 26643 9136 26675
rect 9168 26643 9208 26675
rect 9240 26643 9280 26675
rect 9312 26643 9352 26675
rect 9384 26643 9424 26675
rect 9456 26643 9496 26675
rect 9528 26643 9568 26675
rect 9600 26643 9640 26675
rect 9672 26643 9712 26675
rect 9744 26643 9784 26675
rect 9816 26643 9856 26675
rect 9888 26643 9928 26675
rect 9960 26643 10000 26675
rect 10032 26643 10072 26675
rect 10104 26643 10144 26675
rect 10176 26643 10216 26675
rect 10248 26643 10288 26675
rect 10320 26643 10360 26675
rect 10392 26643 10432 26675
rect 10464 26643 10504 26675
rect 10536 26643 10576 26675
rect 10608 26643 10648 26675
rect 10680 26643 10720 26675
rect 10752 26643 10792 26675
rect 10824 26643 10864 26675
rect 10896 26643 10936 26675
rect 10968 26643 11008 26675
rect 11040 26643 11080 26675
rect 11112 26643 11152 26675
rect 11184 26643 11224 26675
rect 11256 26643 11296 26675
rect 11328 26643 11368 26675
rect 11400 26643 11440 26675
rect 11472 26643 11512 26675
rect 11544 26643 11584 26675
rect 11616 26643 11656 26675
rect 11688 26643 11728 26675
rect 11760 26643 11800 26675
rect 11832 26643 11872 26675
rect 11904 26643 11944 26675
rect 11976 26643 12016 26675
rect 12048 26643 12088 26675
rect 12120 26643 12160 26675
rect 12192 26643 12232 26675
rect 12264 26643 12304 26675
rect 12336 26643 12376 26675
rect 12408 26643 12448 26675
rect 12480 26643 12520 26675
rect 12552 26643 12592 26675
rect 12624 26643 12664 26675
rect 12696 26643 12736 26675
rect 12768 26643 12808 26675
rect 12840 26643 12880 26675
rect 12912 26643 12952 26675
rect 12984 26643 13024 26675
rect 13056 26643 13096 26675
rect 13128 26643 13168 26675
rect 13200 26643 13240 26675
rect 13272 26643 13312 26675
rect 13344 26643 13384 26675
rect 13416 26643 13456 26675
rect 13488 26643 13528 26675
rect 13560 26643 13600 26675
rect 13632 26643 13672 26675
rect 13704 26643 13744 26675
rect 13776 26643 13816 26675
rect 13848 26643 13888 26675
rect 13920 26643 13960 26675
rect 13992 26643 14032 26675
rect 14064 26643 14104 26675
rect 14136 26643 14176 26675
rect 14208 26643 14248 26675
rect 14280 26643 14320 26675
rect 14352 26643 14392 26675
rect 14424 26643 14464 26675
rect 14496 26643 14536 26675
rect 14568 26643 14608 26675
rect 14640 26643 14680 26675
rect 14712 26643 14752 26675
rect 14784 26643 14824 26675
rect 14856 26643 14896 26675
rect 14928 26643 14968 26675
rect 15000 26643 15040 26675
rect 15072 26643 15112 26675
rect 15144 26643 15184 26675
rect 15216 26643 15256 26675
rect 15288 26643 15328 26675
rect 15360 26643 15400 26675
rect 15432 26643 15472 26675
rect 15504 26643 15544 26675
rect 15576 26643 15616 26675
rect 15648 26643 15688 26675
rect 15720 26643 15760 26675
rect 15792 26643 15832 26675
rect 15864 26643 15904 26675
rect 15936 26643 16000 26675
rect 91 26617 149 26643
rect 189 26617 247 26643
rect 287 26617 345 26643
rect 385 26617 443 26643
rect 483 26617 541 26643
rect 581 26617 639 26643
rect 679 26617 737 26643
rect 777 26617 835 26643
rect 875 26617 933 26643
rect 973 26617 1031 26643
rect 1071 26617 1129 26643
rect 1169 26617 16000 26643
rect 0 26603 16000 26617
rect 0 26571 64 26603
rect 96 26571 136 26603
rect 168 26571 208 26603
rect 240 26571 280 26603
rect 312 26571 352 26603
rect 384 26571 424 26603
rect 456 26571 496 26603
rect 528 26571 568 26603
rect 600 26571 640 26603
rect 672 26571 712 26603
rect 744 26571 784 26603
rect 816 26571 856 26603
rect 888 26571 928 26603
rect 960 26571 1000 26603
rect 1032 26571 1072 26603
rect 1104 26571 1144 26603
rect 1176 26571 1216 26603
rect 1248 26571 1288 26603
rect 1320 26571 1360 26603
rect 1392 26571 1432 26603
rect 1464 26571 1504 26603
rect 1536 26571 1576 26603
rect 1608 26571 1648 26603
rect 1680 26571 1720 26603
rect 1752 26571 1792 26603
rect 1824 26571 1864 26603
rect 1896 26571 1936 26603
rect 1968 26571 2008 26603
rect 2040 26571 2080 26603
rect 2112 26571 2152 26603
rect 2184 26571 2224 26603
rect 2256 26571 2296 26603
rect 2328 26571 2368 26603
rect 2400 26571 2440 26603
rect 2472 26571 2512 26603
rect 2544 26571 2584 26603
rect 2616 26571 2656 26603
rect 2688 26571 2728 26603
rect 2760 26571 2800 26603
rect 2832 26571 2872 26603
rect 2904 26571 2944 26603
rect 2976 26571 3016 26603
rect 3048 26571 3088 26603
rect 3120 26571 3160 26603
rect 3192 26571 3232 26603
rect 3264 26571 3304 26603
rect 3336 26571 3376 26603
rect 3408 26571 3448 26603
rect 3480 26571 3520 26603
rect 3552 26571 3592 26603
rect 3624 26571 3664 26603
rect 3696 26571 3736 26603
rect 3768 26571 3808 26603
rect 3840 26571 3880 26603
rect 3912 26571 3952 26603
rect 3984 26571 4024 26603
rect 4056 26571 4096 26603
rect 4128 26571 4168 26603
rect 4200 26571 4240 26603
rect 4272 26571 4312 26603
rect 4344 26571 4384 26603
rect 4416 26571 4456 26603
rect 4488 26571 4528 26603
rect 4560 26571 4600 26603
rect 4632 26571 4672 26603
rect 4704 26571 4744 26603
rect 4776 26571 4816 26603
rect 4848 26571 4888 26603
rect 4920 26571 4960 26603
rect 4992 26571 5032 26603
rect 5064 26571 5104 26603
rect 5136 26571 5176 26603
rect 5208 26571 5248 26603
rect 5280 26571 5320 26603
rect 5352 26571 5392 26603
rect 5424 26571 5464 26603
rect 5496 26571 5536 26603
rect 5568 26571 5608 26603
rect 5640 26571 5680 26603
rect 5712 26571 5752 26603
rect 5784 26571 5824 26603
rect 5856 26571 5896 26603
rect 5928 26571 5968 26603
rect 6000 26571 6040 26603
rect 6072 26571 6112 26603
rect 6144 26571 6184 26603
rect 6216 26571 6256 26603
rect 6288 26571 6328 26603
rect 6360 26571 6400 26603
rect 6432 26571 6472 26603
rect 6504 26571 6544 26603
rect 6576 26571 6616 26603
rect 6648 26571 6688 26603
rect 6720 26571 6760 26603
rect 6792 26571 6832 26603
rect 6864 26571 6904 26603
rect 6936 26571 6976 26603
rect 7008 26571 7048 26603
rect 7080 26571 7120 26603
rect 7152 26571 7192 26603
rect 7224 26571 7264 26603
rect 7296 26571 7336 26603
rect 7368 26571 7408 26603
rect 7440 26571 7480 26603
rect 7512 26571 7552 26603
rect 7584 26571 7624 26603
rect 7656 26571 7696 26603
rect 7728 26571 7768 26603
rect 7800 26571 7840 26603
rect 7872 26571 7912 26603
rect 7944 26571 7984 26603
rect 8016 26571 8056 26603
rect 8088 26571 8128 26603
rect 8160 26571 8200 26603
rect 8232 26571 8272 26603
rect 8304 26571 8344 26603
rect 8376 26571 8416 26603
rect 8448 26571 8488 26603
rect 8520 26571 8560 26603
rect 8592 26571 8632 26603
rect 8664 26571 8704 26603
rect 8736 26571 8776 26603
rect 8808 26571 8848 26603
rect 8880 26571 8920 26603
rect 8952 26571 8992 26603
rect 9024 26571 9064 26603
rect 9096 26571 9136 26603
rect 9168 26571 9208 26603
rect 9240 26571 9280 26603
rect 9312 26571 9352 26603
rect 9384 26571 9424 26603
rect 9456 26571 9496 26603
rect 9528 26571 9568 26603
rect 9600 26571 9640 26603
rect 9672 26571 9712 26603
rect 9744 26571 9784 26603
rect 9816 26571 9856 26603
rect 9888 26571 9928 26603
rect 9960 26571 10000 26603
rect 10032 26571 10072 26603
rect 10104 26571 10144 26603
rect 10176 26571 10216 26603
rect 10248 26571 10288 26603
rect 10320 26571 10360 26603
rect 10392 26571 10432 26603
rect 10464 26571 10504 26603
rect 10536 26571 10576 26603
rect 10608 26571 10648 26603
rect 10680 26571 10720 26603
rect 10752 26571 10792 26603
rect 10824 26571 10864 26603
rect 10896 26571 10936 26603
rect 10968 26571 11008 26603
rect 11040 26571 11080 26603
rect 11112 26571 11152 26603
rect 11184 26571 11224 26603
rect 11256 26571 11296 26603
rect 11328 26571 11368 26603
rect 11400 26571 11440 26603
rect 11472 26571 11512 26603
rect 11544 26571 11584 26603
rect 11616 26571 11656 26603
rect 11688 26571 11728 26603
rect 11760 26571 11800 26603
rect 11832 26571 11872 26603
rect 11904 26571 11944 26603
rect 11976 26571 12016 26603
rect 12048 26571 12088 26603
rect 12120 26571 12160 26603
rect 12192 26571 12232 26603
rect 12264 26571 12304 26603
rect 12336 26571 12376 26603
rect 12408 26571 12448 26603
rect 12480 26571 12520 26603
rect 12552 26571 12592 26603
rect 12624 26571 12664 26603
rect 12696 26571 12736 26603
rect 12768 26571 12808 26603
rect 12840 26571 12880 26603
rect 12912 26571 12952 26603
rect 12984 26571 13024 26603
rect 13056 26571 13096 26603
rect 13128 26571 13168 26603
rect 13200 26571 13240 26603
rect 13272 26571 13312 26603
rect 13344 26571 13384 26603
rect 13416 26571 13456 26603
rect 13488 26571 13528 26603
rect 13560 26571 13600 26603
rect 13632 26571 13672 26603
rect 13704 26571 13744 26603
rect 13776 26571 13816 26603
rect 13848 26571 13888 26603
rect 13920 26571 13960 26603
rect 13992 26571 14032 26603
rect 14064 26571 14104 26603
rect 14136 26571 14176 26603
rect 14208 26571 14248 26603
rect 14280 26571 14320 26603
rect 14352 26571 14392 26603
rect 14424 26571 14464 26603
rect 14496 26571 14536 26603
rect 14568 26571 14608 26603
rect 14640 26571 14680 26603
rect 14712 26571 14752 26603
rect 14784 26571 14824 26603
rect 14856 26571 14896 26603
rect 14928 26571 14968 26603
rect 15000 26571 15040 26603
rect 15072 26571 15112 26603
rect 15144 26571 15184 26603
rect 15216 26571 15256 26603
rect 15288 26571 15328 26603
rect 15360 26571 15400 26603
rect 15432 26571 15472 26603
rect 15504 26571 15544 26603
rect 15576 26571 15616 26603
rect 15648 26571 15688 26603
rect 15720 26571 15760 26603
rect 15792 26571 15832 26603
rect 15864 26571 15904 26603
rect 15936 26571 16000 26603
rect 0 26559 16000 26571
rect 0 26519 51 26559
rect 91 26531 149 26559
rect 189 26531 247 26559
rect 287 26531 345 26559
rect 385 26531 443 26559
rect 483 26531 541 26559
rect 581 26531 639 26559
rect 679 26531 737 26559
rect 777 26531 835 26559
rect 875 26531 933 26559
rect 973 26531 1031 26559
rect 1071 26531 1129 26559
rect 1169 26531 16000 26559
rect 0 26499 64 26519
rect 96 26499 136 26531
rect 189 26519 208 26531
rect 168 26499 208 26519
rect 240 26519 247 26531
rect 312 26519 345 26531
rect 385 26519 424 26531
rect 483 26519 496 26531
rect 240 26499 280 26519
rect 312 26499 352 26519
rect 384 26499 424 26519
rect 456 26499 496 26519
rect 528 26519 541 26531
rect 600 26519 639 26531
rect 679 26519 712 26531
rect 777 26519 784 26531
rect 528 26499 568 26519
rect 600 26499 640 26519
rect 672 26499 712 26519
rect 744 26499 784 26519
rect 816 26519 835 26531
rect 816 26499 856 26519
rect 888 26499 928 26531
rect 973 26519 1000 26531
rect 1071 26519 1072 26531
rect 960 26499 1000 26519
rect 1032 26499 1072 26519
rect 1104 26519 1129 26531
rect 1104 26499 1144 26519
rect 1176 26499 1216 26531
rect 1248 26499 1288 26531
rect 1320 26499 1360 26531
rect 1392 26499 1432 26531
rect 1464 26499 1504 26531
rect 1536 26499 1576 26531
rect 1608 26499 1648 26531
rect 1680 26499 1720 26531
rect 1752 26499 1792 26531
rect 1824 26499 1864 26531
rect 1896 26499 1936 26531
rect 1968 26499 2008 26531
rect 2040 26499 2080 26531
rect 2112 26499 2152 26531
rect 2184 26499 2224 26531
rect 2256 26499 2296 26531
rect 2328 26499 2368 26531
rect 2400 26499 2440 26531
rect 2472 26499 2512 26531
rect 2544 26499 2584 26531
rect 2616 26499 2656 26531
rect 2688 26499 2728 26531
rect 2760 26499 2800 26531
rect 2832 26499 2872 26531
rect 2904 26499 2944 26531
rect 2976 26499 3016 26531
rect 3048 26499 3088 26531
rect 3120 26499 3160 26531
rect 3192 26499 3232 26531
rect 3264 26499 3304 26531
rect 3336 26499 3376 26531
rect 3408 26499 3448 26531
rect 3480 26499 3520 26531
rect 3552 26499 3592 26531
rect 3624 26499 3664 26531
rect 3696 26499 3736 26531
rect 3768 26499 3808 26531
rect 3840 26499 3880 26531
rect 3912 26499 3952 26531
rect 3984 26499 4024 26531
rect 4056 26499 4096 26531
rect 4128 26499 4168 26531
rect 4200 26499 4240 26531
rect 4272 26499 4312 26531
rect 4344 26499 4384 26531
rect 4416 26499 4456 26531
rect 4488 26499 4528 26531
rect 4560 26499 4600 26531
rect 4632 26499 4672 26531
rect 4704 26499 4744 26531
rect 4776 26499 4816 26531
rect 4848 26499 4888 26531
rect 4920 26499 4960 26531
rect 4992 26499 5032 26531
rect 5064 26499 5104 26531
rect 5136 26499 5176 26531
rect 5208 26499 5248 26531
rect 5280 26499 5320 26531
rect 5352 26499 5392 26531
rect 5424 26499 5464 26531
rect 5496 26499 5536 26531
rect 5568 26499 5608 26531
rect 5640 26499 5680 26531
rect 5712 26499 5752 26531
rect 5784 26499 5824 26531
rect 5856 26499 5896 26531
rect 5928 26499 5968 26531
rect 6000 26499 6040 26531
rect 6072 26499 6112 26531
rect 6144 26499 6184 26531
rect 6216 26499 6256 26531
rect 6288 26499 6328 26531
rect 6360 26499 6400 26531
rect 6432 26499 6472 26531
rect 6504 26499 6544 26531
rect 6576 26499 6616 26531
rect 6648 26499 6688 26531
rect 6720 26499 6760 26531
rect 6792 26499 6832 26531
rect 6864 26499 6904 26531
rect 6936 26499 6976 26531
rect 7008 26499 7048 26531
rect 7080 26499 7120 26531
rect 7152 26499 7192 26531
rect 7224 26499 7264 26531
rect 7296 26499 7336 26531
rect 7368 26499 7408 26531
rect 7440 26499 7480 26531
rect 7512 26499 7552 26531
rect 7584 26499 7624 26531
rect 7656 26499 7696 26531
rect 7728 26499 7768 26531
rect 7800 26499 7840 26531
rect 7872 26499 7912 26531
rect 7944 26499 7984 26531
rect 8016 26499 8056 26531
rect 8088 26499 8128 26531
rect 8160 26499 8200 26531
rect 8232 26499 8272 26531
rect 8304 26499 8344 26531
rect 8376 26499 8416 26531
rect 8448 26499 8488 26531
rect 8520 26499 8560 26531
rect 8592 26499 8632 26531
rect 8664 26499 8704 26531
rect 8736 26499 8776 26531
rect 8808 26499 8848 26531
rect 8880 26499 8920 26531
rect 8952 26499 8992 26531
rect 9024 26499 9064 26531
rect 9096 26499 9136 26531
rect 9168 26499 9208 26531
rect 9240 26499 9280 26531
rect 9312 26499 9352 26531
rect 9384 26499 9424 26531
rect 9456 26499 9496 26531
rect 9528 26499 9568 26531
rect 9600 26499 9640 26531
rect 9672 26499 9712 26531
rect 9744 26499 9784 26531
rect 9816 26499 9856 26531
rect 9888 26499 9928 26531
rect 9960 26499 10000 26531
rect 10032 26499 10072 26531
rect 10104 26499 10144 26531
rect 10176 26499 10216 26531
rect 10248 26499 10288 26531
rect 10320 26499 10360 26531
rect 10392 26499 10432 26531
rect 10464 26499 10504 26531
rect 10536 26499 10576 26531
rect 10608 26499 10648 26531
rect 10680 26499 10720 26531
rect 10752 26499 10792 26531
rect 10824 26499 10864 26531
rect 10896 26499 10936 26531
rect 10968 26499 11008 26531
rect 11040 26499 11080 26531
rect 11112 26499 11152 26531
rect 11184 26499 11224 26531
rect 11256 26499 11296 26531
rect 11328 26499 11368 26531
rect 11400 26499 11440 26531
rect 11472 26499 11512 26531
rect 11544 26499 11584 26531
rect 11616 26499 11656 26531
rect 11688 26499 11728 26531
rect 11760 26499 11800 26531
rect 11832 26499 11872 26531
rect 11904 26499 11944 26531
rect 11976 26499 12016 26531
rect 12048 26499 12088 26531
rect 12120 26499 12160 26531
rect 12192 26499 12232 26531
rect 12264 26499 12304 26531
rect 12336 26499 12376 26531
rect 12408 26499 12448 26531
rect 12480 26499 12520 26531
rect 12552 26499 12592 26531
rect 12624 26499 12664 26531
rect 12696 26499 12736 26531
rect 12768 26499 12808 26531
rect 12840 26499 12880 26531
rect 12912 26499 12952 26531
rect 12984 26499 13024 26531
rect 13056 26499 13096 26531
rect 13128 26499 13168 26531
rect 13200 26499 13240 26531
rect 13272 26499 13312 26531
rect 13344 26499 13384 26531
rect 13416 26499 13456 26531
rect 13488 26499 13528 26531
rect 13560 26499 13600 26531
rect 13632 26499 13672 26531
rect 13704 26499 13744 26531
rect 13776 26499 13816 26531
rect 13848 26499 13888 26531
rect 13920 26499 13960 26531
rect 13992 26499 14032 26531
rect 14064 26499 14104 26531
rect 14136 26499 14176 26531
rect 14208 26499 14248 26531
rect 14280 26499 14320 26531
rect 14352 26499 14392 26531
rect 14424 26499 14464 26531
rect 14496 26499 14536 26531
rect 14568 26499 14608 26531
rect 14640 26499 14680 26531
rect 14712 26499 14752 26531
rect 14784 26499 14824 26531
rect 14856 26499 14896 26531
rect 14928 26499 14968 26531
rect 15000 26499 15040 26531
rect 15072 26499 15112 26531
rect 15144 26499 15184 26531
rect 15216 26499 15256 26531
rect 15288 26499 15328 26531
rect 15360 26499 15400 26531
rect 15432 26499 15472 26531
rect 15504 26499 15544 26531
rect 15576 26499 15616 26531
rect 15648 26499 15688 26531
rect 15720 26499 15760 26531
rect 15792 26499 15832 26531
rect 15864 26499 15904 26531
rect 15936 26499 16000 26531
rect 0 26461 16000 26499
rect 0 26421 51 26461
rect 91 26459 149 26461
rect 189 26459 247 26461
rect 287 26459 345 26461
rect 385 26459 443 26461
rect 483 26459 541 26461
rect 581 26459 639 26461
rect 679 26459 737 26461
rect 777 26459 835 26461
rect 875 26459 933 26461
rect 973 26459 1031 26461
rect 1071 26459 1129 26461
rect 1169 26459 16000 26461
rect 96 26427 136 26459
rect 189 26427 208 26459
rect 240 26427 247 26459
rect 312 26427 345 26459
rect 385 26427 424 26459
rect 483 26427 496 26459
rect 528 26427 541 26459
rect 600 26427 639 26459
rect 679 26427 712 26459
rect 777 26427 784 26459
rect 816 26427 835 26459
rect 888 26427 928 26459
rect 973 26427 1000 26459
rect 1071 26427 1072 26459
rect 1104 26427 1129 26459
rect 1176 26427 1216 26459
rect 1248 26427 1288 26459
rect 1320 26427 1360 26459
rect 1392 26427 1432 26459
rect 1464 26427 1504 26459
rect 1536 26427 1576 26459
rect 1608 26427 1648 26459
rect 1680 26427 1720 26459
rect 1752 26427 1792 26459
rect 1824 26427 1864 26459
rect 1896 26427 1936 26459
rect 1968 26427 2008 26459
rect 2040 26427 2080 26459
rect 2112 26427 2152 26459
rect 2184 26427 2224 26459
rect 2256 26427 2296 26459
rect 2328 26427 2368 26459
rect 2400 26427 2440 26459
rect 2472 26427 2512 26459
rect 2544 26427 2584 26459
rect 2616 26427 2656 26459
rect 2688 26427 2728 26459
rect 2760 26427 2800 26459
rect 2832 26427 2872 26459
rect 2904 26427 2944 26459
rect 2976 26427 3016 26459
rect 3048 26427 3088 26459
rect 3120 26427 3160 26459
rect 3192 26427 3232 26459
rect 3264 26427 3304 26459
rect 3336 26427 3376 26459
rect 3408 26427 3448 26459
rect 3480 26427 3520 26459
rect 3552 26427 3592 26459
rect 3624 26427 3664 26459
rect 3696 26427 3736 26459
rect 3768 26427 3808 26459
rect 3840 26427 3880 26459
rect 3912 26427 3952 26459
rect 3984 26427 4024 26459
rect 4056 26427 4096 26459
rect 4128 26427 4168 26459
rect 4200 26427 4240 26459
rect 4272 26427 4312 26459
rect 4344 26427 4384 26459
rect 4416 26427 4456 26459
rect 4488 26427 4528 26459
rect 4560 26427 4600 26459
rect 4632 26427 4672 26459
rect 4704 26427 4744 26459
rect 4776 26427 4816 26459
rect 4848 26427 4888 26459
rect 4920 26427 4960 26459
rect 4992 26427 5032 26459
rect 5064 26427 5104 26459
rect 5136 26427 5176 26459
rect 5208 26427 5248 26459
rect 5280 26427 5320 26459
rect 5352 26427 5392 26459
rect 5424 26427 5464 26459
rect 5496 26427 5536 26459
rect 5568 26427 5608 26459
rect 5640 26427 5680 26459
rect 5712 26427 5752 26459
rect 5784 26427 5824 26459
rect 5856 26427 5896 26459
rect 5928 26427 5968 26459
rect 6000 26427 6040 26459
rect 6072 26427 6112 26459
rect 6144 26427 6184 26459
rect 6216 26427 6256 26459
rect 6288 26427 6328 26459
rect 6360 26427 6400 26459
rect 6432 26427 6472 26459
rect 6504 26427 6544 26459
rect 6576 26427 6616 26459
rect 6648 26427 6688 26459
rect 6720 26427 6760 26459
rect 6792 26427 6832 26459
rect 6864 26427 6904 26459
rect 6936 26427 6976 26459
rect 7008 26427 7048 26459
rect 7080 26427 7120 26459
rect 7152 26427 7192 26459
rect 7224 26427 7264 26459
rect 7296 26427 7336 26459
rect 7368 26427 7408 26459
rect 7440 26427 7480 26459
rect 7512 26427 7552 26459
rect 7584 26427 7624 26459
rect 7656 26427 7696 26459
rect 7728 26427 7768 26459
rect 7800 26427 7840 26459
rect 7872 26427 7912 26459
rect 7944 26427 7984 26459
rect 8016 26427 8056 26459
rect 8088 26427 8128 26459
rect 8160 26427 8200 26459
rect 8232 26427 8272 26459
rect 8304 26427 8344 26459
rect 8376 26427 8416 26459
rect 8448 26427 8488 26459
rect 8520 26427 8560 26459
rect 8592 26427 8632 26459
rect 8664 26427 8704 26459
rect 8736 26427 8776 26459
rect 8808 26427 8848 26459
rect 8880 26427 8920 26459
rect 8952 26427 8992 26459
rect 9024 26427 9064 26459
rect 9096 26427 9136 26459
rect 9168 26427 9208 26459
rect 9240 26427 9280 26459
rect 9312 26427 9352 26459
rect 9384 26427 9424 26459
rect 9456 26427 9496 26459
rect 9528 26427 9568 26459
rect 9600 26427 9640 26459
rect 9672 26427 9712 26459
rect 9744 26427 9784 26459
rect 9816 26427 9856 26459
rect 9888 26427 9928 26459
rect 9960 26427 10000 26459
rect 10032 26427 10072 26459
rect 10104 26427 10144 26459
rect 10176 26427 10216 26459
rect 10248 26427 10288 26459
rect 10320 26427 10360 26459
rect 10392 26427 10432 26459
rect 10464 26427 10504 26459
rect 10536 26427 10576 26459
rect 10608 26427 10648 26459
rect 10680 26427 10720 26459
rect 10752 26427 10792 26459
rect 10824 26427 10864 26459
rect 10896 26427 10936 26459
rect 10968 26427 11008 26459
rect 11040 26427 11080 26459
rect 11112 26427 11152 26459
rect 11184 26427 11224 26459
rect 11256 26427 11296 26459
rect 11328 26427 11368 26459
rect 11400 26427 11440 26459
rect 11472 26427 11512 26459
rect 11544 26427 11584 26459
rect 11616 26427 11656 26459
rect 11688 26427 11728 26459
rect 11760 26427 11800 26459
rect 11832 26427 11872 26459
rect 11904 26427 11944 26459
rect 11976 26427 12016 26459
rect 12048 26427 12088 26459
rect 12120 26427 12160 26459
rect 12192 26427 12232 26459
rect 12264 26427 12304 26459
rect 12336 26427 12376 26459
rect 12408 26427 12448 26459
rect 12480 26427 12520 26459
rect 12552 26427 12592 26459
rect 12624 26427 12664 26459
rect 12696 26427 12736 26459
rect 12768 26427 12808 26459
rect 12840 26427 12880 26459
rect 12912 26427 12952 26459
rect 12984 26427 13024 26459
rect 13056 26427 13096 26459
rect 13128 26427 13168 26459
rect 13200 26427 13240 26459
rect 13272 26427 13312 26459
rect 13344 26427 13384 26459
rect 13416 26427 13456 26459
rect 13488 26427 13528 26459
rect 13560 26427 13600 26459
rect 13632 26427 13672 26459
rect 13704 26427 13744 26459
rect 13776 26427 13816 26459
rect 13848 26427 13888 26459
rect 13920 26427 13960 26459
rect 13992 26427 14032 26459
rect 14064 26427 14104 26459
rect 14136 26427 14176 26459
rect 14208 26427 14248 26459
rect 14280 26427 14320 26459
rect 14352 26427 14392 26459
rect 14424 26427 14464 26459
rect 14496 26427 14536 26459
rect 14568 26427 14608 26459
rect 14640 26427 14680 26459
rect 14712 26427 14752 26459
rect 14784 26427 14824 26459
rect 14856 26427 14896 26459
rect 14928 26427 14968 26459
rect 15000 26427 15040 26459
rect 15072 26427 15112 26459
rect 15144 26427 15184 26459
rect 15216 26427 15256 26459
rect 15288 26427 15328 26459
rect 15360 26427 15400 26459
rect 15432 26427 15472 26459
rect 15504 26427 15544 26459
rect 15576 26427 15616 26459
rect 15648 26427 15688 26459
rect 15720 26427 15760 26459
rect 15792 26427 15832 26459
rect 15864 26427 15904 26459
rect 15936 26427 16000 26459
rect 91 26421 149 26427
rect 189 26421 247 26427
rect 287 26421 345 26427
rect 385 26421 443 26427
rect 483 26421 541 26427
rect 581 26421 639 26427
rect 679 26421 737 26427
rect 777 26421 835 26427
rect 875 26421 933 26427
rect 973 26421 1031 26427
rect 1071 26421 1129 26427
rect 1169 26421 16000 26427
rect 0 26387 16000 26421
rect 0 26363 64 26387
rect 0 26323 51 26363
rect 96 26355 136 26387
rect 168 26363 208 26387
rect 189 26355 208 26363
rect 240 26363 280 26387
rect 312 26363 352 26387
rect 384 26363 424 26387
rect 456 26363 496 26387
rect 240 26355 247 26363
rect 312 26355 345 26363
rect 385 26355 424 26363
rect 483 26355 496 26363
rect 528 26363 568 26387
rect 600 26363 640 26387
rect 672 26363 712 26387
rect 744 26363 784 26387
rect 528 26355 541 26363
rect 600 26355 639 26363
rect 679 26355 712 26363
rect 777 26355 784 26363
rect 816 26363 856 26387
rect 816 26355 835 26363
rect 888 26355 928 26387
rect 960 26363 1000 26387
rect 1032 26363 1072 26387
rect 973 26355 1000 26363
rect 1071 26355 1072 26363
rect 1104 26363 1144 26387
rect 1104 26355 1129 26363
rect 1176 26355 1216 26387
rect 1248 26355 1288 26387
rect 1320 26355 1360 26387
rect 1392 26355 1432 26387
rect 1464 26355 1504 26387
rect 1536 26355 1576 26387
rect 1608 26355 1648 26387
rect 1680 26355 1720 26387
rect 1752 26355 1792 26387
rect 1824 26355 1864 26387
rect 1896 26355 1936 26387
rect 1968 26355 2008 26387
rect 2040 26355 2080 26387
rect 2112 26355 2152 26387
rect 2184 26355 2224 26387
rect 2256 26355 2296 26387
rect 2328 26355 2368 26387
rect 2400 26355 2440 26387
rect 2472 26355 2512 26387
rect 2544 26355 2584 26387
rect 2616 26355 2656 26387
rect 2688 26355 2728 26387
rect 2760 26355 2800 26387
rect 2832 26355 2872 26387
rect 2904 26355 2944 26387
rect 2976 26355 3016 26387
rect 3048 26355 3088 26387
rect 3120 26355 3160 26387
rect 3192 26355 3232 26387
rect 3264 26355 3304 26387
rect 3336 26355 3376 26387
rect 3408 26355 3448 26387
rect 3480 26355 3520 26387
rect 3552 26355 3592 26387
rect 3624 26355 3664 26387
rect 3696 26355 3736 26387
rect 3768 26355 3808 26387
rect 3840 26355 3880 26387
rect 3912 26355 3952 26387
rect 3984 26355 4024 26387
rect 4056 26355 4096 26387
rect 4128 26355 4168 26387
rect 4200 26355 4240 26387
rect 4272 26355 4312 26387
rect 4344 26355 4384 26387
rect 4416 26355 4456 26387
rect 4488 26355 4528 26387
rect 4560 26355 4600 26387
rect 4632 26355 4672 26387
rect 4704 26355 4744 26387
rect 4776 26355 4816 26387
rect 4848 26355 4888 26387
rect 4920 26355 4960 26387
rect 4992 26355 5032 26387
rect 5064 26355 5104 26387
rect 5136 26355 5176 26387
rect 5208 26355 5248 26387
rect 5280 26355 5320 26387
rect 5352 26355 5392 26387
rect 5424 26355 5464 26387
rect 5496 26355 5536 26387
rect 5568 26355 5608 26387
rect 5640 26355 5680 26387
rect 5712 26355 5752 26387
rect 5784 26355 5824 26387
rect 5856 26355 5896 26387
rect 5928 26355 5968 26387
rect 6000 26355 6040 26387
rect 6072 26355 6112 26387
rect 6144 26355 6184 26387
rect 6216 26355 6256 26387
rect 6288 26355 6328 26387
rect 6360 26355 6400 26387
rect 6432 26355 6472 26387
rect 6504 26355 6544 26387
rect 6576 26355 6616 26387
rect 6648 26355 6688 26387
rect 6720 26355 6760 26387
rect 6792 26355 6832 26387
rect 6864 26355 6904 26387
rect 6936 26355 6976 26387
rect 7008 26355 7048 26387
rect 7080 26355 7120 26387
rect 7152 26355 7192 26387
rect 7224 26355 7264 26387
rect 7296 26355 7336 26387
rect 7368 26355 7408 26387
rect 7440 26355 7480 26387
rect 7512 26355 7552 26387
rect 7584 26355 7624 26387
rect 7656 26355 7696 26387
rect 7728 26355 7768 26387
rect 7800 26355 7840 26387
rect 7872 26355 7912 26387
rect 7944 26355 7984 26387
rect 8016 26355 8056 26387
rect 8088 26355 8128 26387
rect 8160 26355 8200 26387
rect 8232 26355 8272 26387
rect 8304 26355 8344 26387
rect 8376 26355 8416 26387
rect 8448 26355 8488 26387
rect 8520 26355 8560 26387
rect 8592 26355 8632 26387
rect 8664 26355 8704 26387
rect 8736 26355 8776 26387
rect 8808 26355 8848 26387
rect 8880 26355 8920 26387
rect 8952 26355 8992 26387
rect 9024 26355 9064 26387
rect 9096 26355 9136 26387
rect 9168 26355 9208 26387
rect 9240 26355 9280 26387
rect 9312 26355 9352 26387
rect 9384 26355 9424 26387
rect 9456 26355 9496 26387
rect 9528 26355 9568 26387
rect 9600 26355 9640 26387
rect 9672 26355 9712 26387
rect 9744 26355 9784 26387
rect 9816 26355 9856 26387
rect 9888 26355 9928 26387
rect 9960 26355 10000 26387
rect 10032 26355 10072 26387
rect 10104 26355 10144 26387
rect 10176 26355 10216 26387
rect 10248 26355 10288 26387
rect 10320 26355 10360 26387
rect 10392 26355 10432 26387
rect 10464 26355 10504 26387
rect 10536 26355 10576 26387
rect 10608 26355 10648 26387
rect 10680 26355 10720 26387
rect 10752 26355 10792 26387
rect 10824 26355 10864 26387
rect 10896 26355 10936 26387
rect 10968 26355 11008 26387
rect 11040 26355 11080 26387
rect 11112 26355 11152 26387
rect 11184 26355 11224 26387
rect 11256 26355 11296 26387
rect 11328 26355 11368 26387
rect 11400 26355 11440 26387
rect 11472 26355 11512 26387
rect 11544 26355 11584 26387
rect 11616 26355 11656 26387
rect 11688 26355 11728 26387
rect 11760 26355 11800 26387
rect 11832 26355 11872 26387
rect 11904 26355 11944 26387
rect 11976 26355 12016 26387
rect 12048 26355 12088 26387
rect 12120 26355 12160 26387
rect 12192 26355 12232 26387
rect 12264 26355 12304 26387
rect 12336 26355 12376 26387
rect 12408 26355 12448 26387
rect 12480 26355 12520 26387
rect 12552 26355 12592 26387
rect 12624 26355 12664 26387
rect 12696 26355 12736 26387
rect 12768 26355 12808 26387
rect 12840 26355 12880 26387
rect 12912 26355 12952 26387
rect 12984 26355 13024 26387
rect 13056 26355 13096 26387
rect 13128 26355 13168 26387
rect 13200 26355 13240 26387
rect 13272 26355 13312 26387
rect 13344 26355 13384 26387
rect 13416 26355 13456 26387
rect 13488 26355 13528 26387
rect 13560 26355 13600 26387
rect 13632 26355 13672 26387
rect 13704 26355 13744 26387
rect 13776 26355 13816 26387
rect 13848 26355 13888 26387
rect 13920 26355 13960 26387
rect 13992 26355 14032 26387
rect 14064 26355 14104 26387
rect 14136 26355 14176 26387
rect 14208 26355 14248 26387
rect 14280 26355 14320 26387
rect 14352 26355 14392 26387
rect 14424 26355 14464 26387
rect 14496 26355 14536 26387
rect 14568 26355 14608 26387
rect 14640 26355 14680 26387
rect 14712 26355 14752 26387
rect 14784 26355 14824 26387
rect 14856 26355 14896 26387
rect 14928 26355 14968 26387
rect 15000 26355 15040 26387
rect 15072 26355 15112 26387
rect 15144 26355 15184 26387
rect 15216 26355 15256 26387
rect 15288 26355 15328 26387
rect 15360 26355 15400 26387
rect 15432 26355 15472 26387
rect 15504 26355 15544 26387
rect 15576 26355 15616 26387
rect 15648 26355 15688 26387
rect 15720 26355 15760 26387
rect 15792 26355 15832 26387
rect 15864 26355 15904 26387
rect 15936 26355 16000 26387
rect 91 26323 149 26355
rect 189 26323 247 26355
rect 287 26323 345 26355
rect 385 26323 443 26355
rect 483 26323 541 26355
rect 581 26323 639 26355
rect 679 26323 737 26355
rect 777 26323 835 26355
rect 875 26323 933 26355
rect 973 26323 1031 26355
rect 1071 26323 1129 26355
rect 1169 26323 16000 26355
rect 0 26315 16000 26323
rect 0 26283 64 26315
rect 96 26283 136 26315
rect 168 26283 208 26315
rect 240 26283 280 26315
rect 312 26283 352 26315
rect 384 26283 424 26315
rect 456 26283 496 26315
rect 528 26283 568 26315
rect 600 26283 640 26315
rect 672 26283 712 26315
rect 744 26283 784 26315
rect 816 26283 856 26315
rect 888 26283 928 26315
rect 960 26283 1000 26315
rect 1032 26283 1072 26315
rect 1104 26283 1144 26315
rect 1176 26283 1216 26315
rect 1248 26283 1288 26315
rect 1320 26283 1360 26315
rect 1392 26283 1432 26315
rect 1464 26283 1504 26315
rect 1536 26283 1576 26315
rect 1608 26283 1648 26315
rect 1680 26283 1720 26315
rect 1752 26283 1792 26315
rect 1824 26283 1864 26315
rect 1896 26283 1936 26315
rect 1968 26283 2008 26315
rect 2040 26283 2080 26315
rect 2112 26283 2152 26315
rect 2184 26283 2224 26315
rect 2256 26283 2296 26315
rect 2328 26283 2368 26315
rect 2400 26283 2440 26315
rect 2472 26283 2512 26315
rect 2544 26283 2584 26315
rect 2616 26283 2656 26315
rect 2688 26283 2728 26315
rect 2760 26283 2800 26315
rect 2832 26283 2872 26315
rect 2904 26283 2944 26315
rect 2976 26283 3016 26315
rect 3048 26283 3088 26315
rect 3120 26283 3160 26315
rect 3192 26283 3232 26315
rect 3264 26283 3304 26315
rect 3336 26283 3376 26315
rect 3408 26283 3448 26315
rect 3480 26283 3520 26315
rect 3552 26283 3592 26315
rect 3624 26283 3664 26315
rect 3696 26283 3736 26315
rect 3768 26283 3808 26315
rect 3840 26283 3880 26315
rect 3912 26283 3952 26315
rect 3984 26283 4024 26315
rect 4056 26283 4096 26315
rect 4128 26283 4168 26315
rect 4200 26283 4240 26315
rect 4272 26283 4312 26315
rect 4344 26283 4384 26315
rect 4416 26283 4456 26315
rect 4488 26283 4528 26315
rect 4560 26283 4600 26315
rect 4632 26283 4672 26315
rect 4704 26283 4744 26315
rect 4776 26283 4816 26315
rect 4848 26283 4888 26315
rect 4920 26283 4960 26315
rect 4992 26283 5032 26315
rect 5064 26283 5104 26315
rect 5136 26283 5176 26315
rect 5208 26283 5248 26315
rect 5280 26283 5320 26315
rect 5352 26283 5392 26315
rect 5424 26283 5464 26315
rect 5496 26283 5536 26315
rect 5568 26283 5608 26315
rect 5640 26283 5680 26315
rect 5712 26283 5752 26315
rect 5784 26283 5824 26315
rect 5856 26283 5896 26315
rect 5928 26283 5968 26315
rect 6000 26283 6040 26315
rect 6072 26283 6112 26315
rect 6144 26283 6184 26315
rect 6216 26283 6256 26315
rect 6288 26283 6328 26315
rect 6360 26283 6400 26315
rect 6432 26283 6472 26315
rect 6504 26283 6544 26315
rect 6576 26283 6616 26315
rect 6648 26283 6688 26315
rect 6720 26283 6760 26315
rect 6792 26283 6832 26315
rect 6864 26283 6904 26315
rect 6936 26283 6976 26315
rect 7008 26283 7048 26315
rect 7080 26283 7120 26315
rect 7152 26283 7192 26315
rect 7224 26283 7264 26315
rect 7296 26283 7336 26315
rect 7368 26283 7408 26315
rect 7440 26283 7480 26315
rect 7512 26283 7552 26315
rect 7584 26283 7624 26315
rect 7656 26283 7696 26315
rect 7728 26283 7768 26315
rect 7800 26283 7840 26315
rect 7872 26283 7912 26315
rect 7944 26283 7984 26315
rect 8016 26283 8056 26315
rect 8088 26283 8128 26315
rect 8160 26283 8200 26315
rect 8232 26283 8272 26315
rect 8304 26283 8344 26315
rect 8376 26283 8416 26315
rect 8448 26283 8488 26315
rect 8520 26283 8560 26315
rect 8592 26283 8632 26315
rect 8664 26283 8704 26315
rect 8736 26283 8776 26315
rect 8808 26283 8848 26315
rect 8880 26283 8920 26315
rect 8952 26283 8992 26315
rect 9024 26283 9064 26315
rect 9096 26283 9136 26315
rect 9168 26283 9208 26315
rect 9240 26283 9280 26315
rect 9312 26283 9352 26315
rect 9384 26283 9424 26315
rect 9456 26283 9496 26315
rect 9528 26283 9568 26315
rect 9600 26283 9640 26315
rect 9672 26283 9712 26315
rect 9744 26283 9784 26315
rect 9816 26283 9856 26315
rect 9888 26283 9928 26315
rect 9960 26283 10000 26315
rect 10032 26283 10072 26315
rect 10104 26283 10144 26315
rect 10176 26283 10216 26315
rect 10248 26283 10288 26315
rect 10320 26283 10360 26315
rect 10392 26283 10432 26315
rect 10464 26283 10504 26315
rect 10536 26283 10576 26315
rect 10608 26283 10648 26315
rect 10680 26283 10720 26315
rect 10752 26283 10792 26315
rect 10824 26283 10864 26315
rect 10896 26283 10936 26315
rect 10968 26283 11008 26315
rect 11040 26283 11080 26315
rect 11112 26283 11152 26315
rect 11184 26283 11224 26315
rect 11256 26283 11296 26315
rect 11328 26283 11368 26315
rect 11400 26283 11440 26315
rect 11472 26283 11512 26315
rect 11544 26283 11584 26315
rect 11616 26283 11656 26315
rect 11688 26283 11728 26315
rect 11760 26283 11800 26315
rect 11832 26283 11872 26315
rect 11904 26283 11944 26315
rect 11976 26283 12016 26315
rect 12048 26283 12088 26315
rect 12120 26283 12160 26315
rect 12192 26283 12232 26315
rect 12264 26283 12304 26315
rect 12336 26283 12376 26315
rect 12408 26283 12448 26315
rect 12480 26283 12520 26315
rect 12552 26283 12592 26315
rect 12624 26283 12664 26315
rect 12696 26283 12736 26315
rect 12768 26283 12808 26315
rect 12840 26283 12880 26315
rect 12912 26283 12952 26315
rect 12984 26283 13024 26315
rect 13056 26283 13096 26315
rect 13128 26283 13168 26315
rect 13200 26283 13240 26315
rect 13272 26283 13312 26315
rect 13344 26283 13384 26315
rect 13416 26283 13456 26315
rect 13488 26283 13528 26315
rect 13560 26283 13600 26315
rect 13632 26283 13672 26315
rect 13704 26283 13744 26315
rect 13776 26283 13816 26315
rect 13848 26283 13888 26315
rect 13920 26283 13960 26315
rect 13992 26283 14032 26315
rect 14064 26283 14104 26315
rect 14136 26283 14176 26315
rect 14208 26283 14248 26315
rect 14280 26283 14320 26315
rect 14352 26283 14392 26315
rect 14424 26283 14464 26315
rect 14496 26283 14536 26315
rect 14568 26283 14608 26315
rect 14640 26283 14680 26315
rect 14712 26283 14752 26315
rect 14784 26283 14824 26315
rect 14856 26283 14896 26315
rect 14928 26283 14968 26315
rect 15000 26283 15040 26315
rect 15072 26283 15112 26315
rect 15144 26283 15184 26315
rect 15216 26283 15256 26315
rect 15288 26283 15328 26315
rect 15360 26283 15400 26315
rect 15432 26283 15472 26315
rect 15504 26283 15544 26315
rect 15576 26283 15616 26315
rect 15648 26283 15688 26315
rect 15720 26283 15760 26315
rect 15792 26283 15832 26315
rect 15864 26283 15904 26315
rect 15936 26283 16000 26315
rect 0 26265 16000 26283
rect 0 26225 51 26265
rect 91 26243 149 26265
rect 189 26243 247 26265
rect 287 26243 345 26265
rect 385 26243 443 26265
rect 483 26243 541 26265
rect 581 26243 639 26265
rect 679 26243 737 26265
rect 777 26243 835 26265
rect 875 26243 933 26265
rect 973 26243 1031 26265
rect 1071 26243 1129 26265
rect 1169 26243 16000 26265
rect 0 26211 64 26225
rect 96 26211 136 26243
rect 189 26225 208 26243
rect 168 26211 208 26225
rect 240 26225 247 26243
rect 312 26225 345 26243
rect 385 26225 424 26243
rect 483 26225 496 26243
rect 240 26211 280 26225
rect 312 26211 352 26225
rect 384 26211 424 26225
rect 456 26211 496 26225
rect 528 26225 541 26243
rect 600 26225 639 26243
rect 679 26225 712 26243
rect 777 26225 784 26243
rect 528 26211 568 26225
rect 600 26211 640 26225
rect 672 26211 712 26225
rect 744 26211 784 26225
rect 816 26225 835 26243
rect 816 26211 856 26225
rect 888 26211 928 26243
rect 973 26225 1000 26243
rect 1071 26225 1072 26243
rect 960 26211 1000 26225
rect 1032 26211 1072 26225
rect 1104 26225 1129 26243
rect 1104 26211 1144 26225
rect 1176 26211 1216 26243
rect 1248 26211 1288 26243
rect 1320 26211 1360 26243
rect 1392 26211 1432 26243
rect 1464 26211 1504 26243
rect 1536 26211 1576 26243
rect 1608 26211 1648 26243
rect 1680 26211 1720 26243
rect 1752 26211 1792 26243
rect 1824 26211 1864 26243
rect 1896 26211 1936 26243
rect 1968 26211 2008 26243
rect 2040 26211 2080 26243
rect 2112 26211 2152 26243
rect 2184 26211 2224 26243
rect 2256 26211 2296 26243
rect 2328 26211 2368 26243
rect 2400 26211 2440 26243
rect 2472 26211 2512 26243
rect 2544 26211 2584 26243
rect 2616 26211 2656 26243
rect 2688 26211 2728 26243
rect 2760 26211 2800 26243
rect 2832 26211 2872 26243
rect 2904 26211 2944 26243
rect 2976 26211 3016 26243
rect 3048 26211 3088 26243
rect 3120 26211 3160 26243
rect 3192 26211 3232 26243
rect 3264 26211 3304 26243
rect 3336 26211 3376 26243
rect 3408 26211 3448 26243
rect 3480 26211 3520 26243
rect 3552 26211 3592 26243
rect 3624 26211 3664 26243
rect 3696 26211 3736 26243
rect 3768 26211 3808 26243
rect 3840 26211 3880 26243
rect 3912 26211 3952 26243
rect 3984 26211 4024 26243
rect 4056 26211 4096 26243
rect 4128 26211 4168 26243
rect 4200 26211 4240 26243
rect 4272 26211 4312 26243
rect 4344 26211 4384 26243
rect 4416 26211 4456 26243
rect 4488 26211 4528 26243
rect 4560 26211 4600 26243
rect 4632 26211 4672 26243
rect 4704 26211 4744 26243
rect 4776 26211 4816 26243
rect 4848 26211 4888 26243
rect 4920 26211 4960 26243
rect 4992 26211 5032 26243
rect 5064 26211 5104 26243
rect 5136 26211 5176 26243
rect 5208 26211 5248 26243
rect 5280 26211 5320 26243
rect 5352 26211 5392 26243
rect 5424 26211 5464 26243
rect 5496 26211 5536 26243
rect 5568 26211 5608 26243
rect 5640 26211 5680 26243
rect 5712 26211 5752 26243
rect 5784 26211 5824 26243
rect 5856 26211 5896 26243
rect 5928 26211 5968 26243
rect 6000 26211 6040 26243
rect 6072 26211 6112 26243
rect 6144 26211 6184 26243
rect 6216 26211 6256 26243
rect 6288 26211 6328 26243
rect 6360 26211 6400 26243
rect 6432 26211 6472 26243
rect 6504 26211 6544 26243
rect 6576 26211 6616 26243
rect 6648 26211 6688 26243
rect 6720 26211 6760 26243
rect 6792 26211 6832 26243
rect 6864 26211 6904 26243
rect 6936 26211 6976 26243
rect 7008 26211 7048 26243
rect 7080 26211 7120 26243
rect 7152 26211 7192 26243
rect 7224 26211 7264 26243
rect 7296 26211 7336 26243
rect 7368 26211 7408 26243
rect 7440 26211 7480 26243
rect 7512 26211 7552 26243
rect 7584 26211 7624 26243
rect 7656 26211 7696 26243
rect 7728 26211 7768 26243
rect 7800 26211 7840 26243
rect 7872 26211 7912 26243
rect 7944 26211 7984 26243
rect 8016 26211 8056 26243
rect 8088 26211 8128 26243
rect 8160 26211 8200 26243
rect 8232 26211 8272 26243
rect 8304 26211 8344 26243
rect 8376 26211 8416 26243
rect 8448 26211 8488 26243
rect 8520 26211 8560 26243
rect 8592 26211 8632 26243
rect 8664 26211 8704 26243
rect 8736 26211 8776 26243
rect 8808 26211 8848 26243
rect 8880 26211 8920 26243
rect 8952 26211 8992 26243
rect 9024 26211 9064 26243
rect 9096 26211 9136 26243
rect 9168 26211 9208 26243
rect 9240 26211 9280 26243
rect 9312 26211 9352 26243
rect 9384 26211 9424 26243
rect 9456 26211 9496 26243
rect 9528 26211 9568 26243
rect 9600 26211 9640 26243
rect 9672 26211 9712 26243
rect 9744 26211 9784 26243
rect 9816 26211 9856 26243
rect 9888 26211 9928 26243
rect 9960 26211 10000 26243
rect 10032 26211 10072 26243
rect 10104 26211 10144 26243
rect 10176 26211 10216 26243
rect 10248 26211 10288 26243
rect 10320 26211 10360 26243
rect 10392 26211 10432 26243
rect 10464 26211 10504 26243
rect 10536 26211 10576 26243
rect 10608 26211 10648 26243
rect 10680 26211 10720 26243
rect 10752 26211 10792 26243
rect 10824 26211 10864 26243
rect 10896 26211 10936 26243
rect 10968 26211 11008 26243
rect 11040 26211 11080 26243
rect 11112 26211 11152 26243
rect 11184 26211 11224 26243
rect 11256 26211 11296 26243
rect 11328 26211 11368 26243
rect 11400 26211 11440 26243
rect 11472 26211 11512 26243
rect 11544 26211 11584 26243
rect 11616 26211 11656 26243
rect 11688 26211 11728 26243
rect 11760 26211 11800 26243
rect 11832 26211 11872 26243
rect 11904 26211 11944 26243
rect 11976 26211 12016 26243
rect 12048 26211 12088 26243
rect 12120 26211 12160 26243
rect 12192 26211 12232 26243
rect 12264 26211 12304 26243
rect 12336 26211 12376 26243
rect 12408 26211 12448 26243
rect 12480 26211 12520 26243
rect 12552 26211 12592 26243
rect 12624 26211 12664 26243
rect 12696 26211 12736 26243
rect 12768 26211 12808 26243
rect 12840 26211 12880 26243
rect 12912 26211 12952 26243
rect 12984 26211 13024 26243
rect 13056 26211 13096 26243
rect 13128 26211 13168 26243
rect 13200 26211 13240 26243
rect 13272 26211 13312 26243
rect 13344 26211 13384 26243
rect 13416 26211 13456 26243
rect 13488 26211 13528 26243
rect 13560 26211 13600 26243
rect 13632 26211 13672 26243
rect 13704 26211 13744 26243
rect 13776 26211 13816 26243
rect 13848 26211 13888 26243
rect 13920 26211 13960 26243
rect 13992 26211 14032 26243
rect 14064 26211 14104 26243
rect 14136 26211 14176 26243
rect 14208 26211 14248 26243
rect 14280 26211 14320 26243
rect 14352 26211 14392 26243
rect 14424 26211 14464 26243
rect 14496 26211 14536 26243
rect 14568 26211 14608 26243
rect 14640 26211 14680 26243
rect 14712 26211 14752 26243
rect 14784 26211 14824 26243
rect 14856 26211 14896 26243
rect 14928 26211 14968 26243
rect 15000 26211 15040 26243
rect 15072 26211 15112 26243
rect 15144 26211 15184 26243
rect 15216 26211 15256 26243
rect 15288 26211 15328 26243
rect 15360 26211 15400 26243
rect 15432 26211 15472 26243
rect 15504 26211 15544 26243
rect 15576 26211 15616 26243
rect 15648 26211 15688 26243
rect 15720 26211 15760 26243
rect 15792 26211 15832 26243
rect 15864 26211 15904 26243
rect 15936 26211 16000 26243
rect 0 26171 16000 26211
rect 0 26167 64 26171
rect 0 26127 51 26167
rect 96 26139 136 26171
rect 168 26167 208 26171
rect 189 26139 208 26167
rect 240 26167 280 26171
rect 312 26167 352 26171
rect 384 26167 424 26171
rect 456 26167 496 26171
rect 240 26139 247 26167
rect 312 26139 345 26167
rect 385 26139 424 26167
rect 483 26139 496 26167
rect 528 26167 568 26171
rect 600 26167 640 26171
rect 672 26167 712 26171
rect 744 26167 784 26171
rect 528 26139 541 26167
rect 600 26139 639 26167
rect 679 26139 712 26167
rect 777 26139 784 26167
rect 816 26167 856 26171
rect 816 26139 835 26167
rect 888 26139 928 26171
rect 960 26167 1000 26171
rect 1032 26167 1072 26171
rect 973 26139 1000 26167
rect 1071 26139 1072 26167
rect 1104 26167 1144 26171
rect 1104 26139 1129 26167
rect 1176 26139 1216 26171
rect 1248 26139 1288 26171
rect 1320 26139 1360 26171
rect 1392 26139 1432 26171
rect 1464 26139 1504 26171
rect 1536 26139 1576 26171
rect 1608 26139 1648 26171
rect 1680 26139 1720 26171
rect 1752 26139 1792 26171
rect 1824 26139 1864 26171
rect 1896 26139 1936 26171
rect 1968 26139 2008 26171
rect 2040 26139 2080 26171
rect 2112 26139 2152 26171
rect 2184 26139 2224 26171
rect 2256 26139 2296 26171
rect 2328 26139 2368 26171
rect 2400 26139 2440 26171
rect 2472 26139 2512 26171
rect 2544 26139 2584 26171
rect 2616 26139 2656 26171
rect 2688 26139 2728 26171
rect 2760 26139 2800 26171
rect 2832 26139 2872 26171
rect 2904 26139 2944 26171
rect 2976 26139 3016 26171
rect 3048 26139 3088 26171
rect 3120 26139 3160 26171
rect 3192 26139 3232 26171
rect 3264 26139 3304 26171
rect 3336 26139 3376 26171
rect 3408 26139 3448 26171
rect 3480 26139 3520 26171
rect 3552 26139 3592 26171
rect 3624 26139 3664 26171
rect 3696 26139 3736 26171
rect 3768 26139 3808 26171
rect 3840 26139 3880 26171
rect 3912 26139 3952 26171
rect 3984 26139 4024 26171
rect 4056 26139 4096 26171
rect 4128 26139 4168 26171
rect 4200 26139 4240 26171
rect 4272 26139 4312 26171
rect 4344 26139 4384 26171
rect 4416 26139 4456 26171
rect 4488 26139 4528 26171
rect 4560 26139 4600 26171
rect 4632 26139 4672 26171
rect 4704 26139 4744 26171
rect 4776 26139 4816 26171
rect 4848 26139 4888 26171
rect 4920 26139 4960 26171
rect 4992 26139 5032 26171
rect 5064 26139 5104 26171
rect 5136 26139 5176 26171
rect 5208 26139 5248 26171
rect 5280 26139 5320 26171
rect 5352 26139 5392 26171
rect 5424 26139 5464 26171
rect 5496 26139 5536 26171
rect 5568 26139 5608 26171
rect 5640 26139 5680 26171
rect 5712 26139 5752 26171
rect 5784 26139 5824 26171
rect 5856 26139 5896 26171
rect 5928 26139 5968 26171
rect 6000 26139 6040 26171
rect 6072 26139 6112 26171
rect 6144 26139 6184 26171
rect 6216 26139 6256 26171
rect 6288 26139 6328 26171
rect 6360 26139 6400 26171
rect 6432 26139 6472 26171
rect 6504 26139 6544 26171
rect 6576 26139 6616 26171
rect 6648 26139 6688 26171
rect 6720 26139 6760 26171
rect 6792 26139 6832 26171
rect 6864 26139 6904 26171
rect 6936 26139 6976 26171
rect 7008 26139 7048 26171
rect 7080 26139 7120 26171
rect 7152 26139 7192 26171
rect 7224 26139 7264 26171
rect 7296 26139 7336 26171
rect 7368 26139 7408 26171
rect 7440 26139 7480 26171
rect 7512 26139 7552 26171
rect 7584 26139 7624 26171
rect 7656 26139 7696 26171
rect 7728 26139 7768 26171
rect 7800 26139 7840 26171
rect 7872 26139 7912 26171
rect 7944 26139 7984 26171
rect 8016 26139 8056 26171
rect 8088 26139 8128 26171
rect 8160 26139 8200 26171
rect 8232 26139 8272 26171
rect 8304 26139 8344 26171
rect 8376 26139 8416 26171
rect 8448 26139 8488 26171
rect 8520 26139 8560 26171
rect 8592 26139 8632 26171
rect 8664 26139 8704 26171
rect 8736 26139 8776 26171
rect 8808 26139 8848 26171
rect 8880 26139 8920 26171
rect 8952 26139 8992 26171
rect 9024 26139 9064 26171
rect 9096 26139 9136 26171
rect 9168 26139 9208 26171
rect 9240 26139 9280 26171
rect 9312 26139 9352 26171
rect 9384 26139 9424 26171
rect 9456 26139 9496 26171
rect 9528 26139 9568 26171
rect 9600 26139 9640 26171
rect 9672 26139 9712 26171
rect 9744 26139 9784 26171
rect 9816 26139 9856 26171
rect 9888 26139 9928 26171
rect 9960 26139 10000 26171
rect 10032 26139 10072 26171
rect 10104 26139 10144 26171
rect 10176 26139 10216 26171
rect 10248 26139 10288 26171
rect 10320 26139 10360 26171
rect 10392 26139 10432 26171
rect 10464 26139 10504 26171
rect 10536 26139 10576 26171
rect 10608 26139 10648 26171
rect 10680 26139 10720 26171
rect 10752 26139 10792 26171
rect 10824 26139 10864 26171
rect 10896 26139 10936 26171
rect 10968 26139 11008 26171
rect 11040 26139 11080 26171
rect 11112 26139 11152 26171
rect 11184 26139 11224 26171
rect 11256 26139 11296 26171
rect 11328 26139 11368 26171
rect 11400 26139 11440 26171
rect 11472 26139 11512 26171
rect 11544 26139 11584 26171
rect 11616 26139 11656 26171
rect 11688 26139 11728 26171
rect 11760 26139 11800 26171
rect 11832 26139 11872 26171
rect 11904 26139 11944 26171
rect 11976 26139 12016 26171
rect 12048 26139 12088 26171
rect 12120 26139 12160 26171
rect 12192 26139 12232 26171
rect 12264 26139 12304 26171
rect 12336 26139 12376 26171
rect 12408 26139 12448 26171
rect 12480 26139 12520 26171
rect 12552 26139 12592 26171
rect 12624 26139 12664 26171
rect 12696 26139 12736 26171
rect 12768 26139 12808 26171
rect 12840 26139 12880 26171
rect 12912 26139 12952 26171
rect 12984 26139 13024 26171
rect 13056 26139 13096 26171
rect 13128 26139 13168 26171
rect 13200 26139 13240 26171
rect 13272 26139 13312 26171
rect 13344 26139 13384 26171
rect 13416 26139 13456 26171
rect 13488 26139 13528 26171
rect 13560 26139 13600 26171
rect 13632 26139 13672 26171
rect 13704 26139 13744 26171
rect 13776 26139 13816 26171
rect 13848 26139 13888 26171
rect 13920 26139 13960 26171
rect 13992 26139 14032 26171
rect 14064 26139 14104 26171
rect 14136 26139 14176 26171
rect 14208 26139 14248 26171
rect 14280 26139 14320 26171
rect 14352 26139 14392 26171
rect 14424 26139 14464 26171
rect 14496 26139 14536 26171
rect 14568 26139 14608 26171
rect 14640 26139 14680 26171
rect 14712 26139 14752 26171
rect 14784 26139 14824 26171
rect 14856 26139 14896 26171
rect 14928 26139 14968 26171
rect 15000 26139 15040 26171
rect 15072 26139 15112 26171
rect 15144 26139 15184 26171
rect 15216 26139 15256 26171
rect 15288 26139 15328 26171
rect 15360 26139 15400 26171
rect 15432 26139 15472 26171
rect 15504 26139 15544 26171
rect 15576 26139 15616 26171
rect 15648 26139 15688 26171
rect 15720 26139 15760 26171
rect 15792 26139 15832 26171
rect 15864 26139 15904 26171
rect 15936 26139 16000 26171
rect 91 26127 149 26139
rect 189 26127 247 26139
rect 287 26127 345 26139
rect 385 26127 443 26139
rect 483 26127 541 26139
rect 581 26127 639 26139
rect 679 26127 737 26139
rect 777 26127 835 26139
rect 875 26127 933 26139
rect 973 26127 1031 26139
rect 1071 26127 1129 26139
rect 1169 26127 16000 26139
rect 0 26099 16000 26127
rect 0 26069 64 26099
rect 0 26029 51 26069
rect 96 26067 136 26099
rect 168 26069 208 26099
rect 189 26067 208 26069
rect 240 26069 280 26099
rect 312 26069 352 26099
rect 384 26069 424 26099
rect 456 26069 496 26099
rect 240 26067 247 26069
rect 312 26067 345 26069
rect 385 26067 424 26069
rect 483 26067 496 26069
rect 528 26069 568 26099
rect 600 26069 640 26099
rect 672 26069 712 26099
rect 744 26069 784 26099
rect 528 26067 541 26069
rect 600 26067 639 26069
rect 679 26067 712 26069
rect 777 26067 784 26069
rect 816 26069 856 26099
rect 816 26067 835 26069
rect 888 26067 928 26099
rect 960 26069 1000 26099
rect 1032 26069 1072 26099
rect 973 26067 1000 26069
rect 1071 26067 1072 26069
rect 1104 26069 1144 26099
rect 1104 26067 1129 26069
rect 1176 26067 1216 26099
rect 1248 26067 1288 26099
rect 1320 26067 1360 26099
rect 1392 26067 1432 26099
rect 1464 26067 1504 26099
rect 1536 26067 1576 26099
rect 1608 26067 1648 26099
rect 1680 26067 1720 26099
rect 1752 26067 1792 26099
rect 1824 26067 1864 26099
rect 1896 26067 1936 26099
rect 1968 26067 2008 26099
rect 2040 26067 2080 26099
rect 2112 26067 2152 26099
rect 2184 26067 2224 26099
rect 2256 26067 2296 26099
rect 2328 26067 2368 26099
rect 2400 26067 2440 26099
rect 2472 26067 2512 26099
rect 2544 26067 2584 26099
rect 2616 26067 2656 26099
rect 2688 26067 2728 26099
rect 2760 26067 2800 26099
rect 2832 26067 2872 26099
rect 2904 26067 2944 26099
rect 2976 26067 3016 26099
rect 3048 26067 3088 26099
rect 3120 26067 3160 26099
rect 3192 26067 3232 26099
rect 3264 26067 3304 26099
rect 3336 26067 3376 26099
rect 3408 26067 3448 26099
rect 3480 26067 3520 26099
rect 3552 26067 3592 26099
rect 3624 26067 3664 26099
rect 3696 26067 3736 26099
rect 3768 26067 3808 26099
rect 3840 26067 3880 26099
rect 3912 26067 3952 26099
rect 3984 26067 4024 26099
rect 4056 26067 4096 26099
rect 4128 26067 4168 26099
rect 4200 26067 4240 26099
rect 4272 26067 4312 26099
rect 4344 26067 4384 26099
rect 4416 26067 4456 26099
rect 4488 26067 4528 26099
rect 4560 26067 4600 26099
rect 4632 26067 4672 26099
rect 4704 26067 4744 26099
rect 4776 26067 4816 26099
rect 4848 26067 4888 26099
rect 4920 26067 4960 26099
rect 4992 26067 5032 26099
rect 5064 26067 5104 26099
rect 5136 26067 5176 26099
rect 5208 26067 5248 26099
rect 5280 26067 5320 26099
rect 5352 26067 5392 26099
rect 5424 26067 5464 26099
rect 5496 26067 5536 26099
rect 5568 26067 5608 26099
rect 5640 26067 5680 26099
rect 5712 26067 5752 26099
rect 5784 26067 5824 26099
rect 5856 26067 5896 26099
rect 5928 26067 5968 26099
rect 6000 26067 6040 26099
rect 6072 26067 6112 26099
rect 6144 26067 6184 26099
rect 6216 26067 6256 26099
rect 6288 26067 6328 26099
rect 6360 26067 6400 26099
rect 6432 26067 6472 26099
rect 6504 26067 6544 26099
rect 6576 26067 6616 26099
rect 6648 26067 6688 26099
rect 6720 26067 6760 26099
rect 6792 26067 6832 26099
rect 6864 26067 6904 26099
rect 6936 26067 6976 26099
rect 7008 26067 7048 26099
rect 7080 26067 7120 26099
rect 7152 26067 7192 26099
rect 7224 26067 7264 26099
rect 7296 26067 7336 26099
rect 7368 26067 7408 26099
rect 7440 26067 7480 26099
rect 7512 26067 7552 26099
rect 7584 26067 7624 26099
rect 7656 26067 7696 26099
rect 7728 26067 7768 26099
rect 7800 26067 7840 26099
rect 7872 26067 7912 26099
rect 7944 26067 7984 26099
rect 8016 26067 8056 26099
rect 8088 26067 8128 26099
rect 8160 26067 8200 26099
rect 8232 26067 8272 26099
rect 8304 26067 8344 26099
rect 8376 26067 8416 26099
rect 8448 26067 8488 26099
rect 8520 26067 8560 26099
rect 8592 26067 8632 26099
rect 8664 26067 8704 26099
rect 8736 26067 8776 26099
rect 8808 26067 8848 26099
rect 8880 26067 8920 26099
rect 8952 26067 8992 26099
rect 9024 26067 9064 26099
rect 9096 26067 9136 26099
rect 9168 26067 9208 26099
rect 9240 26067 9280 26099
rect 9312 26067 9352 26099
rect 9384 26067 9424 26099
rect 9456 26067 9496 26099
rect 9528 26067 9568 26099
rect 9600 26067 9640 26099
rect 9672 26067 9712 26099
rect 9744 26067 9784 26099
rect 9816 26067 9856 26099
rect 9888 26067 9928 26099
rect 9960 26067 10000 26099
rect 10032 26067 10072 26099
rect 10104 26067 10144 26099
rect 10176 26067 10216 26099
rect 10248 26067 10288 26099
rect 10320 26067 10360 26099
rect 10392 26067 10432 26099
rect 10464 26067 10504 26099
rect 10536 26067 10576 26099
rect 10608 26067 10648 26099
rect 10680 26067 10720 26099
rect 10752 26067 10792 26099
rect 10824 26067 10864 26099
rect 10896 26067 10936 26099
rect 10968 26067 11008 26099
rect 11040 26067 11080 26099
rect 11112 26067 11152 26099
rect 11184 26067 11224 26099
rect 11256 26067 11296 26099
rect 11328 26067 11368 26099
rect 11400 26067 11440 26099
rect 11472 26067 11512 26099
rect 11544 26067 11584 26099
rect 11616 26067 11656 26099
rect 11688 26067 11728 26099
rect 11760 26067 11800 26099
rect 11832 26067 11872 26099
rect 11904 26067 11944 26099
rect 11976 26067 12016 26099
rect 12048 26067 12088 26099
rect 12120 26067 12160 26099
rect 12192 26067 12232 26099
rect 12264 26067 12304 26099
rect 12336 26067 12376 26099
rect 12408 26067 12448 26099
rect 12480 26067 12520 26099
rect 12552 26067 12592 26099
rect 12624 26067 12664 26099
rect 12696 26067 12736 26099
rect 12768 26067 12808 26099
rect 12840 26067 12880 26099
rect 12912 26067 12952 26099
rect 12984 26067 13024 26099
rect 13056 26067 13096 26099
rect 13128 26067 13168 26099
rect 13200 26067 13240 26099
rect 13272 26067 13312 26099
rect 13344 26067 13384 26099
rect 13416 26067 13456 26099
rect 13488 26067 13528 26099
rect 13560 26067 13600 26099
rect 13632 26067 13672 26099
rect 13704 26067 13744 26099
rect 13776 26067 13816 26099
rect 13848 26067 13888 26099
rect 13920 26067 13960 26099
rect 13992 26067 14032 26099
rect 14064 26067 14104 26099
rect 14136 26067 14176 26099
rect 14208 26067 14248 26099
rect 14280 26067 14320 26099
rect 14352 26067 14392 26099
rect 14424 26067 14464 26099
rect 14496 26067 14536 26099
rect 14568 26067 14608 26099
rect 14640 26067 14680 26099
rect 14712 26067 14752 26099
rect 14784 26067 14824 26099
rect 14856 26067 14896 26099
rect 14928 26067 14968 26099
rect 15000 26067 15040 26099
rect 15072 26067 15112 26099
rect 15144 26067 15184 26099
rect 15216 26067 15256 26099
rect 15288 26067 15328 26099
rect 15360 26067 15400 26099
rect 15432 26067 15472 26099
rect 15504 26067 15544 26099
rect 15576 26067 15616 26099
rect 15648 26067 15688 26099
rect 15720 26067 15760 26099
rect 15792 26067 15832 26099
rect 15864 26067 15904 26099
rect 15936 26067 16000 26099
rect 91 26029 149 26067
rect 189 26029 247 26067
rect 287 26029 345 26067
rect 385 26029 443 26067
rect 483 26029 541 26067
rect 581 26029 639 26067
rect 679 26029 737 26067
rect 777 26029 835 26067
rect 875 26029 933 26067
rect 973 26029 1031 26067
rect 1071 26029 1129 26067
rect 1169 26029 16000 26067
rect 0 26027 16000 26029
rect 0 25995 64 26027
rect 96 25995 136 26027
rect 168 25995 208 26027
rect 240 25995 280 26027
rect 312 25995 352 26027
rect 384 25995 424 26027
rect 456 25995 496 26027
rect 528 25995 568 26027
rect 600 25995 640 26027
rect 672 25995 712 26027
rect 744 25995 784 26027
rect 816 25995 856 26027
rect 888 25995 928 26027
rect 960 25995 1000 26027
rect 1032 25995 1072 26027
rect 1104 25995 1144 26027
rect 1176 25995 1216 26027
rect 1248 25995 1288 26027
rect 1320 25995 1360 26027
rect 1392 25995 1432 26027
rect 1464 25995 1504 26027
rect 1536 25995 1576 26027
rect 1608 25995 1648 26027
rect 1680 25995 1720 26027
rect 1752 25995 1792 26027
rect 1824 25995 1864 26027
rect 1896 25995 1936 26027
rect 1968 25995 2008 26027
rect 2040 25995 2080 26027
rect 2112 25995 2152 26027
rect 2184 25995 2224 26027
rect 2256 25995 2296 26027
rect 2328 25995 2368 26027
rect 2400 25995 2440 26027
rect 2472 25995 2512 26027
rect 2544 25995 2584 26027
rect 2616 25995 2656 26027
rect 2688 25995 2728 26027
rect 2760 25995 2800 26027
rect 2832 25995 2872 26027
rect 2904 25995 2944 26027
rect 2976 25995 3016 26027
rect 3048 25995 3088 26027
rect 3120 25995 3160 26027
rect 3192 25995 3232 26027
rect 3264 25995 3304 26027
rect 3336 25995 3376 26027
rect 3408 25995 3448 26027
rect 3480 25995 3520 26027
rect 3552 25995 3592 26027
rect 3624 25995 3664 26027
rect 3696 25995 3736 26027
rect 3768 25995 3808 26027
rect 3840 25995 3880 26027
rect 3912 25995 3952 26027
rect 3984 25995 4024 26027
rect 4056 25995 4096 26027
rect 4128 25995 4168 26027
rect 4200 25995 4240 26027
rect 4272 25995 4312 26027
rect 4344 25995 4384 26027
rect 4416 25995 4456 26027
rect 4488 25995 4528 26027
rect 4560 25995 4600 26027
rect 4632 25995 4672 26027
rect 4704 25995 4744 26027
rect 4776 25995 4816 26027
rect 4848 25995 4888 26027
rect 4920 25995 4960 26027
rect 4992 25995 5032 26027
rect 5064 25995 5104 26027
rect 5136 25995 5176 26027
rect 5208 25995 5248 26027
rect 5280 25995 5320 26027
rect 5352 25995 5392 26027
rect 5424 25995 5464 26027
rect 5496 25995 5536 26027
rect 5568 25995 5608 26027
rect 5640 25995 5680 26027
rect 5712 25995 5752 26027
rect 5784 25995 5824 26027
rect 5856 25995 5896 26027
rect 5928 25995 5968 26027
rect 6000 25995 6040 26027
rect 6072 25995 6112 26027
rect 6144 25995 6184 26027
rect 6216 25995 6256 26027
rect 6288 25995 6328 26027
rect 6360 25995 6400 26027
rect 6432 25995 6472 26027
rect 6504 25995 6544 26027
rect 6576 25995 6616 26027
rect 6648 25995 6688 26027
rect 6720 25995 6760 26027
rect 6792 25995 6832 26027
rect 6864 25995 6904 26027
rect 6936 25995 6976 26027
rect 7008 25995 7048 26027
rect 7080 25995 7120 26027
rect 7152 25995 7192 26027
rect 7224 25995 7264 26027
rect 7296 25995 7336 26027
rect 7368 25995 7408 26027
rect 7440 25995 7480 26027
rect 7512 25995 7552 26027
rect 7584 25995 7624 26027
rect 7656 25995 7696 26027
rect 7728 25995 7768 26027
rect 7800 25995 7840 26027
rect 7872 25995 7912 26027
rect 7944 25995 7984 26027
rect 8016 25995 8056 26027
rect 8088 25995 8128 26027
rect 8160 25995 8200 26027
rect 8232 25995 8272 26027
rect 8304 25995 8344 26027
rect 8376 25995 8416 26027
rect 8448 25995 8488 26027
rect 8520 25995 8560 26027
rect 8592 25995 8632 26027
rect 8664 25995 8704 26027
rect 8736 25995 8776 26027
rect 8808 25995 8848 26027
rect 8880 25995 8920 26027
rect 8952 25995 8992 26027
rect 9024 25995 9064 26027
rect 9096 25995 9136 26027
rect 9168 25995 9208 26027
rect 9240 25995 9280 26027
rect 9312 25995 9352 26027
rect 9384 25995 9424 26027
rect 9456 25995 9496 26027
rect 9528 25995 9568 26027
rect 9600 25995 9640 26027
rect 9672 25995 9712 26027
rect 9744 25995 9784 26027
rect 9816 25995 9856 26027
rect 9888 25995 9928 26027
rect 9960 25995 10000 26027
rect 10032 25995 10072 26027
rect 10104 25995 10144 26027
rect 10176 25995 10216 26027
rect 10248 25995 10288 26027
rect 10320 25995 10360 26027
rect 10392 25995 10432 26027
rect 10464 25995 10504 26027
rect 10536 25995 10576 26027
rect 10608 25995 10648 26027
rect 10680 25995 10720 26027
rect 10752 25995 10792 26027
rect 10824 25995 10864 26027
rect 10896 25995 10936 26027
rect 10968 25995 11008 26027
rect 11040 25995 11080 26027
rect 11112 25995 11152 26027
rect 11184 25995 11224 26027
rect 11256 25995 11296 26027
rect 11328 25995 11368 26027
rect 11400 25995 11440 26027
rect 11472 25995 11512 26027
rect 11544 25995 11584 26027
rect 11616 25995 11656 26027
rect 11688 25995 11728 26027
rect 11760 25995 11800 26027
rect 11832 25995 11872 26027
rect 11904 25995 11944 26027
rect 11976 25995 12016 26027
rect 12048 25995 12088 26027
rect 12120 25995 12160 26027
rect 12192 25995 12232 26027
rect 12264 25995 12304 26027
rect 12336 25995 12376 26027
rect 12408 25995 12448 26027
rect 12480 25995 12520 26027
rect 12552 25995 12592 26027
rect 12624 25995 12664 26027
rect 12696 25995 12736 26027
rect 12768 25995 12808 26027
rect 12840 25995 12880 26027
rect 12912 25995 12952 26027
rect 12984 25995 13024 26027
rect 13056 25995 13096 26027
rect 13128 25995 13168 26027
rect 13200 25995 13240 26027
rect 13272 25995 13312 26027
rect 13344 25995 13384 26027
rect 13416 25995 13456 26027
rect 13488 25995 13528 26027
rect 13560 25995 13600 26027
rect 13632 25995 13672 26027
rect 13704 25995 13744 26027
rect 13776 25995 13816 26027
rect 13848 25995 13888 26027
rect 13920 25995 13960 26027
rect 13992 25995 14032 26027
rect 14064 25995 14104 26027
rect 14136 25995 14176 26027
rect 14208 25995 14248 26027
rect 14280 25995 14320 26027
rect 14352 25995 14392 26027
rect 14424 25995 14464 26027
rect 14496 25995 14536 26027
rect 14568 25995 14608 26027
rect 14640 25995 14680 26027
rect 14712 25995 14752 26027
rect 14784 25995 14824 26027
rect 14856 25995 14896 26027
rect 14928 25995 14968 26027
rect 15000 25995 15040 26027
rect 15072 25995 15112 26027
rect 15144 25995 15184 26027
rect 15216 25995 15256 26027
rect 15288 25995 15328 26027
rect 15360 25995 15400 26027
rect 15432 25995 15472 26027
rect 15504 25995 15544 26027
rect 15576 25995 15616 26027
rect 15648 25995 15688 26027
rect 15720 25995 15760 26027
rect 15792 25995 15832 26027
rect 15864 25995 15904 26027
rect 15936 25995 16000 26027
rect 0 25971 16000 25995
rect 0 25931 51 25971
rect 91 25955 149 25971
rect 189 25955 247 25971
rect 287 25955 345 25971
rect 385 25955 443 25971
rect 483 25955 541 25971
rect 581 25955 639 25971
rect 679 25955 737 25971
rect 777 25955 835 25971
rect 875 25955 933 25971
rect 973 25955 1031 25971
rect 1071 25955 1129 25971
rect 1169 25955 16000 25971
rect 0 25923 64 25931
rect 96 25923 136 25955
rect 189 25931 208 25955
rect 168 25923 208 25931
rect 240 25931 247 25955
rect 312 25931 345 25955
rect 385 25931 424 25955
rect 483 25931 496 25955
rect 240 25923 280 25931
rect 312 25923 352 25931
rect 384 25923 424 25931
rect 456 25923 496 25931
rect 528 25931 541 25955
rect 600 25931 639 25955
rect 679 25931 712 25955
rect 777 25931 784 25955
rect 528 25923 568 25931
rect 600 25923 640 25931
rect 672 25923 712 25931
rect 744 25923 784 25931
rect 816 25931 835 25955
rect 816 25923 856 25931
rect 888 25923 928 25955
rect 973 25931 1000 25955
rect 1071 25931 1072 25955
rect 960 25923 1000 25931
rect 1032 25923 1072 25931
rect 1104 25931 1129 25955
rect 1104 25923 1144 25931
rect 1176 25923 1216 25955
rect 1248 25923 1288 25955
rect 1320 25923 1360 25955
rect 1392 25923 1432 25955
rect 1464 25923 1504 25955
rect 1536 25923 1576 25955
rect 1608 25923 1648 25955
rect 1680 25923 1720 25955
rect 1752 25923 1792 25955
rect 1824 25923 1864 25955
rect 1896 25923 1936 25955
rect 1968 25923 2008 25955
rect 2040 25923 2080 25955
rect 2112 25923 2152 25955
rect 2184 25923 2224 25955
rect 2256 25923 2296 25955
rect 2328 25923 2368 25955
rect 2400 25923 2440 25955
rect 2472 25923 2512 25955
rect 2544 25923 2584 25955
rect 2616 25923 2656 25955
rect 2688 25923 2728 25955
rect 2760 25923 2800 25955
rect 2832 25923 2872 25955
rect 2904 25923 2944 25955
rect 2976 25923 3016 25955
rect 3048 25923 3088 25955
rect 3120 25923 3160 25955
rect 3192 25923 3232 25955
rect 3264 25923 3304 25955
rect 3336 25923 3376 25955
rect 3408 25923 3448 25955
rect 3480 25923 3520 25955
rect 3552 25923 3592 25955
rect 3624 25923 3664 25955
rect 3696 25923 3736 25955
rect 3768 25923 3808 25955
rect 3840 25923 3880 25955
rect 3912 25923 3952 25955
rect 3984 25923 4024 25955
rect 4056 25923 4096 25955
rect 4128 25923 4168 25955
rect 4200 25923 4240 25955
rect 4272 25923 4312 25955
rect 4344 25923 4384 25955
rect 4416 25923 4456 25955
rect 4488 25923 4528 25955
rect 4560 25923 4600 25955
rect 4632 25923 4672 25955
rect 4704 25923 4744 25955
rect 4776 25923 4816 25955
rect 4848 25923 4888 25955
rect 4920 25923 4960 25955
rect 4992 25923 5032 25955
rect 5064 25923 5104 25955
rect 5136 25923 5176 25955
rect 5208 25923 5248 25955
rect 5280 25923 5320 25955
rect 5352 25923 5392 25955
rect 5424 25923 5464 25955
rect 5496 25923 5536 25955
rect 5568 25923 5608 25955
rect 5640 25923 5680 25955
rect 5712 25923 5752 25955
rect 5784 25923 5824 25955
rect 5856 25923 5896 25955
rect 5928 25923 5968 25955
rect 6000 25923 6040 25955
rect 6072 25923 6112 25955
rect 6144 25923 6184 25955
rect 6216 25923 6256 25955
rect 6288 25923 6328 25955
rect 6360 25923 6400 25955
rect 6432 25923 6472 25955
rect 6504 25923 6544 25955
rect 6576 25923 6616 25955
rect 6648 25923 6688 25955
rect 6720 25923 6760 25955
rect 6792 25923 6832 25955
rect 6864 25923 6904 25955
rect 6936 25923 6976 25955
rect 7008 25923 7048 25955
rect 7080 25923 7120 25955
rect 7152 25923 7192 25955
rect 7224 25923 7264 25955
rect 7296 25923 7336 25955
rect 7368 25923 7408 25955
rect 7440 25923 7480 25955
rect 7512 25923 7552 25955
rect 7584 25923 7624 25955
rect 7656 25923 7696 25955
rect 7728 25923 7768 25955
rect 7800 25923 7840 25955
rect 7872 25923 7912 25955
rect 7944 25923 7984 25955
rect 8016 25923 8056 25955
rect 8088 25923 8128 25955
rect 8160 25923 8200 25955
rect 8232 25923 8272 25955
rect 8304 25923 8344 25955
rect 8376 25923 8416 25955
rect 8448 25923 8488 25955
rect 8520 25923 8560 25955
rect 8592 25923 8632 25955
rect 8664 25923 8704 25955
rect 8736 25923 8776 25955
rect 8808 25923 8848 25955
rect 8880 25923 8920 25955
rect 8952 25923 8992 25955
rect 9024 25923 9064 25955
rect 9096 25923 9136 25955
rect 9168 25923 9208 25955
rect 9240 25923 9280 25955
rect 9312 25923 9352 25955
rect 9384 25923 9424 25955
rect 9456 25923 9496 25955
rect 9528 25923 9568 25955
rect 9600 25923 9640 25955
rect 9672 25923 9712 25955
rect 9744 25923 9784 25955
rect 9816 25923 9856 25955
rect 9888 25923 9928 25955
rect 9960 25923 10000 25955
rect 10032 25923 10072 25955
rect 10104 25923 10144 25955
rect 10176 25923 10216 25955
rect 10248 25923 10288 25955
rect 10320 25923 10360 25955
rect 10392 25923 10432 25955
rect 10464 25923 10504 25955
rect 10536 25923 10576 25955
rect 10608 25923 10648 25955
rect 10680 25923 10720 25955
rect 10752 25923 10792 25955
rect 10824 25923 10864 25955
rect 10896 25923 10936 25955
rect 10968 25923 11008 25955
rect 11040 25923 11080 25955
rect 11112 25923 11152 25955
rect 11184 25923 11224 25955
rect 11256 25923 11296 25955
rect 11328 25923 11368 25955
rect 11400 25923 11440 25955
rect 11472 25923 11512 25955
rect 11544 25923 11584 25955
rect 11616 25923 11656 25955
rect 11688 25923 11728 25955
rect 11760 25923 11800 25955
rect 11832 25923 11872 25955
rect 11904 25923 11944 25955
rect 11976 25923 12016 25955
rect 12048 25923 12088 25955
rect 12120 25923 12160 25955
rect 12192 25923 12232 25955
rect 12264 25923 12304 25955
rect 12336 25923 12376 25955
rect 12408 25923 12448 25955
rect 12480 25923 12520 25955
rect 12552 25923 12592 25955
rect 12624 25923 12664 25955
rect 12696 25923 12736 25955
rect 12768 25923 12808 25955
rect 12840 25923 12880 25955
rect 12912 25923 12952 25955
rect 12984 25923 13024 25955
rect 13056 25923 13096 25955
rect 13128 25923 13168 25955
rect 13200 25923 13240 25955
rect 13272 25923 13312 25955
rect 13344 25923 13384 25955
rect 13416 25923 13456 25955
rect 13488 25923 13528 25955
rect 13560 25923 13600 25955
rect 13632 25923 13672 25955
rect 13704 25923 13744 25955
rect 13776 25923 13816 25955
rect 13848 25923 13888 25955
rect 13920 25923 13960 25955
rect 13992 25923 14032 25955
rect 14064 25923 14104 25955
rect 14136 25923 14176 25955
rect 14208 25923 14248 25955
rect 14280 25923 14320 25955
rect 14352 25923 14392 25955
rect 14424 25923 14464 25955
rect 14496 25923 14536 25955
rect 14568 25923 14608 25955
rect 14640 25923 14680 25955
rect 14712 25923 14752 25955
rect 14784 25923 14824 25955
rect 14856 25923 14896 25955
rect 14928 25923 14968 25955
rect 15000 25923 15040 25955
rect 15072 25923 15112 25955
rect 15144 25923 15184 25955
rect 15216 25923 15256 25955
rect 15288 25923 15328 25955
rect 15360 25923 15400 25955
rect 15432 25923 15472 25955
rect 15504 25923 15544 25955
rect 15576 25923 15616 25955
rect 15648 25923 15688 25955
rect 15720 25923 15760 25955
rect 15792 25923 15832 25955
rect 15864 25923 15904 25955
rect 15936 25923 16000 25955
rect 0 25883 16000 25923
rect 0 25873 64 25883
rect 0 25833 51 25873
rect 96 25851 136 25883
rect 168 25873 208 25883
rect 189 25851 208 25873
rect 240 25873 280 25883
rect 312 25873 352 25883
rect 384 25873 424 25883
rect 456 25873 496 25883
rect 240 25851 247 25873
rect 312 25851 345 25873
rect 385 25851 424 25873
rect 483 25851 496 25873
rect 528 25873 568 25883
rect 600 25873 640 25883
rect 672 25873 712 25883
rect 744 25873 784 25883
rect 528 25851 541 25873
rect 600 25851 639 25873
rect 679 25851 712 25873
rect 777 25851 784 25873
rect 816 25873 856 25883
rect 816 25851 835 25873
rect 888 25851 928 25883
rect 960 25873 1000 25883
rect 1032 25873 1072 25883
rect 973 25851 1000 25873
rect 1071 25851 1072 25873
rect 1104 25873 1144 25883
rect 1104 25851 1129 25873
rect 1176 25851 1216 25883
rect 1248 25851 1288 25883
rect 1320 25851 1360 25883
rect 1392 25851 1432 25883
rect 1464 25851 1504 25883
rect 1536 25851 1576 25883
rect 1608 25851 1648 25883
rect 1680 25851 1720 25883
rect 1752 25851 1792 25883
rect 1824 25851 1864 25883
rect 1896 25851 1936 25883
rect 1968 25851 2008 25883
rect 2040 25851 2080 25883
rect 2112 25851 2152 25883
rect 2184 25851 2224 25883
rect 2256 25851 2296 25883
rect 2328 25851 2368 25883
rect 2400 25851 2440 25883
rect 2472 25851 2512 25883
rect 2544 25851 2584 25883
rect 2616 25851 2656 25883
rect 2688 25851 2728 25883
rect 2760 25851 2800 25883
rect 2832 25851 2872 25883
rect 2904 25851 2944 25883
rect 2976 25851 3016 25883
rect 3048 25851 3088 25883
rect 3120 25851 3160 25883
rect 3192 25851 3232 25883
rect 3264 25851 3304 25883
rect 3336 25851 3376 25883
rect 3408 25851 3448 25883
rect 3480 25851 3520 25883
rect 3552 25851 3592 25883
rect 3624 25851 3664 25883
rect 3696 25851 3736 25883
rect 3768 25851 3808 25883
rect 3840 25851 3880 25883
rect 3912 25851 3952 25883
rect 3984 25851 4024 25883
rect 4056 25851 4096 25883
rect 4128 25851 4168 25883
rect 4200 25851 4240 25883
rect 4272 25851 4312 25883
rect 4344 25851 4384 25883
rect 4416 25851 4456 25883
rect 4488 25851 4528 25883
rect 4560 25851 4600 25883
rect 4632 25851 4672 25883
rect 4704 25851 4744 25883
rect 4776 25851 4816 25883
rect 4848 25851 4888 25883
rect 4920 25851 4960 25883
rect 4992 25851 5032 25883
rect 5064 25851 5104 25883
rect 5136 25851 5176 25883
rect 5208 25851 5248 25883
rect 5280 25851 5320 25883
rect 5352 25851 5392 25883
rect 5424 25851 5464 25883
rect 5496 25851 5536 25883
rect 5568 25851 5608 25883
rect 5640 25851 5680 25883
rect 5712 25851 5752 25883
rect 5784 25851 5824 25883
rect 5856 25851 5896 25883
rect 5928 25851 5968 25883
rect 6000 25851 6040 25883
rect 6072 25851 6112 25883
rect 6144 25851 6184 25883
rect 6216 25851 6256 25883
rect 6288 25851 6328 25883
rect 6360 25851 6400 25883
rect 6432 25851 6472 25883
rect 6504 25851 6544 25883
rect 6576 25851 6616 25883
rect 6648 25851 6688 25883
rect 6720 25851 6760 25883
rect 6792 25851 6832 25883
rect 6864 25851 6904 25883
rect 6936 25851 6976 25883
rect 7008 25851 7048 25883
rect 7080 25851 7120 25883
rect 7152 25851 7192 25883
rect 7224 25851 7264 25883
rect 7296 25851 7336 25883
rect 7368 25851 7408 25883
rect 7440 25851 7480 25883
rect 7512 25851 7552 25883
rect 7584 25851 7624 25883
rect 7656 25851 7696 25883
rect 7728 25851 7768 25883
rect 7800 25851 7840 25883
rect 7872 25851 7912 25883
rect 7944 25851 7984 25883
rect 8016 25851 8056 25883
rect 8088 25851 8128 25883
rect 8160 25851 8200 25883
rect 8232 25851 8272 25883
rect 8304 25851 8344 25883
rect 8376 25851 8416 25883
rect 8448 25851 8488 25883
rect 8520 25851 8560 25883
rect 8592 25851 8632 25883
rect 8664 25851 8704 25883
rect 8736 25851 8776 25883
rect 8808 25851 8848 25883
rect 8880 25851 8920 25883
rect 8952 25851 8992 25883
rect 9024 25851 9064 25883
rect 9096 25851 9136 25883
rect 9168 25851 9208 25883
rect 9240 25851 9280 25883
rect 9312 25851 9352 25883
rect 9384 25851 9424 25883
rect 9456 25851 9496 25883
rect 9528 25851 9568 25883
rect 9600 25851 9640 25883
rect 9672 25851 9712 25883
rect 9744 25851 9784 25883
rect 9816 25851 9856 25883
rect 9888 25851 9928 25883
rect 9960 25851 10000 25883
rect 10032 25851 10072 25883
rect 10104 25851 10144 25883
rect 10176 25851 10216 25883
rect 10248 25851 10288 25883
rect 10320 25851 10360 25883
rect 10392 25851 10432 25883
rect 10464 25851 10504 25883
rect 10536 25851 10576 25883
rect 10608 25851 10648 25883
rect 10680 25851 10720 25883
rect 10752 25851 10792 25883
rect 10824 25851 10864 25883
rect 10896 25851 10936 25883
rect 10968 25851 11008 25883
rect 11040 25851 11080 25883
rect 11112 25851 11152 25883
rect 11184 25851 11224 25883
rect 11256 25851 11296 25883
rect 11328 25851 11368 25883
rect 11400 25851 11440 25883
rect 11472 25851 11512 25883
rect 11544 25851 11584 25883
rect 11616 25851 11656 25883
rect 11688 25851 11728 25883
rect 11760 25851 11800 25883
rect 11832 25851 11872 25883
rect 11904 25851 11944 25883
rect 11976 25851 12016 25883
rect 12048 25851 12088 25883
rect 12120 25851 12160 25883
rect 12192 25851 12232 25883
rect 12264 25851 12304 25883
rect 12336 25851 12376 25883
rect 12408 25851 12448 25883
rect 12480 25851 12520 25883
rect 12552 25851 12592 25883
rect 12624 25851 12664 25883
rect 12696 25851 12736 25883
rect 12768 25851 12808 25883
rect 12840 25851 12880 25883
rect 12912 25851 12952 25883
rect 12984 25851 13024 25883
rect 13056 25851 13096 25883
rect 13128 25851 13168 25883
rect 13200 25851 13240 25883
rect 13272 25851 13312 25883
rect 13344 25851 13384 25883
rect 13416 25851 13456 25883
rect 13488 25851 13528 25883
rect 13560 25851 13600 25883
rect 13632 25851 13672 25883
rect 13704 25851 13744 25883
rect 13776 25851 13816 25883
rect 13848 25851 13888 25883
rect 13920 25851 13960 25883
rect 13992 25851 14032 25883
rect 14064 25851 14104 25883
rect 14136 25851 14176 25883
rect 14208 25851 14248 25883
rect 14280 25851 14320 25883
rect 14352 25851 14392 25883
rect 14424 25851 14464 25883
rect 14496 25851 14536 25883
rect 14568 25851 14608 25883
rect 14640 25851 14680 25883
rect 14712 25851 14752 25883
rect 14784 25851 14824 25883
rect 14856 25851 14896 25883
rect 14928 25851 14968 25883
rect 15000 25851 15040 25883
rect 15072 25851 15112 25883
rect 15144 25851 15184 25883
rect 15216 25851 15256 25883
rect 15288 25851 15328 25883
rect 15360 25851 15400 25883
rect 15432 25851 15472 25883
rect 15504 25851 15544 25883
rect 15576 25851 15616 25883
rect 15648 25851 15688 25883
rect 15720 25851 15760 25883
rect 15792 25851 15832 25883
rect 15864 25851 15904 25883
rect 15936 25851 16000 25883
rect 91 25833 149 25851
rect 189 25833 247 25851
rect 287 25833 345 25851
rect 385 25833 443 25851
rect 483 25833 541 25851
rect 581 25833 639 25851
rect 679 25833 737 25851
rect 777 25833 835 25851
rect 875 25833 933 25851
rect 973 25833 1031 25851
rect 1071 25833 1129 25851
rect 1169 25833 16000 25851
rect 0 25811 16000 25833
rect 0 25779 64 25811
rect 96 25779 136 25811
rect 168 25779 208 25811
rect 240 25779 280 25811
rect 312 25779 352 25811
rect 384 25779 424 25811
rect 456 25779 496 25811
rect 528 25779 568 25811
rect 600 25779 640 25811
rect 672 25779 712 25811
rect 744 25779 784 25811
rect 816 25779 856 25811
rect 888 25779 928 25811
rect 960 25779 1000 25811
rect 1032 25779 1072 25811
rect 1104 25779 1144 25811
rect 1176 25779 1216 25811
rect 1248 25779 1288 25811
rect 1320 25779 1360 25811
rect 1392 25779 1432 25811
rect 1464 25779 1504 25811
rect 1536 25779 1576 25811
rect 1608 25779 1648 25811
rect 1680 25779 1720 25811
rect 1752 25779 1792 25811
rect 1824 25779 1864 25811
rect 1896 25779 1936 25811
rect 1968 25779 2008 25811
rect 2040 25779 2080 25811
rect 2112 25779 2152 25811
rect 2184 25779 2224 25811
rect 2256 25779 2296 25811
rect 2328 25779 2368 25811
rect 2400 25779 2440 25811
rect 2472 25779 2512 25811
rect 2544 25779 2584 25811
rect 2616 25779 2656 25811
rect 2688 25779 2728 25811
rect 2760 25779 2800 25811
rect 2832 25779 2872 25811
rect 2904 25779 2944 25811
rect 2976 25779 3016 25811
rect 3048 25779 3088 25811
rect 3120 25779 3160 25811
rect 3192 25779 3232 25811
rect 3264 25779 3304 25811
rect 3336 25779 3376 25811
rect 3408 25779 3448 25811
rect 3480 25779 3520 25811
rect 3552 25779 3592 25811
rect 3624 25779 3664 25811
rect 3696 25779 3736 25811
rect 3768 25779 3808 25811
rect 3840 25779 3880 25811
rect 3912 25779 3952 25811
rect 3984 25779 4024 25811
rect 4056 25779 4096 25811
rect 4128 25779 4168 25811
rect 4200 25779 4240 25811
rect 4272 25779 4312 25811
rect 4344 25779 4384 25811
rect 4416 25779 4456 25811
rect 4488 25779 4528 25811
rect 4560 25779 4600 25811
rect 4632 25779 4672 25811
rect 4704 25779 4744 25811
rect 4776 25779 4816 25811
rect 4848 25779 4888 25811
rect 4920 25779 4960 25811
rect 4992 25779 5032 25811
rect 5064 25779 5104 25811
rect 5136 25779 5176 25811
rect 5208 25779 5248 25811
rect 5280 25779 5320 25811
rect 5352 25779 5392 25811
rect 5424 25779 5464 25811
rect 5496 25779 5536 25811
rect 5568 25779 5608 25811
rect 5640 25779 5680 25811
rect 5712 25779 5752 25811
rect 5784 25779 5824 25811
rect 5856 25779 5896 25811
rect 5928 25779 5968 25811
rect 6000 25779 6040 25811
rect 6072 25779 6112 25811
rect 6144 25779 6184 25811
rect 6216 25779 6256 25811
rect 6288 25779 6328 25811
rect 6360 25779 6400 25811
rect 6432 25779 6472 25811
rect 6504 25779 6544 25811
rect 6576 25779 6616 25811
rect 6648 25779 6688 25811
rect 6720 25779 6760 25811
rect 6792 25779 6832 25811
rect 6864 25779 6904 25811
rect 6936 25779 6976 25811
rect 7008 25779 7048 25811
rect 7080 25779 7120 25811
rect 7152 25779 7192 25811
rect 7224 25779 7264 25811
rect 7296 25779 7336 25811
rect 7368 25779 7408 25811
rect 7440 25779 7480 25811
rect 7512 25779 7552 25811
rect 7584 25779 7624 25811
rect 7656 25779 7696 25811
rect 7728 25779 7768 25811
rect 7800 25779 7840 25811
rect 7872 25779 7912 25811
rect 7944 25779 7984 25811
rect 8016 25779 8056 25811
rect 8088 25779 8128 25811
rect 8160 25779 8200 25811
rect 8232 25779 8272 25811
rect 8304 25779 8344 25811
rect 8376 25779 8416 25811
rect 8448 25779 8488 25811
rect 8520 25779 8560 25811
rect 8592 25779 8632 25811
rect 8664 25779 8704 25811
rect 8736 25779 8776 25811
rect 8808 25779 8848 25811
rect 8880 25779 8920 25811
rect 8952 25779 8992 25811
rect 9024 25779 9064 25811
rect 9096 25779 9136 25811
rect 9168 25779 9208 25811
rect 9240 25779 9280 25811
rect 9312 25779 9352 25811
rect 9384 25779 9424 25811
rect 9456 25779 9496 25811
rect 9528 25779 9568 25811
rect 9600 25779 9640 25811
rect 9672 25779 9712 25811
rect 9744 25779 9784 25811
rect 9816 25779 9856 25811
rect 9888 25779 9928 25811
rect 9960 25779 10000 25811
rect 10032 25779 10072 25811
rect 10104 25779 10144 25811
rect 10176 25779 10216 25811
rect 10248 25779 10288 25811
rect 10320 25779 10360 25811
rect 10392 25779 10432 25811
rect 10464 25779 10504 25811
rect 10536 25779 10576 25811
rect 10608 25779 10648 25811
rect 10680 25779 10720 25811
rect 10752 25779 10792 25811
rect 10824 25779 10864 25811
rect 10896 25779 10936 25811
rect 10968 25779 11008 25811
rect 11040 25779 11080 25811
rect 11112 25779 11152 25811
rect 11184 25779 11224 25811
rect 11256 25779 11296 25811
rect 11328 25779 11368 25811
rect 11400 25779 11440 25811
rect 11472 25779 11512 25811
rect 11544 25779 11584 25811
rect 11616 25779 11656 25811
rect 11688 25779 11728 25811
rect 11760 25779 11800 25811
rect 11832 25779 11872 25811
rect 11904 25779 11944 25811
rect 11976 25779 12016 25811
rect 12048 25779 12088 25811
rect 12120 25779 12160 25811
rect 12192 25779 12232 25811
rect 12264 25779 12304 25811
rect 12336 25779 12376 25811
rect 12408 25779 12448 25811
rect 12480 25779 12520 25811
rect 12552 25779 12592 25811
rect 12624 25779 12664 25811
rect 12696 25779 12736 25811
rect 12768 25779 12808 25811
rect 12840 25779 12880 25811
rect 12912 25779 12952 25811
rect 12984 25779 13024 25811
rect 13056 25779 13096 25811
rect 13128 25779 13168 25811
rect 13200 25779 13240 25811
rect 13272 25779 13312 25811
rect 13344 25779 13384 25811
rect 13416 25779 13456 25811
rect 13488 25779 13528 25811
rect 13560 25779 13600 25811
rect 13632 25779 13672 25811
rect 13704 25779 13744 25811
rect 13776 25779 13816 25811
rect 13848 25779 13888 25811
rect 13920 25779 13960 25811
rect 13992 25779 14032 25811
rect 14064 25779 14104 25811
rect 14136 25779 14176 25811
rect 14208 25779 14248 25811
rect 14280 25779 14320 25811
rect 14352 25779 14392 25811
rect 14424 25779 14464 25811
rect 14496 25779 14536 25811
rect 14568 25779 14608 25811
rect 14640 25779 14680 25811
rect 14712 25779 14752 25811
rect 14784 25779 14824 25811
rect 14856 25779 14896 25811
rect 14928 25779 14968 25811
rect 15000 25779 15040 25811
rect 15072 25779 15112 25811
rect 15144 25779 15184 25811
rect 15216 25779 15256 25811
rect 15288 25779 15328 25811
rect 15360 25779 15400 25811
rect 15432 25779 15472 25811
rect 15504 25779 15544 25811
rect 15576 25779 15616 25811
rect 15648 25779 15688 25811
rect 15720 25779 15760 25811
rect 15792 25779 15832 25811
rect 15864 25779 15904 25811
rect 15936 25779 16000 25811
rect 0 25775 16000 25779
rect 0 25735 51 25775
rect 91 25739 149 25775
rect 189 25739 247 25775
rect 287 25739 345 25775
rect 385 25739 443 25775
rect 483 25739 541 25775
rect 581 25739 639 25775
rect 679 25739 737 25775
rect 777 25739 835 25775
rect 875 25739 933 25775
rect 973 25739 1031 25775
rect 1071 25739 1129 25775
rect 1169 25739 16000 25775
rect 0 25707 64 25735
rect 96 25707 136 25739
rect 189 25735 208 25739
rect 168 25707 208 25735
rect 240 25735 247 25739
rect 312 25735 345 25739
rect 385 25735 424 25739
rect 483 25735 496 25739
rect 240 25707 280 25735
rect 312 25707 352 25735
rect 384 25707 424 25735
rect 456 25707 496 25735
rect 528 25735 541 25739
rect 600 25735 639 25739
rect 679 25735 712 25739
rect 777 25735 784 25739
rect 528 25707 568 25735
rect 600 25707 640 25735
rect 672 25707 712 25735
rect 744 25707 784 25735
rect 816 25735 835 25739
rect 816 25707 856 25735
rect 888 25707 928 25739
rect 973 25735 1000 25739
rect 1071 25735 1072 25739
rect 960 25707 1000 25735
rect 1032 25707 1072 25735
rect 1104 25735 1129 25739
rect 1104 25707 1144 25735
rect 1176 25707 1216 25739
rect 1248 25707 1288 25739
rect 1320 25707 1360 25739
rect 1392 25707 1432 25739
rect 1464 25707 1504 25739
rect 1536 25707 1576 25739
rect 1608 25707 1648 25739
rect 1680 25707 1720 25739
rect 1752 25707 1792 25739
rect 1824 25707 1864 25739
rect 1896 25707 1936 25739
rect 1968 25707 2008 25739
rect 2040 25707 2080 25739
rect 2112 25707 2152 25739
rect 2184 25707 2224 25739
rect 2256 25707 2296 25739
rect 2328 25707 2368 25739
rect 2400 25707 2440 25739
rect 2472 25707 2512 25739
rect 2544 25707 2584 25739
rect 2616 25707 2656 25739
rect 2688 25707 2728 25739
rect 2760 25707 2800 25739
rect 2832 25707 2872 25739
rect 2904 25707 2944 25739
rect 2976 25707 3016 25739
rect 3048 25707 3088 25739
rect 3120 25707 3160 25739
rect 3192 25707 3232 25739
rect 3264 25707 3304 25739
rect 3336 25707 3376 25739
rect 3408 25707 3448 25739
rect 3480 25707 3520 25739
rect 3552 25707 3592 25739
rect 3624 25707 3664 25739
rect 3696 25707 3736 25739
rect 3768 25707 3808 25739
rect 3840 25707 3880 25739
rect 3912 25707 3952 25739
rect 3984 25707 4024 25739
rect 4056 25707 4096 25739
rect 4128 25707 4168 25739
rect 4200 25707 4240 25739
rect 4272 25707 4312 25739
rect 4344 25707 4384 25739
rect 4416 25707 4456 25739
rect 4488 25707 4528 25739
rect 4560 25707 4600 25739
rect 4632 25707 4672 25739
rect 4704 25707 4744 25739
rect 4776 25707 4816 25739
rect 4848 25707 4888 25739
rect 4920 25707 4960 25739
rect 4992 25707 5032 25739
rect 5064 25707 5104 25739
rect 5136 25707 5176 25739
rect 5208 25707 5248 25739
rect 5280 25707 5320 25739
rect 5352 25707 5392 25739
rect 5424 25707 5464 25739
rect 5496 25707 5536 25739
rect 5568 25707 5608 25739
rect 5640 25707 5680 25739
rect 5712 25707 5752 25739
rect 5784 25707 5824 25739
rect 5856 25707 5896 25739
rect 5928 25707 5968 25739
rect 6000 25707 6040 25739
rect 6072 25707 6112 25739
rect 6144 25707 6184 25739
rect 6216 25707 6256 25739
rect 6288 25707 6328 25739
rect 6360 25707 6400 25739
rect 6432 25707 6472 25739
rect 6504 25707 6544 25739
rect 6576 25707 6616 25739
rect 6648 25707 6688 25739
rect 6720 25707 6760 25739
rect 6792 25707 6832 25739
rect 6864 25707 6904 25739
rect 6936 25707 6976 25739
rect 7008 25707 7048 25739
rect 7080 25707 7120 25739
rect 7152 25707 7192 25739
rect 7224 25707 7264 25739
rect 7296 25707 7336 25739
rect 7368 25707 7408 25739
rect 7440 25707 7480 25739
rect 7512 25707 7552 25739
rect 7584 25707 7624 25739
rect 7656 25707 7696 25739
rect 7728 25707 7768 25739
rect 7800 25707 7840 25739
rect 7872 25707 7912 25739
rect 7944 25707 7984 25739
rect 8016 25707 8056 25739
rect 8088 25707 8128 25739
rect 8160 25707 8200 25739
rect 8232 25707 8272 25739
rect 8304 25707 8344 25739
rect 8376 25707 8416 25739
rect 8448 25707 8488 25739
rect 8520 25707 8560 25739
rect 8592 25707 8632 25739
rect 8664 25707 8704 25739
rect 8736 25707 8776 25739
rect 8808 25707 8848 25739
rect 8880 25707 8920 25739
rect 8952 25707 8992 25739
rect 9024 25707 9064 25739
rect 9096 25707 9136 25739
rect 9168 25707 9208 25739
rect 9240 25707 9280 25739
rect 9312 25707 9352 25739
rect 9384 25707 9424 25739
rect 9456 25707 9496 25739
rect 9528 25707 9568 25739
rect 9600 25707 9640 25739
rect 9672 25707 9712 25739
rect 9744 25707 9784 25739
rect 9816 25707 9856 25739
rect 9888 25707 9928 25739
rect 9960 25707 10000 25739
rect 10032 25707 10072 25739
rect 10104 25707 10144 25739
rect 10176 25707 10216 25739
rect 10248 25707 10288 25739
rect 10320 25707 10360 25739
rect 10392 25707 10432 25739
rect 10464 25707 10504 25739
rect 10536 25707 10576 25739
rect 10608 25707 10648 25739
rect 10680 25707 10720 25739
rect 10752 25707 10792 25739
rect 10824 25707 10864 25739
rect 10896 25707 10936 25739
rect 10968 25707 11008 25739
rect 11040 25707 11080 25739
rect 11112 25707 11152 25739
rect 11184 25707 11224 25739
rect 11256 25707 11296 25739
rect 11328 25707 11368 25739
rect 11400 25707 11440 25739
rect 11472 25707 11512 25739
rect 11544 25707 11584 25739
rect 11616 25707 11656 25739
rect 11688 25707 11728 25739
rect 11760 25707 11800 25739
rect 11832 25707 11872 25739
rect 11904 25707 11944 25739
rect 11976 25707 12016 25739
rect 12048 25707 12088 25739
rect 12120 25707 12160 25739
rect 12192 25707 12232 25739
rect 12264 25707 12304 25739
rect 12336 25707 12376 25739
rect 12408 25707 12448 25739
rect 12480 25707 12520 25739
rect 12552 25707 12592 25739
rect 12624 25707 12664 25739
rect 12696 25707 12736 25739
rect 12768 25707 12808 25739
rect 12840 25707 12880 25739
rect 12912 25707 12952 25739
rect 12984 25707 13024 25739
rect 13056 25707 13096 25739
rect 13128 25707 13168 25739
rect 13200 25707 13240 25739
rect 13272 25707 13312 25739
rect 13344 25707 13384 25739
rect 13416 25707 13456 25739
rect 13488 25707 13528 25739
rect 13560 25707 13600 25739
rect 13632 25707 13672 25739
rect 13704 25707 13744 25739
rect 13776 25707 13816 25739
rect 13848 25707 13888 25739
rect 13920 25707 13960 25739
rect 13992 25707 14032 25739
rect 14064 25707 14104 25739
rect 14136 25707 14176 25739
rect 14208 25707 14248 25739
rect 14280 25707 14320 25739
rect 14352 25707 14392 25739
rect 14424 25707 14464 25739
rect 14496 25707 14536 25739
rect 14568 25707 14608 25739
rect 14640 25707 14680 25739
rect 14712 25707 14752 25739
rect 14784 25707 14824 25739
rect 14856 25707 14896 25739
rect 14928 25707 14968 25739
rect 15000 25707 15040 25739
rect 15072 25707 15112 25739
rect 15144 25707 15184 25739
rect 15216 25707 15256 25739
rect 15288 25707 15328 25739
rect 15360 25707 15400 25739
rect 15432 25707 15472 25739
rect 15504 25707 15544 25739
rect 15576 25707 15616 25739
rect 15648 25707 15688 25739
rect 15720 25707 15760 25739
rect 15792 25707 15832 25739
rect 15864 25707 15904 25739
rect 15936 25707 16000 25739
rect 0 25677 16000 25707
rect 0 25637 51 25677
rect 91 25667 149 25677
rect 189 25667 247 25677
rect 287 25667 345 25677
rect 385 25667 443 25677
rect 483 25667 541 25677
rect 581 25667 639 25677
rect 679 25667 737 25677
rect 777 25667 835 25677
rect 875 25667 933 25677
rect 973 25667 1031 25677
rect 1071 25667 1129 25677
rect 1169 25667 16000 25677
rect 0 25635 64 25637
rect 96 25635 136 25667
rect 189 25637 208 25667
rect 168 25635 208 25637
rect 240 25637 247 25667
rect 312 25637 345 25667
rect 385 25637 424 25667
rect 483 25637 496 25667
rect 240 25635 280 25637
rect 312 25635 352 25637
rect 384 25635 424 25637
rect 456 25635 496 25637
rect 528 25637 541 25667
rect 600 25637 639 25667
rect 679 25637 712 25667
rect 777 25637 784 25667
rect 528 25635 568 25637
rect 600 25635 640 25637
rect 672 25635 712 25637
rect 744 25635 784 25637
rect 816 25637 835 25667
rect 816 25635 856 25637
rect 888 25635 928 25667
rect 973 25637 1000 25667
rect 1071 25637 1072 25667
rect 960 25635 1000 25637
rect 1032 25635 1072 25637
rect 1104 25637 1129 25667
rect 1104 25635 1144 25637
rect 1176 25635 1216 25667
rect 1248 25635 1288 25667
rect 1320 25635 1360 25667
rect 1392 25635 1432 25667
rect 1464 25635 1504 25667
rect 1536 25635 1576 25667
rect 1608 25635 1648 25667
rect 1680 25635 1720 25667
rect 1752 25635 1792 25667
rect 1824 25635 1864 25667
rect 1896 25635 1936 25667
rect 1968 25635 2008 25667
rect 2040 25635 2080 25667
rect 2112 25635 2152 25667
rect 2184 25635 2224 25667
rect 2256 25635 2296 25667
rect 2328 25635 2368 25667
rect 2400 25635 2440 25667
rect 2472 25635 2512 25667
rect 2544 25635 2584 25667
rect 2616 25635 2656 25667
rect 2688 25635 2728 25667
rect 2760 25635 2800 25667
rect 2832 25635 2872 25667
rect 2904 25635 2944 25667
rect 2976 25635 3016 25667
rect 3048 25635 3088 25667
rect 3120 25635 3160 25667
rect 3192 25635 3232 25667
rect 3264 25635 3304 25667
rect 3336 25635 3376 25667
rect 3408 25635 3448 25667
rect 3480 25635 3520 25667
rect 3552 25635 3592 25667
rect 3624 25635 3664 25667
rect 3696 25635 3736 25667
rect 3768 25635 3808 25667
rect 3840 25635 3880 25667
rect 3912 25635 3952 25667
rect 3984 25635 4024 25667
rect 4056 25635 4096 25667
rect 4128 25635 4168 25667
rect 4200 25635 4240 25667
rect 4272 25635 4312 25667
rect 4344 25635 4384 25667
rect 4416 25635 4456 25667
rect 4488 25635 4528 25667
rect 4560 25635 4600 25667
rect 4632 25635 4672 25667
rect 4704 25635 4744 25667
rect 4776 25635 4816 25667
rect 4848 25635 4888 25667
rect 4920 25635 4960 25667
rect 4992 25635 5032 25667
rect 5064 25635 5104 25667
rect 5136 25635 5176 25667
rect 5208 25635 5248 25667
rect 5280 25635 5320 25667
rect 5352 25635 5392 25667
rect 5424 25635 5464 25667
rect 5496 25635 5536 25667
rect 5568 25635 5608 25667
rect 5640 25635 5680 25667
rect 5712 25635 5752 25667
rect 5784 25635 5824 25667
rect 5856 25635 5896 25667
rect 5928 25635 5968 25667
rect 6000 25635 6040 25667
rect 6072 25635 6112 25667
rect 6144 25635 6184 25667
rect 6216 25635 6256 25667
rect 6288 25635 6328 25667
rect 6360 25635 6400 25667
rect 6432 25635 6472 25667
rect 6504 25635 6544 25667
rect 6576 25635 6616 25667
rect 6648 25635 6688 25667
rect 6720 25635 6760 25667
rect 6792 25635 6832 25667
rect 6864 25635 6904 25667
rect 6936 25635 6976 25667
rect 7008 25635 7048 25667
rect 7080 25635 7120 25667
rect 7152 25635 7192 25667
rect 7224 25635 7264 25667
rect 7296 25635 7336 25667
rect 7368 25635 7408 25667
rect 7440 25635 7480 25667
rect 7512 25635 7552 25667
rect 7584 25635 7624 25667
rect 7656 25635 7696 25667
rect 7728 25635 7768 25667
rect 7800 25635 7840 25667
rect 7872 25635 7912 25667
rect 7944 25635 7984 25667
rect 8016 25635 8056 25667
rect 8088 25635 8128 25667
rect 8160 25635 8200 25667
rect 8232 25635 8272 25667
rect 8304 25635 8344 25667
rect 8376 25635 8416 25667
rect 8448 25635 8488 25667
rect 8520 25635 8560 25667
rect 8592 25635 8632 25667
rect 8664 25635 8704 25667
rect 8736 25635 8776 25667
rect 8808 25635 8848 25667
rect 8880 25635 8920 25667
rect 8952 25635 8992 25667
rect 9024 25635 9064 25667
rect 9096 25635 9136 25667
rect 9168 25635 9208 25667
rect 9240 25635 9280 25667
rect 9312 25635 9352 25667
rect 9384 25635 9424 25667
rect 9456 25635 9496 25667
rect 9528 25635 9568 25667
rect 9600 25635 9640 25667
rect 9672 25635 9712 25667
rect 9744 25635 9784 25667
rect 9816 25635 9856 25667
rect 9888 25635 9928 25667
rect 9960 25635 10000 25667
rect 10032 25635 10072 25667
rect 10104 25635 10144 25667
rect 10176 25635 10216 25667
rect 10248 25635 10288 25667
rect 10320 25635 10360 25667
rect 10392 25635 10432 25667
rect 10464 25635 10504 25667
rect 10536 25635 10576 25667
rect 10608 25635 10648 25667
rect 10680 25635 10720 25667
rect 10752 25635 10792 25667
rect 10824 25635 10864 25667
rect 10896 25635 10936 25667
rect 10968 25635 11008 25667
rect 11040 25635 11080 25667
rect 11112 25635 11152 25667
rect 11184 25635 11224 25667
rect 11256 25635 11296 25667
rect 11328 25635 11368 25667
rect 11400 25635 11440 25667
rect 11472 25635 11512 25667
rect 11544 25635 11584 25667
rect 11616 25635 11656 25667
rect 11688 25635 11728 25667
rect 11760 25635 11800 25667
rect 11832 25635 11872 25667
rect 11904 25635 11944 25667
rect 11976 25635 12016 25667
rect 12048 25635 12088 25667
rect 12120 25635 12160 25667
rect 12192 25635 12232 25667
rect 12264 25635 12304 25667
rect 12336 25635 12376 25667
rect 12408 25635 12448 25667
rect 12480 25635 12520 25667
rect 12552 25635 12592 25667
rect 12624 25635 12664 25667
rect 12696 25635 12736 25667
rect 12768 25635 12808 25667
rect 12840 25635 12880 25667
rect 12912 25635 12952 25667
rect 12984 25635 13024 25667
rect 13056 25635 13096 25667
rect 13128 25635 13168 25667
rect 13200 25635 13240 25667
rect 13272 25635 13312 25667
rect 13344 25635 13384 25667
rect 13416 25635 13456 25667
rect 13488 25635 13528 25667
rect 13560 25635 13600 25667
rect 13632 25635 13672 25667
rect 13704 25635 13744 25667
rect 13776 25635 13816 25667
rect 13848 25635 13888 25667
rect 13920 25635 13960 25667
rect 13992 25635 14032 25667
rect 14064 25635 14104 25667
rect 14136 25635 14176 25667
rect 14208 25635 14248 25667
rect 14280 25635 14320 25667
rect 14352 25635 14392 25667
rect 14424 25635 14464 25667
rect 14496 25635 14536 25667
rect 14568 25635 14608 25667
rect 14640 25635 14680 25667
rect 14712 25635 14752 25667
rect 14784 25635 14824 25667
rect 14856 25635 14896 25667
rect 14928 25635 14968 25667
rect 15000 25635 15040 25667
rect 15072 25635 15112 25667
rect 15144 25635 15184 25667
rect 15216 25635 15256 25667
rect 15288 25635 15328 25667
rect 15360 25635 15400 25667
rect 15432 25635 15472 25667
rect 15504 25635 15544 25667
rect 15576 25635 15616 25667
rect 15648 25635 15688 25667
rect 15720 25635 15760 25667
rect 15792 25635 15832 25667
rect 15864 25635 15904 25667
rect 15936 25635 16000 25667
rect 0 25595 16000 25635
rect 0 25579 64 25595
rect 0 25539 51 25579
rect 96 25563 136 25595
rect 168 25579 208 25595
rect 189 25563 208 25579
rect 240 25579 280 25595
rect 312 25579 352 25595
rect 384 25579 424 25595
rect 456 25579 496 25595
rect 240 25563 247 25579
rect 312 25563 345 25579
rect 385 25563 424 25579
rect 483 25563 496 25579
rect 528 25579 568 25595
rect 600 25579 640 25595
rect 672 25579 712 25595
rect 744 25579 784 25595
rect 528 25563 541 25579
rect 600 25563 639 25579
rect 679 25563 712 25579
rect 777 25563 784 25579
rect 816 25579 856 25595
rect 816 25563 835 25579
rect 888 25563 928 25595
rect 960 25579 1000 25595
rect 1032 25579 1072 25595
rect 973 25563 1000 25579
rect 1071 25563 1072 25579
rect 1104 25579 1144 25595
rect 1104 25563 1129 25579
rect 1176 25563 1216 25595
rect 1248 25563 1288 25595
rect 1320 25563 1360 25595
rect 1392 25563 1432 25595
rect 1464 25563 1504 25595
rect 1536 25563 1576 25595
rect 1608 25563 1648 25595
rect 1680 25563 1720 25595
rect 1752 25563 1792 25595
rect 1824 25563 1864 25595
rect 1896 25563 1936 25595
rect 1968 25563 2008 25595
rect 2040 25563 2080 25595
rect 2112 25563 2152 25595
rect 2184 25563 2224 25595
rect 2256 25563 2296 25595
rect 2328 25563 2368 25595
rect 2400 25563 2440 25595
rect 2472 25563 2512 25595
rect 2544 25563 2584 25595
rect 2616 25563 2656 25595
rect 2688 25563 2728 25595
rect 2760 25563 2800 25595
rect 2832 25563 2872 25595
rect 2904 25563 2944 25595
rect 2976 25563 3016 25595
rect 3048 25563 3088 25595
rect 3120 25563 3160 25595
rect 3192 25563 3232 25595
rect 3264 25563 3304 25595
rect 3336 25563 3376 25595
rect 3408 25563 3448 25595
rect 3480 25563 3520 25595
rect 3552 25563 3592 25595
rect 3624 25563 3664 25595
rect 3696 25563 3736 25595
rect 3768 25563 3808 25595
rect 3840 25563 3880 25595
rect 3912 25563 3952 25595
rect 3984 25563 4024 25595
rect 4056 25563 4096 25595
rect 4128 25563 4168 25595
rect 4200 25563 4240 25595
rect 4272 25563 4312 25595
rect 4344 25563 4384 25595
rect 4416 25563 4456 25595
rect 4488 25563 4528 25595
rect 4560 25563 4600 25595
rect 4632 25563 4672 25595
rect 4704 25563 4744 25595
rect 4776 25563 4816 25595
rect 4848 25563 4888 25595
rect 4920 25563 4960 25595
rect 4992 25563 5032 25595
rect 5064 25563 5104 25595
rect 5136 25563 5176 25595
rect 5208 25563 5248 25595
rect 5280 25563 5320 25595
rect 5352 25563 5392 25595
rect 5424 25563 5464 25595
rect 5496 25563 5536 25595
rect 5568 25563 5608 25595
rect 5640 25563 5680 25595
rect 5712 25563 5752 25595
rect 5784 25563 5824 25595
rect 5856 25563 5896 25595
rect 5928 25563 5968 25595
rect 6000 25563 6040 25595
rect 6072 25563 6112 25595
rect 6144 25563 6184 25595
rect 6216 25563 6256 25595
rect 6288 25563 6328 25595
rect 6360 25563 6400 25595
rect 6432 25563 6472 25595
rect 6504 25563 6544 25595
rect 6576 25563 6616 25595
rect 6648 25563 6688 25595
rect 6720 25563 6760 25595
rect 6792 25563 6832 25595
rect 6864 25563 6904 25595
rect 6936 25563 6976 25595
rect 7008 25563 7048 25595
rect 7080 25563 7120 25595
rect 7152 25563 7192 25595
rect 7224 25563 7264 25595
rect 7296 25563 7336 25595
rect 7368 25563 7408 25595
rect 7440 25563 7480 25595
rect 7512 25563 7552 25595
rect 7584 25563 7624 25595
rect 7656 25563 7696 25595
rect 7728 25563 7768 25595
rect 7800 25563 7840 25595
rect 7872 25563 7912 25595
rect 7944 25563 7984 25595
rect 8016 25563 8056 25595
rect 8088 25563 8128 25595
rect 8160 25563 8200 25595
rect 8232 25563 8272 25595
rect 8304 25563 8344 25595
rect 8376 25563 8416 25595
rect 8448 25563 8488 25595
rect 8520 25563 8560 25595
rect 8592 25563 8632 25595
rect 8664 25563 8704 25595
rect 8736 25563 8776 25595
rect 8808 25563 8848 25595
rect 8880 25563 8920 25595
rect 8952 25563 8992 25595
rect 9024 25563 9064 25595
rect 9096 25563 9136 25595
rect 9168 25563 9208 25595
rect 9240 25563 9280 25595
rect 9312 25563 9352 25595
rect 9384 25563 9424 25595
rect 9456 25563 9496 25595
rect 9528 25563 9568 25595
rect 9600 25563 9640 25595
rect 9672 25563 9712 25595
rect 9744 25563 9784 25595
rect 9816 25563 9856 25595
rect 9888 25563 9928 25595
rect 9960 25563 10000 25595
rect 10032 25563 10072 25595
rect 10104 25563 10144 25595
rect 10176 25563 10216 25595
rect 10248 25563 10288 25595
rect 10320 25563 10360 25595
rect 10392 25563 10432 25595
rect 10464 25563 10504 25595
rect 10536 25563 10576 25595
rect 10608 25563 10648 25595
rect 10680 25563 10720 25595
rect 10752 25563 10792 25595
rect 10824 25563 10864 25595
rect 10896 25563 10936 25595
rect 10968 25563 11008 25595
rect 11040 25563 11080 25595
rect 11112 25563 11152 25595
rect 11184 25563 11224 25595
rect 11256 25563 11296 25595
rect 11328 25563 11368 25595
rect 11400 25563 11440 25595
rect 11472 25563 11512 25595
rect 11544 25563 11584 25595
rect 11616 25563 11656 25595
rect 11688 25563 11728 25595
rect 11760 25563 11800 25595
rect 11832 25563 11872 25595
rect 11904 25563 11944 25595
rect 11976 25563 12016 25595
rect 12048 25563 12088 25595
rect 12120 25563 12160 25595
rect 12192 25563 12232 25595
rect 12264 25563 12304 25595
rect 12336 25563 12376 25595
rect 12408 25563 12448 25595
rect 12480 25563 12520 25595
rect 12552 25563 12592 25595
rect 12624 25563 12664 25595
rect 12696 25563 12736 25595
rect 12768 25563 12808 25595
rect 12840 25563 12880 25595
rect 12912 25563 12952 25595
rect 12984 25563 13024 25595
rect 13056 25563 13096 25595
rect 13128 25563 13168 25595
rect 13200 25563 13240 25595
rect 13272 25563 13312 25595
rect 13344 25563 13384 25595
rect 13416 25563 13456 25595
rect 13488 25563 13528 25595
rect 13560 25563 13600 25595
rect 13632 25563 13672 25595
rect 13704 25563 13744 25595
rect 13776 25563 13816 25595
rect 13848 25563 13888 25595
rect 13920 25563 13960 25595
rect 13992 25563 14032 25595
rect 14064 25563 14104 25595
rect 14136 25563 14176 25595
rect 14208 25563 14248 25595
rect 14280 25563 14320 25595
rect 14352 25563 14392 25595
rect 14424 25563 14464 25595
rect 14496 25563 14536 25595
rect 14568 25563 14608 25595
rect 14640 25563 14680 25595
rect 14712 25563 14752 25595
rect 14784 25563 14824 25595
rect 14856 25563 14896 25595
rect 14928 25563 14968 25595
rect 15000 25563 15040 25595
rect 15072 25563 15112 25595
rect 15144 25563 15184 25595
rect 15216 25563 15256 25595
rect 15288 25563 15328 25595
rect 15360 25563 15400 25595
rect 15432 25563 15472 25595
rect 15504 25563 15544 25595
rect 15576 25563 15616 25595
rect 15648 25563 15688 25595
rect 15720 25563 15760 25595
rect 15792 25563 15832 25595
rect 15864 25563 15904 25595
rect 15936 25563 16000 25595
rect 91 25539 149 25563
rect 189 25539 247 25563
rect 287 25539 345 25563
rect 385 25539 443 25563
rect 483 25539 541 25563
rect 581 25539 639 25563
rect 679 25539 737 25563
rect 777 25539 835 25563
rect 875 25539 933 25563
rect 973 25539 1031 25563
rect 1071 25539 1129 25563
rect 1169 25539 16000 25563
rect 0 25523 16000 25539
rect 0 25491 64 25523
rect 96 25491 136 25523
rect 168 25491 208 25523
rect 240 25491 280 25523
rect 312 25491 352 25523
rect 384 25491 424 25523
rect 456 25491 496 25523
rect 528 25491 568 25523
rect 600 25491 640 25523
rect 672 25491 712 25523
rect 744 25491 784 25523
rect 816 25491 856 25523
rect 888 25491 928 25523
rect 960 25491 1000 25523
rect 1032 25491 1072 25523
rect 1104 25491 1144 25523
rect 1176 25491 1216 25523
rect 1248 25491 1288 25523
rect 1320 25491 1360 25523
rect 1392 25491 1432 25523
rect 1464 25491 1504 25523
rect 1536 25491 1576 25523
rect 1608 25491 1648 25523
rect 1680 25491 1720 25523
rect 1752 25491 1792 25523
rect 1824 25491 1864 25523
rect 1896 25491 1936 25523
rect 1968 25491 2008 25523
rect 2040 25491 2080 25523
rect 2112 25491 2152 25523
rect 2184 25491 2224 25523
rect 2256 25491 2296 25523
rect 2328 25491 2368 25523
rect 2400 25491 2440 25523
rect 2472 25491 2512 25523
rect 2544 25491 2584 25523
rect 2616 25491 2656 25523
rect 2688 25491 2728 25523
rect 2760 25491 2800 25523
rect 2832 25491 2872 25523
rect 2904 25491 2944 25523
rect 2976 25491 3016 25523
rect 3048 25491 3088 25523
rect 3120 25491 3160 25523
rect 3192 25491 3232 25523
rect 3264 25491 3304 25523
rect 3336 25491 3376 25523
rect 3408 25491 3448 25523
rect 3480 25491 3520 25523
rect 3552 25491 3592 25523
rect 3624 25491 3664 25523
rect 3696 25491 3736 25523
rect 3768 25491 3808 25523
rect 3840 25491 3880 25523
rect 3912 25491 3952 25523
rect 3984 25491 4024 25523
rect 4056 25491 4096 25523
rect 4128 25491 4168 25523
rect 4200 25491 4240 25523
rect 4272 25491 4312 25523
rect 4344 25491 4384 25523
rect 4416 25491 4456 25523
rect 4488 25491 4528 25523
rect 4560 25491 4600 25523
rect 4632 25491 4672 25523
rect 4704 25491 4744 25523
rect 4776 25491 4816 25523
rect 4848 25491 4888 25523
rect 4920 25491 4960 25523
rect 4992 25491 5032 25523
rect 5064 25491 5104 25523
rect 5136 25491 5176 25523
rect 5208 25491 5248 25523
rect 5280 25491 5320 25523
rect 5352 25491 5392 25523
rect 5424 25491 5464 25523
rect 5496 25491 5536 25523
rect 5568 25491 5608 25523
rect 5640 25491 5680 25523
rect 5712 25491 5752 25523
rect 5784 25491 5824 25523
rect 5856 25491 5896 25523
rect 5928 25491 5968 25523
rect 6000 25491 6040 25523
rect 6072 25491 6112 25523
rect 6144 25491 6184 25523
rect 6216 25491 6256 25523
rect 6288 25491 6328 25523
rect 6360 25491 6400 25523
rect 6432 25491 6472 25523
rect 6504 25491 6544 25523
rect 6576 25491 6616 25523
rect 6648 25491 6688 25523
rect 6720 25491 6760 25523
rect 6792 25491 6832 25523
rect 6864 25491 6904 25523
rect 6936 25491 6976 25523
rect 7008 25491 7048 25523
rect 7080 25491 7120 25523
rect 7152 25491 7192 25523
rect 7224 25491 7264 25523
rect 7296 25491 7336 25523
rect 7368 25491 7408 25523
rect 7440 25491 7480 25523
rect 7512 25491 7552 25523
rect 7584 25491 7624 25523
rect 7656 25491 7696 25523
rect 7728 25491 7768 25523
rect 7800 25491 7840 25523
rect 7872 25491 7912 25523
rect 7944 25491 7984 25523
rect 8016 25491 8056 25523
rect 8088 25491 8128 25523
rect 8160 25491 8200 25523
rect 8232 25491 8272 25523
rect 8304 25491 8344 25523
rect 8376 25491 8416 25523
rect 8448 25491 8488 25523
rect 8520 25491 8560 25523
rect 8592 25491 8632 25523
rect 8664 25491 8704 25523
rect 8736 25491 8776 25523
rect 8808 25491 8848 25523
rect 8880 25491 8920 25523
rect 8952 25491 8992 25523
rect 9024 25491 9064 25523
rect 9096 25491 9136 25523
rect 9168 25491 9208 25523
rect 9240 25491 9280 25523
rect 9312 25491 9352 25523
rect 9384 25491 9424 25523
rect 9456 25491 9496 25523
rect 9528 25491 9568 25523
rect 9600 25491 9640 25523
rect 9672 25491 9712 25523
rect 9744 25491 9784 25523
rect 9816 25491 9856 25523
rect 9888 25491 9928 25523
rect 9960 25491 10000 25523
rect 10032 25491 10072 25523
rect 10104 25491 10144 25523
rect 10176 25491 10216 25523
rect 10248 25491 10288 25523
rect 10320 25491 10360 25523
rect 10392 25491 10432 25523
rect 10464 25491 10504 25523
rect 10536 25491 10576 25523
rect 10608 25491 10648 25523
rect 10680 25491 10720 25523
rect 10752 25491 10792 25523
rect 10824 25491 10864 25523
rect 10896 25491 10936 25523
rect 10968 25491 11008 25523
rect 11040 25491 11080 25523
rect 11112 25491 11152 25523
rect 11184 25491 11224 25523
rect 11256 25491 11296 25523
rect 11328 25491 11368 25523
rect 11400 25491 11440 25523
rect 11472 25491 11512 25523
rect 11544 25491 11584 25523
rect 11616 25491 11656 25523
rect 11688 25491 11728 25523
rect 11760 25491 11800 25523
rect 11832 25491 11872 25523
rect 11904 25491 11944 25523
rect 11976 25491 12016 25523
rect 12048 25491 12088 25523
rect 12120 25491 12160 25523
rect 12192 25491 12232 25523
rect 12264 25491 12304 25523
rect 12336 25491 12376 25523
rect 12408 25491 12448 25523
rect 12480 25491 12520 25523
rect 12552 25491 12592 25523
rect 12624 25491 12664 25523
rect 12696 25491 12736 25523
rect 12768 25491 12808 25523
rect 12840 25491 12880 25523
rect 12912 25491 12952 25523
rect 12984 25491 13024 25523
rect 13056 25491 13096 25523
rect 13128 25491 13168 25523
rect 13200 25491 13240 25523
rect 13272 25491 13312 25523
rect 13344 25491 13384 25523
rect 13416 25491 13456 25523
rect 13488 25491 13528 25523
rect 13560 25491 13600 25523
rect 13632 25491 13672 25523
rect 13704 25491 13744 25523
rect 13776 25491 13816 25523
rect 13848 25491 13888 25523
rect 13920 25491 13960 25523
rect 13992 25491 14032 25523
rect 14064 25491 14104 25523
rect 14136 25491 14176 25523
rect 14208 25491 14248 25523
rect 14280 25491 14320 25523
rect 14352 25491 14392 25523
rect 14424 25491 14464 25523
rect 14496 25491 14536 25523
rect 14568 25491 14608 25523
rect 14640 25491 14680 25523
rect 14712 25491 14752 25523
rect 14784 25491 14824 25523
rect 14856 25491 14896 25523
rect 14928 25491 14968 25523
rect 15000 25491 15040 25523
rect 15072 25491 15112 25523
rect 15144 25491 15184 25523
rect 15216 25491 15256 25523
rect 15288 25491 15328 25523
rect 15360 25491 15400 25523
rect 15432 25491 15472 25523
rect 15504 25491 15544 25523
rect 15576 25491 15616 25523
rect 15648 25491 15688 25523
rect 15720 25491 15760 25523
rect 15792 25491 15832 25523
rect 15864 25491 15904 25523
rect 15936 25491 16000 25523
rect 0 25481 16000 25491
rect 0 25441 51 25481
rect 91 25451 149 25481
rect 189 25451 247 25481
rect 287 25451 345 25481
rect 385 25451 443 25481
rect 483 25451 541 25481
rect 581 25451 639 25481
rect 679 25451 737 25481
rect 777 25451 835 25481
rect 875 25451 933 25481
rect 973 25451 1031 25481
rect 1071 25451 1129 25481
rect 1169 25451 16000 25481
rect 0 25419 64 25441
rect 96 25419 136 25451
rect 189 25441 208 25451
rect 168 25419 208 25441
rect 240 25441 247 25451
rect 312 25441 345 25451
rect 385 25441 424 25451
rect 483 25441 496 25451
rect 240 25419 280 25441
rect 312 25419 352 25441
rect 384 25419 424 25441
rect 456 25419 496 25441
rect 528 25441 541 25451
rect 600 25441 639 25451
rect 679 25441 712 25451
rect 777 25441 784 25451
rect 528 25419 568 25441
rect 600 25419 640 25441
rect 672 25419 712 25441
rect 744 25419 784 25441
rect 816 25441 835 25451
rect 816 25419 856 25441
rect 888 25419 928 25451
rect 973 25441 1000 25451
rect 1071 25441 1072 25451
rect 960 25419 1000 25441
rect 1032 25419 1072 25441
rect 1104 25441 1129 25451
rect 1104 25419 1144 25441
rect 1176 25419 1216 25451
rect 1248 25419 1288 25451
rect 1320 25419 1360 25451
rect 1392 25419 1432 25451
rect 1464 25419 1504 25451
rect 1536 25419 1576 25451
rect 1608 25419 1648 25451
rect 1680 25419 1720 25451
rect 1752 25419 1792 25451
rect 1824 25419 1864 25451
rect 1896 25419 1936 25451
rect 1968 25419 2008 25451
rect 2040 25419 2080 25451
rect 2112 25419 2152 25451
rect 2184 25419 2224 25451
rect 2256 25419 2296 25451
rect 2328 25419 2368 25451
rect 2400 25419 2440 25451
rect 2472 25419 2512 25451
rect 2544 25419 2584 25451
rect 2616 25419 2656 25451
rect 2688 25419 2728 25451
rect 2760 25419 2800 25451
rect 2832 25419 2872 25451
rect 2904 25419 2944 25451
rect 2976 25419 3016 25451
rect 3048 25419 3088 25451
rect 3120 25419 3160 25451
rect 3192 25419 3232 25451
rect 3264 25419 3304 25451
rect 3336 25419 3376 25451
rect 3408 25419 3448 25451
rect 3480 25419 3520 25451
rect 3552 25419 3592 25451
rect 3624 25419 3664 25451
rect 3696 25419 3736 25451
rect 3768 25419 3808 25451
rect 3840 25419 3880 25451
rect 3912 25419 3952 25451
rect 3984 25419 4024 25451
rect 4056 25419 4096 25451
rect 4128 25419 4168 25451
rect 4200 25419 4240 25451
rect 4272 25419 4312 25451
rect 4344 25419 4384 25451
rect 4416 25419 4456 25451
rect 4488 25419 4528 25451
rect 4560 25419 4600 25451
rect 4632 25419 4672 25451
rect 4704 25419 4744 25451
rect 4776 25419 4816 25451
rect 4848 25419 4888 25451
rect 4920 25419 4960 25451
rect 4992 25419 5032 25451
rect 5064 25419 5104 25451
rect 5136 25419 5176 25451
rect 5208 25419 5248 25451
rect 5280 25419 5320 25451
rect 5352 25419 5392 25451
rect 5424 25419 5464 25451
rect 5496 25419 5536 25451
rect 5568 25419 5608 25451
rect 5640 25419 5680 25451
rect 5712 25419 5752 25451
rect 5784 25419 5824 25451
rect 5856 25419 5896 25451
rect 5928 25419 5968 25451
rect 6000 25419 6040 25451
rect 6072 25419 6112 25451
rect 6144 25419 6184 25451
rect 6216 25419 6256 25451
rect 6288 25419 6328 25451
rect 6360 25419 6400 25451
rect 6432 25419 6472 25451
rect 6504 25419 6544 25451
rect 6576 25419 6616 25451
rect 6648 25419 6688 25451
rect 6720 25419 6760 25451
rect 6792 25419 6832 25451
rect 6864 25419 6904 25451
rect 6936 25419 6976 25451
rect 7008 25419 7048 25451
rect 7080 25419 7120 25451
rect 7152 25419 7192 25451
rect 7224 25419 7264 25451
rect 7296 25419 7336 25451
rect 7368 25419 7408 25451
rect 7440 25419 7480 25451
rect 7512 25419 7552 25451
rect 7584 25419 7624 25451
rect 7656 25419 7696 25451
rect 7728 25419 7768 25451
rect 7800 25419 7840 25451
rect 7872 25419 7912 25451
rect 7944 25419 7984 25451
rect 8016 25419 8056 25451
rect 8088 25419 8128 25451
rect 8160 25419 8200 25451
rect 8232 25419 8272 25451
rect 8304 25419 8344 25451
rect 8376 25419 8416 25451
rect 8448 25419 8488 25451
rect 8520 25419 8560 25451
rect 8592 25419 8632 25451
rect 8664 25419 8704 25451
rect 8736 25419 8776 25451
rect 8808 25419 8848 25451
rect 8880 25419 8920 25451
rect 8952 25419 8992 25451
rect 9024 25419 9064 25451
rect 9096 25419 9136 25451
rect 9168 25419 9208 25451
rect 9240 25419 9280 25451
rect 9312 25419 9352 25451
rect 9384 25419 9424 25451
rect 9456 25419 9496 25451
rect 9528 25419 9568 25451
rect 9600 25419 9640 25451
rect 9672 25419 9712 25451
rect 9744 25419 9784 25451
rect 9816 25419 9856 25451
rect 9888 25419 9928 25451
rect 9960 25419 10000 25451
rect 10032 25419 10072 25451
rect 10104 25419 10144 25451
rect 10176 25419 10216 25451
rect 10248 25419 10288 25451
rect 10320 25419 10360 25451
rect 10392 25419 10432 25451
rect 10464 25419 10504 25451
rect 10536 25419 10576 25451
rect 10608 25419 10648 25451
rect 10680 25419 10720 25451
rect 10752 25419 10792 25451
rect 10824 25419 10864 25451
rect 10896 25419 10936 25451
rect 10968 25419 11008 25451
rect 11040 25419 11080 25451
rect 11112 25419 11152 25451
rect 11184 25419 11224 25451
rect 11256 25419 11296 25451
rect 11328 25419 11368 25451
rect 11400 25419 11440 25451
rect 11472 25419 11512 25451
rect 11544 25419 11584 25451
rect 11616 25419 11656 25451
rect 11688 25419 11728 25451
rect 11760 25419 11800 25451
rect 11832 25419 11872 25451
rect 11904 25419 11944 25451
rect 11976 25419 12016 25451
rect 12048 25419 12088 25451
rect 12120 25419 12160 25451
rect 12192 25419 12232 25451
rect 12264 25419 12304 25451
rect 12336 25419 12376 25451
rect 12408 25419 12448 25451
rect 12480 25419 12520 25451
rect 12552 25419 12592 25451
rect 12624 25419 12664 25451
rect 12696 25419 12736 25451
rect 12768 25419 12808 25451
rect 12840 25419 12880 25451
rect 12912 25419 12952 25451
rect 12984 25419 13024 25451
rect 13056 25419 13096 25451
rect 13128 25419 13168 25451
rect 13200 25419 13240 25451
rect 13272 25419 13312 25451
rect 13344 25419 13384 25451
rect 13416 25419 13456 25451
rect 13488 25419 13528 25451
rect 13560 25419 13600 25451
rect 13632 25419 13672 25451
rect 13704 25419 13744 25451
rect 13776 25419 13816 25451
rect 13848 25419 13888 25451
rect 13920 25419 13960 25451
rect 13992 25419 14032 25451
rect 14064 25419 14104 25451
rect 14136 25419 14176 25451
rect 14208 25419 14248 25451
rect 14280 25419 14320 25451
rect 14352 25419 14392 25451
rect 14424 25419 14464 25451
rect 14496 25419 14536 25451
rect 14568 25419 14608 25451
rect 14640 25419 14680 25451
rect 14712 25419 14752 25451
rect 14784 25419 14824 25451
rect 14856 25419 14896 25451
rect 14928 25419 14968 25451
rect 15000 25419 15040 25451
rect 15072 25419 15112 25451
rect 15144 25419 15184 25451
rect 15216 25419 15256 25451
rect 15288 25419 15328 25451
rect 15360 25419 15400 25451
rect 15432 25419 15472 25451
rect 15504 25419 15544 25451
rect 15576 25419 15616 25451
rect 15648 25419 15688 25451
rect 15720 25419 15760 25451
rect 15792 25419 15832 25451
rect 15864 25419 15904 25451
rect 15936 25419 16000 25451
rect 0 25383 16000 25419
rect 0 25343 51 25383
rect 91 25379 149 25383
rect 189 25379 247 25383
rect 287 25379 345 25383
rect 385 25379 443 25383
rect 483 25379 541 25383
rect 581 25379 639 25383
rect 679 25379 737 25383
rect 777 25379 835 25383
rect 875 25379 933 25383
rect 973 25379 1031 25383
rect 1071 25379 1129 25383
rect 1169 25379 16000 25383
rect 96 25347 136 25379
rect 189 25347 208 25379
rect 240 25347 247 25379
rect 312 25347 345 25379
rect 385 25347 424 25379
rect 483 25347 496 25379
rect 528 25347 541 25379
rect 600 25347 639 25379
rect 679 25347 712 25379
rect 777 25347 784 25379
rect 816 25347 835 25379
rect 888 25347 928 25379
rect 973 25347 1000 25379
rect 1071 25347 1072 25379
rect 1104 25347 1129 25379
rect 1176 25347 1216 25379
rect 1248 25347 1288 25379
rect 1320 25347 1360 25379
rect 1392 25347 1432 25379
rect 1464 25347 1504 25379
rect 1536 25347 1576 25379
rect 1608 25347 1648 25379
rect 1680 25347 1720 25379
rect 1752 25347 1792 25379
rect 1824 25347 1864 25379
rect 1896 25347 1936 25379
rect 1968 25347 2008 25379
rect 2040 25347 2080 25379
rect 2112 25347 2152 25379
rect 2184 25347 2224 25379
rect 2256 25347 2296 25379
rect 2328 25347 2368 25379
rect 2400 25347 2440 25379
rect 2472 25347 2512 25379
rect 2544 25347 2584 25379
rect 2616 25347 2656 25379
rect 2688 25347 2728 25379
rect 2760 25347 2800 25379
rect 2832 25347 2872 25379
rect 2904 25347 2944 25379
rect 2976 25347 3016 25379
rect 3048 25347 3088 25379
rect 3120 25347 3160 25379
rect 3192 25347 3232 25379
rect 3264 25347 3304 25379
rect 3336 25347 3376 25379
rect 3408 25347 3448 25379
rect 3480 25347 3520 25379
rect 3552 25347 3592 25379
rect 3624 25347 3664 25379
rect 3696 25347 3736 25379
rect 3768 25347 3808 25379
rect 3840 25347 3880 25379
rect 3912 25347 3952 25379
rect 3984 25347 4024 25379
rect 4056 25347 4096 25379
rect 4128 25347 4168 25379
rect 4200 25347 4240 25379
rect 4272 25347 4312 25379
rect 4344 25347 4384 25379
rect 4416 25347 4456 25379
rect 4488 25347 4528 25379
rect 4560 25347 4600 25379
rect 4632 25347 4672 25379
rect 4704 25347 4744 25379
rect 4776 25347 4816 25379
rect 4848 25347 4888 25379
rect 4920 25347 4960 25379
rect 4992 25347 5032 25379
rect 5064 25347 5104 25379
rect 5136 25347 5176 25379
rect 5208 25347 5248 25379
rect 5280 25347 5320 25379
rect 5352 25347 5392 25379
rect 5424 25347 5464 25379
rect 5496 25347 5536 25379
rect 5568 25347 5608 25379
rect 5640 25347 5680 25379
rect 5712 25347 5752 25379
rect 5784 25347 5824 25379
rect 5856 25347 5896 25379
rect 5928 25347 5968 25379
rect 6000 25347 6040 25379
rect 6072 25347 6112 25379
rect 6144 25347 6184 25379
rect 6216 25347 6256 25379
rect 6288 25347 6328 25379
rect 6360 25347 6400 25379
rect 6432 25347 6472 25379
rect 6504 25347 6544 25379
rect 6576 25347 6616 25379
rect 6648 25347 6688 25379
rect 6720 25347 6760 25379
rect 6792 25347 6832 25379
rect 6864 25347 6904 25379
rect 6936 25347 6976 25379
rect 7008 25347 7048 25379
rect 7080 25347 7120 25379
rect 7152 25347 7192 25379
rect 7224 25347 7264 25379
rect 7296 25347 7336 25379
rect 7368 25347 7408 25379
rect 7440 25347 7480 25379
rect 7512 25347 7552 25379
rect 7584 25347 7624 25379
rect 7656 25347 7696 25379
rect 7728 25347 7768 25379
rect 7800 25347 7840 25379
rect 7872 25347 7912 25379
rect 7944 25347 7984 25379
rect 8016 25347 8056 25379
rect 8088 25347 8128 25379
rect 8160 25347 8200 25379
rect 8232 25347 8272 25379
rect 8304 25347 8344 25379
rect 8376 25347 8416 25379
rect 8448 25347 8488 25379
rect 8520 25347 8560 25379
rect 8592 25347 8632 25379
rect 8664 25347 8704 25379
rect 8736 25347 8776 25379
rect 8808 25347 8848 25379
rect 8880 25347 8920 25379
rect 8952 25347 8992 25379
rect 9024 25347 9064 25379
rect 9096 25347 9136 25379
rect 9168 25347 9208 25379
rect 9240 25347 9280 25379
rect 9312 25347 9352 25379
rect 9384 25347 9424 25379
rect 9456 25347 9496 25379
rect 9528 25347 9568 25379
rect 9600 25347 9640 25379
rect 9672 25347 9712 25379
rect 9744 25347 9784 25379
rect 9816 25347 9856 25379
rect 9888 25347 9928 25379
rect 9960 25347 10000 25379
rect 10032 25347 10072 25379
rect 10104 25347 10144 25379
rect 10176 25347 10216 25379
rect 10248 25347 10288 25379
rect 10320 25347 10360 25379
rect 10392 25347 10432 25379
rect 10464 25347 10504 25379
rect 10536 25347 10576 25379
rect 10608 25347 10648 25379
rect 10680 25347 10720 25379
rect 10752 25347 10792 25379
rect 10824 25347 10864 25379
rect 10896 25347 10936 25379
rect 10968 25347 11008 25379
rect 11040 25347 11080 25379
rect 11112 25347 11152 25379
rect 11184 25347 11224 25379
rect 11256 25347 11296 25379
rect 11328 25347 11368 25379
rect 11400 25347 11440 25379
rect 11472 25347 11512 25379
rect 11544 25347 11584 25379
rect 11616 25347 11656 25379
rect 11688 25347 11728 25379
rect 11760 25347 11800 25379
rect 11832 25347 11872 25379
rect 11904 25347 11944 25379
rect 11976 25347 12016 25379
rect 12048 25347 12088 25379
rect 12120 25347 12160 25379
rect 12192 25347 12232 25379
rect 12264 25347 12304 25379
rect 12336 25347 12376 25379
rect 12408 25347 12448 25379
rect 12480 25347 12520 25379
rect 12552 25347 12592 25379
rect 12624 25347 12664 25379
rect 12696 25347 12736 25379
rect 12768 25347 12808 25379
rect 12840 25347 12880 25379
rect 12912 25347 12952 25379
rect 12984 25347 13024 25379
rect 13056 25347 13096 25379
rect 13128 25347 13168 25379
rect 13200 25347 13240 25379
rect 13272 25347 13312 25379
rect 13344 25347 13384 25379
rect 13416 25347 13456 25379
rect 13488 25347 13528 25379
rect 13560 25347 13600 25379
rect 13632 25347 13672 25379
rect 13704 25347 13744 25379
rect 13776 25347 13816 25379
rect 13848 25347 13888 25379
rect 13920 25347 13960 25379
rect 13992 25347 14032 25379
rect 14064 25347 14104 25379
rect 14136 25347 14176 25379
rect 14208 25347 14248 25379
rect 14280 25347 14320 25379
rect 14352 25347 14392 25379
rect 14424 25347 14464 25379
rect 14496 25347 14536 25379
rect 14568 25347 14608 25379
rect 14640 25347 14680 25379
rect 14712 25347 14752 25379
rect 14784 25347 14824 25379
rect 14856 25347 14896 25379
rect 14928 25347 14968 25379
rect 15000 25347 15040 25379
rect 15072 25347 15112 25379
rect 15144 25347 15184 25379
rect 15216 25347 15256 25379
rect 15288 25347 15328 25379
rect 15360 25347 15400 25379
rect 15432 25347 15472 25379
rect 15504 25347 15544 25379
rect 15576 25347 15616 25379
rect 15648 25347 15688 25379
rect 15720 25347 15760 25379
rect 15792 25347 15832 25379
rect 15864 25347 15904 25379
rect 15936 25347 16000 25379
rect 91 25343 149 25347
rect 189 25343 247 25347
rect 287 25343 345 25347
rect 385 25343 443 25347
rect 483 25343 541 25347
rect 581 25343 639 25347
rect 679 25343 737 25347
rect 777 25343 835 25347
rect 875 25343 933 25347
rect 973 25343 1031 25347
rect 1071 25343 1129 25347
rect 1169 25343 16000 25347
rect 0 25307 16000 25343
rect 0 25285 64 25307
rect 0 25245 51 25285
rect 96 25275 136 25307
rect 168 25285 208 25307
rect 189 25275 208 25285
rect 240 25285 280 25307
rect 312 25285 352 25307
rect 384 25285 424 25307
rect 456 25285 496 25307
rect 240 25275 247 25285
rect 312 25275 345 25285
rect 385 25275 424 25285
rect 483 25275 496 25285
rect 528 25285 568 25307
rect 600 25285 640 25307
rect 672 25285 712 25307
rect 744 25285 784 25307
rect 528 25275 541 25285
rect 600 25275 639 25285
rect 679 25275 712 25285
rect 777 25275 784 25285
rect 816 25285 856 25307
rect 816 25275 835 25285
rect 888 25275 928 25307
rect 960 25285 1000 25307
rect 1032 25285 1072 25307
rect 973 25275 1000 25285
rect 1071 25275 1072 25285
rect 1104 25285 1144 25307
rect 1104 25275 1129 25285
rect 1176 25275 1216 25307
rect 1248 25275 1288 25307
rect 1320 25275 1360 25307
rect 1392 25275 1432 25307
rect 1464 25275 1504 25307
rect 1536 25275 1576 25307
rect 1608 25275 1648 25307
rect 1680 25275 1720 25307
rect 1752 25275 1792 25307
rect 1824 25275 1864 25307
rect 1896 25275 1936 25307
rect 1968 25275 2008 25307
rect 2040 25275 2080 25307
rect 2112 25275 2152 25307
rect 2184 25275 2224 25307
rect 2256 25275 2296 25307
rect 2328 25275 2368 25307
rect 2400 25275 2440 25307
rect 2472 25275 2512 25307
rect 2544 25275 2584 25307
rect 2616 25275 2656 25307
rect 2688 25275 2728 25307
rect 2760 25275 2800 25307
rect 2832 25275 2872 25307
rect 2904 25275 2944 25307
rect 2976 25275 3016 25307
rect 3048 25275 3088 25307
rect 3120 25275 3160 25307
rect 3192 25275 3232 25307
rect 3264 25275 3304 25307
rect 3336 25275 3376 25307
rect 3408 25275 3448 25307
rect 3480 25275 3520 25307
rect 3552 25275 3592 25307
rect 3624 25275 3664 25307
rect 3696 25275 3736 25307
rect 3768 25275 3808 25307
rect 3840 25275 3880 25307
rect 3912 25275 3952 25307
rect 3984 25275 4024 25307
rect 4056 25275 4096 25307
rect 4128 25275 4168 25307
rect 4200 25275 4240 25307
rect 4272 25275 4312 25307
rect 4344 25275 4384 25307
rect 4416 25275 4456 25307
rect 4488 25275 4528 25307
rect 4560 25275 4600 25307
rect 4632 25275 4672 25307
rect 4704 25275 4744 25307
rect 4776 25275 4816 25307
rect 4848 25275 4888 25307
rect 4920 25275 4960 25307
rect 4992 25275 5032 25307
rect 5064 25275 5104 25307
rect 5136 25275 5176 25307
rect 5208 25275 5248 25307
rect 5280 25275 5320 25307
rect 5352 25275 5392 25307
rect 5424 25275 5464 25307
rect 5496 25275 5536 25307
rect 5568 25275 5608 25307
rect 5640 25275 5680 25307
rect 5712 25275 5752 25307
rect 5784 25275 5824 25307
rect 5856 25275 5896 25307
rect 5928 25275 5968 25307
rect 6000 25275 6040 25307
rect 6072 25275 6112 25307
rect 6144 25275 6184 25307
rect 6216 25275 6256 25307
rect 6288 25275 6328 25307
rect 6360 25275 6400 25307
rect 6432 25275 6472 25307
rect 6504 25275 6544 25307
rect 6576 25275 6616 25307
rect 6648 25275 6688 25307
rect 6720 25275 6760 25307
rect 6792 25275 6832 25307
rect 6864 25275 6904 25307
rect 6936 25275 6976 25307
rect 7008 25275 7048 25307
rect 7080 25275 7120 25307
rect 7152 25275 7192 25307
rect 7224 25275 7264 25307
rect 7296 25275 7336 25307
rect 7368 25275 7408 25307
rect 7440 25275 7480 25307
rect 7512 25275 7552 25307
rect 7584 25275 7624 25307
rect 7656 25275 7696 25307
rect 7728 25275 7768 25307
rect 7800 25275 7840 25307
rect 7872 25275 7912 25307
rect 7944 25275 7984 25307
rect 8016 25275 8056 25307
rect 8088 25275 8128 25307
rect 8160 25275 8200 25307
rect 8232 25275 8272 25307
rect 8304 25275 8344 25307
rect 8376 25275 8416 25307
rect 8448 25275 8488 25307
rect 8520 25275 8560 25307
rect 8592 25275 8632 25307
rect 8664 25275 8704 25307
rect 8736 25275 8776 25307
rect 8808 25275 8848 25307
rect 8880 25275 8920 25307
rect 8952 25275 8992 25307
rect 9024 25275 9064 25307
rect 9096 25275 9136 25307
rect 9168 25275 9208 25307
rect 9240 25275 9280 25307
rect 9312 25275 9352 25307
rect 9384 25275 9424 25307
rect 9456 25275 9496 25307
rect 9528 25275 9568 25307
rect 9600 25275 9640 25307
rect 9672 25275 9712 25307
rect 9744 25275 9784 25307
rect 9816 25275 9856 25307
rect 9888 25275 9928 25307
rect 9960 25275 10000 25307
rect 10032 25275 10072 25307
rect 10104 25275 10144 25307
rect 10176 25275 10216 25307
rect 10248 25275 10288 25307
rect 10320 25275 10360 25307
rect 10392 25275 10432 25307
rect 10464 25275 10504 25307
rect 10536 25275 10576 25307
rect 10608 25275 10648 25307
rect 10680 25275 10720 25307
rect 10752 25275 10792 25307
rect 10824 25275 10864 25307
rect 10896 25275 10936 25307
rect 10968 25275 11008 25307
rect 11040 25275 11080 25307
rect 11112 25275 11152 25307
rect 11184 25275 11224 25307
rect 11256 25275 11296 25307
rect 11328 25275 11368 25307
rect 11400 25275 11440 25307
rect 11472 25275 11512 25307
rect 11544 25275 11584 25307
rect 11616 25275 11656 25307
rect 11688 25275 11728 25307
rect 11760 25275 11800 25307
rect 11832 25275 11872 25307
rect 11904 25275 11944 25307
rect 11976 25275 12016 25307
rect 12048 25275 12088 25307
rect 12120 25275 12160 25307
rect 12192 25275 12232 25307
rect 12264 25275 12304 25307
rect 12336 25275 12376 25307
rect 12408 25275 12448 25307
rect 12480 25275 12520 25307
rect 12552 25275 12592 25307
rect 12624 25275 12664 25307
rect 12696 25275 12736 25307
rect 12768 25275 12808 25307
rect 12840 25275 12880 25307
rect 12912 25275 12952 25307
rect 12984 25275 13024 25307
rect 13056 25275 13096 25307
rect 13128 25275 13168 25307
rect 13200 25275 13240 25307
rect 13272 25275 13312 25307
rect 13344 25275 13384 25307
rect 13416 25275 13456 25307
rect 13488 25275 13528 25307
rect 13560 25275 13600 25307
rect 13632 25275 13672 25307
rect 13704 25275 13744 25307
rect 13776 25275 13816 25307
rect 13848 25275 13888 25307
rect 13920 25275 13960 25307
rect 13992 25275 14032 25307
rect 14064 25275 14104 25307
rect 14136 25275 14176 25307
rect 14208 25275 14248 25307
rect 14280 25275 14320 25307
rect 14352 25275 14392 25307
rect 14424 25275 14464 25307
rect 14496 25275 14536 25307
rect 14568 25275 14608 25307
rect 14640 25275 14680 25307
rect 14712 25275 14752 25307
rect 14784 25275 14824 25307
rect 14856 25275 14896 25307
rect 14928 25275 14968 25307
rect 15000 25275 15040 25307
rect 15072 25275 15112 25307
rect 15144 25275 15184 25307
rect 15216 25275 15256 25307
rect 15288 25275 15328 25307
rect 15360 25275 15400 25307
rect 15432 25275 15472 25307
rect 15504 25275 15544 25307
rect 15576 25275 15616 25307
rect 15648 25275 15688 25307
rect 15720 25275 15760 25307
rect 15792 25275 15832 25307
rect 15864 25275 15904 25307
rect 15936 25275 16000 25307
rect 91 25245 149 25275
rect 189 25245 247 25275
rect 287 25245 345 25275
rect 385 25245 443 25275
rect 483 25245 541 25275
rect 581 25245 639 25275
rect 679 25245 737 25275
rect 777 25245 835 25275
rect 875 25245 933 25275
rect 973 25245 1031 25275
rect 1071 25245 1129 25275
rect 1169 25245 16000 25275
rect 0 25235 16000 25245
rect 0 25203 64 25235
rect 96 25203 136 25235
rect 168 25203 208 25235
rect 240 25203 280 25235
rect 312 25203 352 25235
rect 384 25203 424 25235
rect 456 25203 496 25235
rect 528 25203 568 25235
rect 600 25203 640 25235
rect 672 25203 712 25235
rect 744 25203 784 25235
rect 816 25203 856 25235
rect 888 25203 928 25235
rect 960 25203 1000 25235
rect 1032 25203 1072 25235
rect 1104 25203 1144 25235
rect 1176 25203 1216 25235
rect 1248 25203 1288 25235
rect 1320 25203 1360 25235
rect 1392 25203 1432 25235
rect 1464 25203 1504 25235
rect 1536 25203 1576 25235
rect 1608 25203 1648 25235
rect 1680 25203 1720 25235
rect 1752 25203 1792 25235
rect 1824 25203 1864 25235
rect 1896 25203 1936 25235
rect 1968 25203 2008 25235
rect 2040 25203 2080 25235
rect 2112 25203 2152 25235
rect 2184 25203 2224 25235
rect 2256 25203 2296 25235
rect 2328 25203 2368 25235
rect 2400 25203 2440 25235
rect 2472 25203 2512 25235
rect 2544 25203 2584 25235
rect 2616 25203 2656 25235
rect 2688 25203 2728 25235
rect 2760 25203 2800 25235
rect 2832 25203 2872 25235
rect 2904 25203 2944 25235
rect 2976 25203 3016 25235
rect 3048 25203 3088 25235
rect 3120 25203 3160 25235
rect 3192 25203 3232 25235
rect 3264 25203 3304 25235
rect 3336 25203 3376 25235
rect 3408 25203 3448 25235
rect 3480 25203 3520 25235
rect 3552 25203 3592 25235
rect 3624 25203 3664 25235
rect 3696 25203 3736 25235
rect 3768 25203 3808 25235
rect 3840 25203 3880 25235
rect 3912 25203 3952 25235
rect 3984 25203 4024 25235
rect 4056 25203 4096 25235
rect 4128 25203 4168 25235
rect 4200 25203 4240 25235
rect 4272 25203 4312 25235
rect 4344 25203 4384 25235
rect 4416 25203 4456 25235
rect 4488 25203 4528 25235
rect 4560 25203 4600 25235
rect 4632 25203 4672 25235
rect 4704 25203 4744 25235
rect 4776 25203 4816 25235
rect 4848 25203 4888 25235
rect 4920 25203 4960 25235
rect 4992 25203 5032 25235
rect 5064 25203 5104 25235
rect 5136 25203 5176 25235
rect 5208 25203 5248 25235
rect 5280 25203 5320 25235
rect 5352 25203 5392 25235
rect 5424 25203 5464 25235
rect 5496 25203 5536 25235
rect 5568 25203 5608 25235
rect 5640 25203 5680 25235
rect 5712 25203 5752 25235
rect 5784 25203 5824 25235
rect 5856 25203 5896 25235
rect 5928 25203 5968 25235
rect 6000 25203 6040 25235
rect 6072 25203 6112 25235
rect 6144 25203 6184 25235
rect 6216 25203 6256 25235
rect 6288 25203 6328 25235
rect 6360 25203 6400 25235
rect 6432 25203 6472 25235
rect 6504 25203 6544 25235
rect 6576 25203 6616 25235
rect 6648 25203 6688 25235
rect 6720 25203 6760 25235
rect 6792 25203 6832 25235
rect 6864 25203 6904 25235
rect 6936 25203 6976 25235
rect 7008 25203 7048 25235
rect 7080 25203 7120 25235
rect 7152 25203 7192 25235
rect 7224 25203 7264 25235
rect 7296 25203 7336 25235
rect 7368 25203 7408 25235
rect 7440 25203 7480 25235
rect 7512 25203 7552 25235
rect 7584 25203 7624 25235
rect 7656 25203 7696 25235
rect 7728 25203 7768 25235
rect 7800 25203 7840 25235
rect 7872 25203 7912 25235
rect 7944 25203 7984 25235
rect 8016 25203 8056 25235
rect 8088 25203 8128 25235
rect 8160 25203 8200 25235
rect 8232 25203 8272 25235
rect 8304 25203 8344 25235
rect 8376 25203 8416 25235
rect 8448 25203 8488 25235
rect 8520 25203 8560 25235
rect 8592 25203 8632 25235
rect 8664 25203 8704 25235
rect 8736 25203 8776 25235
rect 8808 25203 8848 25235
rect 8880 25203 8920 25235
rect 8952 25203 8992 25235
rect 9024 25203 9064 25235
rect 9096 25203 9136 25235
rect 9168 25203 9208 25235
rect 9240 25203 9280 25235
rect 9312 25203 9352 25235
rect 9384 25203 9424 25235
rect 9456 25203 9496 25235
rect 9528 25203 9568 25235
rect 9600 25203 9640 25235
rect 9672 25203 9712 25235
rect 9744 25203 9784 25235
rect 9816 25203 9856 25235
rect 9888 25203 9928 25235
rect 9960 25203 10000 25235
rect 10032 25203 10072 25235
rect 10104 25203 10144 25235
rect 10176 25203 10216 25235
rect 10248 25203 10288 25235
rect 10320 25203 10360 25235
rect 10392 25203 10432 25235
rect 10464 25203 10504 25235
rect 10536 25203 10576 25235
rect 10608 25203 10648 25235
rect 10680 25203 10720 25235
rect 10752 25203 10792 25235
rect 10824 25203 10864 25235
rect 10896 25203 10936 25235
rect 10968 25203 11008 25235
rect 11040 25203 11080 25235
rect 11112 25203 11152 25235
rect 11184 25203 11224 25235
rect 11256 25203 11296 25235
rect 11328 25203 11368 25235
rect 11400 25203 11440 25235
rect 11472 25203 11512 25235
rect 11544 25203 11584 25235
rect 11616 25203 11656 25235
rect 11688 25203 11728 25235
rect 11760 25203 11800 25235
rect 11832 25203 11872 25235
rect 11904 25203 11944 25235
rect 11976 25203 12016 25235
rect 12048 25203 12088 25235
rect 12120 25203 12160 25235
rect 12192 25203 12232 25235
rect 12264 25203 12304 25235
rect 12336 25203 12376 25235
rect 12408 25203 12448 25235
rect 12480 25203 12520 25235
rect 12552 25203 12592 25235
rect 12624 25203 12664 25235
rect 12696 25203 12736 25235
rect 12768 25203 12808 25235
rect 12840 25203 12880 25235
rect 12912 25203 12952 25235
rect 12984 25203 13024 25235
rect 13056 25203 13096 25235
rect 13128 25203 13168 25235
rect 13200 25203 13240 25235
rect 13272 25203 13312 25235
rect 13344 25203 13384 25235
rect 13416 25203 13456 25235
rect 13488 25203 13528 25235
rect 13560 25203 13600 25235
rect 13632 25203 13672 25235
rect 13704 25203 13744 25235
rect 13776 25203 13816 25235
rect 13848 25203 13888 25235
rect 13920 25203 13960 25235
rect 13992 25203 14032 25235
rect 14064 25203 14104 25235
rect 14136 25203 14176 25235
rect 14208 25203 14248 25235
rect 14280 25203 14320 25235
rect 14352 25203 14392 25235
rect 14424 25203 14464 25235
rect 14496 25203 14536 25235
rect 14568 25203 14608 25235
rect 14640 25203 14680 25235
rect 14712 25203 14752 25235
rect 14784 25203 14824 25235
rect 14856 25203 14896 25235
rect 14928 25203 14968 25235
rect 15000 25203 15040 25235
rect 15072 25203 15112 25235
rect 15144 25203 15184 25235
rect 15216 25203 15256 25235
rect 15288 25203 15328 25235
rect 15360 25203 15400 25235
rect 15432 25203 15472 25235
rect 15504 25203 15544 25235
rect 15576 25203 15616 25235
rect 15648 25203 15688 25235
rect 15720 25203 15760 25235
rect 15792 25203 15832 25235
rect 15864 25203 15904 25235
rect 15936 25203 16000 25235
rect 0 25163 16000 25203
rect 0 25131 64 25163
rect 96 25131 136 25163
rect 168 25131 208 25163
rect 240 25131 280 25163
rect 312 25131 352 25163
rect 384 25131 424 25163
rect 456 25131 496 25163
rect 528 25131 568 25163
rect 600 25131 640 25163
rect 672 25131 712 25163
rect 744 25131 784 25163
rect 816 25131 856 25163
rect 888 25131 928 25163
rect 960 25131 1000 25163
rect 1032 25131 1072 25163
rect 1104 25131 1144 25163
rect 1176 25131 1216 25163
rect 1248 25131 1288 25163
rect 1320 25131 1360 25163
rect 1392 25131 1432 25163
rect 1464 25131 1504 25163
rect 1536 25131 1576 25163
rect 1608 25131 1648 25163
rect 1680 25131 1720 25163
rect 1752 25131 1792 25163
rect 1824 25131 1864 25163
rect 1896 25131 1936 25163
rect 1968 25131 2008 25163
rect 2040 25131 2080 25163
rect 2112 25131 2152 25163
rect 2184 25131 2224 25163
rect 2256 25131 2296 25163
rect 2328 25131 2368 25163
rect 2400 25131 2440 25163
rect 2472 25131 2512 25163
rect 2544 25131 2584 25163
rect 2616 25131 2656 25163
rect 2688 25131 2728 25163
rect 2760 25131 2800 25163
rect 2832 25131 2872 25163
rect 2904 25131 2944 25163
rect 2976 25131 3016 25163
rect 3048 25131 3088 25163
rect 3120 25131 3160 25163
rect 3192 25131 3232 25163
rect 3264 25131 3304 25163
rect 3336 25131 3376 25163
rect 3408 25131 3448 25163
rect 3480 25131 3520 25163
rect 3552 25131 3592 25163
rect 3624 25131 3664 25163
rect 3696 25131 3736 25163
rect 3768 25131 3808 25163
rect 3840 25131 3880 25163
rect 3912 25131 3952 25163
rect 3984 25131 4024 25163
rect 4056 25131 4096 25163
rect 4128 25131 4168 25163
rect 4200 25131 4240 25163
rect 4272 25131 4312 25163
rect 4344 25131 4384 25163
rect 4416 25131 4456 25163
rect 4488 25131 4528 25163
rect 4560 25131 4600 25163
rect 4632 25131 4672 25163
rect 4704 25131 4744 25163
rect 4776 25131 4816 25163
rect 4848 25131 4888 25163
rect 4920 25131 4960 25163
rect 4992 25131 5032 25163
rect 5064 25131 5104 25163
rect 5136 25131 5176 25163
rect 5208 25131 5248 25163
rect 5280 25131 5320 25163
rect 5352 25131 5392 25163
rect 5424 25131 5464 25163
rect 5496 25131 5536 25163
rect 5568 25131 5608 25163
rect 5640 25131 5680 25163
rect 5712 25131 5752 25163
rect 5784 25131 5824 25163
rect 5856 25131 5896 25163
rect 5928 25131 5968 25163
rect 6000 25131 6040 25163
rect 6072 25131 6112 25163
rect 6144 25131 6184 25163
rect 6216 25131 6256 25163
rect 6288 25131 6328 25163
rect 6360 25131 6400 25163
rect 6432 25131 6472 25163
rect 6504 25131 6544 25163
rect 6576 25131 6616 25163
rect 6648 25131 6688 25163
rect 6720 25131 6760 25163
rect 6792 25131 6832 25163
rect 6864 25131 6904 25163
rect 6936 25131 6976 25163
rect 7008 25131 7048 25163
rect 7080 25131 7120 25163
rect 7152 25131 7192 25163
rect 7224 25131 7264 25163
rect 7296 25131 7336 25163
rect 7368 25131 7408 25163
rect 7440 25131 7480 25163
rect 7512 25131 7552 25163
rect 7584 25131 7624 25163
rect 7656 25131 7696 25163
rect 7728 25131 7768 25163
rect 7800 25131 7840 25163
rect 7872 25131 7912 25163
rect 7944 25131 7984 25163
rect 8016 25131 8056 25163
rect 8088 25131 8128 25163
rect 8160 25131 8200 25163
rect 8232 25131 8272 25163
rect 8304 25131 8344 25163
rect 8376 25131 8416 25163
rect 8448 25131 8488 25163
rect 8520 25131 8560 25163
rect 8592 25131 8632 25163
rect 8664 25131 8704 25163
rect 8736 25131 8776 25163
rect 8808 25131 8848 25163
rect 8880 25131 8920 25163
rect 8952 25131 8992 25163
rect 9024 25131 9064 25163
rect 9096 25131 9136 25163
rect 9168 25131 9208 25163
rect 9240 25131 9280 25163
rect 9312 25131 9352 25163
rect 9384 25131 9424 25163
rect 9456 25131 9496 25163
rect 9528 25131 9568 25163
rect 9600 25131 9640 25163
rect 9672 25131 9712 25163
rect 9744 25131 9784 25163
rect 9816 25131 9856 25163
rect 9888 25131 9928 25163
rect 9960 25131 10000 25163
rect 10032 25131 10072 25163
rect 10104 25131 10144 25163
rect 10176 25131 10216 25163
rect 10248 25131 10288 25163
rect 10320 25131 10360 25163
rect 10392 25131 10432 25163
rect 10464 25131 10504 25163
rect 10536 25131 10576 25163
rect 10608 25131 10648 25163
rect 10680 25131 10720 25163
rect 10752 25131 10792 25163
rect 10824 25131 10864 25163
rect 10896 25131 10936 25163
rect 10968 25131 11008 25163
rect 11040 25131 11080 25163
rect 11112 25131 11152 25163
rect 11184 25131 11224 25163
rect 11256 25131 11296 25163
rect 11328 25131 11368 25163
rect 11400 25131 11440 25163
rect 11472 25131 11512 25163
rect 11544 25131 11584 25163
rect 11616 25131 11656 25163
rect 11688 25131 11728 25163
rect 11760 25131 11800 25163
rect 11832 25131 11872 25163
rect 11904 25131 11944 25163
rect 11976 25131 12016 25163
rect 12048 25131 12088 25163
rect 12120 25131 12160 25163
rect 12192 25131 12232 25163
rect 12264 25131 12304 25163
rect 12336 25131 12376 25163
rect 12408 25131 12448 25163
rect 12480 25131 12520 25163
rect 12552 25131 12592 25163
rect 12624 25131 12664 25163
rect 12696 25131 12736 25163
rect 12768 25131 12808 25163
rect 12840 25131 12880 25163
rect 12912 25131 12952 25163
rect 12984 25131 13024 25163
rect 13056 25131 13096 25163
rect 13128 25131 13168 25163
rect 13200 25131 13240 25163
rect 13272 25131 13312 25163
rect 13344 25131 13384 25163
rect 13416 25131 13456 25163
rect 13488 25131 13528 25163
rect 13560 25131 13600 25163
rect 13632 25131 13672 25163
rect 13704 25131 13744 25163
rect 13776 25131 13816 25163
rect 13848 25131 13888 25163
rect 13920 25131 13960 25163
rect 13992 25131 14032 25163
rect 14064 25131 14104 25163
rect 14136 25131 14176 25163
rect 14208 25131 14248 25163
rect 14280 25131 14320 25163
rect 14352 25131 14392 25163
rect 14424 25131 14464 25163
rect 14496 25131 14536 25163
rect 14568 25131 14608 25163
rect 14640 25131 14680 25163
rect 14712 25131 14752 25163
rect 14784 25131 14824 25163
rect 14856 25131 14896 25163
rect 14928 25131 14968 25163
rect 15000 25131 15040 25163
rect 15072 25131 15112 25163
rect 15144 25131 15184 25163
rect 15216 25131 15256 25163
rect 15288 25131 15328 25163
rect 15360 25131 15400 25163
rect 15432 25131 15472 25163
rect 15504 25131 15544 25163
rect 15576 25131 15616 25163
rect 15648 25131 15688 25163
rect 15720 25131 15760 25163
rect 15792 25131 15832 25163
rect 15864 25131 15904 25163
rect 15936 25131 16000 25163
rect 0 25091 16000 25131
rect 0 25059 64 25091
rect 96 25059 136 25091
rect 168 25059 208 25091
rect 240 25059 280 25091
rect 312 25059 352 25091
rect 384 25059 424 25091
rect 456 25059 496 25091
rect 528 25059 568 25091
rect 600 25059 640 25091
rect 672 25059 712 25091
rect 744 25059 784 25091
rect 816 25059 856 25091
rect 888 25059 928 25091
rect 960 25059 1000 25091
rect 1032 25059 1072 25091
rect 1104 25059 1144 25091
rect 1176 25059 1216 25091
rect 1248 25059 1288 25091
rect 1320 25059 1360 25091
rect 1392 25059 1432 25091
rect 1464 25059 1504 25091
rect 1536 25059 1576 25091
rect 1608 25059 1648 25091
rect 1680 25059 1720 25091
rect 1752 25059 1792 25091
rect 1824 25059 1864 25091
rect 1896 25059 1936 25091
rect 1968 25059 2008 25091
rect 2040 25059 2080 25091
rect 2112 25059 2152 25091
rect 2184 25059 2224 25091
rect 2256 25059 2296 25091
rect 2328 25059 2368 25091
rect 2400 25059 2440 25091
rect 2472 25059 2512 25091
rect 2544 25059 2584 25091
rect 2616 25059 2656 25091
rect 2688 25059 2728 25091
rect 2760 25059 2800 25091
rect 2832 25059 2872 25091
rect 2904 25059 2944 25091
rect 2976 25059 3016 25091
rect 3048 25059 3088 25091
rect 3120 25059 3160 25091
rect 3192 25059 3232 25091
rect 3264 25059 3304 25091
rect 3336 25059 3376 25091
rect 3408 25059 3448 25091
rect 3480 25059 3520 25091
rect 3552 25059 3592 25091
rect 3624 25059 3664 25091
rect 3696 25059 3736 25091
rect 3768 25059 3808 25091
rect 3840 25059 3880 25091
rect 3912 25059 3952 25091
rect 3984 25059 4024 25091
rect 4056 25059 4096 25091
rect 4128 25059 4168 25091
rect 4200 25059 4240 25091
rect 4272 25059 4312 25091
rect 4344 25059 4384 25091
rect 4416 25059 4456 25091
rect 4488 25059 4528 25091
rect 4560 25059 4600 25091
rect 4632 25059 4672 25091
rect 4704 25059 4744 25091
rect 4776 25059 4816 25091
rect 4848 25059 4888 25091
rect 4920 25059 4960 25091
rect 4992 25059 5032 25091
rect 5064 25059 5104 25091
rect 5136 25059 5176 25091
rect 5208 25059 5248 25091
rect 5280 25059 5320 25091
rect 5352 25059 5392 25091
rect 5424 25059 5464 25091
rect 5496 25059 5536 25091
rect 5568 25059 5608 25091
rect 5640 25059 5680 25091
rect 5712 25059 5752 25091
rect 5784 25059 5824 25091
rect 5856 25059 5896 25091
rect 5928 25059 5968 25091
rect 6000 25059 6040 25091
rect 6072 25059 6112 25091
rect 6144 25059 6184 25091
rect 6216 25059 6256 25091
rect 6288 25059 6328 25091
rect 6360 25059 6400 25091
rect 6432 25059 6472 25091
rect 6504 25059 6544 25091
rect 6576 25059 6616 25091
rect 6648 25059 6688 25091
rect 6720 25059 6760 25091
rect 6792 25059 6832 25091
rect 6864 25059 6904 25091
rect 6936 25059 6976 25091
rect 7008 25059 7048 25091
rect 7080 25059 7120 25091
rect 7152 25059 7192 25091
rect 7224 25059 7264 25091
rect 7296 25059 7336 25091
rect 7368 25059 7408 25091
rect 7440 25059 7480 25091
rect 7512 25059 7552 25091
rect 7584 25059 7624 25091
rect 7656 25059 7696 25091
rect 7728 25059 7768 25091
rect 7800 25059 7840 25091
rect 7872 25059 7912 25091
rect 7944 25059 7984 25091
rect 8016 25059 8056 25091
rect 8088 25059 8128 25091
rect 8160 25059 8200 25091
rect 8232 25059 8272 25091
rect 8304 25059 8344 25091
rect 8376 25059 8416 25091
rect 8448 25059 8488 25091
rect 8520 25059 8560 25091
rect 8592 25059 8632 25091
rect 8664 25059 8704 25091
rect 8736 25059 8776 25091
rect 8808 25059 8848 25091
rect 8880 25059 8920 25091
rect 8952 25059 8992 25091
rect 9024 25059 9064 25091
rect 9096 25059 9136 25091
rect 9168 25059 9208 25091
rect 9240 25059 9280 25091
rect 9312 25059 9352 25091
rect 9384 25059 9424 25091
rect 9456 25059 9496 25091
rect 9528 25059 9568 25091
rect 9600 25059 9640 25091
rect 9672 25059 9712 25091
rect 9744 25059 9784 25091
rect 9816 25059 9856 25091
rect 9888 25059 9928 25091
rect 9960 25059 10000 25091
rect 10032 25059 10072 25091
rect 10104 25059 10144 25091
rect 10176 25059 10216 25091
rect 10248 25059 10288 25091
rect 10320 25059 10360 25091
rect 10392 25059 10432 25091
rect 10464 25059 10504 25091
rect 10536 25059 10576 25091
rect 10608 25059 10648 25091
rect 10680 25059 10720 25091
rect 10752 25059 10792 25091
rect 10824 25059 10864 25091
rect 10896 25059 10936 25091
rect 10968 25059 11008 25091
rect 11040 25059 11080 25091
rect 11112 25059 11152 25091
rect 11184 25059 11224 25091
rect 11256 25059 11296 25091
rect 11328 25059 11368 25091
rect 11400 25059 11440 25091
rect 11472 25059 11512 25091
rect 11544 25059 11584 25091
rect 11616 25059 11656 25091
rect 11688 25059 11728 25091
rect 11760 25059 11800 25091
rect 11832 25059 11872 25091
rect 11904 25059 11944 25091
rect 11976 25059 12016 25091
rect 12048 25059 12088 25091
rect 12120 25059 12160 25091
rect 12192 25059 12232 25091
rect 12264 25059 12304 25091
rect 12336 25059 12376 25091
rect 12408 25059 12448 25091
rect 12480 25059 12520 25091
rect 12552 25059 12592 25091
rect 12624 25059 12664 25091
rect 12696 25059 12736 25091
rect 12768 25059 12808 25091
rect 12840 25059 12880 25091
rect 12912 25059 12952 25091
rect 12984 25059 13024 25091
rect 13056 25059 13096 25091
rect 13128 25059 13168 25091
rect 13200 25059 13240 25091
rect 13272 25059 13312 25091
rect 13344 25059 13384 25091
rect 13416 25059 13456 25091
rect 13488 25059 13528 25091
rect 13560 25059 13600 25091
rect 13632 25059 13672 25091
rect 13704 25059 13744 25091
rect 13776 25059 13816 25091
rect 13848 25059 13888 25091
rect 13920 25059 13960 25091
rect 13992 25059 14032 25091
rect 14064 25059 14104 25091
rect 14136 25059 14176 25091
rect 14208 25059 14248 25091
rect 14280 25059 14320 25091
rect 14352 25059 14392 25091
rect 14424 25059 14464 25091
rect 14496 25059 14536 25091
rect 14568 25059 14608 25091
rect 14640 25059 14680 25091
rect 14712 25059 14752 25091
rect 14784 25059 14824 25091
rect 14856 25059 14896 25091
rect 14928 25059 14968 25091
rect 15000 25059 15040 25091
rect 15072 25059 15112 25091
rect 15144 25059 15184 25091
rect 15216 25059 15256 25091
rect 15288 25059 15328 25091
rect 15360 25059 15400 25091
rect 15432 25059 15472 25091
rect 15504 25059 15544 25091
rect 15576 25059 15616 25091
rect 15648 25059 15688 25091
rect 15720 25059 15760 25091
rect 15792 25059 15832 25091
rect 15864 25059 15904 25091
rect 15936 25059 16000 25091
rect 0 25019 16000 25059
rect 0 24987 64 25019
rect 96 24987 136 25019
rect 168 24987 208 25019
rect 240 24987 280 25019
rect 312 24987 352 25019
rect 384 24987 424 25019
rect 456 24987 496 25019
rect 528 24987 568 25019
rect 600 24987 640 25019
rect 672 24987 712 25019
rect 744 24987 784 25019
rect 816 24987 856 25019
rect 888 24987 928 25019
rect 960 24987 1000 25019
rect 1032 24987 1072 25019
rect 1104 24987 1144 25019
rect 1176 24987 1216 25019
rect 1248 24987 1288 25019
rect 1320 24987 1360 25019
rect 1392 24987 1432 25019
rect 1464 24987 1504 25019
rect 1536 24987 1576 25019
rect 1608 24987 1648 25019
rect 1680 24987 1720 25019
rect 1752 24987 1792 25019
rect 1824 24987 1864 25019
rect 1896 24987 1936 25019
rect 1968 24987 2008 25019
rect 2040 24987 2080 25019
rect 2112 24987 2152 25019
rect 2184 24987 2224 25019
rect 2256 24987 2296 25019
rect 2328 24987 2368 25019
rect 2400 24987 2440 25019
rect 2472 24987 2512 25019
rect 2544 24987 2584 25019
rect 2616 24987 2656 25019
rect 2688 24987 2728 25019
rect 2760 24987 2800 25019
rect 2832 24987 2872 25019
rect 2904 24987 2944 25019
rect 2976 24987 3016 25019
rect 3048 24987 3088 25019
rect 3120 24987 3160 25019
rect 3192 24987 3232 25019
rect 3264 24987 3304 25019
rect 3336 24987 3376 25019
rect 3408 24987 3448 25019
rect 3480 24987 3520 25019
rect 3552 24987 3592 25019
rect 3624 24987 3664 25019
rect 3696 24987 3736 25019
rect 3768 24987 3808 25019
rect 3840 24987 3880 25019
rect 3912 24987 3952 25019
rect 3984 24987 4024 25019
rect 4056 24987 4096 25019
rect 4128 24987 4168 25019
rect 4200 24987 4240 25019
rect 4272 24987 4312 25019
rect 4344 24987 4384 25019
rect 4416 24987 4456 25019
rect 4488 24987 4528 25019
rect 4560 24987 4600 25019
rect 4632 24987 4672 25019
rect 4704 24987 4744 25019
rect 4776 24987 4816 25019
rect 4848 24987 4888 25019
rect 4920 24987 4960 25019
rect 4992 24987 5032 25019
rect 5064 24987 5104 25019
rect 5136 24987 5176 25019
rect 5208 24987 5248 25019
rect 5280 24987 5320 25019
rect 5352 24987 5392 25019
rect 5424 24987 5464 25019
rect 5496 24987 5536 25019
rect 5568 24987 5608 25019
rect 5640 24987 5680 25019
rect 5712 24987 5752 25019
rect 5784 24987 5824 25019
rect 5856 24987 5896 25019
rect 5928 24987 5968 25019
rect 6000 24987 6040 25019
rect 6072 24987 6112 25019
rect 6144 24987 6184 25019
rect 6216 24987 6256 25019
rect 6288 24987 6328 25019
rect 6360 24987 6400 25019
rect 6432 24987 6472 25019
rect 6504 24987 6544 25019
rect 6576 24987 6616 25019
rect 6648 24987 6688 25019
rect 6720 24987 6760 25019
rect 6792 24987 6832 25019
rect 6864 24987 6904 25019
rect 6936 24987 6976 25019
rect 7008 24987 7048 25019
rect 7080 24987 7120 25019
rect 7152 24987 7192 25019
rect 7224 24987 7264 25019
rect 7296 24987 7336 25019
rect 7368 24987 7408 25019
rect 7440 24987 7480 25019
rect 7512 24987 7552 25019
rect 7584 24987 7624 25019
rect 7656 24987 7696 25019
rect 7728 24987 7768 25019
rect 7800 24987 7840 25019
rect 7872 24987 7912 25019
rect 7944 24987 7984 25019
rect 8016 24987 8056 25019
rect 8088 24987 8128 25019
rect 8160 24987 8200 25019
rect 8232 24987 8272 25019
rect 8304 24987 8344 25019
rect 8376 24987 8416 25019
rect 8448 24987 8488 25019
rect 8520 24987 8560 25019
rect 8592 24987 8632 25019
rect 8664 24987 8704 25019
rect 8736 24987 8776 25019
rect 8808 24987 8848 25019
rect 8880 24987 8920 25019
rect 8952 24987 8992 25019
rect 9024 24987 9064 25019
rect 9096 24987 9136 25019
rect 9168 24987 9208 25019
rect 9240 24987 9280 25019
rect 9312 24987 9352 25019
rect 9384 24987 9424 25019
rect 9456 24987 9496 25019
rect 9528 24987 9568 25019
rect 9600 24987 9640 25019
rect 9672 24987 9712 25019
rect 9744 24987 9784 25019
rect 9816 24987 9856 25019
rect 9888 24987 9928 25019
rect 9960 24987 10000 25019
rect 10032 24987 10072 25019
rect 10104 24987 10144 25019
rect 10176 24987 10216 25019
rect 10248 24987 10288 25019
rect 10320 24987 10360 25019
rect 10392 24987 10432 25019
rect 10464 24987 10504 25019
rect 10536 24987 10576 25019
rect 10608 24987 10648 25019
rect 10680 24987 10720 25019
rect 10752 24987 10792 25019
rect 10824 24987 10864 25019
rect 10896 24987 10936 25019
rect 10968 24987 11008 25019
rect 11040 24987 11080 25019
rect 11112 24987 11152 25019
rect 11184 24987 11224 25019
rect 11256 24987 11296 25019
rect 11328 24987 11368 25019
rect 11400 24987 11440 25019
rect 11472 24987 11512 25019
rect 11544 24987 11584 25019
rect 11616 24987 11656 25019
rect 11688 24987 11728 25019
rect 11760 24987 11800 25019
rect 11832 24987 11872 25019
rect 11904 24987 11944 25019
rect 11976 24987 12016 25019
rect 12048 24987 12088 25019
rect 12120 24987 12160 25019
rect 12192 24987 12232 25019
rect 12264 24987 12304 25019
rect 12336 24987 12376 25019
rect 12408 24987 12448 25019
rect 12480 24987 12520 25019
rect 12552 24987 12592 25019
rect 12624 24987 12664 25019
rect 12696 24987 12736 25019
rect 12768 24987 12808 25019
rect 12840 24987 12880 25019
rect 12912 24987 12952 25019
rect 12984 24987 13024 25019
rect 13056 24987 13096 25019
rect 13128 24987 13168 25019
rect 13200 24987 13240 25019
rect 13272 24987 13312 25019
rect 13344 24987 13384 25019
rect 13416 24987 13456 25019
rect 13488 24987 13528 25019
rect 13560 24987 13600 25019
rect 13632 24987 13672 25019
rect 13704 24987 13744 25019
rect 13776 24987 13816 25019
rect 13848 24987 13888 25019
rect 13920 24987 13960 25019
rect 13992 24987 14032 25019
rect 14064 24987 14104 25019
rect 14136 24987 14176 25019
rect 14208 24987 14248 25019
rect 14280 24987 14320 25019
rect 14352 24987 14392 25019
rect 14424 24987 14464 25019
rect 14496 24987 14536 25019
rect 14568 24987 14608 25019
rect 14640 24987 14680 25019
rect 14712 24987 14752 25019
rect 14784 24987 14824 25019
rect 14856 24987 14896 25019
rect 14928 24987 14968 25019
rect 15000 24987 15040 25019
rect 15072 24987 15112 25019
rect 15144 24987 15184 25019
rect 15216 24987 15256 25019
rect 15288 24987 15328 25019
rect 15360 24987 15400 25019
rect 15432 24987 15472 25019
rect 15504 24987 15544 25019
rect 15576 24987 15616 25019
rect 15648 24987 15688 25019
rect 15720 24987 15760 25019
rect 15792 24987 15832 25019
rect 15864 24987 15904 25019
rect 15936 24987 16000 25019
rect 0 24947 16000 24987
rect 0 24915 64 24947
rect 96 24915 136 24947
rect 168 24915 208 24947
rect 240 24915 280 24947
rect 312 24915 352 24947
rect 384 24915 424 24947
rect 456 24915 496 24947
rect 528 24915 568 24947
rect 600 24915 640 24947
rect 672 24915 712 24947
rect 744 24915 784 24947
rect 816 24915 856 24947
rect 888 24915 928 24947
rect 960 24915 1000 24947
rect 1032 24915 1072 24947
rect 1104 24915 1144 24947
rect 1176 24915 1216 24947
rect 1248 24915 1288 24947
rect 1320 24915 1360 24947
rect 1392 24915 1432 24947
rect 1464 24915 1504 24947
rect 1536 24915 1576 24947
rect 1608 24915 1648 24947
rect 1680 24915 1720 24947
rect 1752 24915 1792 24947
rect 1824 24915 1864 24947
rect 1896 24915 1936 24947
rect 1968 24915 2008 24947
rect 2040 24915 2080 24947
rect 2112 24915 2152 24947
rect 2184 24915 2224 24947
rect 2256 24915 2296 24947
rect 2328 24915 2368 24947
rect 2400 24915 2440 24947
rect 2472 24915 2512 24947
rect 2544 24915 2584 24947
rect 2616 24915 2656 24947
rect 2688 24915 2728 24947
rect 2760 24915 2800 24947
rect 2832 24915 2872 24947
rect 2904 24915 2944 24947
rect 2976 24915 3016 24947
rect 3048 24915 3088 24947
rect 3120 24915 3160 24947
rect 3192 24915 3232 24947
rect 3264 24915 3304 24947
rect 3336 24915 3376 24947
rect 3408 24915 3448 24947
rect 3480 24915 3520 24947
rect 3552 24915 3592 24947
rect 3624 24915 3664 24947
rect 3696 24915 3736 24947
rect 3768 24915 3808 24947
rect 3840 24915 3880 24947
rect 3912 24915 3952 24947
rect 3984 24915 4024 24947
rect 4056 24915 4096 24947
rect 4128 24915 4168 24947
rect 4200 24915 4240 24947
rect 4272 24915 4312 24947
rect 4344 24915 4384 24947
rect 4416 24915 4456 24947
rect 4488 24915 4528 24947
rect 4560 24915 4600 24947
rect 4632 24915 4672 24947
rect 4704 24915 4744 24947
rect 4776 24915 4816 24947
rect 4848 24915 4888 24947
rect 4920 24915 4960 24947
rect 4992 24915 5032 24947
rect 5064 24915 5104 24947
rect 5136 24915 5176 24947
rect 5208 24915 5248 24947
rect 5280 24915 5320 24947
rect 5352 24915 5392 24947
rect 5424 24915 5464 24947
rect 5496 24915 5536 24947
rect 5568 24915 5608 24947
rect 5640 24915 5680 24947
rect 5712 24915 5752 24947
rect 5784 24915 5824 24947
rect 5856 24915 5896 24947
rect 5928 24915 5968 24947
rect 6000 24915 6040 24947
rect 6072 24915 6112 24947
rect 6144 24915 6184 24947
rect 6216 24915 6256 24947
rect 6288 24915 6328 24947
rect 6360 24915 6400 24947
rect 6432 24915 6472 24947
rect 6504 24915 6544 24947
rect 6576 24915 6616 24947
rect 6648 24915 6688 24947
rect 6720 24915 6760 24947
rect 6792 24915 6832 24947
rect 6864 24915 6904 24947
rect 6936 24915 6976 24947
rect 7008 24915 7048 24947
rect 7080 24915 7120 24947
rect 7152 24915 7192 24947
rect 7224 24915 7264 24947
rect 7296 24915 7336 24947
rect 7368 24915 7408 24947
rect 7440 24915 7480 24947
rect 7512 24915 7552 24947
rect 7584 24915 7624 24947
rect 7656 24915 7696 24947
rect 7728 24915 7768 24947
rect 7800 24915 7840 24947
rect 7872 24915 7912 24947
rect 7944 24915 7984 24947
rect 8016 24915 8056 24947
rect 8088 24915 8128 24947
rect 8160 24915 8200 24947
rect 8232 24915 8272 24947
rect 8304 24915 8344 24947
rect 8376 24915 8416 24947
rect 8448 24915 8488 24947
rect 8520 24915 8560 24947
rect 8592 24915 8632 24947
rect 8664 24915 8704 24947
rect 8736 24915 8776 24947
rect 8808 24915 8848 24947
rect 8880 24915 8920 24947
rect 8952 24915 8992 24947
rect 9024 24915 9064 24947
rect 9096 24915 9136 24947
rect 9168 24915 9208 24947
rect 9240 24915 9280 24947
rect 9312 24915 9352 24947
rect 9384 24915 9424 24947
rect 9456 24915 9496 24947
rect 9528 24915 9568 24947
rect 9600 24915 9640 24947
rect 9672 24915 9712 24947
rect 9744 24915 9784 24947
rect 9816 24915 9856 24947
rect 9888 24915 9928 24947
rect 9960 24915 10000 24947
rect 10032 24915 10072 24947
rect 10104 24915 10144 24947
rect 10176 24915 10216 24947
rect 10248 24915 10288 24947
rect 10320 24915 10360 24947
rect 10392 24915 10432 24947
rect 10464 24915 10504 24947
rect 10536 24915 10576 24947
rect 10608 24915 10648 24947
rect 10680 24915 10720 24947
rect 10752 24915 10792 24947
rect 10824 24915 10864 24947
rect 10896 24915 10936 24947
rect 10968 24915 11008 24947
rect 11040 24915 11080 24947
rect 11112 24915 11152 24947
rect 11184 24915 11224 24947
rect 11256 24915 11296 24947
rect 11328 24915 11368 24947
rect 11400 24915 11440 24947
rect 11472 24915 11512 24947
rect 11544 24915 11584 24947
rect 11616 24915 11656 24947
rect 11688 24915 11728 24947
rect 11760 24915 11800 24947
rect 11832 24915 11872 24947
rect 11904 24915 11944 24947
rect 11976 24915 12016 24947
rect 12048 24915 12088 24947
rect 12120 24915 12160 24947
rect 12192 24915 12232 24947
rect 12264 24915 12304 24947
rect 12336 24915 12376 24947
rect 12408 24915 12448 24947
rect 12480 24915 12520 24947
rect 12552 24915 12592 24947
rect 12624 24915 12664 24947
rect 12696 24915 12736 24947
rect 12768 24915 12808 24947
rect 12840 24915 12880 24947
rect 12912 24915 12952 24947
rect 12984 24915 13024 24947
rect 13056 24915 13096 24947
rect 13128 24915 13168 24947
rect 13200 24915 13240 24947
rect 13272 24915 13312 24947
rect 13344 24915 13384 24947
rect 13416 24915 13456 24947
rect 13488 24915 13528 24947
rect 13560 24915 13600 24947
rect 13632 24915 13672 24947
rect 13704 24915 13744 24947
rect 13776 24915 13816 24947
rect 13848 24915 13888 24947
rect 13920 24915 13960 24947
rect 13992 24915 14032 24947
rect 14064 24915 14104 24947
rect 14136 24915 14176 24947
rect 14208 24915 14248 24947
rect 14280 24915 14320 24947
rect 14352 24915 14392 24947
rect 14424 24915 14464 24947
rect 14496 24915 14536 24947
rect 14568 24915 14608 24947
rect 14640 24915 14680 24947
rect 14712 24915 14752 24947
rect 14784 24915 14824 24947
rect 14856 24915 14896 24947
rect 14928 24915 14968 24947
rect 15000 24915 15040 24947
rect 15072 24915 15112 24947
rect 15144 24915 15184 24947
rect 15216 24915 15256 24947
rect 15288 24915 15328 24947
rect 15360 24915 15400 24947
rect 15432 24915 15472 24947
rect 15504 24915 15544 24947
rect 15576 24915 15616 24947
rect 15648 24915 15688 24947
rect 15720 24915 15760 24947
rect 15792 24915 15832 24947
rect 15864 24915 15904 24947
rect 15936 24915 16000 24947
rect 0 24875 16000 24915
rect 0 24843 64 24875
rect 96 24843 136 24875
rect 168 24843 208 24875
rect 240 24843 280 24875
rect 312 24843 352 24875
rect 384 24843 424 24875
rect 456 24843 496 24875
rect 528 24843 568 24875
rect 600 24843 640 24875
rect 672 24843 712 24875
rect 744 24843 784 24875
rect 816 24843 856 24875
rect 888 24843 928 24875
rect 960 24843 1000 24875
rect 1032 24843 1072 24875
rect 1104 24843 1144 24875
rect 1176 24843 1216 24875
rect 1248 24843 1288 24875
rect 1320 24843 1360 24875
rect 1392 24843 1432 24875
rect 1464 24843 1504 24875
rect 1536 24843 1576 24875
rect 1608 24843 1648 24875
rect 1680 24843 1720 24875
rect 1752 24843 1792 24875
rect 1824 24843 1864 24875
rect 1896 24843 1936 24875
rect 1968 24843 2008 24875
rect 2040 24843 2080 24875
rect 2112 24843 2152 24875
rect 2184 24843 2224 24875
rect 2256 24843 2296 24875
rect 2328 24843 2368 24875
rect 2400 24843 2440 24875
rect 2472 24843 2512 24875
rect 2544 24843 2584 24875
rect 2616 24843 2656 24875
rect 2688 24843 2728 24875
rect 2760 24843 2800 24875
rect 2832 24843 2872 24875
rect 2904 24843 2944 24875
rect 2976 24843 3016 24875
rect 3048 24843 3088 24875
rect 3120 24843 3160 24875
rect 3192 24843 3232 24875
rect 3264 24843 3304 24875
rect 3336 24843 3376 24875
rect 3408 24843 3448 24875
rect 3480 24843 3520 24875
rect 3552 24843 3592 24875
rect 3624 24843 3664 24875
rect 3696 24843 3736 24875
rect 3768 24843 3808 24875
rect 3840 24843 3880 24875
rect 3912 24843 3952 24875
rect 3984 24843 4024 24875
rect 4056 24843 4096 24875
rect 4128 24843 4168 24875
rect 4200 24843 4240 24875
rect 4272 24843 4312 24875
rect 4344 24843 4384 24875
rect 4416 24843 4456 24875
rect 4488 24843 4528 24875
rect 4560 24843 4600 24875
rect 4632 24843 4672 24875
rect 4704 24843 4744 24875
rect 4776 24843 4816 24875
rect 4848 24843 4888 24875
rect 4920 24843 4960 24875
rect 4992 24843 5032 24875
rect 5064 24843 5104 24875
rect 5136 24843 5176 24875
rect 5208 24843 5248 24875
rect 5280 24843 5320 24875
rect 5352 24843 5392 24875
rect 5424 24843 5464 24875
rect 5496 24843 5536 24875
rect 5568 24843 5608 24875
rect 5640 24843 5680 24875
rect 5712 24843 5752 24875
rect 5784 24843 5824 24875
rect 5856 24843 5896 24875
rect 5928 24843 5968 24875
rect 6000 24843 6040 24875
rect 6072 24843 6112 24875
rect 6144 24843 6184 24875
rect 6216 24843 6256 24875
rect 6288 24843 6328 24875
rect 6360 24843 6400 24875
rect 6432 24843 6472 24875
rect 6504 24843 6544 24875
rect 6576 24843 6616 24875
rect 6648 24843 6688 24875
rect 6720 24843 6760 24875
rect 6792 24843 6832 24875
rect 6864 24843 6904 24875
rect 6936 24843 6976 24875
rect 7008 24843 7048 24875
rect 7080 24843 7120 24875
rect 7152 24843 7192 24875
rect 7224 24843 7264 24875
rect 7296 24843 7336 24875
rect 7368 24843 7408 24875
rect 7440 24843 7480 24875
rect 7512 24843 7552 24875
rect 7584 24843 7624 24875
rect 7656 24843 7696 24875
rect 7728 24843 7768 24875
rect 7800 24843 7840 24875
rect 7872 24843 7912 24875
rect 7944 24843 7984 24875
rect 8016 24843 8056 24875
rect 8088 24843 8128 24875
rect 8160 24843 8200 24875
rect 8232 24843 8272 24875
rect 8304 24843 8344 24875
rect 8376 24843 8416 24875
rect 8448 24843 8488 24875
rect 8520 24843 8560 24875
rect 8592 24843 8632 24875
rect 8664 24843 8704 24875
rect 8736 24843 8776 24875
rect 8808 24843 8848 24875
rect 8880 24843 8920 24875
rect 8952 24843 8992 24875
rect 9024 24843 9064 24875
rect 9096 24843 9136 24875
rect 9168 24843 9208 24875
rect 9240 24843 9280 24875
rect 9312 24843 9352 24875
rect 9384 24843 9424 24875
rect 9456 24843 9496 24875
rect 9528 24843 9568 24875
rect 9600 24843 9640 24875
rect 9672 24843 9712 24875
rect 9744 24843 9784 24875
rect 9816 24843 9856 24875
rect 9888 24843 9928 24875
rect 9960 24843 10000 24875
rect 10032 24843 10072 24875
rect 10104 24843 10144 24875
rect 10176 24843 10216 24875
rect 10248 24843 10288 24875
rect 10320 24843 10360 24875
rect 10392 24843 10432 24875
rect 10464 24843 10504 24875
rect 10536 24843 10576 24875
rect 10608 24843 10648 24875
rect 10680 24843 10720 24875
rect 10752 24843 10792 24875
rect 10824 24843 10864 24875
rect 10896 24843 10936 24875
rect 10968 24843 11008 24875
rect 11040 24843 11080 24875
rect 11112 24843 11152 24875
rect 11184 24843 11224 24875
rect 11256 24843 11296 24875
rect 11328 24843 11368 24875
rect 11400 24843 11440 24875
rect 11472 24843 11512 24875
rect 11544 24843 11584 24875
rect 11616 24843 11656 24875
rect 11688 24843 11728 24875
rect 11760 24843 11800 24875
rect 11832 24843 11872 24875
rect 11904 24843 11944 24875
rect 11976 24843 12016 24875
rect 12048 24843 12088 24875
rect 12120 24843 12160 24875
rect 12192 24843 12232 24875
rect 12264 24843 12304 24875
rect 12336 24843 12376 24875
rect 12408 24843 12448 24875
rect 12480 24843 12520 24875
rect 12552 24843 12592 24875
rect 12624 24843 12664 24875
rect 12696 24843 12736 24875
rect 12768 24843 12808 24875
rect 12840 24843 12880 24875
rect 12912 24843 12952 24875
rect 12984 24843 13024 24875
rect 13056 24843 13096 24875
rect 13128 24843 13168 24875
rect 13200 24843 13240 24875
rect 13272 24843 13312 24875
rect 13344 24843 13384 24875
rect 13416 24843 13456 24875
rect 13488 24843 13528 24875
rect 13560 24843 13600 24875
rect 13632 24843 13672 24875
rect 13704 24843 13744 24875
rect 13776 24843 13816 24875
rect 13848 24843 13888 24875
rect 13920 24843 13960 24875
rect 13992 24843 14032 24875
rect 14064 24843 14104 24875
rect 14136 24843 14176 24875
rect 14208 24843 14248 24875
rect 14280 24843 14320 24875
rect 14352 24843 14392 24875
rect 14424 24843 14464 24875
rect 14496 24843 14536 24875
rect 14568 24843 14608 24875
rect 14640 24843 14680 24875
rect 14712 24843 14752 24875
rect 14784 24843 14824 24875
rect 14856 24843 14896 24875
rect 14928 24843 14968 24875
rect 15000 24843 15040 24875
rect 15072 24843 15112 24875
rect 15144 24843 15184 24875
rect 15216 24843 15256 24875
rect 15288 24843 15328 24875
rect 15360 24843 15400 24875
rect 15432 24843 15472 24875
rect 15504 24843 15544 24875
rect 15576 24843 15616 24875
rect 15648 24843 15688 24875
rect 15720 24843 15760 24875
rect 15792 24843 15832 24875
rect 15864 24843 15904 24875
rect 15936 24843 16000 24875
rect 0 24803 16000 24843
rect 0 24771 64 24803
rect 96 24771 136 24803
rect 168 24771 208 24803
rect 240 24771 280 24803
rect 312 24771 352 24803
rect 384 24771 424 24803
rect 456 24771 496 24803
rect 528 24771 568 24803
rect 600 24771 640 24803
rect 672 24771 712 24803
rect 744 24771 784 24803
rect 816 24771 856 24803
rect 888 24771 928 24803
rect 960 24771 1000 24803
rect 1032 24771 1072 24803
rect 1104 24771 1144 24803
rect 1176 24771 1216 24803
rect 1248 24771 1288 24803
rect 1320 24771 1360 24803
rect 1392 24771 1432 24803
rect 1464 24771 1504 24803
rect 1536 24771 1576 24803
rect 1608 24771 1648 24803
rect 1680 24771 1720 24803
rect 1752 24771 1792 24803
rect 1824 24771 1864 24803
rect 1896 24771 1936 24803
rect 1968 24771 2008 24803
rect 2040 24771 2080 24803
rect 2112 24771 2152 24803
rect 2184 24771 2224 24803
rect 2256 24771 2296 24803
rect 2328 24771 2368 24803
rect 2400 24771 2440 24803
rect 2472 24771 2512 24803
rect 2544 24771 2584 24803
rect 2616 24771 2656 24803
rect 2688 24771 2728 24803
rect 2760 24771 2800 24803
rect 2832 24771 2872 24803
rect 2904 24771 2944 24803
rect 2976 24771 3016 24803
rect 3048 24771 3088 24803
rect 3120 24771 3160 24803
rect 3192 24771 3232 24803
rect 3264 24771 3304 24803
rect 3336 24771 3376 24803
rect 3408 24771 3448 24803
rect 3480 24771 3520 24803
rect 3552 24771 3592 24803
rect 3624 24771 3664 24803
rect 3696 24771 3736 24803
rect 3768 24771 3808 24803
rect 3840 24771 3880 24803
rect 3912 24771 3952 24803
rect 3984 24771 4024 24803
rect 4056 24771 4096 24803
rect 4128 24771 4168 24803
rect 4200 24771 4240 24803
rect 4272 24771 4312 24803
rect 4344 24771 4384 24803
rect 4416 24771 4456 24803
rect 4488 24771 4528 24803
rect 4560 24771 4600 24803
rect 4632 24771 4672 24803
rect 4704 24771 4744 24803
rect 4776 24771 4816 24803
rect 4848 24771 4888 24803
rect 4920 24771 4960 24803
rect 4992 24771 5032 24803
rect 5064 24771 5104 24803
rect 5136 24771 5176 24803
rect 5208 24771 5248 24803
rect 5280 24771 5320 24803
rect 5352 24771 5392 24803
rect 5424 24771 5464 24803
rect 5496 24771 5536 24803
rect 5568 24771 5608 24803
rect 5640 24771 5680 24803
rect 5712 24771 5752 24803
rect 5784 24771 5824 24803
rect 5856 24771 5896 24803
rect 5928 24771 5968 24803
rect 6000 24771 6040 24803
rect 6072 24771 6112 24803
rect 6144 24771 6184 24803
rect 6216 24771 6256 24803
rect 6288 24771 6328 24803
rect 6360 24771 6400 24803
rect 6432 24771 6472 24803
rect 6504 24771 6544 24803
rect 6576 24771 6616 24803
rect 6648 24771 6688 24803
rect 6720 24771 6760 24803
rect 6792 24771 6832 24803
rect 6864 24771 6904 24803
rect 6936 24771 6976 24803
rect 7008 24771 7048 24803
rect 7080 24771 7120 24803
rect 7152 24771 7192 24803
rect 7224 24771 7264 24803
rect 7296 24771 7336 24803
rect 7368 24771 7408 24803
rect 7440 24771 7480 24803
rect 7512 24771 7552 24803
rect 7584 24771 7624 24803
rect 7656 24771 7696 24803
rect 7728 24771 7768 24803
rect 7800 24771 7840 24803
rect 7872 24771 7912 24803
rect 7944 24771 7984 24803
rect 8016 24771 8056 24803
rect 8088 24771 8128 24803
rect 8160 24771 8200 24803
rect 8232 24771 8272 24803
rect 8304 24771 8344 24803
rect 8376 24771 8416 24803
rect 8448 24771 8488 24803
rect 8520 24771 8560 24803
rect 8592 24771 8632 24803
rect 8664 24771 8704 24803
rect 8736 24771 8776 24803
rect 8808 24771 8848 24803
rect 8880 24771 8920 24803
rect 8952 24771 8992 24803
rect 9024 24771 9064 24803
rect 9096 24771 9136 24803
rect 9168 24771 9208 24803
rect 9240 24771 9280 24803
rect 9312 24771 9352 24803
rect 9384 24771 9424 24803
rect 9456 24771 9496 24803
rect 9528 24771 9568 24803
rect 9600 24771 9640 24803
rect 9672 24771 9712 24803
rect 9744 24771 9784 24803
rect 9816 24771 9856 24803
rect 9888 24771 9928 24803
rect 9960 24771 10000 24803
rect 10032 24771 10072 24803
rect 10104 24771 10144 24803
rect 10176 24771 10216 24803
rect 10248 24771 10288 24803
rect 10320 24771 10360 24803
rect 10392 24771 10432 24803
rect 10464 24771 10504 24803
rect 10536 24771 10576 24803
rect 10608 24771 10648 24803
rect 10680 24771 10720 24803
rect 10752 24771 10792 24803
rect 10824 24771 10864 24803
rect 10896 24771 10936 24803
rect 10968 24771 11008 24803
rect 11040 24771 11080 24803
rect 11112 24771 11152 24803
rect 11184 24771 11224 24803
rect 11256 24771 11296 24803
rect 11328 24771 11368 24803
rect 11400 24771 11440 24803
rect 11472 24771 11512 24803
rect 11544 24771 11584 24803
rect 11616 24771 11656 24803
rect 11688 24771 11728 24803
rect 11760 24771 11800 24803
rect 11832 24771 11872 24803
rect 11904 24771 11944 24803
rect 11976 24771 12016 24803
rect 12048 24771 12088 24803
rect 12120 24771 12160 24803
rect 12192 24771 12232 24803
rect 12264 24771 12304 24803
rect 12336 24771 12376 24803
rect 12408 24771 12448 24803
rect 12480 24771 12520 24803
rect 12552 24771 12592 24803
rect 12624 24771 12664 24803
rect 12696 24771 12736 24803
rect 12768 24771 12808 24803
rect 12840 24771 12880 24803
rect 12912 24771 12952 24803
rect 12984 24771 13024 24803
rect 13056 24771 13096 24803
rect 13128 24771 13168 24803
rect 13200 24771 13240 24803
rect 13272 24771 13312 24803
rect 13344 24771 13384 24803
rect 13416 24771 13456 24803
rect 13488 24771 13528 24803
rect 13560 24771 13600 24803
rect 13632 24771 13672 24803
rect 13704 24771 13744 24803
rect 13776 24771 13816 24803
rect 13848 24771 13888 24803
rect 13920 24771 13960 24803
rect 13992 24771 14032 24803
rect 14064 24771 14104 24803
rect 14136 24771 14176 24803
rect 14208 24771 14248 24803
rect 14280 24771 14320 24803
rect 14352 24771 14392 24803
rect 14424 24771 14464 24803
rect 14496 24771 14536 24803
rect 14568 24771 14608 24803
rect 14640 24771 14680 24803
rect 14712 24771 14752 24803
rect 14784 24771 14824 24803
rect 14856 24771 14896 24803
rect 14928 24771 14968 24803
rect 15000 24771 15040 24803
rect 15072 24771 15112 24803
rect 15144 24771 15184 24803
rect 15216 24771 15256 24803
rect 15288 24771 15328 24803
rect 15360 24771 15400 24803
rect 15432 24771 15472 24803
rect 15504 24771 15544 24803
rect 15576 24771 15616 24803
rect 15648 24771 15688 24803
rect 15720 24771 15760 24803
rect 15792 24771 15832 24803
rect 15864 24771 15904 24803
rect 15936 24771 16000 24803
rect 0 24731 16000 24771
rect 0 24699 64 24731
rect 96 24699 136 24731
rect 168 24699 208 24731
rect 240 24699 280 24731
rect 312 24699 352 24731
rect 384 24699 424 24731
rect 456 24699 496 24731
rect 528 24699 568 24731
rect 600 24699 640 24731
rect 672 24699 712 24731
rect 744 24699 784 24731
rect 816 24699 856 24731
rect 888 24699 928 24731
rect 960 24699 1000 24731
rect 1032 24699 1072 24731
rect 1104 24699 1144 24731
rect 1176 24699 1216 24731
rect 1248 24699 1288 24731
rect 1320 24699 1360 24731
rect 1392 24699 1432 24731
rect 1464 24699 1504 24731
rect 1536 24699 1576 24731
rect 1608 24699 1648 24731
rect 1680 24699 1720 24731
rect 1752 24699 1792 24731
rect 1824 24699 1864 24731
rect 1896 24699 1936 24731
rect 1968 24699 2008 24731
rect 2040 24699 2080 24731
rect 2112 24699 2152 24731
rect 2184 24699 2224 24731
rect 2256 24699 2296 24731
rect 2328 24699 2368 24731
rect 2400 24699 2440 24731
rect 2472 24699 2512 24731
rect 2544 24699 2584 24731
rect 2616 24699 2656 24731
rect 2688 24699 2728 24731
rect 2760 24699 2800 24731
rect 2832 24699 2872 24731
rect 2904 24699 2944 24731
rect 2976 24699 3016 24731
rect 3048 24699 3088 24731
rect 3120 24699 3160 24731
rect 3192 24699 3232 24731
rect 3264 24699 3304 24731
rect 3336 24699 3376 24731
rect 3408 24699 3448 24731
rect 3480 24699 3520 24731
rect 3552 24699 3592 24731
rect 3624 24699 3664 24731
rect 3696 24699 3736 24731
rect 3768 24699 3808 24731
rect 3840 24699 3880 24731
rect 3912 24699 3952 24731
rect 3984 24699 4024 24731
rect 4056 24699 4096 24731
rect 4128 24699 4168 24731
rect 4200 24699 4240 24731
rect 4272 24699 4312 24731
rect 4344 24699 4384 24731
rect 4416 24699 4456 24731
rect 4488 24699 4528 24731
rect 4560 24699 4600 24731
rect 4632 24699 4672 24731
rect 4704 24699 4744 24731
rect 4776 24699 4816 24731
rect 4848 24699 4888 24731
rect 4920 24699 4960 24731
rect 4992 24699 5032 24731
rect 5064 24699 5104 24731
rect 5136 24699 5176 24731
rect 5208 24699 5248 24731
rect 5280 24699 5320 24731
rect 5352 24699 5392 24731
rect 5424 24699 5464 24731
rect 5496 24699 5536 24731
rect 5568 24699 5608 24731
rect 5640 24699 5680 24731
rect 5712 24699 5752 24731
rect 5784 24699 5824 24731
rect 5856 24699 5896 24731
rect 5928 24699 5968 24731
rect 6000 24699 6040 24731
rect 6072 24699 6112 24731
rect 6144 24699 6184 24731
rect 6216 24699 6256 24731
rect 6288 24699 6328 24731
rect 6360 24699 6400 24731
rect 6432 24699 6472 24731
rect 6504 24699 6544 24731
rect 6576 24699 6616 24731
rect 6648 24699 6688 24731
rect 6720 24699 6760 24731
rect 6792 24699 6832 24731
rect 6864 24699 6904 24731
rect 6936 24699 6976 24731
rect 7008 24699 7048 24731
rect 7080 24699 7120 24731
rect 7152 24699 7192 24731
rect 7224 24699 7264 24731
rect 7296 24699 7336 24731
rect 7368 24699 7408 24731
rect 7440 24699 7480 24731
rect 7512 24699 7552 24731
rect 7584 24699 7624 24731
rect 7656 24699 7696 24731
rect 7728 24699 7768 24731
rect 7800 24699 7840 24731
rect 7872 24699 7912 24731
rect 7944 24699 7984 24731
rect 8016 24699 8056 24731
rect 8088 24699 8128 24731
rect 8160 24699 8200 24731
rect 8232 24699 8272 24731
rect 8304 24699 8344 24731
rect 8376 24699 8416 24731
rect 8448 24699 8488 24731
rect 8520 24699 8560 24731
rect 8592 24699 8632 24731
rect 8664 24699 8704 24731
rect 8736 24699 8776 24731
rect 8808 24699 8848 24731
rect 8880 24699 8920 24731
rect 8952 24699 8992 24731
rect 9024 24699 9064 24731
rect 9096 24699 9136 24731
rect 9168 24699 9208 24731
rect 9240 24699 9280 24731
rect 9312 24699 9352 24731
rect 9384 24699 9424 24731
rect 9456 24699 9496 24731
rect 9528 24699 9568 24731
rect 9600 24699 9640 24731
rect 9672 24699 9712 24731
rect 9744 24699 9784 24731
rect 9816 24699 9856 24731
rect 9888 24699 9928 24731
rect 9960 24699 10000 24731
rect 10032 24699 10072 24731
rect 10104 24699 10144 24731
rect 10176 24699 10216 24731
rect 10248 24699 10288 24731
rect 10320 24699 10360 24731
rect 10392 24699 10432 24731
rect 10464 24699 10504 24731
rect 10536 24699 10576 24731
rect 10608 24699 10648 24731
rect 10680 24699 10720 24731
rect 10752 24699 10792 24731
rect 10824 24699 10864 24731
rect 10896 24699 10936 24731
rect 10968 24699 11008 24731
rect 11040 24699 11080 24731
rect 11112 24699 11152 24731
rect 11184 24699 11224 24731
rect 11256 24699 11296 24731
rect 11328 24699 11368 24731
rect 11400 24699 11440 24731
rect 11472 24699 11512 24731
rect 11544 24699 11584 24731
rect 11616 24699 11656 24731
rect 11688 24699 11728 24731
rect 11760 24699 11800 24731
rect 11832 24699 11872 24731
rect 11904 24699 11944 24731
rect 11976 24699 12016 24731
rect 12048 24699 12088 24731
rect 12120 24699 12160 24731
rect 12192 24699 12232 24731
rect 12264 24699 12304 24731
rect 12336 24699 12376 24731
rect 12408 24699 12448 24731
rect 12480 24699 12520 24731
rect 12552 24699 12592 24731
rect 12624 24699 12664 24731
rect 12696 24699 12736 24731
rect 12768 24699 12808 24731
rect 12840 24699 12880 24731
rect 12912 24699 12952 24731
rect 12984 24699 13024 24731
rect 13056 24699 13096 24731
rect 13128 24699 13168 24731
rect 13200 24699 13240 24731
rect 13272 24699 13312 24731
rect 13344 24699 13384 24731
rect 13416 24699 13456 24731
rect 13488 24699 13528 24731
rect 13560 24699 13600 24731
rect 13632 24699 13672 24731
rect 13704 24699 13744 24731
rect 13776 24699 13816 24731
rect 13848 24699 13888 24731
rect 13920 24699 13960 24731
rect 13992 24699 14032 24731
rect 14064 24699 14104 24731
rect 14136 24699 14176 24731
rect 14208 24699 14248 24731
rect 14280 24699 14320 24731
rect 14352 24699 14392 24731
rect 14424 24699 14464 24731
rect 14496 24699 14536 24731
rect 14568 24699 14608 24731
rect 14640 24699 14680 24731
rect 14712 24699 14752 24731
rect 14784 24699 14824 24731
rect 14856 24699 14896 24731
rect 14928 24699 14968 24731
rect 15000 24699 15040 24731
rect 15072 24699 15112 24731
rect 15144 24699 15184 24731
rect 15216 24699 15256 24731
rect 15288 24699 15328 24731
rect 15360 24699 15400 24731
rect 15432 24699 15472 24731
rect 15504 24699 15544 24731
rect 15576 24699 15616 24731
rect 15648 24699 15688 24731
rect 15720 24699 15760 24731
rect 15792 24699 15832 24731
rect 15864 24699 15904 24731
rect 15936 24699 16000 24731
rect 0 24659 16000 24699
rect 0 24627 64 24659
rect 96 24627 136 24659
rect 168 24627 208 24659
rect 240 24627 280 24659
rect 312 24627 352 24659
rect 384 24627 424 24659
rect 456 24627 496 24659
rect 528 24627 568 24659
rect 600 24627 640 24659
rect 672 24627 712 24659
rect 744 24627 784 24659
rect 816 24627 856 24659
rect 888 24627 928 24659
rect 960 24627 1000 24659
rect 1032 24627 1072 24659
rect 1104 24627 1144 24659
rect 1176 24627 1216 24659
rect 1248 24627 1288 24659
rect 1320 24627 1360 24659
rect 1392 24627 1432 24659
rect 1464 24627 1504 24659
rect 1536 24627 1576 24659
rect 1608 24627 1648 24659
rect 1680 24627 1720 24659
rect 1752 24627 1792 24659
rect 1824 24627 1864 24659
rect 1896 24627 1936 24659
rect 1968 24627 2008 24659
rect 2040 24627 2080 24659
rect 2112 24627 2152 24659
rect 2184 24627 2224 24659
rect 2256 24627 2296 24659
rect 2328 24627 2368 24659
rect 2400 24627 2440 24659
rect 2472 24627 2512 24659
rect 2544 24627 2584 24659
rect 2616 24627 2656 24659
rect 2688 24627 2728 24659
rect 2760 24627 2800 24659
rect 2832 24627 2872 24659
rect 2904 24627 2944 24659
rect 2976 24627 3016 24659
rect 3048 24627 3088 24659
rect 3120 24627 3160 24659
rect 3192 24627 3232 24659
rect 3264 24627 3304 24659
rect 3336 24627 3376 24659
rect 3408 24627 3448 24659
rect 3480 24627 3520 24659
rect 3552 24627 3592 24659
rect 3624 24627 3664 24659
rect 3696 24627 3736 24659
rect 3768 24627 3808 24659
rect 3840 24627 3880 24659
rect 3912 24627 3952 24659
rect 3984 24627 4024 24659
rect 4056 24627 4096 24659
rect 4128 24627 4168 24659
rect 4200 24627 4240 24659
rect 4272 24627 4312 24659
rect 4344 24627 4384 24659
rect 4416 24627 4456 24659
rect 4488 24627 4528 24659
rect 4560 24627 4600 24659
rect 4632 24627 4672 24659
rect 4704 24627 4744 24659
rect 4776 24627 4816 24659
rect 4848 24627 4888 24659
rect 4920 24627 4960 24659
rect 4992 24627 5032 24659
rect 5064 24627 5104 24659
rect 5136 24627 5176 24659
rect 5208 24627 5248 24659
rect 5280 24627 5320 24659
rect 5352 24627 5392 24659
rect 5424 24627 5464 24659
rect 5496 24627 5536 24659
rect 5568 24627 5608 24659
rect 5640 24627 5680 24659
rect 5712 24627 5752 24659
rect 5784 24627 5824 24659
rect 5856 24627 5896 24659
rect 5928 24627 5968 24659
rect 6000 24627 6040 24659
rect 6072 24627 6112 24659
rect 6144 24627 6184 24659
rect 6216 24627 6256 24659
rect 6288 24627 6328 24659
rect 6360 24627 6400 24659
rect 6432 24627 6472 24659
rect 6504 24627 6544 24659
rect 6576 24627 6616 24659
rect 6648 24627 6688 24659
rect 6720 24627 6760 24659
rect 6792 24627 6832 24659
rect 6864 24627 6904 24659
rect 6936 24627 6976 24659
rect 7008 24627 7048 24659
rect 7080 24627 7120 24659
rect 7152 24627 7192 24659
rect 7224 24627 7264 24659
rect 7296 24627 7336 24659
rect 7368 24627 7408 24659
rect 7440 24627 7480 24659
rect 7512 24627 7552 24659
rect 7584 24627 7624 24659
rect 7656 24627 7696 24659
rect 7728 24627 7768 24659
rect 7800 24627 7840 24659
rect 7872 24627 7912 24659
rect 7944 24627 7984 24659
rect 8016 24627 8056 24659
rect 8088 24627 8128 24659
rect 8160 24627 8200 24659
rect 8232 24627 8272 24659
rect 8304 24627 8344 24659
rect 8376 24627 8416 24659
rect 8448 24627 8488 24659
rect 8520 24627 8560 24659
rect 8592 24627 8632 24659
rect 8664 24627 8704 24659
rect 8736 24627 8776 24659
rect 8808 24627 8848 24659
rect 8880 24627 8920 24659
rect 8952 24627 8992 24659
rect 9024 24627 9064 24659
rect 9096 24627 9136 24659
rect 9168 24627 9208 24659
rect 9240 24627 9280 24659
rect 9312 24627 9352 24659
rect 9384 24627 9424 24659
rect 9456 24627 9496 24659
rect 9528 24627 9568 24659
rect 9600 24627 9640 24659
rect 9672 24627 9712 24659
rect 9744 24627 9784 24659
rect 9816 24627 9856 24659
rect 9888 24627 9928 24659
rect 9960 24627 10000 24659
rect 10032 24627 10072 24659
rect 10104 24627 10144 24659
rect 10176 24627 10216 24659
rect 10248 24627 10288 24659
rect 10320 24627 10360 24659
rect 10392 24627 10432 24659
rect 10464 24627 10504 24659
rect 10536 24627 10576 24659
rect 10608 24627 10648 24659
rect 10680 24627 10720 24659
rect 10752 24627 10792 24659
rect 10824 24627 10864 24659
rect 10896 24627 10936 24659
rect 10968 24627 11008 24659
rect 11040 24627 11080 24659
rect 11112 24627 11152 24659
rect 11184 24627 11224 24659
rect 11256 24627 11296 24659
rect 11328 24627 11368 24659
rect 11400 24627 11440 24659
rect 11472 24627 11512 24659
rect 11544 24627 11584 24659
rect 11616 24627 11656 24659
rect 11688 24627 11728 24659
rect 11760 24627 11800 24659
rect 11832 24627 11872 24659
rect 11904 24627 11944 24659
rect 11976 24627 12016 24659
rect 12048 24627 12088 24659
rect 12120 24627 12160 24659
rect 12192 24627 12232 24659
rect 12264 24627 12304 24659
rect 12336 24627 12376 24659
rect 12408 24627 12448 24659
rect 12480 24627 12520 24659
rect 12552 24627 12592 24659
rect 12624 24627 12664 24659
rect 12696 24627 12736 24659
rect 12768 24627 12808 24659
rect 12840 24627 12880 24659
rect 12912 24627 12952 24659
rect 12984 24627 13024 24659
rect 13056 24627 13096 24659
rect 13128 24627 13168 24659
rect 13200 24627 13240 24659
rect 13272 24627 13312 24659
rect 13344 24627 13384 24659
rect 13416 24627 13456 24659
rect 13488 24627 13528 24659
rect 13560 24627 13600 24659
rect 13632 24627 13672 24659
rect 13704 24627 13744 24659
rect 13776 24627 13816 24659
rect 13848 24627 13888 24659
rect 13920 24627 13960 24659
rect 13992 24627 14032 24659
rect 14064 24627 14104 24659
rect 14136 24627 14176 24659
rect 14208 24627 14248 24659
rect 14280 24627 14320 24659
rect 14352 24627 14392 24659
rect 14424 24627 14464 24659
rect 14496 24627 14536 24659
rect 14568 24627 14608 24659
rect 14640 24627 14680 24659
rect 14712 24627 14752 24659
rect 14784 24627 14824 24659
rect 14856 24627 14896 24659
rect 14928 24627 14968 24659
rect 15000 24627 15040 24659
rect 15072 24627 15112 24659
rect 15144 24627 15184 24659
rect 15216 24627 15256 24659
rect 15288 24627 15328 24659
rect 15360 24627 15400 24659
rect 15432 24627 15472 24659
rect 15504 24627 15544 24659
rect 15576 24627 15616 24659
rect 15648 24627 15688 24659
rect 15720 24627 15760 24659
rect 15792 24627 15832 24659
rect 15864 24627 15904 24659
rect 15936 24627 16000 24659
rect 0 24587 16000 24627
rect 0 24555 64 24587
rect 96 24555 136 24587
rect 168 24555 208 24587
rect 240 24555 280 24587
rect 312 24555 352 24587
rect 384 24555 424 24587
rect 456 24555 496 24587
rect 528 24555 568 24587
rect 600 24555 640 24587
rect 672 24555 712 24587
rect 744 24555 784 24587
rect 816 24555 856 24587
rect 888 24555 928 24587
rect 960 24555 1000 24587
rect 1032 24555 1072 24587
rect 1104 24555 1144 24587
rect 1176 24555 1216 24587
rect 1248 24555 1288 24587
rect 1320 24555 1360 24587
rect 1392 24555 1432 24587
rect 1464 24555 1504 24587
rect 1536 24555 1576 24587
rect 1608 24555 1648 24587
rect 1680 24555 1720 24587
rect 1752 24555 1792 24587
rect 1824 24555 1864 24587
rect 1896 24555 1936 24587
rect 1968 24555 2008 24587
rect 2040 24555 2080 24587
rect 2112 24555 2152 24587
rect 2184 24555 2224 24587
rect 2256 24555 2296 24587
rect 2328 24555 2368 24587
rect 2400 24555 2440 24587
rect 2472 24555 2512 24587
rect 2544 24555 2584 24587
rect 2616 24555 2656 24587
rect 2688 24555 2728 24587
rect 2760 24555 2800 24587
rect 2832 24555 2872 24587
rect 2904 24555 2944 24587
rect 2976 24555 3016 24587
rect 3048 24555 3088 24587
rect 3120 24555 3160 24587
rect 3192 24555 3232 24587
rect 3264 24555 3304 24587
rect 3336 24555 3376 24587
rect 3408 24555 3448 24587
rect 3480 24555 3520 24587
rect 3552 24555 3592 24587
rect 3624 24555 3664 24587
rect 3696 24555 3736 24587
rect 3768 24555 3808 24587
rect 3840 24555 3880 24587
rect 3912 24555 3952 24587
rect 3984 24555 4024 24587
rect 4056 24555 4096 24587
rect 4128 24555 4168 24587
rect 4200 24555 4240 24587
rect 4272 24555 4312 24587
rect 4344 24555 4384 24587
rect 4416 24555 4456 24587
rect 4488 24555 4528 24587
rect 4560 24555 4600 24587
rect 4632 24555 4672 24587
rect 4704 24555 4744 24587
rect 4776 24555 4816 24587
rect 4848 24555 4888 24587
rect 4920 24555 4960 24587
rect 4992 24555 5032 24587
rect 5064 24555 5104 24587
rect 5136 24555 5176 24587
rect 5208 24555 5248 24587
rect 5280 24555 5320 24587
rect 5352 24555 5392 24587
rect 5424 24555 5464 24587
rect 5496 24555 5536 24587
rect 5568 24555 5608 24587
rect 5640 24555 5680 24587
rect 5712 24555 5752 24587
rect 5784 24555 5824 24587
rect 5856 24555 5896 24587
rect 5928 24555 5968 24587
rect 6000 24555 6040 24587
rect 6072 24555 6112 24587
rect 6144 24555 6184 24587
rect 6216 24555 6256 24587
rect 6288 24555 6328 24587
rect 6360 24555 6400 24587
rect 6432 24555 6472 24587
rect 6504 24555 6544 24587
rect 6576 24555 6616 24587
rect 6648 24555 6688 24587
rect 6720 24555 6760 24587
rect 6792 24555 6832 24587
rect 6864 24555 6904 24587
rect 6936 24555 6976 24587
rect 7008 24555 7048 24587
rect 7080 24555 7120 24587
rect 7152 24555 7192 24587
rect 7224 24555 7264 24587
rect 7296 24555 7336 24587
rect 7368 24555 7408 24587
rect 7440 24555 7480 24587
rect 7512 24555 7552 24587
rect 7584 24555 7624 24587
rect 7656 24555 7696 24587
rect 7728 24555 7768 24587
rect 7800 24555 7840 24587
rect 7872 24555 7912 24587
rect 7944 24555 7984 24587
rect 8016 24555 8056 24587
rect 8088 24555 8128 24587
rect 8160 24555 8200 24587
rect 8232 24555 8272 24587
rect 8304 24555 8344 24587
rect 8376 24555 8416 24587
rect 8448 24555 8488 24587
rect 8520 24555 8560 24587
rect 8592 24555 8632 24587
rect 8664 24555 8704 24587
rect 8736 24555 8776 24587
rect 8808 24555 8848 24587
rect 8880 24555 8920 24587
rect 8952 24555 8992 24587
rect 9024 24555 9064 24587
rect 9096 24555 9136 24587
rect 9168 24555 9208 24587
rect 9240 24555 9280 24587
rect 9312 24555 9352 24587
rect 9384 24555 9424 24587
rect 9456 24555 9496 24587
rect 9528 24555 9568 24587
rect 9600 24555 9640 24587
rect 9672 24555 9712 24587
rect 9744 24555 9784 24587
rect 9816 24555 9856 24587
rect 9888 24555 9928 24587
rect 9960 24555 10000 24587
rect 10032 24555 10072 24587
rect 10104 24555 10144 24587
rect 10176 24555 10216 24587
rect 10248 24555 10288 24587
rect 10320 24555 10360 24587
rect 10392 24555 10432 24587
rect 10464 24555 10504 24587
rect 10536 24555 10576 24587
rect 10608 24555 10648 24587
rect 10680 24555 10720 24587
rect 10752 24555 10792 24587
rect 10824 24555 10864 24587
rect 10896 24555 10936 24587
rect 10968 24555 11008 24587
rect 11040 24555 11080 24587
rect 11112 24555 11152 24587
rect 11184 24555 11224 24587
rect 11256 24555 11296 24587
rect 11328 24555 11368 24587
rect 11400 24555 11440 24587
rect 11472 24555 11512 24587
rect 11544 24555 11584 24587
rect 11616 24555 11656 24587
rect 11688 24555 11728 24587
rect 11760 24555 11800 24587
rect 11832 24555 11872 24587
rect 11904 24555 11944 24587
rect 11976 24555 12016 24587
rect 12048 24555 12088 24587
rect 12120 24555 12160 24587
rect 12192 24555 12232 24587
rect 12264 24555 12304 24587
rect 12336 24555 12376 24587
rect 12408 24555 12448 24587
rect 12480 24555 12520 24587
rect 12552 24555 12592 24587
rect 12624 24555 12664 24587
rect 12696 24555 12736 24587
rect 12768 24555 12808 24587
rect 12840 24555 12880 24587
rect 12912 24555 12952 24587
rect 12984 24555 13024 24587
rect 13056 24555 13096 24587
rect 13128 24555 13168 24587
rect 13200 24555 13240 24587
rect 13272 24555 13312 24587
rect 13344 24555 13384 24587
rect 13416 24555 13456 24587
rect 13488 24555 13528 24587
rect 13560 24555 13600 24587
rect 13632 24555 13672 24587
rect 13704 24555 13744 24587
rect 13776 24555 13816 24587
rect 13848 24555 13888 24587
rect 13920 24555 13960 24587
rect 13992 24555 14032 24587
rect 14064 24555 14104 24587
rect 14136 24555 14176 24587
rect 14208 24555 14248 24587
rect 14280 24555 14320 24587
rect 14352 24555 14392 24587
rect 14424 24555 14464 24587
rect 14496 24555 14536 24587
rect 14568 24555 14608 24587
rect 14640 24555 14680 24587
rect 14712 24555 14752 24587
rect 14784 24555 14824 24587
rect 14856 24555 14896 24587
rect 14928 24555 14968 24587
rect 15000 24555 15040 24587
rect 15072 24555 15112 24587
rect 15144 24555 15184 24587
rect 15216 24555 15256 24587
rect 15288 24555 15328 24587
rect 15360 24555 15400 24587
rect 15432 24555 15472 24587
rect 15504 24555 15544 24587
rect 15576 24555 15616 24587
rect 15648 24555 15688 24587
rect 15720 24555 15760 24587
rect 15792 24555 15832 24587
rect 15864 24555 15904 24587
rect 15936 24555 16000 24587
rect 0 24515 16000 24555
rect 0 24483 64 24515
rect 96 24483 136 24515
rect 168 24483 208 24515
rect 240 24483 280 24515
rect 312 24483 352 24515
rect 384 24483 424 24515
rect 456 24483 496 24515
rect 528 24483 568 24515
rect 600 24483 640 24515
rect 672 24483 712 24515
rect 744 24483 784 24515
rect 816 24483 856 24515
rect 888 24483 928 24515
rect 960 24483 1000 24515
rect 1032 24483 1072 24515
rect 1104 24483 1144 24515
rect 1176 24483 1216 24515
rect 1248 24483 1288 24515
rect 1320 24483 1360 24515
rect 1392 24483 1432 24515
rect 1464 24483 1504 24515
rect 1536 24483 1576 24515
rect 1608 24483 1648 24515
rect 1680 24483 1720 24515
rect 1752 24483 1792 24515
rect 1824 24483 1864 24515
rect 1896 24483 1936 24515
rect 1968 24483 2008 24515
rect 2040 24483 2080 24515
rect 2112 24483 2152 24515
rect 2184 24483 2224 24515
rect 2256 24483 2296 24515
rect 2328 24483 2368 24515
rect 2400 24483 2440 24515
rect 2472 24483 2512 24515
rect 2544 24483 2584 24515
rect 2616 24483 2656 24515
rect 2688 24483 2728 24515
rect 2760 24483 2800 24515
rect 2832 24483 2872 24515
rect 2904 24483 2944 24515
rect 2976 24483 3016 24515
rect 3048 24483 3088 24515
rect 3120 24483 3160 24515
rect 3192 24483 3232 24515
rect 3264 24483 3304 24515
rect 3336 24483 3376 24515
rect 3408 24483 3448 24515
rect 3480 24483 3520 24515
rect 3552 24483 3592 24515
rect 3624 24483 3664 24515
rect 3696 24483 3736 24515
rect 3768 24483 3808 24515
rect 3840 24483 3880 24515
rect 3912 24483 3952 24515
rect 3984 24483 4024 24515
rect 4056 24483 4096 24515
rect 4128 24483 4168 24515
rect 4200 24483 4240 24515
rect 4272 24483 4312 24515
rect 4344 24483 4384 24515
rect 4416 24483 4456 24515
rect 4488 24483 4528 24515
rect 4560 24483 4600 24515
rect 4632 24483 4672 24515
rect 4704 24483 4744 24515
rect 4776 24483 4816 24515
rect 4848 24483 4888 24515
rect 4920 24483 4960 24515
rect 4992 24483 5032 24515
rect 5064 24483 5104 24515
rect 5136 24483 5176 24515
rect 5208 24483 5248 24515
rect 5280 24483 5320 24515
rect 5352 24483 5392 24515
rect 5424 24483 5464 24515
rect 5496 24483 5536 24515
rect 5568 24483 5608 24515
rect 5640 24483 5680 24515
rect 5712 24483 5752 24515
rect 5784 24483 5824 24515
rect 5856 24483 5896 24515
rect 5928 24483 5968 24515
rect 6000 24483 6040 24515
rect 6072 24483 6112 24515
rect 6144 24483 6184 24515
rect 6216 24483 6256 24515
rect 6288 24483 6328 24515
rect 6360 24483 6400 24515
rect 6432 24483 6472 24515
rect 6504 24483 6544 24515
rect 6576 24483 6616 24515
rect 6648 24483 6688 24515
rect 6720 24483 6760 24515
rect 6792 24483 6832 24515
rect 6864 24483 6904 24515
rect 6936 24483 6976 24515
rect 7008 24483 7048 24515
rect 7080 24483 7120 24515
rect 7152 24483 7192 24515
rect 7224 24483 7264 24515
rect 7296 24483 7336 24515
rect 7368 24483 7408 24515
rect 7440 24483 7480 24515
rect 7512 24483 7552 24515
rect 7584 24483 7624 24515
rect 7656 24483 7696 24515
rect 7728 24483 7768 24515
rect 7800 24483 7840 24515
rect 7872 24483 7912 24515
rect 7944 24483 7984 24515
rect 8016 24483 8056 24515
rect 8088 24483 8128 24515
rect 8160 24483 8200 24515
rect 8232 24483 8272 24515
rect 8304 24483 8344 24515
rect 8376 24483 8416 24515
rect 8448 24483 8488 24515
rect 8520 24483 8560 24515
rect 8592 24483 8632 24515
rect 8664 24483 8704 24515
rect 8736 24483 8776 24515
rect 8808 24483 8848 24515
rect 8880 24483 8920 24515
rect 8952 24483 8992 24515
rect 9024 24483 9064 24515
rect 9096 24483 9136 24515
rect 9168 24483 9208 24515
rect 9240 24483 9280 24515
rect 9312 24483 9352 24515
rect 9384 24483 9424 24515
rect 9456 24483 9496 24515
rect 9528 24483 9568 24515
rect 9600 24483 9640 24515
rect 9672 24483 9712 24515
rect 9744 24483 9784 24515
rect 9816 24483 9856 24515
rect 9888 24483 9928 24515
rect 9960 24483 10000 24515
rect 10032 24483 10072 24515
rect 10104 24483 10144 24515
rect 10176 24483 10216 24515
rect 10248 24483 10288 24515
rect 10320 24483 10360 24515
rect 10392 24483 10432 24515
rect 10464 24483 10504 24515
rect 10536 24483 10576 24515
rect 10608 24483 10648 24515
rect 10680 24483 10720 24515
rect 10752 24483 10792 24515
rect 10824 24483 10864 24515
rect 10896 24483 10936 24515
rect 10968 24483 11008 24515
rect 11040 24483 11080 24515
rect 11112 24483 11152 24515
rect 11184 24483 11224 24515
rect 11256 24483 11296 24515
rect 11328 24483 11368 24515
rect 11400 24483 11440 24515
rect 11472 24483 11512 24515
rect 11544 24483 11584 24515
rect 11616 24483 11656 24515
rect 11688 24483 11728 24515
rect 11760 24483 11800 24515
rect 11832 24483 11872 24515
rect 11904 24483 11944 24515
rect 11976 24483 12016 24515
rect 12048 24483 12088 24515
rect 12120 24483 12160 24515
rect 12192 24483 12232 24515
rect 12264 24483 12304 24515
rect 12336 24483 12376 24515
rect 12408 24483 12448 24515
rect 12480 24483 12520 24515
rect 12552 24483 12592 24515
rect 12624 24483 12664 24515
rect 12696 24483 12736 24515
rect 12768 24483 12808 24515
rect 12840 24483 12880 24515
rect 12912 24483 12952 24515
rect 12984 24483 13024 24515
rect 13056 24483 13096 24515
rect 13128 24483 13168 24515
rect 13200 24483 13240 24515
rect 13272 24483 13312 24515
rect 13344 24483 13384 24515
rect 13416 24483 13456 24515
rect 13488 24483 13528 24515
rect 13560 24483 13600 24515
rect 13632 24483 13672 24515
rect 13704 24483 13744 24515
rect 13776 24483 13816 24515
rect 13848 24483 13888 24515
rect 13920 24483 13960 24515
rect 13992 24483 14032 24515
rect 14064 24483 14104 24515
rect 14136 24483 14176 24515
rect 14208 24483 14248 24515
rect 14280 24483 14320 24515
rect 14352 24483 14392 24515
rect 14424 24483 14464 24515
rect 14496 24483 14536 24515
rect 14568 24483 14608 24515
rect 14640 24483 14680 24515
rect 14712 24483 14752 24515
rect 14784 24483 14824 24515
rect 14856 24483 14896 24515
rect 14928 24483 14968 24515
rect 15000 24483 15040 24515
rect 15072 24483 15112 24515
rect 15144 24483 15184 24515
rect 15216 24483 15256 24515
rect 15288 24483 15328 24515
rect 15360 24483 15400 24515
rect 15432 24483 15472 24515
rect 15504 24483 15544 24515
rect 15576 24483 15616 24515
rect 15648 24483 15688 24515
rect 15720 24483 15760 24515
rect 15792 24483 15832 24515
rect 15864 24483 15904 24515
rect 15936 24483 16000 24515
rect 0 24443 16000 24483
rect 0 24411 64 24443
rect 96 24411 136 24443
rect 168 24411 208 24443
rect 240 24411 280 24443
rect 312 24411 352 24443
rect 384 24411 424 24443
rect 456 24411 496 24443
rect 528 24411 568 24443
rect 600 24411 640 24443
rect 672 24411 712 24443
rect 744 24411 784 24443
rect 816 24411 856 24443
rect 888 24411 928 24443
rect 960 24411 1000 24443
rect 1032 24411 1072 24443
rect 1104 24411 1144 24443
rect 1176 24411 1216 24443
rect 1248 24411 1288 24443
rect 1320 24411 1360 24443
rect 1392 24411 1432 24443
rect 1464 24411 1504 24443
rect 1536 24411 1576 24443
rect 1608 24411 1648 24443
rect 1680 24411 1720 24443
rect 1752 24411 1792 24443
rect 1824 24411 1864 24443
rect 1896 24411 1936 24443
rect 1968 24411 2008 24443
rect 2040 24411 2080 24443
rect 2112 24411 2152 24443
rect 2184 24411 2224 24443
rect 2256 24411 2296 24443
rect 2328 24411 2368 24443
rect 2400 24411 2440 24443
rect 2472 24411 2512 24443
rect 2544 24411 2584 24443
rect 2616 24411 2656 24443
rect 2688 24411 2728 24443
rect 2760 24411 2800 24443
rect 2832 24411 2872 24443
rect 2904 24411 2944 24443
rect 2976 24411 3016 24443
rect 3048 24411 3088 24443
rect 3120 24411 3160 24443
rect 3192 24411 3232 24443
rect 3264 24411 3304 24443
rect 3336 24411 3376 24443
rect 3408 24411 3448 24443
rect 3480 24411 3520 24443
rect 3552 24411 3592 24443
rect 3624 24411 3664 24443
rect 3696 24411 3736 24443
rect 3768 24411 3808 24443
rect 3840 24411 3880 24443
rect 3912 24411 3952 24443
rect 3984 24411 4024 24443
rect 4056 24411 4096 24443
rect 4128 24411 4168 24443
rect 4200 24411 4240 24443
rect 4272 24411 4312 24443
rect 4344 24411 4384 24443
rect 4416 24411 4456 24443
rect 4488 24411 4528 24443
rect 4560 24411 4600 24443
rect 4632 24411 4672 24443
rect 4704 24411 4744 24443
rect 4776 24411 4816 24443
rect 4848 24411 4888 24443
rect 4920 24411 4960 24443
rect 4992 24411 5032 24443
rect 5064 24411 5104 24443
rect 5136 24411 5176 24443
rect 5208 24411 5248 24443
rect 5280 24411 5320 24443
rect 5352 24411 5392 24443
rect 5424 24411 5464 24443
rect 5496 24411 5536 24443
rect 5568 24411 5608 24443
rect 5640 24411 5680 24443
rect 5712 24411 5752 24443
rect 5784 24411 5824 24443
rect 5856 24411 5896 24443
rect 5928 24411 5968 24443
rect 6000 24411 6040 24443
rect 6072 24411 6112 24443
rect 6144 24411 6184 24443
rect 6216 24411 6256 24443
rect 6288 24411 6328 24443
rect 6360 24411 6400 24443
rect 6432 24411 6472 24443
rect 6504 24411 6544 24443
rect 6576 24411 6616 24443
rect 6648 24411 6688 24443
rect 6720 24411 6760 24443
rect 6792 24411 6832 24443
rect 6864 24411 6904 24443
rect 6936 24411 6976 24443
rect 7008 24411 7048 24443
rect 7080 24411 7120 24443
rect 7152 24411 7192 24443
rect 7224 24411 7264 24443
rect 7296 24411 7336 24443
rect 7368 24411 7408 24443
rect 7440 24411 7480 24443
rect 7512 24411 7552 24443
rect 7584 24411 7624 24443
rect 7656 24411 7696 24443
rect 7728 24411 7768 24443
rect 7800 24411 7840 24443
rect 7872 24411 7912 24443
rect 7944 24411 7984 24443
rect 8016 24411 8056 24443
rect 8088 24411 8128 24443
rect 8160 24411 8200 24443
rect 8232 24411 8272 24443
rect 8304 24411 8344 24443
rect 8376 24411 8416 24443
rect 8448 24411 8488 24443
rect 8520 24411 8560 24443
rect 8592 24411 8632 24443
rect 8664 24411 8704 24443
rect 8736 24411 8776 24443
rect 8808 24411 8848 24443
rect 8880 24411 8920 24443
rect 8952 24411 8992 24443
rect 9024 24411 9064 24443
rect 9096 24411 9136 24443
rect 9168 24411 9208 24443
rect 9240 24411 9280 24443
rect 9312 24411 9352 24443
rect 9384 24411 9424 24443
rect 9456 24411 9496 24443
rect 9528 24411 9568 24443
rect 9600 24411 9640 24443
rect 9672 24411 9712 24443
rect 9744 24411 9784 24443
rect 9816 24411 9856 24443
rect 9888 24411 9928 24443
rect 9960 24411 10000 24443
rect 10032 24411 10072 24443
rect 10104 24411 10144 24443
rect 10176 24411 10216 24443
rect 10248 24411 10288 24443
rect 10320 24411 10360 24443
rect 10392 24411 10432 24443
rect 10464 24411 10504 24443
rect 10536 24411 10576 24443
rect 10608 24411 10648 24443
rect 10680 24411 10720 24443
rect 10752 24411 10792 24443
rect 10824 24411 10864 24443
rect 10896 24411 10936 24443
rect 10968 24411 11008 24443
rect 11040 24411 11080 24443
rect 11112 24411 11152 24443
rect 11184 24411 11224 24443
rect 11256 24411 11296 24443
rect 11328 24411 11368 24443
rect 11400 24411 11440 24443
rect 11472 24411 11512 24443
rect 11544 24411 11584 24443
rect 11616 24411 11656 24443
rect 11688 24411 11728 24443
rect 11760 24411 11800 24443
rect 11832 24411 11872 24443
rect 11904 24411 11944 24443
rect 11976 24411 12016 24443
rect 12048 24411 12088 24443
rect 12120 24411 12160 24443
rect 12192 24411 12232 24443
rect 12264 24411 12304 24443
rect 12336 24411 12376 24443
rect 12408 24411 12448 24443
rect 12480 24411 12520 24443
rect 12552 24411 12592 24443
rect 12624 24411 12664 24443
rect 12696 24411 12736 24443
rect 12768 24411 12808 24443
rect 12840 24411 12880 24443
rect 12912 24411 12952 24443
rect 12984 24411 13024 24443
rect 13056 24411 13096 24443
rect 13128 24411 13168 24443
rect 13200 24411 13240 24443
rect 13272 24411 13312 24443
rect 13344 24411 13384 24443
rect 13416 24411 13456 24443
rect 13488 24411 13528 24443
rect 13560 24411 13600 24443
rect 13632 24411 13672 24443
rect 13704 24411 13744 24443
rect 13776 24411 13816 24443
rect 13848 24411 13888 24443
rect 13920 24411 13960 24443
rect 13992 24411 14032 24443
rect 14064 24411 14104 24443
rect 14136 24411 14176 24443
rect 14208 24411 14248 24443
rect 14280 24411 14320 24443
rect 14352 24411 14392 24443
rect 14424 24411 14464 24443
rect 14496 24411 14536 24443
rect 14568 24411 14608 24443
rect 14640 24411 14680 24443
rect 14712 24411 14752 24443
rect 14784 24411 14824 24443
rect 14856 24411 14896 24443
rect 14928 24411 14968 24443
rect 15000 24411 15040 24443
rect 15072 24411 15112 24443
rect 15144 24411 15184 24443
rect 15216 24411 15256 24443
rect 15288 24411 15328 24443
rect 15360 24411 15400 24443
rect 15432 24411 15472 24443
rect 15504 24411 15544 24443
rect 15576 24411 15616 24443
rect 15648 24411 15688 24443
rect 15720 24411 15760 24443
rect 15792 24411 15832 24443
rect 15864 24411 15904 24443
rect 15936 24411 16000 24443
rect 0 24371 16000 24411
rect 0 24339 64 24371
rect 96 24339 136 24371
rect 168 24339 208 24371
rect 240 24339 280 24371
rect 312 24339 352 24371
rect 384 24339 424 24371
rect 456 24339 496 24371
rect 528 24339 568 24371
rect 600 24339 640 24371
rect 672 24339 712 24371
rect 744 24339 784 24371
rect 816 24339 856 24371
rect 888 24339 928 24371
rect 960 24339 1000 24371
rect 1032 24339 1072 24371
rect 1104 24339 1144 24371
rect 1176 24339 1216 24371
rect 1248 24339 1288 24371
rect 1320 24339 1360 24371
rect 1392 24339 1432 24371
rect 1464 24339 1504 24371
rect 1536 24339 1576 24371
rect 1608 24339 1648 24371
rect 1680 24339 1720 24371
rect 1752 24339 1792 24371
rect 1824 24339 1864 24371
rect 1896 24339 1936 24371
rect 1968 24339 2008 24371
rect 2040 24339 2080 24371
rect 2112 24339 2152 24371
rect 2184 24339 2224 24371
rect 2256 24339 2296 24371
rect 2328 24339 2368 24371
rect 2400 24339 2440 24371
rect 2472 24339 2512 24371
rect 2544 24339 2584 24371
rect 2616 24339 2656 24371
rect 2688 24339 2728 24371
rect 2760 24339 2800 24371
rect 2832 24339 2872 24371
rect 2904 24339 2944 24371
rect 2976 24339 3016 24371
rect 3048 24339 3088 24371
rect 3120 24339 3160 24371
rect 3192 24339 3232 24371
rect 3264 24339 3304 24371
rect 3336 24339 3376 24371
rect 3408 24339 3448 24371
rect 3480 24339 3520 24371
rect 3552 24339 3592 24371
rect 3624 24339 3664 24371
rect 3696 24339 3736 24371
rect 3768 24339 3808 24371
rect 3840 24339 3880 24371
rect 3912 24339 3952 24371
rect 3984 24339 4024 24371
rect 4056 24339 4096 24371
rect 4128 24339 4168 24371
rect 4200 24339 4240 24371
rect 4272 24339 4312 24371
rect 4344 24339 4384 24371
rect 4416 24339 4456 24371
rect 4488 24339 4528 24371
rect 4560 24339 4600 24371
rect 4632 24339 4672 24371
rect 4704 24339 4744 24371
rect 4776 24339 4816 24371
rect 4848 24339 4888 24371
rect 4920 24339 4960 24371
rect 4992 24339 5032 24371
rect 5064 24339 5104 24371
rect 5136 24339 5176 24371
rect 5208 24339 5248 24371
rect 5280 24339 5320 24371
rect 5352 24339 5392 24371
rect 5424 24339 5464 24371
rect 5496 24339 5536 24371
rect 5568 24339 5608 24371
rect 5640 24339 5680 24371
rect 5712 24339 5752 24371
rect 5784 24339 5824 24371
rect 5856 24339 5896 24371
rect 5928 24339 5968 24371
rect 6000 24339 6040 24371
rect 6072 24339 6112 24371
rect 6144 24339 6184 24371
rect 6216 24339 6256 24371
rect 6288 24339 6328 24371
rect 6360 24339 6400 24371
rect 6432 24339 6472 24371
rect 6504 24339 6544 24371
rect 6576 24339 6616 24371
rect 6648 24339 6688 24371
rect 6720 24339 6760 24371
rect 6792 24339 6832 24371
rect 6864 24339 6904 24371
rect 6936 24339 6976 24371
rect 7008 24339 7048 24371
rect 7080 24339 7120 24371
rect 7152 24339 7192 24371
rect 7224 24339 7264 24371
rect 7296 24339 7336 24371
rect 7368 24339 7408 24371
rect 7440 24339 7480 24371
rect 7512 24339 7552 24371
rect 7584 24339 7624 24371
rect 7656 24339 7696 24371
rect 7728 24339 7768 24371
rect 7800 24339 7840 24371
rect 7872 24339 7912 24371
rect 7944 24339 7984 24371
rect 8016 24339 8056 24371
rect 8088 24339 8128 24371
rect 8160 24339 8200 24371
rect 8232 24339 8272 24371
rect 8304 24339 8344 24371
rect 8376 24339 8416 24371
rect 8448 24339 8488 24371
rect 8520 24339 8560 24371
rect 8592 24339 8632 24371
rect 8664 24339 8704 24371
rect 8736 24339 8776 24371
rect 8808 24339 8848 24371
rect 8880 24339 8920 24371
rect 8952 24339 8992 24371
rect 9024 24339 9064 24371
rect 9096 24339 9136 24371
rect 9168 24339 9208 24371
rect 9240 24339 9280 24371
rect 9312 24339 9352 24371
rect 9384 24339 9424 24371
rect 9456 24339 9496 24371
rect 9528 24339 9568 24371
rect 9600 24339 9640 24371
rect 9672 24339 9712 24371
rect 9744 24339 9784 24371
rect 9816 24339 9856 24371
rect 9888 24339 9928 24371
rect 9960 24339 10000 24371
rect 10032 24339 10072 24371
rect 10104 24339 10144 24371
rect 10176 24339 10216 24371
rect 10248 24339 10288 24371
rect 10320 24339 10360 24371
rect 10392 24339 10432 24371
rect 10464 24339 10504 24371
rect 10536 24339 10576 24371
rect 10608 24339 10648 24371
rect 10680 24339 10720 24371
rect 10752 24339 10792 24371
rect 10824 24339 10864 24371
rect 10896 24339 10936 24371
rect 10968 24339 11008 24371
rect 11040 24339 11080 24371
rect 11112 24339 11152 24371
rect 11184 24339 11224 24371
rect 11256 24339 11296 24371
rect 11328 24339 11368 24371
rect 11400 24339 11440 24371
rect 11472 24339 11512 24371
rect 11544 24339 11584 24371
rect 11616 24339 11656 24371
rect 11688 24339 11728 24371
rect 11760 24339 11800 24371
rect 11832 24339 11872 24371
rect 11904 24339 11944 24371
rect 11976 24339 12016 24371
rect 12048 24339 12088 24371
rect 12120 24339 12160 24371
rect 12192 24339 12232 24371
rect 12264 24339 12304 24371
rect 12336 24339 12376 24371
rect 12408 24339 12448 24371
rect 12480 24339 12520 24371
rect 12552 24339 12592 24371
rect 12624 24339 12664 24371
rect 12696 24339 12736 24371
rect 12768 24339 12808 24371
rect 12840 24339 12880 24371
rect 12912 24339 12952 24371
rect 12984 24339 13024 24371
rect 13056 24339 13096 24371
rect 13128 24339 13168 24371
rect 13200 24339 13240 24371
rect 13272 24339 13312 24371
rect 13344 24339 13384 24371
rect 13416 24339 13456 24371
rect 13488 24339 13528 24371
rect 13560 24339 13600 24371
rect 13632 24339 13672 24371
rect 13704 24339 13744 24371
rect 13776 24339 13816 24371
rect 13848 24339 13888 24371
rect 13920 24339 13960 24371
rect 13992 24339 14032 24371
rect 14064 24339 14104 24371
rect 14136 24339 14176 24371
rect 14208 24339 14248 24371
rect 14280 24339 14320 24371
rect 14352 24339 14392 24371
rect 14424 24339 14464 24371
rect 14496 24339 14536 24371
rect 14568 24339 14608 24371
rect 14640 24339 14680 24371
rect 14712 24339 14752 24371
rect 14784 24339 14824 24371
rect 14856 24339 14896 24371
rect 14928 24339 14968 24371
rect 15000 24339 15040 24371
rect 15072 24339 15112 24371
rect 15144 24339 15184 24371
rect 15216 24339 15256 24371
rect 15288 24339 15328 24371
rect 15360 24339 15400 24371
rect 15432 24339 15472 24371
rect 15504 24339 15544 24371
rect 15576 24339 15616 24371
rect 15648 24339 15688 24371
rect 15720 24339 15760 24371
rect 15792 24339 15832 24371
rect 15864 24339 15904 24371
rect 15936 24339 16000 24371
rect 0 24299 16000 24339
rect 0 24267 64 24299
rect 96 24267 136 24299
rect 168 24267 208 24299
rect 240 24267 280 24299
rect 312 24267 352 24299
rect 384 24267 424 24299
rect 456 24267 496 24299
rect 528 24267 568 24299
rect 600 24267 640 24299
rect 672 24267 712 24299
rect 744 24267 784 24299
rect 816 24267 856 24299
rect 888 24267 928 24299
rect 960 24267 1000 24299
rect 1032 24267 1072 24299
rect 1104 24267 1144 24299
rect 1176 24267 1216 24299
rect 1248 24267 1288 24299
rect 1320 24267 1360 24299
rect 1392 24267 1432 24299
rect 1464 24267 1504 24299
rect 1536 24267 1576 24299
rect 1608 24267 1648 24299
rect 1680 24267 1720 24299
rect 1752 24267 1792 24299
rect 1824 24267 1864 24299
rect 1896 24267 1936 24299
rect 1968 24267 2008 24299
rect 2040 24267 2080 24299
rect 2112 24267 2152 24299
rect 2184 24267 2224 24299
rect 2256 24267 2296 24299
rect 2328 24267 2368 24299
rect 2400 24267 2440 24299
rect 2472 24267 2512 24299
rect 2544 24267 2584 24299
rect 2616 24267 2656 24299
rect 2688 24267 2728 24299
rect 2760 24267 2800 24299
rect 2832 24267 2872 24299
rect 2904 24267 2944 24299
rect 2976 24267 3016 24299
rect 3048 24267 3088 24299
rect 3120 24267 3160 24299
rect 3192 24267 3232 24299
rect 3264 24267 3304 24299
rect 3336 24267 3376 24299
rect 3408 24267 3448 24299
rect 3480 24267 3520 24299
rect 3552 24267 3592 24299
rect 3624 24267 3664 24299
rect 3696 24267 3736 24299
rect 3768 24267 3808 24299
rect 3840 24267 3880 24299
rect 3912 24267 3952 24299
rect 3984 24267 4024 24299
rect 4056 24267 4096 24299
rect 4128 24267 4168 24299
rect 4200 24267 4240 24299
rect 4272 24267 4312 24299
rect 4344 24267 4384 24299
rect 4416 24267 4456 24299
rect 4488 24267 4528 24299
rect 4560 24267 4600 24299
rect 4632 24267 4672 24299
rect 4704 24267 4744 24299
rect 4776 24267 4816 24299
rect 4848 24267 4888 24299
rect 4920 24267 4960 24299
rect 4992 24267 5032 24299
rect 5064 24267 5104 24299
rect 5136 24267 5176 24299
rect 5208 24267 5248 24299
rect 5280 24267 5320 24299
rect 5352 24267 5392 24299
rect 5424 24267 5464 24299
rect 5496 24267 5536 24299
rect 5568 24267 5608 24299
rect 5640 24267 5680 24299
rect 5712 24267 5752 24299
rect 5784 24267 5824 24299
rect 5856 24267 5896 24299
rect 5928 24267 5968 24299
rect 6000 24267 6040 24299
rect 6072 24267 6112 24299
rect 6144 24267 6184 24299
rect 6216 24267 6256 24299
rect 6288 24267 6328 24299
rect 6360 24267 6400 24299
rect 6432 24267 6472 24299
rect 6504 24267 6544 24299
rect 6576 24267 6616 24299
rect 6648 24267 6688 24299
rect 6720 24267 6760 24299
rect 6792 24267 6832 24299
rect 6864 24267 6904 24299
rect 6936 24267 6976 24299
rect 7008 24267 7048 24299
rect 7080 24267 7120 24299
rect 7152 24267 7192 24299
rect 7224 24267 7264 24299
rect 7296 24267 7336 24299
rect 7368 24267 7408 24299
rect 7440 24267 7480 24299
rect 7512 24267 7552 24299
rect 7584 24267 7624 24299
rect 7656 24267 7696 24299
rect 7728 24267 7768 24299
rect 7800 24267 7840 24299
rect 7872 24267 7912 24299
rect 7944 24267 7984 24299
rect 8016 24267 8056 24299
rect 8088 24267 8128 24299
rect 8160 24267 8200 24299
rect 8232 24267 8272 24299
rect 8304 24267 8344 24299
rect 8376 24267 8416 24299
rect 8448 24267 8488 24299
rect 8520 24267 8560 24299
rect 8592 24267 8632 24299
rect 8664 24267 8704 24299
rect 8736 24267 8776 24299
rect 8808 24267 8848 24299
rect 8880 24267 8920 24299
rect 8952 24267 8992 24299
rect 9024 24267 9064 24299
rect 9096 24267 9136 24299
rect 9168 24267 9208 24299
rect 9240 24267 9280 24299
rect 9312 24267 9352 24299
rect 9384 24267 9424 24299
rect 9456 24267 9496 24299
rect 9528 24267 9568 24299
rect 9600 24267 9640 24299
rect 9672 24267 9712 24299
rect 9744 24267 9784 24299
rect 9816 24267 9856 24299
rect 9888 24267 9928 24299
rect 9960 24267 10000 24299
rect 10032 24267 10072 24299
rect 10104 24267 10144 24299
rect 10176 24267 10216 24299
rect 10248 24267 10288 24299
rect 10320 24267 10360 24299
rect 10392 24267 10432 24299
rect 10464 24267 10504 24299
rect 10536 24267 10576 24299
rect 10608 24267 10648 24299
rect 10680 24267 10720 24299
rect 10752 24267 10792 24299
rect 10824 24267 10864 24299
rect 10896 24267 10936 24299
rect 10968 24267 11008 24299
rect 11040 24267 11080 24299
rect 11112 24267 11152 24299
rect 11184 24267 11224 24299
rect 11256 24267 11296 24299
rect 11328 24267 11368 24299
rect 11400 24267 11440 24299
rect 11472 24267 11512 24299
rect 11544 24267 11584 24299
rect 11616 24267 11656 24299
rect 11688 24267 11728 24299
rect 11760 24267 11800 24299
rect 11832 24267 11872 24299
rect 11904 24267 11944 24299
rect 11976 24267 12016 24299
rect 12048 24267 12088 24299
rect 12120 24267 12160 24299
rect 12192 24267 12232 24299
rect 12264 24267 12304 24299
rect 12336 24267 12376 24299
rect 12408 24267 12448 24299
rect 12480 24267 12520 24299
rect 12552 24267 12592 24299
rect 12624 24267 12664 24299
rect 12696 24267 12736 24299
rect 12768 24267 12808 24299
rect 12840 24267 12880 24299
rect 12912 24267 12952 24299
rect 12984 24267 13024 24299
rect 13056 24267 13096 24299
rect 13128 24267 13168 24299
rect 13200 24267 13240 24299
rect 13272 24267 13312 24299
rect 13344 24267 13384 24299
rect 13416 24267 13456 24299
rect 13488 24267 13528 24299
rect 13560 24267 13600 24299
rect 13632 24267 13672 24299
rect 13704 24267 13744 24299
rect 13776 24267 13816 24299
rect 13848 24267 13888 24299
rect 13920 24267 13960 24299
rect 13992 24267 14032 24299
rect 14064 24267 14104 24299
rect 14136 24267 14176 24299
rect 14208 24267 14248 24299
rect 14280 24267 14320 24299
rect 14352 24267 14392 24299
rect 14424 24267 14464 24299
rect 14496 24267 14536 24299
rect 14568 24267 14608 24299
rect 14640 24267 14680 24299
rect 14712 24267 14752 24299
rect 14784 24267 14824 24299
rect 14856 24267 14896 24299
rect 14928 24267 14968 24299
rect 15000 24267 15040 24299
rect 15072 24267 15112 24299
rect 15144 24267 15184 24299
rect 15216 24267 15256 24299
rect 15288 24267 15328 24299
rect 15360 24267 15400 24299
rect 15432 24267 15472 24299
rect 15504 24267 15544 24299
rect 15576 24267 15616 24299
rect 15648 24267 15688 24299
rect 15720 24267 15760 24299
rect 15792 24267 15832 24299
rect 15864 24267 15904 24299
rect 15936 24267 16000 24299
rect 0 24227 16000 24267
rect 0 24195 64 24227
rect 96 24195 136 24227
rect 168 24195 208 24227
rect 240 24195 280 24227
rect 312 24195 352 24227
rect 384 24195 424 24227
rect 456 24195 496 24227
rect 528 24195 568 24227
rect 600 24195 640 24227
rect 672 24195 712 24227
rect 744 24195 784 24227
rect 816 24195 856 24227
rect 888 24195 928 24227
rect 960 24195 1000 24227
rect 1032 24195 1072 24227
rect 1104 24195 1144 24227
rect 1176 24195 1216 24227
rect 1248 24195 1288 24227
rect 1320 24195 1360 24227
rect 1392 24195 1432 24227
rect 1464 24195 1504 24227
rect 1536 24195 1576 24227
rect 1608 24195 1648 24227
rect 1680 24195 1720 24227
rect 1752 24195 1792 24227
rect 1824 24195 1864 24227
rect 1896 24195 1936 24227
rect 1968 24195 2008 24227
rect 2040 24195 2080 24227
rect 2112 24195 2152 24227
rect 2184 24195 2224 24227
rect 2256 24195 2296 24227
rect 2328 24195 2368 24227
rect 2400 24195 2440 24227
rect 2472 24195 2512 24227
rect 2544 24195 2584 24227
rect 2616 24195 2656 24227
rect 2688 24195 2728 24227
rect 2760 24195 2800 24227
rect 2832 24195 2872 24227
rect 2904 24195 2944 24227
rect 2976 24195 3016 24227
rect 3048 24195 3088 24227
rect 3120 24195 3160 24227
rect 3192 24195 3232 24227
rect 3264 24195 3304 24227
rect 3336 24195 3376 24227
rect 3408 24195 3448 24227
rect 3480 24195 3520 24227
rect 3552 24195 3592 24227
rect 3624 24195 3664 24227
rect 3696 24195 3736 24227
rect 3768 24195 3808 24227
rect 3840 24195 3880 24227
rect 3912 24195 3952 24227
rect 3984 24195 4024 24227
rect 4056 24195 4096 24227
rect 4128 24195 4168 24227
rect 4200 24195 4240 24227
rect 4272 24195 4312 24227
rect 4344 24195 4384 24227
rect 4416 24195 4456 24227
rect 4488 24195 4528 24227
rect 4560 24195 4600 24227
rect 4632 24195 4672 24227
rect 4704 24195 4744 24227
rect 4776 24195 4816 24227
rect 4848 24195 4888 24227
rect 4920 24195 4960 24227
rect 4992 24195 5032 24227
rect 5064 24195 5104 24227
rect 5136 24195 5176 24227
rect 5208 24195 5248 24227
rect 5280 24195 5320 24227
rect 5352 24195 5392 24227
rect 5424 24195 5464 24227
rect 5496 24195 5536 24227
rect 5568 24195 5608 24227
rect 5640 24195 5680 24227
rect 5712 24195 5752 24227
rect 5784 24195 5824 24227
rect 5856 24195 5896 24227
rect 5928 24195 5968 24227
rect 6000 24195 6040 24227
rect 6072 24195 6112 24227
rect 6144 24195 6184 24227
rect 6216 24195 6256 24227
rect 6288 24195 6328 24227
rect 6360 24195 6400 24227
rect 6432 24195 6472 24227
rect 6504 24195 6544 24227
rect 6576 24195 6616 24227
rect 6648 24195 6688 24227
rect 6720 24195 6760 24227
rect 6792 24195 6832 24227
rect 6864 24195 6904 24227
rect 6936 24195 6976 24227
rect 7008 24195 7048 24227
rect 7080 24195 7120 24227
rect 7152 24195 7192 24227
rect 7224 24195 7264 24227
rect 7296 24195 7336 24227
rect 7368 24195 7408 24227
rect 7440 24195 7480 24227
rect 7512 24195 7552 24227
rect 7584 24195 7624 24227
rect 7656 24195 7696 24227
rect 7728 24195 7768 24227
rect 7800 24195 7840 24227
rect 7872 24195 7912 24227
rect 7944 24195 7984 24227
rect 8016 24195 8056 24227
rect 8088 24195 8128 24227
rect 8160 24195 8200 24227
rect 8232 24195 8272 24227
rect 8304 24195 8344 24227
rect 8376 24195 8416 24227
rect 8448 24195 8488 24227
rect 8520 24195 8560 24227
rect 8592 24195 8632 24227
rect 8664 24195 8704 24227
rect 8736 24195 8776 24227
rect 8808 24195 8848 24227
rect 8880 24195 8920 24227
rect 8952 24195 8992 24227
rect 9024 24195 9064 24227
rect 9096 24195 9136 24227
rect 9168 24195 9208 24227
rect 9240 24195 9280 24227
rect 9312 24195 9352 24227
rect 9384 24195 9424 24227
rect 9456 24195 9496 24227
rect 9528 24195 9568 24227
rect 9600 24195 9640 24227
rect 9672 24195 9712 24227
rect 9744 24195 9784 24227
rect 9816 24195 9856 24227
rect 9888 24195 9928 24227
rect 9960 24195 10000 24227
rect 10032 24195 10072 24227
rect 10104 24195 10144 24227
rect 10176 24195 10216 24227
rect 10248 24195 10288 24227
rect 10320 24195 10360 24227
rect 10392 24195 10432 24227
rect 10464 24195 10504 24227
rect 10536 24195 10576 24227
rect 10608 24195 10648 24227
rect 10680 24195 10720 24227
rect 10752 24195 10792 24227
rect 10824 24195 10864 24227
rect 10896 24195 10936 24227
rect 10968 24195 11008 24227
rect 11040 24195 11080 24227
rect 11112 24195 11152 24227
rect 11184 24195 11224 24227
rect 11256 24195 11296 24227
rect 11328 24195 11368 24227
rect 11400 24195 11440 24227
rect 11472 24195 11512 24227
rect 11544 24195 11584 24227
rect 11616 24195 11656 24227
rect 11688 24195 11728 24227
rect 11760 24195 11800 24227
rect 11832 24195 11872 24227
rect 11904 24195 11944 24227
rect 11976 24195 12016 24227
rect 12048 24195 12088 24227
rect 12120 24195 12160 24227
rect 12192 24195 12232 24227
rect 12264 24195 12304 24227
rect 12336 24195 12376 24227
rect 12408 24195 12448 24227
rect 12480 24195 12520 24227
rect 12552 24195 12592 24227
rect 12624 24195 12664 24227
rect 12696 24195 12736 24227
rect 12768 24195 12808 24227
rect 12840 24195 12880 24227
rect 12912 24195 12952 24227
rect 12984 24195 13024 24227
rect 13056 24195 13096 24227
rect 13128 24195 13168 24227
rect 13200 24195 13240 24227
rect 13272 24195 13312 24227
rect 13344 24195 13384 24227
rect 13416 24195 13456 24227
rect 13488 24195 13528 24227
rect 13560 24195 13600 24227
rect 13632 24195 13672 24227
rect 13704 24195 13744 24227
rect 13776 24195 13816 24227
rect 13848 24195 13888 24227
rect 13920 24195 13960 24227
rect 13992 24195 14032 24227
rect 14064 24195 14104 24227
rect 14136 24195 14176 24227
rect 14208 24195 14248 24227
rect 14280 24195 14320 24227
rect 14352 24195 14392 24227
rect 14424 24195 14464 24227
rect 14496 24195 14536 24227
rect 14568 24195 14608 24227
rect 14640 24195 14680 24227
rect 14712 24195 14752 24227
rect 14784 24195 14824 24227
rect 14856 24195 14896 24227
rect 14928 24195 14968 24227
rect 15000 24195 15040 24227
rect 15072 24195 15112 24227
rect 15144 24195 15184 24227
rect 15216 24195 15256 24227
rect 15288 24195 15328 24227
rect 15360 24195 15400 24227
rect 15432 24195 15472 24227
rect 15504 24195 15544 24227
rect 15576 24195 15616 24227
rect 15648 24195 15688 24227
rect 15720 24195 15760 24227
rect 15792 24195 15832 24227
rect 15864 24195 15904 24227
rect 15936 24195 16000 24227
rect 0 24155 16000 24195
rect 0 24123 64 24155
rect 96 24123 136 24155
rect 168 24123 208 24155
rect 240 24123 280 24155
rect 312 24123 352 24155
rect 384 24123 424 24155
rect 456 24123 496 24155
rect 528 24123 568 24155
rect 600 24123 640 24155
rect 672 24123 712 24155
rect 744 24123 784 24155
rect 816 24123 856 24155
rect 888 24123 928 24155
rect 960 24123 1000 24155
rect 1032 24123 1072 24155
rect 1104 24123 1144 24155
rect 1176 24123 1216 24155
rect 1248 24123 1288 24155
rect 1320 24123 1360 24155
rect 1392 24123 1432 24155
rect 1464 24123 1504 24155
rect 1536 24123 1576 24155
rect 1608 24123 1648 24155
rect 1680 24123 1720 24155
rect 1752 24123 1792 24155
rect 1824 24123 1864 24155
rect 1896 24123 1936 24155
rect 1968 24123 2008 24155
rect 2040 24123 2080 24155
rect 2112 24123 2152 24155
rect 2184 24123 2224 24155
rect 2256 24123 2296 24155
rect 2328 24123 2368 24155
rect 2400 24123 2440 24155
rect 2472 24123 2512 24155
rect 2544 24123 2584 24155
rect 2616 24123 2656 24155
rect 2688 24123 2728 24155
rect 2760 24123 2800 24155
rect 2832 24123 2872 24155
rect 2904 24123 2944 24155
rect 2976 24123 3016 24155
rect 3048 24123 3088 24155
rect 3120 24123 3160 24155
rect 3192 24123 3232 24155
rect 3264 24123 3304 24155
rect 3336 24123 3376 24155
rect 3408 24123 3448 24155
rect 3480 24123 3520 24155
rect 3552 24123 3592 24155
rect 3624 24123 3664 24155
rect 3696 24123 3736 24155
rect 3768 24123 3808 24155
rect 3840 24123 3880 24155
rect 3912 24123 3952 24155
rect 3984 24123 4024 24155
rect 4056 24123 4096 24155
rect 4128 24123 4168 24155
rect 4200 24123 4240 24155
rect 4272 24123 4312 24155
rect 4344 24123 4384 24155
rect 4416 24123 4456 24155
rect 4488 24123 4528 24155
rect 4560 24123 4600 24155
rect 4632 24123 4672 24155
rect 4704 24123 4744 24155
rect 4776 24123 4816 24155
rect 4848 24123 4888 24155
rect 4920 24123 4960 24155
rect 4992 24123 5032 24155
rect 5064 24123 5104 24155
rect 5136 24123 5176 24155
rect 5208 24123 5248 24155
rect 5280 24123 5320 24155
rect 5352 24123 5392 24155
rect 5424 24123 5464 24155
rect 5496 24123 5536 24155
rect 5568 24123 5608 24155
rect 5640 24123 5680 24155
rect 5712 24123 5752 24155
rect 5784 24123 5824 24155
rect 5856 24123 5896 24155
rect 5928 24123 5968 24155
rect 6000 24123 6040 24155
rect 6072 24123 6112 24155
rect 6144 24123 6184 24155
rect 6216 24123 6256 24155
rect 6288 24123 6328 24155
rect 6360 24123 6400 24155
rect 6432 24123 6472 24155
rect 6504 24123 6544 24155
rect 6576 24123 6616 24155
rect 6648 24123 6688 24155
rect 6720 24123 6760 24155
rect 6792 24123 6832 24155
rect 6864 24123 6904 24155
rect 6936 24123 6976 24155
rect 7008 24123 7048 24155
rect 7080 24123 7120 24155
rect 7152 24123 7192 24155
rect 7224 24123 7264 24155
rect 7296 24123 7336 24155
rect 7368 24123 7408 24155
rect 7440 24123 7480 24155
rect 7512 24123 7552 24155
rect 7584 24123 7624 24155
rect 7656 24123 7696 24155
rect 7728 24123 7768 24155
rect 7800 24123 7840 24155
rect 7872 24123 7912 24155
rect 7944 24123 7984 24155
rect 8016 24123 8056 24155
rect 8088 24123 8128 24155
rect 8160 24123 8200 24155
rect 8232 24123 8272 24155
rect 8304 24123 8344 24155
rect 8376 24123 8416 24155
rect 8448 24123 8488 24155
rect 8520 24123 8560 24155
rect 8592 24123 8632 24155
rect 8664 24123 8704 24155
rect 8736 24123 8776 24155
rect 8808 24123 8848 24155
rect 8880 24123 8920 24155
rect 8952 24123 8992 24155
rect 9024 24123 9064 24155
rect 9096 24123 9136 24155
rect 9168 24123 9208 24155
rect 9240 24123 9280 24155
rect 9312 24123 9352 24155
rect 9384 24123 9424 24155
rect 9456 24123 9496 24155
rect 9528 24123 9568 24155
rect 9600 24123 9640 24155
rect 9672 24123 9712 24155
rect 9744 24123 9784 24155
rect 9816 24123 9856 24155
rect 9888 24123 9928 24155
rect 9960 24123 10000 24155
rect 10032 24123 10072 24155
rect 10104 24123 10144 24155
rect 10176 24123 10216 24155
rect 10248 24123 10288 24155
rect 10320 24123 10360 24155
rect 10392 24123 10432 24155
rect 10464 24123 10504 24155
rect 10536 24123 10576 24155
rect 10608 24123 10648 24155
rect 10680 24123 10720 24155
rect 10752 24123 10792 24155
rect 10824 24123 10864 24155
rect 10896 24123 10936 24155
rect 10968 24123 11008 24155
rect 11040 24123 11080 24155
rect 11112 24123 11152 24155
rect 11184 24123 11224 24155
rect 11256 24123 11296 24155
rect 11328 24123 11368 24155
rect 11400 24123 11440 24155
rect 11472 24123 11512 24155
rect 11544 24123 11584 24155
rect 11616 24123 11656 24155
rect 11688 24123 11728 24155
rect 11760 24123 11800 24155
rect 11832 24123 11872 24155
rect 11904 24123 11944 24155
rect 11976 24123 12016 24155
rect 12048 24123 12088 24155
rect 12120 24123 12160 24155
rect 12192 24123 12232 24155
rect 12264 24123 12304 24155
rect 12336 24123 12376 24155
rect 12408 24123 12448 24155
rect 12480 24123 12520 24155
rect 12552 24123 12592 24155
rect 12624 24123 12664 24155
rect 12696 24123 12736 24155
rect 12768 24123 12808 24155
rect 12840 24123 12880 24155
rect 12912 24123 12952 24155
rect 12984 24123 13024 24155
rect 13056 24123 13096 24155
rect 13128 24123 13168 24155
rect 13200 24123 13240 24155
rect 13272 24123 13312 24155
rect 13344 24123 13384 24155
rect 13416 24123 13456 24155
rect 13488 24123 13528 24155
rect 13560 24123 13600 24155
rect 13632 24123 13672 24155
rect 13704 24123 13744 24155
rect 13776 24123 13816 24155
rect 13848 24123 13888 24155
rect 13920 24123 13960 24155
rect 13992 24123 14032 24155
rect 14064 24123 14104 24155
rect 14136 24123 14176 24155
rect 14208 24123 14248 24155
rect 14280 24123 14320 24155
rect 14352 24123 14392 24155
rect 14424 24123 14464 24155
rect 14496 24123 14536 24155
rect 14568 24123 14608 24155
rect 14640 24123 14680 24155
rect 14712 24123 14752 24155
rect 14784 24123 14824 24155
rect 14856 24123 14896 24155
rect 14928 24123 14968 24155
rect 15000 24123 15040 24155
rect 15072 24123 15112 24155
rect 15144 24123 15184 24155
rect 15216 24123 15256 24155
rect 15288 24123 15328 24155
rect 15360 24123 15400 24155
rect 15432 24123 15472 24155
rect 15504 24123 15544 24155
rect 15576 24123 15616 24155
rect 15648 24123 15688 24155
rect 15720 24123 15760 24155
rect 15792 24123 15832 24155
rect 15864 24123 15904 24155
rect 15936 24123 16000 24155
rect 0 24083 16000 24123
rect 0 24051 64 24083
rect 96 24051 136 24083
rect 168 24051 208 24083
rect 240 24051 280 24083
rect 312 24051 352 24083
rect 384 24051 424 24083
rect 456 24051 496 24083
rect 528 24051 568 24083
rect 600 24051 640 24083
rect 672 24051 712 24083
rect 744 24051 784 24083
rect 816 24051 856 24083
rect 888 24051 928 24083
rect 960 24051 1000 24083
rect 1032 24051 1072 24083
rect 1104 24051 1144 24083
rect 1176 24051 1216 24083
rect 1248 24051 1288 24083
rect 1320 24051 1360 24083
rect 1392 24051 1432 24083
rect 1464 24051 1504 24083
rect 1536 24051 1576 24083
rect 1608 24051 1648 24083
rect 1680 24051 1720 24083
rect 1752 24051 1792 24083
rect 1824 24051 1864 24083
rect 1896 24051 1936 24083
rect 1968 24051 2008 24083
rect 2040 24051 2080 24083
rect 2112 24051 2152 24083
rect 2184 24051 2224 24083
rect 2256 24051 2296 24083
rect 2328 24051 2368 24083
rect 2400 24051 2440 24083
rect 2472 24051 2512 24083
rect 2544 24051 2584 24083
rect 2616 24051 2656 24083
rect 2688 24051 2728 24083
rect 2760 24051 2800 24083
rect 2832 24051 2872 24083
rect 2904 24051 2944 24083
rect 2976 24051 3016 24083
rect 3048 24051 3088 24083
rect 3120 24051 3160 24083
rect 3192 24051 3232 24083
rect 3264 24051 3304 24083
rect 3336 24051 3376 24083
rect 3408 24051 3448 24083
rect 3480 24051 3520 24083
rect 3552 24051 3592 24083
rect 3624 24051 3664 24083
rect 3696 24051 3736 24083
rect 3768 24051 3808 24083
rect 3840 24051 3880 24083
rect 3912 24051 3952 24083
rect 3984 24051 4024 24083
rect 4056 24051 4096 24083
rect 4128 24051 4168 24083
rect 4200 24051 4240 24083
rect 4272 24051 4312 24083
rect 4344 24051 4384 24083
rect 4416 24051 4456 24083
rect 4488 24051 4528 24083
rect 4560 24051 4600 24083
rect 4632 24051 4672 24083
rect 4704 24051 4744 24083
rect 4776 24051 4816 24083
rect 4848 24051 4888 24083
rect 4920 24051 4960 24083
rect 4992 24051 5032 24083
rect 5064 24051 5104 24083
rect 5136 24051 5176 24083
rect 5208 24051 5248 24083
rect 5280 24051 5320 24083
rect 5352 24051 5392 24083
rect 5424 24051 5464 24083
rect 5496 24051 5536 24083
rect 5568 24051 5608 24083
rect 5640 24051 5680 24083
rect 5712 24051 5752 24083
rect 5784 24051 5824 24083
rect 5856 24051 5896 24083
rect 5928 24051 5968 24083
rect 6000 24051 6040 24083
rect 6072 24051 6112 24083
rect 6144 24051 6184 24083
rect 6216 24051 6256 24083
rect 6288 24051 6328 24083
rect 6360 24051 6400 24083
rect 6432 24051 6472 24083
rect 6504 24051 6544 24083
rect 6576 24051 6616 24083
rect 6648 24051 6688 24083
rect 6720 24051 6760 24083
rect 6792 24051 6832 24083
rect 6864 24051 6904 24083
rect 6936 24051 6976 24083
rect 7008 24051 7048 24083
rect 7080 24051 7120 24083
rect 7152 24051 7192 24083
rect 7224 24051 7264 24083
rect 7296 24051 7336 24083
rect 7368 24051 7408 24083
rect 7440 24051 7480 24083
rect 7512 24051 7552 24083
rect 7584 24051 7624 24083
rect 7656 24051 7696 24083
rect 7728 24051 7768 24083
rect 7800 24051 7840 24083
rect 7872 24051 7912 24083
rect 7944 24051 7984 24083
rect 8016 24051 8056 24083
rect 8088 24051 8128 24083
rect 8160 24051 8200 24083
rect 8232 24051 8272 24083
rect 8304 24051 8344 24083
rect 8376 24051 8416 24083
rect 8448 24051 8488 24083
rect 8520 24051 8560 24083
rect 8592 24051 8632 24083
rect 8664 24051 8704 24083
rect 8736 24051 8776 24083
rect 8808 24051 8848 24083
rect 8880 24051 8920 24083
rect 8952 24051 8992 24083
rect 9024 24051 9064 24083
rect 9096 24051 9136 24083
rect 9168 24051 9208 24083
rect 9240 24051 9280 24083
rect 9312 24051 9352 24083
rect 9384 24051 9424 24083
rect 9456 24051 9496 24083
rect 9528 24051 9568 24083
rect 9600 24051 9640 24083
rect 9672 24051 9712 24083
rect 9744 24051 9784 24083
rect 9816 24051 9856 24083
rect 9888 24051 9928 24083
rect 9960 24051 10000 24083
rect 10032 24051 10072 24083
rect 10104 24051 10144 24083
rect 10176 24051 10216 24083
rect 10248 24051 10288 24083
rect 10320 24051 10360 24083
rect 10392 24051 10432 24083
rect 10464 24051 10504 24083
rect 10536 24051 10576 24083
rect 10608 24051 10648 24083
rect 10680 24051 10720 24083
rect 10752 24051 10792 24083
rect 10824 24051 10864 24083
rect 10896 24051 10936 24083
rect 10968 24051 11008 24083
rect 11040 24051 11080 24083
rect 11112 24051 11152 24083
rect 11184 24051 11224 24083
rect 11256 24051 11296 24083
rect 11328 24051 11368 24083
rect 11400 24051 11440 24083
rect 11472 24051 11512 24083
rect 11544 24051 11584 24083
rect 11616 24051 11656 24083
rect 11688 24051 11728 24083
rect 11760 24051 11800 24083
rect 11832 24051 11872 24083
rect 11904 24051 11944 24083
rect 11976 24051 12016 24083
rect 12048 24051 12088 24083
rect 12120 24051 12160 24083
rect 12192 24051 12232 24083
rect 12264 24051 12304 24083
rect 12336 24051 12376 24083
rect 12408 24051 12448 24083
rect 12480 24051 12520 24083
rect 12552 24051 12592 24083
rect 12624 24051 12664 24083
rect 12696 24051 12736 24083
rect 12768 24051 12808 24083
rect 12840 24051 12880 24083
rect 12912 24051 12952 24083
rect 12984 24051 13024 24083
rect 13056 24051 13096 24083
rect 13128 24051 13168 24083
rect 13200 24051 13240 24083
rect 13272 24051 13312 24083
rect 13344 24051 13384 24083
rect 13416 24051 13456 24083
rect 13488 24051 13528 24083
rect 13560 24051 13600 24083
rect 13632 24051 13672 24083
rect 13704 24051 13744 24083
rect 13776 24051 13816 24083
rect 13848 24051 13888 24083
rect 13920 24051 13960 24083
rect 13992 24051 14032 24083
rect 14064 24051 14104 24083
rect 14136 24051 14176 24083
rect 14208 24051 14248 24083
rect 14280 24051 14320 24083
rect 14352 24051 14392 24083
rect 14424 24051 14464 24083
rect 14496 24051 14536 24083
rect 14568 24051 14608 24083
rect 14640 24051 14680 24083
rect 14712 24051 14752 24083
rect 14784 24051 14824 24083
rect 14856 24051 14896 24083
rect 14928 24051 14968 24083
rect 15000 24051 15040 24083
rect 15072 24051 15112 24083
rect 15144 24051 15184 24083
rect 15216 24051 15256 24083
rect 15288 24051 15328 24083
rect 15360 24051 15400 24083
rect 15432 24051 15472 24083
rect 15504 24051 15544 24083
rect 15576 24051 15616 24083
rect 15648 24051 15688 24083
rect 15720 24051 15760 24083
rect 15792 24051 15832 24083
rect 15864 24051 15904 24083
rect 15936 24051 16000 24083
rect 0 24011 16000 24051
rect 0 23979 64 24011
rect 96 23979 136 24011
rect 168 23979 208 24011
rect 240 23979 280 24011
rect 312 23979 352 24011
rect 384 23979 424 24011
rect 456 23979 496 24011
rect 528 23979 568 24011
rect 600 23979 640 24011
rect 672 23979 712 24011
rect 744 23979 784 24011
rect 816 23979 856 24011
rect 888 23979 928 24011
rect 960 23979 1000 24011
rect 1032 23979 1072 24011
rect 1104 23979 1144 24011
rect 1176 23979 1216 24011
rect 1248 23979 1288 24011
rect 1320 23979 1360 24011
rect 1392 23979 1432 24011
rect 1464 23979 1504 24011
rect 1536 23979 1576 24011
rect 1608 23979 1648 24011
rect 1680 23979 1720 24011
rect 1752 23979 1792 24011
rect 1824 23979 1864 24011
rect 1896 23979 1936 24011
rect 1968 23979 2008 24011
rect 2040 23979 2080 24011
rect 2112 23979 2152 24011
rect 2184 23979 2224 24011
rect 2256 23979 2296 24011
rect 2328 23979 2368 24011
rect 2400 23979 2440 24011
rect 2472 23979 2512 24011
rect 2544 23979 2584 24011
rect 2616 23979 2656 24011
rect 2688 23979 2728 24011
rect 2760 23979 2800 24011
rect 2832 23979 2872 24011
rect 2904 23979 2944 24011
rect 2976 23979 3016 24011
rect 3048 23979 3088 24011
rect 3120 23979 3160 24011
rect 3192 23979 3232 24011
rect 3264 23979 3304 24011
rect 3336 23979 3376 24011
rect 3408 23979 3448 24011
rect 3480 23979 3520 24011
rect 3552 23979 3592 24011
rect 3624 23979 3664 24011
rect 3696 23979 3736 24011
rect 3768 23979 3808 24011
rect 3840 23979 3880 24011
rect 3912 23979 3952 24011
rect 3984 23979 4024 24011
rect 4056 23979 4096 24011
rect 4128 23979 4168 24011
rect 4200 23979 4240 24011
rect 4272 23979 4312 24011
rect 4344 23979 4384 24011
rect 4416 23979 4456 24011
rect 4488 23979 4528 24011
rect 4560 23979 4600 24011
rect 4632 23979 4672 24011
rect 4704 23979 4744 24011
rect 4776 23979 4816 24011
rect 4848 23979 4888 24011
rect 4920 23979 4960 24011
rect 4992 23979 5032 24011
rect 5064 23979 5104 24011
rect 5136 23979 5176 24011
rect 5208 23979 5248 24011
rect 5280 23979 5320 24011
rect 5352 23979 5392 24011
rect 5424 23979 5464 24011
rect 5496 23979 5536 24011
rect 5568 23979 5608 24011
rect 5640 23979 5680 24011
rect 5712 23979 5752 24011
rect 5784 23979 5824 24011
rect 5856 23979 5896 24011
rect 5928 23979 5968 24011
rect 6000 23979 6040 24011
rect 6072 23979 6112 24011
rect 6144 23979 6184 24011
rect 6216 23979 6256 24011
rect 6288 23979 6328 24011
rect 6360 23979 6400 24011
rect 6432 23979 6472 24011
rect 6504 23979 6544 24011
rect 6576 23979 6616 24011
rect 6648 23979 6688 24011
rect 6720 23979 6760 24011
rect 6792 23979 6832 24011
rect 6864 23979 6904 24011
rect 6936 23979 6976 24011
rect 7008 23979 7048 24011
rect 7080 23979 7120 24011
rect 7152 23979 7192 24011
rect 7224 23979 7264 24011
rect 7296 23979 7336 24011
rect 7368 23979 7408 24011
rect 7440 23979 7480 24011
rect 7512 23979 7552 24011
rect 7584 23979 7624 24011
rect 7656 23979 7696 24011
rect 7728 23979 7768 24011
rect 7800 23979 7840 24011
rect 7872 23979 7912 24011
rect 7944 23979 7984 24011
rect 8016 23979 8056 24011
rect 8088 23979 8128 24011
rect 8160 23979 8200 24011
rect 8232 23979 8272 24011
rect 8304 23979 8344 24011
rect 8376 23979 8416 24011
rect 8448 23979 8488 24011
rect 8520 23979 8560 24011
rect 8592 23979 8632 24011
rect 8664 23979 8704 24011
rect 8736 23979 8776 24011
rect 8808 23979 8848 24011
rect 8880 23979 8920 24011
rect 8952 23979 8992 24011
rect 9024 23979 9064 24011
rect 9096 23979 9136 24011
rect 9168 23979 9208 24011
rect 9240 23979 9280 24011
rect 9312 23979 9352 24011
rect 9384 23979 9424 24011
rect 9456 23979 9496 24011
rect 9528 23979 9568 24011
rect 9600 23979 9640 24011
rect 9672 23979 9712 24011
rect 9744 23979 9784 24011
rect 9816 23979 9856 24011
rect 9888 23979 9928 24011
rect 9960 23979 10000 24011
rect 10032 23979 10072 24011
rect 10104 23979 10144 24011
rect 10176 23979 10216 24011
rect 10248 23979 10288 24011
rect 10320 23979 10360 24011
rect 10392 23979 10432 24011
rect 10464 23979 10504 24011
rect 10536 23979 10576 24011
rect 10608 23979 10648 24011
rect 10680 23979 10720 24011
rect 10752 23979 10792 24011
rect 10824 23979 10864 24011
rect 10896 23979 10936 24011
rect 10968 23979 11008 24011
rect 11040 23979 11080 24011
rect 11112 23979 11152 24011
rect 11184 23979 11224 24011
rect 11256 23979 11296 24011
rect 11328 23979 11368 24011
rect 11400 23979 11440 24011
rect 11472 23979 11512 24011
rect 11544 23979 11584 24011
rect 11616 23979 11656 24011
rect 11688 23979 11728 24011
rect 11760 23979 11800 24011
rect 11832 23979 11872 24011
rect 11904 23979 11944 24011
rect 11976 23979 12016 24011
rect 12048 23979 12088 24011
rect 12120 23979 12160 24011
rect 12192 23979 12232 24011
rect 12264 23979 12304 24011
rect 12336 23979 12376 24011
rect 12408 23979 12448 24011
rect 12480 23979 12520 24011
rect 12552 23979 12592 24011
rect 12624 23979 12664 24011
rect 12696 23979 12736 24011
rect 12768 23979 12808 24011
rect 12840 23979 12880 24011
rect 12912 23979 12952 24011
rect 12984 23979 13024 24011
rect 13056 23979 13096 24011
rect 13128 23979 13168 24011
rect 13200 23979 13240 24011
rect 13272 23979 13312 24011
rect 13344 23979 13384 24011
rect 13416 23979 13456 24011
rect 13488 23979 13528 24011
rect 13560 23979 13600 24011
rect 13632 23979 13672 24011
rect 13704 23979 13744 24011
rect 13776 23979 13816 24011
rect 13848 23979 13888 24011
rect 13920 23979 13960 24011
rect 13992 23979 14032 24011
rect 14064 23979 14104 24011
rect 14136 23979 14176 24011
rect 14208 23979 14248 24011
rect 14280 23979 14320 24011
rect 14352 23979 14392 24011
rect 14424 23979 14464 24011
rect 14496 23979 14536 24011
rect 14568 23979 14608 24011
rect 14640 23979 14680 24011
rect 14712 23979 14752 24011
rect 14784 23979 14824 24011
rect 14856 23979 14896 24011
rect 14928 23979 14968 24011
rect 15000 23979 15040 24011
rect 15072 23979 15112 24011
rect 15144 23979 15184 24011
rect 15216 23979 15256 24011
rect 15288 23979 15328 24011
rect 15360 23979 15400 24011
rect 15432 23979 15472 24011
rect 15504 23979 15544 24011
rect 15576 23979 15616 24011
rect 15648 23979 15688 24011
rect 15720 23979 15760 24011
rect 15792 23979 15832 24011
rect 15864 23979 15904 24011
rect 15936 23979 16000 24011
rect 0 23939 16000 23979
rect 0 23907 64 23939
rect 96 23907 136 23939
rect 168 23907 208 23939
rect 240 23907 280 23939
rect 312 23907 352 23939
rect 384 23907 424 23939
rect 456 23907 496 23939
rect 528 23907 568 23939
rect 600 23907 640 23939
rect 672 23907 712 23939
rect 744 23907 784 23939
rect 816 23907 856 23939
rect 888 23907 928 23939
rect 960 23907 1000 23939
rect 1032 23907 1072 23939
rect 1104 23907 1144 23939
rect 1176 23907 1216 23939
rect 1248 23907 1288 23939
rect 1320 23907 1360 23939
rect 1392 23907 1432 23939
rect 1464 23907 1504 23939
rect 1536 23907 1576 23939
rect 1608 23907 1648 23939
rect 1680 23907 1720 23939
rect 1752 23907 1792 23939
rect 1824 23907 1864 23939
rect 1896 23907 1936 23939
rect 1968 23907 2008 23939
rect 2040 23907 2080 23939
rect 2112 23907 2152 23939
rect 2184 23907 2224 23939
rect 2256 23907 2296 23939
rect 2328 23907 2368 23939
rect 2400 23907 2440 23939
rect 2472 23907 2512 23939
rect 2544 23907 2584 23939
rect 2616 23907 2656 23939
rect 2688 23907 2728 23939
rect 2760 23907 2800 23939
rect 2832 23907 2872 23939
rect 2904 23907 2944 23939
rect 2976 23907 3016 23939
rect 3048 23907 3088 23939
rect 3120 23907 3160 23939
rect 3192 23907 3232 23939
rect 3264 23907 3304 23939
rect 3336 23907 3376 23939
rect 3408 23907 3448 23939
rect 3480 23907 3520 23939
rect 3552 23907 3592 23939
rect 3624 23907 3664 23939
rect 3696 23907 3736 23939
rect 3768 23907 3808 23939
rect 3840 23907 3880 23939
rect 3912 23907 3952 23939
rect 3984 23907 4024 23939
rect 4056 23907 4096 23939
rect 4128 23907 4168 23939
rect 4200 23907 4240 23939
rect 4272 23907 4312 23939
rect 4344 23907 4384 23939
rect 4416 23907 4456 23939
rect 4488 23907 4528 23939
rect 4560 23907 4600 23939
rect 4632 23907 4672 23939
rect 4704 23907 4744 23939
rect 4776 23907 4816 23939
rect 4848 23907 4888 23939
rect 4920 23907 4960 23939
rect 4992 23907 5032 23939
rect 5064 23907 5104 23939
rect 5136 23907 5176 23939
rect 5208 23907 5248 23939
rect 5280 23907 5320 23939
rect 5352 23907 5392 23939
rect 5424 23907 5464 23939
rect 5496 23907 5536 23939
rect 5568 23907 5608 23939
rect 5640 23907 5680 23939
rect 5712 23907 5752 23939
rect 5784 23907 5824 23939
rect 5856 23907 5896 23939
rect 5928 23907 5968 23939
rect 6000 23907 6040 23939
rect 6072 23907 6112 23939
rect 6144 23907 6184 23939
rect 6216 23907 6256 23939
rect 6288 23907 6328 23939
rect 6360 23907 6400 23939
rect 6432 23907 6472 23939
rect 6504 23907 6544 23939
rect 6576 23907 6616 23939
rect 6648 23907 6688 23939
rect 6720 23907 6760 23939
rect 6792 23907 6832 23939
rect 6864 23907 6904 23939
rect 6936 23907 6976 23939
rect 7008 23907 7048 23939
rect 7080 23907 7120 23939
rect 7152 23907 7192 23939
rect 7224 23907 7264 23939
rect 7296 23907 7336 23939
rect 7368 23907 7408 23939
rect 7440 23907 7480 23939
rect 7512 23907 7552 23939
rect 7584 23907 7624 23939
rect 7656 23907 7696 23939
rect 7728 23907 7768 23939
rect 7800 23907 7840 23939
rect 7872 23907 7912 23939
rect 7944 23907 7984 23939
rect 8016 23907 8056 23939
rect 8088 23907 8128 23939
rect 8160 23907 8200 23939
rect 8232 23907 8272 23939
rect 8304 23907 8344 23939
rect 8376 23907 8416 23939
rect 8448 23907 8488 23939
rect 8520 23907 8560 23939
rect 8592 23907 8632 23939
rect 8664 23907 8704 23939
rect 8736 23907 8776 23939
rect 8808 23907 8848 23939
rect 8880 23907 8920 23939
rect 8952 23907 8992 23939
rect 9024 23907 9064 23939
rect 9096 23907 9136 23939
rect 9168 23907 9208 23939
rect 9240 23907 9280 23939
rect 9312 23907 9352 23939
rect 9384 23907 9424 23939
rect 9456 23907 9496 23939
rect 9528 23907 9568 23939
rect 9600 23907 9640 23939
rect 9672 23907 9712 23939
rect 9744 23907 9784 23939
rect 9816 23907 9856 23939
rect 9888 23907 9928 23939
rect 9960 23907 10000 23939
rect 10032 23907 10072 23939
rect 10104 23907 10144 23939
rect 10176 23907 10216 23939
rect 10248 23907 10288 23939
rect 10320 23907 10360 23939
rect 10392 23907 10432 23939
rect 10464 23907 10504 23939
rect 10536 23907 10576 23939
rect 10608 23907 10648 23939
rect 10680 23907 10720 23939
rect 10752 23907 10792 23939
rect 10824 23907 10864 23939
rect 10896 23907 10936 23939
rect 10968 23907 11008 23939
rect 11040 23907 11080 23939
rect 11112 23907 11152 23939
rect 11184 23907 11224 23939
rect 11256 23907 11296 23939
rect 11328 23907 11368 23939
rect 11400 23907 11440 23939
rect 11472 23907 11512 23939
rect 11544 23907 11584 23939
rect 11616 23907 11656 23939
rect 11688 23907 11728 23939
rect 11760 23907 11800 23939
rect 11832 23907 11872 23939
rect 11904 23907 11944 23939
rect 11976 23907 12016 23939
rect 12048 23907 12088 23939
rect 12120 23907 12160 23939
rect 12192 23907 12232 23939
rect 12264 23907 12304 23939
rect 12336 23907 12376 23939
rect 12408 23907 12448 23939
rect 12480 23907 12520 23939
rect 12552 23907 12592 23939
rect 12624 23907 12664 23939
rect 12696 23907 12736 23939
rect 12768 23907 12808 23939
rect 12840 23907 12880 23939
rect 12912 23907 12952 23939
rect 12984 23907 13024 23939
rect 13056 23907 13096 23939
rect 13128 23907 13168 23939
rect 13200 23907 13240 23939
rect 13272 23907 13312 23939
rect 13344 23907 13384 23939
rect 13416 23907 13456 23939
rect 13488 23907 13528 23939
rect 13560 23907 13600 23939
rect 13632 23907 13672 23939
rect 13704 23907 13744 23939
rect 13776 23907 13816 23939
rect 13848 23907 13888 23939
rect 13920 23907 13960 23939
rect 13992 23907 14032 23939
rect 14064 23907 14104 23939
rect 14136 23907 14176 23939
rect 14208 23907 14248 23939
rect 14280 23907 14320 23939
rect 14352 23907 14392 23939
rect 14424 23907 14464 23939
rect 14496 23907 14536 23939
rect 14568 23907 14608 23939
rect 14640 23907 14680 23939
rect 14712 23907 14752 23939
rect 14784 23907 14824 23939
rect 14856 23907 14896 23939
rect 14928 23907 14968 23939
rect 15000 23907 15040 23939
rect 15072 23907 15112 23939
rect 15144 23907 15184 23939
rect 15216 23907 15256 23939
rect 15288 23907 15328 23939
rect 15360 23907 15400 23939
rect 15432 23907 15472 23939
rect 15504 23907 15544 23939
rect 15576 23907 15616 23939
rect 15648 23907 15688 23939
rect 15720 23907 15760 23939
rect 15792 23907 15832 23939
rect 15864 23907 15904 23939
rect 15936 23907 16000 23939
rect 0 23867 16000 23907
rect 0 23835 64 23867
rect 96 23835 136 23867
rect 168 23835 208 23867
rect 240 23835 280 23867
rect 312 23835 352 23867
rect 384 23835 424 23867
rect 456 23835 496 23867
rect 528 23835 568 23867
rect 600 23835 640 23867
rect 672 23835 712 23867
rect 744 23835 784 23867
rect 816 23835 856 23867
rect 888 23835 928 23867
rect 960 23835 1000 23867
rect 1032 23835 1072 23867
rect 1104 23835 1144 23867
rect 1176 23835 1216 23867
rect 1248 23835 1288 23867
rect 1320 23835 1360 23867
rect 1392 23835 1432 23867
rect 1464 23835 1504 23867
rect 1536 23835 1576 23867
rect 1608 23835 1648 23867
rect 1680 23835 1720 23867
rect 1752 23835 1792 23867
rect 1824 23835 1864 23867
rect 1896 23835 1936 23867
rect 1968 23835 2008 23867
rect 2040 23835 2080 23867
rect 2112 23835 2152 23867
rect 2184 23835 2224 23867
rect 2256 23835 2296 23867
rect 2328 23835 2368 23867
rect 2400 23835 2440 23867
rect 2472 23835 2512 23867
rect 2544 23835 2584 23867
rect 2616 23835 2656 23867
rect 2688 23835 2728 23867
rect 2760 23835 2800 23867
rect 2832 23835 2872 23867
rect 2904 23835 2944 23867
rect 2976 23835 3016 23867
rect 3048 23835 3088 23867
rect 3120 23835 3160 23867
rect 3192 23835 3232 23867
rect 3264 23835 3304 23867
rect 3336 23835 3376 23867
rect 3408 23835 3448 23867
rect 3480 23835 3520 23867
rect 3552 23835 3592 23867
rect 3624 23835 3664 23867
rect 3696 23835 3736 23867
rect 3768 23835 3808 23867
rect 3840 23835 3880 23867
rect 3912 23835 3952 23867
rect 3984 23835 4024 23867
rect 4056 23835 4096 23867
rect 4128 23835 4168 23867
rect 4200 23835 4240 23867
rect 4272 23835 4312 23867
rect 4344 23835 4384 23867
rect 4416 23835 4456 23867
rect 4488 23835 4528 23867
rect 4560 23835 4600 23867
rect 4632 23835 4672 23867
rect 4704 23835 4744 23867
rect 4776 23835 4816 23867
rect 4848 23835 4888 23867
rect 4920 23835 4960 23867
rect 4992 23835 5032 23867
rect 5064 23835 5104 23867
rect 5136 23835 5176 23867
rect 5208 23835 5248 23867
rect 5280 23835 5320 23867
rect 5352 23835 5392 23867
rect 5424 23835 5464 23867
rect 5496 23835 5536 23867
rect 5568 23835 5608 23867
rect 5640 23835 5680 23867
rect 5712 23835 5752 23867
rect 5784 23835 5824 23867
rect 5856 23835 5896 23867
rect 5928 23835 5968 23867
rect 6000 23835 6040 23867
rect 6072 23835 6112 23867
rect 6144 23835 6184 23867
rect 6216 23835 6256 23867
rect 6288 23835 6328 23867
rect 6360 23835 6400 23867
rect 6432 23835 6472 23867
rect 6504 23835 6544 23867
rect 6576 23835 6616 23867
rect 6648 23835 6688 23867
rect 6720 23835 6760 23867
rect 6792 23835 6832 23867
rect 6864 23835 6904 23867
rect 6936 23835 6976 23867
rect 7008 23835 7048 23867
rect 7080 23835 7120 23867
rect 7152 23835 7192 23867
rect 7224 23835 7264 23867
rect 7296 23835 7336 23867
rect 7368 23835 7408 23867
rect 7440 23835 7480 23867
rect 7512 23835 7552 23867
rect 7584 23835 7624 23867
rect 7656 23835 7696 23867
rect 7728 23835 7768 23867
rect 7800 23835 7840 23867
rect 7872 23835 7912 23867
rect 7944 23835 7984 23867
rect 8016 23835 8056 23867
rect 8088 23835 8128 23867
rect 8160 23835 8200 23867
rect 8232 23835 8272 23867
rect 8304 23835 8344 23867
rect 8376 23835 8416 23867
rect 8448 23835 8488 23867
rect 8520 23835 8560 23867
rect 8592 23835 8632 23867
rect 8664 23835 8704 23867
rect 8736 23835 8776 23867
rect 8808 23835 8848 23867
rect 8880 23835 8920 23867
rect 8952 23835 8992 23867
rect 9024 23835 9064 23867
rect 9096 23835 9136 23867
rect 9168 23835 9208 23867
rect 9240 23835 9280 23867
rect 9312 23835 9352 23867
rect 9384 23835 9424 23867
rect 9456 23835 9496 23867
rect 9528 23835 9568 23867
rect 9600 23835 9640 23867
rect 9672 23835 9712 23867
rect 9744 23835 9784 23867
rect 9816 23835 9856 23867
rect 9888 23835 9928 23867
rect 9960 23835 10000 23867
rect 10032 23835 10072 23867
rect 10104 23835 10144 23867
rect 10176 23835 10216 23867
rect 10248 23835 10288 23867
rect 10320 23835 10360 23867
rect 10392 23835 10432 23867
rect 10464 23835 10504 23867
rect 10536 23835 10576 23867
rect 10608 23835 10648 23867
rect 10680 23835 10720 23867
rect 10752 23835 10792 23867
rect 10824 23835 10864 23867
rect 10896 23835 10936 23867
rect 10968 23835 11008 23867
rect 11040 23835 11080 23867
rect 11112 23835 11152 23867
rect 11184 23835 11224 23867
rect 11256 23835 11296 23867
rect 11328 23835 11368 23867
rect 11400 23835 11440 23867
rect 11472 23835 11512 23867
rect 11544 23835 11584 23867
rect 11616 23835 11656 23867
rect 11688 23835 11728 23867
rect 11760 23835 11800 23867
rect 11832 23835 11872 23867
rect 11904 23835 11944 23867
rect 11976 23835 12016 23867
rect 12048 23835 12088 23867
rect 12120 23835 12160 23867
rect 12192 23835 12232 23867
rect 12264 23835 12304 23867
rect 12336 23835 12376 23867
rect 12408 23835 12448 23867
rect 12480 23835 12520 23867
rect 12552 23835 12592 23867
rect 12624 23835 12664 23867
rect 12696 23835 12736 23867
rect 12768 23835 12808 23867
rect 12840 23835 12880 23867
rect 12912 23835 12952 23867
rect 12984 23835 13024 23867
rect 13056 23835 13096 23867
rect 13128 23835 13168 23867
rect 13200 23835 13240 23867
rect 13272 23835 13312 23867
rect 13344 23835 13384 23867
rect 13416 23835 13456 23867
rect 13488 23835 13528 23867
rect 13560 23835 13600 23867
rect 13632 23835 13672 23867
rect 13704 23835 13744 23867
rect 13776 23835 13816 23867
rect 13848 23835 13888 23867
rect 13920 23835 13960 23867
rect 13992 23835 14032 23867
rect 14064 23835 14104 23867
rect 14136 23835 14176 23867
rect 14208 23835 14248 23867
rect 14280 23835 14320 23867
rect 14352 23835 14392 23867
rect 14424 23835 14464 23867
rect 14496 23835 14536 23867
rect 14568 23835 14608 23867
rect 14640 23835 14680 23867
rect 14712 23835 14752 23867
rect 14784 23835 14824 23867
rect 14856 23835 14896 23867
rect 14928 23835 14968 23867
rect 15000 23835 15040 23867
rect 15072 23835 15112 23867
rect 15144 23835 15184 23867
rect 15216 23835 15256 23867
rect 15288 23835 15328 23867
rect 15360 23835 15400 23867
rect 15432 23835 15472 23867
rect 15504 23835 15544 23867
rect 15576 23835 15616 23867
rect 15648 23835 15688 23867
rect 15720 23835 15760 23867
rect 15792 23835 15832 23867
rect 15864 23835 15904 23867
rect 15936 23835 16000 23867
rect 0 23795 16000 23835
rect 0 23763 64 23795
rect 96 23763 136 23795
rect 168 23763 208 23795
rect 240 23763 280 23795
rect 312 23763 352 23795
rect 384 23763 424 23795
rect 456 23763 496 23795
rect 528 23763 568 23795
rect 600 23763 640 23795
rect 672 23763 712 23795
rect 744 23763 784 23795
rect 816 23763 856 23795
rect 888 23763 928 23795
rect 960 23763 1000 23795
rect 1032 23763 1072 23795
rect 1104 23763 1144 23795
rect 1176 23763 1216 23795
rect 1248 23763 1288 23795
rect 1320 23763 1360 23795
rect 1392 23763 1432 23795
rect 1464 23763 1504 23795
rect 1536 23763 1576 23795
rect 1608 23763 1648 23795
rect 1680 23763 1720 23795
rect 1752 23763 1792 23795
rect 1824 23763 1864 23795
rect 1896 23763 1936 23795
rect 1968 23763 2008 23795
rect 2040 23763 2080 23795
rect 2112 23763 2152 23795
rect 2184 23763 2224 23795
rect 2256 23763 2296 23795
rect 2328 23763 2368 23795
rect 2400 23763 2440 23795
rect 2472 23763 2512 23795
rect 2544 23763 2584 23795
rect 2616 23763 2656 23795
rect 2688 23763 2728 23795
rect 2760 23763 2800 23795
rect 2832 23763 2872 23795
rect 2904 23763 2944 23795
rect 2976 23763 3016 23795
rect 3048 23763 3088 23795
rect 3120 23763 3160 23795
rect 3192 23763 3232 23795
rect 3264 23763 3304 23795
rect 3336 23763 3376 23795
rect 3408 23763 3448 23795
rect 3480 23763 3520 23795
rect 3552 23763 3592 23795
rect 3624 23763 3664 23795
rect 3696 23763 3736 23795
rect 3768 23763 3808 23795
rect 3840 23763 3880 23795
rect 3912 23763 3952 23795
rect 3984 23763 4024 23795
rect 4056 23763 4096 23795
rect 4128 23763 4168 23795
rect 4200 23763 4240 23795
rect 4272 23763 4312 23795
rect 4344 23763 4384 23795
rect 4416 23763 4456 23795
rect 4488 23763 4528 23795
rect 4560 23763 4600 23795
rect 4632 23763 4672 23795
rect 4704 23763 4744 23795
rect 4776 23763 4816 23795
rect 4848 23763 4888 23795
rect 4920 23763 4960 23795
rect 4992 23763 5032 23795
rect 5064 23763 5104 23795
rect 5136 23763 5176 23795
rect 5208 23763 5248 23795
rect 5280 23763 5320 23795
rect 5352 23763 5392 23795
rect 5424 23763 5464 23795
rect 5496 23763 5536 23795
rect 5568 23763 5608 23795
rect 5640 23763 5680 23795
rect 5712 23763 5752 23795
rect 5784 23763 5824 23795
rect 5856 23763 5896 23795
rect 5928 23763 5968 23795
rect 6000 23763 6040 23795
rect 6072 23763 6112 23795
rect 6144 23763 6184 23795
rect 6216 23763 6256 23795
rect 6288 23763 6328 23795
rect 6360 23763 6400 23795
rect 6432 23763 6472 23795
rect 6504 23763 6544 23795
rect 6576 23763 6616 23795
rect 6648 23763 6688 23795
rect 6720 23763 6760 23795
rect 6792 23763 6832 23795
rect 6864 23763 6904 23795
rect 6936 23763 6976 23795
rect 7008 23763 7048 23795
rect 7080 23763 7120 23795
rect 7152 23763 7192 23795
rect 7224 23763 7264 23795
rect 7296 23763 7336 23795
rect 7368 23763 7408 23795
rect 7440 23763 7480 23795
rect 7512 23763 7552 23795
rect 7584 23763 7624 23795
rect 7656 23763 7696 23795
rect 7728 23763 7768 23795
rect 7800 23763 7840 23795
rect 7872 23763 7912 23795
rect 7944 23763 7984 23795
rect 8016 23763 8056 23795
rect 8088 23763 8128 23795
rect 8160 23763 8200 23795
rect 8232 23763 8272 23795
rect 8304 23763 8344 23795
rect 8376 23763 8416 23795
rect 8448 23763 8488 23795
rect 8520 23763 8560 23795
rect 8592 23763 8632 23795
rect 8664 23763 8704 23795
rect 8736 23763 8776 23795
rect 8808 23763 8848 23795
rect 8880 23763 8920 23795
rect 8952 23763 8992 23795
rect 9024 23763 9064 23795
rect 9096 23763 9136 23795
rect 9168 23763 9208 23795
rect 9240 23763 9280 23795
rect 9312 23763 9352 23795
rect 9384 23763 9424 23795
rect 9456 23763 9496 23795
rect 9528 23763 9568 23795
rect 9600 23763 9640 23795
rect 9672 23763 9712 23795
rect 9744 23763 9784 23795
rect 9816 23763 9856 23795
rect 9888 23763 9928 23795
rect 9960 23763 10000 23795
rect 10032 23763 10072 23795
rect 10104 23763 10144 23795
rect 10176 23763 10216 23795
rect 10248 23763 10288 23795
rect 10320 23763 10360 23795
rect 10392 23763 10432 23795
rect 10464 23763 10504 23795
rect 10536 23763 10576 23795
rect 10608 23763 10648 23795
rect 10680 23763 10720 23795
rect 10752 23763 10792 23795
rect 10824 23763 10864 23795
rect 10896 23763 10936 23795
rect 10968 23763 11008 23795
rect 11040 23763 11080 23795
rect 11112 23763 11152 23795
rect 11184 23763 11224 23795
rect 11256 23763 11296 23795
rect 11328 23763 11368 23795
rect 11400 23763 11440 23795
rect 11472 23763 11512 23795
rect 11544 23763 11584 23795
rect 11616 23763 11656 23795
rect 11688 23763 11728 23795
rect 11760 23763 11800 23795
rect 11832 23763 11872 23795
rect 11904 23763 11944 23795
rect 11976 23763 12016 23795
rect 12048 23763 12088 23795
rect 12120 23763 12160 23795
rect 12192 23763 12232 23795
rect 12264 23763 12304 23795
rect 12336 23763 12376 23795
rect 12408 23763 12448 23795
rect 12480 23763 12520 23795
rect 12552 23763 12592 23795
rect 12624 23763 12664 23795
rect 12696 23763 12736 23795
rect 12768 23763 12808 23795
rect 12840 23763 12880 23795
rect 12912 23763 12952 23795
rect 12984 23763 13024 23795
rect 13056 23763 13096 23795
rect 13128 23763 13168 23795
rect 13200 23763 13240 23795
rect 13272 23763 13312 23795
rect 13344 23763 13384 23795
rect 13416 23763 13456 23795
rect 13488 23763 13528 23795
rect 13560 23763 13600 23795
rect 13632 23763 13672 23795
rect 13704 23763 13744 23795
rect 13776 23763 13816 23795
rect 13848 23763 13888 23795
rect 13920 23763 13960 23795
rect 13992 23763 14032 23795
rect 14064 23763 14104 23795
rect 14136 23763 14176 23795
rect 14208 23763 14248 23795
rect 14280 23763 14320 23795
rect 14352 23763 14392 23795
rect 14424 23763 14464 23795
rect 14496 23763 14536 23795
rect 14568 23763 14608 23795
rect 14640 23763 14680 23795
rect 14712 23763 14752 23795
rect 14784 23763 14824 23795
rect 14856 23763 14896 23795
rect 14928 23763 14968 23795
rect 15000 23763 15040 23795
rect 15072 23763 15112 23795
rect 15144 23763 15184 23795
rect 15216 23763 15256 23795
rect 15288 23763 15328 23795
rect 15360 23763 15400 23795
rect 15432 23763 15472 23795
rect 15504 23763 15544 23795
rect 15576 23763 15616 23795
rect 15648 23763 15688 23795
rect 15720 23763 15760 23795
rect 15792 23763 15832 23795
rect 15864 23763 15904 23795
rect 15936 23763 16000 23795
rect 0 23723 16000 23763
rect 0 23691 64 23723
rect 96 23691 136 23723
rect 168 23691 208 23723
rect 240 23691 280 23723
rect 312 23691 352 23723
rect 384 23691 424 23723
rect 456 23691 496 23723
rect 528 23691 568 23723
rect 600 23691 640 23723
rect 672 23691 712 23723
rect 744 23691 784 23723
rect 816 23691 856 23723
rect 888 23691 928 23723
rect 960 23691 1000 23723
rect 1032 23691 1072 23723
rect 1104 23691 1144 23723
rect 1176 23691 1216 23723
rect 1248 23691 1288 23723
rect 1320 23691 1360 23723
rect 1392 23691 1432 23723
rect 1464 23691 1504 23723
rect 1536 23691 1576 23723
rect 1608 23691 1648 23723
rect 1680 23691 1720 23723
rect 1752 23691 1792 23723
rect 1824 23691 1864 23723
rect 1896 23691 1936 23723
rect 1968 23691 2008 23723
rect 2040 23691 2080 23723
rect 2112 23691 2152 23723
rect 2184 23691 2224 23723
rect 2256 23691 2296 23723
rect 2328 23691 2368 23723
rect 2400 23691 2440 23723
rect 2472 23691 2512 23723
rect 2544 23691 2584 23723
rect 2616 23691 2656 23723
rect 2688 23691 2728 23723
rect 2760 23691 2800 23723
rect 2832 23691 2872 23723
rect 2904 23691 2944 23723
rect 2976 23691 3016 23723
rect 3048 23691 3088 23723
rect 3120 23691 3160 23723
rect 3192 23691 3232 23723
rect 3264 23691 3304 23723
rect 3336 23691 3376 23723
rect 3408 23691 3448 23723
rect 3480 23691 3520 23723
rect 3552 23691 3592 23723
rect 3624 23691 3664 23723
rect 3696 23691 3736 23723
rect 3768 23691 3808 23723
rect 3840 23691 3880 23723
rect 3912 23691 3952 23723
rect 3984 23691 4024 23723
rect 4056 23691 4096 23723
rect 4128 23691 4168 23723
rect 4200 23691 4240 23723
rect 4272 23691 4312 23723
rect 4344 23691 4384 23723
rect 4416 23691 4456 23723
rect 4488 23691 4528 23723
rect 4560 23691 4600 23723
rect 4632 23691 4672 23723
rect 4704 23691 4744 23723
rect 4776 23691 4816 23723
rect 4848 23691 4888 23723
rect 4920 23691 4960 23723
rect 4992 23691 5032 23723
rect 5064 23691 5104 23723
rect 5136 23691 5176 23723
rect 5208 23691 5248 23723
rect 5280 23691 5320 23723
rect 5352 23691 5392 23723
rect 5424 23691 5464 23723
rect 5496 23691 5536 23723
rect 5568 23691 5608 23723
rect 5640 23691 5680 23723
rect 5712 23691 5752 23723
rect 5784 23691 5824 23723
rect 5856 23691 5896 23723
rect 5928 23691 5968 23723
rect 6000 23691 6040 23723
rect 6072 23691 6112 23723
rect 6144 23691 6184 23723
rect 6216 23691 6256 23723
rect 6288 23691 6328 23723
rect 6360 23691 6400 23723
rect 6432 23691 6472 23723
rect 6504 23691 6544 23723
rect 6576 23691 6616 23723
rect 6648 23691 6688 23723
rect 6720 23691 6760 23723
rect 6792 23691 6832 23723
rect 6864 23691 6904 23723
rect 6936 23691 6976 23723
rect 7008 23691 7048 23723
rect 7080 23691 7120 23723
rect 7152 23691 7192 23723
rect 7224 23691 7264 23723
rect 7296 23691 7336 23723
rect 7368 23691 7408 23723
rect 7440 23691 7480 23723
rect 7512 23691 7552 23723
rect 7584 23691 7624 23723
rect 7656 23691 7696 23723
rect 7728 23691 7768 23723
rect 7800 23691 7840 23723
rect 7872 23691 7912 23723
rect 7944 23691 7984 23723
rect 8016 23691 8056 23723
rect 8088 23691 8128 23723
rect 8160 23691 8200 23723
rect 8232 23691 8272 23723
rect 8304 23691 8344 23723
rect 8376 23691 8416 23723
rect 8448 23691 8488 23723
rect 8520 23691 8560 23723
rect 8592 23691 8632 23723
rect 8664 23691 8704 23723
rect 8736 23691 8776 23723
rect 8808 23691 8848 23723
rect 8880 23691 8920 23723
rect 8952 23691 8992 23723
rect 9024 23691 9064 23723
rect 9096 23691 9136 23723
rect 9168 23691 9208 23723
rect 9240 23691 9280 23723
rect 9312 23691 9352 23723
rect 9384 23691 9424 23723
rect 9456 23691 9496 23723
rect 9528 23691 9568 23723
rect 9600 23691 9640 23723
rect 9672 23691 9712 23723
rect 9744 23691 9784 23723
rect 9816 23691 9856 23723
rect 9888 23691 9928 23723
rect 9960 23691 10000 23723
rect 10032 23691 10072 23723
rect 10104 23691 10144 23723
rect 10176 23691 10216 23723
rect 10248 23691 10288 23723
rect 10320 23691 10360 23723
rect 10392 23691 10432 23723
rect 10464 23691 10504 23723
rect 10536 23691 10576 23723
rect 10608 23691 10648 23723
rect 10680 23691 10720 23723
rect 10752 23691 10792 23723
rect 10824 23691 10864 23723
rect 10896 23691 10936 23723
rect 10968 23691 11008 23723
rect 11040 23691 11080 23723
rect 11112 23691 11152 23723
rect 11184 23691 11224 23723
rect 11256 23691 11296 23723
rect 11328 23691 11368 23723
rect 11400 23691 11440 23723
rect 11472 23691 11512 23723
rect 11544 23691 11584 23723
rect 11616 23691 11656 23723
rect 11688 23691 11728 23723
rect 11760 23691 11800 23723
rect 11832 23691 11872 23723
rect 11904 23691 11944 23723
rect 11976 23691 12016 23723
rect 12048 23691 12088 23723
rect 12120 23691 12160 23723
rect 12192 23691 12232 23723
rect 12264 23691 12304 23723
rect 12336 23691 12376 23723
rect 12408 23691 12448 23723
rect 12480 23691 12520 23723
rect 12552 23691 12592 23723
rect 12624 23691 12664 23723
rect 12696 23691 12736 23723
rect 12768 23691 12808 23723
rect 12840 23691 12880 23723
rect 12912 23691 12952 23723
rect 12984 23691 13024 23723
rect 13056 23691 13096 23723
rect 13128 23691 13168 23723
rect 13200 23691 13240 23723
rect 13272 23691 13312 23723
rect 13344 23691 13384 23723
rect 13416 23691 13456 23723
rect 13488 23691 13528 23723
rect 13560 23691 13600 23723
rect 13632 23691 13672 23723
rect 13704 23691 13744 23723
rect 13776 23691 13816 23723
rect 13848 23691 13888 23723
rect 13920 23691 13960 23723
rect 13992 23691 14032 23723
rect 14064 23691 14104 23723
rect 14136 23691 14176 23723
rect 14208 23691 14248 23723
rect 14280 23691 14320 23723
rect 14352 23691 14392 23723
rect 14424 23691 14464 23723
rect 14496 23691 14536 23723
rect 14568 23691 14608 23723
rect 14640 23691 14680 23723
rect 14712 23691 14752 23723
rect 14784 23691 14824 23723
rect 14856 23691 14896 23723
rect 14928 23691 14968 23723
rect 15000 23691 15040 23723
rect 15072 23691 15112 23723
rect 15144 23691 15184 23723
rect 15216 23691 15256 23723
rect 15288 23691 15328 23723
rect 15360 23691 15400 23723
rect 15432 23691 15472 23723
rect 15504 23691 15544 23723
rect 15576 23691 15616 23723
rect 15648 23691 15688 23723
rect 15720 23691 15760 23723
rect 15792 23691 15832 23723
rect 15864 23691 15904 23723
rect 15936 23691 16000 23723
rect 0 23651 16000 23691
rect 0 23619 64 23651
rect 96 23619 136 23651
rect 168 23619 208 23651
rect 240 23619 280 23651
rect 312 23619 352 23651
rect 384 23619 424 23651
rect 456 23619 496 23651
rect 528 23619 568 23651
rect 600 23619 640 23651
rect 672 23619 712 23651
rect 744 23619 784 23651
rect 816 23619 856 23651
rect 888 23619 928 23651
rect 960 23619 1000 23651
rect 1032 23619 1072 23651
rect 1104 23619 1144 23651
rect 1176 23619 1216 23651
rect 1248 23619 1288 23651
rect 1320 23619 1360 23651
rect 1392 23619 1432 23651
rect 1464 23619 1504 23651
rect 1536 23619 1576 23651
rect 1608 23619 1648 23651
rect 1680 23619 1720 23651
rect 1752 23619 1792 23651
rect 1824 23619 1864 23651
rect 1896 23619 1936 23651
rect 1968 23619 2008 23651
rect 2040 23619 2080 23651
rect 2112 23619 2152 23651
rect 2184 23619 2224 23651
rect 2256 23619 2296 23651
rect 2328 23619 2368 23651
rect 2400 23619 2440 23651
rect 2472 23619 2512 23651
rect 2544 23619 2584 23651
rect 2616 23619 2656 23651
rect 2688 23619 2728 23651
rect 2760 23619 2800 23651
rect 2832 23619 2872 23651
rect 2904 23619 2944 23651
rect 2976 23619 3016 23651
rect 3048 23619 3088 23651
rect 3120 23619 3160 23651
rect 3192 23619 3232 23651
rect 3264 23619 3304 23651
rect 3336 23619 3376 23651
rect 3408 23619 3448 23651
rect 3480 23619 3520 23651
rect 3552 23619 3592 23651
rect 3624 23619 3664 23651
rect 3696 23619 3736 23651
rect 3768 23619 3808 23651
rect 3840 23619 3880 23651
rect 3912 23619 3952 23651
rect 3984 23619 4024 23651
rect 4056 23619 4096 23651
rect 4128 23619 4168 23651
rect 4200 23619 4240 23651
rect 4272 23619 4312 23651
rect 4344 23619 4384 23651
rect 4416 23619 4456 23651
rect 4488 23619 4528 23651
rect 4560 23619 4600 23651
rect 4632 23619 4672 23651
rect 4704 23619 4744 23651
rect 4776 23619 4816 23651
rect 4848 23619 4888 23651
rect 4920 23619 4960 23651
rect 4992 23619 5032 23651
rect 5064 23619 5104 23651
rect 5136 23619 5176 23651
rect 5208 23619 5248 23651
rect 5280 23619 5320 23651
rect 5352 23619 5392 23651
rect 5424 23619 5464 23651
rect 5496 23619 5536 23651
rect 5568 23619 5608 23651
rect 5640 23619 5680 23651
rect 5712 23619 5752 23651
rect 5784 23619 5824 23651
rect 5856 23619 5896 23651
rect 5928 23619 5968 23651
rect 6000 23619 6040 23651
rect 6072 23619 6112 23651
rect 6144 23619 6184 23651
rect 6216 23619 6256 23651
rect 6288 23619 6328 23651
rect 6360 23619 6400 23651
rect 6432 23619 6472 23651
rect 6504 23619 6544 23651
rect 6576 23619 6616 23651
rect 6648 23619 6688 23651
rect 6720 23619 6760 23651
rect 6792 23619 6832 23651
rect 6864 23619 6904 23651
rect 6936 23619 6976 23651
rect 7008 23619 7048 23651
rect 7080 23619 7120 23651
rect 7152 23619 7192 23651
rect 7224 23619 7264 23651
rect 7296 23619 7336 23651
rect 7368 23619 7408 23651
rect 7440 23619 7480 23651
rect 7512 23619 7552 23651
rect 7584 23619 7624 23651
rect 7656 23619 7696 23651
rect 7728 23619 7768 23651
rect 7800 23619 7840 23651
rect 7872 23619 7912 23651
rect 7944 23619 7984 23651
rect 8016 23619 8056 23651
rect 8088 23619 8128 23651
rect 8160 23619 8200 23651
rect 8232 23619 8272 23651
rect 8304 23619 8344 23651
rect 8376 23619 8416 23651
rect 8448 23619 8488 23651
rect 8520 23619 8560 23651
rect 8592 23619 8632 23651
rect 8664 23619 8704 23651
rect 8736 23619 8776 23651
rect 8808 23619 8848 23651
rect 8880 23619 8920 23651
rect 8952 23619 8992 23651
rect 9024 23619 9064 23651
rect 9096 23619 9136 23651
rect 9168 23619 9208 23651
rect 9240 23619 9280 23651
rect 9312 23619 9352 23651
rect 9384 23619 9424 23651
rect 9456 23619 9496 23651
rect 9528 23619 9568 23651
rect 9600 23619 9640 23651
rect 9672 23619 9712 23651
rect 9744 23619 9784 23651
rect 9816 23619 9856 23651
rect 9888 23619 9928 23651
rect 9960 23619 10000 23651
rect 10032 23619 10072 23651
rect 10104 23619 10144 23651
rect 10176 23619 10216 23651
rect 10248 23619 10288 23651
rect 10320 23619 10360 23651
rect 10392 23619 10432 23651
rect 10464 23619 10504 23651
rect 10536 23619 10576 23651
rect 10608 23619 10648 23651
rect 10680 23619 10720 23651
rect 10752 23619 10792 23651
rect 10824 23619 10864 23651
rect 10896 23619 10936 23651
rect 10968 23619 11008 23651
rect 11040 23619 11080 23651
rect 11112 23619 11152 23651
rect 11184 23619 11224 23651
rect 11256 23619 11296 23651
rect 11328 23619 11368 23651
rect 11400 23619 11440 23651
rect 11472 23619 11512 23651
rect 11544 23619 11584 23651
rect 11616 23619 11656 23651
rect 11688 23619 11728 23651
rect 11760 23619 11800 23651
rect 11832 23619 11872 23651
rect 11904 23619 11944 23651
rect 11976 23619 12016 23651
rect 12048 23619 12088 23651
rect 12120 23619 12160 23651
rect 12192 23619 12232 23651
rect 12264 23619 12304 23651
rect 12336 23619 12376 23651
rect 12408 23619 12448 23651
rect 12480 23619 12520 23651
rect 12552 23619 12592 23651
rect 12624 23619 12664 23651
rect 12696 23619 12736 23651
rect 12768 23619 12808 23651
rect 12840 23619 12880 23651
rect 12912 23619 12952 23651
rect 12984 23619 13024 23651
rect 13056 23619 13096 23651
rect 13128 23619 13168 23651
rect 13200 23619 13240 23651
rect 13272 23619 13312 23651
rect 13344 23619 13384 23651
rect 13416 23619 13456 23651
rect 13488 23619 13528 23651
rect 13560 23619 13600 23651
rect 13632 23619 13672 23651
rect 13704 23619 13744 23651
rect 13776 23619 13816 23651
rect 13848 23619 13888 23651
rect 13920 23619 13960 23651
rect 13992 23619 14032 23651
rect 14064 23619 14104 23651
rect 14136 23619 14176 23651
rect 14208 23619 14248 23651
rect 14280 23619 14320 23651
rect 14352 23619 14392 23651
rect 14424 23619 14464 23651
rect 14496 23619 14536 23651
rect 14568 23619 14608 23651
rect 14640 23619 14680 23651
rect 14712 23619 14752 23651
rect 14784 23619 14824 23651
rect 14856 23619 14896 23651
rect 14928 23619 14968 23651
rect 15000 23619 15040 23651
rect 15072 23619 15112 23651
rect 15144 23619 15184 23651
rect 15216 23619 15256 23651
rect 15288 23619 15328 23651
rect 15360 23619 15400 23651
rect 15432 23619 15472 23651
rect 15504 23619 15544 23651
rect 15576 23619 15616 23651
rect 15648 23619 15688 23651
rect 15720 23619 15760 23651
rect 15792 23619 15832 23651
rect 15864 23619 15904 23651
rect 15936 23619 16000 23651
rect 0 23579 16000 23619
rect 0 23547 64 23579
rect 96 23547 136 23579
rect 168 23547 208 23579
rect 240 23547 280 23579
rect 312 23547 352 23579
rect 384 23547 424 23579
rect 456 23547 496 23579
rect 528 23547 568 23579
rect 600 23547 640 23579
rect 672 23547 712 23579
rect 744 23547 784 23579
rect 816 23547 856 23579
rect 888 23547 928 23579
rect 960 23547 1000 23579
rect 1032 23547 1072 23579
rect 1104 23547 1144 23579
rect 1176 23547 1216 23579
rect 1248 23547 1288 23579
rect 1320 23547 1360 23579
rect 1392 23547 1432 23579
rect 1464 23547 1504 23579
rect 1536 23547 1576 23579
rect 1608 23547 1648 23579
rect 1680 23547 1720 23579
rect 1752 23547 1792 23579
rect 1824 23547 1864 23579
rect 1896 23547 1936 23579
rect 1968 23547 2008 23579
rect 2040 23547 2080 23579
rect 2112 23547 2152 23579
rect 2184 23547 2224 23579
rect 2256 23547 2296 23579
rect 2328 23547 2368 23579
rect 2400 23547 2440 23579
rect 2472 23547 2512 23579
rect 2544 23547 2584 23579
rect 2616 23547 2656 23579
rect 2688 23547 2728 23579
rect 2760 23547 2800 23579
rect 2832 23547 2872 23579
rect 2904 23547 2944 23579
rect 2976 23547 3016 23579
rect 3048 23547 3088 23579
rect 3120 23547 3160 23579
rect 3192 23547 3232 23579
rect 3264 23547 3304 23579
rect 3336 23547 3376 23579
rect 3408 23547 3448 23579
rect 3480 23547 3520 23579
rect 3552 23547 3592 23579
rect 3624 23547 3664 23579
rect 3696 23547 3736 23579
rect 3768 23547 3808 23579
rect 3840 23547 3880 23579
rect 3912 23547 3952 23579
rect 3984 23547 4024 23579
rect 4056 23547 4096 23579
rect 4128 23547 4168 23579
rect 4200 23547 4240 23579
rect 4272 23547 4312 23579
rect 4344 23547 4384 23579
rect 4416 23547 4456 23579
rect 4488 23547 4528 23579
rect 4560 23547 4600 23579
rect 4632 23547 4672 23579
rect 4704 23547 4744 23579
rect 4776 23547 4816 23579
rect 4848 23547 4888 23579
rect 4920 23547 4960 23579
rect 4992 23547 5032 23579
rect 5064 23547 5104 23579
rect 5136 23547 5176 23579
rect 5208 23547 5248 23579
rect 5280 23547 5320 23579
rect 5352 23547 5392 23579
rect 5424 23547 5464 23579
rect 5496 23547 5536 23579
rect 5568 23547 5608 23579
rect 5640 23547 5680 23579
rect 5712 23547 5752 23579
rect 5784 23547 5824 23579
rect 5856 23547 5896 23579
rect 5928 23547 5968 23579
rect 6000 23547 6040 23579
rect 6072 23547 6112 23579
rect 6144 23547 6184 23579
rect 6216 23547 6256 23579
rect 6288 23547 6328 23579
rect 6360 23547 6400 23579
rect 6432 23547 6472 23579
rect 6504 23547 6544 23579
rect 6576 23547 6616 23579
rect 6648 23547 6688 23579
rect 6720 23547 6760 23579
rect 6792 23547 6832 23579
rect 6864 23547 6904 23579
rect 6936 23547 6976 23579
rect 7008 23547 7048 23579
rect 7080 23547 7120 23579
rect 7152 23547 7192 23579
rect 7224 23547 7264 23579
rect 7296 23547 7336 23579
rect 7368 23547 7408 23579
rect 7440 23547 7480 23579
rect 7512 23547 7552 23579
rect 7584 23547 7624 23579
rect 7656 23547 7696 23579
rect 7728 23547 7768 23579
rect 7800 23547 7840 23579
rect 7872 23547 7912 23579
rect 7944 23547 7984 23579
rect 8016 23547 8056 23579
rect 8088 23547 8128 23579
rect 8160 23547 8200 23579
rect 8232 23547 8272 23579
rect 8304 23547 8344 23579
rect 8376 23547 8416 23579
rect 8448 23547 8488 23579
rect 8520 23547 8560 23579
rect 8592 23547 8632 23579
rect 8664 23547 8704 23579
rect 8736 23547 8776 23579
rect 8808 23547 8848 23579
rect 8880 23547 8920 23579
rect 8952 23547 8992 23579
rect 9024 23547 9064 23579
rect 9096 23547 9136 23579
rect 9168 23547 9208 23579
rect 9240 23547 9280 23579
rect 9312 23547 9352 23579
rect 9384 23547 9424 23579
rect 9456 23547 9496 23579
rect 9528 23547 9568 23579
rect 9600 23547 9640 23579
rect 9672 23547 9712 23579
rect 9744 23547 9784 23579
rect 9816 23547 9856 23579
rect 9888 23547 9928 23579
rect 9960 23547 10000 23579
rect 10032 23547 10072 23579
rect 10104 23547 10144 23579
rect 10176 23547 10216 23579
rect 10248 23547 10288 23579
rect 10320 23547 10360 23579
rect 10392 23547 10432 23579
rect 10464 23547 10504 23579
rect 10536 23547 10576 23579
rect 10608 23547 10648 23579
rect 10680 23547 10720 23579
rect 10752 23547 10792 23579
rect 10824 23547 10864 23579
rect 10896 23547 10936 23579
rect 10968 23547 11008 23579
rect 11040 23547 11080 23579
rect 11112 23547 11152 23579
rect 11184 23547 11224 23579
rect 11256 23547 11296 23579
rect 11328 23547 11368 23579
rect 11400 23547 11440 23579
rect 11472 23547 11512 23579
rect 11544 23547 11584 23579
rect 11616 23547 11656 23579
rect 11688 23547 11728 23579
rect 11760 23547 11800 23579
rect 11832 23547 11872 23579
rect 11904 23547 11944 23579
rect 11976 23547 12016 23579
rect 12048 23547 12088 23579
rect 12120 23547 12160 23579
rect 12192 23547 12232 23579
rect 12264 23547 12304 23579
rect 12336 23547 12376 23579
rect 12408 23547 12448 23579
rect 12480 23547 12520 23579
rect 12552 23547 12592 23579
rect 12624 23547 12664 23579
rect 12696 23547 12736 23579
rect 12768 23547 12808 23579
rect 12840 23547 12880 23579
rect 12912 23547 12952 23579
rect 12984 23547 13024 23579
rect 13056 23547 13096 23579
rect 13128 23547 13168 23579
rect 13200 23547 13240 23579
rect 13272 23547 13312 23579
rect 13344 23547 13384 23579
rect 13416 23547 13456 23579
rect 13488 23547 13528 23579
rect 13560 23547 13600 23579
rect 13632 23547 13672 23579
rect 13704 23547 13744 23579
rect 13776 23547 13816 23579
rect 13848 23547 13888 23579
rect 13920 23547 13960 23579
rect 13992 23547 14032 23579
rect 14064 23547 14104 23579
rect 14136 23547 14176 23579
rect 14208 23547 14248 23579
rect 14280 23547 14320 23579
rect 14352 23547 14392 23579
rect 14424 23547 14464 23579
rect 14496 23547 14536 23579
rect 14568 23547 14608 23579
rect 14640 23547 14680 23579
rect 14712 23547 14752 23579
rect 14784 23547 14824 23579
rect 14856 23547 14896 23579
rect 14928 23547 14968 23579
rect 15000 23547 15040 23579
rect 15072 23547 15112 23579
rect 15144 23547 15184 23579
rect 15216 23547 15256 23579
rect 15288 23547 15328 23579
rect 15360 23547 15400 23579
rect 15432 23547 15472 23579
rect 15504 23547 15544 23579
rect 15576 23547 15616 23579
rect 15648 23547 15688 23579
rect 15720 23547 15760 23579
rect 15792 23547 15832 23579
rect 15864 23547 15904 23579
rect 15936 23547 16000 23579
rect 0 23507 16000 23547
rect 0 23475 64 23507
rect 96 23475 136 23507
rect 168 23475 208 23507
rect 240 23475 280 23507
rect 312 23475 352 23507
rect 384 23475 424 23507
rect 456 23475 496 23507
rect 528 23475 568 23507
rect 600 23475 640 23507
rect 672 23475 712 23507
rect 744 23475 784 23507
rect 816 23475 856 23507
rect 888 23475 928 23507
rect 960 23475 1000 23507
rect 1032 23475 1072 23507
rect 1104 23475 1144 23507
rect 1176 23475 1216 23507
rect 1248 23475 1288 23507
rect 1320 23475 1360 23507
rect 1392 23475 1432 23507
rect 1464 23475 1504 23507
rect 1536 23475 1576 23507
rect 1608 23475 1648 23507
rect 1680 23475 1720 23507
rect 1752 23475 1792 23507
rect 1824 23475 1864 23507
rect 1896 23475 1936 23507
rect 1968 23475 2008 23507
rect 2040 23475 2080 23507
rect 2112 23475 2152 23507
rect 2184 23475 2224 23507
rect 2256 23475 2296 23507
rect 2328 23475 2368 23507
rect 2400 23475 2440 23507
rect 2472 23475 2512 23507
rect 2544 23475 2584 23507
rect 2616 23475 2656 23507
rect 2688 23475 2728 23507
rect 2760 23475 2800 23507
rect 2832 23475 2872 23507
rect 2904 23475 2944 23507
rect 2976 23475 3016 23507
rect 3048 23475 3088 23507
rect 3120 23475 3160 23507
rect 3192 23475 3232 23507
rect 3264 23475 3304 23507
rect 3336 23475 3376 23507
rect 3408 23475 3448 23507
rect 3480 23475 3520 23507
rect 3552 23475 3592 23507
rect 3624 23475 3664 23507
rect 3696 23475 3736 23507
rect 3768 23475 3808 23507
rect 3840 23475 3880 23507
rect 3912 23475 3952 23507
rect 3984 23475 4024 23507
rect 4056 23475 4096 23507
rect 4128 23475 4168 23507
rect 4200 23475 4240 23507
rect 4272 23475 4312 23507
rect 4344 23475 4384 23507
rect 4416 23475 4456 23507
rect 4488 23475 4528 23507
rect 4560 23475 4600 23507
rect 4632 23475 4672 23507
rect 4704 23475 4744 23507
rect 4776 23475 4816 23507
rect 4848 23475 4888 23507
rect 4920 23475 4960 23507
rect 4992 23475 5032 23507
rect 5064 23475 5104 23507
rect 5136 23475 5176 23507
rect 5208 23475 5248 23507
rect 5280 23475 5320 23507
rect 5352 23475 5392 23507
rect 5424 23475 5464 23507
rect 5496 23475 5536 23507
rect 5568 23475 5608 23507
rect 5640 23475 5680 23507
rect 5712 23475 5752 23507
rect 5784 23475 5824 23507
rect 5856 23475 5896 23507
rect 5928 23475 5968 23507
rect 6000 23475 6040 23507
rect 6072 23475 6112 23507
rect 6144 23475 6184 23507
rect 6216 23475 6256 23507
rect 6288 23475 6328 23507
rect 6360 23475 6400 23507
rect 6432 23475 6472 23507
rect 6504 23475 6544 23507
rect 6576 23475 6616 23507
rect 6648 23475 6688 23507
rect 6720 23475 6760 23507
rect 6792 23475 6832 23507
rect 6864 23475 6904 23507
rect 6936 23475 6976 23507
rect 7008 23475 7048 23507
rect 7080 23475 7120 23507
rect 7152 23475 7192 23507
rect 7224 23475 7264 23507
rect 7296 23475 7336 23507
rect 7368 23475 7408 23507
rect 7440 23475 7480 23507
rect 7512 23475 7552 23507
rect 7584 23475 7624 23507
rect 7656 23475 7696 23507
rect 7728 23475 7768 23507
rect 7800 23475 7840 23507
rect 7872 23475 7912 23507
rect 7944 23475 7984 23507
rect 8016 23475 8056 23507
rect 8088 23475 8128 23507
rect 8160 23475 8200 23507
rect 8232 23475 8272 23507
rect 8304 23475 8344 23507
rect 8376 23475 8416 23507
rect 8448 23475 8488 23507
rect 8520 23475 8560 23507
rect 8592 23475 8632 23507
rect 8664 23475 8704 23507
rect 8736 23475 8776 23507
rect 8808 23475 8848 23507
rect 8880 23475 8920 23507
rect 8952 23475 8992 23507
rect 9024 23475 9064 23507
rect 9096 23475 9136 23507
rect 9168 23475 9208 23507
rect 9240 23475 9280 23507
rect 9312 23475 9352 23507
rect 9384 23475 9424 23507
rect 9456 23475 9496 23507
rect 9528 23475 9568 23507
rect 9600 23475 9640 23507
rect 9672 23475 9712 23507
rect 9744 23475 9784 23507
rect 9816 23475 9856 23507
rect 9888 23475 9928 23507
rect 9960 23475 10000 23507
rect 10032 23475 10072 23507
rect 10104 23475 10144 23507
rect 10176 23475 10216 23507
rect 10248 23475 10288 23507
rect 10320 23475 10360 23507
rect 10392 23475 10432 23507
rect 10464 23475 10504 23507
rect 10536 23475 10576 23507
rect 10608 23475 10648 23507
rect 10680 23475 10720 23507
rect 10752 23475 10792 23507
rect 10824 23475 10864 23507
rect 10896 23475 10936 23507
rect 10968 23475 11008 23507
rect 11040 23475 11080 23507
rect 11112 23475 11152 23507
rect 11184 23475 11224 23507
rect 11256 23475 11296 23507
rect 11328 23475 11368 23507
rect 11400 23475 11440 23507
rect 11472 23475 11512 23507
rect 11544 23475 11584 23507
rect 11616 23475 11656 23507
rect 11688 23475 11728 23507
rect 11760 23475 11800 23507
rect 11832 23475 11872 23507
rect 11904 23475 11944 23507
rect 11976 23475 12016 23507
rect 12048 23475 12088 23507
rect 12120 23475 12160 23507
rect 12192 23475 12232 23507
rect 12264 23475 12304 23507
rect 12336 23475 12376 23507
rect 12408 23475 12448 23507
rect 12480 23475 12520 23507
rect 12552 23475 12592 23507
rect 12624 23475 12664 23507
rect 12696 23475 12736 23507
rect 12768 23475 12808 23507
rect 12840 23475 12880 23507
rect 12912 23475 12952 23507
rect 12984 23475 13024 23507
rect 13056 23475 13096 23507
rect 13128 23475 13168 23507
rect 13200 23475 13240 23507
rect 13272 23475 13312 23507
rect 13344 23475 13384 23507
rect 13416 23475 13456 23507
rect 13488 23475 13528 23507
rect 13560 23475 13600 23507
rect 13632 23475 13672 23507
rect 13704 23475 13744 23507
rect 13776 23475 13816 23507
rect 13848 23475 13888 23507
rect 13920 23475 13960 23507
rect 13992 23475 14032 23507
rect 14064 23475 14104 23507
rect 14136 23475 14176 23507
rect 14208 23475 14248 23507
rect 14280 23475 14320 23507
rect 14352 23475 14392 23507
rect 14424 23475 14464 23507
rect 14496 23475 14536 23507
rect 14568 23475 14608 23507
rect 14640 23475 14680 23507
rect 14712 23475 14752 23507
rect 14784 23475 14824 23507
rect 14856 23475 14896 23507
rect 14928 23475 14968 23507
rect 15000 23475 15040 23507
rect 15072 23475 15112 23507
rect 15144 23475 15184 23507
rect 15216 23475 15256 23507
rect 15288 23475 15328 23507
rect 15360 23475 15400 23507
rect 15432 23475 15472 23507
rect 15504 23475 15544 23507
rect 15576 23475 15616 23507
rect 15648 23475 15688 23507
rect 15720 23475 15760 23507
rect 15792 23475 15832 23507
rect 15864 23475 15904 23507
rect 15936 23475 16000 23507
rect 0 23435 16000 23475
rect 0 23403 64 23435
rect 96 23403 136 23435
rect 168 23403 208 23435
rect 240 23403 280 23435
rect 312 23403 352 23435
rect 384 23403 424 23435
rect 456 23403 496 23435
rect 528 23403 568 23435
rect 600 23403 640 23435
rect 672 23403 712 23435
rect 744 23403 784 23435
rect 816 23403 856 23435
rect 888 23403 928 23435
rect 960 23403 1000 23435
rect 1032 23403 1072 23435
rect 1104 23403 1144 23435
rect 1176 23403 1216 23435
rect 1248 23403 1288 23435
rect 1320 23403 1360 23435
rect 1392 23403 1432 23435
rect 1464 23403 1504 23435
rect 1536 23403 1576 23435
rect 1608 23403 1648 23435
rect 1680 23403 1720 23435
rect 1752 23403 1792 23435
rect 1824 23403 1864 23435
rect 1896 23403 1936 23435
rect 1968 23403 2008 23435
rect 2040 23403 2080 23435
rect 2112 23403 2152 23435
rect 2184 23403 2224 23435
rect 2256 23403 2296 23435
rect 2328 23403 2368 23435
rect 2400 23403 2440 23435
rect 2472 23403 2512 23435
rect 2544 23403 2584 23435
rect 2616 23403 2656 23435
rect 2688 23403 2728 23435
rect 2760 23403 2800 23435
rect 2832 23403 2872 23435
rect 2904 23403 2944 23435
rect 2976 23403 3016 23435
rect 3048 23403 3088 23435
rect 3120 23403 3160 23435
rect 3192 23403 3232 23435
rect 3264 23403 3304 23435
rect 3336 23403 3376 23435
rect 3408 23403 3448 23435
rect 3480 23403 3520 23435
rect 3552 23403 3592 23435
rect 3624 23403 3664 23435
rect 3696 23403 3736 23435
rect 3768 23403 3808 23435
rect 3840 23403 3880 23435
rect 3912 23403 3952 23435
rect 3984 23403 4024 23435
rect 4056 23403 4096 23435
rect 4128 23403 4168 23435
rect 4200 23403 4240 23435
rect 4272 23403 4312 23435
rect 4344 23403 4384 23435
rect 4416 23403 4456 23435
rect 4488 23403 4528 23435
rect 4560 23403 4600 23435
rect 4632 23403 4672 23435
rect 4704 23403 4744 23435
rect 4776 23403 4816 23435
rect 4848 23403 4888 23435
rect 4920 23403 4960 23435
rect 4992 23403 5032 23435
rect 5064 23403 5104 23435
rect 5136 23403 5176 23435
rect 5208 23403 5248 23435
rect 5280 23403 5320 23435
rect 5352 23403 5392 23435
rect 5424 23403 5464 23435
rect 5496 23403 5536 23435
rect 5568 23403 5608 23435
rect 5640 23403 5680 23435
rect 5712 23403 5752 23435
rect 5784 23403 5824 23435
rect 5856 23403 5896 23435
rect 5928 23403 5968 23435
rect 6000 23403 6040 23435
rect 6072 23403 6112 23435
rect 6144 23403 6184 23435
rect 6216 23403 6256 23435
rect 6288 23403 6328 23435
rect 6360 23403 6400 23435
rect 6432 23403 6472 23435
rect 6504 23403 6544 23435
rect 6576 23403 6616 23435
rect 6648 23403 6688 23435
rect 6720 23403 6760 23435
rect 6792 23403 6832 23435
rect 6864 23403 6904 23435
rect 6936 23403 6976 23435
rect 7008 23403 7048 23435
rect 7080 23403 7120 23435
rect 7152 23403 7192 23435
rect 7224 23403 7264 23435
rect 7296 23403 7336 23435
rect 7368 23403 7408 23435
rect 7440 23403 7480 23435
rect 7512 23403 7552 23435
rect 7584 23403 7624 23435
rect 7656 23403 7696 23435
rect 7728 23403 7768 23435
rect 7800 23403 7840 23435
rect 7872 23403 7912 23435
rect 7944 23403 7984 23435
rect 8016 23403 8056 23435
rect 8088 23403 8128 23435
rect 8160 23403 8200 23435
rect 8232 23403 8272 23435
rect 8304 23403 8344 23435
rect 8376 23403 8416 23435
rect 8448 23403 8488 23435
rect 8520 23403 8560 23435
rect 8592 23403 8632 23435
rect 8664 23403 8704 23435
rect 8736 23403 8776 23435
rect 8808 23403 8848 23435
rect 8880 23403 8920 23435
rect 8952 23403 8992 23435
rect 9024 23403 9064 23435
rect 9096 23403 9136 23435
rect 9168 23403 9208 23435
rect 9240 23403 9280 23435
rect 9312 23403 9352 23435
rect 9384 23403 9424 23435
rect 9456 23403 9496 23435
rect 9528 23403 9568 23435
rect 9600 23403 9640 23435
rect 9672 23403 9712 23435
rect 9744 23403 9784 23435
rect 9816 23403 9856 23435
rect 9888 23403 9928 23435
rect 9960 23403 10000 23435
rect 10032 23403 10072 23435
rect 10104 23403 10144 23435
rect 10176 23403 10216 23435
rect 10248 23403 10288 23435
rect 10320 23403 10360 23435
rect 10392 23403 10432 23435
rect 10464 23403 10504 23435
rect 10536 23403 10576 23435
rect 10608 23403 10648 23435
rect 10680 23403 10720 23435
rect 10752 23403 10792 23435
rect 10824 23403 10864 23435
rect 10896 23403 10936 23435
rect 10968 23403 11008 23435
rect 11040 23403 11080 23435
rect 11112 23403 11152 23435
rect 11184 23403 11224 23435
rect 11256 23403 11296 23435
rect 11328 23403 11368 23435
rect 11400 23403 11440 23435
rect 11472 23403 11512 23435
rect 11544 23403 11584 23435
rect 11616 23403 11656 23435
rect 11688 23403 11728 23435
rect 11760 23403 11800 23435
rect 11832 23403 11872 23435
rect 11904 23403 11944 23435
rect 11976 23403 12016 23435
rect 12048 23403 12088 23435
rect 12120 23403 12160 23435
rect 12192 23403 12232 23435
rect 12264 23403 12304 23435
rect 12336 23403 12376 23435
rect 12408 23403 12448 23435
rect 12480 23403 12520 23435
rect 12552 23403 12592 23435
rect 12624 23403 12664 23435
rect 12696 23403 12736 23435
rect 12768 23403 12808 23435
rect 12840 23403 12880 23435
rect 12912 23403 12952 23435
rect 12984 23403 13024 23435
rect 13056 23403 13096 23435
rect 13128 23403 13168 23435
rect 13200 23403 13240 23435
rect 13272 23403 13312 23435
rect 13344 23403 13384 23435
rect 13416 23403 13456 23435
rect 13488 23403 13528 23435
rect 13560 23403 13600 23435
rect 13632 23403 13672 23435
rect 13704 23403 13744 23435
rect 13776 23403 13816 23435
rect 13848 23403 13888 23435
rect 13920 23403 13960 23435
rect 13992 23403 14032 23435
rect 14064 23403 14104 23435
rect 14136 23403 14176 23435
rect 14208 23403 14248 23435
rect 14280 23403 14320 23435
rect 14352 23403 14392 23435
rect 14424 23403 14464 23435
rect 14496 23403 14536 23435
rect 14568 23403 14608 23435
rect 14640 23403 14680 23435
rect 14712 23403 14752 23435
rect 14784 23403 14824 23435
rect 14856 23403 14896 23435
rect 14928 23403 14968 23435
rect 15000 23403 15040 23435
rect 15072 23403 15112 23435
rect 15144 23403 15184 23435
rect 15216 23403 15256 23435
rect 15288 23403 15328 23435
rect 15360 23403 15400 23435
rect 15432 23403 15472 23435
rect 15504 23403 15544 23435
rect 15576 23403 15616 23435
rect 15648 23403 15688 23435
rect 15720 23403 15760 23435
rect 15792 23403 15832 23435
rect 15864 23403 15904 23435
rect 15936 23403 16000 23435
rect 0 23363 16000 23403
rect 0 23331 64 23363
rect 96 23331 136 23363
rect 168 23331 208 23363
rect 240 23331 280 23363
rect 312 23331 352 23363
rect 384 23331 424 23363
rect 456 23331 496 23363
rect 528 23331 568 23363
rect 600 23331 640 23363
rect 672 23331 712 23363
rect 744 23331 784 23363
rect 816 23331 856 23363
rect 888 23331 928 23363
rect 960 23331 1000 23363
rect 1032 23331 1072 23363
rect 1104 23331 1144 23363
rect 1176 23331 1216 23363
rect 1248 23331 1288 23363
rect 1320 23331 1360 23363
rect 1392 23331 1432 23363
rect 1464 23331 1504 23363
rect 1536 23331 1576 23363
rect 1608 23331 1648 23363
rect 1680 23331 1720 23363
rect 1752 23331 1792 23363
rect 1824 23331 1864 23363
rect 1896 23331 1936 23363
rect 1968 23331 2008 23363
rect 2040 23331 2080 23363
rect 2112 23331 2152 23363
rect 2184 23331 2224 23363
rect 2256 23331 2296 23363
rect 2328 23331 2368 23363
rect 2400 23331 2440 23363
rect 2472 23331 2512 23363
rect 2544 23331 2584 23363
rect 2616 23331 2656 23363
rect 2688 23331 2728 23363
rect 2760 23331 2800 23363
rect 2832 23331 2872 23363
rect 2904 23331 2944 23363
rect 2976 23331 3016 23363
rect 3048 23331 3088 23363
rect 3120 23331 3160 23363
rect 3192 23331 3232 23363
rect 3264 23331 3304 23363
rect 3336 23331 3376 23363
rect 3408 23331 3448 23363
rect 3480 23331 3520 23363
rect 3552 23331 3592 23363
rect 3624 23331 3664 23363
rect 3696 23331 3736 23363
rect 3768 23331 3808 23363
rect 3840 23331 3880 23363
rect 3912 23331 3952 23363
rect 3984 23331 4024 23363
rect 4056 23331 4096 23363
rect 4128 23331 4168 23363
rect 4200 23331 4240 23363
rect 4272 23331 4312 23363
rect 4344 23331 4384 23363
rect 4416 23331 4456 23363
rect 4488 23331 4528 23363
rect 4560 23331 4600 23363
rect 4632 23331 4672 23363
rect 4704 23331 4744 23363
rect 4776 23331 4816 23363
rect 4848 23331 4888 23363
rect 4920 23331 4960 23363
rect 4992 23331 5032 23363
rect 5064 23331 5104 23363
rect 5136 23331 5176 23363
rect 5208 23331 5248 23363
rect 5280 23331 5320 23363
rect 5352 23331 5392 23363
rect 5424 23331 5464 23363
rect 5496 23331 5536 23363
rect 5568 23331 5608 23363
rect 5640 23331 5680 23363
rect 5712 23331 5752 23363
rect 5784 23331 5824 23363
rect 5856 23331 5896 23363
rect 5928 23331 5968 23363
rect 6000 23331 6040 23363
rect 6072 23331 6112 23363
rect 6144 23331 6184 23363
rect 6216 23331 6256 23363
rect 6288 23331 6328 23363
rect 6360 23331 6400 23363
rect 6432 23331 6472 23363
rect 6504 23331 6544 23363
rect 6576 23331 6616 23363
rect 6648 23331 6688 23363
rect 6720 23331 6760 23363
rect 6792 23331 6832 23363
rect 6864 23331 6904 23363
rect 6936 23331 6976 23363
rect 7008 23331 7048 23363
rect 7080 23331 7120 23363
rect 7152 23331 7192 23363
rect 7224 23331 7264 23363
rect 7296 23331 7336 23363
rect 7368 23331 7408 23363
rect 7440 23331 7480 23363
rect 7512 23331 7552 23363
rect 7584 23331 7624 23363
rect 7656 23331 7696 23363
rect 7728 23331 7768 23363
rect 7800 23331 7840 23363
rect 7872 23331 7912 23363
rect 7944 23331 7984 23363
rect 8016 23331 8056 23363
rect 8088 23331 8128 23363
rect 8160 23331 8200 23363
rect 8232 23331 8272 23363
rect 8304 23331 8344 23363
rect 8376 23331 8416 23363
rect 8448 23331 8488 23363
rect 8520 23331 8560 23363
rect 8592 23331 8632 23363
rect 8664 23331 8704 23363
rect 8736 23331 8776 23363
rect 8808 23331 8848 23363
rect 8880 23331 8920 23363
rect 8952 23331 8992 23363
rect 9024 23331 9064 23363
rect 9096 23331 9136 23363
rect 9168 23331 9208 23363
rect 9240 23331 9280 23363
rect 9312 23331 9352 23363
rect 9384 23331 9424 23363
rect 9456 23331 9496 23363
rect 9528 23331 9568 23363
rect 9600 23331 9640 23363
rect 9672 23331 9712 23363
rect 9744 23331 9784 23363
rect 9816 23331 9856 23363
rect 9888 23331 9928 23363
rect 9960 23331 10000 23363
rect 10032 23331 10072 23363
rect 10104 23331 10144 23363
rect 10176 23331 10216 23363
rect 10248 23331 10288 23363
rect 10320 23331 10360 23363
rect 10392 23331 10432 23363
rect 10464 23331 10504 23363
rect 10536 23331 10576 23363
rect 10608 23331 10648 23363
rect 10680 23331 10720 23363
rect 10752 23331 10792 23363
rect 10824 23331 10864 23363
rect 10896 23331 10936 23363
rect 10968 23331 11008 23363
rect 11040 23331 11080 23363
rect 11112 23331 11152 23363
rect 11184 23331 11224 23363
rect 11256 23331 11296 23363
rect 11328 23331 11368 23363
rect 11400 23331 11440 23363
rect 11472 23331 11512 23363
rect 11544 23331 11584 23363
rect 11616 23331 11656 23363
rect 11688 23331 11728 23363
rect 11760 23331 11800 23363
rect 11832 23331 11872 23363
rect 11904 23331 11944 23363
rect 11976 23331 12016 23363
rect 12048 23331 12088 23363
rect 12120 23331 12160 23363
rect 12192 23331 12232 23363
rect 12264 23331 12304 23363
rect 12336 23331 12376 23363
rect 12408 23331 12448 23363
rect 12480 23331 12520 23363
rect 12552 23331 12592 23363
rect 12624 23331 12664 23363
rect 12696 23331 12736 23363
rect 12768 23331 12808 23363
rect 12840 23331 12880 23363
rect 12912 23331 12952 23363
rect 12984 23331 13024 23363
rect 13056 23331 13096 23363
rect 13128 23331 13168 23363
rect 13200 23331 13240 23363
rect 13272 23331 13312 23363
rect 13344 23331 13384 23363
rect 13416 23331 13456 23363
rect 13488 23331 13528 23363
rect 13560 23331 13600 23363
rect 13632 23331 13672 23363
rect 13704 23331 13744 23363
rect 13776 23331 13816 23363
rect 13848 23331 13888 23363
rect 13920 23331 13960 23363
rect 13992 23331 14032 23363
rect 14064 23331 14104 23363
rect 14136 23331 14176 23363
rect 14208 23331 14248 23363
rect 14280 23331 14320 23363
rect 14352 23331 14392 23363
rect 14424 23331 14464 23363
rect 14496 23331 14536 23363
rect 14568 23331 14608 23363
rect 14640 23331 14680 23363
rect 14712 23331 14752 23363
rect 14784 23331 14824 23363
rect 14856 23331 14896 23363
rect 14928 23331 14968 23363
rect 15000 23331 15040 23363
rect 15072 23331 15112 23363
rect 15144 23331 15184 23363
rect 15216 23331 15256 23363
rect 15288 23331 15328 23363
rect 15360 23331 15400 23363
rect 15432 23331 15472 23363
rect 15504 23331 15544 23363
rect 15576 23331 15616 23363
rect 15648 23331 15688 23363
rect 15720 23331 15760 23363
rect 15792 23331 15832 23363
rect 15864 23331 15904 23363
rect 15936 23331 16000 23363
rect 0 23291 16000 23331
rect 0 23259 64 23291
rect 96 23259 136 23291
rect 168 23259 208 23291
rect 240 23259 280 23291
rect 312 23259 352 23291
rect 384 23259 424 23291
rect 456 23259 496 23291
rect 528 23259 568 23291
rect 600 23259 640 23291
rect 672 23259 712 23291
rect 744 23259 784 23291
rect 816 23259 856 23291
rect 888 23259 928 23291
rect 960 23259 1000 23291
rect 1032 23259 1072 23291
rect 1104 23259 1144 23291
rect 1176 23259 1216 23291
rect 1248 23259 1288 23291
rect 1320 23259 1360 23291
rect 1392 23259 1432 23291
rect 1464 23259 1504 23291
rect 1536 23259 1576 23291
rect 1608 23259 1648 23291
rect 1680 23259 1720 23291
rect 1752 23259 1792 23291
rect 1824 23259 1864 23291
rect 1896 23259 1936 23291
rect 1968 23259 2008 23291
rect 2040 23259 2080 23291
rect 2112 23259 2152 23291
rect 2184 23259 2224 23291
rect 2256 23259 2296 23291
rect 2328 23259 2368 23291
rect 2400 23259 2440 23291
rect 2472 23259 2512 23291
rect 2544 23259 2584 23291
rect 2616 23259 2656 23291
rect 2688 23259 2728 23291
rect 2760 23259 2800 23291
rect 2832 23259 2872 23291
rect 2904 23259 2944 23291
rect 2976 23259 3016 23291
rect 3048 23259 3088 23291
rect 3120 23259 3160 23291
rect 3192 23259 3232 23291
rect 3264 23259 3304 23291
rect 3336 23259 3376 23291
rect 3408 23259 3448 23291
rect 3480 23259 3520 23291
rect 3552 23259 3592 23291
rect 3624 23259 3664 23291
rect 3696 23259 3736 23291
rect 3768 23259 3808 23291
rect 3840 23259 3880 23291
rect 3912 23259 3952 23291
rect 3984 23259 4024 23291
rect 4056 23259 4096 23291
rect 4128 23259 4168 23291
rect 4200 23259 4240 23291
rect 4272 23259 4312 23291
rect 4344 23259 4384 23291
rect 4416 23259 4456 23291
rect 4488 23259 4528 23291
rect 4560 23259 4600 23291
rect 4632 23259 4672 23291
rect 4704 23259 4744 23291
rect 4776 23259 4816 23291
rect 4848 23259 4888 23291
rect 4920 23259 4960 23291
rect 4992 23259 5032 23291
rect 5064 23259 5104 23291
rect 5136 23259 5176 23291
rect 5208 23259 5248 23291
rect 5280 23259 5320 23291
rect 5352 23259 5392 23291
rect 5424 23259 5464 23291
rect 5496 23259 5536 23291
rect 5568 23259 5608 23291
rect 5640 23259 5680 23291
rect 5712 23259 5752 23291
rect 5784 23259 5824 23291
rect 5856 23259 5896 23291
rect 5928 23259 5968 23291
rect 6000 23259 6040 23291
rect 6072 23259 6112 23291
rect 6144 23259 6184 23291
rect 6216 23259 6256 23291
rect 6288 23259 6328 23291
rect 6360 23259 6400 23291
rect 6432 23259 6472 23291
rect 6504 23259 6544 23291
rect 6576 23259 6616 23291
rect 6648 23259 6688 23291
rect 6720 23259 6760 23291
rect 6792 23259 6832 23291
rect 6864 23259 6904 23291
rect 6936 23259 6976 23291
rect 7008 23259 7048 23291
rect 7080 23259 7120 23291
rect 7152 23259 7192 23291
rect 7224 23259 7264 23291
rect 7296 23259 7336 23291
rect 7368 23259 7408 23291
rect 7440 23259 7480 23291
rect 7512 23259 7552 23291
rect 7584 23259 7624 23291
rect 7656 23259 7696 23291
rect 7728 23259 7768 23291
rect 7800 23259 7840 23291
rect 7872 23259 7912 23291
rect 7944 23259 7984 23291
rect 8016 23259 8056 23291
rect 8088 23259 8128 23291
rect 8160 23259 8200 23291
rect 8232 23259 8272 23291
rect 8304 23259 8344 23291
rect 8376 23259 8416 23291
rect 8448 23259 8488 23291
rect 8520 23259 8560 23291
rect 8592 23259 8632 23291
rect 8664 23259 8704 23291
rect 8736 23259 8776 23291
rect 8808 23259 8848 23291
rect 8880 23259 8920 23291
rect 8952 23259 8992 23291
rect 9024 23259 9064 23291
rect 9096 23259 9136 23291
rect 9168 23259 9208 23291
rect 9240 23259 9280 23291
rect 9312 23259 9352 23291
rect 9384 23259 9424 23291
rect 9456 23259 9496 23291
rect 9528 23259 9568 23291
rect 9600 23259 9640 23291
rect 9672 23259 9712 23291
rect 9744 23259 9784 23291
rect 9816 23259 9856 23291
rect 9888 23259 9928 23291
rect 9960 23259 10000 23291
rect 10032 23259 10072 23291
rect 10104 23259 10144 23291
rect 10176 23259 10216 23291
rect 10248 23259 10288 23291
rect 10320 23259 10360 23291
rect 10392 23259 10432 23291
rect 10464 23259 10504 23291
rect 10536 23259 10576 23291
rect 10608 23259 10648 23291
rect 10680 23259 10720 23291
rect 10752 23259 10792 23291
rect 10824 23259 10864 23291
rect 10896 23259 10936 23291
rect 10968 23259 11008 23291
rect 11040 23259 11080 23291
rect 11112 23259 11152 23291
rect 11184 23259 11224 23291
rect 11256 23259 11296 23291
rect 11328 23259 11368 23291
rect 11400 23259 11440 23291
rect 11472 23259 11512 23291
rect 11544 23259 11584 23291
rect 11616 23259 11656 23291
rect 11688 23259 11728 23291
rect 11760 23259 11800 23291
rect 11832 23259 11872 23291
rect 11904 23259 11944 23291
rect 11976 23259 12016 23291
rect 12048 23259 12088 23291
rect 12120 23259 12160 23291
rect 12192 23259 12232 23291
rect 12264 23259 12304 23291
rect 12336 23259 12376 23291
rect 12408 23259 12448 23291
rect 12480 23259 12520 23291
rect 12552 23259 12592 23291
rect 12624 23259 12664 23291
rect 12696 23259 12736 23291
rect 12768 23259 12808 23291
rect 12840 23259 12880 23291
rect 12912 23259 12952 23291
rect 12984 23259 13024 23291
rect 13056 23259 13096 23291
rect 13128 23259 13168 23291
rect 13200 23259 13240 23291
rect 13272 23259 13312 23291
rect 13344 23259 13384 23291
rect 13416 23259 13456 23291
rect 13488 23259 13528 23291
rect 13560 23259 13600 23291
rect 13632 23259 13672 23291
rect 13704 23259 13744 23291
rect 13776 23259 13816 23291
rect 13848 23259 13888 23291
rect 13920 23259 13960 23291
rect 13992 23259 14032 23291
rect 14064 23259 14104 23291
rect 14136 23259 14176 23291
rect 14208 23259 14248 23291
rect 14280 23259 14320 23291
rect 14352 23259 14392 23291
rect 14424 23259 14464 23291
rect 14496 23259 14536 23291
rect 14568 23259 14608 23291
rect 14640 23259 14680 23291
rect 14712 23259 14752 23291
rect 14784 23259 14824 23291
rect 14856 23259 14896 23291
rect 14928 23259 14968 23291
rect 15000 23259 15040 23291
rect 15072 23259 15112 23291
rect 15144 23259 15184 23291
rect 15216 23259 15256 23291
rect 15288 23259 15328 23291
rect 15360 23259 15400 23291
rect 15432 23259 15472 23291
rect 15504 23259 15544 23291
rect 15576 23259 15616 23291
rect 15648 23259 15688 23291
rect 15720 23259 15760 23291
rect 15792 23259 15832 23291
rect 15864 23259 15904 23291
rect 15936 23259 16000 23291
rect 0 23219 16000 23259
rect 0 23187 64 23219
rect 96 23187 136 23219
rect 168 23187 208 23219
rect 240 23187 280 23219
rect 312 23187 352 23219
rect 384 23187 424 23219
rect 456 23187 496 23219
rect 528 23187 568 23219
rect 600 23187 640 23219
rect 672 23187 712 23219
rect 744 23187 784 23219
rect 816 23187 856 23219
rect 888 23187 928 23219
rect 960 23187 1000 23219
rect 1032 23187 1072 23219
rect 1104 23187 1144 23219
rect 1176 23187 1216 23219
rect 1248 23187 1288 23219
rect 1320 23187 1360 23219
rect 1392 23187 1432 23219
rect 1464 23187 1504 23219
rect 1536 23187 1576 23219
rect 1608 23187 1648 23219
rect 1680 23187 1720 23219
rect 1752 23187 1792 23219
rect 1824 23187 1864 23219
rect 1896 23187 1936 23219
rect 1968 23187 2008 23219
rect 2040 23187 2080 23219
rect 2112 23187 2152 23219
rect 2184 23187 2224 23219
rect 2256 23187 2296 23219
rect 2328 23187 2368 23219
rect 2400 23187 2440 23219
rect 2472 23187 2512 23219
rect 2544 23187 2584 23219
rect 2616 23187 2656 23219
rect 2688 23187 2728 23219
rect 2760 23187 2800 23219
rect 2832 23187 2872 23219
rect 2904 23187 2944 23219
rect 2976 23187 3016 23219
rect 3048 23187 3088 23219
rect 3120 23187 3160 23219
rect 3192 23187 3232 23219
rect 3264 23187 3304 23219
rect 3336 23187 3376 23219
rect 3408 23187 3448 23219
rect 3480 23187 3520 23219
rect 3552 23187 3592 23219
rect 3624 23187 3664 23219
rect 3696 23187 3736 23219
rect 3768 23187 3808 23219
rect 3840 23187 3880 23219
rect 3912 23187 3952 23219
rect 3984 23187 4024 23219
rect 4056 23187 4096 23219
rect 4128 23187 4168 23219
rect 4200 23187 4240 23219
rect 4272 23187 4312 23219
rect 4344 23187 4384 23219
rect 4416 23187 4456 23219
rect 4488 23187 4528 23219
rect 4560 23187 4600 23219
rect 4632 23187 4672 23219
rect 4704 23187 4744 23219
rect 4776 23187 4816 23219
rect 4848 23187 4888 23219
rect 4920 23187 4960 23219
rect 4992 23187 5032 23219
rect 5064 23187 5104 23219
rect 5136 23187 5176 23219
rect 5208 23187 5248 23219
rect 5280 23187 5320 23219
rect 5352 23187 5392 23219
rect 5424 23187 5464 23219
rect 5496 23187 5536 23219
rect 5568 23187 5608 23219
rect 5640 23187 5680 23219
rect 5712 23187 5752 23219
rect 5784 23187 5824 23219
rect 5856 23187 5896 23219
rect 5928 23187 5968 23219
rect 6000 23187 6040 23219
rect 6072 23187 6112 23219
rect 6144 23187 6184 23219
rect 6216 23187 6256 23219
rect 6288 23187 6328 23219
rect 6360 23187 6400 23219
rect 6432 23187 6472 23219
rect 6504 23187 6544 23219
rect 6576 23187 6616 23219
rect 6648 23187 6688 23219
rect 6720 23187 6760 23219
rect 6792 23187 6832 23219
rect 6864 23187 6904 23219
rect 6936 23187 6976 23219
rect 7008 23187 7048 23219
rect 7080 23187 7120 23219
rect 7152 23187 7192 23219
rect 7224 23187 7264 23219
rect 7296 23187 7336 23219
rect 7368 23187 7408 23219
rect 7440 23187 7480 23219
rect 7512 23187 7552 23219
rect 7584 23187 7624 23219
rect 7656 23187 7696 23219
rect 7728 23187 7768 23219
rect 7800 23187 7840 23219
rect 7872 23187 7912 23219
rect 7944 23187 7984 23219
rect 8016 23187 8056 23219
rect 8088 23187 8128 23219
rect 8160 23187 8200 23219
rect 8232 23187 8272 23219
rect 8304 23187 8344 23219
rect 8376 23187 8416 23219
rect 8448 23187 8488 23219
rect 8520 23187 8560 23219
rect 8592 23187 8632 23219
rect 8664 23187 8704 23219
rect 8736 23187 8776 23219
rect 8808 23187 8848 23219
rect 8880 23187 8920 23219
rect 8952 23187 8992 23219
rect 9024 23187 9064 23219
rect 9096 23187 9136 23219
rect 9168 23187 9208 23219
rect 9240 23187 9280 23219
rect 9312 23187 9352 23219
rect 9384 23187 9424 23219
rect 9456 23187 9496 23219
rect 9528 23187 9568 23219
rect 9600 23187 9640 23219
rect 9672 23187 9712 23219
rect 9744 23187 9784 23219
rect 9816 23187 9856 23219
rect 9888 23187 9928 23219
rect 9960 23187 10000 23219
rect 10032 23187 10072 23219
rect 10104 23187 10144 23219
rect 10176 23187 10216 23219
rect 10248 23187 10288 23219
rect 10320 23187 10360 23219
rect 10392 23187 10432 23219
rect 10464 23187 10504 23219
rect 10536 23187 10576 23219
rect 10608 23187 10648 23219
rect 10680 23187 10720 23219
rect 10752 23187 10792 23219
rect 10824 23187 10864 23219
rect 10896 23187 10936 23219
rect 10968 23187 11008 23219
rect 11040 23187 11080 23219
rect 11112 23187 11152 23219
rect 11184 23187 11224 23219
rect 11256 23187 11296 23219
rect 11328 23187 11368 23219
rect 11400 23187 11440 23219
rect 11472 23187 11512 23219
rect 11544 23187 11584 23219
rect 11616 23187 11656 23219
rect 11688 23187 11728 23219
rect 11760 23187 11800 23219
rect 11832 23187 11872 23219
rect 11904 23187 11944 23219
rect 11976 23187 12016 23219
rect 12048 23187 12088 23219
rect 12120 23187 12160 23219
rect 12192 23187 12232 23219
rect 12264 23187 12304 23219
rect 12336 23187 12376 23219
rect 12408 23187 12448 23219
rect 12480 23187 12520 23219
rect 12552 23187 12592 23219
rect 12624 23187 12664 23219
rect 12696 23187 12736 23219
rect 12768 23187 12808 23219
rect 12840 23187 12880 23219
rect 12912 23187 12952 23219
rect 12984 23187 13024 23219
rect 13056 23187 13096 23219
rect 13128 23187 13168 23219
rect 13200 23187 13240 23219
rect 13272 23187 13312 23219
rect 13344 23187 13384 23219
rect 13416 23187 13456 23219
rect 13488 23187 13528 23219
rect 13560 23187 13600 23219
rect 13632 23187 13672 23219
rect 13704 23187 13744 23219
rect 13776 23187 13816 23219
rect 13848 23187 13888 23219
rect 13920 23187 13960 23219
rect 13992 23187 14032 23219
rect 14064 23187 14104 23219
rect 14136 23187 14176 23219
rect 14208 23187 14248 23219
rect 14280 23187 14320 23219
rect 14352 23187 14392 23219
rect 14424 23187 14464 23219
rect 14496 23187 14536 23219
rect 14568 23187 14608 23219
rect 14640 23187 14680 23219
rect 14712 23187 14752 23219
rect 14784 23187 14824 23219
rect 14856 23187 14896 23219
rect 14928 23187 14968 23219
rect 15000 23187 15040 23219
rect 15072 23187 15112 23219
rect 15144 23187 15184 23219
rect 15216 23187 15256 23219
rect 15288 23187 15328 23219
rect 15360 23187 15400 23219
rect 15432 23187 15472 23219
rect 15504 23187 15544 23219
rect 15576 23187 15616 23219
rect 15648 23187 15688 23219
rect 15720 23187 15760 23219
rect 15792 23187 15832 23219
rect 15864 23187 15904 23219
rect 15936 23187 16000 23219
rect 0 23124 16000 23187
rect 0 23121 68 23124
rect 0 23089 18 23121
rect 50 23089 68 23121
rect 0 23053 68 23089
rect 0 23021 18 23053
rect 50 23021 68 23053
rect 0 22984 68 23021
rect 0 22952 18 22984
rect 50 22952 68 22984
rect 0 22915 68 22952
rect 0 22883 18 22915
rect 50 22883 68 22915
rect 0 22846 68 22883
rect 0 22814 18 22846
rect 50 22814 68 22846
rect 0 22777 68 22814
rect 0 22745 18 22777
rect 50 22745 68 22777
rect 0 22708 68 22745
rect 0 22676 18 22708
rect 50 22676 68 22708
rect 0 22639 68 22676
rect 0 22607 18 22639
rect 50 22607 68 22639
rect 0 22570 68 22607
rect 0 22538 18 22570
rect 50 22538 68 22570
rect 0 22501 68 22538
rect 0 22469 18 22501
rect 50 22469 68 22501
rect 0 22432 68 22469
rect 0 22400 18 22432
rect 50 22400 68 22432
rect 0 22363 68 22400
rect 0 22331 18 22363
rect 50 22331 68 22363
rect 0 22294 68 22331
rect 0 22262 18 22294
rect 50 22262 68 22294
rect 0 22225 68 22262
rect 0 22193 18 22225
rect 50 22193 68 22225
rect 0 22156 68 22193
rect 0 22124 18 22156
rect 50 22124 68 22156
rect 0 22087 68 22124
rect 0 22055 18 22087
rect 50 22055 68 22087
rect 0 22018 68 22055
rect 0 21986 18 22018
rect 50 21986 68 22018
rect 0 21949 68 21986
rect 0 21917 18 21949
rect 50 21917 68 21949
rect 0 21880 68 21917
rect 0 21848 18 21880
rect 50 21848 68 21880
rect 0 21811 68 21848
rect 0 21779 18 21811
rect 50 21779 68 21811
rect 0 21742 68 21779
rect 0 21710 18 21742
rect 50 21710 68 21742
rect 0 21673 68 21710
rect 0 21641 18 21673
rect 50 21641 68 21673
rect 0 21604 68 21641
rect 0 21572 18 21604
rect 50 21572 68 21604
rect 0 21535 68 21572
rect 0 21503 18 21535
rect 50 21503 68 21535
rect 0 21466 68 21503
rect 0 21434 18 21466
rect 50 21434 68 21466
rect 0 21397 68 21434
rect 0 21365 18 21397
rect 50 21365 68 21397
rect 0 21328 68 21365
rect 0 21296 18 21328
rect 50 21296 68 21328
rect 0 21259 68 21296
rect 0 21227 18 21259
rect 50 21227 68 21259
rect 0 21190 68 21227
rect 0 21158 18 21190
rect 50 21158 68 21190
rect 0 21121 68 21158
rect 0 21089 18 21121
rect 50 21089 68 21121
rect 0 21052 68 21089
rect 0 21020 18 21052
rect 50 21020 68 21052
rect 0 20983 68 21020
rect 0 20951 18 20983
rect 50 20951 68 20983
rect 0 20914 68 20951
rect 0 20882 18 20914
rect 50 20882 68 20914
rect 0 20845 68 20882
rect 0 20813 18 20845
rect 50 20813 68 20845
rect 0 20776 68 20813
rect 0 20744 18 20776
rect 50 20744 68 20776
rect 0 20707 68 20744
rect 0 20675 18 20707
rect 50 20675 68 20707
rect 0 20638 68 20675
rect 0 20606 18 20638
rect 50 20606 68 20638
rect 0 20569 68 20606
rect 0 20537 18 20569
rect 50 20537 68 20569
rect 0 20500 68 20537
rect 0 20468 18 20500
rect 50 20468 68 20500
rect 0 20431 68 20468
rect 0 20399 18 20431
rect 50 20399 68 20431
rect 0 20362 68 20399
rect 0 20330 18 20362
rect 50 20330 68 20362
rect 0 20293 68 20330
rect 0 20261 18 20293
rect 50 20261 68 20293
rect 0 20224 68 20261
rect 0 20192 18 20224
rect 50 20192 68 20224
rect 0 20155 68 20192
rect 0 20123 18 20155
rect 50 20123 68 20155
rect 0 20086 68 20123
rect 0 20054 18 20086
rect 50 20054 68 20086
rect 15934 23110 16000 23124
rect 15934 23078 15951 23110
rect 15983 23078 16000 23110
rect 15934 23042 16000 23078
rect 15934 23010 15951 23042
rect 15983 23010 16000 23042
rect 15934 22974 16000 23010
rect 15934 22942 15951 22974
rect 15983 22942 16000 22974
rect 15934 22906 16000 22942
rect 15934 22874 15951 22906
rect 15983 22874 16000 22906
rect 15934 22838 16000 22874
rect 15934 22806 15951 22838
rect 15983 22806 16000 22838
rect 15934 22770 16000 22806
rect 15934 22738 15951 22770
rect 15983 22738 16000 22770
rect 15934 22702 16000 22738
rect 15934 22670 15951 22702
rect 15983 22670 16000 22702
rect 15934 22634 16000 22670
rect 15934 22602 15951 22634
rect 15983 22602 16000 22634
rect 15934 22566 16000 22602
rect 15934 22534 15951 22566
rect 15983 22534 16000 22566
rect 15934 22498 16000 22534
rect 15934 22466 15951 22498
rect 15983 22466 16000 22498
rect 15934 22430 16000 22466
rect 15934 22398 15951 22430
rect 15983 22398 16000 22430
rect 15934 22362 16000 22398
rect 15934 22330 15951 22362
rect 15983 22330 16000 22362
rect 15934 22294 16000 22330
rect 15934 22262 15951 22294
rect 15983 22262 16000 22294
rect 15934 22226 16000 22262
rect 15934 22194 15951 22226
rect 15983 22194 16000 22226
rect 15934 22158 16000 22194
rect 15934 22126 15951 22158
rect 15983 22126 16000 22158
rect 15934 22090 16000 22126
rect 15934 22058 15951 22090
rect 15983 22058 16000 22090
rect 15934 22022 16000 22058
rect 15934 21990 15951 22022
rect 15983 21990 16000 22022
rect 15934 21954 16000 21990
rect 15934 21922 15951 21954
rect 15983 21922 16000 21954
rect 15934 21886 16000 21922
rect 15934 21854 15951 21886
rect 15983 21854 16000 21886
rect 15934 21818 16000 21854
rect 15934 21786 15951 21818
rect 15983 21786 16000 21818
rect 15934 21750 16000 21786
rect 15934 21718 15951 21750
rect 15983 21718 16000 21750
rect 15934 21682 16000 21718
rect 15934 21650 15951 21682
rect 15983 21650 16000 21682
rect 15934 21614 16000 21650
rect 15934 21582 15951 21614
rect 15983 21582 16000 21614
rect 15934 21546 16000 21582
rect 15934 21514 15951 21546
rect 15983 21514 16000 21546
rect 15934 21478 16000 21514
rect 15934 21446 15951 21478
rect 15983 21446 16000 21478
rect 15934 21410 16000 21446
rect 15934 21378 15951 21410
rect 15983 21378 16000 21410
rect 15934 21342 16000 21378
rect 15934 21310 15951 21342
rect 15983 21310 16000 21342
rect 15934 21274 16000 21310
rect 15934 21242 15951 21274
rect 15983 21242 16000 21274
rect 15934 21206 16000 21242
rect 15934 21174 15951 21206
rect 15983 21174 16000 21206
rect 15934 21138 16000 21174
rect 15934 21106 15951 21138
rect 15983 21106 16000 21138
rect 15934 21070 16000 21106
rect 15934 21038 15951 21070
rect 15983 21038 16000 21070
rect 15934 21002 16000 21038
rect 15934 20970 15951 21002
rect 15983 20970 16000 21002
rect 15934 20934 16000 20970
rect 15934 20902 15951 20934
rect 15983 20902 16000 20934
rect 15934 20866 16000 20902
rect 15934 20834 15951 20866
rect 15983 20834 16000 20866
rect 15934 20798 16000 20834
rect 15934 20766 15951 20798
rect 15983 20766 16000 20798
rect 15934 20730 16000 20766
rect 15934 20698 15951 20730
rect 15983 20698 16000 20730
rect 15934 20662 16000 20698
rect 15934 20630 15951 20662
rect 15983 20630 16000 20662
rect 15934 20594 16000 20630
rect 15934 20562 15951 20594
rect 15983 20562 16000 20594
rect 15934 20526 16000 20562
rect 15934 20494 15951 20526
rect 15983 20494 16000 20526
rect 15934 20458 16000 20494
rect 15934 20426 15951 20458
rect 15983 20426 16000 20458
rect 15934 20390 16000 20426
rect 15934 20358 15951 20390
rect 15983 20358 16000 20390
rect 15934 20322 16000 20358
rect 15934 20290 15951 20322
rect 15983 20290 16000 20322
rect 15934 20254 16000 20290
rect 15934 20222 15951 20254
rect 15983 20222 16000 20254
rect 15934 20186 16000 20222
rect 15934 20154 15951 20186
rect 15983 20154 16000 20186
rect 15934 20118 16000 20154
rect 15934 20086 15951 20118
rect 15983 20086 16000 20118
rect 0 20017 68 20054
rect 3264 20071 12736 20080
rect 3264 20031 3306 20071
rect 12694 20031 12736 20071
rect 3264 20022 12736 20031
rect 15934 20050 16000 20086
rect 0 19985 18 20017
rect 50 19985 68 20017
rect 0 19948 68 19985
rect 0 19916 18 19948
rect 50 19916 68 19948
rect 0 19879 68 19916
rect 0 19847 18 19879
rect 50 19847 68 19879
rect 0 19810 68 19847
rect 0 19778 18 19810
rect 50 19778 68 19810
rect 0 19741 68 19778
rect 0 19709 18 19741
rect 50 19709 68 19741
rect 0 19672 68 19709
rect 0 19640 18 19672
rect 50 19640 68 19672
rect 0 19603 68 19640
rect 0 19571 18 19603
rect 50 19571 68 19603
rect 0 19534 68 19571
rect 0 19502 18 19534
rect 50 19502 68 19534
rect 0 19465 68 19502
rect 0 19433 18 19465
rect 50 19433 68 19465
rect 0 19396 68 19433
rect 0 19364 18 19396
rect 50 19364 68 19396
rect 0 19327 68 19364
rect 0 19295 18 19327
rect 50 19295 68 19327
rect 0 19258 68 19295
rect 0 19226 18 19258
rect 50 19226 68 19258
rect 0 19189 68 19226
rect 0 19157 18 19189
rect 50 19157 68 19189
rect 0 19120 68 19157
rect 0 19088 18 19120
rect 50 19088 68 19120
rect 0 19051 68 19088
rect 0 19019 18 19051
rect 50 19019 68 19051
rect 0 18982 68 19019
rect 0 18950 18 18982
rect 50 18950 68 18982
rect 0 18913 68 18950
rect 0 18881 18 18913
rect 50 18881 68 18913
rect 0 18844 68 18881
rect 0 18812 18 18844
rect 50 18812 68 18844
rect 0 18775 68 18812
rect 0 18743 18 18775
rect 50 18743 68 18775
rect 0 18706 68 18743
rect 0 18674 18 18706
rect 50 18674 68 18706
rect 0 18637 68 18674
rect 0 18605 18 18637
rect 50 18605 68 18637
rect 0 18568 68 18605
rect 0 18536 18 18568
rect 50 18536 68 18568
rect 0 18499 68 18536
rect 0 18467 18 18499
rect 50 18467 68 18499
rect 0 18430 68 18467
rect 0 18398 18 18430
rect 50 18398 68 18430
rect 0 18361 68 18398
rect 0 18329 18 18361
rect 50 18329 68 18361
rect 0 18292 68 18329
rect 0 18260 18 18292
rect 50 18260 68 18292
rect 0 18223 68 18260
rect 0 18191 18 18223
rect 50 18191 68 18223
rect 0 18154 68 18191
rect 0 18122 18 18154
rect 50 18122 68 18154
rect 0 18085 68 18122
rect 0 18053 18 18085
rect 50 18053 68 18085
rect 0 18016 68 18053
rect 0 17984 18 18016
rect 50 17984 68 18016
rect 0 17947 68 17984
rect 0 17915 18 17947
rect 50 17915 68 17947
rect 0 17878 68 17915
rect 0 17846 18 17878
rect 50 17846 68 17878
rect 0 17809 68 17846
rect 0 17777 18 17809
rect 50 17777 68 17809
rect 0 17740 68 17777
rect 0 17708 18 17740
rect 50 17708 68 17740
rect 0 17671 68 17708
rect 0 17639 18 17671
rect 50 17639 68 17671
rect 0 17602 68 17639
rect 0 17570 18 17602
rect 50 17570 68 17602
rect 0 17534 68 17570
rect 0 17502 18 17534
rect 50 17502 68 17534
rect 0 13000 68 17502
rect 15934 20018 15951 20050
rect 15983 20018 16000 20050
rect 15934 19982 16000 20018
rect 15934 19950 15951 19982
rect 15983 19950 16000 19982
rect 15934 19914 16000 19950
rect 15934 19882 15951 19914
rect 15983 19882 16000 19914
rect 15934 19846 16000 19882
rect 15934 19814 15951 19846
rect 15983 19814 16000 19846
rect 15934 19778 16000 19814
rect 15934 19746 15951 19778
rect 15983 19746 16000 19778
rect 15934 19710 16000 19746
rect 15934 19678 15951 19710
rect 15983 19678 16000 19710
rect 15934 19642 16000 19678
rect 15934 19610 15951 19642
rect 15983 19610 16000 19642
rect 15934 19574 16000 19610
rect 15934 19542 15951 19574
rect 15983 19542 16000 19574
rect 15934 19506 16000 19542
rect 15934 19474 15951 19506
rect 15983 19474 16000 19506
rect 15934 19438 16000 19474
rect 15934 19406 15951 19438
rect 15983 19406 16000 19438
rect 15934 19370 16000 19406
rect 15934 19338 15951 19370
rect 15983 19338 16000 19370
rect 15934 19302 16000 19338
rect 15934 19270 15951 19302
rect 15983 19270 16000 19302
rect 15934 19234 16000 19270
rect 15934 19202 15951 19234
rect 15983 19202 16000 19234
rect 15934 19166 16000 19202
rect 15934 19134 15951 19166
rect 15983 19134 16000 19166
rect 15934 19098 16000 19134
rect 15934 19066 15951 19098
rect 15983 19066 16000 19098
rect 15934 19030 16000 19066
rect 15934 18998 15951 19030
rect 15983 18998 16000 19030
rect 15934 18962 16000 18998
rect 15934 18930 15951 18962
rect 15983 18930 16000 18962
rect 15934 18894 16000 18930
rect 15934 18862 15951 18894
rect 15983 18862 16000 18894
rect 15934 18826 16000 18862
rect 15934 18794 15951 18826
rect 15983 18794 16000 18826
rect 15934 18758 16000 18794
rect 15934 18726 15951 18758
rect 15983 18726 16000 18758
rect 15934 18690 16000 18726
rect 15934 18658 15951 18690
rect 15983 18658 16000 18690
rect 15934 18622 16000 18658
rect 15934 18590 15951 18622
rect 15983 18590 16000 18622
rect 15934 18554 16000 18590
rect 15934 18522 15951 18554
rect 15983 18522 16000 18554
rect 15934 18486 16000 18522
rect 15934 18454 15951 18486
rect 15983 18454 16000 18486
rect 15934 18418 16000 18454
rect 15934 18386 15951 18418
rect 15983 18386 16000 18418
rect 15934 18350 16000 18386
rect 15934 18318 15951 18350
rect 15983 18318 16000 18350
rect 15934 18282 16000 18318
rect 15934 18250 15951 18282
rect 15983 18250 16000 18282
rect 15934 18214 16000 18250
rect 15934 18182 15951 18214
rect 15983 18182 16000 18214
rect 15934 18146 16000 18182
rect 15934 18114 15951 18146
rect 15983 18114 16000 18146
rect 15934 18078 16000 18114
rect 15934 18046 15951 18078
rect 15983 18046 16000 18078
rect 15934 18010 16000 18046
rect 15934 17978 15951 18010
rect 15983 17978 16000 18010
rect 15934 17942 16000 17978
rect 15934 17910 15951 17942
rect 15983 17910 16000 17942
rect 15934 17874 16000 17910
rect 15934 17842 15951 17874
rect 15983 17842 16000 17874
rect 15934 17806 16000 17842
rect 15934 17774 15951 17806
rect 15983 17774 16000 17806
rect 15934 17738 16000 17774
rect 15934 17706 15951 17738
rect 15983 17706 16000 17738
rect 15934 17670 16000 17706
rect 15934 17638 15951 17670
rect 15983 17638 16000 17670
rect 15934 17602 16000 17638
rect 15934 17570 15951 17602
rect 15983 17570 16000 17602
rect 15934 17534 16000 17570
rect 15934 17502 15951 17534
rect 15983 17502 16000 17534
rect 15934 13000 16000 17502
rect 0 12690 16000 12708
rect 0 12658 28 12690
rect 60 12658 96 12690
rect 128 12658 164 12690
rect 196 12658 232 12690
rect 264 12658 300 12690
rect 332 12658 368 12690
rect 400 12658 436 12690
rect 468 12658 504 12690
rect 536 12658 572 12690
rect 604 12658 640 12690
rect 672 12658 708 12690
rect 740 12658 776 12690
rect 808 12658 844 12690
rect 876 12658 912 12690
rect 944 12658 980 12690
rect 1012 12658 1048 12690
rect 1080 12658 1116 12690
rect 1148 12658 1184 12690
rect 1216 12658 1252 12690
rect 1284 12658 1320 12690
rect 1352 12658 1388 12690
rect 1420 12658 1456 12690
rect 1488 12658 1524 12690
rect 1556 12658 1592 12690
rect 1624 12658 1660 12690
rect 1692 12658 1728 12690
rect 1760 12658 1796 12690
rect 1828 12658 1864 12690
rect 1896 12658 1932 12690
rect 1964 12658 2000 12690
rect 2032 12658 2068 12690
rect 2100 12658 2136 12690
rect 2168 12658 2204 12690
rect 2236 12658 2272 12690
rect 2304 12658 2340 12690
rect 2372 12658 2408 12690
rect 2440 12658 2476 12690
rect 2508 12658 2544 12690
rect 2576 12658 2612 12690
rect 2644 12658 2680 12690
rect 2712 12658 2748 12690
rect 2780 12658 2816 12690
rect 2848 12658 2884 12690
rect 2916 12658 2952 12690
rect 2984 12658 3020 12690
rect 3052 12658 3088 12690
rect 3120 12658 3156 12690
rect 3188 12658 3224 12690
rect 3256 12658 3292 12690
rect 3324 12658 3360 12690
rect 3392 12658 3428 12690
rect 3460 12658 3496 12690
rect 3528 12658 3564 12690
rect 3596 12658 3632 12690
rect 3664 12658 3700 12690
rect 3732 12658 3768 12690
rect 3800 12658 3836 12690
rect 3868 12658 3904 12690
rect 3936 12658 3972 12690
rect 4004 12658 4040 12690
rect 4072 12658 4108 12690
rect 4140 12658 4176 12690
rect 4208 12658 4244 12690
rect 4276 12658 4312 12690
rect 4344 12658 4380 12690
rect 4412 12658 4448 12690
rect 4480 12658 4516 12690
rect 4548 12658 4584 12690
rect 4616 12658 4652 12690
rect 4684 12658 4720 12690
rect 4752 12658 4788 12690
rect 4820 12658 4856 12690
rect 4888 12658 4924 12690
rect 4956 12658 4992 12690
rect 5024 12658 5060 12690
rect 5092 12658 5128 12690
rect 5160 12658 5196 12690
rect 5228 12658 5264 12690
rect 5296 12658 5332 12690
rect 5364 12658 5400 12690
rect 5432 12658 5468 12690
rect 5500 12658 5536 12690
rect 5568 12658 5604 12690
rect 5636 12658 5672 12690
rect 5704 12658 5740 12690
rect 5772 12658 5808 12690
rect 5840 12658 5876 12690
rect 5908 12658 5944 12690
rect 5976 12658 6012 12690
rect 6044 12658 6080 12690
rect 6112 12658 6148 12690
rect 6180 12658 6216 12690
rect 6248 12658 6284 12690
rect 6316 12658 6352 12690
rect 6384 12658 6420 12690
rect 6452 12658 6488 12690
rect 6520 12658 6556 12690
rect 6588 12658 6624 12690
rect 6656 12658 6692 12690
rect 6724 12658 6760 12690
rect 6792 12658 6828 12690
rect 6860 12658 6896 12690
rect 6928 12658 6964 12690
rect 6996 12658 7032 12690
rect 7064 12658 7100 12690
rect 7132 12658 7168 12690
rect 7200 12658 7236 12690
rect 7268 12658 7304 12690
rect 7336 12658 7372 12690
rect 7404 12658 7440 12690
rect 7472 12658 7508 12690
rect 7540 12658 7576 12690
rect 7608 12658 7644 12690
rect 7676 12658 7712 12690
rect 7744 12658 7780 12690
rect 7812 12658 7848 12690
rect 7880 12658 7916 12690
rect 7948 12658 7984 12690
rect 8016 12658 8052 12690
rect 8084 12658 8120 12690
rect 8152 12658 8188 12690
rect 8220 12658 8256 12690
rect 8288 12658 8324 12690
rect 8356 12658 8392 12690
rect 8424 12658 8460 12690
rect 8492 12658 8528 12690
rect 8560 12658 8596 12690
rect 8628 12658 8664 12690
rect 8696 12658 8732 12690
rect 8764 12658 8800 12690
rect 8832 12658 8868 12690
rect 8900 12658 8936 12690
rect 8968 12658 9004 12690
rect 9036 12658 9072 12690
rect 9104 12658 9140 12690
rect 9172 12658 9208 12690
rect 9240 12658 9276 12690
rect 9308 12658 9344 12690
rect 9376 12658 9412 12690
rect 9444 12658 9480 12690
rect 9512 12658 9548 12690
rect 9580 12658 9616 12690
rect 9648 12658 9684 12690
rect 9716 12658 9752 12690
rect 9784 12658 9820 12690
rect 9852 12658 9888 12690
rect 9920 12658 9956 12690
rect 9988 12658 10024 12690
rect 10056 12658 10092 12690
rect 10124 12658 10160 12690
rect 10192 12658 10228 12690
rect 10260 12658 10296 12690
rect 10328 12658 10364 12690
rect 10396 12658 10432 12690
rect 10464 12658 10500 12690
rect 10532 12658 10568 12690
rect 10600 12658 10636 12690
rect 10668 12658 10704 12690
rect 10736 12658 10772 12690
rect 10804 12658 10840 12690
rect 10872 12658 10908 12690
rect 10940 12658 10976 12690
rect 11008 12658 11044 12690
rect 11076 12658 11112 12690
rect 11144 12658 11180 12690
rect 11212 12658 11248 12690
rect 11280 12658 11316 12690
rect 11348 12658 11384 12690
rect 11416 12658 11452 12690
rect 11484 12658 11520 12690
rect 11552 12658 11588 12690
rect 11620 12658 11656 12690
rect 11688 12658 11724 12690
rect 11756 12658 11792 12690
rect 11824 12658 11860 12690
rect 11892 12658 11928 12690
rect 11960 12658 11996 12690
rect 12028 12658 12064 12690
rect 12096 12658 12132 12690
rect 12164 12658 12200 12690
rect 12232 12658 12268 12690
rect 12300 12658 12336 12690
rect 12368 12658 12404 12690
rect 12436 12658 12472 12690
rect 12504 12658 12540 12690
rect 12572 12658 12608 12690
rect 12640 12658 12676 12690
rect 12708 12658 12744 12690
rect 12776 12658 12812 12690
rect 12844 12658 12880 12690
rect 12912 12658 12948 12690
rect 12980 12658 13016 12690
rect 13048 12658 13084 12690
rect 13116 12658 13152 12690
rect 13184 12658 13220 12690
rect 13252 12658 13288 12690
rect 13320 12658 13356 12690
rect 13388 12658 13424 12690
rect 13456 12658 13492 12690
rect 13524 12658 13560 12690
rect 13592 12658 13628 12690
rect 13660 12658 13696 12690
rect 13728 12658 13764 12690
rect 13796 12658 13832 12690
rect 13864 12658 13900 12690
rect 13932 12658 13968 12690
rect 14000 12658 14036 12690
rect 14068 12658 14104 12690
rect 14136 12658 14172 12690
rect 14204 12658 14240 12690
rect 14272 12658 14308 12690
rect 14340 12658 14376 12690
rect 14408 12658 14444 12690
rect 14476 12658 14512 12690
rect 14544 12658 14580 12690
rect 14612 12658 14648 12690
rect 14680 12658 14716 12690
rect 14748 12658 14784 12690
rect 14816 12658 14852 12690
rect 14884 12658 14920 12690
rect 14952 12658 14988 12690
rect 15020 12658 15056 12690
rect 15088 12658 15124 12690
rect 15156 12658 15192 12690
rect 15224 12658 15260 12690
rect 15292 12658 15328 12690
rect 15360 12658 15396 12690
rect 15428 12658 15464 12690
rect 15496 12658 15532 12690
rect 15564 12658 15600 12690
rect 15632 12658 15668 12690
rect 15700 12658 15736 12690
rect 15768 12658 15804 12690
rect 15836 12658 15872 12690
rect 15904 12658 15940 12690
rect 15972 12658 16000 12690
rect 0 12640 16000 12658
rect 0 12574 68 12640
rect 0 12542 18 12574
rect 50 12542 68 12574
rect 15932 12574 16000 12640
rect 0 12506 68 12542
rect 0 12474 18 12506
rect 50 12474 68 12506
rect 0 12438 68 12474
rect 0 12406 18 12438
rect 50 12406 68 12438
rect 0 12370 68 12406
rect 0 12338 18 12370
rect 50 12338 68 12370
rect 0 12302 68 12338
rect 0 12270 18 12302
rect 50 12270 68 12302
rect 0 12234 68 12270
rect 0 12202 18 12234
rect 50 12202 68 12234
rect 0 12166 68 12202
rect 0 12134 18 12166
rect 50 12134 68 12166
rect 0 12098 68 12134
rect 0 12066 18 12098
rect 50 12066 68 12098
rect 0 12030 68 12066
rect 0 11998 18 12030
rect 50 11998 68 12030
rect 0 11962 68 11998
rect 0 11930 18 11962
rect 50 11930 68 11962
rect 0 11894 68 11930
rect 0 11862 18 11894
rect 50 11862 68 11894
rect 0 11826 68 11862
rect 0 11794 18 11826
rect 50 11794 68 11826
rect 0 11758 68 11794
rect 0 11726 18 11758
rect 50 11726 68 11758
rect 0 11690 68 11726
rect 0 11658 18 11690
rect 50 11658 68 11690
rect 0 11622 68 11658
rect 12041 12559 15406 12568
rect 12041 12519 12064 12559
rect 15384 12519 15406 12559
rect 12041 12510 15406 12519
rect 15932 12542 15950 12574
rect 15982 12542 16000 12574
rect 0 11590 18 11622
rect 50 11590 68 11622
rect 0 11554 68 11590
rect 3835 11618 3959 11627
rect 3835 11578 3836 11618
rect 3958 11578 3959 11618
rect 3835 11569 3959 11578
rect 12041 11566 12209 12510
rect 15932 12506 16000 12542
rect 15932 12474 15950 12506
rect 15982 12474 16000 12506
rect 15932 12438 16000 12474
rect 15932 12406 15950 12438
rect 15982 12406 16000 12438
rect 15932 12370 16000 12406
rect 15932 12338 15950 12370
rect 15982 12338 16000 12370
rect 15932 12302 16000 12338
rect 15932 12270 15950 12302
rect 15982 12270 16000 12302
rect 15932 12234 16000 12270
rect 15932 12202 15950 12234
rect 15982 12202 16000 12234
rect 15932 12166 16000 12202
rect 15932 12134 15950 12166
rect 15982 12134 16000 12166
rect 15932 12098 16000 12134
rect 15932 12066 15950 12098
rect 15982 12066 16000 12098
rect 15932 12030 16000 12066
rect 15932 11998 15950 12030
rect 15982 11998 16000 12030
rect 15932 11962 16000 11998
rect 15932 11930 15950 11962
rect 15982 11930 16000 11962
rect 15932 11894 16000 11930
rect 15932 11862 15950 11894
rect 15982 11862 16000 11894
rect 15932 11826 16000 11862
rect 15932 11794 15950 11826
rect 15982 11794 16000 11826
rect 15932 11758 16000 11794
rect 15932 11726 15950 11758
rect 15982 11726 16000 11758
rect 15932 11690 16000 11726
rect 15932 11658 15950 11690
rect 15982 11658 16000 11690
rect 15932 11622 16000 11658
rect 15932 11590 15950 11622
rect 15982 11590 16000 11622
rect 0 11522 18 11554
rect 50 11522 68 11554
rect 0 11486 68 11522
rect 0 11454 18 11486
rect 50 11454 68 11486
rect 0 11418 68 11454
rect 0 11386 18 11418
rect 50 11386 68 11418
rect 0 11350 68 11386
rect 0 11318 18 11350
rect 50 11318 68 11350
rect 0 11282 68 11318
rect 0 11250 18 11282
rect 50 11250 68 11282
rect 0 11214 68 11250
rect 0 11182 18 11214
rect 50 11182 68 11214
rect 0 11146 68 11182
rect 0 11114 18 11146
rect 50 11114 68 11146
rect 0 11078 68 11114
rect 0 11046 18 11078
rect 50 11046 68 11078
rect 0 11010 68 11046
rect 0 10978 18 11010
rect 50 10978 68 11010
rect 0 10942 68 10978
rect 0 10910 18 10942
rect 50 10910 68 10942
rect 0 10874 68 10910
rect 0 10842 18 10874
rect 50 10842 68 10874
rect 0 10806 68 10842
rect 0 10774 18 10806
rect 50 10774 68 10806
rect 0 10738 68 10774
rect 0 10706 18 10738
rect 50 10706 68 10738
rect 0 10670 68 10706
rect 0 10638 18 10670
rect 50 10638 68 10670
rect 0 10602 68 10638
rect 0 10570 18 10602
rect 50 10570 68 10602
rect 0 10534 68 10570
rect 0 10502 18 10534
rect 50 10502 68 10534
rect 0 10466 68 10502
rect 0 10434 18 10466
rect 50 10434 68 10466
rect 0 10398 68 10434
rect 0 10366 18 10398
rect 50 10366 68 10398
rect 0 10330 68 10366
rect 0 10298 18 10330
rect 50 10298 68 10330
rect 0 10262 68 10298
rect 0 10230 18 10262
rect 50 10230 68 10262
rect 0 10194 68 10230
rect 0 10162 18 10194
rect 50 10162 68 10194
rect 0 10126 68 10162
rect 0 10094 18 10126
rect 50 10094 68 10126
rect 0 10058 68 10094
rect 0 10026 18 10058
rect 50 10026 68 10058
rect 0 9990 68 10026
rect 0 9958 18 9990
rect 50 9958 68 9990
rect 0 9922 68 9958
rect 0 9890 18 9922
rect 50 9890 68 9922
rect 0 9854 68 9890
rect 0 9822 18 9854
rect 50 9822 68 9854
rect 0 9786 68 9822
rect 0 9754 18 9786
rect 50 9754 68 9786
rect 0 9718 68 9754
rect 0 9686 18 9718
rect 50 9686 68 9718
rect 0 9650 68 9686
rect 0 9618 18 9650
rect 50 9618 68 9650
rect 0 9582 68 9618
rect 0 9550 18 9582
rect 50 9550 68 9582
rect 0 9514 68 9550
rect 0 9482 18 9514
rect 50 9482 68 9514
rect 0 9446 68 9482
rect 0 9414 18 9446
rect 50 9414 68 9446
rect 0 9378 68 9414
rect 0 9346 18 9378
rect 50 9346 68 9378
rect 0 9310 68 9346
rect 0 9278 18 9310
rect 50 9278 68 9310
rect 0 9242 68 9278
rect 0 9210 18 9242
rect 50 9210 68 9242
rect 0 9174 68 9210
rect 0 9142 18 9174
rect 50 9142 68 9174
rect 0 9106 68 9142
rect 0 9074 18 9106
rect 50 9074 68 9106
rect 0 9038 68 9074
rect 0 9006 18 9038
rect 50 9006 68 9038
rect 0 8970 68 9006
rect 0 8938 18 8970
rect 50 8938 68 8970
rect 0 8902 68 8938
rect 0 8870 18 8902
rect 50 8870 68 8902
rect 0 8834 68 8870
rect 0 8802 18 8834
rect 50 8802 68 8834
rect 0 8766 68 8802
rect 0 8734 18 8766
rect 50 8734 68 8766
rect 0 8698 68 8734
rect 0 8666 18 8698
rect 50 8666 68 8698
rect 0 8630 68 8666
rect 0 8598 18 8630
rect 50 8598 68 8630
rect 0 8562 68 8598
rect 0 8530 18 8562
rect 50 8530 68 8562
rect 0 8494 68 8530
rect 0 8462 18 8494
rect 50 8462 68 8494
rect 0 8426 68 8462
rect 0 8394 18 8426
rect 50 8394 68 8426
rect 0 8358 68 8394
rect 0 8326 18 8358
rect 50 8326 68 8358
rect 0 8290 68 8326
rect 0 8258 18 8290
rect 50 8258 68 8290
rect 0 8222 68 8258
rect 0 8190 18 8222
rect 50 8190 68 8222
rect 0 8154 68 8190
rect 0 8122 18 8154
rect 50 8122 68 8154
rect 0 8086 68 8122
rect 0 8054 18 8086
rect 50 8054 68 8086
rect 0 8018 68 8054
rect 0 7986 18 8018
rect 50 7986 68 8018
rect 0 7950 68 7986
rect 0 7918 18 7950
rect 50 7918 68 7950
rect 0 7882 68 7918
rect 0 7850 18 7882
rect 50 7850 68 7882
rect 0 7814 68 7850
rect 0 7782 18 7814
rect 50 7782 68 7814
rect 0 7746 68 7782
rect 0 7714 18 7746
rect 50 7714 68 7746
rect 0 7678 68 7714
rect 0 7646 18 7678
rect 50 7646 68 7678
rect 0 7610 68 7646
rect 0 7578 18 7610
rect 50 7578 68 7610
rect 0 7542 68 7578
rect 0 7510 18 7542
rect 50 7510 68 7542
rect 0 7474 68 7510
rect 0 7442 18 7474
rect 50 7442 68 7474
rect 0 7406 68 7442
rect 0 7374 18 7406
rect 50 7374 68 7406
rect 0 7338 68 7374
rect 0 7306 18 7338
rect 50 7306 68 7338
rect 0 7270 68 7306
rect 0 7238 18 7270
rect 50 7238 68 7270
rect 0 7202 68 7238
rect 0 7170 18 7202
rect 50 7170 68 7202
rect 0 7134 68 7170
rect 0 7102 18 7134
rect 50 7102 68 7134
rect 0 7066 68 7102
rect 0 7034 18 7066
rect 50 7034 68 7066
rect 0 6998 68 7034
rect 0 6966 18 6998
rect 50 6966 68 6998
rect 0 6930 68 6966
rect 0 6898 18 6930
rect 50 6898 68 6930
rect 0 6862 68 6898
rect 0 6830 18 6862
rect 50 6830 68 6862
rect 0 6794 68 6830
rect 0 6762 18 6794
rect 50 6762 68 6794
rect 0 6726 68 6762
rect 0 6694 18 6726
rect 50 6694 68 6726
rect 0 6658 68 6694
rect 0 6626 18 6658
rect 50 6626 68 6658
rect 0 6590 68 6626
rect 0 6558 18 6590
rect 50 6558 68 6590
rect 0 6522 68 6558
rect 0 6490 18 6522
rect 50 6490 68 6522
rect 0 6454 68 6490
rect 0 6422 18 6454
rect 50 6422 68 6454
rect 0 6386 68 6422
rect 0 6354 18 6386
rect 50 6354 68 6386
rect 0 6318 68 6354
rect 0 6286 18 6318
rect 50 6286 68 6318
rect 0 6250 68 6286
rect 0 6218 18 6250
rect 50 6218 68 6250
rect 0 6152 68 6218
rect 15932 11554 16000 11590
rect 15932 11522 15950 11554
rect 15982 11522 16000 11554
rect 15932 11486 16000 11522
rect 15932 11454 15950 11486
rect 15982 11454 16000 11486
rect 15932 11418 16000 11454
rect 15932 11386 15950 11418
rect 15982 11386 16000 11418
rect 15932 11350 16000 11386
rect 15932 11318 15950 11350
rect 15982 11318 16000 11350
rect 15932 11282 16000 11318
rect 15932 11250 15950 11282
rect 15982 11250 16000 11282
rect 15932 11214 16000 11250
rect 15932 11182 15950 11214
rect 15982 11182 16000 11214
rect 15932 11146 16000 11182
rect 15932 11114 15950 11146
rect 15982 11114 16000 11146
rect 15932 11078 16000 11114
rect 15932 11046 15950 11078
rect 15982 11046 16000 11078
rect 15932 11010 16000 11046
rect 15932 10978 15950 11010
rect 15982 10978 16000 11010
rect 15932 10942 16000 10978
rect 15932 10910 15950 10942
rect 15982 10910 16000 10942
rect 15932 10874 16000 10910
rect 15932 10842 15950 10874
rect 15982 10842 16000 10874
rect 15932 10806 16000 10842
rect 15932 10774 15950 10806
rect 15982 10774 16000 10806
rect 15932 10738 16000 10774
rect 15932 10706 15950 10738
rect 15982 10706 16000 10738
rect 15932 10670 16000 10706
rect 15932 10638 15950 10670
rect 15982 10638 16000 10670
rect 15932 10602 16000 10638
rect 15932 10570 15950 10602
rect 15982 10570 16000 10602
rect 15932 10534 16000 10570
rect 15932 10502 15950 10534
rect 15982 10502 16000 10534
rect 15932 10466 16000 10502
rect 15932 10434 15950 10466
rect 15982 10434 16000 10466
rect 15932 10398 16000 10434
rect 15932 10366 15950 10398
rect 15982 10366 16000 10398
rect 15932 10330 16000 10366
rect 15932 10298 15950 10330
rect 15982 10298 16000 10330
rect 15932 10262 16000 10298
rect 15932 10230 15950 10262
rect 15982 10230 16000 10262
rect 15932 10194 16000 10230
rect 15932 10162 15950 10194
rect 15982 10162 16000 10194
rect 15932 10126 16000 10162
rect 15932 10094 15950 10126
rect 15982 10094 16000 10126
rect 15932 10058 16000 10094
rect 15932 10026 15950 10058
rect 15982 10026 16000 10058
rect 15932 9990 16000 10026
rect 15932 9958 15950 9990
rect 15982 9958 16000 9990
rect 15932 9922 16000 9958
rect 15932 9890 15950 9922
rect 15982 9890 16000 9922
rect 15932 9854 16000 9890
rect 15932 9822 15950 9854
rect 15982 9822 16000 9854
rect 15932 9786 16000 9822
rect 15932 9754 15950 9786
rect 15982 9754 16000 9786
rect 15932 9718 16000 9754
rect 15932 9686 15950 9718
rect 15982 9686 16000 9718
rect 15932 9650 16000 9686
rect 15932 9618 15950 9650
rect 15982 9618 16000 9650
rect 15932 9582 16000 9618
rect 15932 9550 15950 9582
rect 15982 9550 16000 9582
rect 15932 9514 16000 9550
rect 15932 9482 15950 9514
rect 15982 9482 16000 9514
rect 15932 9446 16000 9482
rect 15932 9414 15950 9446
rect 15982 9414 16000 9446
rect 15932 9378 16000 9414
rect 15932 9346 15950 9378
rect 15982 9346 16000 9378
rect 15932 9310 16000 9346
rect 15932 9278 15950 9310
rect 15982 9278 16000 9310
rect 15932 9242 16000 9278
rect 15932 9210 15950 9242
rect 15982 9210 16000 9242
rect 15932 9174 16000 9210
rect 15932 9142 15950 9174
rect 15982 9142 16000 9174
rect 15932 9106 16000 9142
rect 15932 9074 15950 9106
rect 15982 9074 16000 9106
rect 15932 9038 16000 9074
rect 15932 9006 15950 9038
rect 15982 9006 16000 9038
rect 15932 8970 16000 9006
rect 15932 8938 15950 8970
rect 15982 8938 16000 8970
rect 15932 8902 16000 8938
rect 15932 8870 15950 8902
rect 15982 8870 16000 8902
rect 15932 8834 16000 8870
rect 15932 8802 15950 8834
rect 15982 8802 16000 8834
rect 15932 8766 16000 8802
rect 15932 8734 15950 8766
rect 15982 8734 16000 8766
rect 15932 8698 16000 8734
rect 15932 8666 15950 8698
rect 15982 8666 16000 8698
rect 15932 8630 16000 8666
rect 15932 8598 15950 8630
rect 15982 8598 16000 8630
rect 15932 8562 16000 8598
rect 15932 8530 15950 8562
rect 15982 8530 16000 8562
rect 15932 8494 16000 8530
rect 15932 8462 15950 8494
rect 15982 8462 16000 8494
rect 15932 8426 16000 8462
rect 15932 8394 15950 8426
rect 15982 8394 16000 8426
rect 15932 8358 16000 8394
rect 15932 8326 15950 8358
rect 15982 8326 16000 8358
rect 15932 8290 16000 8326
rect 15932 8258 15950 8290
rect 15982 8258 16000 8290
rect 15932 8222 16000 8258
rect 15932 8190 15950 8222
rect 15982 8190 16000 8222
rect 15932 8154 16000 8190
rect 15932 8122 15950 8154
rect 15982 8122 16000 8154
rect 15932 8086 16000 8122
rect 15932 8054 15950 8086
rect 15982 8054 16000 8086
rect 15932 8018 16000 8054
rect 15932 7986 15950 8018
rect 15982 7986 16000 8018
rect 15932 7950 16000 7986
rect 15932 7918 15950 7950
rect 15982 7918 16000 7950
rect 15932 7882 16000 7918
rect 15932 7850 15950 7882
rect 15982 7850 16000 7882
rect 15932 7814 16000 7850
rect 15932 7782 15950 7814
rect 15982 7782 16000 7814
rect 15932 7746 16000 7782
rect 15932 7714 15950 7746
rect 15982 7714 16000 7746
rect 15932 7678 16000 7714
rect 15932 7646 15950 7678
rect 15982 7646 16000 7678
rect 15932 7610 16000 7646
rect 15932 7578 15950 7610
rect 15982 7578 16000 7610
rect 15932 7542 16000 7578
rect 15932 7510 15950 7542
rect 15982 7510 16000 7542
rect 15932 7474 16000 7510
rect 15932 7442 15950 7474
rect 15982 7442 16000 7474
rect 15932 7406 16000 7442
rect 15932 7374 15950 7406
rect 15982 7374 16000 7406
rect 15932 7338 16000 7374
rect 15932 7306 15950 7338
rect 15982 7306 16000 7338
rect 15932 7270 16000 7306
rect 15932 7238 15950 7270
rect 15982 7238 16000 7270
rect 15932 7202 16000 7238
rect 15932 7170 15950 7202
rect 15982 7170 16000 7202
rect 15932 7134 16000 7170
rect 15932 7102 15950 7134
rect 15982 7102 16000 7134
rect 15932 7066 16000 7102
rect 15932 7034 15950 7066
rect 15982 7034 16000 7066
rect 15932 6998 16000 7034
rect 15932 6966 15950 6998
rect 15982 6966 16000 6998
rect 15932 6930 16000 6966
rect 15932 6898 15950 6930
rect 15982 6898 16000 6930
rect 15932 6862 16000 6898
rect 15932 6830 15950 6862
rect 15982 6830 16000 6862
rect 15932 6794 16000 6830
rect 15932 6762 15950 6794
rect 15982 6762 16000 6794
rect 15932 6726 16000 6762
rect 15932 6694 15950 6726
rect 15982 6694 16000 6726
rect 15932 6658 16000 6694
rect 15932 6626 15950 6658
rect 15982 6626 16000 6658
rect 15932 6590 16000 6626
rect 15932 6558 15950 6590
rect 15982 6558 16000 6590
rect 15932 6522 16000 6558
rect 15932 6490 15950 6522
rect 15982 6490 16000 6522
rect 15932 6454 16000 6490
rect 15932 6422 15950 6454
rect 15982 6422 16000 6454
rect 15932 6386 16000 6422
rect 15932 6354 15950 6386
rect 15982 6354 16000 6386
rect 15932 6318 16000 6354
rect 15932 6286 15950 6318
rect 15982 6286 16000 6318
rect 15932 6250 16000 6286
rect 15932 6218 15950 6250
rect 15982 6218 16000 6250
rect 15932 6152 16000 6218
rect 0 6134 16000 6152
rect 0 6102 28 6134
rect 60 6102 96 6134
rect 128 6102 164 6134
rect 196 6102 232 6134
rect 264 6102 300 6134
rect 332 6102 368 6134
rect 400 6102 436 6134
rect 468 6102 504 6134
rect 536 6102 572 6134
rect 604 6102 640 6134
rect 672 6102 708 6134
rect 740 6102 776 6134
rect 808 6102 844 6134
rect 876 6102 912 6134
rect 944 6102 980 6134
rect 1012 6102 1048 6134
rect 1080 6102 1116 6134
rect 1148 6102 1184 6134
rect 1216 6102 1252 6134
rect 1284 6102 1320 6134
rect 1352 6102 1388 6134
rect 1420 6102 1456 6134
rect 1488 6102 1524 6134
rect 1556 6102 1592 6134
rect 1624 6102 1660 6134
rect 1692 6102 1728 6134
rect 1760 6104 1796 6134
rect 1828 6104 1864 6134
rect 1760 6102 1789 6104
rect 1829 6102 1864 6104
rect 1896 6102 1932 6134
rect 1964 6102 2000 6134
rect 2032 6102 2068 6134
rect 2100 6102 2136 6134
rect 2168 6102 2204 6134
rect 2236 6102 2272 6134
rect 2304 6102 2340 6134
rect 2372 6104 2408 6134
rect 2372 6102 2393 6104
rect 2440 6102 2476 6134
rect 2508 6102 2544 6134
rect 2576 6102 2612 6134
rect 2644 6102 2680 6134
rect 2712 6102 2748 6134
rect 2780 6102 2816 6134
rect 2848 6102 2884 6134
rect 2916 6102 2952 6134
rect 2984 6104 3020 6134
rect 2984 6102 2997 6104
rect 3052 6102 3088 6134
rect 3120 6102 3156 6134
rect 3188 6102 3224 6134
rect 3256 6102 3292 6134
rect 3324 6102 3360 6134
rect 3392 6102 3428 6134
rect 3460 6102 3496 6134
rect 3528 6102 3564 6134
rect 3596 6104 3632 6134
rect 3596 6102 3601 6104
rect 3664 6102 3700 6134
rect 3732 6102 3768 6134
rect 3800 6102 3836 6134
rect 3868 6102 3904 6134
rect 3936 6102 3972 6134
rect 4004 6102 4040 6134
rect 4072 6102 4108 6134
rect 4140 6102 4176 6134
rect 4208 6104 4244 6134
rect 4276 6102 4312 6134
rect 4344 6102 4380 6134
rect 4412 6102 4448 6134
rect 4480 6102 4516 6134
rect 4548 6102 4584 6134
rect 4616 6102 4652 6134
rect 4684 6102 4720 6134
rect 4752 6102 4788 6134
rect 4820 6104 4856 6134
rect 4849 6102 4856 6104
rect 4888 6102 4924 6134
rect 4956 6102 4992 6134
rect 5024 6102 5060 6134
rect 5092 6102 5128 6134
rect 5160 6102 5196 6134
rect 5228 6102 5264 6134
rect 5296 6102 5332 6134
rect 5364 6102 5400 6134
rect 5432 6104 5468 6134
rect 5453 6102 5468 6104
rect 5500 6102 5536 6134
rect 5568 6102 5604 6134
rect 5636 6102 5672 6134
rect 5704 6102 5740 6134
rect 5772 6102 5808 6134
rect 5840 6102 5876 6134
rect 5908 6102 5944 6134
rect 5976 6102 6012 6134
rect 6044 6104 6080 6134
rect 6057 6102 6080 6104
rect 6112 6102 6148 6134
rect 6180 6102 6216 6134
rect 6248 6102 6284 6134
rect 6316 6102 6352 6134
rect 6384 6102 6420 6134
rect 6452 6102 6488 6134
rect 6520 6102 6556 6134
rect 6588 6104 6624 6134
rect 6656 6104 6692 6134
rect 6588 6102 6621 6104
rect 6661 6102 6692 6104
rect 6724 6102 6760 6134
rect 6792 6102 6828 6134
rect 6860 6102 6896 6134
rect 6928 6102 6964 6134
rect 6996 6102 7032 6134
rect 7064 6102 7100 6134
rect 7132 6102 7168 6134
rect 7200 6104 7236 6134
rect 7200 6102 7225 6104
rect 7268 6102 7304 6134
rect 7336 6102 7372 6134
rect 7404 6102 7440 6134
rect 7472 6102 7508 6134
rect 7540 6102 7576 6134
rect 7608 6102 7644 6134
rect 7676 6102 7712 6134
rect 7744 6102 7780 6134
rect 7812 6104 7848 6134
rect 7812 6102 7829 6104
rect 7880 6102 7916 6134
rect 7948 6102 7984 6134
rect 8016 6102 8052 6134
rect 8084 6102 8120 6134
rect 8152 6102 8188 6134
rect 8220 6102 8256 6134
rect 8288 6102 8324 6134
rect 8356 6102 8392 6134
rect 8424 6104 8460 6134
rect 8424 6102 8433 6104
rect 8492 6102 8528 6134
rect 8560 6102 8596 6134
rect 8628 6102 8664 6134
rect 8696 6102 8732 6134
rect 8764 6102 8800 6134
rect 8832 6102 8868 6134
rect 8900 6102 8936 6134
rect 8968 6102 9004 6134
rect 9036 6104 9072 6134
rect 9036 6102 9037 6104
rect 9104 6102 9140 6134
rect 9172 6102 9208 6134
rect 9240 6102 9276 6134
rect 9308 6102 9344 6134
rect 9376 6102 9412 6134
rect 9444 6102 9480 6134
rect 9512 6102 9548 6134
rect 9580 6102 9616 6134
rect 9648 6104 9684 6134
rect 9681 6102 9684 6104
rect 9716 6102 9752 6134
rect 9784 6102 9820 6134
rect 9852 6102 9888 6134
rect 9920 6102 9956 6134
rect 9988 6102 10024 6134
rect 10056 6102 10092 6134
rect 10124 6102 10160 6134
rect 10192 6102 10228 6134
rect 10260 6104 10296 6134
rect 10285 6102 10296 6104
rect 10328 6102 10364 6134
rect 10396 6102 10432 6134
rect 10464 6102 10500 6134
rect 10532 6102 10568 6134
rect 10600 6102 10636 6134
rect 10668 6102 10704 6134
rect 10736 6102 10772 6134
rect 10804 6102 10840 6134
rect 10872 6104 10908 6134
rect 10889 6102 10908 6104
rect 10940 6102 10976 6134
rect 11008 6102 11044 6134
rect 11076 6102 11112 6134
rect 11144 6102 11180 6134
rect 11212 6102 11248 6134
rect 11280 6102 11316 6134
rect 11348 6102 11384 6134
rect 11416 6102 11452 6134
rect 11484 6104 11520 6134
rect 11493 6102 11520 6104
rect 11552 6102 11588 6134
rect 11620 6102 11656 6134
rect 11688 6102 11724 6134
rect 11756 6102 11792 6134
rect 11824 6102 11860 6134
rect 11892 6102 11928 6134
rect 11960 6102 11996 6134
rect 12028 6104 12064 6134
rect 12096 6104 12132 6134
rect 12028 6102 12057 6104
rect 12097 6102 12132 6104
rect 12164 6102 12200 6134
rect 12232 6102 12268 6134
rect 12300 6102 12336 6134
rect 12368 6102 12404 6134
rect 12436 6102 12472 6134
rect 12504 6102 12540 6134
rect 12572 6102 12608 6134
rect 12640 6104 12676 6134
rect 12640 6102 12661 6104
rect 12708 6102 12744 6134
rect 12776 6102 12812 6134
rect 12844 6102 12880 6134
rect 12912 6102 12948 6134
rect 12980 6102 13016 6134
rect 13048 6102 13084 6134
rect 13116 6102 13152 6134
rect 13184 6102 13220 6134
rect 13252 6104 13288 6134
rect 13252 6102 13265 6104
rect 13320 6102 13356 6134
rect 13388 6102 13424 6134
rect 13456 6102 13492 6134
rect 13524 6102 13560 6134
rect 13592 6102 13628 6134
rect 13660 6102 13696 6134
rect 13728 6102 13764 6134
rect 13796 6102 13832 6134
rect 13864 6104 13900 6134
rect 13864 6102 13869 6104
rect 13932 6102 13968 6134
rect 14000 6102 14036 6134
rect 14068 6102 14104 6134
rect 14136 6102 14172 6134
rect 14204 6102 14240 6134
rect 14272 6102 14308 6134
rect 14340 6102 14376 6134
rect 14408 6102 14444 6134
rect 14476 6104 14512 6134
rect 14544 6102 14580 6134
rect 14612 6102 14648 6134
rect 14680 6102 14716 6134
rect 14748 6102 14784 6134
rect 14816 6102 14852 6134
rect 14884 6102 14920 6134
rect 14952 6102 14988 6134
rect 15020 6102 15056 6134
rect 15088 6102 15124 6134
rect 15156 6102 15192 6134
rect 15224 6102 15260 6134
rect 15292 6102 15328 6134
rect 15360 6102 15396 6134
rect 15428 6102 15464 6134
rect 15496 6102 15532 6134
rect 15564 6102 15600 6134
rect 15632 6102 15668 6134
rect 15700 6102 15736 6134
rect 15768 6102 15804 6134
rect 15836 6102 15872 6134
rect 15904 6102 15940 6134
rect 15972 6102 16000 6134
rect 0 6084 1789 6102
rect 0 1200 32 6084
rect 1748 6064 1789 6084
rect 1829 6084 2393 6102
rect 1829 6064 1870 6084
rect 1748 6055 1870 6064
rect 2352 6064 2393 6084
rect 2433 6084 2997 6102
rect 2433 6064 2474 6084
rect 2352 6055 2474 6064
rect 2956 6064 2997 6084
rect 3037 6084 3601 6102
rect 3037 6064 3078 6084
rect 2956 6055 3078 6064
rect 3560 6064 3601 6084
rect 3641 6084 4205 6102
rect 3641 6064 3682 6084
rect 3560 6055 3682 6064
rect 4164 6064 4205 6084
rect 4245 6084 4809 6102
rect 4245 6064 4286 6084
rect 4164 6055 4286 6064
rect 4768 6064 4809 6084
rect 4849 6084 5413 6102
rect 4849 6064 4890 6084
rect 4768 6055 4890 6064
rect 5372 6064 5413 6084
rect 5453 6084 6017 6102
rect 5453 6064 5494 6084
rect 5372 6055 5494 6064
rect 5976 6064 6017 6084
rect 6057 6084 6621 6102
rect 6057 6064 6098 6084
rect 5976 6055 6098 6064
rect 6580 6064 6621 6084
rect 6661 6084 7225 6102
rect 6661 6064 6702 6084
rect 6580 6055 6702 6064
rect 7184 6064 7225 6084
rect 7265 6084 7829 6102
rect 7265 6064 7306 6084
rect 7184 6055 7306 6064
rect 7788 6064 7829 6084
rect 7869 6084 8433 6102
rect 7869 6064 7910 6084
rect 7788 6055 7910 6064
rect 8392 6064 8433 6084
rect 8473 6084 9037 6102
rect 8473 6064 8514 6084
rect 8392 6055 8514 6064
rect 8996 6064 9037 6084
rect 9077 6084 9641 6102
rect 9077 6064 9118 6084
rect 8996 6055 9118 6064
rect 9600 6064 9641 6084
rect 9681 6084 10245 6102
rect 9681 6064 9722 6084
rect 9600 6055 9722 6064
rect 10204 6064 10245 6084
rect 10285 6084 10849 6102
rect 10285 6064 10326 6084
rect 10204 6055 10326 6064
rect 10808 6064 10849 6084
rect 10889 6084 11453 6102
rect 10889 6064 10930 6084
rect 10808 6055 10930 6064
rect 11412 6064 11453 6084
rect 11493 6084 12057 6102
rect 11493 6064 11534 6084
rect 11412 6055 11534 6064
rect 12016 6064 12057 6084
rect 12097 6084 12661 6102
rect 12097 6064 12138 6084
rect 12016 6055 12138 6064
rect 12620 6064 12661 6084
rect 12701 6084 13265 6102
rect 12701 6064 12742 6084
rect 12620 6055 12742 6064
rect 13224 6064 13265 6084
rect 13305 6084 13869 6102
rect 13305 6064 13346 6084
rect 13224 6055 13346 6064
rect 13828 6064 13869 6084
rect 13909 6084 14473 6102
rect 13909 6064 13950 6084
rect 13828 6055 13950 6064
rect 14432 6064 14473 6084
rect 14513 6084 16000 6102
rect 14513 6064 14554 6084
rect 14432 6055 14554 6064
rect 15968 1200 16000 6084
<< via1 >>
rect 42 33416 656 33420
rect 15344 33416 15958 33420
rect 42 33384 50 33416
rect 50 33384 82 33416
rect 82 33384 118 33416
rect 118 33384 150 33416
rect 150 33384 186 33416
rect 186 33384 218 33416
rect 218 33384 254 33416
rect 254 33384 286 33416
rect 286 33384 322 33416
rect 322 33384 354 33416
rect 354 33384 390 33416
rect 390 33384 422 33416
rect 422 33384 458 33416
rect 458 33384 490 33416
rect 490 33384 526 33416
rect 526 33384 558 33416
rect 558 33384 594 33416
rect 594 33384 626 33416
rect 626 33384 656 33416
rect 15344 33384 15350 33416
rect 15350 33384 15382 33416
rect 15382 33384 15442 33416
rect 15442 33384 15474 33416
rect 15474 33384 15510 33416
rect 15510 33384 15542 33416
rect 15542 33384 15578 33416
rect 15578 33384 15610 33416
rect 15610 33384 15646 33416
rect 15646 33384 15678 33416
rect 15678 33384 15714 33416
rect 15714 33384 15746 33416
rect 15746 33384 15782 33416
rect 15782 33384 15814 33416
rect 15814 33384 15850 33416
rect 15850 33384 15882 33416
rect 15882 33384 15918 33416
rect 15918 33384 15950 33416
rect 15950 33384 15958 33416
rect 42 33380 656 33384
rect 15344 33380 15958 33384
rect 42 31416 656 31420
rect 15344 31416 15958 31420
rect 42 31384 50 31416
rect 50 31384 82 31416
rect 82 31384 118 31416
rect 118 31384 150 31416
rect 150 31384 186 31416
rect 186 31384 218 31416
rect 218 31384 254 31416
rect 254 31384 286 31416
rect 286 31384 322 31416
rect 322 31384 354 31416
rect 354 31384 390 31416
rect 390 31384 422 31416
rect 422 31384 458 31416
rect 458 31384 490 31416
rect 490 31384 526 31416
rect 526 31384 558 31416
rect 558 31384 594 31416
rect 594 31384 626 31416
rect 626 31384 656 31416
rect 15344 31384 15350 31416
rect 15350 31384 15382 31416
rect 15382 31384 15442 31416
rect 15442 31384 15474 31416
rect 15474 31384 15510 31416
rect 15510 31384 15542 31416
rect 15542 31384 15578 31416
rect 15578 31384 15610 31416
rect 15610 31384 15646 31416
rect 15646 31384 15678 31416
rect 15678 31384 15714 31416
rect 15714 31384 15746 31416
rect 15746 31384 15782 31416
rect 15782 31384 15814 31416
rect 15814 31384 15850 31416
rect 15850 31384 15882 31416
rect 15882 31384 15918 31416
rect 15918 31384 15950 31416
rect 15950 31384 15958 31416
rect 42 31380 656 31384
rect 15344 31380 15958 31384
rect 15836 29716 15958 29720
rect 15836 29684 15850 29716
rect 15850 29684 15882 29716
rect 15882 29684 15918 29716
rect 15918 29684 15950 29716
rect 15950 29684 15958 29716
rect 15836 29680 15958 29684
rect 51 26747 91 26755
rect 149 26747 189 26755
rect 247 26747 287 26755
rect 345 26747 385 26755
rect 443 26747 483 26755
rect 541 26747 581 26755
rect 639 26747 679 26755
rect 737 26747 777 26755
rect 835 26747 875 26755
rect 933 26747 973 26755
rect 1031 26747 1071 26755
rect 1129 26747 1169 26755
rect 51 26715 64 26747
rect 64 26715 91 26747
rect 149 26715 168 26747
rect 168 26715 189 26747
rect 247 26715 280 26747
rect 280 26715 287 26747
rect 345 26715 352 26747
rect 352 26715 384 26747
rect 384 26715 385 26747
rect 443 26715 456 26747
rect 456 26715 483 26747
rect 541 26715 568 26747
rect 568 26715 581 26747
rect 639 26715 640 26747
rect 640 26715 672 26747
rect 672 26715 679 26747
rect 737 26715 744 26747
rect 744 26715 777 26747
rect 835 26715 856 26747
rect 856 26715 875 26747
rect 933 26715 960 26747
rect 960 26715 973 26747
rect 1031 26715 1032 26747
rect 1032 26715 1071 26747
rect 1129 26715 1144 26747
rect 1144 26715 1169 26747
rect 51 26643 64 26657
rect 64 26643 91 26657
rect 149 26643 168 26657
rect 168 26643 189 26657
rect 247 26643 280 26657
rect 280 26643 287 26657
rect 345 26643 352 26657
rect 352 26643 384 26657
rect 384 26643 385 26657
rect 443 26643 456 26657
rect 456 26643 483 26657
rect 541 26643 568 26657
rect 568 26643 581 26657
rect 639 26643 640 26657
rect 640 26643 672 26657
rect 672 26643 679 26657
rect 737 26643 744 26657
rect 744 26643 777 26657
rect 835 26643 856 26657
rect 856 26643 875 26657
rect 933 26643 960 26657
rect 960 26643 973 26657
rect 1031 26643 1032 26657
rect 1032 26643 1071 26657
rect 1129 26643 1144 26657
rect 1144 26643 1169 26657
rect 51 26617 91 26643
rect 149 26617 189 26643
rect 247 26617 287 26643
rect 345 26617 385 26643
rect 443 26617 483 26643
rect 541 26617 581 26643
rect 639 26617 679 26643
rect 737 26617 777 26643
rect 835 26617 875 26643
rect 933 26617 973 26643
rect 1031 26617 1071 26643
rect 1129 26617 1169 26643
rect 51 26531 91 26559
rect 149 26531 189 26559
rect 247 26531 287 26559
rect 345 26531 385 26559
rect 443 26531 483 26559
rect 541 26531 581 26559
rect 639 26531 679 26559
rect 737 26531 777 26559
rect 835 26531 875 26559
rect 933 26531 973 26559
rect 1031 26531 1071 26559
rect 1129 26531 1169 26559
rect 51 26519 64 26531
rect 64 26519 91 26531
rect 149 26519 168 26531
rect 168 26519 189 26531
rect 247 26519 280 26531
rect 280 26519 287 26531
rect 345 26519 352 26531
rect 352 26519 384 26531
rect 384 26519 385 26531
rect 443 26519 456 26531
rect 456 26519 483 26531
rect 541 26519 568 26531
rect 568 26519 581 26531
rect 639 26519 640 26531
rect 640 26519 672 26531
rect 672 26519 679 26531
rect 737 26519 744 26531
rect 744 26519 777 26531
rect 835 26519 856 26531
rect 856 26519 875 26531
rect 933 26519 960 26531
rect 960 26519 973 26531
rect 1031 26519 1032 26531
rect 1032 26519 1071 26531
rect 1129 26519 1144 26531
rect 1144 26519 1169 26531
rect 51 26459 91 26461
rect 149 26459 189 26461
rect 247 26459 287 26461
rect 345 26459 385 26461
rect 443 26459 483 26461
rect 541 26459 581 26461
rect 639 26459 679 26461
rect 737 26459 777 26461
rect 835 26459 875 26461
rect 933 26459 973 26461
rect 1031 26459 1071 26461
rect 1129 26459 1169 26461
rect 51 26427 64 26459
rect 64 26427 91 26459
rect 149 26427 168 26459
rect 168 26427 189 26459
rect 247 26427 280 26459
rect 280 26427 287 26459
rect 345 26427 352 26459
rect 352 26427 384 26459
rect 384 26427 385 26459
rect 443 26427 456 26459
rect 456 26427 483 26459
rect 541 26427 568 26459
rect 568 26427 581 26459
rect 639 26427 640 26459
rect 640 26427 672 26459
rect 672 26427 679 26459
rect 737 26427 744 26459
rect 744 26427 777 26459
rect 835 26427 856 26459
rect 856 26427 875 26459
rect 933 26427 960 26459
rect 960 26427 973 26459
rect 1031 26427 1032 26459
rect 1032 26427 1071 26459
rect 1129 26427 1144 26459
rect 1144 26427 1169 26459
rect 51 26421 91 26427
rect 149 26421 189 26427
rect 247 26421 287 26427
rect 345 26421 385 26427
rect 443 26421 483 26427
rect 541 26421 581 26427
rect 639 26421 679 26427
rect 737 26421 777 26427
rect 835 26421 875 26427
rect 933 26421 973 26427
rect 1031 26421 1071 26427
rect 1129 26421 1169 26427
rect 51 26355 64 26363
rect 64 26355 91 26363
rect 149 26355 168 26363
rect 168 26355 189 26363
rect 247 26355 280 26363
rect 280 26355 287 26363
rect 345 26355 352 26363
rect 352 26355 384 26363
rect 384 26355 385 26363
rect 443 26355 456 26363
rect 456 26355 483 26363
rect 541 26355 568 26363
rect 568 26355 581 26363
rect 639 26355 640 26363
rect 640 26355 672 26363
rect 672 26355 679 26363
rect 737 26355 744 26363
rect 744 26355 777 26363
rect 835 26355 856 26363
rect 856 26355 875 26363
rect 933 26355 960 26363
rect 960 26355 973 26363
rect 1031 26355 1032 26363
rect 1032 26355 1071 26363
rect 1129 26355 1144 26363
rect 1144 26355 1169 26363
rect 51 26323 91 26355
rect 149 26323 189 26355
rect 247 26323 287 26355
rect 345 26323 385 26355
rect 443 26323 483 26355
rect 541 26323 581 26355
rect 639 26323 679 26355
rect 737 26323 777 26355
rect 835 26323 875 26355
rect 933 26323 973 26355
rect 1031 26323 1071 26355
rect 1129 26323 1169 26355
rect 51 26243 91 26265
rect 149 26243 189 26265
rect 247 26243 287 26265
rect 345 26243 385 26265
rect 443 26243 483 26265
rect 541 26243 581 26265
rect 639 26243 679 26265
rect 737 26243 777 26265
rect 835 26243 875 26265
rect 933 26243 973 26265
rect 1031 26243 1071 26265
rect 1129 26243 1169 26265
rect 51 26225 64 26243
rect 64 26225 91 26243
rect 149 26225 168 26243
rect 168 26225 189 26243
rect 247 26225 280 26243
rect 280 26225 287 26243
rect 345 26225 352 26243
rect 352 26225 384 26243
rect 384 26225 385 26243
rect 443 26225 456 26243
rect 456 26225 483 26243
rect 541 26225 568 26243
rect 568 26225 581 26243
rect 639 26225 640 26243
rect 640 26225 672 26243
rect 672 26225 679 26243
rect 737 26225 744 26243
rect 744 26225 777 26243
rect 835 26225 856 26243
rect 856 26225 875 26243
rect 933 26225 960 26243
rect 960 26225 973 26243
rect 1031 26225 1032 26243
rect 1032 26225 1071 26243
rect 1129 26225 1144 26243
rect 1144 26225 1169 26243
rect 51 26139 64 26167
rect 64 26139 91 26167
rect 149 26139 168 26167
rect 168 26139 189 26167
rect 247 26139 280 26167
rect 280 26139 287 26167
rect 345 26139 352 26167
rect 352 26139 384 26167
rect 384 26139 385 26167
rect 443 26139 456 26167
rect 456 26139 483 26167
rect 541 26139 568 26167
rect 568 26139 581 26167
rect 639 26139 640 26167
rect 640 26139 672 26167
rect 672 26139 679 26167
rect 737 26139 744 26167
rect 744 26139 777 26167
rect 835 26139 856 26167
rect 856 26139 875 26167
rect 933 26139 960 26167
rect 960 26139 973 26167
rect 1031 26139 1032 26167
rect 1032 26139 1071 26167
rect 1129 26139 1144 26167
rect 1144 26139 1169 26167
rect 51 26127 91 26139
rect 149 26127 189 26139
rect 247 26127 287 26139
rect 345 26127 385 26139
rect 443 26127 483 26139
rect 541 26127 581 26139
rect 639 26127 679 26139
rect 737 26127 777 26139
rect 835 26127 875 26139
rect 933 26127 973 26139
rect 1031 26127 1071 26139
rect 1129 26127 1169 26139
rect 51 26067 64 26069
rect 64 26067 91 26069
rect 149 26067 168 26069
rect 168 26067 189 26069
rect 247 26067 280 26069
rect 280 26067 287 26069
rect 345 26067 352 26069
rect 352 26067 384 26069
rect 384 26067 385 26069
rect 443 26067 456 26069
rect 456 26067 483 26069
rect 541 26067 568 26069
rect 568 26067 581 26069
rect 639 26067 640 26069
rect 640 26067 672 26069
rect 672 26067 679 26069
rect 737 26067 744 26069
rect 744 26067 777 26069
rect 835 26067 856 26069
rect 856 26067 875 26069
rect 933 26067 960 26069
rect 960 26067 973 26069
rect 1031 26067 1032 26069
rect 1032 26067 1071 26069
rect 1129 26067 1144 26069
rect 1144 26067 1169 26069
rect 51 26029 91 26067
rect 149 26029 189 26067
rect 247 26029 287 26067
rect 345 26029 385 26067
rect 443 26029 483 26067
rect 541 26029 581 26067
rect 639 26029 679 26067
rect 737 26029 777 26067
rect 835 26029 875 26067
rect 933 26029 973 26067
rect 1031 26029 1071 26067
rect 1129 26029 1169 26067
rect 51 25955 91 25971
rect 149 25955 189 25971
rect 247 25955 287 25971
rect 345 25955 385 25971
rect 443 25955 483 25971
rect 541 25955 581 25971
rect 639 25955 679 25971
rect 737 25955 777 25971
rect 835 25955 875 25971
rect 933 25955 973 25971
rect 1031 25955 1071 25971
rect 1129 25955 1169 25971
rect 51 25931 64 25955
rect 64 25931 91 25955
rect 149 25931 168 25955
rect 168 25931 189 25955
rect 247 25931 280 25955
rect 280 25931 287 25955
rect 345 25931 352 25955
rect 352 25931 384 25955
rect 384 25931 385 25955
rect 443 25931 456 25955
rect 456 25931 483 25955
rect 541 25931 568 25955
rect 568 25931 581 25955
rect 639 25931 640 25955
rect 640 25931 672 25955
rect 672 25931 679 25955
rect 737 25931 744 25955
rect 744 25931 777 25955
rect 835 25931 856 25955
rect 856 25931 875 25955
rect 933 25931 960 25955
rect 960 25931 973 25955
rect 1031 25931 1032 25955
rect 1032 25931 1071 25955
rect 1129 25931 1144 25955
rect 1144 25931 1169 25955
rect 51 25851 64 25873
rect 64 25851 91 25873
rect 149 25851 168 25873
rect 168 25851 189 25873
rect 247 25851 280 25873
rect 280 25851 287 25873
rect 345 25851 352 25873
rect 352 25851 384 25873
rect 384 25851 385 25873
rect 443 25851 456 25873
rect 456 25851 483 25873
rect 541 25851 568 25873
rect 568 25851 581 25873
rect 639 25851 640 25873
rect 640 25851 672 25873
rect 672 25851 679 25873
rect 737 25851 744 25873
rect 744 25851 777 25873
rect 835 25851 856 25873
rect 856 25851 875 25873
rect 933 25851 960 25873
rect 960 25851 973 25873
rect 1031 25851 1032 25873
rect 1032 25851 1071 25873
rect 1129 25851 1144 25873
rect 1144 25851 1169 25873
rect 51 25833 91 25851
rect 149 25833 189 25851
rect 247 25833 287 25851
rect 345 25833 385 25851
rect 443 25833 483 25851
rect 541 25833 581 25851
rect 639 25833 679 25851
rect 737 25833 777 25851
rect 835 25833 875 25851
rect 933 25833 973 25851
rect 1031 25833 1071 25851
rect 1129 25833 1169 25851
rect 51 25739 91 25775
rect 149 25739 189 25775
rect 247 25739 287 25775
rect 345 25739 385 25775
rect 443 25739 483 25775
rect 541 25739 581 25775
rect 639 25739 679 25775
rect 737 25739 777 25775
rect 835 25739 875 25775
rect 933 25739 973 25775
rect 1031 25739 1071 25775
rect 1129 25739 1169 25775
rect 51 25735 64 25739
rect 64 25735 91 25739
rect 149 25735 168 25739
rect 168 25735 189 25739
rect 247 25735 280 25739
rect 280 25735 287 25739
rect 345 25735 352 25739
rect 352 25735 384 25739
rect 384 25735 385 25739
rect 443 25735 456 25739
rect 456 25735 483 25739
rect 541 25735 568 25739
rect 568 25735 581 25739
rect 639 25735 640 25739
rect 640 25735 672 25739
rect 672 25735 679 25739
rect 737 25735 744 25739
rect 744 25735 777 25739
rect 835 25735 856 25739
rect 856 25735 875 25739
rect 933 25735 960 25739
rect 960 25735 973 25739
rect 1031 25735 1032 25739
rect 1032 25735 1071 25739
rect 1129 25735 1144 25739
rect 1144 25735 1169 25739
rect 51 25667 91 25677
rect 149 25667 189 25677
rect 247 25667 287 25677
rect 345 25667 385 25677
rect 443 25667 483 25677
rect 541 25667 581 25677
rect 639 25667 679 25677
rect 737 25667 777 25677
rect 835 25667 875 25677
rect 933 25667 973 25677
rect 1031 25667 1071 25677
rect 1129 25667 1169 25677
rect 51 25637 64 25667
rect 64 25637 91 25667
rect 149 25637 168 25667
rect 168 25637 189 25667
rect 247 25637 280 25667
rect 280 25637 287 25667
rect 345 25637 352 25667
rect 352 25637 384 25667
rect 384 25637 385 25667
rect 443 25637 456 25667
rect 456 25637 483 25667
rect 541 25637 568 25667
rect 568 25637 581 25667
rect 639 25637 640 25667
rect 640 25637 672 25667
rect 672 25637 679 25667
rect 737 25637 744 25667
rect 744 25637 777 25667
rect 835 25637 856 25667
rect 856 25637 875 25667
rect 933 25637 960 25667
rect 960 25637 973 25667
rect 1031 25637 1032 25667
rect 1032 25637 1071 25667
rect 1129 25637 1144 25667
rect 1144 25637 1169 25667
rect 51 25563 64 25579
rect 64 25563 91 25579
rect 149 25563 168 25579
rect 168 25563 189 25579
rect 247 25563 280 25579
rect 280 25563 287 25579
rect 345 25563 352 25579
rect 352 25563 384 25579
rect 384 25563 385 25579
rect 443 25563 456 25579
rect 456 25563 483 25579
rect 541 25563 568 25579
rect 568 25563 581 25579
rect 639 25563 640 25579
rect 640 25563 672 25579
rect 672 25563 679 25579
rect 737 25563 744 25579
rect 744 25563 777 25579
rect 835 25563 856 25579
rect 856 25563 875 25579
rect 933 25563 960 25579
rect 960 25563 973 25579
rect 1031 25563 1032 25579
rect 1032 25563 1071 25579
rect 1129 25563 1144 25579
rect 1144 25563 1169 25579
rect 51 25539 91 25563
rect 149 25539 189 25563
rect 247 25539 287 25563
rect 345 25539 385 25563
rect 443 25539 483 25563
rect 541 25539 581 25563
rect 639 25539 679 25563
rect 737 25539 777 25563
rect 835 25539 875 25563
rect 933 25539 973 25563
rect 1031 25539 1071 25563
rect 1129 25539 1169 25563
rect 51 25451 91 25481
rect 149 25451 189 25481
rect 247 25451 287 25481
rect 345 25451 385 25481
rect 443 25451 483 25481
rect 541 25451 581 25481
rect 639 25451 679 25481
rect 737 25451 777 25481
rect 835 25451 875 25481
rect 933 25451 973 25481
rect 1031 25451 1071 25481
rect 1129 25451 1169 25481
rect 51 25441 64 25451
rect 64 25441 91 25451
rect 149 25441 168 25451
rect 168 25441 189 25451
rect 247 25441 280 25451
rect 280 25441 287 25451
rect 345 25441 352 25451
rect 352 25441 384 25451
rect 384 25441 385 25451
rect 443 25441 456 25451
rect 456 25441 483 25451
rect 541 25441 568 25451
rect 568 25441 581 25451
rect 639 25441 640 25451
rect 640 25441 672 25451
rect 672 25441 679 25451
rect 737 25441 744 25451
rect 744 25441 777 25451
rect 835 25441 856 25451
rect 856 25441 875 25451
rect 933 25441 960 25451
rect 960 25441 973 25451
rect 1031 25441 1032 25451
rect 1032 25441 1071 25451
rect 1129 25441 1144 25451
rect 1144 25441 1169 25451
rect 51 25379 91 25383
rect 149 25379 189 25383
rect 247 25379 287 25383
rect 345 25379 385 25383
rect 443 25379 483 25383
rect 541 25379 581 25383
rect 639 25379 679 25383
rect 737 25379 777 25383
rect 835 25379 875 25383
rect 933 25379 973 25383
rect 1031 25379 1071 25383
rect 1129 25379 1169 25383
rect 51 25347 64 25379
rect 64 25347 91 25379
rect 149 25347 168 25379
rect 168 25347 189 25379
rect 247 25347 280 25379
rect 280 25347 287 25379
rect 345 25347 352 25379
rect 352 25347 384 25379
rect 384 25347 385 25379
rect 443 25347 456 25379
rect 456 25347 483 25379
rect 541 25347 568 25379
rect 568 25347 581 25379
rect 639 25347 640 25379
rect 640 25347 672 25379
rect 672 25347 679 25379
rect 737 25347 744 25379
rect 744 25347 777 25379
rect 835 25347 856 25379
rect 856 25347 875 25379
rect 933 25347 960 25379
rect 960 25347 973 25379
rect 1031 25347 1032 25379
rect 1032 25347 1071 25379
rect 1129 25347 1144 25379
rect 1144 25347 1169 25379
rect 51 25343 91 25347
rect 149 25343 189 25347
rect 247 25343 287 25347
rect 345 25343 385 25347
rect 443 25343 483 25347
rect 541 25343 581 25347
rect 639 25343 679 25347
rect 737 25343 777 25347
rect 835 25343 875 25347
rect 933 25343 973 25347
rect 1031 25343 1071 25347
rect 1129 25343 1169 25347
rect 51 25275 64 25285
rect 64 25275 91 25285
rect 149 25275 168 25285
rect 168 25275 189 25285
rect 247 25275 280 25285
rect 280 25275 287 25285
rect 345 25275 352 25285
rect 352 25275 384 25285
rect 384 25275 385 25285
rect 443 25275 456 25285
rect 456 25275 483 25285
rect 541 25275 568 25285
rect 568 25275 581 25285
rect 639 25275 640 25285
rect 640 25275 672 25285
rect 672 25275 679 25285
rect 737 25275 744 25285
rect 744 25275 777 25285
rect 835 25275 856 25285
rect 856 25275 875 25285
rect 933 25275 960 25285
rect 960 25275 973 25285
rect 1031 25275 1032 25285
rect 1032 25275 1071 25285
rect 1129 25275 1144 25285
rect 1144 25275 1169 25285
rect 51 25245 91 25275
rect 149 25245 189 25275
rect 247 25245 287 25275
rect 345 25245 385 25275
rect 443 25245 483 25275
rect 541 25245 581 25275
rect 639 25245 679 25275
rect 737 25245 777 25275
rect 835 25245 875 25275
rect 933 25245 973 25275
rect 1031 25245 1071 25275
rect 1129 25245 1169 25275
rect 3306 20031 12694 20071
rect 12064 12519 15384 12559
rect 3836 11578 3958 11618
rect 1789 6102 1796 6104
rect 1796 6102 1828 6104
rect 1828 6102 1829 6104
rect 2393 6102 2408 6104
rect 2408 6102 2433 6104
rect 2997 6102 3020 6104
rect 3020 6102 3037 6104
rect 3601 6102 3632 6104
rect 3632 6102 3641 6104
rect 4205 6102 4208 6104
rect 4208 6102 4244 6104
rect 4244 6102 4245 6104
rect 4809 6102 4820 6104
rect 4820 6102 4849 6104
rect 5413 6102 5432 6104
rect 5432 6102 5453 6104
rect 6017 6102 6044 6104
rect 6044 6102 6057 6104
rect 6621 6102 6624 6104
rect 6624 6102 6656 6104
rect 6656 6102 6661 6104
rect 7225 6102 7236 6104
rect 7236 6102 7265 6104
rect 7829 6102 7848 6104
rect 7848 6102 7869 6104
rect 8433 6102 8460 6104
rect 8460 6102 8473 6104
rect 9037 6102 9072 6104
rect 9072 6102 9077 6104
rect 9641 6102 9648 6104
rect 9648 6102 9681 6104
rect 10245 6102 10260 6104
rect 10260 6102 10285 6104
rect 10849 6102 10872 6104
rect 10872 6102 10889 6104
rect 11453 6102 11484 6104
rect 11484 6102 11493 6104
rect 12057 6102 12064 6104
rect 12064 6102 12096 6104
rect 12096 6102 12097 6104
rect 12661 6102 12676 6104
rect 12676 6102 12701 6104
rect 13265 6102 13288 6104
rect 13288 6102 13305 6104
rect 13869 6102 13900 6104
rect 13900 6102 13909 6104
rect 14473 6102 14476 6104
rect 14476 6102 14512 6104
rect 14512 6102 14513 6104
rect 1789 6064 1829 6102
rect 2393 6064 2433 6102
rect 2997 6064 3037 6102
rect 3601 6064 3641 6102
rect 4205 6064 4245 6102
rect 4809 6064 4849 6102
rect 5413 6064 5453 6102
rect 6017 6064 6057 6102
rect 6621 6064 6661 6102
rect 7225 6064 7265 6102
rect 7829 6064 7869 6102
rect 8433 6064 8473 6102
rect 9037 6064 9077 6102
rect 9641 6064 9681 6102
rect 10245 6064 10285 6102
rect 10849 6064 10889 6102
rect 11453 6064 11493 6102
rect 12057 6064 12097 6102
rect 12661 6064 12701 6102
rect 13265 6064 13305 6102
rect 13869 6064 13909 6102
rect 14473 6064 14513 6102
<< metal2 >>
rect 42 33420 656 33429
rect 42 33371 656 33380
rect 15344 33420 15958 33429
rect 15344 33371 15958 33380
rect 42 31420 656 31429
rect 42 31371 656 31380
rect 15344 31420 15958 31429
rect 15344 31371 15958 31380
rect 15836 29720 15958 29729
rect 42 26755 1178 26800
rect 42 26715 51 26755
rect 91 26715 149 26755
rect 189 26715 247 26755
rect 287 26715 345 26755
rect 385 26715 443 26755
rect 483 26715 541 26755
rect 581 26715 639 26755
rect 679 26715 737 26755
rect 777 26715 835 26755
rect 875 26715 933 26755
rect 973 26715 1031 26755
rect 1071 26715 1129 26755
rect 1169 26715 1178 26755
rect 42 26657 1178 26715
rect 42 26617 51 26657
rect 91 26617 149 26657
rect 189 26617 247 26657
rect 287 26617 345 26657
rect 385 26617 443 26657
rect 483 26617 541 26657
rect 581 26617 639 26657
rect 679 26617 737 26657
rect 777 26617 835 26657
rect 875 26617 933 26657
rect 973 26617 1031 26657
rect 1071 26617 1129 26657
rect 1169 26617 1178 26657
rect 42 26559 1178 26617
rect 42 26519 51 26559
rect 91 26519 149 26559
rect 189 26519 247 26559
rect 287 26519 345 26559
rect 385 26519 443 26559
rect 483 26519 541 26559
rect 581 26519 639 26559
rect 679 26519 737 26559
rect 777 26519 835 26559
rect 875 26519 933 26559
rect 973 26519 1031 26559
rect 1071 26519 1129 26559
rect 1169 26519 1178 26559
rect 42 26461 1178 26519
rect 42 26421 51 26461
rect 91 26421 149 26461
rect 189 26421 247 26461
rect 287 26421 345 26461
rect 385 26421 443 26461
rect 483 26421 541 26461
rect 581 26421 639 26461
rect 679 26421 737 26461
rect 777 26421 835 26461
rect 875 26421 933 26461
rect 973 26421 1031 26461
rect 1071 26421 1129 26461
rect 1169 26421 1178 26461
rect 42 26363 1178 26421
rect 42 26323 51 26363
rect 91 26323 149 26363
rect 189 26323 247 26363
rect 287 26323 345 26363
rect 385 26323 443 26363
rect 483 26323 541 26363
rect 581 26323 639 26363
rect 679 26323 737 26363
rect 777 26323 835 26363
rect 875 26323 933 26363
rect 973 26323 1031 26363
rect 1071 26323 1129 26363
rect 1169 26323 1178 26363
rect 42 26265 1178 26323
rect 42 26225 51 26265
rect 91 26225 149 26265
rect 189 26225 247 26265
rect 287 26225 345 26265
rect 385 26225 443 26265
rect 483 26225 541 26265
rect 581 26225 639 26265
rect 679 26225 737 26265
rect 777 26225 835 26265
rect 875 26225 933 26265
rect 973 26225 1031 26265
rect 1071 26225 1129 26265
rect 1169 26225 1178 26265
rect 42 26167 1178 26225
rect 42 26127 51 26167
rect 91 26127 149 26167
rect 189 26127 247 26167
rect 287 26127 345 26167
rect 385 26127 443 26167
rect 483 26127 541 26167
rect 581 26127 639 26167
rect 679 26127 737 26167
rect 777 26127 835 26167
rect 875 26127 933 26167
rect 973 26127 1031 26167
rect 1071 26127 1129 26167
rect 1169 26127 1178 26167
rect 42 26069 1178 26127
rect 42 26029 51 26069
rect 91 26029 149 26069
rect 189 26029 247 26069
rect 287 26029 345 26069
rect 385 26029 443 26069
rect 483 26029 541 26069
rect 581 26029 639 26069
rect 679 26029 737 26069
rect 777 26029 835 26069
rect 875 26029 933 26069
rect 973 26029 1031 26069
rect 1071 26029 1129 26069
rect 1169 26029 1178 26069
rect 42 25971 1178 26029
rect 42 25931 51 25971
rect 91 25931 149 25971
rect 189 25931 247 25971
rect 287 25931 345 25971
rect 385 25931 443 25971
rect 483 25931 541 25971
rect 581 25931 639 25971
rect 679 25931 737 25971
rect 777 25931 835 25971
rect 875 25931 933 25971
rect 973 25931 1031 25971
rect 1071 25931 1129 25971
rect 1169 25931 1178 25971
rect 42 25873 1178 25931
rect 42 25833 51 25873
rect 91 25833 149 25873
rect 189 25833 247 25873
rect 287 25833 345 25873
rect 385 25833 443 25873
rect 483 25833 541 25873
rect 581 25833 639 25873
rect 679 25833 737 25873
rect 777 25833 835 25873
rect 875 25833 933 25873
rect 973 25833 1031 25873
rect 1071 25833 1129 25873
rect 1169 25833 1178 25873
rect 42 25775 1178 25833
rect 42 25735 51 25775
rect 91 25735 149 25775
rect 189 25735 247 25775
rect 287 25735 345 25775
rect 385 25735 443 25775
rect 483 25735 541 25775
rect 581 25735 639 25775
rect 679 25735 737 25775
rect 777 25735 835 25775
rect 875 25735 933 25775
rect 973 25735 1031 25775
rect 1071 25735 1129 25775
rect 1169 25735 1178 25775
rect 42 25677 1178 25735
rect 42 25637 51 25677
rect 91 25637 149 25677
rect 189 25637 247 25677
rect 287 25637 345 25677
rect 385 25637 443 25677
rect 483 25637 541 25677
rect 581 25637 639 25677
rect 679 25637 737 25677
rect 777 25637 835 25677
rect 875 25637 933 25677
rect 973 25637 1031 25677
rect 1071 25637 1129 25677
rect 1169 25637 1178 25677
rect 42 25579 1178 25637
rect 42 25539 51 25579
rect 91 25539 149 25579
rect 189 25539 247 25579
rect 287 25539 345 25579
rect 385 25539 443 25579
rect 483 25539 541 25579
rect 581 25539 639 25579
rect 679 25539 737 25579
rect 777 25539 835 25579
rect 875 25539 933 25579
rect 973 25539 1031 25579
rect 1071 25539 1129 25579
rect 1169 25539 1178 25579
rect 42 25481 1178 25539
rect 42 25441 51 25481
rect 91 25441 149 25481
rect 189 25441 247 25481
rect 287 25441 345 25481
rect 385 25441 443 25481
rect 483 25441 541 25481
rect 581 25441 639 25481
rect 679 25441 737 25481
rect 777 25441 835 25481
rect 875 25441 933 25481
rect 973 25441 1031 25481
rect 1071 25441 1129 25481
rect 1169 25441 1178 25481
rect 42 25383 1178 25441
rect 42 25343 51 25383
rect 91 25343 149 25383
rect 189 25343 247 25383
rect 287 25343 345 25383
rect 385 25343 443 25383
rect 483 25343 541 25383
rect 581 25343 639 25383
rect 679 25343 737 25383
rect 777 25343 835 25383
rect 875 25343 933 25383
rect 973 25343 1031 25383
rect 1071 25343 1129 25383
rect 1169 25343 1178 25383
rect 42 25285 1178 25343
rect 42 25245 51 25285
rect 91 25245 149 25285
rect 189 25245 247 25285
rect 287 25245 345 25285
rect 385 25245 443 25285
rect 483 25245 541 25285
rect 581 25245 639 25285
rect 679 25245 737 25285
rect 777 25245 835 25285
rect 875 25245 933 25285
rect 973 25245 1031 25285
rect 1071 25245 1129 25285
rect 1169 25245 1178 25285
rect 42 25200 1178 25245
rect 15836 23791 15958 29680
rect 15836 23742 15958 23751
rect 3264 20071 12736 20080
rect 3264 20031 3265 20071
rect 12735 20031 12736 20071
rect 3264 20022 12736 20031
rect 84 13426 1456 19660
rect 84 6084 164 13426
rect 12370 12568 15406 19784
rect 12041 12559 15406 12568
rect 12041 12519 12064 12559
rect 15384 12519 15406 12559
rect 12041 12510 15406 12519
rect 1044 11618 3958 11627
rect 1044 11578 3836 11618
rect 1044 11569 3958 11578
rect 84 5437 973 6084
rect 1044 600 1102 11569
rect 1748 6104 1870 6113
rect 1748 6064 1789 6104
rect 1829 6064 1870 6104
rect 1748 600 1870 6064
rect 2352 6104 2474 6113
rect 2352 6064 2393 6104
rect 2433 6064 2474 6104
rect 2352 600 2474 6064
rect 2956 6104 3078 6113
rect 2956 6064 2997 6104
rect 3037 6064 3078 6104
rect 2956 600 3078 6064
rect 3560 6104 3682 6113
rect 3560 6064 3601 6104
rect 3641 6064 3682 6104
rect 3560 600 3682 6064
rect 4164 6104 4286 6113
rect 4164 6064 4205 6104
rect 4245 6064 4286 6104
rect 4164 600 4286 6064
rect 4768 6104 4890 6113
rect 4768 6064 4809 6104
rect 4849 6064 4890 6104
rect 4768 600 4890 6064
rect 5372 6104 5494 6113
rect 5372 6064 5413 6104
rect 5453 6064 5494 6104
rect 5372 600 5494 6064
rect 5976 6104 6098 6113
rect 5976 6064 6017 6104
rect 6057 6064 6098 6104
rect 5976 600 6098 6064
rect 6580 6104 6702 6113
rect 6580 6064 6621 6104
rect 6661 6064 6702 6104
rect 6580 600 6702 6064
rect 7184 6104 7306 6113
rect 7184 6064 7225 6104
rect 7265 6064 7306 6104
rect 7184 600 7306 6064
rect 7788 6104 7910 6113
rect 7788 6064 7829 6104
rect 7869 6064 7910 6104
rect 7788 600 7910 6064
rect 8392 6104 8514 6113
rect 8392 6064 8433 6104
rect 8473 6064 8514 6104
rect 8392 600 8514 6064
rect 8996 6104 9118 6113
rect 8996 6064 9037 6104
rect 9077 6064 9118 6104
rect 8996 600 9118 6064
rect 9600 6104 9722 6113
rect 9600 6064 9641 6104
rect 9681 6064 9722 6104
rect 9600 600 9722 6064
rect 10204 6104 10326 6113
rect 10204 6064 10245 6104
rect 10285 6064 10326 6104
rect 10204 600 10326 6064
rect 10808 6104 10930 6113
rect 10808 6064 10849 6104
rect 10889 6064 10930 6104
rect 10808 600 10930 6064
rect 11412 6104 11534 6113
rect 11412 6064 11453 6104
rect 11493 6064 11534 6104
rect 11412 600 11534 6064
rect 12016 6104 12138 6113
rect 12016 6064 12057 6104
rect 12097 6064 12138 6104
rect 12016 600 12138 6064
rect 12620 6104 12742 6113
rect 12620 6064 12661 6104
rect 12701 6064 12742 6104
rect 12620 600 12742 6064
rect 13224 6104 13346 6113
rect 13224 6064 13265 6104
rect 13305 6064 13346 6104
rect 13224 600 13346 6064
rect 13828 6104 13950 6113
rect 13828 6064 13869 6104
rect 13909 6064 13950 6104
rect 13828 600 13950 6064
rect 14432 6104 14554 6113
rect 14432 6064 14473 6104
rect 14513 6064 14554 6104
rect 14432 600 14554 6064
rect 1000 565 15000 600
rect 1000 525 1022 565
rect 1062 525 1120 565
rect 1160 525 1218 565
rect 1258 525 1316 565
rect 1356 525 1414 565
rect 1454 525 1512 565
rect 1552 525 1610 565
rect 1650 525 1708 565
rect 1748 525 1806 565
rect 1846 525 1904 565
rect 1944 525 2002 565
rect 2042 525 2100 565
rect 2140 525 2198 565
rect 2238 525 2296 565
rect 2336 525 2394 565
rect 2434 525 2492 565
rect 2532 525 2590 565
rect 2630 525 2688 565
rect 2728 525 2786 565
rect 2826 525 2884 565
rect 2924 525 2982 565
rect 3022 525 3080 565
rect 3120 525 3178 565
rect 3218 525 3276 565
rect 3316 525 3374 565
rect 3414 525 3472 565
rect 3512 525 3570 565
rect 3610 525 3668 565
rect 3708 525 3766 565
rect 3806 525 3864 565
rect 3904 525 3962 565
rect 4002 525 4060 565
rect 4100 525 4158 565
rect 4198 525 4256 565
rect 4296 525 4354 565
rect 4394 525 4452 565
rect 4492 525 4550 565
rect 4590 525 4648 565
rect 4688 525 4746 565
rect 4786 525 4844 565
rect 4884 525 4942 565
rect 4982 525 5040 565
rect 5080 525 5138 565
rect 5178 525 5236 565
rect 5276 525 5334 565
rect 5374 525 5432 565
rect 5472 525 5530 565
rect 5570 525 5628 565
rect 5668 525 5726 565
rect 5766 525 5824 565
rect 5864 525 5922 565
rect 5962 525 6020 565
rect 6060 525 6118 565
rect 6158 525 6216 565
rect 6256 525 6314 565
rect 6354 525 6412 565
rect 6452 525 6510 565
rect 6550 525 6608 565
rect 6648 525 6706 565
rect 6746 525 6804 565
rect 6844 525 6902 565
rect 6942 525 7000 565
rect 7040 525 7098 565
rect 7138 525 7196 565
rect 7236 525 7294 565
rect 7334 525 7392 565
rect 7432 525 7490 565
rect 7530 525 7588 565
rect 7628 525 7686 565
rect 7726 525 7784 565
rect 7824 525 7882 565
rect 7922 525 7980 565
rect 8020 525 8078 565
rect 8118 525 8176 565
rect 8216 525 8274 565
rect 8314 525 8372 565
rect 8412 525 8470 565
rect 8510 525 8568 565
rect 8608 525 8666 565
rect 8706 525 8764 565
rect 8804 525 8862 565
rect 8902 525 8960 565
rect 9000 525 9058 565
rect 9098 525 9156 565
rect 9196 525 9254 565
rect 9294 525 9352 565
rect 9392 525 9450 565
rect 9490 525 9548 565
rect 9588 525 9646 565
rect 9686 525 9744 565
rect 9784 525 9842 565
rect 9882 525 9940 565
rect 9980 525 10038 565
rect 10078 525 10136 565
rect 10176 525 10234 565
rect 10274 525 10332 565
rect 10372 525 10430 565
rect 10470 525 10528 565
rect 10568 525 10626 565
rect 10666 525 10724 565
rect 10764 525 10822 565
rect 10862 525 10920 565
rect 10960 525 11018 565
rect 11058 525 11116 565
rect 11156 525 11214 565
rect 11254 525 11312 565
rect 11352 525 11410 565
rect 11450 525 11508 565
rect 11548 525 11606 565
rect 11646 525 11704 565
rect 11744 525 11802 565
rect 11842 525 11900 565
rect 11940 525 11998 565
rect 12038 525 12096 565
rect 12136 525 12194 565
rect 12234 525 12292 565
rect 12332 525 12390 565
rect 12430 525 12488 565
rect 12528 525 12586 565
rect 12626 525 12684 565
rect 12724 525 12782 565
rect 12822 525 12880 565
rect 12920 525 12978 565
rect 13018 525 13076 565
rect 13116 525 13174 565
rect 13214 525 13272 565
rect 13312 525 13370 565
rect 13410 525 13468 565
rect 13508 525 13566 565
rect 13606 525 13664 565
rect 13704 525 13762 565
rect 13802 525 13860 565
rect 13900 525 13958 565
rect 13998 525 14056 565
rect 14096 525 14154 565
rect 14194 525 14252 565
rect 14292 525 14350 565
rect 14390 525 14448 565
rect 14488 525 14546 565
rect 14586 525 14644 565
rect 14684 525 14742 565
rect 14782 525 14840 565
rect 14880 525 14938 565
rect 14978 525 15000 565
rect 1000 467 15000 525
rect 1000 427 1022 467
rect 1062 427 1120 467
rect 1160 427 1218 467
rect 1258 427 1316 467
rect 1356 427 1414 467
rect 1454 427 1512 467
rect 1552 427 1610 467
rect 1650 427 1708 467
rect 1748 427 1806 467
rect 1846 427 1904 467
rect 1944 427 2002 467
rect 2042 427 2100 467
rect 2140 427 2198 467
rect 2238 427 2296 467
rect 2336 427 2394 467
rect 2434 427 2492 467
rect 2532 427 2590 467
rect 2630 427 2688 467
rect 2728 427 2786 467
rect 2826 427 2884 467
rect 2924 427 2982 467
rect 3022 427 3080 467
rect 3120 427 3178 467
rect 3218 427 3276 467
rect 3316 427 3374 467
rect 3414 427 3472 467
rect 3512 427 3570 467
rect 3610 427 3668 467
rect 3708 427 3766 467
rect 3806 427 3864 467
rect 3904 427 3962 467
rect 4002 427 4060 467
rect 4100 427 4158 467
rect 4198 427 4256 467
rect 4296 427 4354 467
rect 4394 427 4452 467
rect 4492 427 4550 467
rect 4590 427 4648 467
rect 4688 427 4746 467
rect 4786 427 4844 467
rect 4884 427 4942 467
rect 4982 427 5040 467
rect 5080 427 5138 467
rect 5178 427 5236 467
rect 5276 427 5334 467
rect 5374 427 5432 467
rect 5472 427 5530 467
rect 5570 427 5628 467
rect 5668 427 5726 467
rect 5766 427 5824 467
rect 5864 427 5922 467
rect 5962 427 6020 467
rect 6060 427 6118 467
rect 6158 427 6216 467
rect 6256 427 6314 467
rect 6354 427 6412 467
rect 6452 427 6510 467
rect 6550 427 6608 467
rect 6648 427 6706 467
rect 6746 427 6804 467
rect 6844 427 6902 467
rect 6942 427 7000 467
rect 7040 427 7098 467
rect 7138 427 7196 467
rect 7236 427 7294 467
rect 7334 427 7392 467
rect 7432 427 7490 467
rect 7530 427 7588 467
rect 7628 427 7686 467
rect 7726 427 7784 467
rect 7824 427 7882 467
rect 7922 427 7980 467
rect 8020 427 8078 467
rect 8118 427 8176 467
rect 8216 427 8274 467
rect 8314 427 8372 467
rect 8412 427 8470 467
rect 8510 427 8568 467
rect 8608 427 8666 467
rect 8706 427 8764 467
rect 8804 427 8862 467
rect 8902 427 8960 467
rect 9000 427 9058 467
rect 9098 427 9156 467
rect 9196 427 9254 467
rect 9294 427 9352 467
rect 9392 427 9450 467
rect 9490 427 9548 467
rect 9588 427 9646 467
rect 9686 427 9744 467
rect 9784 427 9842 467
rect 9882 427 9940 467
rect 9980 427 10038 467
rect 10078 427 10136 467
rect 10176 427 10234 467
rect 10274 427 10332 467
rect 10372 427 10430 467
rect 10470 427 10528 467
rect 10568 427 10626 467
rect 10666 427 10724 467
rect 10764 427 10822 467
rect 10862 427 10920 467
rect 10960 427 11018 467
rect 11058 427 11116 467
rect 11156 427 11214 467
rect 11254 427 11312 467
rect 11352 427 11410 467
rect 11450 427 11508 467
rect 11548 427 11606 467
rect 11646 427 11704 467
rect 11744 427 11802 467
rect 11842 427 11900 467
rect 11940 427 11998 467
rect 12038 427 12096 467
rect 12136 427 12194 467
rect 12234 427 12292 467
rect 12332 427 12390 467
rect 12430 427 12488 467
rect 12528 427 12586 467
rect 12626 427 12684 467
rect 12724 427 12782 467
rect 12822 427 12880 467
rect 12920 427 12978 467
rect 13018 427 13076 467
rect 13116 427 13174 467
rect 13214 427 13272 467
rect 13312 427 13370 467
rect 13410 427 13468 467
rect 13508 427 13566 467
rect 13606 427 13664 467
rect 13704 427 13762 467
rect 13802 427 13860 467
rect 13900 427 13958 467
rect 13998 427 14056 467
rect 14096 427 14154 467
rect 14194 427 14252 467
rect 14292 427 14350 467
rect 14390 427 14448 467
rect 14488 427 14546 467
rect 14586 427 14644 467
rect 14684 427 14742 467
rect 14782 427 14840 467
rect 14880 427 14938 467
rect 14978 427 15000 467
rect 1000 369 15000 427
rect 1000 329 1022 369
rect 1062 329 1120 369
rect 1160 329 1218 369
rect 1258 329 1316 369
rect 1356 329 1414 369
rect 1454 329 1512 369
rect 1552 329 1610 369
rect 1650 329 1708 369
rect 1748 329 1806 369
rect 1846 329 1904 369
rect 1944 329 2002 369
rect 2042 329 2100 369
rect 2140 329 2198 369
rect 2238 329 2296 369
rect 2336 329 2394 369
rect 2434 329 2492 369
rect 2532 329 2590 369
rect 2630 329 2688 369
rect 2728 329 2786 369
rect 2826 329 2884 369
rect 2924 329 2982 369
rect 3022 329 3080 369
rect 3120 329 3178 369
rect 3218 329 3276 369
rect 3316 329 3374 369
rect 3414 329 3472 369
rect 3512 329 3570 369
rect 3610 329 3668 369
rect 3708 329 3766 369
rect 3806 329 3864 369
rect 3904 329 3962 369
rect 4002 329 4060 369
rect 4100 329 4158 369
rect 4198 329 4256 369
rect 4296 329 4354 369
rect 4394 329 4452 369
rect 4492 329 4550 369
rect 4590 329 4648 369
rect 4688 329 4746 369
rect 4786 329 4844 369
rect 4884 329 4942 369
rect 4982 329 5040 369
rect 5080 329 5138 369
rect 5178 329 5236 369
rect 5276 329 5334 369
rect 5374 329 5432 369
rect 5472 329 5530 369
rect 5570 329 5628 369
rect 5668 329 5726 369
rect 5766 329 5824 369
rect 5864 329 5922 369
rect 5962 329 6020 369
rect 6060 329 6118 369
rect 6158 329 6216 369
rect 6256 329 6314 369
rect 6354 329 6412 369
rect 6452 329 6510 369
rect 6550 329 6608 369
rect 6648 329 6706 369
rect 6746 329 6804 369
rect 6844 329 6902 369
rect 6942 329 7000 369
rect 7040 329 7098 369
rect 7138 329 7196 369
rect 7236 329 7294 369
rect 7334 329 7392 369
rect 7432 329 7490 369
rect 7530 329 7588 369
rect 7628 329 7686 369
rect 7726 329 7784 369
rect 7824 329 7882 369
rect 7922 329 7980 369
rect 8020 329 8078 369
rect 8118 329 8176 369
rect 8216 329 8274 369
rect 8314 329 8372 369
rect 8412 329 8470 369
rect 8510 329 8568 369
rect 8608 329 8666 369
rect 8706 329 8764 369
rect 8804 329 8862 369
rect 8902 329 8960 369
rect 9000 329 9058 369
rect 9098 329 9156 369
rect 9196 329 9254 369
rect 9294 329 9352 369
rect 9392 329 9450 369
rect 9490 329 9548 369
rect 9588 329 9646 369
rect 9686 329 9744 369
rect 9784 329 9842 369
rect 9882 329 9940 369
rect 9980 329 10038 369
rect 10078 329 10136 369
rect 10176 329 10234 369
rect 10274 329 10332 369
rect 10372 329 10430 369
rect 10470 329 10528 369
rect 10568 329 10626 369
rect 10666 329 10724 369
rect 10764 329 10822 369
rect 10862 329 10920 369
rect 10960 329 11018 369
rect 11058 329 11116 369
rect 11156 329 11214 369
rect 11254 329 11312 369
rect 11352 329 11410 369
rect 11450 329 11508 369
rect 11548 329 11606 369
rect 11646 329 11704 369
rect 11744 329 11802 369
rect 11842 329 11900 369
rect 11940 329 11998 369
rect 12038 329 12096 369
rect 12136 329 12194 369
rect 12234 329 12292 369
rect 12332 329 12390 369
rect 12430 329 12488 369
rect 12528 329 12586 369
rect 12626 329 12684 369
rect 12724 329 12782 369
rect 12822 329 12880 369
rect 12920 329 12978 369
rect 13018 329 13076 369
rect 13116 329 13174 369
rect 13214 329 13272 369
rect 13312 329 13370 369
rect 13410 329 13468 369
rect 13508 329 13566 369
rect 13606 329 13664 369
rect 13704 329 13762 369
rect 13802 329 13860 369
rect 13900 329 13958 369
rect 13998 329 14056 369
rect 14096 329 14154 369
rect 14194 329 14252 369
rect 14292 329 14350 369
rect 14390 329 14448 369
rect 14488 329 14546 369
rect 14586 329 14644 369
rect 14684 329 14742 369
rect 14782 329 14840 369
rect 14880 329 14938 369
rect 14978 329 15000 369
rect 1000 271 15000 329
rect 1000 231 1022 271
rect 1062 231 1120 271
rect 1160 231 1218 271
rect 1258 231 1316 271
rect 1356 231 1414 271
rect 1454 231 1512 271
rect 1552 231 1610 271
rect 1650 231 1708 271
rect 1748 231 1806 271
rect 1846 231 1904 271
rect 1944 231 2002 271
rect 2042 231 2100 271
rect 2140 231 2198 271
rect 2238 231 2296 271
rect 2336 231 2394 271
rect 2434 231 2492 271
rect 2532 231 2590 271
rect 2630 231 2688 271
rect 2728 231 2786 271
rect 2826 231 2884 271
rect 2924 231 2982 271
rect 3022 231 3080 271
rect 3120 231 3178 271
rect 3218 231 3276 271
rect 3316 231 3374 271
rect 3414 231 3472 271
rect 3512 231 3570 271
rect 3610 231 3668 271
rect 3708 231 3766 271
rect 3806 231 3864 271
rect 3904 231 3962 271
rect 4002 231 4060 271
rect 4100 231 4158 271
rect 4198 231 4256 271
rect 4296 231 4354 271
rect 4394 231 4452 271
rect 4492 231 4550 271
rect 4590 231 4648 271
rect 4688 231 4746 271
rect 4786 231 4844 271
rect 4884 231 4942 271
rect 4982 231 5040 271
rect 5080 231 5138 271
rect 5178 231 5236 271
rect 5276 231 5334 271
rect 5374 231 5432 271
rect 5472 231 5530 271
rect 5570 231 5628 271
rect 5668 231 5726 271
rect 5766 231 5824 271
rect 5864 231 5922 271
rect 5962 231 6020 271
rect 6060 231 6118 271
rect 6158 231 6216 271
rect 6256 231 6314 271
rect 6354 231 6412 271
rect 6452 231 6510 271
rect 6550 231 6608 271
rect 6648 231 6706 271
rect 6746 231 6804 271
rect 6844 231 6902 271
rect 6942 231 7000 271
rect 7040 231 7098 271
rect 7138 231 7196 271
rect 7236 231 7294 271
rect 7334 231 7392 271
rect 7432 231 7490 271
rect 7530 231 7588 271
rect 7628 231 7686 271
rect 7726 231 7784 271
rect 7824 231 7882 271
rect 7922 231 7980 271
rect 8020 231 8078 271
rect 8118 231 8176 271
rect 8216 231 8274 271
rect 8314 231 8372 271
rect 8412 231 8470 271
rect 8510 231 8568 271
rect 8608 231 8666 271
rect 8706 231 8764 271
rect 8804 231 8862 271
rect 8902 231 8960 271
rect 9000 231 9058 271
rect 9098 231 9156 271
rect 9196 231 9254 271
rect 9294 231 9352 271
rect 9392 231 9450 271
rect 9490 231 9548 271
rect 9588 231 9646 271
rect 9686 231 9744 271
rect 9784 231 9842 271
rect 9882 231 9940 271
rect 9980 231 10038 271
rect 10078 231 10136 271
rect 10176 231 10234 271
rect 10274 231 10332 271
rect 10372 231 10430 271
rect 10470 231 10528 271
rect 10568 231 10626 271
rect 10666 231 10724 271
rect 10764 231 10822 271
rect 10862 231 10920 271
rect 10960 231 11018 271
rect 11058 231 11116 271
rect 11156 231 11214 271
rect 11254 231 11312 271
rect 11352 231 11410 271
rect 11450 231 11508 271
rect 11548 231 11606 271
rect 11646 231 11704 271
rect 11744 231 11802 271
rect 11842 231 11900 271
rect 11940 231 11998 271
rect 12038 231 12096 271
rect 12136 231 12194 271
rect 12234 231 12292 271
rect 12332 231 12390 271
rect 12430 231 12488 271
rect 12528 231 12586 271
rect 12626 231 12684 271
rect 12724 231 12782 271
rect 12822 231 12880 271
rect 12920 231 12978 271
rect 13018 231 13076 271
rect 13116 231 13174 271
rect 13214 231 13272 271
rect 13312 231 13370 271
rect 13410 231 13468 271
rect 13508 231 13566 271
rect 13606 231 13664 271
rect 13704 231 13762 271
rect 13802 231 13860 271
rect 13900 231 13958 271
rect 13998 231 14056 271
rect 14096 231 14154 271
rect 14194 231 14252 271
rect 14292 231 14350 271
rect 14390 231 14448 271
rect 14488 231 14546 271
rect 14586 231 14644 271
rect 14684 231 14742 271
rect 14782 231 14840 271
rect 14880 231 14938 271
rect 14978 231 15000 271
rect 1000 173 15000 231
rect 1000 133 1022 173
rect 1062 133 1120 173
rect 1160 133 1218 173
rect 1258 133 1316 173
rect 1356 133 1414 173
rect 1454 133 1512 173
rect 1552 133 1610 173
rect 1650 133 1708 173
rect 1748 133 1806 173
rect 1846 133 1904 173
rect 1944 133 2002 173
rect 2042 133 2100 173
rect 2140 133 2198 173
rect 2238 133 2296 173
rect 2336 133 2394 173
rect 2434 133 2492 173
rect 2532 133 2590 173
rect 2630 133 2688 173
rect 2728 133 2786 173
rect 2826 133 2884 173
rect 2924 133 2982 173
rect 3022 133 3080 173
rect 3120 133 3178 173
rect 3218 133 3276 173
rect 3316 133 3374 173
rect 3414 133 3472 173
rect 3512 133 3570 173
rect 3610 133 3668 173
rect 3708 133 3766 173
rect 3806 133 3864 173
rect 3904 133 3962 173
rect 4002 133 4060 173
rect 4100 133 4158 173
rect 4198 133 4256 173
rect 4296 133 4354 173
rect 4394 133 4452 173
rect 4492 133 4550 173
rect 4590 133 4648 173
rect 4688 133 4746 173
rect 4786 133 4844 173
rect 4884 133 4942 173
rect 4982 133 5040 173
rect 5080 133 5138 173
rect 5178 133 5236 173
rect 5276 133 5334 173
rect 5374 133 5432 173
rect 5472 133 5530 173
rect 5570 133 5628 173
rect 5668 133 5726 173
rect 5766 133 5824 173
rect 5864 133 5922 173
rect 5962 133 6020 173
rect 6060 133 6118 173
rect 6158 133 6216 173
rect 6256 133 6314 173
rect 6354 133 6412 173
rect 6452 133 6510 173
rect 6550 133 6608 173
rect 6648 133 6706 173
rect 6746 133 6804 173
rect 6844 133 6902 173
rect 6942 133 7000 173
rect 7040 133 7098 173
rect 7138 133 7196 173
rect 7236 133 7294 173
rect 7334 133 7392 173
rect 7432 133 7490 173
rect 7530 133 7588 173
rect 7628 133 7686 173
rect 7726 133 7784 173
rect 7824 133 7882 173
rect 7922 133 7980 173
rect 8020 133 8078 173
rect 8118 133 8176 173
rect 8216 133 8274 173
rect 8314 133 8372 173
rect 8412 133 8470 173
rect 8510 133 8568 173
rect 8608 133 8666 173
rect 8706 133 8764 173
rect 8804 133 8862 173
rect 8902 133 8960 173
rect 9000 133 9058 173
rect 9098 133 9156 173
rect 9196 133 9254 173
rect 9294 133 9352 173
rect 9392 133 9450 173
rect 9490 133 9548 173
rect 9588 133 9646 173
rect 9686 133 9744 173
rect 9784 133 9842 173
rect 9882 133 9940 173
rect 9980 133 10038 173
rect 10078 133 10136 173
rect 10176 133 10234 173
rect 10274 133 10332 173
rect 10372 133 10430 173
rect 10470 133 10528 173
rect 10568 133 10626 173
rect 10666 133 10724 173
rect 10764 133 10822 173
rect 10862 133 10920 173
rect 10960 133 11018 173
rect 11058 133 11116 173
rect 11156 133 11214 173
rect 11254 133 11312 173
rect 11352 133 11410 173
rect 11450 133 11508 173
rect 11548 133 11606 173
rect 11646 133 11704 173
rect 11744 133 11802 173
rect 11842 133 11900 173
rect 11940 133 11998 173
rect 12038 133 12096 173
rect 12136 133 12194 173
rect 12234 133 12292 173
rect 12332 133 12390 173
rect 12430 133 12488 173
rect 12528 133 12586 173
rect 12626 133 12684 173
rect 12724 133 12782 173
rect 12822 133 12880 173
rect 12920 133 12978 173
rect 13018 133 13076 173
rect 13116 133 13174 173
rect 13214 133 13272 173
rect 13312 133 13370 173
rect 13410 133 13468 173
rect 13508 133 13566 173
rect 13606 133 13664 173
rect 13704 133 13762 173
rect 13802 133 13860 173
rect 13900 133 13958 173
rect 13998 133 14056 173
rect 14096 133 14154 173
rect 14194 133 14252 173
rect 14292 133 14350 173
rect 14390 133 14448 173
rect 14488 133 14546 173
rect 14586 133 14644 173
rect 14684 133 14742 173
rect 14782 133 14840 173
rect 14880 133 14938 173
rect 14978 133 15000 173
rect 1000 75 15000 133
rect 1000 35 1022 75
rect 1062 35 1120 75
rect 1160 35 1218 75
rect 1258 35 1316 75
rect 1356 35 1414 75
rect 1454 35 1512 75
rect 1552 35 1610 75
rect 1650 35 1708 75
rect 1748 35 1806 75
rect 1846 35 1904 75
rect 1944 35 2002 75
rect 2042 35 2100 75
rect 2140 35 2198 75
rect 2238 35 2296 75
rect 2336 35 2394 75
rect 2434 35 2492 75
rect 2532 35 2590 75
rect 2630 35 2688 75
rect 2728 35 2786 75
rect 2826 35 2884 75
rect 2924 35 2982 75
rect 3022 35 3080 75
rect 3120 35 3178 75
rect 3218 35 3276 75
rect 3316 35 3374 75
rect 3414 35 3472 75
rect 3512 35 3570 75
rect 3610 35 3668 75
rect 3708 35 3766 75
rect 3806 35 3864 75
rect 3904 35 3962 75
rect 4002 35 4060 75
rect 4100 35 4158 75
rect 4198 35 4256 75
rect 4296 35 4354 75
rect 4394 35 4452 75
rect 4492 35 4550 75
rect 4590 35 4648 75
rect 4688 35 4746 75
rect 4786 35 4844 75
rect 4884 35 4942 75
rect 4982 35 5040 75
rect 5080 35 5138 75
rect 5178 35 5236 75
rect 5276 35 5334 75
rect 5374 35 5432 75
rect 5472 35 5530 75
rect 5570 35 5628 75
rect 5668 35 5726 75
rect 5766 35 5824 75
rect 5864 35 5922 75
rect 5962 35 6020 75
rect 6060 35 6118 75
rect 6158 35 6216 75
rect 6256 35 6314 75
rect 6354 35 6412 75
rect 6452 35 6510 75
rect 6550 35 6608 75
rect 6648 35 6706 75
rect 6746 35 6804 75
rect 6844 35 6902 75
rect 6942 35 7000 75
rect 7040 35 7098 75
rect 7138 35 7196 75
rect 7236 35 7294 75
rect 7334 35 7392 75
rect 7432 35 7490 75
rect 7530 35 7588 75
rect 7628 35 7686 75
rect 7726 35 7784 75
rect 7824 35 7882 75
rect 7922 35 7980 75
rect 8020 35 8078 75
rect 8118 35 8176 75
rect 8216 35 8274 75
rect 8314 35 8372 75
rect 8412 35 8470 75
rect 8510 35 8568 75
rect 8608 35 8666 75
rect 8706 35 8764 75
rect 8804 35 8862 75
rect 8902 35 8960 75
rect 9000 35 9058 75
rect 9098 35 9156 75
rect 9196 35 9254 75
rect 9294 35 9352 75
rect 9392 35 9450 75
rect 9490 35 9548 75
rect 9588 35 9646 75
rect 9686 35 9744 75
rect 9784 35 9842 75
rect 9882 35 9940 75
rect 9980 35 10038 75
rect 10078 35 10136 75
rect 10176 35 10234 75
rect 10274 35 10332 75
rect 10372 35 10430 75
rect 10470 35 10528 75
rect 10568 35 10626 75
rect 10666 35 10724 75
rect 10764 35 10822 75
rect 10862 35 10920 75
rect 10960 35 11018 75
rect 11058 35 11116 75
rect 11156 35 11214 75
rect 11254 35 11312 75
rect 11352 35 11410 75
rect 11450 35 11508 75
rect 11548 35 11606 75
rect 11646 35 11704 75
rect 11744 35 11802 75
rect 11842 35 11900 75
rect 11940 35 11998 75
rect 12038 35 12096 75
rect 12136 35 12194 75
rect 12234 35 12292 75
rect 12332 35 12390 75
rect 12430 35 12488 75
rect 12528 35 12586 75
rect 12626 35 12684 75
rect 12724 35 12782 75
rect 12822 35 12880 75
rect 12920 35 12978 75
rect 13018 35 13076 75
rect 13116 35 13174 75
rect 13214 35 13272 75
rect 13312 35 13370 75
rect 13410 35 13468 75
rect 13508 35 13566 75
rect 13606 35 13664 75
rect 13704 35 13762 75
rect 13802 35 13860 75
rect 13900 35 13958 75
rect 13998 35 14056 75
rect 14096 35 14154 75
rect 14194 35 14252 75
rect 14292 35 14350 75
rect 14390 35 14448 75
rect 14488 35 14546 75
rect 14586 35 14644 75
rect 14684 35 14742 75
rect 14782 35 14840 75
rect 14880 35 14938 75
rect 14978 35 15000 75
rect 1000 0 15000 35
<< via2 >>
rect 42 33380 656 33420
rect 15344 33380 15958 33420
rect 42 31380 656 31420
rect 15344 31380 15958 31420
rect 51 26715 91 26755
rect 149 26715 189 26755
rect 247 26715 287 26755
rect 345 26715 385 26755
rect 443 26715 483 26755
rect 541 26715 581 26755
rect 639 26715 679 26755
rect 737 26715 777 26755
rect 835 26715 875 26755
rect 933 26715 973 26755
rect 1031 26715 1071 26755
rect 1129 26715 1169 26755
rect 51 26617 91 26657
rect 149 26617 189 26657
rect 247 26617 287 26657
rect 345 26617 385 26657
rect 443 26617 483 26657
rect 541 26617 581 26657
rect 639 26617 679 26657
rect 737 26617 777 26657
rect 835 26617 875 26657
rect 933 26617 973 26657
rect 1031 26617 1071 26657
rect 1129 26617 1169 26657
rect 51 26519 91 26559
rect 149 26519 189 26559
rect 247 26519 287 26559
rect 345 26519 385 26559
rect 443 26519 483 26559
rect 541 26519 581 26559
rect 639 26519 679 26559
rect 737 26519 777 26559
rect 835 26519 875 26559
rect 933 26519 973 26559
rect 1031 26519 1071 26559
rect 1129 26519 1169 26559
rect 51 26421 91 26461
rect 149 26421 189 26461
rect 247 26421 287 26461
rect 345 26421 385 26461
rect 443 26421 483 26461
rect 541 26421 581 26461
rect 639 26421 679 26461
rect 737 26421 777 26461
rect 835 26421 875 26461
rect 933 26421 973 26461
rect 1031 26421 1071 26461
rect 1129 26421 1169 26461
rect 51 26323 91 26363
rect 149 26323 189 26363
rect 247 26323 287 26363
rect 345 26323 385 26363
rect 443 26323 483 26363
rect 541 26323 581 26363
rect 639 26323 679 26363
rect 737 26323 777 26363
rect 835 26323 875 26363
rect 933 26323 973 26363
rect 1031 26323 1071 26363
rect 1129 26323 1169 26363
rect 51 26225 91 26265
rect 149 26225 189 26265
rect 247 26225 287 26265
rect 345 26225 385 26265
rect 443 26225 483 26265
rect 541 26225 581 26265
rect 639 26225 679 26265
rect 737 26225 777 26265
rect 835 26225 875 26265
rect 933 26225 973 26265
rect 1031 26225 1071 26265
rect 1129 26225 1169 26265
rect 51 26127 91 26167
rect 149 26127 189 26167
rect 247 26127 287 26167
rect 345 26127 385 26167
rect 443 26127 483 26167
rect 541 26127 581 26167
rect 639 26127 679 26167
rect 737 26127 777 26167
rect 835 26127 875 26167
rect 933 26127 973 26167
rect 1031 26127 1071 26167
rect 1129 26127 1169 26167
rect 51 26029 91 26069
rect 149 26029 189 26069
rect 247 26029 287 26069
rect 345 26029 385 26069
rect 443 26029 483 26069
rect 541 26029 581 26069
rect 639 26029 679 26069
rect 737 26029 777 26069
rect 835 26029 875 26069
rect 933 26029 973 26069
rect 1031 26029 1071 26069
rect 1129 26029 1169 26069
rect 51 25931 91 25971
rect 149 25931 189 25971
rect 247 25931 287 25971
rect 345 25931 385 25971
rect 443 25931 483 25971
rect 541 25931 581 25971
rect 639 25931 679 25971
rect 737 25931 777 25971
rect 835 25931 875 25971
rect 933 25931 973 25971
rect 1031 25931 1071 25971
rect 1129 25931 1169 25971
rect 51 25833 91 25873
rect 149 25833 189 25873
rect 247 25833 287 25873
rect 345 25833 385 25873
rect 443 25833 483 25873
rect 541 25833 581 25873
rect 639 25833 679 25873
rect 737 25833 777 25873
rect 835 25833 875 25873
rect 933 25833 973 25873
rect 1031 25833 1071 25873
rect 1129 25833 1169 25873
rect 51 25735 91 25775
rect 149 25735 189 25775
rect 247 25735 287 25775
rect 345 25735 385 25775
rect 443 25735 483 25775
rect 541 25735 581 25775
rect 639 25735 679 25775
rect 737 25735 777 25775
rect 835 25735 875 25775
rect 933 25735 973 25775
rect 1031 25735 1071 25775
rect 1129 25735 1169 25775
rect 51 25637 91 25677
rect 149 25637 189 25677
rect 247 25637 287 25677
rect 345 25637 385 25677
rect 443 25637 483 25677
rect 541 25637 581 25677
rect 639 25637 679 25677
rect 737 25637 777 25677
rect 835 25637 875 25677
rect 933 25637 973 25677
rect 1031 25637 1071 25677
rect 1129 25637 1169 25677
rect 51 25539 91 25579
rect 149 25539 189 25579
rect 247 25539 287 25579
rect 345 25539 385 25579
rect 443 25539 483 25579
rect 541 25539 581 25579
rect 639 25539 679 25579
rect 737 25539 777 25579
rect 835 25539 875 25579
rect 933 25539 973 25579
rect 1031 25539 1071 25579
rect 1129 25539 1169 25579
rect 51 25441 91 25481
rect 149 25441 189 25481
rect 247 25441 287 25481
rect 345 25441 385 25481
rect 443 25441 483 25481
rect 541 25441 581 25481
rect 639 25441 679 25481
rect 737 25441 777 25481
rect 835 25441 875 25481
rect 933 25441 973 25481
rect 1031 25441 1071 25481
rect 1129 25441 1169 25481
rect 51 25343 91 25383
rect 149 25343 189 25383
rect 247 25343 287 25383
rect 345 25343 385 25383
rect 443 25343 483 25383
rect 541 25343 581 25383
rect 639 25343 679 25383
rect 737 25343 777 25383
rect 835 25343 875 25383
rect 933 25343 973 25383
rect 1031 25343 1071 25383
rect 1129 25343 1169 25383
rect 51 25245 91 25285
rect 149 25245 189 25285
rect 247 25245 287 25285
rect 345 25245 385 25285
rect 443 25245 483 25285
rect 541 25245 581 25285
rect 639 25245 679 25285
rect 737 25245 777 25285
rect 835 25245 875 25285
rect 933 25245 973 25285
rect 1031 25245 1071 25285
rect 1129 25245 1169 25285
rect 15836 23751 15958 23791
rect 3265 20031 3306 20071
rect 3306 20031 12694 20071
rect 12694 20031 12735 20071
rect 1022 525 1062 565
rect 1120 525 1160 565
rect 1218 525 1258 565
rect 1316 525 1356 565
rect 1414 525 1454 565
rect 1512 525 1552 565
rect 1610 525 1650 565
rect 1708 525 1748 565
rect 1806 525 1846 565
rect 1904 525 1944 565
rect 2002 525 2042 565
rect 2100 525 2140 565
rect 2198 525 2238 565
rect 2296 525 2336 565
rect 2394 525 2434 565
rect 2492 525 2532 565
rect 2590 525 2630 565
rect 2688 525 2728 565
rect 2786 525 2826 565
rect 2884 525 2924 565
rect 2982 525 3022 565
rect 3080 525 3120 565
rect 3178 525 3218 565
rect 3276 525 3316 565
rect 3374 525 3414 565
rect 3472 525 3512 565
rect 3570 525 3610 565
rect 3668 525 3708 565
rect 3766 525 3806 565
rect 3864 525 3904 565
rect 3962 525 4002 565
rect 4060 525 4100 565
rect 4158 525 4198 565
rect 4256 525 4296 565
rect 4354 525 4394 565
rect 4452 525 4492 565
rect 4550 525 4590 565
rect 4648 525 4688 565
rect 4746 525 4786 565
rect 4844 525 4884 565
rect 4942 525 4982 565
rect 5040 525 5080 565
rect 5138 525 5178 565
rect 5236 525 5276 565
rect 5334 525 5374 565
rect 5432 525 5472 565
rect 5530 525 5570 565
rect 5628 525 5668 565
rect 5726 525 5766 565
rect 5824 525 5864 565
rect 5922 525 5962 565
rect 6020 525 6060 565
rect 6118 525 6158 565
rect 6216 525 6256 565
rect 6314 525 6354 565
rect 6412 525 6452 565
rect 6510 525 6550 565
rect 6608 525 6648 565
rect 6706 525 6746 565
rect 6804 525 6844 565
rect 6902 525 6942 565
rect 7000 525 7040 565
rect 7098 525 7138 565
rect 7196 525 7236 565
rect 7294 525 7334 565
rect 7392 525 7432 565
rect 7490 525 7530 565
rect 7588 525 7628 565
rect 7686 525 7726 565
rect 7784 525 7824 565
rect 7882 525 7922 565
rect 7980 525 8020 565
rect 8078 525 8118 565
rect 8176 525 8216 565
rect 8274 525 8314 565
rect 8372 525 8412 565
rect 8470 525 8510 565
rect 8568 525 8608 565
rect 8666 525 8706 565
rect 8764 525 8804 565
rect 8862 525 8902 565
rect 8960 525 9000 565
rect 9058 525 9098 565
rect 9156 525 9196 565
rect 9254 525 9294 565
rect 9352 525 9392 565
rect 9450 525 9490 565
rect 9548 525 9588 565
rect 9646 525 9686 565
rect 9744 525 9784 565
rect 9842 525 9882 565
rect 9940 525 9980 565
rect 10038 525 10078 565
rect 10136 525 10176 565
rect 10234 525 10274 565
rect 10332 525 10372 565
rect 10430 525 10470 565
rect 10528 525 10568 565
rect 10626 525 10666 565
rect 10724 525 10764 565
rect 10822 525 10862 565
rect 10920 525 10960 565
rect 11018 525 11058 565
rect 11116 525 11156 565
rect 11214 525 11254 565
rect 11312 525 11352 565
rect 11410 525 11450 565
rect 11508 525 11548 565
rect 11606 525 11646 565
rect 11704 525 11744 565
rect 11802 525 11842 565
rect 11900 525 11940 565
rect 11998 525 12038 565
rect 12096 525 12136 565
rect 12194 525 12234 565
rect 12292 525 12332 565
rect 12390 525 12430 565
rect 12488 525 12528 565
rect 12586 525 12626 565
rect 12684 525 12724 565
rect 12782 525 12822 565
rect 12880 525 12920 565
rect 12978 525 13018 565
rect 13076 525 13116 565
rect 13174 525 13214 565
rect 13272 525 13312 565
rect 13370 525 13410 565
rect 13468 525 13508 565
rect 13566 525 13606 565
rect 13664 525 13704 565
rect 13762 525 13802 565
rect 13860 525 13900 565
rect 13958 525 13998 565
rect 14056 525 14096 565
rect 14154 525 14194 565
rect 14252 525 14292 565
rect 14350 525 14390 565
rect 14448 525 14488 565
rect 14546 525 14586 565
rect 14644 525 14684 565
rect 14742 525 14782 565
rect 14840 525 14880 565
rect 14938 525 14978 565
rect 1022 427 1062 467
rect 1120 427 1160 467
rect 1218 427 1258 467
rect 1316 427 1356 467
rect 1414 427 1454 467
rect 1512 427 1552 467
rect 1610 427 1650 467
rect 1708 427 1748 467
rect 1806 427 1846 467
rect 1904 427 1944 467
rect 2002 427 2042 467
rect 2100 427 2140 467
rect 2198 427 2238 467
rect 2296 427 2336 467
rect 2394 427 2434 467
rect 2492 427 2532 467
rect 2590 427 2630 467
rect 2688 427 2728 467
rect 2786 427 2826 467
rect 2884 427 2924 467
rect 2982 427 3022 467
rect 3080 427 3120 467
rect 3178 427 3218 467
rect 3276 427 3316 467
rect 3374 427 3414 467
rect 3472 427 3512 467
rect 3570 427 3610 467
rect 3668 427 3708 467
rect 3766 427 3806 467
rect 3864 427 3904 467
rect 3962 427 4002 467
rect 4060 427 4100 467
rect 4158 427 4198 467
rect 4256 427 4296 467
rect 4354 427 4394 467
rect 4452 427 4492 467
rect 4550 427 4590 467
rect 4648 427 4688 467
rect 4746 427 4786 467
rect 4844 427 4884 467
rect 4942 427 4982 467
rect 5040 427 5080 467
rect 5138 427 5178 467
rect 5236 427 5276 467
rect 5334 427 5374 467
rect 5432 427 5472 467
rect 5530 427 5570 467
rect 5628 427 5668 467
rect 5726 427 5766 467
rect 5824 427 5864 467
rect 5922 427 5962 467
rect 6020 427 6060 467
rect 6118 427 6158 467
rect 6216 427 6256 467
rect 6314 427 6354 467
rect 6412 427 6452 467
rect 6510 427 6550 467
rect 6608 427 6648 467
rect 6706 427 6746 467
rect 6804 427 6844 467
rect 6902 427 6942 467
rect 7000 427 7040 467
rect 7098 427 7138 467
rect 7196 427 7236 467
rect 7294 427 7334 467
rect 7392 427 7432 467
rect 7490 427 7530 467
rect 7588 427 7628 467
rect 7686 427 7726 467
rect 7784 427 7824 467
rect 7882 427 7922 467
rect 7980 427 8020 467
rect 8078 427 8118 467
rect 8176 427 8216 467
rect 8274 427 8314 467
rect 8372 427 8412 467
rect 8470 427 8510 467
rect 8568 427 8608 467
rect 8666 427 8706 467
rect 8764 427 8804 467
rect 8862 427 8902 467
rect 8960 427 9000 467
rect 9058 427 9098 467
rect 9156 427 9196 467
rect 9254 427 9294 467
rect 9352 427 9392 467
rect 9450 427 9490 467
rect 9548 427 9588 467
rect 9646 427 9686 467
rect 9744 427 9784 467
rect 9842 427 9882 467
rect 9940 427 9980 467
rect 10038 427 10078 467
rect 10136 427 10176 467
rect 10234 427 10274 467
rect 10332 427 10372 467
rect 10430 427 10470 467
rect 10528 427 10568 467
rect 10626 427 10666 467
rect 10724 427 10764 467
rect 10822 427 10862 467
rect 10920 427 10960 467
rect 11018 427 11058 467
rect 11116 427 11156 467
rect 11214 427 11254 467
rect 11312 427 11352 467
rect 11410 427 11450 467
rect 11508 427 11548 467
rect 11606 427 11646 467
rect 11704 427 11744 467
rect 11802 427 11842 467
rect 11900 427 11940 467
rect 11998 427 12038 467
rect 12096 427 12136 467
rect 12194 427 12234 467
rect 12292 427 12332 467
rect 12390 427 12430 467
rect 12488 427 12528 467
rect 12586 427 12626 467
rect 12684 427 12724 467
rect 12782 427 12822 467
rect 12880 427 12920 467
rect 12978 427 13018 467
rect 13076 427 13116 467
rect 13174 427 13214 467
rect 13272 427 13312 467
rect 13370 427 13410 467
rect 13468 427 13508 467
rect 13566 427 13606 467
rect 13664 427 13704 467
rect 13762 427 13802 467
rect 13860 427 13900 467
rect 13958 427 13998 467
rect 14056 427 14096 467
rect 14154 427 14194 467
rect 14252 427 14292 467
rect 14350 427 14390 467
rect 14448 427 14488 467
rect 14546 427 14586 467
rect 14644 427 14684 467
rect 14742 427 14782 467
rect 14840 427 14880 467
rect 14938 427 14978 467
rect 1022 329 1062 369
rect 1120 329 1160 369
rect 1218 329 1258 369
rect 1316 329 1356 369
rect 1414 329 1454 369
rect 1512 329 1552 369
rect 1610 329 1650 369
rect 1708 329 1748 369
rect 1806 329 1846 369
rect 1904 329 1944 369
rect 2002 329 2042 369
rect 2100 329 2140 369
rect 2198 329 2238 369
rect 2296 329 2336 369
rect 2394 329 2434 369
rect 2492 329 2532 369
rect 2590 329 2630 369
rect 2688 329 2728 369
rect 2786 329 2826 369
rect 2884 329 2924 369
rect 2982 329 3022 369
rect 3080 329 3120 369
rect 3178 329 3218 369
rect 3276 329 3316 369
rect 3374 329 3414 369
rect 3472 329 3512 369
rect 3570 329 3610 369
rect 3668 329 3708 369
rect 3766 329 3806 369
rect 3864 329 3904 369
rect 3962 329 4002 369
rect 4060 329 4100 369
rect 4158 329 4198 369
rect 4256 329 4296 369
rect 4354 329 4394 369
rect 4452 329 4492 369
rect 4550 329 4590 369
rect 4648 329 4688 369
rect 4746 329 4786 369
rect 4844 329 4884 369
rect 4942 329 4982 369
rect 5040 329 5080 369
rect 5138 329 5178 369
rect 5236 329 5276 369
rect 5334 329 5374 369
rect 5432 329 5472 369
rect 5530 329 5570 369
rect 5628 329 5668 369
rect 5726 329 5766 369
rect 5824 329 5864 369
rect 5922 329 5962 369
rect 6020 329 6060 369
rect 6118 329 6158 369
rect 6216 329 6256 369
rect 6314 329 6354 369
rect 6412 329 6452 369
rect 6510 329 6550 369
rect 6608 329 6648 369
rect 6706 329 6746 369
rect 6804 329 6844 369
rect 6902 329 6942 369
rect 7000 329 7040 369
rect 7098 329 7138 369
rect 7196 329 7236 369
rect 7294 329 7334 369
rect 7392 329 7432 369
rect 7490 329 7530 369
rect 7588 329 7628 369
rect 7686 329 7726 369
rect 7784 329 7824 369
rect 7882 329 7922 369
rect 7980 329 8020 369
rect 8078 329 8118 369
rect 8176 329 8216 369
rect 8274 329 8314 369
rect 8372 329 8412 369
rect 8470 329 8510 369
rect 8568 329 8608 369
rect 8666 329 8706 369
rect 8764 329 8804 369
rect 8862 329 8902 369
rect 8960 329 9000 369
rect 9058 329 9098 369
rect 9156 329 9196 369
rect 9254 329 9294 369
rect 9352 329 9392 369
rect 9450 329 9490 369
rect 9548 329 9588 369
rect 9646 329 9686 369
rect 9744 329 9784 369
rect 9842 329 9882 369
rect 9940 329 9980 369
rect 10038 329 10078 369
rect 10136 329 10176 369
rect 10234 329 10274 369
rect 10332 329 10372 369
rect 10430 329 10470 369
rect 10528 329 10568 369
rect 10626 329 10666 369
rect 10724 329 10764 369
rect 10822 329 10862 369
rect 10920 329 10960 369
rect 11018 329 11058 369
rect 11116 329 11156 369
rect 11214 329 11254 369
rect 11312 329 11352 369
rect 11410 329 11450 369
rect 11508 329 11548 369
rect 11606 329 11646 369
rect 11704 329 11744 369
rect 11802 329 11842 369
rect 11900 329 11940 369
rect 11998 329 12038 369
rect 12096 329 12136 369
rect 12194 329 12234 369
rect 12292 329 12332 369
rect 12390 329 12430 369
rect 12488 329 12528 369
rect 12586 329 12626 369
rect 12684 329 12724 369
rect 12782 329 12822 369
rect 12880 329 12920 369
rect 12978 329 13018 369
rect 13076 329 13116 369
rect 13174 329 13214 369
rect 13272 329 13312 369
rect 13370 329 13410 369
rect 13468 329 13508 369
rect 13566 329 13606 369
rect 13664 329 13704 369
rect 13762 329 13802 369
rect 13860 329 13900 369
rect 13958 329 13998 369
rect 14056 329 14096 369
rect 14154 329 14194 369
rect 14252 329 14292 369
rect 14350 329 14390 369
rect 14448 329 14488 369
rect 14546 329 14586 369
rect 14644 329 14684 369
rect 14742 329 14782 369
rect 14840 329 14880 369
rect 14938 329 14978 369
rect 1022 231 1062 271
rect 1120 231 1160 271
rect 1218 231 1258 271
rect 1316 231 1356 271
rect 1414 231 1454 271
rect 1512 231 1552 271
rect 1610 231 1650 271
rect 1708 231 1748 271
rect 1806 231 1846 271
rect 1904 231 1944 271
rect 2002 231 2042 271
rect 2100 231 2140 271
rect 2198 231 2238 271
rect 2296 231 2336 271
rect 2394 231 2434 271
rect 2492 231 2532 271
rect 2590 231 2630 271
rect 2688 231 2728 271
rect 2786 231 2826 271
rect 2884 231 2924 271
rect 2982 231 3022 271
rect 3080 231 3120 271
rect 3178 231 3218 271
rect 3276 231 3316 271
rect 3374 231 3414 271
rect 3472 231 3512 271
rect 3570 231 3610 271
rect 3668 231 3708 271
rect 3766 231 3806 271
rect 3864 231 3904 271
rect 3962 231 4002 271
rect 4060 231 4100 271
rect 4158 231 4198 271
rect 4256 231 4296 271
rect 4354 231 4394 271
rect 4452 231 4492 271
rect 4550 231 4590 271
rect 4648 231 4688 271
rect 4746 231 4786 271
rect 4844 231 4884 271
rect 4942 231 4982 271
rect 5040 231 5080 271
rect 5138 231 5178 271
rect 5236 231 5276 271
rect 5334 231 5374 271
rect 5432 231 5472 271
rect 5530 231 5570 271
rect 5628 231 5668 271
rect 5726 231 5766 271
rect 5824 231 5864 271
rect 5922 231 5962 271
rect 6020 231 6060 271
rect 6118 231 6158 271
rect 6216 231 6256 271
rect 6314 231 6354 271
rect 6412 231 6452 271
rect 6510 231 6550 271
rect 6608 231 6648 271
rect 6706 231 6746 271
rect 6804 231 6844 271
rect 6902 231 6942 271
rect 7000 231 7040 271
rect 7098 231 7138 271
rect 7196 231 7236 271
rect 7294 231 7334 271
rect 7392 231 7432 271
rect 7490 231 7530 271
rect 7588 231 7628 271
rect 7686 231 7726 271
rect 7784 231 7824 271
rect 7882 231 7922 271
rect 7980 231 8020 271
rect 8078 231 8118 271
rect 8176 231 8216 271
rect 8274 231 8314 271
rect 8372 231 8412 271
rect 8470 231 8510 271
rect 8568 231 8608 271
rect 8666 231 8706 271
rect 8764 231 8804 271
rect 8862 231 8902 271
rect 8960 231 9000 271
rect 9058 231 9098 271
rect 9156 231 9196 271
rect 9254 231 9294 271
rect 9352 231 9392 271
rect 9450 231 9490 271
rect 9548 231 9588 271
rect 9646 231 9686 271
rect 9744 231 9784 271
rect 9842 231 9882 271
rect 9940 231 9980 271
rect 10038 231 10078 271
rect 10136 231 10176 271
rect 10234 231 10274 271
rect 10332 231 10372 271
rect 10430 231 10470 271
rect 10528 231 10568 271
rect 10626 231 10666 271
rect 10724 231 10764 271
rect 10822 231 10862 271
rect 10920 231 10960 271
rect 11018 231 11058 271
rect 11116 231 11156 271
rect 11214 231 11254 271
rect 11312 231 11352 271
rect 11410 231 11450 271
rect 11508 231 11548 271
rect 11606 231 11646 271
rect 11704 231 11744 271
rect 11802 231 11842 271
rect 11900 231 11940 271
rect 11998 231 12038 271
rect 12096 231 12136 271
rect 12194 231 12234 271
rect 12292 231 12332 271
rect 12390 231 12430 271
rect 12488 231 12528 271
rect 12586 231 12626 271
rect 12684 231 12724 271
rect 12782 231 12822 271
rect 12880 231 12920 271
rect 12978 231 13018 271
rect 13076 231 13116 271
rect 13174 231 13214 271
rect 13272 231 13312 271
rect 13370 231 13410 271
rect 13468 231 13508 271
rect 13566 231 13606 271
rect 13664 231 13704 271
rect 13762 231 13802 271
rect 13860 231 13900 271
rect 13958 231 13998 271
rect 14056 231 14096 271
rect 14154 231 14194 271
rect 14252 231 14292 271
rect 14350 231 14390 271
rect 14448 231 14488 271
rect 14546 231 14586 271
rect 14644 231 14684 271
rect 14742 231 14782 271
rect 14840 231 14880 271
rect 14938 231 14978 271
rect 1022 133 1062 173
rect 1120 133 1160 173
rect 1218 133 1258 173
rect 1316 133 1356 173
rect 1414 133 1454 173
rect 1512 133 1552 173
rect 1610 133 1650 173
rect 1708 133 1748 173
rect 1806 133 1846 173
rect 1904 133 1944 173
rect 2002 133 2042 173
rect 2100 133 2140 173
rect 2198 133 2238 173
rect 2296 133 2336 173
rect 2394 133 2434 173
rect 2492 133 2532 173
rect 2590 133 2630 173
rect 2688 133 2728 173
rect 2786 133 2826 173
rect 2884 133 2924 173
rect 2982 133 3022 173
rect 3080 133 3120 173
rect 3178 133 3218 173
rect 3276 133 3316 173
rect 3374 133 3414 173
rect 3472 133 3512 173
rect 3570 133 3610 173
rect 3668 133 3708 173
rect 3766 133 3806 173
rect 3864 133 3904 173
rect 3962 133 4002 173
rect 4060 133 4100 173
rect 4158 133 4198 173
rect 4256 133 4296 173
rect 4354 133 4394 173
rect 4452 133 4492 173
rect 4550 133 4590 173
rect 4648 133 4688 173
rect 4746 133 4786 173
rect 4844 133 4884 173
rect 4942 133 4982 173
rect 5040 133 5080 173
rect 5138 133 5178 173
rect 5236 133 5276 173
rect 5334 133 5374 173
rect 5432 133 5472 173
rect 5530 133 5570 173
rect 5628 133 5668 173
rect 5726 133 5766 173
rect 5824 133 5864 173
rect 5922 133 5962 173
rect 6020 133 6060 173
rect 6118 133 6158 173
rect 6216 133 6256 173
rect 6314 133 6354 173
rect 6412 133 6452 173
rect 6510 133 6550 173
rect 6608 133 6648 173
rect 6706 133 6746 173
rect 6804 133 6844 173
rect 6902 133 6942 173
rect 7000 133 7040 173
rect 7098 133 7138 173
rect 7196 133 7236 173
rect 7294 133 7334 173
rect 7392 133 7432 173
rect 7490 133 7530 173
rect 7588 133 7628 173
rect 7686 133 7726 173
rect 7784 133 7824 173
rect 7882 133 7922 173
rect 7980 133 8020 173
rect 8078 133 8118 173
rect 8176 133 8216 173
rect 8274 133 8314 173
rect 8372 133 8412 173
rect 8470 133 8510 173
rect 8568 133 8608 173
rect 8666 133 8706 173
rect 8764 133 8804 173
rect 8862 133 8902 173
rect 8960 133 9000 173
rect 9058 133 9098 173
rect 9156 133 9196 173
rect 9254 133 9294 173
rect 9352 133 9392 173
rect 9450 133 9490 173
rect 9548 133 9588 173
rect 9646 133 9686 173
rect 9744 133 9784 173
rect 9842 133 9882 173
rect 9940 133 9980 173
rect 10038 133 10078 173
rect 10136 133 10176 173
rect 10234 133 10274 173
rect 10332 133 10372 173
rect 10430 133 10470 173
rect 10528 133 10568 173
rect 10626 133 10666 173
rect 10724 133 10764 173
rect 10822 133 10862 173
rect 10920 133 10960 173
rect 11018 133 11058 173
rect 11116 133 11156 173
rect 11214 133 11254 173
rect 11312 133 11352 173
rect 11410 133 11450 173
rect 11508 133 11548 173
rect 11606 133 11646 173
rect 11704 133 11744 173
rect 11802 133 11842 173
rect 11900 133 11940 173
rect 11998 133 12038 173
rect 12096 133 12136 173
rect 12194 133 12234 173
rect 12292 133 12332 173
rect 12390 133 12430 173
rect 12488 133 12528 173
rect 12586 133 12626 173
rect 12684 133 12724 173
rect 12782 133 12822 173
rect 12880 133 12920 173
rect 12978 133 13018 173
rect 13076 133 13116 173
rect 13174 133 13214 173
rect 13272 133 13312 173
rect 13370 133 13410 173
rect 13468 133 13508 173
rect 13566 133 13606 173
rect 13664 133 13704 173
rect 13762 133 13802 173
rect 13860 133 13900 173
rect 13958 133 13998 173
rect 14056 133 14096 173
rect 14154 133 14194 173
rect 14252 133 14292 173
rect 14350 133 14390 173
rect 14448 133 14488 173
rect 14546 133 14586 173
rect 14644 133 14684 173
rect 14742 133 14782 173
rect 14840 133 14880 173
rect 14938 133 14978 173
rect 1022 35 1062 75
rect 1120 35 1160 75
rect 1218 35 1258 75
rect 1316 35 1356 75
rect 1414 35 1454 75
rect 1512 35 1552 75
rect 1610 35 1650 75
rect 1708 35 1748 75
rect 1806 35 1846 75
rect 1904 35 1944 75
rect 2002 35 2042 75
rect 2100 35 2140 75
rect 2198 35 2238 75
rect 2296 35 2336 75
rect 2394 35 2434 75
rect 2492 35 2532 75
rect 2590 35 2630 75
rect 2688 35 2728 75
rect 2786 35 2826 75
rect 2884 35 2924 75
rect 2982 35 3022 75
rect 3080 35 3120 75
rect 3178 35 3218 75
rect 3276 35 3316 75
rect 3374 35 3414 75
rect 3472 35 3512 75
rect 3570 35 3610 75
rect 3668 35 3708 75
rect 3766 35 3806 75
rect 3864 35 3904 75
rect 3962 35 4002 75
rect 4060 35 4100 75
rect 4158 35 4198 75
rect 4256 35 4296 75
rect 4354 35 4394 75
rect 4452 35 4492 75
rect 4550 35 4590 75
rect 4648 35 4688 75
rect 4746 35 4786 75
rect 4844 35 4884 75
rect 4942 35 4982 75
rect 5040 35 5080 75
rect 5138 35 5178 75
rect 5236 35 5276 75
rect 5334 35 5374 75
rect 5432 35 5472 75
rect 5530 35 5570 75
rect 5628 35 5668 75
rect 5726 35 5766 75
rect 5824 35 5864 75
rect 5922 35 5962 75
rect 6020 35 6060 75
rect 6118 35 6158 75
rect 6216 35 6256 75
rect 6314 35 6354 75
rect 6412 35 6452 75
rect 6510 35 6550 75
rect 6608 35 6648 75
rect 6706 35 6746 75
rect 6804 35 6844 75
rect 6902 35 6942 75
rect 7000 35 7040 75
rect 7098 35 7138 75
rect 7196 35 7236 75
rect 7294 35 7334 75
rect 7392 35 7432 75
rect 7490 35 7530 75
rect 7588 35 7628 75
rect 7686 35 7726 75
rect 7784 35 7824 75
rect 7882 35 7922 75
rect 7980 35 8020 75
rect 8078 35 8118 75
rect 8176 35 8216 75
rect 8274 35 8314 75
rect 8372 35 8412 75
rect 8470 35 8510 75
rect 8568 35 8608 75
rect 8666 35 8706 75
rect 8764 35 8804 75
rect 8862 35 8902 75
rect 8960 35 9000 75
rect 9058 35 9098 75
rect 9156 35 9196 75
rect 9254 35 9294 75
rect 9352 35 9392 75
rect 9450 35 9490 75
rect 9548 35 9588 75
rect 9646 35 9686 75
rect 9744 35 9784 75
rect 9842 35 9882 75
rect 9940 35 9980 75
rect 10038 35 10078 75
rect 10136 35 10176 75
rect 10234 35 10274 75
rect 10332 35 10372 75
rect 10430 35 10470 75
rect 10528 35 10568 75
rect 10626 35 10666 75
rect 10724 35 10764 75
rect 10822 35 10862 75
rect 10920 35 10960 75
rect 11018 35 11058 75
rect 11116 35 11156 75
rect 11214 35 11254 75
rect 11312 35 11352 75
rect 11410 35 11450 75
rect 11508 35 11548 75
rect 11606 35 11646 75
rect 11704 35 11744 75
rect 11802 35 11842 75
rect 11900 35 11940 75
rect 11998 35 12038 75
rect 12096 35 12136 75
rect 12194 35 12234 75
rect 12292 35 12332 75
rect 12390 35 12430 75
rect 12488 35 12528 75
rect 12586 35 12626 75
rect 12684 35 12724 75
rect 12782 35 12822 75
rect 12880 35 12920 75
rect 12978 35 13018 75
rect 13076 35 13116 75
rect 13174 35 13214 75
rect 13272 35 13312 75
rect 13370 35 13410 75
rect 13468 35 13508 75
rect 13566 35 13606 75
rect 13664 35 13704 75
rect 13762 35 13802 75
rect 13860 35 13900 75
rect 13958 35 13998 75
rect 14056 35 14096 75
rect 14154 35 14194 75
rect 14252 35 14292 75
rect 14350 35 14390 75
rect 14448 35 14488 75
rect 14546 35 14586 75
rect 14644 35 14684 75
rect 14742 35 14782 75
rect 14840 35 14880 75
rect 14938 35 14978 75
<< metal3 >>
rect 0 33420 16000 35600
rect 0 33380 42 33420
rect 656 33380 15344 33420
rect 15958 33380 16000 33420
rect 0 32040 16000 33380
rect 0 32000 249 32040
rect 7751 32000 16000 32040
rect 0 31560 8249 31600
rect 15751 31560 16000 31600
rect 0 31420 16000 31560
rect 0 31380 42 31420
rect 656 31380 15344 31420
rect 15958 31380 16000 31420
rect 0 28000 16000 31380
rect 0 26755 16000 26800
rect 0 26715 51 26755
rect 91 26715 149 26755
rect 189 26715 247 26755
rect 287 26715 345 26755
rect 385 26715 443 26755
rect 483 26715 541 26755
rect 581 26715 639 26755
rect 679 26715 737 26755
rect 777 26715 835 26755
rect 875 26715 933 26755
rect 973 26715 1031 26755
rect 1071 26715 1129 26755
rect 1169 26715 16000 26755
rect 0 26657 16000 26715
rect 0 26617 51 26657
rect 91 26617 149 26657
rect 189 26617 247 26657
rect 287 26617 345 26657
rect 385 26617 443 26657
rect 483 26617 541 26657
rect 581 26617 639 26657
rect 679 26617 737 26657
rect 777 26617 835 26657
rect 875 26617 933 26657
rect 973 26617 1031 26657
rect 1071 26617 1129 26657
rect 1169 26617 16000 26657
rect 0 26559 16000 26617
rect 0 26519 51 26559
rect 91 26519 149 26559
rect 189 26519 247 26559
rect 287 26519 345 26559
rect 385 26519 443 26559
rect 483 26519 541 26559
rect 581 26519 639 26559
rect 679 26519 737 26559
rect 777 26519 835 26559
rect 875 26519 933 26559
rect 973 26519 1031 26559
rect 1071 26519 1129 26559
rect 1169 26519 16000 26559
rect 0 26461 16000 26519
rect 0 26421 51 26461
rect 91 26421 149 26461
rect 189 26421 247 26461
rect 287 26421 345 26461
rect 385 26421 443 26461
rect 483 26421 541 26461
rect 581 26421 639 26461
rect 679 26421 737 26461
rect 777 26421 835 26461
rect 875 26421 933 26461
rect 973 26421 1031 26461
rect 1071 26421 1129 26461
rect 1169 26421 16000 26461
rect 0 26420 16000 26421
rect 0 26380 380 26420
rect 420 26380 780 26420
rect 820 26380 1180 26420
rect 1220 26380 1580 26420
rect 1620 26380 1980 26420
rect 2020 26380 2380 26420
rect 2420 26380 2780 26420
rect 2820 26380 3180 26420
rect 3220 26380 3580 26420
rect 3620 26380 3980 26420
rect 4020 26380 4380 26420
rect 4420 26380 4780 26420
rect 4820 26380 5180 26420
rect 5220 26380 5580 26420
rect 5620 26380 5980 26420
rect 6020 26380 6380 26420
rect 6420 26380 6780 26420
rect 6820 26380 7180 26420
rect 7220 26380 7580 26420
rect 7620 26380 7980 26420
rect 8020 26380 8380 26420
rect 8420 26380 8780 26420
rect 8820 26380 9180 26420
rect 9220 26380 9580 26420
rect 9620 26380 9980 26420
rect 10020 26380 10380 26420
rect 10420 26380 10780 26420
rect 10820 26380 11180 26420
rect 11220 26380 11580 26420
rect 11620 26380 11980 26420
rect 12020 26380 12380 26420
rect 12420 26380 12780 26420
rect 12820 26380 13180 26420
rect 13220 26380 13580 26420
rect 13620 26380 13980 26420
rect 14020 26380 14380 26420
rect 14420 26380 14780 26420
rect 14820 26380 15180 26420
rect 15220 26380 15580 26420
rect 15620 26380 16000 26420
rect 0 26363 16000 26380
rect 0 26323 51 26363
rect 91 26323 149 26363
rect 189 26323 247 26363
rect 287 26323 345 26363
rect 385 26323 443 26363
rect 483 26323 541 26363
rect 581 26323 639 26363
rect 679 26323 737 26363
rect 777 26323 835 26363
rect 875 26323 933 26363
rect 973 26323 1031 26363
rect 1071 26323 1129 26363
rect 1169 26323 16000 26363
rect 0 26265 16000 26323
rect 0 26225 51 26265
rect 91 26225 149 26265
rect 189 26225 247 26265
rect 287 26225 345 26265
rect 385 26225 443 26265
rect 483 26225 541 26265
rect 581 26225 639 26265
rect 679 26225 737 26265
rect 777 26225 835 26265
rect 875 26225 933 26265
rect 973 26225 1031 26265
rect 1071 26225 1129 26265
rect 1169 26225 16000 26265
rect 0 26167 16000 26225
rect 0 26127 51 26167
rect 91 26127 149 26167
rect 189 26127 247 26167
rect 287 26127 345 26167
rect 385 26127 443 26167
rect 483 26127 541 26167
rect 581 26127 639 26167
rect 679 26127 737 26167
rect 777 26127 835 26167
rect 875 26127 933 26167
rect 973 26127 1031 26167
rect 1071 26127 1129 26167
rect 1169 26127 16000 26167
rect 0 26069 16000 26127
rect 0 26029 51 26069
rect 91 26029 149 26069
rect 189 26029 247 26069
rect 287 26029 345 26069
rect 385 26029 443 26069
rect 483 26029 541 26069
rect 581 26029 639 26069
rect 679 26029 737 26069
rect 777 26029 835 26069
rect 875 26029 933 26069
rect 973 26029 1031 26069
rect 1071 26029 1129 26069
rect 1169 26029 16000 26069
rect 0 26020 16000 26029
rect 0 25980 380 26020
rect 420 25980 780 26020
rect 820 25980 1180 26020
rect 1220 25980 1580 26020
rect 1620 25980 1980 26020
rect 2020 25980 2380 26020
rect 2420 25980 2780 26020
rect 2820 25980 3180 26020
rect 3220 25980 3580 26020
rect 3620 25980 3980 26020
rect 4020 25980 4380 26020
rect 4420 25980 4780 26020
rect 4820 25980 5180 26020
rect 5220 25980 5580 26020
rect 5620 25980 5980 26020
rect 6020 25980 6380 26020
rect 6420 25980 6780 26020
rect 6820 25980 7180 26020
rect 7220 25980 7580 26020
rect 7620 25980 7980 26020
rect 8020 25980 8380 26020
rect 8420 25980 8780 26020
rect 8820 25980 9180 26020
rect 9220 25980 9580 26020
rect 9620 25980 9980 26020
rect 10020 25980 10380 26020
rect 10420 25980 10780 26020
rect 10820 25980 11180 26020
rect 11220 25980 11580 26020
rect 11620 25980 11980 26020
rect 12020 25980 12380 26020
rect 12420 25980 12780 26020
rect 12820 25980 13180 26020
rect 13220 25980 13580 26020
rect 13620 25980 13980 26020
rect 14020 25980 14380 26020
rect 14420 25980 14780 26020
rect 14820 25980 15180 26020
rect 15220 25980 15580 26020
rect 15620 25980 16000 26020
rect 0 25971 16000 25980
rect 0 25931 51 25971
rect 91 25931 149 25971
rect 189 25931 247 25971
rect 287 25931 345 25971
rect 385 25931 443 25971
rect 483 25931 541 25971
rect 581 25931 639 25971
rect 679 25931 737 25971
rect 777 25931 835 25971
rect 875 25931 933 25971
rect 973 25931 1031 25971
rect 1071 25931 1129 25971
rect 1169 25931 16000 25971
rect 0 25873 16000 25931
rect 0 25833 51 25873
rect 91 25833 149 25873
rect 189 25833 247 25873
rect 287 25833 345 25873
rect 385 25833 443 25873
rect 483 25833 541 25873
rect 581 25833 639 25873
rect 679 25833 737 25873
rect 777 25833 835 25873
rect 875 25833 933 25873
rect 973 25833 1031 25873
rect 1071 25833 1129 25873
rect 1169 25833 16000 25873
rect 0 25775 16000 25833
rect 0 25735 51 25775
rect 91 25735 149 25775
rect 189 25735 247 25775
rect 287 25735 345 25775
rect 385 25735 443 25775
rect 483 25735 541 25775
rect 581 25735 639 25775
rect 679 25735 737 25775
rect 777 25735 835 25775
rect 875 25735 933 25775
rect 973 25735 1031 25775
rect 1071 25735 1129 25775
rect 1169 25735 16000 25775
rect 0 25677 16000 25735
rect 0 25637 51 25677
rect 91 25637 149 25677
rect 189 25637 247 25677
rect 287 25637 345 25677
rect 385 25637 443 25677
rect 483 25637 541 25677
rect 581 25637 639 25677
rect 679 25637 737 25677
rect 777 25637 835 25677
rect 875 25637 933 25677
rect 973 25637 1031 25677
rect 1071 25637 1129 25677
rect 1169 25637 16000 25677
rect 0 25620 16000 25637
rect 0 25580 380 25620
rect 420 25580 780 25620
rect 820 25580 1180 25620
rect 1220 25580 1580 25620
rect 1620 25580 1980 25620
rect 2020 25580 2380 25620
rect 2420 25580 2780 25620
rect 2820 25580 3180 25620
rect 3220 25580 3580 25620
rect 3620 25580 3980 25620
rect 4020 25580 4380 25620
rect 4420 25580 4780 25620
rect 4820 25580 5180 25620
rect 5220 25580 5580 25620
rect 5620 25580 5980 25620
rect 6020 25580 6380 25620
rect 6420 25580 6780 25620
rect 6820 25580 7180 25620
rect 7220 25580 7580 25620
rect 7620 25580 7980 25620
rect 8020 25580 8380 25620
rect 8420 25580 8780 25620
rect 8820 25580 9180 25620
rect 9220 25580 9580 25620
rect 9620 25580 9980 25620
rect 10020 25580 10380 25620
rect 10420 25580 10780 25620
rect 10820 25580 11180 25620
rect 11220 25580 11580 25620
rect 11620 25580 11980 25620
rect 12020 25580 12380 25620
rect 12420 25580 12780 25620
rect 12820 25580 13180 25620
rect 13220 25580 13580 25620
rect 13620 25580 13980 25620
rect 14020 25580 14380 25620
rect 14420 25580 14780 25620
rect 14820 25580 15180 25620
rect 15220 25580 15580 25620
rect 15620 25580 16000 25620
rect 0 25579 16000 25580
rect 0 25539 51 25579
rect 91 25539 149 25579
rect 189 25539 247 25579
rect 287 25539 345 25579
rect 385 25539 443 25579
rect 483 25539 541 25579
rect 581 25539 639 25579
rect 679 25539 737 25579
rect 777 25539 835 25579
rect 875 25539 933 25579
rect 973 25539 1031 25579
rect 1071 25539 1129 25579
rect 1169 25539 16000 25579
rect 0 25481 16000 25539
rect 0 25441 51 25481
rect 91 25441 149 25481
rect 189 25441 247 25481
rect 287 25441 345 25481
rect 385 25441 443 25481
rect 483 25441 541 25481
rect 581 25441 639 25481
rect 679 25441 737 25481
rect 777 25441 835 25481
rect 875 25441 933 25481
rect 973 25441 1031 25481
rect 1071 25441 1129 25481
rect 1169 25441 16000 25481
rect 0 25383 16000 25441
rect 0 25343 51 25383
rect 91 25343 149 25383
rect 189 25343 247 25383
rect 287 25343 345 25383
rect 385 25343 443 25383
rect 483 25343 541 25383
rect 581 25343 639 25383
rect 679 25343 737 25383
rect 777 25343 835 25383
rect 875 25343 933 25383
rect 973 25343 1031 25383
rect 1071 25343 1129 25383
rect 1169 25343 16000 25383
rect 0 25285 16000 25343
rect 0 25245 51 25285
rect 91 25245 149 25285
rect 189 25245 247 25285
rect 287 25245 345 25285
rect 385 25245 443 25285
rect 483 25245 541 25285
rect 581 25245 639 25285
rect 679 25245 737 25285
rect 777 25245 835 25285
rect 875 25245 933 25285
rect 973 25245 1031 25285
rect 1071 25245 1129 25285
rect 1169 25245 16000 25285
rect 0 25200 16000 25245
rect 0 23791 16000 23800
rect 0 23751 15836 23791
rect 15958 23751 16000 23791
rect 0 23270 16000 23751
rect 0 23230 380 23270
rect 420 23230 780 23270
rect 820 23230 1180 23270
rect 1220 23230 1580 23270
rect 1620 23230 1980 23270
rect 2020 23230 2380 23270
rect 2420 23230 2780 23270
rect 2820 23230 3180 23270
rect 3220 23230 3580 23270
rect 3620 23230 3980 23270
rect 4020 23230 4380 23270
rect 4420 23230 4780 23270
rect 4820 23230 5180 23270
rect 5220 23230 5580 23270
rect 5620 23230 5980 23270
rect 6020 23230 6380 23270
rect 6420 23230 6780 23270
rect 6820 23230 7180 23270
rect 7220 23230 7580 23270
rect 7620 23230 7980 23270
rect 8020 23230 8380 23270
rect 8420 23230 8780 23270
rect 8820 23230 9180 23270
rect 9220 23230 9580 23270
rect 9620 23230 9980 23270
rect 10020 23230 10380 23270
rect 10420 23230 10780 23270
rect 10820 23230 11180 23270
rect 11220 23230 11580 23270
rect 11620 23230 11980 23270
rect 12020 23230 12380 23270
rect 12420 23230 12780 23270
rect 12820 23230 13180 23270
rect 13220 23230 13580 23270
rect 13620 23230 13980 23270
rect 14020 23230 14380 23270
rect 14420 23230 14780 23270
rect 14820 23230 15180 23270
rect 15220 23230 15580 23270
rect 15620 23230 16000 23270
rect 0 22870 16000 23230
rect 0 22830 380 22870
rect 420 22830 780 22870
rect 820 22830 1180 22870
rect 1220 22830 1580 22870
rect 1620 22830 1980 22870
rect 2020 22830 2380 22870
rect 2420 22830 2780 22870
rect 2820 22830 3180 22870
rect 3220 22830 3580 22870
rect 3620 22830 3980 22870
rect 4020 22830 4380 22870
rect 4420 22830 4780 22870
rect 4820 22830 5180 22870
rect 5220 22830 5580 22870
rect 5620 22830 5980 22870
rect 6020 22830 6380 22870
rect 6420 22830 6780 22870
rect 6820 22830 7180 22870
rect 7220 22830 7580 22870
rect 7620 22830 7980 22870
rect 8020 22830 8380 22870
rect 8420 22830 8780 22870
rect 8820 22830 9180 22870
rect 9220 22830 9580 22870
rect 9620 22830 9980 22870
rect 10020 22830 10380 22870
rect 10420 22830 10780 22870
rect 10820 22830 11180 22870
rect 11220 22830 11580 22870
rect 11620 22830 11980 22870
rect 12020 22830 12380 22870
rect 12420 22830 12780 22870
rect 12820 22830 13180 22870
rect 13220 22830 13580 22870
rect 13620 22830 13980 22870
rect 14020 22830 14380 22870
rect 14420 22830 14780 22870
rect 14820 22830 15180 22870
rect 15220 22830 15580 22870
rect 15620 22830 16000 22870
rect 0 22470 16000 22830
rect 0 22430 380 22470
rect 420 22430 780 22470
rect 820 22430 1180 22470
rect 1220 22430 1580 22470
rect 1620 22430 1980 22470
rect 2020 22430 2380 22470
rect 2420 22430 2780 22470
rect 2820 22430 3180 22470
rect 3220 22430 3580 22470
rect 3620 22430 3980 22470
rect 4020 22430 4380 22470
rect 4420 22430 4780 22470
rect 4820 22430 5180 22470
rect 5220 22430 5580 22470
rect 5620 22430 5980 22470
rect 6020 22430 6380 22470
rect 6420 22430 6780 22470
rect 6820 22430 7180 22470
rect 7220 22430 7580 22470
rect 7620 22430 7980 22470
rect 8020 22430 8380 22470
rect 8420 22430 8780 22470
rect 8820 22430 9180 22470
rect 9220 22430 9580 22470
rect 9620 22430 9980 22470
rect 10020 22430 10380 22470
rect 10420 22430 10780 22470
rect 10820 22430 11180 22470
rect 11220 22430 11580 22470
rect 11620 22430 11980 22470
rect 12020 22430 12380 22470
rect 12420 22430 12780 22470
rect 12820 22430 13180 22470
rect 13220 22430 13580 22470
rect 13620 22430 13980 22470
rect 14020 22430 14380 22470
rect 14420 22430 14780 22470
rect 14820 22430 15180 22470
rect 15220 22430 15580 22470
rect 15620 22430 16000 22470
rect 0 22070 16000 22430
rect 0 22030 380 22070
rect 420 22030 780 22070
rect 820 22030 1180 22070
rect 1220 22030 1580 22070
rect 1620 22030 1980 22070
rect 2020 22030 2380 22070
rect 2420 22030 2780 22070
rect 2820 22030 3180 22070
rect 3220 22030 3580 22070
rect 3620 22030 3980 22070
rect 4020 22030 4380 22070
rect 4420 22030 4780 22070
rect 4820 22030 5180 22070
rect 5220 22030 5580 22070
rect 5620 22030 5980 22070
rect 6020 22030 6380 22070
rect 6420 22030 6780 22070
rect 6820 22030 7180 22070
rect 7220 22030 7580 22070
rect 7620 22030 7980 22070
rect 8020 22030 8380 22070
rect 8420 22030 8780 22070
rect 8820 22030 9180 22070
rect 9220 22030 9580 22070
rect 9620 22030 9980 22070
rect 10020 22030 10380 22070
rect 10420 22030 10780 22070
rect 10820 22030 11180 22070
rect 11220 22030 11580 22070
rect 11620 22030 11980 22070
rect 12020 22030 12380 22070
rect 12420 22030 12780 22070
rect 12820 22030 13180 22070
rect 13220 22030 13580 22070
rect 13620 22030 13980 22070
rect 14020 22030 14380 22070
rect 14420 22030 14780 22070
rect 14820 22030 15180 22070
rect 15220 22030 15580 22070
rect 15620 22030 16000 22070
rect 0 21670 16000 22030
rect 0 21630 380 21670
rect 420 21630 780 21670
rect 820 21630 1180 21670
rect 1220 21630 1580 21670
rect 1620 21630 1980 21670
rect 2020 21630 2380 21670
rect 2420 21630 2780 21670
rect 2820 21630 3180 21670
rect 3220 21630 3580 21670
rect 3620 21630 3980 21670
rect 4020 21630 4380 21670
rect 4420 21630 4780 21670
rect 4820 21630 5180 21670
rect 5220 21630 5580 21670
rect 5620 21630 5980 21670
rect 6020 21630 6380 21670
rect 6420 21630 6780 21670
rect 6820 21630 7180 21670
rect 7220 21630 7580 21670
rect 7620 21630 7980 21670
rect 8020 21630 8380 21670
rect 8420 21630 8780 21670
rect 8820 21630 9180 21670
rect 9220 21630 9580 21670
rect 9620 21630 9980 21670
rect 10020 21630 10380 21670
rect 10420 21630 10780 21670
rect 10820 21630 11180 21670
rect 11220 21630 11580 21670
rect 11620 21630 11980 21670
rect 12020 21630 12380 21670
rect 12420 21630 12780 21670
rect 12820 21630 13180 21670
rect 13220 21630 13580 21670
rect 13620 21630 13980 21670
rect 14020 21630 14380 21670
rect 14420 21630 14780 21670
rect 14820 21630 15180 21670
rect 15220 21630 15580 21670
rect 15620 21630 16000 21670
rect 0 21270 16000 21630
rect 0 21230 380 21270
rect 420 21230 780 21270
rect 820 21230 1180 21270
rect 1220 21230 1580 21270
rect 1620 21230 1980 21270
rect 2020 21230 2380 21270
rect 2420 21230 2780 21270
rect 2820 21230 3180 21270
rect 3220 21230 3580 21270
rect 3620 21230 3980 21270
rect 4020 21230 4380 21270
rect 4420 21230 4780 21270
rect 4820 21230 5180 21270
rect 5220 21230 5580 21270
rect 5620 21230 5980 21270
rect 6020 21230 6380 21270
rect 6420 21230 6780 21270
rect 6820 21230 7180 21270
rect 7220 21230 7580 21270
rect 7620 21230 7980 21270
rect 8020 21230 8380 21270
rect 8420 21230 8780 21270
rect 8820 21230 9180 21270
rect 9220 21230 9580 21270
rect 9620 21230 9980 21270
rect 10020 21230 10380 21270
rect 10420 21230 10780 21270
rect 10820 21230 11180 21270
rect 11220 21230 11580 21270
rect 11620 21230 11980 21270
rect 12020 21230 12380 21270
rect 12420 21230 12780 21270
rect 12820 21230 13180 21270
rect 13220 21230 13580 21270
rect 13620 21230 13980 21270
rect 14020 21230 14380 21270
rect 14420 21230 14780 21270
rect 14820 21230 15180 21270
rect 15220 21230 15580 21270
rect 15620 21230 16000 21270
rect 0 20870 16000 21230
rect 0 20830 380 20870
rect 420 20830 780 20870
rect 820 20830 1180 20870
rect 1220 20830 1580 20870
rect 1620 20830 1980 20870
rect 2020 20830 2380 20870
rect 2420 20830 2780 20870
rect 2820 20830 3180 20870
rect 3220 20830 3580 20870
rect 3620 20830 3980 20870
rect 4020 20830 4380 20870
rect 4420 20830 4780 20870
rect 4820 20830 5180 20870
rect 5220 20830 5580 20870
rect 5620 20830 5980 20870
rect 6020 20830 6380 20870
rect 6420 20830 6780 20870
rect 6820 20830 7180 20870
rect 7220 20830 7580 20870
rect 7620 20830 7980 20870
rect 8020 20830 8380 20870
rect 8420 20830 8780 20870
rect 8820 20830 9180 20870
rect 9220 20830 9580 20870
rect 9620 20830 9980 20870
rect 10020 20830 10380 20870
rect 10420 20830 10780 20870
rect 10820 20830 11180 20870
rect 11220 20830 11580 20870
rect 11620 20830 11980 20870
rect 12020 20830 12380 20870
rect 12420 20830 12780 20870
rect 12820 20830 13180 20870
rect 13220 20830 13580 20870
rect 13620 20830 13980 20870
rect 14020 20830 14380 20870
rect 14420 20830 14780 20870
rect 14820 20830 15180 20870
rect 15220 20830 15580 20870
rect 15620 20830 16000 20870
rect 0 20470 16000 20830
rect 0 20430 380 20470
rect 420 20430 780 20470
rect 820 20430 1180 20470
rect 1220 20430 1580 20470
rect 1620 20430 1980 20470
rect 2020 20430 2380 20470
rect 2420 20430 2780 20470
rect 2820 20430 3180 20470
rect 3220 20430 3580 20470
rect 3620 20430 3980 20470
rect 4020 20430 4380 20470
rect 4420 20430 4780 20470
rect 4820 20430 5180 20470
rect 5220 20430 5580 20470
rect 5620 20430 5980 20470
rect 6020 20430 6380 20470
rect 6420 20430 6780 20470
rect 6820 20430 7180 20470
rect 7220 20430 7580 20470
rect 7620 20430 7980 20470
rect 8020 20430 8380 20470
rect 8420 20430 8780 20470
rect 8820 20430 9180 20470
rect 9220 20430 9580 20470
rect 9620 20430 9980 20470
rect 10020 20430 10380 20470
rect 10420 20430 10780 20470
rect 10820 20430 11180 20470
rect 11220 20430 11580 20470
rect 11620 20430 11980 20470
rect 12020 20430 12380 20470
rect 12420 20430 12780 20470
rect 12820 20430 13180 20470
rect 13220 20430 13580 20470
rect 13620 20430 13980 20470
rect 14020 20430 14380 20470
rect 14420 20430 14780 20470
rect 14820 20430 15180 20470
rect 15220 20430 15580 20470
rect 15620 20430 16000 20470
rect 0 20071 16000 20430
rect 0 20070 3265 20071
rect 12735 20070 16000 20071
rect 0 20030 380 20070
rect 420 20030 780 20070
rect 820 20030 1180 20070
rect 1220 20030 1580 20070
rect 1620 20030 1980 20070
rect 2020 20030 2380 20070
rect 2420 20030 2780 20070
rect 2820 20030 3180 20070
rect 3220 20031 3265 20070
rect 12735 20031 12780 20070
rect 3220 20030 3580 20031
rect 3620 20030 3980 20031
rect 4020 20030 4380 20031
rect 4420 20030 4780 20031
rect 4820 20030 5180 20031
rect 5220 20030 5580 20031
rect 5620 20030 5980 20031
rect 6020 20030 6380 20031
rect 6420 20030 6780 20031
rect 6820 20030 7180 20031
rect 7220 20030 7580 20031
rect 7620 20030 7980 20031
rect 8020 20030 8380 20031
rect 8420 20030 8780 20031
rect 8820 20030 9180 20031
rect 9220 20030 9580 20031
rect 9620 20030 9980 20031
rect 10020 20030 10380 20031
rect 10420 20030 10780 20031
rect 10820 20030 11180 20031
rect 11220 20030 11580 20031
rect 11620 20030 11980 20031
rect 12020 20030 12380 20031
rect 12420 20030 12780 20031
rect 12820 20030 13180 20070
rect 13220 20030 13580 20070
rect 13620 20030 13980 20070
rect 14020 20030 14380 20070
rect 14420 20030 14780 20070
rect 14820 20030 15180 20070
rect 15220 20030 15580 20070
rect 15620 20030 16000 20070
rect 0 19670 16000 20030
rect 0 19630 380 19670
rect 420 19630 780 19670
rect 820 19630 1180 19670
rect 1220 19630 1580 19670
rect 1620 19630 1980 19670
rect 2020 19630 2380 19670
rect 2420 19630 2780 19670
rect 2820 19630 3180 19670
rect 3220 19630 3580 19670
rect 3620 19630 3980 19670
rect 4020 19630 4380 19670
rect 4420 19630 4780 19670
rect 4820 19630 5180 19670
rect 5220 19630 5580 19670
rect 5620 19630 5980 19670
rect 6020 19630 6380 19670
rect 6420 19630 6780 19670
rect 6820 19630 7180 19670
rect 7220 19630 7580 19670
rect 7620 19630 7980 19670
rect 8020 19630 8380 19670
rect 8420 19630 8780 19670
rect 8820 19630 9180 19670
rect 9220 19630 9580 19670
rect 9620 19630 9980 19670
rect 10020 19630 10380 19670
rect 10420 19630 10780 19670
rect 10820 19630 11180 19670
rect 11220 19630 11580 19670
rect 11620 19630 11980 19670
rect 12020 19630 12380 19670
rect 12420 19630 12780 19670
rect 12820 19630 13180 19670
rect 13220 19630 13580 19670
rect 13620 19630 13980 19670
rect 14020 19630 14380 19670
rect 14420 19630 14780 19670
rect 14820 19630 15180 19670
rect 15220 19630 15580 19670
rect 15620 19630 16000 19670
rect 0 19270 16000 19630
rect 0 19230 380 19270
rect 420 19230 780 19270
rect 820 19230 1180 19270
rect 1220 19230 1580 19270
rect 1620 19230 1980 19270
rect 2020 19230 2380 19270
rect 2420 19230 2780 19270
rect 2820 19230 3180 19270
rect 3220 19230 3580 19270
rect 3620 19230 3980 19270
rect 4020 19230 4380 19270
rect 4420 19230 4780 19270
rect 4820 19230 5180 19270
rect 5220 19230 5580 19270
rect 5620 19230 5980 19270
rect 6020 19230 6380 19270
rect 6420 19230 6780 19270
rect 6820 19230 7180 19270
rect 7220 19230 7580 19270
rect 7620 19230 7980 19270
rect 8020 19230 8380 19270
rect 8420 19230 8780 19270
rect 8820 19230 9180 19270
rect 9220 19230 9580 19270
rect 9620 19230 9980 19270
rect 10020 19230 10380 19270
rect 10420 19230 10780 19270
rect 10820 19230 11180 19270
rect 11220 19230 11580 19270
rect 11620 19230 11980 19270
rect 12020 19230 12380 19270
rect 12420 19230 12780 19270
rect 12820 19230 13180 19270
rect 13220 19230 13580 19270
rect 13620 19230 13980 19270
rect 14020 19230 14380 19270
rect 14420 19230 14780 19270
rect 14820 19230 15180 19270
rect 15220 19230 15580 19270
rect 15620 19230 16000 19270
rect 0 18700 16000 19230
rect 0 17770 16000 18300
rect 0 17730 380 17770
rect 420 17730 780 17770
rect 820 17730 1180 17770
rect 1220 17730 1580 17770
rect 1620 17730 1980 17770
rect 2020 17730 2380 17770
rect 2420 17730 2780 17770
rect 2820 17730 3180 17770
rect 3220 17730 3580 17770
rect 3620 17730 3980 17770
rect 4020 17730 4380 17770
rect 4420 17730 4780 17770
rect 4820 17730 5180 17770
rect 5220 17730 5580 17770
rect 5620 17730 5980 17770
rect 6020 17730 6380 17770
rect 6420 17730 6780 17770
rect 6820 17730 7180 17770
rect 7220 17730 7580 17770
rect 7620 17730 7980 17770
rect 8020 17730 8380 17770
rect 8420 17730 8780 17770
rect 8820 17730 9180 17770
rect 9220 17730 9580 17770
rect 9620 17730 9980 17770
rect 10020 17730 10380 17770
rect 10420 17730 10780 17770
rect 10820 17730 11180 17770
rect 11220 17730 11580 17770
rect 11620 17730 11980 17770
rect 12020 17730 12380 17770
rect 12420 17730 12780 17770
rect 12820 17730 13180 17770
rect 13220 17730 13580 17770
rect 13620 17730 13980 17770
rect 14020 17730 14380 17770
rect 14420 17730 14780 17770
rect 14820 17730 15180 17770
rect 15220 17730 15580 17770
rect 15620 17730 16000 17770
rect 0 17370 16000 17730
rect 0 17330 380 17370
rect 420 17330 780 17370
rect 820 17330 1180 17370
rect 1220 17330 1580 17370
rect 1620 17330 1980 17370
rect 2020 17330 2380 17370
rect 2420 17330 2780 17370
rect 2820 17330 3180 17370
rect 3220 17330 3580 17370
rect 3620 17330 3980 17370
rect 4020 17330 4380 17370
rect 4420 17330 4780 17370
rect 4820 17330 5180 17370
rect 5220 17330 5580 17370
rect 5620 17330 5980 17370
rect 6020 17330 6380 17370
rect 6420 17330 6780 17370
rect 6820 17330 7180 17370
rect 7220 17330 7580 17370
rect 7620 17330 7980 17370
rect 8020 17330 8380 17370
rect 8420 17330 8780 17370
rect 8820 17330 9180 17370
rect 9220 17330 9580 17370
rect 9620 17330 9980 17370
rect 10020 17330 10380 17370
rect 10420 17330 10780 17370
rect 10820 17330 11180 17370
rect 11220 17330 11580 17370
rect 11620 17330 11980 17370
rect 12020 17330 12380 17370
rect 12420 17330 12780 17370
rect 12820 17330 13180 17370
rect 13220 17330 13580 17370
rect 13620 17330 13980 17370
rect 14020 17330 14380 17370
rect 14420 17330 14780 17370
rect 14820 17330 15180 17370
rect 15220 17330 15580 17370
rect 15620 17330 16000 17370
rect 0 16970 16000 17330
rect 0 16930 380 16970
rect 420 16930 780 16970
rect 820 16930 1180 16970
rect 1220 16930 1580 16970
rect 1620 16930 1980 16970
rect 2020 16930 2380 16970
rect 2420 16930 2780 16970
rect 2820 16930 3180 16970
rect 3220 16930 3580 16970
rect 3620 16930 3980 16970
rect 4020 16930 4380 16970
rect 4420 16930 4780 16970
rect 4820 16930 5180 16970
rect 5220 16930 5580 16970
rect 5620 16930 5980 16970
rect 6020 16930 6380 16970
rect 6420 16930 6780 16970
rect 6820 16930 7180 16970
rect 7220 16930 7580 16970
rect 7620 16930 7980 16970
rect 8020 16930 8380 16970
rect 8420 16930 8780 16970
rect 8820 16930 9180 16970
rect 9220 16930 9580 16970
rect 9620 16930 9980 16970
rect 10020 16930 10380 16970
rect 10420 16930 10780 16970
rect 10820 16930 11180 16970
rect 11220 16930 11580 16970
rect 11620 16930 11980 16970
rect 12020 16930 12380 16970
rect 12420 16930 12780 16970
rect 12820 16930 13180 16970
rect 13220 16930 13580 16970
rect 13620 16930 13980 16970
rect 14020 16930 14380 16970
rect 14420 16930 14780 16970
rect 14820 16930 15180 16970
rect 15220 16930 15580 16970
rect 15620 16930 16000 16970
rect 0 16570 16000 16930
rect 0 16530 380 16570
rect 420 16530 780 16570
rect 820 16530 1180 16570
rect 1220 16530 1580 16570
rect 1620 16530 1980 16570
rect 2020 16530 2380 16570
rect 2420 16530 2780 16570
rect 2820 16530 3180 16570
rect 3220 16530 3580 16570
rect 3620 16530 3980 16570
rect 4020 16530 4380 16570
rect 4420 16530 4780 16570
rect 4820 16530 5180 16570
rect 5220 16530 5580 16570
rect 5620 16530 5980 16570
rect 6020 16530 6380 16570
rect 6420 16530 6780 16570
rect 6820 16530 7180 16570
rect 7220 16530 7580 16570
rect 7620 16530 7980 16570
rect 8020 16530 8380 16570
rect 8420 16530 8780 16570
rect 8820 16530 9180 16570
rect 9220 16530 9580 16570
rect 9620 16530 9980 16570
rect 10020 16530 10380 16570
rect 10420 16530 10780 16570
rect 10820 16530 11180 16570
rect 11220 16530 11580 16570
rect 11620 16530 11980 16570
rect 12020 16530 12380 16570
rect 12420 16530 12780 16570
rect 12820 16530 13180 16570
rect 13220 16530 13580 16570
rect 13620 16530 13980 16570
rect 14020 16530 14380 16570
rect 14420 16530 14780 16570
rect 14820 16530 15180 16570
rect 15220 16530 15580 16570
rect 15620 16530 16000 16570
rect 0 16170 16000 16530
rect 0 16130 380 16170
rect 420 16130 780 16170
rect 820 16130 1180 16170
rect 1220 16130 1580 16170
rect 1620 16130 1980 16170
rect 2020 16130 2380 16170
rect 2420 16130 2780 16170
rect 2820 16130 3180 16170
rect 3220 16130 3580 16170
rect 3620 16130 3980 16170
rect 4020 16130 4380 16170
rect 4420 16130 4780 16170
rect 4820 16130 5180 16170
rect 5220 16130 5580 16170
rect 5620 16130 5980 16170
rect 6020 16130 6380 16170
rect 6420 16130 6780 16170
rect 6820 16130 7180 16170
rect 7220 16130 7580 16170
rect 7620 16130 7980 16170
rect 8020 16130 8380 16170
rect 8420 16130 8780 16170
rect 8820 16130 9180 16170
rect 9220 16130 9580 16170
rect 9620 16130 9980 16170
rect 10020 16130 10380 16170
rect 10420 16130 10780 16170
rect 10820 16130 11180 16170
rect 11220 16130 11580 16170
rect 11620 16130 11980 16170
rect 12020 16130 12380 16170
rect 12420 16130 12780 16170
rect 12820 16130 13180 16170
rect 13220 16130 13580 16170
rect 13620 16130 13980 16170
rect 14020 16130 14380 16170
rect 14420 16130 14780 16170
rect 14820 16130 15180 16170
rect 15220 16130 15580 16170
rect 15620 16130 16000 16170
rect 0 15770 16000 16130
rect 0 15730 380 15770
rect 420 15730 780 15770
rect 820 15730 1180 15770
rect 1220 15730 1580 15770
rect 1620 15730 1980 15770
rect 2020 15730 2380 15770
rect 2420 15730 2780 15770
rect 2820 15730 3180 15770
rect 3220 15730 3580 15770
rect 3620 15730 3980 15770
rect 4020 15730 4380 15770
rect 4420 15730 4780 15770
rect 4820 15730 5180 15770
rect 5220 15730 5580 15770
rect 5620 15730 5980 15770
rect 6020 15730 6380 15770
rect 6420 15730 6780 15770
rect 6820 15730 7180 15770
rect 7220 15730 7580 15770
rect 7620 15730 7980 15770
rect 8020 15730 8380 15770
rect 8420 15730 8780 15770
rect 8820 15730 9180 15770
rect 9220 15730 9580 15770
rect 9620 15730 9980 15770
rect 10020 15730 10380 15770
rect 10420 15730 10780 15770
rect 10820 15730 11180 15770
rect 11220 15730 11580 15770
rect 11620 15730 11980 15770
rect 12020 15730 12380 15770
rect 12420 15730 12780 15770
rect 12820 15730 13180 15770
rect 13220 15730 13580 15770
rect 13620 15730 13980 15770
rect 14020 15730 14380 15770
rect 14420 15730 14780 15770
rect 14820 15730 15180 15770
rect 15220 15730 15580 15770
rect 15620 15730 16000 15770
rect 0 15370 16000 15730
rect 0 15330 380 15370
rect 420 15330 780 15370
rect 820 15330 1180 15370
rect 1220 15330 1580 15370
rect 1620 15330 1980 15370
rect 2020 15330 2380 15370
rect 2420 15330 2780 15370
rect 2820 15330 3180 15370
rect 3220 15330 3580 15370
rect 3620 15330 3980 15370
rect 4020 15330 4380 15370
rect 4420 15330 4780 15370
rect 4820 15330 5180 15370
rect 5220 15330 5580 15370
rect 5620 15330 5980 15370
rect 6020 15330 6380 15370
rect 6420 15330 6780 15370
rect 6820 15330 7180 15370
rect 7220 15330 7580 15370
rect 7620 15330 7980 15370
rect 8020 15330 8380 15370
rect 8420 15330 8780 15370
rect 8820 15330 9180 15370
rect 9220 15330 9580 15370
rect 9620 15330 9980 15370
rect 10020 15330 10380 15370
rect 10420 15330 10780 15370
rect 10820 15330 11180 15370
rect 11220 15330 11580 15370
rect 11620 15330 11980 15370
rect 12020 15330 12380 15370
rect 12420 15330 12780 15370
rect 12820 15330 13180 15370
rect 13220 15330 13580 15370
rect 13620 15330 13980 15370
rect 14020 15330 14380 15370
rect 14420 15330 14780 15370
rect 14820 15330 15180 15370
rect 15220 15330 15580 15370
rect 15620 15330 16000 15370
rect 0 14970 16000 15330
rect 0 14930 380 14970
rect 420 14930 780 14970
rect 820 14930 1180 14970
rect 1220 14930 1580 14970
rect 1620 14930 1980 14970
rect 2020 14930 2380 14970
rect 2420 14930 2780 14970
rect 2820 14930 3180 14970
rect 3220 14930 3580 14970
rect 3620 14930 3980 14970
rect 4020 14930 4380 14970
rect 4420 14930 4780 14970
rect 4820 14930 5180 14970
rect 5220 14930 5580 14970
rect 5620 14930 5980 14970
rect 6020 14930 6380 14970
rect 6420 14930 6780 14970
rect 6820 14930 7180 14970
rect 7220 14930 7580 14970
rect 7620 14930 7980 14970
rect 8020 14930 8380 14970
rect 8420 14930 8780 14970
rect 8820 14930 9180 14970
rect 9220 14930 9580 14970
rect 9620 14930 9980 14970
rect 10020 14930 10380 14970
rect 10420 14930 10780 14970
rect 10820 14930 11180 14970
rect 11220 14930 11580 14970
rect 11620 14930 11980 14970
rect 12020 14930 12380 14970
rect 12420 14930 12780 14970
rect 12820 14930 13180 14970
rect 13220 14930 13580 14970
rect 13620 14930 13980 14970
rect 14020 14930 14380 14970
rect 14420 14930 14780 14970
rect 14820 14930 15180 14970
rect 15220 14930 15580 14970
rect 15620 14930 16000 14970
rect 0 14570 16000 14930
rect 0 14530 380 14570
rect 420 14530 780 14570
rect 820 14530 1180 14570
rect 1220 14530 1580 14570
rect 1620 14530 1980 14570
rect 2020 14530 2380 14570
rect 2420 14530 2780 14570
rect 2820 14530 3180 14570
rect 3220 14530 3580 14570
rect 3620 14530 3980 14570
rect 4020 14530 4380 14570
rect 4420 14530 4780 14570
rect 4820 14530 5180 14570
rect 5220 14530 5580 14570
rect 5620 14530 5980 14570
rect 6020 14530 6380 14570
rect 6420 14530 6780 14570
rect 6820 14530 7180 14570
rect 7220 14530 7580 14570
rect 7620 14530 7980 14570
rect 8020 14530 8380 14570
rect 8420 14530 8780 14570
rect 8820 14530 9180 14570
rect 9220 14530 9580 14570
rect 9620 14530 9980 14570
rect 10020 14530 10380 14570
rect 10420 14530 10780 14570
rect 10820 14530 11180 14570
rect 11220 14530 11580 14570
rect 11620 14530 11980 14570
rect 12020 14530 12380 14570
rect 12420 14530 12780 14570
rect 12820 14530 13180 14570
rect 13220 14530 13580 14570
rect 13620 14530 13980 14570
rect 14020 14530 14380 14570
rect 14420 14530 14780 14570
rect 14820 14530 15180 14570
rect 15220 14530 15580 14570
rect 15620 14530 16000 14570
rect 0 14170 16000 14530
rect 0 14130 380 14170
rect 420 14130 780 14170
rect 820 14130 1180 14170
rect 1220 14130 1580 14170
rect 1620 14130 1980 14170
rect 2020 14130 2380 14170
rect 2420 14130 2780 14170
rect 2820 14130 3180 14170
rect 3220 14130 3580 14170
rect 3620 14130 3980 14170
rect 4020 14130 4380 14170
rect 4420 14130 4780 14170
rect 4820 14130 5180 14170
rect 5220 14130 5580 14170
rect 5620 14130 5980 14170
rect 6020 14130 6380 14170
rect 6420 14130 6780 14170
rect 6820 14130 7180 14170
rect 7220 14130 7580 14170
rect 7620 14130 7980 14170
rect 8020 14130 8380 14170
rect 8420 14130 8780 14170
rect 8820 14130 9180 14170
rect 9220 14130 9580 14170
rect 9620 14130 9980 14170
rect 10020 14130 10380 14170
rect 10420 14130 10780 14170
rect 10820 14130 11180 14170
rect 11220 14130 11580 14170
rect 11620 14130 11980 14170
rect 12020 14130 12380 14170
rect 12420 14130 12780 14170
rect 12820 14130 13180 14170
rect 13220 14130 13580 14170
rect 13620 14130 13980 14170
rect 14020 14130 14380 14170
rect 14420 14130 14780 14170
rect 14820 14130 15180 14170
rect 15220 14130 15580 14170
rect 15620 14130 16000 14170
rect 0 13770 16000 14130
rect 0 13730 380 13770
rect 420 13730 780 13770
rect 820 13730 1180 13770
rect 1220 13730 1580 13770
rect 1620 13730 1980 13770
rect 2020 13730 2380 13770
rect 2420 13730 2780 13770
rect 2820 13730 3180 13770
rect 3220 13730 3580 13770
rect 3620 13730 3980 13770
rect 4020 13730 4380 13770
rect 4420 13730 4780 13770
rect 4820 13730 5180 13770
rect 5220 13730 5580 13770
rect 5620 13730 5980 13770
rect 6020 13730 6380 13770
rect 6420 13730 6780 13770
rect 6820 13730 7180 13770
rect 7220 13730 7580 13770
rect 7620 13730 7980 13770
rect 8020 13730 8380 13770
rect 8420 13730 8780 13770
rect 8820 13730 9180 13770
rect 9220 13730 9580 13770
rect 9620 13730 9980 13770
rect 10020 13730 10380 13770
rect 10420 13730 10780 13770
rect 10820 13730 11180 13770
rect 11220 13730 11580 13770
rect 11620 13730 11980 13770
rect 12020 13730 12380 13770
rect 12420 13730 12780 13770
rect 12820 13730 13180 13770
rect 13220 13730 13580 13770
rect 13620 13730 13980 13770
rect 14020 13730 14380 13770
rect 14420 13730 14780 13770
rect 14820 13730 15180 13770
rect 15220 13730 15580 13770
rect 15620 13730 16000 13770
rect 0 13200 16000 13730
rect 0 11470 16000 12000
rect 0 11430 380 11470
rect 420 11430 780 11470
rect 820 11430 1180 11470
rect 1220 11430 1580 11470
rect 1620 11430 1980 11470
rect 2020 11430 2380 11470
rect 2420 11430 2780 11470
rect 2820 11430 3180 11470
rect 3220 11430 3580 11470
rect 3620 11430 3980 11470
rect 4020 11430 4380 11470
rect 4420 11430 4780 11470
rect 4820 11430 5180 11470
rect 5220 11430 5580 11470
rect 5620 11430 5980 11470
rect 6020 11430 6380 11470
rect 6420 11430 6780 11470
rect 6820 11430 7180 11470
rect 7220 11430 7580 11470
rect 7620 11430 7980 11470
rect 8020 11430 8380 11470
rect 8420 11430 8780 11470
rect 8820 11430 9180 11470
rect 9220 11430 9580 11470
rect 9620 11430 9980 11470
rect 10020 11430 10380 11470
rect 10420 11430 10780 11470
rect 10820 11430 11180 11470
rect 11220 11430 11580 11470
rect 11620 11430 11980 11470
rect 12020 11430 12380 11470
rect 12420 11430 12780 11470
rect 12820 11430 13180 11470
rect 13220 11430 13580 11470
rect 13620 11430 13980 11470
rect 14020 11430 14380 11470
rect 14420 11430 14780 11470
rect 14820 11430 15180 11470
rect 15220 11430 15580 11470
rect 15620 11430 16000 11470
rect 0 11070 16000 11430
rect 0 11030 380 11070
rect 420 11030 780 11070
rect 820 11030 1180 11070
rect 1220 11030 1580 11070
rect 1620 11030 1980 11070
rect 2020 11030 2380 11070
rect 2420 11030 2780 11070
rect 2820 11030 3180 11070
rect 3220 11030 3580 11070
rect 3620 11030 3980 11070
rect 4020 11030 4380 11070
rect 4420 11030 4780 11070
rect 4820 11030 5180 11070
rect 5220 11030 5580 11070
rect 5620 11030 5980 11070
rect 6020 11030 6380 11070
rect 6420 11030 6780 11070
rect 6820 11030 7180 11070
rect 7220 11030 7580 11070
rect 7620 11030 7980 11070
rect 8020 11030 8380 11070
rect 8420 11030 8780 11070
rect 8820 11030 9180 11070
rect 9220 11030 9580 11070
rect 9620 11030 9980 11070
rect 10020 11030 10380 11070
rect 10420 11030 10780 11070
rect 10820 11030 11180 11070
rect 11220 11030 11580 11070
rect 11620 11030 11980 11070
rect 12020 11030 12380 11070
rect 12420 11030 12780 11070
rect 12820 11030 13180 11070
rect 13220 11030 13580 11070
rect 13620 11030 13980 11070
rect 14020 11030 14380 11070
rect 14420 11030 14780 11070
rect 14820 11030 15180 11070
rect 15220 11030 15580 11070
rect 15620 11030 16000 11070
rect 0 10670 16000 11030
rect 0 10630 380 10670
rect 420 10630 780 10670
rect 820 10630 1180 10670
rect 1220 10630 1580 10670
rect 1620 10630 1980 10670
rect 2020 10630 2380 10670
rect 2420 10630 2780 10670
rect 2820 10630 3180 10670
rect 3220 10630 3580 10670
rect 3620 10630 3980 10670
rect 4020 10630 4380 10670
rect 4420 10630 4780 10670
rect 4820 10630 5180 10670
rect 5220 10630 5580 10670
rect 5620 10630 5980 10670
rect 6020 10630 6380 10670
rect 6420 10630 6780 10670
rect 6820 10630 7180 10670
rect 7220 10630 7580 10670
rect 7620 10630 7980 10670
rect 8020 10630 8380 10670
rect 8420 10630 8780 10670
rect 8820 10630 9180 10670
rect 9220 10630 9580 10670
rect 9620 10630 9980 10670
rect 10020 10630 10380 10670
rect 10420 10630 10780 10670
rect 10820 10630 11180 10670
rect 11220 10630 11580 10670
rect 11620 10630 11980 10670
rect 12020 10630 12380 10670
rect 12420 10630 12780 10670
rect 12820 10630 13180 10670
rect 13220 10630 13580 10670
rect 13620 10630 13980 10670
rect 14020 10630 14380 10670
rect 14420 10630 14780 10670
rect 14820 10630 15180 10670
rect 15220 10630 15580 10670
rect 15620 10630 16000 10670
rect 0 10270 16000 10630
rect 0 10230 380 10270
rect 420 10230 780 10270
rect 820 10230 1180 10270
rect 1220 10230 1580 10270
rect 1620 10230 1980 10270
rect 2020 10230 2380 10270
rect 2420 10230 2780 10270
rect 2820 10230 3180 10270
rect 3220 10230 3580 10270
rect 3620 10230 3980 10270
rect 4020 10230 4380 10270
rect 4420 10230 4780 10270
rect 4820 10230 5180 10270
rect 5220 10230 5580 10270
rect 5620 10230 5980 10270
rect 6020 10230 6380 10270
rect 6420 10230 6780 10270
rect 6820 10230 7180 10270
rect 7220 10230 7580 10270
rect 7620 10230 7980 10270
rect 8020 10230 8380 10270
rect 8420 10230 8780 10270
rect 8820 10230 9180 10270
rect 9220 10230 9580 10270
rect 9620 10230 9980 10270
rect 10020 10230 10380 10270
rect 10420 10230 10780 10270
rect 10820 10230 11180 10270
rect 11220 10230 11580 10270
rect 11620 10230 11980 10270
rect 12020 10230 12380 10270
rect 12420 10230 12780 10270
rect 12820 10230 13180 10270
rect 13220 10230 13580 10270
rect 13620 10230 13980 10270
rect 14020 10230 14380 10270
rect 14420 10230 14780 10270
rect 14820 10230 15180 10270
rect 15220 10230 15580 10270
rect 15620 10230 16000 10270
rect 0 9870 16000 10230
rect 0 9830 380 9870
rect 420 9830 780 9870
rect 820 9830 1180 9870
rect 1220 9830 1580 9870
rect 1620 9830 1980 9870
rect 2020 9830 2380 9870
rect 2420 9830 2780 9870
rect 2820 9830 3180 9870
rect 3220 9830 3580 9870
rect 3620 9830 3980 9870
rect 4020 9830 4380 9870
rect 4420 9830 4780 9870
rect 4820 9830 5180 9870
rect 5220 9830 5580 9870
rect 5620 9830 5980 9870
rect 6020 9830 6380 9870
rect 6420 9830 6780 9870
rect 6820 9830 7180 9870
rect 7220 9830 7580 9870
rect 7620 9830 7980 9870
rect 8020 9830 8380 9870
rect 8420 9830 8780 9870
rect 8820 9830 9180 9870
rect 9220 9830 9580 9870
rect 9620 9830 9980 9870
rect 10020 9830 10380 9870
rect 10420 9830 10780 9870
rect 10820 9830 11180 9870
rect 11220 9830 11580 9870
rect 11620 9830 11980 9870
rect 12020 9830 12380 9870
rect 12420 9830 12780 9870
rect 12820 9830 13180 9870
rect 13220 9830 13580 9870
rect 13620 9830 13980 9870
rect 14020 9830 14380 9870
rect 14420 9830 14780 9870
rect 14820 9830 15180 9870
rect 15220 9830 15580 9870
rect 15620 9830 16000 9870
rect 0 9470 16000 9830
rect 0 9430 380 9470
rect 420 9430 780 9470
rect 820 9430 1180 9470
rect 1220 9430 1580 9470
rect 1620 9430 1980 9470
rect 2020 9430 2380 9470
rect 2420 9430 2780 9470
rect 2820 9430 3180 9470
rect 3220 9430 3580 9470
rect 3620 9430 3980 9470
rect 4020 9430 4380 9470
rect 4420 9430 4780 9470
rect 4820 9430 5180 9470
rect 5220 9430 5580 9470
rect 5620 9430 5980 9470
rect 6020 9430 6380 9470
rect 6420 9430 6780 9470
rect 6820 9430 7180 9470
rect 7220 9430 7580 9470
rect 7620 9430 7980 9470
rect 8020 9430 8380 9470
rect 8420 9430 8780 9470
rect 8820 9430 9180 9470
rect 9220 9430 9580 9470
rect 9620 9430 9980 9470
rect 10020 9430 10380 9470
rect 10420 9430 10780 9470
rect 10820 9430 11180 9470
rect 11220 9430 11580 9470
rect 11620 9430 11980 9470
rect 12020 9430 12380 9470
rect 12420 9430 12780 9470
rect 12820 9430 13180 9470
rect 13220 9430 13580 9470
rect 13620 9430 13980 9470
rect 14020 9430 14380 9470
rect 14420 9430 14780 9470
rect 14820 9430 15180 9470
rect 15220 9430 15580 9470
rect 15620 9430 16000 9470
rect 0 9070 16000 9430
rect 0 9030 380 9070
rect 420 9030 780 9070
rect 820 9030 1180 9070
rect 1220 9030 1580 9070
rect 1620 9030 1980 9070
rect 2020 9030 2380 9070
rect 2420 9030 2780 9070
rect 2820 9030 3180 9070
rect 3220 9030 3580 9070
rect 3620 9030 3980 9070
rect 4020 9030 4380 9070
rect 4420 9030 4780 9070
rect 4820 9030 5180 9070
rect 5220 9030 5580 9070
rect 5620 9030 5980 9070
rect 6020 9030 6380 9070
rect 6420 9030 6780 9070
rect 6820 9030 7180 9070
rect 7220 9030 7580 9070
rect 7620 9030 7980 9070
rect 8020 9030 8380 9070
rect 8420 9030 8780 9070
rect 8820 9030 9180 9070
rect 9220 9030 9580 9070
rect 9620 9030 9980 9070
rect 10020 9030 10380 9070
rect 10420 9030 10780 9070
rect 10820 9030 11180 9070
rect 11220 9030 11580 9070
rect 11620 9030 11980 9070
rect 12020 9030 12380 9070
rect 12420 9030 12780 9070
rect 12820 9030 13180 9070
rect 13220 9030 13580 9070
rect 13620 9030 13980 9070
rect 14020 9030 14380 9070
rect 14420 9030 14780 9070
rect 14820 9030 15180 9070
rect 15220 9030 15580 9070
rect 15620 9030 16000 9070
rect 0 8670 16000 9030
rect 0 8630 380 8670
rect 420 8630 780 8670
rect 820 8630 1180 8670
rect 1220 8630 1580 8670
rect 1620 8630 1980 8670
rect 2020 8630 2380 8670
rect 2420 8630 2780 8670
rect 2820 8630 3180 8670
rect 3220 8630 3580 8670
rect 3620 8630 3980 8670
rect 4020 8630 4380 8670
rect 4420 8630 4780 8670
rect 4820 8630 5180 8670
rect 5220 8630 5580 8670
rect 5620 8630 5980 8670
rect 6020 8630 6380 8670
rect 6420 8630 6780 8670
rect 6820 8630 7180 8670
rect 7220 8630 7580 8670
rect 7620 8630 7980 8670
rect 8020 8630 8380 8670
rect 8420 8630 8780 8670
rect 8820 8630 9180 8670
rect 9220 8630 9580 8670
rect 9620 8630 9980 8670
rect 10020 8630 10380 8670
rect 10420 8630 10780 8670
rect 10820 8630 11180 8670
rect 11220 8630 11580 8670
rect 11620 8630 11980 8670
rect 12020 8630 12380 8670
rect 12420 8630 12780 8670
rect 12820 8630 13180 8670
rect 13220 8630 13580 8670
rect 13620 8630 13980 8670
rect 14020 8630 14380 8670
rect 14420 8630 14780 8670
rect 14820 8630 15180 8670
rect 15220 8630 15580 8670
rect 15620 8630 16000 8670
rect 0 8270 16000 8630
rect 0 8230 380 8270
rect 420 8230 780 8270
rect 820 8230 1180 8270
rect 1220 8230 1580 8270
rect 1620 8230 1980 8270
rect 2020 8230 2380 8270
rect 2420 8230 2780 8270
rect 2820 8230 3180 8270
rect 3220 8230 3580 8270
rect 3620 8230 3980 8270
rect 4020 8230 4380 8270
rect 4420 8230 4780 8270
rect 4820 8230 5180 8270
rect 5220 8230 5580 8270
rect 5620 8230 5980 8270
rect 6020 8230 6380 8270
rect 6420 8230 6780 8270
rect 6820 8230 7180 8270
rect 7220 8230 7580 8270
rect 7620 8230 7980 8270
rect 8020 8230 8380 8270
rect 8420 8230 8780 8270
rect 8820 8230 9180 8270
rect 9220 8230 9580 8270
rect 9620 8230 9980 8270
rect 10020 8230 10380 8270
rect 10420 8230 10780 8270
rect 10820 8230 11180 8270
rect 11220 8230 11580 8270
rect 11620 8230 11980 8270
rect 12020 8230 12380 8270
rect 12420 8230 12780 8270
rect 12820 8230 13180 8270
rect 13220 8230 13580 8270
rect 13620 8230 13980 8270
rect 14020 8230 14380 8270
rect 14420 8230 14780 8270
rect 14820 8230 15180 8270
rect 15220 8230 15580 8270
rect 15620 8230 16000 8270
rect 0 7870 16000 8230
rect 0 7830 380 7870
rect 420 7830 780 7870
rect 820 7830 1180 7870
rect 1220 7830 1580 7870
rect 1620 7830 1980 7870
rect 2020 7830 2380 7870
rect 2420 7830 2780 7870
rect 2820 7830 3180 7870
rect 3220 7830 3580 7870
rect 3620 7830 3980 7870
rect 4020 7830 4380 7870
rect 4420 7830 4780 7870
rect 4820 7830 5180 7870
rect 5220 7830 5580 7870
rect 5620 7830 5980 7870
rect 6020 7830 6380 7870
rect 6420 7830 6780 7870
rect 6820 7830 7180 7870
rect 7220 7830 7580 7870
rect 7620 7830 7980 7870
rect 8020 7830 8380 7870
rect 8420 7830 8780 7870
rect 8820 7830 9180 7870
rect 9220 7830 9580 7870
rect 9620 7830 9980 7870
rect 10020 7830 10380 7870
rect 10420 7830 10780 7870
rect 10820 7830 11180 7870
rect 11220 7830 11580 7870
rect 11620 7830 11980 7870
rect 12020 7830 12380 7870
rect 12420 7830 12780 7870
rect 12820 7830 13180 7870
rect 13220 7830 13580 7870
rect 13620 7830 13980 7870
rect 14020 7830 14380 7870
rect 14420 7830 14780 7870
rect 14820 7830 15180 7870
rect 15220 7830 15580 7870
rect 15620 7830 16000 7870
rect 0 7470 16000 7830
rect 0 7430 380 7470
rect 420 7430 780 7470
rect 820 7430 1180 7470
rect 1220 7430 1580 7470
rect 1620 7430 1980 7470
rect 2020 7430 2380 7470
rect 2420 7430 2780 7470
rect 2820 7430 3180 7470
rect 3220 7430 3580 7470
rect 3620 7430 3980 7470
rect 4020 7430 4380 7470
rect 4420 7430 4780 7470
rect 4820 7430 5180 7470
rect 5220 7430 5580 7470
rect 5620 7430 5980 7470
rect 6020 7430 6380 7470
rect 6420 7430 6780 7470
rect 6820 7430 7180 7470
rect 7220 7430 7580 7470
rect 7620 7430 7980 7470
rect 8020 7430 8380 7470
rect 8420 7430 8780 7470
rect 8820 7430 9180 7470
rect 9220 7430 9580 7470
rect 9620 7430 9980 7470
rect 10020 7430 10380 7470
rect 10420 7430 10780 7470
rect 10820 7430 11180 7470
rect 11220 7430 11580 7470
rect 11620 7430 11980 7470
rect 12020 7430 12380 7470
rect 12420 7430 12780 7470
rect 12820 7430 13180 7470
rect 13220 7430 13580 7470
rect 13620 7430 13980 7470
rect 14020 7430 14380 7470
rect 14420 7430 14780 7470
rect 14820 7430 15180 7470
rect 15220 7430 15580 7470
rect 15620 7430 16000 7470
rect 0 6900 16000 7430
rect 0 5970 16000 6500
rect 0 5930 380 5970
rect 420 5930 780 5970
rect 820 5930 1180 5970
rect 1220 5930 1580 5970
rect 1620 5930 1980 5970
rect 2020 5930 2380 5970
rect 2420 5930 2780 5970
rect 2820 5930 3180 5970
rect 3220 5930 3580 5970
rect 3620 5930 3980 5970
rect 4020 5930 4380 5970
rect 4420 5930 4780 5970
rect 4820 5930 5180 5970
rect 5220 5930 5580 5970
rect 5620 5930 5980 5970
rect 6020 5930 6380 5970
rect 6420 5930 6780 5970
rect 6820 5930 7180 5970
rect 7220 5930 7580 5970
rect 7620 5930 7980 5970
rect 8020 5930 8380 5970
rect 8420 5930 8780 5970
rect 8820 5930 9180 5970
rect 9220 5930 9580 5970
rect 9620 5930 9980 5970
rect 10020 5930 10380 5970
rect 10420 5930 10780 5970
rect 10820 5930 11180 5970
rect 11220 5930 11580 5970
rect 11620 5930 11980 5970
rect 12020 5930 12380 5970
rect 12420 5930 12780 5970
rect 12820 5930 13180 5970
rect 13220 5930 13580 5970
rect 13620 5930 13980 5970
rect 14020 5930 14380 5970
rect 14420 5930 14780 5970
rect 14820 5930 15180 5970
rect 15220 5930 15580 5970
rect 15620 5930 16000 5970
rect 0 5570 16000 5930
rect 0 5530 380 5570
rect 420 5530 780 5570
rect 820 5530 1180 5570
rect 1220 5530 1580 5570
rect 1620 5530 1980 5570
rect 2020 5530 2380 5570
rect 2420 5530 2780 5570
rect 2820 5530 3180 5570
rect 3220 5530 3580 5570
rect 3620 5530 3980 5570
rect 4020 5530 4380 5570
rect 4420 5530 4780 5570
rect 4820 5530 5180 5570
rect 5220 5530 5580 5570
rect 5620 5530 5980 5570
rect 6020 5530 6380 5570
rect 6420 5530 6780 5570
rect 6820 5530 7180 5570
rect 7220 5530 7580 5570
rect 7620 5530 7980 5570
rect 8020 5530 8380 5570
rect 8420 5530 8780 5570
rect 8820 5530 9180 5570
rect 9220 5530 9580 5570
rect 9620 5530 9980 5570
rect 10020 5530 10380 5570
rect 10420 5530 10780 5570
rect 10820 5530 11180 5570
rect 11220 5530 11580 5570
rect 11620 5530 11980 5570
rect 12020 5530 12380 5570
rect 12420 5530 12780 5570
rect 12820 5530 13180 5570
rect 13220 5530 13580 5570
rect 13620 5530 13980 5570
rect 14020 5530 14380 5570
rect 14420 5530 14780 5570
rect 14820 5530 15180 5570
rect 15220 5530 15580 5570
rect 15620 5530 16000 5570
rect 0 5170 16000 5530
rect 0 5130 380 5170
rect 420 5130 780 5170
rect 820 5130 1180 5170
rect 1220 5130 1580 5170
rect 1620 5130 1980 5170
rect 2020 5130 2380 5170
rect 2420 5130 2780 5170
rect 2820 5130 3180 5170
rect 3220 5130 3580 5170
rect 3620 5130 3980 5170
rect 4020 5130 4380 5170
rect 4420 5130 4780 5170
rect 4820 5130 5180 5170
rect 5220 5130 5580 5170
rect 5620 5130 5980 5170
rect 6020 5130 6380 5170
rect 6420 5130 6780 5170
rect 6820 5130 7180 5170
rect 7220 5130 7580 5170
rect 7620 5130 7980 5170
rect 8020 5130 8380 5170
rect 8420 5130 8780 5170
rect 8820 5130 9180 5170
rect 9220 5130 9580 5170
rect 9620 5130 9980 5170
rect 10020 5130 10380 5170
rect 10420 5130 10780 5170
rect 10820 5130 11180 5170
rect 11220 5130 11580 5170
rect 11620 5130 11980 5170
rect 12020 5130 12380 5170
rect 12420 5130 12780 5170
rect 12820 5130 13180 5170
rect 13220 5130 13580 5170
rect 13620 5130 13980 5170
rect 14020 5130 14380 5170
rect 14420 5130 14780 5170
rect 14820 5130 15180 5170
rect 15220 5130 15580 5170
rect 15620 5130 16000 5170
rect 0 4770 16000 5130
rect 0 4730 380 4770
rect 420 4730 780 4770
rect 820 4730 1180 4770
rect 1220 4730 1580 4770
rect 1620 4730 1980 4770
rect 2020 4730 2380 4770
rect 2420 4730 2780 4770
rect 2820 4730 3180 4770
rect 3220 4730 3580 4770
rect 3620 4730 3980 4770
rect 4020 4730 4380 4770
rect 4420 4730 4780 4770
rect 4820 4730 5180 4770
rect 5220 4730 5580 4770
rect 5620 4730 5980 4770
rect 6020 4730 6380 4770
rect 6420 4730 6780 4770
rect 6820 4730 7180 4770
rect 7220 4730 7580 4770
rect 7620 4730 7980 4770
rect 8020 4730 8380 4770
rect 8420 4730 8780 4770
rect 8820 4730 9180 4770
rect 9220 4730 9580 4770
rect 9620 4730 9980 4770
rect 10020 4730 10380 4770
rect 10420 4730 10780 4770
rect 10820 4730 11180 4770
rect 11220 4730 11580 4770
rect 11620 4730 11980 4770
rect 12020 4730 12380 4770
rect 12420 4730 12780 4770
rect 12820 4730 13180 4770
rect 13220 4730 13580 4770
rect 13620 4730 13980 4770
rect 14020 4730 14380 4770
rect 14420 4730 14780 4770
rect 14820 4730 15180 4770
rect 15220 4730 15580 4770
rect 15620 4730 16000 4770
rect 0 4370 16000 4730
rect 0 4330 380 4370
rect 420 4330 780 4370
rect 820 4330 1180 4370
rect 1220 4330 1580 4370
rect 1620 4330 1980 4370
rect 2020 4330 2380 4370
rect 2420 4330 2780 4370
rect 2820 4330 3180 4370
rect 3220 4330 3580 4370
rect 3620 4330 3980 4370
rect 4020 4330 4380 4370
rect 4420 4330 4780 4370
rect 4820 4330 5180 4370
rect 5220 4330 5580 4370
rect 5620 4330 5980 4370
rect 6020 4330 6380 4370
rect 6420 4330 6780 4370
rect 6820 4330 7180 4370
rect 7220 4330 7580 4370
rect 7620 4330 7980 4370
rect 8020 4330 8380 4370
rect 8420 4330 8780 4370
rect 8820 4330 9180 4370
rect 9220 4330 9580 4370
rect 9620 4330 9980 4370
rect 10020 4330 10380 4370
rect 10420 4330 10780 4370
rect 10820 4330 11180 4370
rect 11220 4330 11580 4370
rect 11620 4330 11980 4370
rect 12020 4330 12380 4370
rect 12420 4330 12780 4370
rect 12820 4330 13180 4370
rect 13220 4330 13580 4370
rect 13620 4330 13980 4370
rect 14020 4330 14380 4370
rect 14420 4330 14780 4370
rect 14820 4330 15180 4370
rect 15220 4330 15580 4370
rect 15620 4330 16000 4370
rect 0 3970 16000 4330
rect 0 3930 380 3970
rect 420 3930 780 3970
rect 820 3930 1180 3970
rect 1220 3930 1580 3970
rect 1620 3930 1980 3970
rect 2020 3930 2380 3970
rect 2420 3930 2780 3970
rect 2820 3930 3180 3970
rect 3220 3930 3580 3970
rect 3620 3930 3980 3970
rect 4020 3930 4380 3970
rect 4420 3930 4780 3970
rect 4820 3930 5180 3970
rect 5220 3930 5580 3970
rect 5620 3930 5980 3970
rect 6020 3930 6380 3970
rect 6420 3930 6780 3970
rect 6820 3930 7180 3970
rect 7220 3930 7580 3970
rect 7620 3930 7980 3970
rect 8020 3930 8380 3970
rect 8420 3930 8780 3970
rect 8820 3930 9180 3970
rect 9220 3930 9580 3970
rect 9620 3930 9980 3970
rect 10020 3930 10380 3970
rect 10420 3930 10780 3970
rect 10820 3930 11180 3970
rect 11220 3930 11580 3970
rect 11620 3930 11980 3970
rect 12020 3930 12380 3970
rect 12420 3930 12780 3970
rect 12820 3930 13180 3970
rect 13220 3930 13580 3970
rect 13620 3930 13980 3970
rect 14020 3930 14380 3970
rect 14420 3930 14780 3970
rect 14820 3930 15180 3970
rect 15220 3930 15580 3970
rect 15620 3930 16000 3970
rect 0 3570 16000 3930
rect 0 3530 380 3570
rect 420 3530 780 3570
rect 820 3530 1180 3570
rect 1220 3530 1580 3570
rect 1620 3530 1980 3570
rect 2020 3530 2380 3570
rect 2420 3530 2780 3570
rect 2820 3530 3180 3570
rect 3220 3530 3580 3570
rect 3620 3530 3980 3570
rect 4020 3530 4380 3570
rect 4420 3530 4780 3570
rect 4820 3530 5180 3570
rect 5220 3530 5580 3570
rect 5620 3530 5980 3570
rect 6020 3530 6380 3570
rect 6420 3530 6780 3570
rect 6820 3530 7180 3570
rect 7220 3530 7580 3570
rect 7620 3530 7980 3570
rect 8020 3530 8380 3570
rect 8420 3530 8780 3570
rect 8820 3530 9180 3570
rect 9220 3530 9580 3570
rect 9620 3530 9980 3570
rect 10020 3530 10380 3570
rect 10420 3530 10780 3570
rect 10820 3530 11180 3570
rect 11220 3530 11580 3570
rect 11620 3530 11980 3570
rect 12020 3530 12380 3570
rect 12420 3530 12780 3570
rect 12820 3530 13180 3570
rect 13220 3530 13580 3570
rect 13620 3530 13980 3570
rect 14020 3530 14380 3570
rect 14420 3530 14780 3570
rect 14820 3530 15180 3570
rect 15220 3530 15580 3570
rect 15620 3530 16000 3570
rect 0 3170 16000 3530
rect 0 3130 380 3170
rect 420 3130 780 3170
rect 820 3130 1180 3170
rect 1220 3130 1580 3170
rect 1620 3130 1980 3170
rect 2020 3130 2380 3170
rect 2420 3130 2780 3170
rect 2820 3130 3180 3170
rect 3220 3130 3580 3170
rect 3620 3130 3980 3170
rect 4020 3130 4380 3170
rect 4420 3130 4780 3170
rect 4820 3130 5180 3170
rect 5220 3130 5580 3170
rect 5620 3130 5980 3170
rect 6020 3130 6380 3170
rect 6420 3130 6780 3170
rect 6820 3130 7180 3170
rect 7220 3130 7580 3170
rect 7620 3130 7980 3170
rect 8020 3130 8380 3170
rect 8420 3130 8780 3170
rect 8820 3130 9180 3170
rect 9220 3130 9580 3170
rect 9620 3130 9980 3170
rect 10020 3130 10380 3170
rect 10420 3130 10780 3170
rect 10820 3130 11180 3170
rect 11220 3130 11580 3170
rect 11620 3130 11980 3170
rect 12020 3130 12380 3170
rect 12420 3130 12780 3170
rect 12820 3130 13180 3170
rect 13220 3130 13580 3170
rect 13620 3130 13980 3170
rect 14020 3130 14380 3170
rect 14420 3130 14780 3170
rect 14820 3130 15180 3170
rect 15220 3130 15580 3170
rect 15620 3130 16000 3170
rect 0 2770 16000 3130
rect 0 2730 380 2770
rect 420 2730 780 2770
rect 820 2730 1180 2770
rect 1220 2730 1580 2770
rect 1620 2730 1980 2770
rect 2020 2730 2380 2770
rect 2420 2730 2780 2770
rect 2820 2730 3180 2770
rect 3220 2730 3580 2770
rect 3620 2730 3980 2770
rect 4020 2730 4380 2770
rect 4420 2730 4780 2770
rect 4820 2730 5180 2770
rect 5220 2730 5580 2770
rect 5620 2730 5980 2770
rect 6020 2730 6380 2770
rect 6420 2730 6780 2770
rect 6820 2730 7180 2770
rect 7220 2730 7580 2770
rect 7620 2730 7980 2770
rect 8020 2730 8380 2770
rect 8420 2730 8780 2770
rect 8820 2730 9180 2770
rect 9220 2730 9580 2770
rect 9620 2730 9980 2770
rect 10020 2730 10380 2770
rect 10420 2730 10780 2770
rect 10820 2730 11180 2770
rect 11220 2730 11580 2770
rect 11620 2730 11980 2770
rect 12020 2730 12380 2770
rect 12420 2730 12780 2770
rect 12820 2730 13180 2770
rect 13220 2730 13580 2770
rect 13620 2730 13980 2770
rect 14020 2730 14380 2770
rect 14420 2730 14780 2770
rect 14820 2730 15180 2770
rect 15220 2730 15580 2770
rect 15620 2730 16000 2770
rect 0 2370 16000 2730
rect 0 2330 380 2370
rect 420 2330 780 2370
rect 820 2330 1180 2370
rect 1220 2330 1580 2370
rect 1620 2330 1980 2370
rect 2020 2330 2380 2370
rect 2420 2330 2780 2370
rect 2820 2330 3180 2370
rect 3220 2330 3580 2370
rect 3620 2330 3980 2370
rect 4020 2330 4380 2370
rect 4420 2330 4780 2370
rect 4820 2330 5180 2370
rect 5220 2330 5580 2370
rect 5620 2330 5980 2370
rect 6020 2330 6380 2370
rect 6420 2330 6780 2370
rect 6820 2330 7180 2370
rect 7220 2330 7580 2370
rect 7620 2330 7980 2370
rect 8020 2330 8380 2370
rect 8420 2330 8780 2370
rect 8820 2330 9180 2370
rect 9220 2330 9580 2370
rect 9620 2330 9980 2370
rect 10020 2330 10380 2370
rect 10420 2330 10780 2370
rect 10820 2330 11180 2370
rect 11220 2330 11580 2370
rect 11620 2330 11980 2370
rect 12020 2330 12380 2370
rect 12420 2330 12780 2370
rect 12820 2330 13180 2370
rect 13220 2330 13580 2370
rect 13620 2330 13980 2370
rect 14020 2330 14380 2370
rect 14420 2330 14780 2370
rect 14820 2330 15180 2370
rect 15220 2330 15580 2370
rect 15620 2330 16000 2370
rect 0 1970 16000 2330
rect 0 1930 380 1970
rect 420 1930 780 1970
rect 820 1930 1180 1970
rect 1220 1930 1580 1970
rect 1620 1930 1980 1970
rect 2020 1930 2380 1970
rect 2420 1930 2780 1970
rect 2820 1930 3180 1970
rect 3220 1930 3580 1970
rect 3620 1930 3980 1970
rect 4020 1930 4380 1970
rect 4420 1930 4780 1970
rect 4820 1930 5180 1970
rect 5220 1930 5580 1970
rect 5620 1930 5980 1970
rect 6020 1930 6380 1970
rect 6420 1930 6780 1970
rect 6820 1930 7180 1970
rect 7220 1930 7580 1970
rect 7620 1930 7980 1970
rect 8020 1930 8380 1970
rect 8420 1930 8780 1970
rect 8820 1930 9180 1970
rect 9220 1930 9580 1970
rect 9620 1930 9980 1970
rect 10020 1930 10380 1970
rect 10420 1930 10780 1970
rect 10820 1930 11180 1970
rect 11220 1930 11580 1970
rect 11620 1930 11980 1970
rect 12020 1930 12380 1970
rect 12420 1930 12780 1970
rect 12820 1930 13180 1970
rect 13220 1930 13580 1970
rect 13620 1930 13980 1970
rect 14020 1930 14380 1970
rect 14420 1930 14780 1970
rect 14820 1930 15180 1970
rect 15220 1930 15580 1970
rect 15620 1930 16000 1970
rect 0 1400 16000 1930
rect 1000 565 15000 600
rect 1000 525 1022 565
rect 1062 525 1120 565
rect 1160 525 1218 565
rect 1258 525 1316 565
rect 1356 525 1414 565
rect 1454 525 1512 565
rect 1552 525 1610 565
rect 1650 525 1708 565
rect 1748 525 1806 565
rect 1846 525 1904 565
rect 1944 525 2002 565
rect 2042 525 2100 565
rect 2140 525 2198 565
rect 2238 525 2296 565
rect 2336 525 2394 565
rect 2434 525 2492 565
rect 2532 525 2590 565
rect 2630 525 2688 565
rect 2728 525 2786 565
rect 2826 525 2884 565
rect 2924 525 2982 565
rect 3022 525 3080 565
rect 3120 525 3178 565
rect 3218 525 3276 565
rect 3316 525 3374 565
rect 3414 525 3472 565
rect 3512 525 3570 565
rect 3610 525 3668 565
rect 3708 525 3766 565
rect 3806 525 3864 565
rect 3904 525 3962 565
rect 4002 525 4060 565
rect 4100 525 4158 565
rect 4198 525 4256 565
rect 4296 525 4354 565
rect 4394 525 4452 565
rect 4492 525 4550 565
rect 4590 525 4648 565
rect 4688 525 4746 565
rect 4786 525 4844 565
rect 4884 525 4942 565
rect 4982 525 5040 565
rect 5080 525 5138 565
rect 5178 525 5236 565
rect 5276 525 5334 565
rect 5374 525 5432 565
rect 5472 525 5530 565
rect 5570 525 5628 565
rect 5668 525 5726 565
rect 5766 525 5824 565
rect 5864 525 5922 565
rect 5962 525 6020 565
rect 6060 525 6118 565
rect 6158 525 6216 565
rect 6256 525 6314 565
rect 6354 525 6412 565
rect 6452 525 6510 565
rect 6550 525 6608 565
rect 6648 525 6706 565
rect 6746 525 6804 565
rect 6844 525 6902 565
rect 6942 525 7000 565
rect 7040 525 7098 565
rect 7138 525 7196 565
rect 7236 525 7294 565
rect 7334 525 7392 565
rect 7432 525 7490 565
rect 7530 525 7588 565
rect 7628 525 7686 565
rect 7726 525 7784 565
rect 7824 525 7882 565
rect 7922 525 7980 565
rect 8020 525 8078 565
rect 8118 525 8176 565
rect 8216 525 8274 565
rect 8314 525 8372 565
rect 8412 525 8470 565
rect 8510 525 8568 565
rect 8608 525 8666 565
rect 8706 525 8764 565
rect 8804 525 8862 565
rect 8902 525 8960 565
rect 9000 525 9058 565
rect 9098 525 9156 565
rect 9196 525 9254 565
rect 9294 525 9352 565
rect 9392 525 9450 565
rect 9490 525 9548 565
rect 9588 525 9646 565
rect 9686 525 9744 565
rect 9784 525 9842 565
rect 9882 525 9940 565
rect 9980 525 10038 565
rect 10078 525 10136 565
rect 10176 525 10234 565
rect 10274 525 10332 565
rect 10372 525 10430 565
rect 10470 525 10528 565
rect 10568 525 10626 565
rect 10666 525 10724 565
rect 10764 525 10822 565
rect 10862 525 10920 565
rect 10960 525 11018 565
rect 11058 525 11116 565
rect 11156 525 11214 565
rect 11254 525 11312 565
rect 11352 525 11410 565
rect 11450 525 11508 565
rect 11548 525 11606 565
rect 11646 525 11704 565
rect 11744 525 11802 565
rect 11842 525 11900 565
rect 11940 525 11998 565
rect 12038 525 12096 565
rect 12136 525 12194 565
rect 12234 525 12292 565
rect 12332 525 12390 565
rect 12430 525 12488 565
rect 12528 525 12586 565
rect 12626 525 12684 565
rect 12724 525 12782 565
rect 12822 525 12880 565
rect 12920 525 12978 565
rect 13018 525 13076 565
rect 13116 525 13174 565
rect 13214 525 13272 565
rect 13312 525 13370 565
rect 13410 525 13468 565
rect 13508 525 13566 565
rect 13606 525 13664 565
rect 13704 525 13762 565
rect 13802 525 13860 565
rect 13900 525 13958 565
rect 13998 525 14056 565
rect 14096 525 14154 565
rect 14194 525 14252 565
rect 14292 525 14350 565
rect 14390 525 14448 565
rect 14488 525 14546 565
rect 14586 525 14644 565
rect 14684 525 14742 565
rect 14782 525 14840 565
rect 14880 525 14938 565
rect 14978 525 15000 565
rect 1000 520 15000 525
rect 1000 480 1180 520
rect 1220 480 1580 520
rect 1620 480 1980 520
rect 2020 480 2380 520
rect 2420 480 2780 520
rect 2820 480 3180 520
rect 3220 480 3580 520
rect 3620 480 3980 520
rect 4020 480 4380 520
rect 4420 480 4780 520
rect 4820 480 5180 520
rect 5220 480 5580 520
rect 5620 480 5980 520
rect 6020 480 6380 520
rect 6420 480 6780 520
rect 6820 480 7180 520
rect 7220 480 7580 520
rect 7620 480 7980 520
rect 8020 480 8380 520
rect 8420 480 8780 520
rect 8820 480 9180 520
rect 9220 480 9580 520
rect 9620 480 9980 520
rect 10020 480 10380 520
rect 10420 480 10780 520
rect 10820 480 11180 520
rect 11220 480 11580 520
rect 11620 480 11980 520
rect 12020 480 12380 520
rect 12420 480 12780 520
rect 12820 480 13180 520
rect 13220 480 13580 520
rect 13620 480 13980 520
rect 14020 480 14380 520
rect 14420 480 14780 520
rect 14820 480 15000 520
rect 1000 467 15000 480
rect 1000 427 1022 467
rect 1062 427 1120 467
rect 1160 427 1218 467
rect 1258 427 1316 467
rect 1356 427 1414 467
rect 1454 427 1512 467
rect 1552 427 1610 467
rect 1650 427 1708 467
rect 1748 427 1806 467
rect 1846 427 1904 467
rect 1944 427 2002 467
rect 2042 427 2100 467
rect 2140 427 2198 467
rect 2238 427 2296 467
rect 2336 427 2394 467
rect 2434 427 2492 467
rect 2532 427 2590 467
rect 2630 427 2688 467
rect 2728 427 2786 467
rect 2826 427 2884 467
rect 2924 427 2982 467
rect 3022 427 3080 467
rect 3120 427 3178 467
rect 3218 427 3276 467
rect 3316 427 3374 467
rect 3414 427 3472 467
rect 3512 427 3570 467
rect 3610 427 3668 467
rect 3708 427 3766 467
rect 3806 427 3864 467
rect 3904 427 3962 467
rect 4002 427 4060 467
rect 4100 427 4158 467
rect 4198 427 4256 467
rect 4296 427 4354 467
rect 4394 427 4452 467
rect 4492 427 4550 467
rect 4590 427 4648 467
rect 4688 427 4746 467
rect 4786 427 4844 467
rect 4884 427 4942 467
rect 4982 427 5040 467
rect 5080 427 5138 467
rect 5178 427 5236 467
rect 5276 427 5334 467
rect 5374 427 5432 467
rect 5472 427 5530 467
rect 5570 427 5628 467
rect 5668 427 5726 467
rect 5766 427 5824 467
rect 5864 427 5922 467
rect 5962 427 6020 467
rect 6060 427 6118 467
rect 6158 427 6216 467
rect 6256 427 6314 467
rect 6354 427 6412 467
rect 6452 427 6510 467
rect 6550 427 6608 467
rect 6648 427 6706 467
rect 6746 427 6804 467
rect 6844 427 6902 467
rect 6942 427 7000 467
rect 7040 427 7098 467
rect 7138 427 7196 467
rect 7236 427 7294 467
rect 7334 427 7392 467
rect 7432 427 7490 467
rect 7530 427 7588 467
rect 7628 427 7686 467
rect 7726 427 7784 467
rect 7824 427 7882 467
rect 7922 427 7980 467
rect 8020 427 8078 467
rect 8118 427 8176 467
rect 8216 427 8274 467
rect 8314 427 8372 467
rect 8412 427 8470 467
rect 8510 427 8568 467
rect 8608 427 8666 467
rect 8706 427 8764 467
rect 8804 427 8862 467
rect 8902 427 8960 467
rect 9000 427 9058 467
rect 9098 427 9156 467
rect 9196 427 9254 467
rect 9294 427 9352 467
rect 9392 427 9450 467
rect 9490 427 9548 467
rect 9588 427 9646 467
rect 9686 427 9744 467
rect 9784 427 9842 467
rect 9882 427 9940 467
rect 9980 427 10038 467
rect 10078 427 10136 467
rect 10176 427 10234 467
rect 10274 427 10332 467
rect 10372 427 10430 467
rect 10470 427 10528 467
rect 10568 427 10626 467
rect 10666 427 10724 467
rect 10764 427 10822 467
rect 10862 427 10920 467
rect 10960 427 11018 467
rect 11058 427 11116 467
rect 11156 427 11214 467
rect 11254 427 11312 467
rect 11352 427 11410 467
rect 11450 427 11508 467
rect 11548 427 11606 467
rect 11646 427 11704 467
rect 11744 427 11802 467
rect 11842 427 11900 467
rect 11940 427 11998 467
rect 12038 427 12096 467
rect 12136 427 12194 467
rect 12234 427 12292 467
rect 12332 427 12390 467
rect 12430 427 12488 467
rect 12528 427 12586 467
rect 12626 427 12684 467
rect 12724 427 12782 467
rect 12822 427 12880 467
rect 12920 427 12978 467
rect 13018 427 13076 467
rect 13116 427 13174 467
rect 13214 427 13272 467
rect 13312 427 13370 467
rect 13410 427 13468 467
rect 13508 427 13566 467
rect 13606 427 13664 467
rect 13704 427 13762 467
rect 13802 427 13860 467
rect 13900 427 13958 467
rect 13998 427 14056 467
rect 14096 427 14154 467
rect 14194 427 14252 467
rect 14292 427 14350 467
rect 14390 427 14448 467
rect 14488 427 14546 467
rect 14586 427 14644 467
rect 14684 427 14742 467
rect 14782 427 14840 467
rect 14880 427 14938 467
rect 14978 427 15000 467
rect 1000 369 15000 427
rect 1000 329 1022 369
rect 1062 329 1120 369
rect 1160 329 1218 369
rect 1258 329 1316 369
rect 1356 329 1414 369
rect 1454 329 1512 369
rect 1552 329 1610 369
rect 1650 329 1708 369
rect 1748 329 1806 369
rect 1846 329 1904 369
rect 1944 329 2002 369
rect 2042 329 2100 369
rect 2140 329 2198 369
rect 2238 329 2296 369
rect 2336 329 2394 369
rect 2434 329 2492 369
rect 2532 329 2590 369
rect 2630 329 2688 369
rect 2728 329 2786 369
rect 2826 329 2884 369
rect 2924 329 2982 369
rect 3022 329 3080 369
rect 3120 329 3178 369
rect 3218 329 3276 369
rect 3316 329 3374 369
rect 3414 329 3472 369
rect 3512 329 3570 369
rect 3610 329 3668 369
rect 3708 329 3766 369
rect 3806 329 3864 369
rect 3904 329 3962 369
rect 4002 329 4060 369
rect 4100 329 4158 369
rect 4198 329 4256 369
rect 4296 329 4354 369
rect 4394 329 4452 369
rect 4492 329 4550 369
rect 4590 329 4648 369
rect 4688 329 4746 369
rect 4786 329 4844 369
rect 4884 329 4942 369
rect 4982 329 5040 369
rect 5080 329 5138 369
rect 5178 329 5236 369
rect 5276 329 5334 369
rect 5374 329 5432 369
rect 5472 329 5530 369
rect 5570 329 5628 369
rect 5668 329 5726 369
rect 5766 329 5824 369
rect 5864 329 5922 369
rect 5962 329 6020 369
rect 6060 329 6118 369
rect 6158 329 6216 369
rect 6256 329 6314 369
rect 6354 329 6412 369
rect 6452 329 6510 369
rect 6550 329 6608 369
rect 6648 329 6706 369
rect 6746 329 6804 369
rect 6844 329 6902 369
rect 6942 329 7000 369
rect 7040 329 7098 369
rect 7138 329 7196 369
rect 7236 329 7294 369
rect 7334 329 7392 369
rect 7432 329 7490 369
rect 7530 329 7588 369
rect 7628 329 7686 369
rect 7726 329 7784 369
rect 7824 329 7882 369
rect 7922 329 7980 369
rect 8020 329 8078 369
rect 8118 329 8176 369
rect 8216 329 8274 369
rect 8314 329 8372 369
rect 8412 329 8470 369
rect 8510 329 8568 369
rect 8608 329 8666 369
rect 8706 329 8764 369
rect 8804 329 8862 369
rect 8902 329 8960 369
rect 9000 329 9058 369
rect 9098 329 9156 369
rect 9196 329 9254 369
rect 9294 329 9352 369
rect 9392 329 9450 369
rect 9490 329 9548 369
rect 9588 329 9646 369
rect 9686 329 9744 369
rect 9784 329 9842 369
rect 9882 329 9940 369
rect 9980 329 10038 369
rect 10078 329 10136 369
rect 10176 329 10234 369
rect 10274 329 10332 369
rect 10372 329 10430 369
rect 10470 329 10528 369
rect 10568 329 10626 369
rect 10666 329 10724 369
rect 10764 329 10822 369
rect 10862 329 10920 369
rect 10960 329 11018 369
rect 11058 329 11116 369
rect 11156 329 11214 369
rect 11254 329 11312 369
rect 11352 329 11410 369
rect 11450 329 11508 369
rect 11548 329 11606 369
rect 11646 329 11704 369
rect 11744 329 11802 369
rect 11842 329 11900 369
rect 11940 329 11998 369
rect 12038 329 12096 369
rect 12136 329 12194 369
rect 12234 329 12292 369
rect 12332 329 12390 369
rect 12430 329 12488 369
rect 12528 329 12586 369
rect 12626 329 12684 369
rect 12724 329 12782 369
rect 12822 329 12880 369
rect 12920 329 12978 369
rect 13018 329 13076 369
rect 13116 329 13174 369
rect 13214 329 13272 369
rect 13312 329 13370 369
rect 13410 329 13468 369
rect 13508 329 13566 369
rect 13606 329 13664 369
rect 13704 329 13762 369
rect 13802 329 13860 369
rect 13900 329 13958 369
rect 13998 329 14056 369
rect 14096 329 14154 369
rect 14194 329 14252 369
rect 14292 329 14350 369
rect 14390 329 14448 369
rect 14488 329 14546 369
rect 14586 329 14644 369
rect 14684 329 14742 369
rect 14782 329 14840 369
rect 14880 329 14938 369
rect 14978 329 15000 369
rect 1000 271 15000 329
rect 1000 231 1022 271
rect 1062 231 1120 271
rect 1160 231 1218 271
rect 1258 231 1316 271
rect 1356 231 1414 271
rect 1454 231 1512 271
rect 1552 231 1610 271
rect 1650 231 1708 271
rect 1748 231 1806 271
rect 1846 231 1904 271
rect 1944 231 2002 271
rect 2042 231 2100 271
rect 2140 231 2198 271
rect 2238 231 2296 271
rect 2336 231 2394 271
rect 2434 231 2492 271
rect 2532 231 2590 271
rect 2630 231 2688 271
rect 2728 231 2786 271
rect 2826 231 2884 271
rect 2924 231 2982 271
rect 3022 231 3080 271
rect 3120 231 3178 271
rect 3218 231 3276 271
rect 3316 231 3374 271
rect 3414 231 3472 271
rect 3512 231 3570 271
rect 3610 231 3668 271
rect 3708 231 3766 271
rect 3806 231 3864 271
rect 3904 231 3962 271
rect 4002 231 4060 271
rect 4100 231 4158 271
rect 4198 231 4256 271
rect 4296 231 4354 271
rect 4394 231 4452 271
rect 4492 231 4550 271
rect 4590 231 4648 271
rect 4688 231 4746 271
rect 4786 231 4844 271
rect 4884 231 4942 271
rect 4982 231 5040 271
rect 5080 231 5138 271
rect 5178 231 5236 271
rect 5276 231 5334 271
rect 5374 231 5432 271
rect 5472 231 5530 271
rect 5570 231 5628 271
rect 5668 231 5726 271
rect 5766 231 5824 271
rect 5864 231 5922 271
rect 5962 231 6020 271
rect 6060 231 6118 271
rect 6158 231 6216 271
rect 6256 231 6314 271
rect 6354 231 6412 271
rect 6452 231 6510 271
rect 6550 231 6608 271
rect 6648 231 6706 271
rect 6746 231 6804 271
rect 6844 231 6902 271
rect 6942 231 7000 271
rect 7040 231 7098 271
rect 7138 231 7196 271
rect 7236 231 7294 271
rect 7334 231 7392 271
rect 7432 231 7490 271
rect 7530 231 7588 271
rect 7628 231 7686 271
rect 7726 231 7784 271
rect 7824 231 7882 271
rect 7922 231 7980 271
rect 8020 231 8078 271
rect 8118 231 8176 271
rect 8216 231 8274 271
rect 8314 231 8372 271
rect 8412 231 8470 271
rect 8510 231 8568 271
rect 8608 231 8666 271
rect 8706 231 8764 271
rect 8804 231 8862 271
rect 8902 231 8960 271
rect 9000 231 9058 271
rect 9098 231 9156 271
rect 9196 231 9254 271
rect 9294 231 9352 271
rect 9392 231 9450 271
rect 9490 231 9548 271
rect 9588 231 9646 271
rect 9686 231 9744 271
rect 9784 231 9842 271
rect 9882 231 9940 271
rect 9980 231 10038 271
rect 10078 231 10136 271
rect 10176 231 10234 271
rect 10274 231 10332 271
rect 10372 231 10430 271
rect 10470 231 10528 271
rect 10568 231 10626 271
rect 10666 231 10724 271
rect 10764 231 10822 271
rect 10862 231 10920 271
rect 10960 231 11018 271
rect 11058 231 11116 271
rect 11156 231 11214 271
rect 11254 231 11312 271
rect 11352 231 11410 271
rect 11450 231 11508 271
rect 11548 231 11606 271
rect 11646 231 11704 271
rect 11744 231 11802 271
rect 11842 231 11900 271
rect 11940 231 11998 271
rect 12038 231 12096 271
rect 12136 231 12194 271
rect 12234 231 12292 271
rect 12332 231 12390 271
rect 12430 231 12488 271
rect 12528 231 12586 271
rect 12626 231 12684 271
rect 12724 231 12782 271
rect 12822 231 12880 271
rect 12920 231 12978 271
rect 13018 231 13076 271
rect 13116 231 13174 271
rect 13214 231 13272 271
rect 13312 231 13370 271
rect 13410 231 13468 271
rect 13508 231 13566 271
rect 13606 231 13664 271
rect 13704 231 13762 271
rect 13802 231 13860 271
rect 13900 231 13958 271
rect 13998 231 14056 271
rect 14096 231 14154 271
rect 14194 231 14252 271
rect 14292 231 14350 271
rect 14390 231 14448 271
rect 14488 231 14546 271
rect 14586 231 14644 271
rect 14684 231 14742 271
rect 14782 231 14840 271
rect 14880 231 14938 271
rect 14978 231 15000 271
rect 1000 173 15000 231
rect 1000 133 1022 173
rect 1062 133 1120 173
rect 1160 133 1218 173
rect 1258 133 1316 173
rect 1356 133 1414 173
rect 1454 133 1512 173
rect 1552 133 1610 173
rect 1650 133 1708 173
rect 1748 133 1806 173
rect 1846 133 1904 173
rect 1944 133 2002 173
rect 2042 133 2100 173
rect 2140 133 2198 173
rect 2238 133 2296 173
rect 2336 133 2394 173
rect 2434 133 2492 173
rect 2532 133 2590 173
rect 2630 133 2688 173
rect 2728 133 2786 173
rect 2826 133 2884 173
rect 2924 133 2982 173
rect 3022 133 3080 173
rect 3120 133 3178 173
rect 3218 133 3276 173
rect 3316 133 3374 173
rect 3414 133 3472 173
rect 3512 133 3570 173
rect 3610 133 3668 173
rect 3708 133 3766 173
rect 3806 133 3864 173
rect 3904 133 3962 173
rect 4002 133 4060 173
rect 4100 133 4158 173
rect 4198 133 4256 173
rect 4296 133 4354 173
rect 4394 133 4452 173
rect 4492 133 4550 173
rect 4590 133 4648 173
rect 4688 133 4746 173
rect 4786 133 4844 173
rect 4884 133 4942 173
rect 4982 133 5040 173
rect 5080 133 5138 173
rect 5178 133 5236 173
rect 5276 133 5334 173
rect 5374 133 5432 173
rect 5472 133 5530 173
rect 5570 133 5628 173
rect 5668 133 5726 173
rect 5766 133 5824 173
rect 5864 133 5922 173
rect 5962 133 6020 173
rect 6060 133 6118 173
rect 6158 133 6216 173
rect 6256 133 6314 173
rect 6354 133 6412 173
rect 6452 133 6510 173
rect 6550 133 6608 173
rect 6648 133 6706 173
rect 6746 133 6804 173
rect 6844 133 6902 173
rect 6942 133 7000 173
rect 7040 133 7098 173
rect 7138 133 7196 173
rect 7236 133 7294 173
rect 7334 133 7392 173
rect 7432 133 7490 173
rect 7530 133 7588 173
rect 7628 133 7686 173
rect 7726 133 7784 173
rect 7824 133 7882 173
rect 7922 133 7980 173
rect 8020 133 8078 173
rect 8118 133 8176 173
rect 8216 133 8274 173
rect 8314 133 8372 173
rect 8412 133 8470 173
rect 8510 133 8568 173
rect 8608 133 8666 173
rect 8706 133 8764 173
rect 8804 133 8862 173
rect 8902 133 8960 173
rect 9000 133 9058 173
rect 9098 133 9156 173
rect 9196 133 9254 173
rect 9294 133 9352 173
rect 9392 133 9450 173
rect 9490 133 9548 173
rect 9588 133 9646 173
rect 9686 133 9744 173
rect 9784 133 9842 173
rect 9882 133 9940 173
rect 9980 133 10038 173
rect 10078 133 10136 173
rect 10176 133 10234 173
rect 10274 133 10332 173
rect 10372 133 10430 173
rect 10470 133 10528 173
rect 10568 133 10626 173
rect 10666 133 10724 173
rect 10764 133 10822 173
rect 10862 133 10920 173
rect 10960 133 11018 173
rect 11058 133 11116 173
rect 11156 133 11214 173
rect 11254 133 11312 173
rect 11352 133 11410 173
rect 11450 133 11508 173
rect 11548 133 11606 173
rect 11646 133 11704 173
rect 11744 133 11802 173
rect 11842 133 11900 173
rect 11940 133 11998 173
rect 12038 133 12096 173
rect 12136 133 12194 173
rect 12234 133 12292 173
rect 12332 133 12390 173
rect 12430 133 12488 173
rect 12528 133 12586 173
rect 12626 133 12684 173
rect 12724 133 12782 173
rect 12822 133 12880 173
rect 12920 133 12978 173
rect 13018 133 13076 173
rect 13116 133 13174 173
rect 13214 133 13272 173
rect 13312 133 13370 173
rect 13410 133 13468 173
rect 13508 133 13566 173
rect 13606 133 13664 173
rect 13704 133 13762 173
rect 13802 133 13860 173
rect 13900 133 13958 173
rect 13998 133 14056 173
rect 14096 133 14154 173
rect 14194 133 14252 173
rect 14292 133 14350 173
rect 14390 133 14448 173
rect 14488 133 14546 173
rect 14586 133 14644 173
rect 14684 133 14742 173
rect 14782 133 14840 173
rect 14880 133 14938 173
rect 14978 133 15000 173
rect 1000 120 15000 133
rect 1000 80 1180 120
rect 1220 80 1580 120
rect 1620 80 1980 120
rect 2020 80 2380 120
rect 2420 80 2780 120
rect 2820 80 3180 120
rect 3220 80 3580 120
rect 3620 80 3980 120
rect 4020 80 4380 120
rect 4420 80 4780 120
rect 4820 80 5180 120
rect 5220 80 5580 120
rect 5620 80 5980 120
rect 6020 80 6380 120
rect 6420 80 6780 120
rect 6820 80 7180 120
rect 7220 80 7580 120
rect 7620 80 7980 120
rect 8020 80 8380 120
rect 8420 80 8780 120
rect 8820 80 9180 120
rect 9220 80 9580 120
rect 9620 80 9980 120
rect 10020 80 10380 120
rect 10420 80 10780 120
rect 10820 80 11180 120
rect 11220 80 11580 120
rect 11620 80 11980 120
rect 12020 80 12380 120
rect 12420 80 12780 120
rect 12820 80 13180 120
rect 13220 80 13580 120
rect 13620 80 13980 120
rect 14020 80 14380 120
rect 14420 80 14780 120
rect 14820 80 15000 120
rect 1000 75 15000 80
rect 1000 35 1022 75
rect 1062 35 1120 75
rect 1160 35 1218 75
rect 1258 35 1316 75
rect 1356 35 1414 75
rect 1454 35 1512 75
rect 1552 35 1610 75
rect 1650 35 1708 75
rect 1748 35 1806 75
rect 1846 35 1904 75
rect 1944 35 2002 75
rect 2042 35 2100 75
rect 2140 35 2198 75
rect 2238 35 2296 75
rect 2336 35 2394 75
rect 2434 35 2492 75
rect 2532 35 2590 75
rect 2630 35 2688 75
rect 2728 35 2786 75
rect 2826 35 2884 75
rect 2924 35 2982 75
rect 3022 35 3080 75
rect 3120 35 3178 75
rect 3218 35 3276 75
rect 3316 35 3374 75
rect 3414 35 3472 75
rect 3512 35 3570 75
rect 3610 35 3668 75
rect 3708 35 3766 75
rect 3806 35 3864 75
rect 3904 35 3962 75
rect 4002 35 4060 75
rect 4100 35 4158 75
rect 4198 35 4256 75
rect 4296 35 4354 75
rect 4394 35 4452 75
rect 4492 35 4550 75
rect 4590 35 4648 75
rect 4688 35 4746 75
rect 4786 35 4844 75
rect 4884 35 4942 75
rect 4982 35 5040 75
rect 5080 35 5138 75
rect 5178 35 5236 75
rect 5276 35 5334 75
rect 5374 35 5432 75
rect 5472 35 5530 75
rect 5570 35 5628 75
rect 5668 35 5726 75
rect 5766 35 5824 75
rect 5864 35 5922 75
rect 5962 35 6020 75
rect 6060 35 6118 75
rect 6158 35 6216 75
rect 6256 35 6314 75
rect 6354 35 6412 75
rect 6452 35 6510 75
rect 6550 35 6608 75
rect 6648 35 6706 75
rect 6746 35 6804 75
rect 6844 35 6902 75
rect 6942 35 7000 75
rect 7040 35 7098 75
rect 7138 35 7196 75
rect 7236 35 7294 75
rect 7334 35 7392 75
rect 7432 35 7490 75
rect 7530 35 7588 75
rect 7628 35 7686 75
rect 7726 35 7784 75
rect 7824 35 7882 75
rect 7922 35 7980 75
rect 8020 35 8078 75
rect 8118 35 8176 75
rect 8216 35 8274 75
rect 8314 35 8372 75
rect 8412 35 8470 75
rect 8510 35 8568 75
rect 8608 35 8666 75
rect 8706 35 8764 75
rect 8804 35 8862 75
rect 8902 35 8960 75
rect 9000 35 9058 75
rect 9098 35 9156 75
rect 9196 35 9254 75
rect 9294 35 9352 75
rect 9392 35 9450 75
rect 9490 35 9548 75
rect 9588 35 9646 75
rect 9686 35 9744 75
rect 9784 35 9842 75
rect 9882 35 9940 75
rect 9980 35 10038 75
rect 10078 35 10136 75
rect 10176 35 10234 75
rect 10274 35 10332 75
rect 10372 35 10430 75
rect 10470 35 10528 75
rect 10568 35 10626 75
rect 10666 35 10724 75
rect 10764 35 10822 75
rect 10862 35 10920 75
rect 10960 35 11018 75
rect 11058 35 11116 75
rect 11156 35 11214 75
rect 11254 35 11312 75
rect 11352 35 11410 75
rect 11450 35 11508 75
rect 11548 35 11606 75
rect 11646 35 11704 75
rect 11744 35 11802 75
rect 11842 35 11900 75
rect 11940 35 11998 75
rect 12038 35 12096 75
rect 12136 35 12194 75
rect 12234 35 12292 75
rect 12332 35 12390 75
rect 12430 35 12488 75
rect 12528 35 12586 75
rect 12626 35 12684 75
rect 12724 35 12782 75
rect 12822 35 12880 75
rect 12920 35 12978 75
rect 13018 35 13076 75
rect 13116 35 13174 75
rect 13214 35 13272 75
rect 13312 35 13370 75
rect 13410 35 13468 75
rect 13508 35 13566 75
rect 13606 35 13664 75
rect 13704 35 13762 75
rect 13802 35 13860 75
rect 13900 35 13958 75
rect 13998 35 14056 75
rect 14096 35 14154 75
rect 14194 35 14252 75
rect 14292 35 14350 75
rect 14390 35 14448 75
rect 14488 35 14546 75
rect 14586 35 14644 75
rect 14684 35 14742 75
rect 14782 35 14840 75
rect 14880 35 14938 75
rect 14978 35 15000 75
rect 1000 0 15000 35
<< via3 >>
rect 249 32000 7751 32040
rect 8249 31560 15751 31600
rect 380 26380 420 26420
rect 780 26380 820 26420
rect 1180 26380 1220 26420
rect 1580 26380 1620 26420
rect 1980 26380 2020 26420
rect 2380 26380 2420 26420
rect 2780 26380 2820 26420
rect 3180 26380 3220 26420
rect 3580 26380 3620 26420
rect 3980 26380 4020 26420
rect 4380 26380 4420 26420
rect 4780 26380 4820 26420
rect 5180 26380 5220 26420
rect 5580 26380 5620 26420
rect 5980 26380 6020 26420
rect 6380 26380 6420 26420
rect 6780 26380 6820 26420
rect 7180 26380 7220 26420
rect 7580 26380 7620 26420
rect 7980 26380 8020 26420
rect 8380 26380 8420 26420
rect 8780 26380 8820 26420
rect 9180 26380 9220 26420
rect 9580 26380 9620 26420
rect 9980 26380 10020 26420
rect 10380 26380 10420 26420
rect 10780 26380 10820 26420
rect 11180 26380 11220 26420
rect 11580 26380 11620 26420
rect 11980 26380 12020 26420
rect 12380 26380 12420 26420
rect 12780 26380 12820 26420
rect 13180 26380 13220 26420
rect 13580 26380 13620 26420
rect 13980 26380 14020 26420
rect 14380 26380 14420 26420
rect 14780 26380 14820 26420
rect 15180 26380 15220 26420
rect 15580 26380 15620 26420
rect 380 25980 420 26020
rect 780 25980 820 26020
rect 1180 25980 1220 26020
rect 1580 25980 1620 26020
rect 1980 25980 2020 26020
rect 2380 25980 2420 26020
rect 2780 25980 2820 26020
rect 3180 25980 3220 26020
rect 3580 25980 3620 26020
rect 3980 25980 4020 26020
rect 4380 25980 4420 26020
rect 4780 25980 4820 26020
rect 5180 25980 5220 26020
rect 5580 25980 5620 26020
rect 5980 25980 6020 26020
rect 6380 25980 6420 26020
rect 6780 25980 6820 26020
rect 7180 25980 7220 26020
rect 7580 25980 7620 26020
rect 7980 25980 8020 26020
rect 8380 25980 8420 26020
rect 8780 25980 8820 26020
rect 9180 25980 9220 26020
rect 9580 25980 9620 26020
rect 9980 25980 10020 26020
rect 10380 25980 10420 26020
rect 10780 25980 10820 26020
rect 11180 25980 11220 26020
rect 11580 25980 11620 26020
rect 11980 25980 12020 26020
rect 12380 25980 12420 26020
rect 12780 25980 12820 26020
rect 13180 25980 13220 26020
rect 13580 25980 13620 26020
rect 13980 25980 14020 26020
rect 14380 25980 14420 26020
rect 14780 25980 14820 26020
rect 15180 25980 15220 26020
rect 15580 25980 15620 26020
rect 380 25580 420 25620
rect 780 25580 820 25620
rect 1180 25580 1220 25620
rect 1580 25580 1620 25620
rect 1980 25580 2020 25620
rect 2380 25580 2420 25620
rect 2780 25580 2820 25620
rect 3180 25580 3220 25620
rect 3580 25580 3620 25620
rect 3980 25580 4020 25620
rect 4380 25580 4420 25620
rect 4780 25580 4820 25620
rect 5180 25580 5220 25620
rect 5580 25580 5620 25620
rect 5980 25580 6020 25620
rect 6380 25580 6420 25620
rect 6780 25580 6820 25620
rect 7180 25580 7220 25620
rect 7580 25580 7620 25620
rect 7980 25580 8020 25620
rect 8380 25580 8420 25620
rect 8780 25580 8820 25620
rect 9180 25580 9220 25620
rect 9580 25580 9620 25620
rect 9980 25580 10020 25620
rect 10380 25580 10420 25620
rect 10780 25580 10820 25620
rect 11180 25580 11220 25620
rect 11580 25580 11620 25620
rect 11980 25580 12020 25620
rect 12380 25580 12420 25620
rect 12780 25580 12820 25620
rect 13180 25580 13220 25620
rect 13580 25580 13620 25620
rect 13980 25580 14020 25620
rect 14380 25580 14420 25620
rect 14780 25580 14820 25620
rect 15180 25580 15220 25620
rect 15580 25580 15620 25620
rect 380 23230 420 23270
rect 780 23230 820 23270
rect 1180 23230 1220 23270
rect 1580 23230 1620 23270
rect 1980 23230 2020 23270
rect 2380 23230 2420 23270
rect 2780 23230 2820 23270
rect 3180 23230 3220 23270
rect 3580 23230 3620 23270
rect 3980 23230 4020 23270
rect 4380 23230 4420 23270
rect 4780 23230 4820 23270
rect 5180 23230 5220 23270
rect 5580 23230 5620 23270
rect 5980 23230 6020 23270
rect 6380 23230 6420 23270
rect 6780 23230 6820 23270
rect 7180 23230 7220 23270
rect 7580 23230 7620 23270
rect 7980 23230 8020 23270
rect 8380 23230 8420 23270
rect 8780 23230 8820 23270
rect 9180 23230 9220 23270
rect 9580 23230 9620 23270
rect 9980 23230 10020 23270
rect 10380 23230 10420 23270
rect 10780 23230 10820 23270
rect 11180 23230 11220 23270
rect 11580 23230 11620 23270
rect 11980 23230 12020 23270
rect 12380 23230 12420 23270
rect 12780 23230 12820 23270
rect 13180 23230 13220 23270
rect 13580 23230 13620 23270
rect 13980 23230 14020 23270
rect 14380 23230 14420 23270
rect 14780 23230 14820 23270
rect 15180 23230 15220 23270
rect 15580 23230 15620 23270
rect 380 22830 420 22870
rect 780 22830 820 22870
rect 1180 22830 1220 22870
rect 1580 22830 1620 22870
rect 1980 22830 2020 22870
rect 2380 22830 2420 22870
rect 2780 22830 2820 22870
rect 3180 22830 3220 22870
rect 3580 22830 3620 22870
rect 3980 22830 4020 22870
rect 4380 22830 4420 22870
rect 4780 22830 4820 22870
rect 5180 22830 5220 22870
rect 5580 22830 5620 22870
rect 5980 22830 6020 22870
rect 6380 22830 6420 22870
rect 6780 22830 6820 22870
rect 7180 22830 7220 22870
rect 7580 22830 7620 22870
rect 7980 22830 8020 22870
rect 8380 22830 8420 22870
rect 8780 22830 8820 22870
rect 9180 22830 9220 22870
rect 9580 22830 9620 22870
rect 9980 22830 10020 22870
rect 10380 22830 10420 22870
rect 10780 22830 10820 22870
rect 11180 22830 11220 22870
rect 11580 22830 11620 22870
rect 11980 22830 12020 22870
rect 12380 22830 12420 22870
rect 12780 22830 12820 22870
rect 13180 22830 13220 22870
rect 13580 22830 13620 22870
rect 13980 22830 14020 22870
rect 14380 22830 14420 22870
rect 14780 22830 14820 22870
rect 15180 22830 15220 22870
rect 15580 22830 15620 22870
rect 380 22430 420 22470
rect 780 22430 820 22470
rect 1180 22430 1220 22470
rect 1580 22430 1620 22470
rect 1980 22430 2020 22470
rect 2380 22430 2420 22470
rect 2780 22430 2820 22470
rect 3180 22430 3220 22470
rect 3580 22430 3620 22470
rect 3980 22430 4020 22470
rect 4380 22430 4420 22470
rect 4780 22430 4820 22470
rect 5180 22430 5220 22470
rect 5580 22430 5620 22470
rect 5980 22430 6020 22470
rect 6380 22430 6420 22470
rect 6780 22430 6820 22470
rect 7180 22430 7220 22470
rect 7580 22430 7620 22470
rect 7980 22430 8020 22470
rect 8380 22430 8420 22470
rect 8780 22430 8820 22470
rect 9180 22430 9220 22470
rect 9580 22430 9620 22470
rect 9980 22430 10020 22470
rect 10380 22430 10420 22470
rect 10780 22430 10820 22470
rect 11180 22430 11220 22470
rect 11580 22430 11620 22470
rect 11980 22430 12020 22470
rect 12380 22430 12420 22470
rect 12780 22430 12820 22470
rect 13180 22430 13220 22470
rect 13580 22430 13620 22470
rect 13980 22430 14020 22470
rect 14380 22430 14420 22470
rect 14780 22430 14820 22470
rect 15180 22430 15220 22470
rect 15580 22430 15620 22470
rect 380 22030 420 22070
rect 780 22030 820 22070
rect 1180 22030 1220 22070
rect 1580 22030 1620 22070
rect 1980 22030 2020 22070
rect 2380 22030 2420 22070
rect 2780 22030 2820 22070
rect 3180 22030 3220 22070
rect 3580 22030 3620 22070
rect 3980 22030 4020 22070
rect 4380 22030 4420 22070
rect 4780 22030 4820 22070
rect 5180 22030 5220 22070
rect 5580 22030 5620 22070
rect 5980 22030 6020 22070
rect 6380 22030 6420 22070
rect 6780 22030 6820 22070
rect 7180 22030 7220 22070
rect 7580 22030 7620 22070
rect 7980 22030 8020 22070
rect 8380 22030 8420 22070
rect 8780 22030 8820 22070
rect 9180 22030 9220 22070
rect 9580 22030 9620 22070
rect 9980 22030 10020 22070
rect 10380 22030 10420 22070
rect 10780 22030 10820 22070
rect 11180 22030 11220 22070
rect 11580 22030 11620 22070
rect 11980 22030 12020 22070
rect 12380 22030 12420 22070
rect 12780 22030 12820 22070
rect 13180 22030 13220 22070
rect 13580 22030 13620 22070
rect 13980 22030 14020 22070
rect 14380 22030 14420 22070
rect 14780 22030 14820 22070
rect 15180 22030 15220 22070
rect 15580 22030 15620 22070
rect 380 21630 420 21670
rect 780 21630 820 21670
rect 1180 21630 1220 21670
rect 1580 21630 1620 21670
rect 1980 21630 2020 21670
rect 2380 21630 2420 21670
rect 2780 21630 2820 21670
rect 3180 21630 3220 21670
rect 3580 21630 3620 21670
rect 3980 21630 4020 21670
rect 4380 21630 4420 21670
rect 4780 21630 4820 21670
rect 5180 21630 5220 21670
rect 5580 21630 5620 21670
rect 5980 21630 6020 21670
rect 6380 21630 6420 21670
rect 6780 21630 6820 21670
rect 7180 21630 7220 21670
rect 7580 21630 7620 21670
rect 7980 21630 8020 21670
rect 8380 21630 8420 21670
rect 8780 21630 8820 21670
rect 9180 21630 9220 21670
rect 9580 21630 9620 21670
rect 9980 21630 10020 21670
rect 10380 21630 10420 21670
rect 10780 21630 10820 21670
rect 11180 21630 11220 21670
rect 11580 21630 11620 21670
rect 11980 21630 12020 21670
rect 12380 21630 12420 21670
rect 12780 21630 12820 21670
rect 13180 21630 13220 21670
rect 13580 21630 13620 21670
rect 13980 21630 14020 21670
rect 14380 21630 14420 21670
rect 14780 21630 14820 21670
rect 15180 21630 15220 21670
rect 15580 21630 15620 21670
rect 380 21230 420 21270
rect 780 21230 820 21270
rect 1180 21230 1220 21270
rect 1580 21230 1620 21270
rect 1980 21230 2020 21270
rect 2380 21230 2420 21270
rect 2780 21230 2820 21270
rect 3180 21230 3220 21270
rect 3580 21230 3620 21270
rect 3980 21230 4020 21270
rect 4380 21230 4420 21270
rect 4780 21230 4820 21270
rect 5180 21230 5220 21270
rect 5580 21230 5620 21270
rect 5980 21230 6020 21270
rect 6380 21230 6420 21270
rect 6780 21230 6820 21270
rect 7180 21230 7220 21270
rect 7580 21230 7620 21270
rect 7980 21230 8020 21270
rect 8380 21230 8420 21270
rect 8780 21230 8820 21270
rect 9180 21230 9220 21270
rect 9580 21230 9620 21270
rect 9980 21230 10020 21270
rect 10380 21230 10420 21270
rect 10780 21230 10820 21270
rect 11180 21230 11220 21270
rect 11580 21230 11620 21270
rect 11980 21230 12020 21270
rect 12380 21230 12420 21270
rect 12780 21230 12820 21270
rect 13180 21230 13220 21270
rect 13580 21230 13620 21270
rect 13980 21230 14020 21270
rect 14380 21230 14420 21270
rect 14780 21230 14820 21270
rect 15180 21230 15220 21270
rect 15580 21230 15620 21270
rect 380 20830 420 20870
rect 780 20830 820 20870
rect 1180 20830 1220 20870
rect 1580 20830 1620 20870
rect 1980 20830 2020 20870
rect 2380 20830 2420 20870
rect 2780 20830 2820 20870
rect 3180 20830 3220 20870
rect 3580 20830 3620 20870
rect 3980 20830 4020 20870
rect 4380 20830 4420 20870
rect 4780 20830 4820 20870
rect 5180 20830 5220 20870
rect 5580 20830 5620 20870
rect 5980 20830 6020 20870
rect 6380 20830 6420 20870
rect 6780 20830 6820 20870
rect 7180 20830 7220 20870
rect 7580 20830 7620 20870
rect 7980 20830 8020 20870
rect 8380 20830 8420 20870
rect 8780 20830 8820 20870
rect 9180 20830 9220 20870
rect 9580 20830 9620 20870
rect 9980 20830 10020 20870
rect 10380 20830 10420 20870
rect 10780 20830 10820 20870
rect 11180 20830 11220 20870
rect 11580 20830 11620 20870
rect 11980 20830 12020 20870
rect 12380 20830 12420 20870
rect 12780 20830 12820 20870
rect 13180 20830 13220 20870
rect 13580 20830 13620 20870
rect 13980 20830 14020 20870
rect 14380 20830 14420 20870
rect 14780 20830 14820 20870
rect 15180 20830 15220 20870
rect 15580 20830 15620 20870
rect 380 20430 420 20470
rect 780 20430 820 20470
rect 1180 20430 1220 20470
rect 1580 20430 1620 20470
rect 1980 20430 2020 20470
rect 2380 20430 2420 20470
rect 2780 20430 2820 20470
rect 3180 20430 3220 20470
rect 3580 20430 3620 20470
rect 3980 20430 4020 20470
rect 4380 20430 4420 20470
rect 4780 20430 4820 20470
rect 5180 20430 5220 20470
rect 5580 20430 5620 20470
rect 5980 20430 6020 20470
rect 6380 20430 6420 20470
rect 6780 20430 6820 20470
rect 7180 20430 7220 20470
rect 7580 20430 7620 20470
rect 7980 20430 8020 20470
rect 8380 20430 8420 20470
rect 8780 20430 8820 20470
rect 9180 20430 9220 20470
rect 9580 20430 9620 20470
rect 9980 20430 10020 20470
rect 10380 20430 10420 20470
rect 10780 20430 10820 20470
rect 11180 20430 11220 20470
rect 11580 20430 11620 20470
rect 11980 20430 12020 20470
rect 12380 20430 12420 20470
rect 12780 20430 12820 20470
rect 13180 20430 13220 20470
rect 13580 20430 13620 20470
rect 13980 20430 14020 20470
rect 14380 20430 14420 20470
rect 14780 20430 14820 20470
rect 15180 20430 15220 20470
rect 15580 20430 15620 20470
rect 380 20030 420 20070
rect 780 20030 820 20070
rect 1180 20030 1220 20070
rect 1580 20030 1620 20070
rect 1980 20030 2020 20070
rect 2380 20030 2420 20070
rect 2780 20030 2820 20070
rect 3180 20030 3220 20070
rect 3580 20031 3620 20070
rect 3980 20031 4020 20070
rect 4380 20031 4420 20070
rect 4780 20031 4820 20070
rect 5180 20031 5220 20070
rect 5580 20031 5620 20070
rect 5980 20031 6020 20070
rect 6380 20031 6420 20070
rect 6780 20031 6820 20070
rect 7180 20031 7220 20070
rect 7580 20031 7620 20070
rect 7980 20031 8020 20070
rect 8380 20031 8420 20070
rect 8780 20031 8820 20070
rect 9180 20031 9220 20070
rect 9580 20031 9620 20070
rect 9980 20031 10020 20070
rect 10380 20031 10420 20070
rect 10780 20031 10820 20070
rect 11180 20031 11220 20070
rect 11580 20031 11620 20070
rect 11980 20031 12020 20070
rect 12380 20031 12420 20070
rect 3580 20030 3620 20031
rect 3980 20030 4020 20031
rect 4380 20030 4420 20031
rect 4780 20030 4820 20031
rect 5180 20030 5220 20031
rect 5580 20030 5620 20031
rect 5980 20030 6020 20031
rect 6380 20030 6420 20031
rect 6780 20030 6820 20031
rect 7180 20030 7220 20031
rect 7580 20030 7620 20031
rect 7980 20030 8020 20031
rect 8380 20030 8420 20031
rect 8780 20030 8820 20031
rect 9180 20030 9220 20031
rect 9580 20030 9620 20031
rect 9980 20030 10020 20031
rect 10380 20030 10420 20031
rect 10780 20030 10820 20031
rect 11180 20030 11220 20031
rect 11580 20030 11620 20031
rect 11980 20030 12020 20031
rect 12380 20030 12420 20031
rect 12780 20030 12820 20070
rect 13180 20030 13220 20070
rect 13580 20030 13620 20070
rect 13980 20030 14020 20070
rect 14380 20030 14420 20070
rect 14780 20030 14820 20070
rect 15180 20030 15220 20070
rect 15580 20030 15620 20070
rect 380 19630 420 19670
rect 780 19630 820 19670
rect 1180 19630 1220 19670
rect 1580 19630 1620 19670
rect 1980 19630 2020 19670
rect 2380 19630 2420 19670
rect 2780 19630 2820 19670
rect 3180 19630 3220 19670
rect 3580 19630 3620 19670
rect 3980 19630 4020 19670
rect 4380 19630 4420 19670
rect 4780 19630 4820 19670
rect 5180 19630 5220 19670
rect 5580 19630 5620 19670
rect 5980 19630 6020 19670
rect 6380 19630 6420 19670
rect 6780 19630 6820 19670
rect 7180 19630 7220 19670
rect 7580 19630 7620 19670
rect 7980 19630 8020 19670
rect 8380 19630 8420 19670
rect 8780 19630 8820 19670
rect 9180 19630 9220 19670
rect 9580 19630 9620 19670
rect 9980 19630 10020 19670
rect 10380 19630 10420 19670
rect 10780 19630 10820 19670
rect 11180 19630 11220 19670
rect 11580 19630 11620 19670
rect 11980 19630 12020 19670
rect 12380 19630 12420 19670
rect 12780 19630 12820 19670
rect 13180 19630 13220 19670
rect 13580 19630 13620 19670
rect 13980 19630 14020 19670
rect 14380 19630 14420 19670
rect 14780 19630 14820 19670
rect 15180 19630 15220 19670
rect 15580 19630 15620 19670
rect 380 19230 420 19270
rect 780 19230 820 19270
rect 1180 19230 1220 19270
rect 1580 19230 1620 19270
rect 1980 19230 2020 19270
rect 2380 19230 2420 19270
rect 2780 19230 2820 19270
rect 3180 19230 3220 19270
rect 3580 19230 3620 19270
rect 3980 19230 4020 19270
rect 4380 19230 4420 19270
rect 4780 19230 4820 19270
rect 5180 19230 5220 19270
rect 5580 19230 5620 19270
rect 5980 19230 6020 19270
rect 6380 19230 6420 19270
rect 6780 19230 6820 19270
rect 7180 19230 7220 19270
rect 7580 19230 7620 19270
rect 7980 19230 8020 19270
rect 8380 19230 8420 19270
rect 8780 19230 8820 19270
rect 9180 19230 9220 19270
rect 9580 19230 9620 19270
rect 9980 19230 10020 19270
rect 10380 19230 10420 19270
rect 10780 19230 10820 19270
rect 11180 19230 11220 19270
rect 11580 19230 11620 19270
rect 11980 19230 12020 19270
rect 12380 19230 12420 19270
rect 12780 19230 12820 19270
rect 13180 19230 13220 19270
rect 13580 19230 13620 19270
rect 13980 19230 14020 19270
rect 14380 19230 14420 19270
rect 14780 19230 14820 19270
rect 15180 19230 15220 19270
rect 15580 19230 15620 19270
rect 380 17730 420 17770
rect 780 17730 820 17770
rect 1180 17730 1220 17770
rect 1580 17730 1620 17770
rect 1980 17730 2020 17770
rect 2380 17730 2420 17770
rect 2780 17730 2820 17770
rect 3180 17730 3220 17770
rect 3580 17730 3620 17770
rect 3980 17730 4020 17770
rect 4380 17730 4420 17770
rect 4780 17730 4820 17770
rect 5180 17730 5220 17770
rect 5580 17730 5620 17770
rect 5980 17730 6020 17770
rect 6380 17730 6420 17770
rect 6780 17730 6820 17770
rect 7180 17730 7220 17770
rect 7580 17730 7620 17770
rect 7980 17730 8020 17770
rect 8380 17730 8420 17770
rect 8780 17730 8820 17770
rect 9180 17730 9220 17770
rect 9580 17730 9620 17770
rect 9980 17730 10020 17770
rect 10380 17730 10420 17770
rect 10780 17730 10820 17770
rect 11180 17730 11220 17770
rect 11580 17730 11620 17770
rect 11980 17730 12020 17770
rect 12380 17730 12420 17770
rect 12780 17730 12820 17770
rect 13180 17730 13220 17770
rect 13580 17730 13620 17770
rect 13980 17730 14020 17770
rect 14380 17730 14420 17770
rect 14780 17730 14820 17770
rect 15180 17730 15220 17770
rect 15580 17730 15620 17770
rect 380 17330 420 17370
rect 780 17330 820 17370
rect 1180 17330 1220 17370
rect 1580 17330 1620 17370
rect 1980 17330 2020 17370
rect 2380 17330 2420 17370
rect 2780 17330 2820 17370
rect 3180 17330 3220 17370
rect 3580 17330 3620 17370
rect 3980 17330 4020 17370
rect 4380 17330 4420 17370
rect 4780 17330 4820 17370
rect 5180 17330 5220 17370
rect 5580 17330 5620 17370
rect 5980 17330 6020 17370
rect 6380 17330 6420 17370
rect 6780 17330 6820 17370
rect 7180 17330 7220 17370
rect 7580 17330 7620 17370
rect 7980 17330 8020 17370
rect 8380 17330 8420 17370
rect 8780 17330 8820 17370
rect 9180 17330 9220 17370
rect 9580 17330 9620 17370
rect 9980 17330 10020 17370
rect 10380 17330 10420 17370
rect 10780 17330 10820 17370
rect 11180 17330 11220 17370
rect 11580 17330 11620 17370
rect 11980 17330 12020 17370
rect 12380 17330 12420 17370
rect 12780 17330 12820 17370
rect 13180 17330 13220 17370
rect 13580 17330 13620 17370
rect 13980 17330 14020 17370
rect 14380 17330 14420 17370
rect 14780 17330 14820 17370
rect 15180 17330 15220 17370
rect 15580 17330 15620 17370
rect 380 16930 420 16970
rect 780 16930 820 16970
rect 1180 16930 1220 16970
rect 1580 16930 1620 16970
rect 1980 16930 2020 16970
rect 2380 16930 2420 16970
rect 2780 16930 2820 16970
rect 3180 16930 3220 16970
rect 3580 16930 3620 16970
rect 3980 16930 4020 16970
rect 4380 16930 4420 16970
rect 4780 16930 4820 16970
rect 5180 16930 5220 16970
rect 5580 16930 5620 16970
rect 5980 16930 6020 16970
rect 6380 16930 6420 16970
rect 6780 16930 6820 16970
rect 7180 16930 7220 16970
rect 7580 16930 7620 16970
rect 7980 16930 8020 16970
rect 8380 16930 8420 16970
rect 8780 16930 8820 16970
rect 9180 16930 9220 16970
rect 9580 16930 9620 16970
rect 9980 16930 10020 16970
rect 10380 16930 10420 16970
rect 10780 16930 10820 16970
rect 11180 16930 11220 16970
rect 11580 16930 11620 16970
rect 11980 16930 12020 16970
rect 12380 16930 12420 16970
rect 12780 16930 12820 16970
rect 13180 16930 13220 16970
rect 13580 16930 13620 16970
rect 13980 16930 14020 16970
rect 14380 16930 14420 16970
rect 14780 16930 14820 16970
rect 15180 16930 15220 16970
rect 15580 16930 15620 16970
rect 380 16530 420 16570
rect 780 16530 820 16570
rect 1180 16530 1220 16570
rect 1580 16530 1620 16570
rect 1980 16530 2020 16570
rect 2380 16530 2420 16570
rect 2780 16530 2820 16570
rect 3180 16530 3220 16570
rect 3580 16530 3620 16570
rect 3980 16530 4020 16570
rect 4380 16530 4420 16570
rect 4780 16530 4820 16570
rect 5180 16530 5220 16570
rect 5580 16530 5620 16570
rect 5980 16530 6020 16570
rect 6380 16530 6420 16570
rect 6780 16530 6820 16570
rect 7180 16530 7220 16570
rect 7580 16530 7620 16570
rect 7980 16530 8020 16570
rect 8380 16530 8420 16570
rect 8780 16530 8820 16570
rect 9180 16530 9220 16570
rect 9580 16530 9620 16570
rect 9980 16530 10020 16570
rect 10380 16530 10420 16570
rect 10780 16530 10820 16570
rect 11180 16530 11220 16570
rect 11580 16530 11620 16570
rect 11980 16530 12020 16570
rect 12380 16530 12420 16570
rect 12780 16530 12820 16570
rect 13180 16530 13220 16570
rect 13580 16530 13620 16570
rect 13980 16530 14020 16570
rect 14380 16530 14420 16570
rect 14780 16530 14820 16570
rect 15180 16530 15220 16570
rect 15580 16530 15620 16570
rect 380 16130 420 16170
rect 780 16130 820 16170
rect 1180 16130 1220 16170
rect 1580 16130 1620 16170
rect 1980 16130 2020 16170
rect 2380 16130 2420 16170
rect 2780 16130 2820 16170
rect 3180 16130 3220 16170
rect 3580 16130 3620 16170
rect 3980 16130 4020 16170
rect 4380 16130 4420 16170
rect 4780 16130 4820 16170
rect 5180 16130 5220 16170
rect 5580 16130 5620 16170
rect 5980 16130 6020 16170
rect 6380 16130 6420 16170
rect 6780 16130 6820 16170
rect 7180 16130 7220 16170
rect 7580 16130 7620 16170
rect 7980 16130 8020 16170
rect 8380 16130 8420 16170
rect 8780 16130 8820 16170
rect 9180 16130 9220 16170
rect 9580 16130 9620 16170
rect 9980 16130 10020 16170
rect 10380 16130 10420 16170
rect 10780 16130 10820 16170
rect 11180 16130 11220 16170
rect 11580 16130 11620 16170
rect 11980 16130 12020 16170
rect 12380 16130 12420 16170
rect 12780 16130 12820 16170
rect 13180 16130 13220 16170
rect 13580 16130 13620 16170
rect 13980 16130 14020 16170
rect 14380 16130 14420 16170
rect 14780 16130 14820 16170
rect 15180 16130 15220 16170
rect 15580 16130 15620 16170
rect 380 15730 420 15770
rect 780 15730 820 15770
rect 1180 15730 1220 15770
rect 1580 15730 1620 15770
rect 1980 15730 2020 15770
rect 2380 15730 2420 15770
rect 2780 15730 2820 15770
rect 3180 15730 3220 15770
rect 3580 15730 3620 15770
rect 3980 15730 4020 15770
rect 4380 15730 4420 15770
rect 4780 15730 4820 15770
rect 5180 15730 5220 15770
rect 5580 15730 5620 15770
rect 5980 15730 6020 15770
rect 6380 15730 6420 15770
rect 6780 15730 6820 15770
rect 7180 15730 7220 15770
rect 7580 15730 7620 15770
rect 7980 15730 8020 15770
rect 8380 15730 8420 15770
rect 8780 15730 8820 15770
rect 9180 15730 9220 15770
rect 9580 15730 9620 15770
rect 9980 15730 10020 15770
rect 10380 15730 10420 15770
rect 10780 15730 10820 15770
rect 11180 15730 11220 15770
rect 11580 15730 11620 15770
rect 11980 15730 12020 15770
rect 12380 15730 12420 15770
rect 12780 15730 12820 15770
rect 13180 15730 13220 15770
rect 13580 15730 13620 15770
rect 13980 15730 14020 15770
rect 14380 15730 14420 15770
rect 14780 15730 14820 15770
rect 15180 15730 15220 15770
rect 15580 15730 15620 15770
rect 380 15330 420 15370
rect 780 15330 820 15370
rect 1180 15330 1220 15370
rect 1580 15330 1620 15370
rect 1980 15330 2020 15370
rect 2380 15330 2420 15370
rect 2780 15330 2820 15370
rect 3180 15330 3220 15370
rect 3580 15330 3620 15370
rect 3980 15330 4020 15370
rect 4380 15330 4420 15370
rect 4780 15330 4820 15370
rect 5180 15330 5220 15370
rect 5580 15330 5620 15370
rect 5980 15330 6020 15370
rect 6380 15330 6420 15370
rect 6780 15330 6820 15370
rect 7180 15330 7220 15370
rect 7580 15330 7620 15370
rect 7980 15330 8020 15370
rect 8380 15330 8420 15370
rect 8780 15330 8820 15370
rect 9180 15330 9220 15370
rect 9580 15330 9620 15370
rect 9980 15330 10020 15370
rect 10380 15330 10420 15370
rect 10780 15330 10820 15370
rect 11180 15330 11220 15370
rect 11580 15330 11620 15370
rect 11980 15330 12020 15370
rect 12380 15330 12420 15370
rect 12780 15330 12820 15370
rect 13180 15330 13220 15370
rect 13580 15330 13620 15370
rect 13980 15330 14020 15370
rect 14380 15330 14420 15370
rect 14780 15330 14820 15370
rect 15180 15330 15220 15370
rect 15580 15330 15620 15370
rect 380 14930 420 14970
rect 780 14930 820 14970
rect 1180 14930 1220 14970
rect 1580 14930 1620 14970
rect 1980 14930 2020 14970
rect 2380 14930 2420 14970
rect 2780 14930 2820 14970
rect 3180 14930 3220 14970
rect 3580 14930 3620 14970
rect 3980 14930 4020 14970
rect 4380 14930 4420 14970
rect 4780 14930 4820 14970
rect 5180 14930 5220 14970
rect 5580 14930 5620 14970
rect 5980 14930 6020 14970
rect 6380 14930 6420 14970
rect 6780 14930 6820 14970
rect 7180 14930 7220 14970
rect 7580 14930 7620 14970
rect 7980 14930 8020 14970
rect 8380 14930 8420 14970
rect 8780 14930 8820 14970
rect 9180 14930 9220 14970
rect 9580 14930 9620 14970
rect 9980 14930 10020 14970
rect 10380 14930 10420 14970
rect 10780 14930 10820 14970
rect 11180 14930 11220 14970
rect 11580 14930 11620 14970
rect 11980 14930 12020 14970
rect 12380 14930 12420 14970
rect 12780 14930 12820 14970
rect 13180 14930 13220 14970
rect 13580 14930 13620 14970
rect 13980 14930 14020 14970
rect 14380 14930 14420 14970
rect 14780 14930 14820 14970
rect 15180 14930 15220 14970
rect 15580 14930 15620 14970
rect 380 14530 420 14570
rect 780 14530 820 14570
rect 1180 14530 1220 14570
rect 1580 14530 1620 14570
rect 1980 14530 2020 14570
rect 2380 14530 2420 14570
rect 2780 14530 2820 14570
rect 3180 14530 3220 14570
rect 3580 14530 3620 14570
rect 3980 14530 4020 14570
rect 4380 14530 4420 14570
rect 4780 14530 4820 14570
rect 5180 14530 5220 14570
rect 5580 14530 5620 14570
rect 5980 14530 6020 14570
rect 6380 14530 6420 14570
rect 6780 14530 6820 14570
rect 7180 14530 7220 14570
rect 7580 14530 7620 14570
rect 7980 14530 8020 14570
rect 8380 14530 8420 14570
rect 8780 14530 8820 14570
rect 9180 14530 9220 14570
rect 9580 14530 9620 14570
rect 9980 14530 10020 14570
rect 10380 14530 10420 14570
rect 10780 14530 10820 14570
rect 11180 14530 11220 14570
rect 11580 14530 11620 14570
rect 11980 14530 12020 14570
rect 12380 14530 12420 14570
rect 12780 14530 12820 14570
rect 13180 14530 13220 14570
rect 13580 14530 13620 14570
rect 13980 14530 14020 14570
rect 14380 14530 14420 14570
rect 14780 14530 14820 14570
rect 15180 14530 15220 14570
rect 15580 14530 15620 14570
rect 380 14130 420 14170
rect 780 14130 820 14170
rect 1180 14130 1220 14170
rect 1580 14130 1620 14170
rect 1980 14130 2020 14170
rect 2380 14130 2420 14170
rect 2780 14130 2820 14170
rect 3180 14130 3220 14170
rect 3580 14130 3620 14170
rect 3980 14130 4020 14170
rect 4380 14130 4420 14170
rect 4780 14130 4820 14170
rect 5180 14130 5220 14170
rect 5580 14130 5620 14170
rect 5980 14130 6020 14170
rect 6380 14130 6420 14170
rect 6780 14130 6820 14170
rect 7180 14130 7220 14170
rect 7580 14130 7620 14170
rect 7980 14130 8020 14170
rect 8380 14130 8420 14170
rect 8780 14130 8820 14170
rect 9180 14130 9220 14170
rect 9580 14130 9620 14170
rect 9980 14130 10020 14170
rect 10380 14130 10420 14170
rect 10780 14130 10820 14170
rect 11180 14130 11220 14170
rect 11580 14130 11620 14170
rect 11980 14130 12020 14170
rect 12380 14130 12420 14170
rect 12780 14130 12820 14170
rect 13180 14130 13220 14170
rect 13580 14130 13620 14170
rect 13980 14130 14020 14170
rect 14380 14130 14420 14170
rect 14780 14130 14820 14170
rect 15180 14130 15220 14170
rect 15580 14130 15620 14170
rect 380 13730 420 13770
rect 780 13730 820 13770
rect 1180 13730 1220 13770
rect 1580 13730 1620 13770
rect 1980 13730 2020 13770
rect 2380 13730 2420 13770
rect 2780 13730 2820 13770
rect 3180 13730 3220 13770
rect 3580 13730 3620 13770
rect 3980 13730 4020 13770
rect 4380 13730 4420 13770
rect 4780 13730 4820 13770
rect 5180 13730 5220 13770
rect 5580 13730 5620 13770
rect 5980 13730 6020 13770
rect 6380 13730 6420 13770
rect 6780 13730 6820 13770
rect 7180 13730 7220 13770
rect 7580 13730 7620 13770
rect 7980 13730 8020 13770
rect 8380 13730 8420 13770
rect 8780 13730 8820 13770
rect 9180 13730 9220 13770
rect 9580 13730 9620 13770
rect 9980 13730 10020 13770
rect 10380 13730 10420 13770
rect 10780 13730 10820 13770
rect 11180 13730 11220 13770
rect 11580 13730 11620 13770
rect 11980 13730 12020 13770
rect 12380 13730 12420 13770
rect 12780 13730 12820 13770
rect 13180 13730 13220 13770
rect 13580 13730 13620 13770
rect 13980 13730 14020 13770
rect 14380 13730 14420 13770
rect 14780 13730 14820 13770
rect 15180 13730 15220 13770
rect 15580 13730 15620 13770
rect 380 11430 420 11470
rect 780 11430 820 11470
rect 1180 11430 1220 11470
rect 1580 11430 1620 11470
rect 1980 11430 2020 11470
rect 2380 11430 2420 11470
rect 2780 11430 2820 11470
rect 3180 11430 3220 11470
rect 3580 11430 3620 11470
rect 3980 11430 4020 11470
rect 4380 11430 4420 11470
rect 4780 11430 4820 11470
rect 5180 11430 5220 11470
rect 5580 11430 5620 11470
rect 5980 11430 6020 11470
rect 6380 11430 6420 11470
rect 6780 11430 6820 11470
rect 7180 11430 7220 11470
rect 7580 11430 7620 11470
rect 7980 11430 8020 11470
rect 8380 11430 8420 11470
rect 8780 11430 8820 11470
rect 9180 11430 9220 11470
rect 9580 11430 9620 11470
rect 9980 11430 10020 11470
rect 10380 11430 10420 11470
rect 10780 11430 10820 11470
rect 11180 11430 11220 11470
rect 11580 11430 11620 11470
rect 11980 11430 12020 11470
rect 12380 11430 12420 11470
rect 12780 11430 12820 11470
rect 13180 11430 13220 11470
rect 13580 11430 13620 11470
rect 13980 11430 14020 11470
rect 14380 11430 14420 11470
rect 14780 11430 14820 11470
rect 15180 11430 15220 11470
rect 15580 11430 15620 11470
rect 380 11030 420 11070
rect 780 11030 820 11070
rect 1180 11030 1220 11070
rect 1580 11030 1620 11070
rect 1980 11030 2020 11070
rect 2380 11030 2420 11070
rect 2780 11030 2820 11070
rect 3180 11030 3220 11070
rect 3580 11030 3620 11070
rect 3980 11030 4020 11070
rect 4380 11030 4420 11070
rect 4780 11030 4820 11070
rect 5180 11030 5220 11070
rect 5580 11030 5620 11070
rect 5980 11030 6020 11070
rect 6380 11030 6420 11070
rect 6780 11030 6820 11070
rect 7180 11030 7220 11070
rect 7580 11030 7620 11070
rect 7980 11030 8020 11070
rect 8380 11030 8420 11070
rect 8780 11030 8820 11070
rect 9180 11030 9220 11070
rect 9580 11030 9620 11070
rect 9980 11030 10020 11070
rect 10380 11030 10420 11070
rect 10780 11030 10820 11070
rect 11180 11030 11220 11070
rect 11580 11030 11620 11070
rect 11980 11030 12020 11070
rect 12380 11030 12420 11070
rect 12780 11030 12820 11070
rect 13180 11030 13220 11070
rect 13580 11030 13620 11070
rect 13980 11030 14020 11070
rect 14380 11030 14420 11070
rect 14780 11030 14820 11070
rect 15180 11030 15220 11070
rect 15580 11030 15620 11070
rect 380 10630 420 10670
rect 780 10630 820 10670
rect 1180 10630 1220 10670
rect 1580 10630 1620 10670
rect 1980 10630 2020 10670
rect 2380 10630 2420 10670
rect 2780 10630 2820 10670
rect 3180 10630 3220 10670
rect 3580 10630 3620 10670
rect 3980 10630 4020 10670
rect 4380 10630 4420 10670
rect 4780 10630 4820 10670
rect 5180 10630 5220 10670
rect 5580 10630 5620 10670
rect 5980 10630 6020 10670
rect 6380 10630 6420 10670
rect 6780 10630 6820 10670
rect 7180 10630 7220 10670
rect 7580 10630 7620 10670
rect 7980 10630 8020 10670
rect 8380 10630 8420 10670
rect 8780 10630 8820 10670
rect 9180 10630 9220 10670
rect 9580 10630 9620 10670
rect 9980 10630 10020 10670
rect 10380 10630 10420 10670
rect 10780 10630 10820 10670
rect 11180 10630 11220 10670
rect 11580 10630 11620 10670
rect 11980 10630 12020 10670
rect 12380 10630 12420 10670
rect 12780 10630 12820 10670
rect 13180 10630 13220 10670
rect 13580 10630 13620 10670
rect 13980 10630 14020 10670
rect 14380 10630 14420 10670
rect 14780 10630 14820 10670
rect 15180 10630 15220 10670
rect 15580 10630 15620 10670
rect 380 10230 420 10270
rect 780 10230 820 10270
rect 1180 10230 1220 10270
rect 1580 10230 1620 10270
rect 1980 10230 2020 10270
rect 2380 10230 2420 10270
rect 2780 10230 2820 10270
rect 3180 10230 3220 10270
rect 3580 10230 3620 10270
rect 3980 10230 4020 10270
rect 4380 10230 4420 10270
rect 4780 10230 4820 10270
rect 5180 10230 5220 10270
rect 5580 10230 5620 10270
rect 5980 10230 6020 10270
rect 6380 10230 6420 10270
rect 6780 10230 6820 10270
rect 7180 10230 7220 10270
rect 7580 10230 7620 10270
rect 7980 10230 8020 10270
rect 8380 10230 8420 10270
rect 8780 10230 8820 10270
rect 9180 10230 9220 10270
rect 9580 10230 9620 10270
rect 9980 10230 10020 10270
rect 10380 10230 10420 10270
rect 10780 10230 10820 10270
rect 11180 10230 11220 10270
rect 11580 10230 11620 10270
rect 11980 10230 12020 10270
rect 12380 10230 12420 10270
rect 12780 10230 12820 10270
rect 13180 10230 13220 10270
rect 13580 10230 13620 10270
rect 13980 10230 14020 10270
rect 14380 10230 14420 10270
rect 14780 10230 14820 10270
rect 15180 10230 15220 10270
rect 15580 10230 15620 10270
rect 380 9830 420 9870
rect 780 9830 820 9870
rect 1180 9830 1220 9870
rect 1580 9830 1620 9870
rect 1980 9830 2020 9870
rect 2380 9830 2420 9870
rect 2780 9830 2820 9870
rect 3180 9830 3220 9870
rect 3580 9830 3620 9870
rect 3980 9830 4020 9870
rect 4380 9830 4420 9870
rect 4780 9830 4820 9870
rect 5180 9830 5220 9870
rect 5580 9830 5620 9870
rect 5980 9830 6020 9870
rect 6380 9830 6420 9870
rect 6780 9830 6820 9870
rect 7180 9830 7220 9870
rect 7580 9830 7620 9870
rect 7980 9830 8020 9870
rect 8380 9830 8420 9870
rect 8780 9830 8820 9870
rect 9180 9830 9220 9870
rect 9580 9830 9620 9870
rect 9980 9830 10020 9870
rect 10380 9830 10420 9870
rect 10780 9830 10820 9870
rect 11180 9830 11220 9870
rect 11580 9830 11620 9870
rect 11980 9830 12020 9870
rect 12380 9830 12420 9870
rect 12780 9830 12820 9870
rect 13180 9830 13220 9870
rect 13580 9830 13620 9870
rect 13980 9830 14020 9870
rect 14380 9830 14420 9870
rect 14780 9830 14820 9870
rect 15180 9830 15220 9870
rect 15580 9830 15620 9870
rect 380 9430 420 9470
rect 780 9430 820 9470
rect 1180 9430 1220 9470
rect 1580 9430 1620 9470
rect 1980 9430 2020 9470
rect 2380 9430 2420 9470
rect 2780 9430 2820 9470
rect 3180 9430 3220 9470
rect 3580 9430 3620 9470
rect 3980 9430 4020 9470
rect 4380 9430 4420 9470
rect 4780 9430 4820 9470
rect 5180 9430 5220 9470
rect 5580 9430 5620 9470
rect 5980 9430 6020 9470
rect 6380 9430 6420 9470
rect 6780 9430 6820 9470
rect 7180 9430 7220 9470
rect 7580 9430 7620 9470
rect 7980 9430 8020 9470
rect 8380 9430 8420 9470
rect 8780 9430 8820 9470
rect 9180 9430 9220 9470
rect 9580 9430 9620 9470
rect 9980 9430 10020 9470
rect 10380 9430 10420 9470
rect 10780 9430 10820 9470
rect 11180 9430 11220 9470
rect 11580 9430 11620 9470
rect 11980 9430 12020 9470
rect 12380 9430 12420 9470
rect 12780 9430 12820 9470
rect 13180 9430 13220 9470
rect 13580 9430 13620 9470
rect 13980 9430 14020 9470
rect 14380 9430 14420 9470
rect 14780 9430 14820 9470
rect 15180 9430 15220 9470
rect 15580 9430 15620 9470
rect 380 9030 420 9070
rect 780 9030 820 9070
rect 1180 9030 1220 9070
rect 1580 9030 1620 9070
rect 1980 9030 2020 9070
rect 2380 9030 2420 9070
rect 2780 9030 2820 9070
rect 3180 9030 3220 9070
rect 3580 9030 3620 9070
rect 3980 9030 4020 9070
rect 4380 9030 4420 9070
rect 4780 9030 4820 9070
rect 5180 9030 5220 9070
rect 5580 9030 5620 9070
rect 5980 9030 6020 9070
rect 6380 9030 6420 9070
rect 6780 9030 6820 9070
rect 7180 9030 7220 9070
rect 7580 9030 7620 9070
rect 7980 9030 8020 9070
rect 8380 9030 8420 9070
rect 8780 9030 8820 9070
rect 9180 9030 9220 9070
rect 9580 9030 9620 9070
rect 9980 9030 10020 9070
rect 10380 9030 10420 9070
rect 10780 9030 10820 9070
rect 11180 9030 11220 9070
rect 11580 9030 11620 9070
rect 11980 9030 12020 9070
rect 12380 9030 12420 9070
rect 12780 9030 12820 9070
rect 13180 9030 13220 9070
rect 13580 9030 13620 9070
rect 13980 9030 14020 9070
rect 14380 9030 14420 9070
rect 14780 9030 14820 9070
rect 15180 9030 15220 9070
rect 15580 9030 15620 9070
rect 380 8630 420 8670
rect 780 8630 820 8670
rect 1180 8630 1220 8670
rect 1580 8630 1620 8670
rect 1980 8630 2020 8670
rect 2380 8630 2420 8670
rect 2780 8630 2820 8670
rect 3180 8630 3220 8670
rect 3580 8630 3620 8670
rect 3980 8630 4020 8670
rect 4380 8630 4420 8670
rect 4780 8630 4820 8670
rect 5180 8630 5220 8670
rect 5580 8630 5620 8670
rect 5980 8630 6020 8670
rect 6380 8630 6420 8670
rect 6780 8630 6820 8670
rect 7180 8630 7220 8670
rect 7580 8630 7620 8670
rect 7980 8630 8020 8670
rect 8380 8630 8420 8670
rect 8780 8630 8820 8670
rect 9180 8630 9220 8670
rect 9580 8630 9620 8670
rect 9980 8630 10020 8670
rect 10380 8630 10420 8670
rect 10780 8630 10820 8670
rect 11180 8630 11220 8670
rect 11580 8630 11620 8670
rect 11980 8630 12020 8670
rect 12380 8630 12420 8670
rect 12780 8630 12820 8670
rect 13180 8630 13220 8670
rect 13580 8630 13620 8670
rect 13980 8630 14020 8670
rect 14380 8630 14420 8670
rect 14780 8630 14820 8670
rect 15180 8630 15220 8670
rect 15580 8630 15620 8670
rect 380 8230 420 8270
rect 780 8230 820 8270
rect 1180 8230 1220 8270
rect 1580 8230 1620 8270
rect 1980 8230 2020 8270
rect 2380 8230 2420 8270
rect 2780 8230 2820 8270
rect 3180 8230 3220 8270
rect 3580 8230 3620 8270
rect 3980 8230 4020 8270
rect 4380 8230 4420 8270
rect 4780 8230 4820 8270
rect 5180 8230 5220 8270
rect 5580 8230 5620 8270
rect 5980 8230 6020 8270
rect 6380 8230 6420 8270
rect 6780 8230 6820 8270
rect 7180 8230 7220 8270
rect 7580 8230 7620 8270
rect 7980 8230 8020 8270
rect 8380 8230 8420 8270
rect 8780 8230 8820 8270
rect 9180 8230 9220 8270
rect 9580 8230 9620 8270
rect 9980 8230 10020 8270
rect 10380 8230 10420 8270
rect 10780 8230 10820 8270
rect 11180 8230 11220 8270
rect 11580 8230 11620 8270
rect 11980 8230 12020 8270
rect 12380 8230 12420 8270
rect 12780 8230 12820 8270
rect 13180 8230 13220 8270
rect 13580 8230 13620 8270
rect 13980 8230 14020 8270
rect 14380 8230 14420 8270
rect 14780 8230 14820 8270
rect 15180 8230 15220 8270
rect 15580 8230 15620 8270
rect 380 7830 420 7870
rect 780 7830 820 7870
rect 1180 7830 1220 7870
rect 1580 7830 1620 7870
rect 1980 7830 2020 7870
rect 2380 7830 2420 7870
rect 2780 7830 2820 7870
rect 3180 7830 3220 7870
rect 3580 7830 3620 7870
rect 3980 7830 4020 7870
rect 4380 7830 4420 7870
rect 4780 7830 4820 7870
rect 5180 7830 5220 7870
rect 5580 7830 5620 7870
rect 5980 7830 6020 7870
rect 6380 7830 6420 7870
rect 6780 7830 6820 7870
rect 7180 7830 7220 7870
rect 7580 7830 7620 7870
rect 7980 7830 8020 7870
rect 8380 7830 8420 7870
rect 8780 7830 8820 7870
rect 9180 7830 9220 7870
rect 9580 7830 9620 7870
rect 9980 7830 10020 7870
rect 10380 7830 10420 7870
rect 10780 7830 10820 7870
rect 11180 7830 11220 7870
rect 11580 7830 11620 7870
rect 11980 7830 12020 7870
rect 12380 7830 12420 7870
rect 12780 7830 12820 7870
rect 13180 7830 13220 7870
rect 13580 7830 13620 7870
rect 13980 7830 14020 7870
rect 14380 7830 14420 7870
rect 14780 7830 14820 7870
rect 15180 7830 15220 7870
rect 15580 7830 15620 7870
rect 380 7430 420 7470
rect 780 7430 820 7470
rect 1180 7430 1220 7470
rect 1580 7430 1620 7470
rect 1980 7430 2020 7470
rect 2380 7430 2420 7470
rect 2780 7430 2820 7470
rect 3180 7430 3220 7470
rect 3580 7430 3620 7470
rect 3980 7430 4020 7470
rect 4380 7430 4420 7470
rect 4780 7430 4820 7470
rect 5180 7430 5220 7470
rect 5580 7430 5620 7470
rect 5980 7430 6020 7470
rect 6380 7430 6420 7470
rect 6780 7430 6820 7470
rect 7180 7430 7220 7470
rect 7580 7430 7620 7470
rect 7980 7430 8020 7470
rect 8380 7430 8420 7470
rect 8780 7430 8820 7470
rect 9180 7430 9220 7470
rect 9580 7430 9620 7470
rect 9980 7430 10020 7470
rect 10380 7430 10420 7470
rect 10780 7430 10820 7470
rect 11180 7430 11220 7470
rect 11580 7430 11620 7470
rect 11980 7430 12020 7470
rect 12380 7430 12420 7470
rect 12780 7430 12820 7470
rect 13180 7430 13220 7470
rect 13580 7430 13620 7470
rect 13980 7430 14020 7470
rect 14380 7430 14420 7470
rect 14780 7430 14820 7470
rect 15180 7430 15220 7470
rect 15580 7430 15620 7470
rect 380 5930 420 5970
rect 780 5930 820 5970
rect 1180 5930 1220 5970
rect 1580 5930 1620 5970
rect 1980 5930 2020 5970
rect 2380 5930 2420 5970
rect 2780 5930 2820 5970
rect 3180 5930 3220 5970
rect 3580 5930 3620 5970
rect 3980 5930 4020 5970
rect 4380 5930 4420 5970
rect 4780 5930 4820 5970
rect 5180 5930 5220 5970
rect 5580 5930 5620 5970
rect 5980 5930 6020 5970
rect 6380 5930 6420 5970
rect 6780 5930 6820 5970
rect 7180 5930 7220 5970
rect 7580 5930 7620 5970
rect 7980 5930 8020 5970
rect 8380 5930 8420 5970
rect 8780 5930 8820 5970
rect 9180 5930 9220 5970
rect 9580 5930 9620 5970
rect 9980 5930 10020 5970
rect 10380 5930 10420 5970
rect 10780 5930 10820 5970
rect 11180 5930 11220 5970
rect 11580 5930 11620 5970
rect 11980 5930 12020 5970
rect 12380 5930 12420 5970
rect 12780 5930 12820 5970
rect 13180 5930 13220 5970
rect 13580 5930 13620 5970
rect 13980 5930 14020 5970
rect 14380 5930 14420 5970
rect 14780 5930 14820 5970
rect 15180 5930 15220 5970
rect 15580 5930 15620 5970
rect 380 5530 420 5570
rect 780 5530 820 5570
rect 1180 5530 1220 5570
rect 1580 5530 1620 5570
rect 1980 5530 2020 5570
rect 2380 5530 2420 5570
rect 2780 5530 2820 5570
rect 3180 5530 3220 5570
rect 3580 5530 3620 5570
rect 3980 5530 4020 5570
rect 4380 5530 4420 5570
rect 4780 5530 4820 5570
rect 5180 5530 5220 5570
rect 5580 5530 5620 5570
rect 5980 5530 6020 5570
rect 6380 5530 6420 5570
rect 6780 5530 6820 5570
rect 7180 5530 7220 5570
rect 7580 5530 7620 5570
rect 7980 5530 8020 5570
rect 8380 5530 8420 5570
rect 8780 5530 8820 5570
rect 9180 5530 9220 5570
rect 9580 5530 9620 5570
rect 9980 5530 10020 5570
rect 10380 5530 10420 5570
rect 10780 5530 10820 5570
rect 11180 5530 11220 5570
rect 11580 5530 11620 5570
rect 11980 5530 12020 5570
rect 12380 5530 12420 5570
rect 12780 5530 12820 5570
rect 13180 5530 13220 5570
rect 13580 5530 13620 5570
rect 13980 5530 14020 5570
rect 14380 5530 14420 5570
rect 14780 5530 14820 5570
rect 15180 5530 15220 5570
rect 15580 5530 15620 5570
rect 380 5130 420 5170
rect 780 5130 820 5170
rect 1180 5130 1220 5170
rect 1580 5130 1620 5170
rect 1980 5130 2020 5170
rect 2380 5130 2420 5170
rect 2780 5130 2820 5170
rect 3180 5130 3220 5170
rect 3580 5130 3620 5170
rect 3980 5130 4020 5170
rect 4380 5130 4420 5170
rect 4780 5130 4820 5170
rect 5180 5130 5220 5170
rect 5580 5130 5620 5170
rect 5980 5130 6020 5170
rect 6380 5130 6420 5170
rect 6780 5130 6820 5170
rect 7180 5130 7220 5170
rect 7580 5130 7620 5170
rect 7980 5130 8020 5170
rect 8380 5130 8420 5170
rect 8780 5130 8820 5170
rect 9180 5130 9220 5170
rect 9580 5130 9620 5170
rect 9980 5130 10020 5170
rect 10380 5130 10420 5170
rect 10780 5130 10820 5170
rect 11180 5130 11220 5170
rect 11580 5130 11620 5170
rect 11980 5130 12020 5170
rect 12380 5130 12420 5170
rect 12780 5130 12820 5170
rect 13180 5130 13220 5170
rect 13580 5130 13620 5170
rect 13980 5130 14020 5170
rect 14380 5130 14420 5170
rect 14780 5130 14820 5170
rect 15180 5130 15220 5170
rect 15580 5130 15620 5170
rect 380 4730 420 4770
rect 780 4730 820 4770
rect 1180 4730 1220 4770
rect 1580 4730 1620 4770
rect 1980 4730 2020 4770
rect 2380 4730 2420 4770
rect 2780 4730 2820 4770
rect 3180 4730 3220 4770
rect 3580 4730 3620 4770
rect 3980 4730 4020 4770
rect 4380 4730 4420 4770
rect 4780 4730 4820 4770
rect 5180 4730 5220 4770
rect 5580 4730 5620 4770
rect 5980 4730 6020 4770
rect 6380 4730 6420 4770
rect 6780 4730 6820 4770
rect 7180 4730 7220 4770
rect 7580 4730 7620 4770
rect 7980 4730 8020 4770
rect 8380 4730 8420 4770
rect 8780 4730 8820 4770
rect 9180 4730 9220 4770
rect 9580 4730 9620 4770
rect 9980 4730 10020 4770
rect 10380 4730 10420 4770
rect 10780 4730 10820 4770
rect 11180 4730 11220 4770
rect 11580 4730 11620 4770
rect 11980 4730 12020 4770
rect 12380 4730 12420 4770
rect 12780 4730 12820 4770
rect 13180 4730 13220 4770
rect 13580 4730 13620 4770
rect 13980 4730 14020 4770
rect 14380 4730 14420 4770
rect 14780 4730 14820 4770
rect 15180 4730 15220 4770
rect 15580 4730 15620 4770
rect 380 4330 420 4370
rect 780 4330 820 4370
rect 1180 4330 1220 4370
rect 1580 4330 1620 4370
rect 1980 4330 2020 4370
rect 2380 4330 2420 4370
rect 2780 4330 2820 4370
rect 3180 4330 3220 4370
rect 3580 4330 3620 4370
rect 3980 4330 4020 4370
rect 4380 4330 4420 4370
rect 4780 4330 4820 4370
rect 5180 4330 5220 4370
rect 5580 4330 5620 4370
rect 5980 4330 6020 4370
rect 6380 4330 6420 4370
rect 6780 4330 6820 4370
rect 7180 4330 7220 4370
rect 7580 4330 7620 4370
rect 7980 4330 8020 4370
rect 8380 4330 8420 4370
rect 8780 4330 8820 4370
rect 9180 4330 9220 4370
rect 9580 4330 9620 4370
rect 9980 4330 10020 4370
rect 10380 4330 10420 4370
rect 10780 4330 10820 4370
rect 11180 4330 11220 4370
rect 11580 4330 11620 4370
rect 11980 4330 12020 4370
rect 12380 4330 12420 4370
rect 12780 4330 12820 4370
rect 13180 4330 13220 4370
rect 13580 4330 13620 4370
rect 13980 4330 14020 4370
rect 14380 4330 14420 4370
rect 14780 4330 14820 4370
rect 15180 4330 15220 4370
rect 15580 4330 15620 4370
rect 380 3930 420 3970
rect 780 3930 820 3970
rect 1180 3930 1220 3970
rect 1580 3930 1620 3970
rect 1980 3930 2020 3970
rect 2380 3930 2420 3970
rect 2780 3930 2820 3970
rect 3180 3930 3220 3970
rect 3580 3930 3620 3970
rect 3980 3930 4020 3970
rect 4380 3930 4420 3970
rect 4780 3930 4820 3970
rect 5180 3930 5220 3970
rect 5580 3930 5620 3970
rect 5980 3930 6020 3970
rect 6380 3930 6420 3970
rect 6780 3930 6820 3970
rect 7180 3930 7220 3970
rect 7580 3930 7620 3970
rect 7980 3930 8020 3970
rect 8380 3930 8420 3970
rect 8780 3930 8820 3970
rect 9180 3930 9220 3970
rect 9580 3930 9620 3970
rect 9980 3930 10020 3970
rect 10380 3930 10420 3970
rect 10780 3930 10820 3970
rect 11180 3930 11220 3970
rect 11580 3930 11620 3970
rect 11980 3930 12020 3970
rect 12380 3930 12420 3970
rect 12780 3930 12820 3970
rect 13180 3930 13220 3970
rect 13580 3930 13620 3970
rect 13980 3930 14020 3970
rect 14380 3930 14420 3970
rect 14780 3930 14820 3970
rect 15180 3930 15220 3970
rect 15580 3930 15620 3970
rect 380 3530 420 3570
rect 780 3530 820 3570
rect 1180 3530 1220 3570
rect 1580 3530 1620 3570
rect 1980 3530 2020 3570
rect 2380 3530 2420 3570
rect 2780 3530 2820 3570
rect 3180 3530 3220 3570
rect 3580 3530 3620 3570
rect 3980 3530 4020 3570
rect 4380 3530 4420 3570
rect 4780 3530 4820 3570
rect 5180 3530 5220 3570
rect 5580 3530 5620 3570
rect 5980 3530 6020 3570
rect 6380 3530 6420 3570
rect 6780 3530 6820 3570
rect 7180 3530 7220 3570
rect 7580 3530 7620 3570
rect 7980 3530 8020 3570
rect 8380 3530 8420 3570
rect 8780 3530 8820 3570
rect 9180 3530 9220 3570
rect 9580 3530 9620 3570
rect 9980 3530 10020 3570
rect 10380 3530 10420 3570
rect 10780 3530 10820 3570
rect 11180 3530 11220 3570
rect 11580 3530 11620 3570
rect 11980 3530 12020 3570
rect 12380 3530 12420 3570
rect 12780 3530 12820 3570
rect 13180 3530 13220 3570
rect 13580 3530 13620 3570
rect 13980 3530 14020 3570
rect 14380 3530 14420 3570
rect 14780 3530 14820 3570
rect 15180 3530 15220 3570
rect 15580 3530 15620 3570
rect 380 3130 420 3170
rect 780 3130 820 3170
rect 1180 3130 1220 3170
rect 1580 3130 1620 3170
rect 1980 3130 2020 3170
rect 2380 3130 2420 3170
rect 2780 3130 2820 3170
rect 3180 3130 3220 3170
rect 3580 3130 3620 3170
rect 3980 3130 4020 3170
rect 4380 3130 4420 3170
rect 4780 3130 4820 3170
rect 5180 3130 5220 3170
rect 5580 3130 5620 3170
rect 5980 3130 6020 3170
rect 6380 3130 6420 3170
rect 6780 3130 6820 3170
rect 7180 3130 7220 3170
rect 7580 3130 7620 3170
rect 7980 3130 8020 3170
rect 8380 3130 8420 3170
rect 8780 3130 8820 3170
rect 9180 3130 9220 3170
rect 9580 3130 9620 3170
rect 9980 3130 10020 3170
rect 10380 3130 10420 3170
rect 10780 3130 10820 3170
rect 11180 3130 11220 3170
rect 11580 3130 11620 3170
rect 11980 3130 12020 3170
rect 12380 3130 12420 3170
rect 12780 3130 12820 3170
rect 13180 3130 13220 3170
rect 13580 3130 13620 3170
rect 13980 3130 14020 3170
rect 14380 3130 14420 3170
rect 14780 3130 14820 3170
rect 15180 3130 15220 3170
rect 15580 3130 15620 3170
rect 380 2730 420 2770
rect 780 2730 820 2770
rect 1180 2730 1220 2770
rect 1580 2730 1620 2770
rect 1980 2730 2020 2770
rect 2380 2730 2420 2770
rect 2780 2730 2820 2770
rect 3180 2730 3220 2770
rect 3580 2730 3620 2770
rect 3980 2730 4020 2770
rect 4380 2730 4420 2770
rect 4780 2730 4820 2770
rect 5180 2730 5220 2770
rect 5580 2730 5620 2770
rect 5980 2730 6020 2770
rect 6380 2730 6420 2770
rect 6780 2730 6820 2770
rect 7180 2730 7220 2770
rect 7580 2730 7620 2770
rect 7980 2730 8020 2770
rect 8380 2730 8420 2770
rect 8780 2730 8820 2770
rect 9180 2730 9220 2770
rect 9580 2730 9620 2770
rect 9980 2730 10020 2770
rect 10380 2730 10420 2770
rect 10780 2730 10820 2770
rect 11180 2730 11220 2770
rect 11580 2730 11620 2770
rect 11980 2730 12020 2770
rect 12380 2730 12420 2770
rect 12780 2730 12820 2770
rect 13180 2730 13220 2770
rect 13580 2730 13620 2770
rect 13980 2730 14020 2770
rect 14380 2730 14420 2770
rect 14780 2730 14820 2770
rect 15180 2730 15220 2770
rect 15580 2730 15620 2770
rect 380 2330 420 2370
rect 780 2330 820 2370
rect 1180 2330 1220 2370
rect 1580 2330 1620 2370
rect 1980 2330 2020 2370
rect 2380 2330 2420 2370
rect 2780 2330 2820 2370
rect 3180 2330 3220 2370
rect 3580 2330 3620 2370
rect 3980 2330 4020 2370
rect 4380 2330 4420 2370
rect 4780 2330 4820 2370
rect 5180 2330 5220 2370
rect 5580 2330 5620 2370
rect 5980 2330 6020 2370
rect 6380 2330 6420 2370
rect 6780 2330 6820 2370
rect 7180 2330 7220 2370
rect 7580 2330 7620 2370
rect 7980 2330 8020 2370
rect 8380 2330 8420 2370
rect 8780 2330 8820 2370
rect 9180 2330 9220 2370
rect 9580 2330 9620 2370
rect 9980 2330 10020 2370
rect 10380 2330 10420 2370
rect 10780 2330 10820 2370
rect 11180 2330 11220 2370
rect 11580 2330 11620 2370
rect 11980 2330 12020 2370
rect 12380 2330 12420 2370
rect 12780 2330 12820 2370
rect 13180 2330 13220 2370
rect 13580 2330 13620 2370
rect 13980 2330 14020 2370
rect 14380 2330 14420 2370
rect 14780 2330 14820 2370
rect 15180 2330 15220 2370
rect 15580 2330 15620 2370
rect 380 1930 420 1970
rect 780 1930 820 1970
rect 1180 1930 1220 1970
rect 1580 1930 1620 1970
rect 1980 1930 2020 1970
rect 2380 1930 2420 1970
rect 2780 1930 2820 1970
rect 3180 1930 3220 1970
rect 3580 1930 3620 1970
rect 3980 1930 4020 1970
rect 4380 1930 4420 1970
rect 4780 1930 4820 1970
rect 5180 1930 5220 1970
rect 5580 1930 5620 1970
rect 5980 1930 6020 1970
rect 6380 1930 6420 1970
rect 6780 1930 6820 1970
rect 7180 1930 7220 1970
rect 7580 1930 7620 1970
rect 7980 1930 8020 1970
rect 8380 1930 8420 1970
rect 8780 1930 8820 1970
rect 9180 1930 9220 1970
rect 9580 1930 9620 1970
rect 9980 1930 10020 1970
rect 10380 1930 10420 1970
rect 10780 1930 10820 1970
rect 11180 1930 11220 1970
rect 11580 1930 11620 1970
rect 11980 1930 12020 1970
rect 12380 1930 12420 1970
rect 12780 1930 12820 1970
rect 13180 1930 13220 1970
rect 13580 1930 13620 1970
rect 13980 1930 14020 1970
rect 14380 1930 14420 1970
rect 14780 1930 14820 1970
rect 15180 1930 15220 1970
rect 15580 1930 15620 1970
rect 1180 480 1220 520
rect 1580 480 1620 520
rect 1980 480 2020 520
rect 2380 480 2420 520
rect 2780 480 2820 520
rect 3180 480 3220 520
rect 3580 480 3620 520
rect 3980 480 4020 520
rect 4380 480 4420 520
rect 4780 480 4820 520
rect 5180 480 5220 520
rect 5580 480 5620 520
rect 5980 480 6020 520
rect 6380 480 6420 520
rect 6780 480 6820 520
rect 7180 480 7220 520
rect 7580 480 7620 520
rect 7980 480 8020 520
rect 8380 480 8420 520
rect 8780 480 8820 520
rect 9180 480 9220 520
rect 9580 480 9620 520
rect 9980 480 10020 520
rect 10380 480 10420 520
rect 10780 480 10820 520
rect 11180 480 11220 520
rect 11580 480 11620 520
rect 11980 480 12020 520
rect 12380 480 12420 520
rect 12780 480 12820 520
rect 13180 480 13220 520
rect 13580 480 13620 520
rect 13980 480 14020 520
rect 14380 480 14420 520
rect 14780 480 14820 520
rect 1180 80 1220 120
rect 1580 80 1620 120
rect 1980 80 2020 120
rect 2380 80 2420 120
rect 2780 80 2820 120
rect 3180 80 3220 120
rect 3580 80 3620 120
rect 3980 80 4020 120
rect 4380 80 4420 120
rect 4780 80 4820 120
rect 5180 80 5220 120
rect 5580 80 5620 120
rect 5980 80 6020 120
rect 6380 80 6420 120
rect 6780 80 6820 120
rect 7180 80 7220 120
rect 7580 80 7620 120
rect 7980 80 8020 120
rect 8380 80 8420 120
rect 8780 80 8820 120
rect 9180 80 9220 120
rect 9580 80 9620 120
rect 9980 80 10020 120
rect 10380 80 10420 120
rect 10780 80 10820 120
rect 11180 80 11220 120
rect 11580 80 11620 120
rect 11980 80 12020 120
rect 12380 80 12420 120
rect 12780 80 12820 120
rect 13180 80 13220 120
rect 13580 80 13620 120
rect 13980 80 14020 120
rect 14380 80 14420 120
rect 14780 80 14820 120
<< metal4 >>
rect 0 35040 16000 35600
rect 0 35000 380 35040
rect 420 35000 780 35040
rect 820 35000 1180 35040
rect 1220 35000 1580 35040
rect 1620 35000 1980 35040
rect 2020 35000 2380 35040
rect 2420 35000 2780 35040
rect 2820 35000 3180 35040
rect 3220 35000 3580 35040
rect 3620 35000 3980 35040
rect 4020 35000 4380 35040
rect 4420 35000 4780 35040
rect 4820 35000 5180 35040
rect 5220 35000 5580 35040
rect 5620 35000 5980 35040
rect 6020 35000 6380 35040
rect 6420 35000 6780 35040
rect 6820 35000 7180 35040
rect 7220 35000 7580 35040
rect 7620 35000 7980 35040
rect 8020 35000 8380 35040
rect 8420 35000 8780 35040
rect 8820 35000 9180 35040
rect 9220 35000 9580 35040
rect 9620 35000 9980 35040
rect 10020 35000 10380 35040
rect 10420 35000 10780 35040
rect 10820 35000 11180 35040
rect 11220 35000 11580 35040
rect 11620 35000 11980 35040
rect 12020 35000 12380 35040
rect 12420 35000 12780 35040
rect 12820 35000 13180 35040
rect 13220 35000 13580 35040
rect 13620 35000 13980 35040
rect 14020 35000 14380 35040
rect 14420 35000 14780 35040
rect 14820 35000 15180 35040
rect 15220 35000 15580 35040
rect 15620 35000 16000 35040
rect 0 34640 16000 35000
rect 0 34600 380 34640
rect 420 34600 780 34640
rect 820 34600 1180 34640
rect 1220 34600 1580 34640
rect 1620 34600 1980 34640
rect 2020 34600 2380 34640
rect 2420 34600 2780 34640
rect 2820 34600 3180 34640
rect 3220 34600 3580 34640
rect 3620 34600 3980 34640
rect 4020 34600 4380 34640
rect 4420 34600 4780 34640
rect 4820 34600 5180 34640
rect 5220 34600 5580 34640
rect 5620 34600 5980 34640
rect 6020 34600 6380 34640
rect 6420 34600 6780 34640
rect 6820 34600 7180 34640
rect 7220 34600 7580 34640
rect 7620 34600 7980 34640
rect 8020 34600 8380 34640
rect 8420 34600 8780 34640
rect 8820 34600 9180 34640
rect 9220 34600 9580 34640
rect 9620 34600 9980 34640
rect 10020 34600 10380 34640
rect 10420 34600 10780 34640
rect 10820 34600 11180 34640
rect 11220 34600 11580 34640
rect 11620 34600 11980 34640
rect 12020 34600 12380 34640
rect 12420 34600 12780 34640
rect 12820 34600 13180 34640
rect 13220 34600 13580 34640
rect 13620 34600 13980 34640
rect 14020 34600 14380 34640
rect 14420 34600 14780 34640
rect 14820 34600 15180 34640
rect 15220 34600 15580 34640
rect 15620 34600 16000 34640
rect 0 34240 16000 34600
rect 0 34200 380 34240
rect 420 34200 780 34240
rect 820 34200 1180 34240
rect 1220 34200 1580 34240
rect 1620 34200 1980 34240
rect 2020 34200 2380 34240
rect 2420 34200 2780 34240
rect 2820 34200 3180 34240
rect 3220 34200 3580 34240
rect 3620 34200 3980 34240
rect 4020 34200 4380 34240
rect 4420 34200 4780 34240
rect 4820 34200 5180 34240
rect 5220 34200 5580 34240
rect 5620 34200 5980 34240
rect 6020 34200 6380 34240
rect 6420 34200 6780 34240
rect 6820 34200 7180 34240
rect 7220 34200 7580 34240
rect 7620 34200 7980 34240
rect 8020 34200 8380 34240
rect 8420 34200 8780 34240
rect 8820 34200 9180 34240
rect 9220 34200 9580 34240
rect 9620 34200 9980 34240
rect 10020 34200 10380 34240
rect 10420 34200 10780 34240
rect 10820 34200 11180 34240
rect 11220 34200 11580 34240
rect 11620 34200 11980 34240
rect 12020 34200 12380 34240
rect 12420 34200 12780 34240
rect 12820 34200 13180 34240
rect 13220 34200 13580 34240
rect 13620 34200 13980 34240
rect 14020 34200 14380 34240
rect 14420 34200 14780 34240
rect 14820 34200 15180 34240
rect 15220 34200 15580 34240
rect 15620 34200 16000 34240
rect 0 33840 16000 34200
rect 0 33800 380 33840
rect 420 33800 780 33840
rect 820 33800 1180 33840
rect 1220 33800 1580 33840
rect 1620 33800 1980 33840
rect 2020 33800 2380 33840
rect 2420 33800 2780 33840
rect 2820 33800 3180 33840
rect 3220 33800 3580 33840
rect 3620 33800 3980 33840
rect 4020 33800 4380 33840
rect 4420 33800 4780 33840
rect 4820 33800 5180 33840
rect 5220 33800 5580 33840
rect 5620 33800 5980 33840
rect 6020 33800 6380 33840
rect 6420 33800 6780 33840
rect 6820 33800 7180 33840
rect 7220 33800 7580 33840
rect 7620 33800 7980 33840
rect 8020 33800 8380 33840
rect 8420 33800 8780 33840
rect 8820 33800 9180 33840
rect 9220 33800 9580 33840
rect 9620 33800 9980 33840
rect 10020 33800 10380 33840
rect 10420 33800 10780 33840
rect 10820 33800 11180 33840
rect 11220 33800 11580 33840
rect 11620 33800 11980 33840
rect 12020 33800 12380 33840
rect 12420 33800 12780 33840
rect 12820 33800 13180 33840
rect 13220 33800 13580 33840
rect 13620 33800 13980 33840
rect 14020 33800 14380 33840
rect 14420 33800 14780 33840
rect 14820 33800 15180 33840
rect 15220 33800 15580 33840
rect 15620 33800 16000 33840
rect 0 33440 16000 33800
rect 0 33400 380 33440
rect 420 33400 780 33440
rect 820 33400 1180 33440
rect 1220 33400 1580 33440
rect 1620 33400 1980 33440
rect 2020 33400 2380 33440
rect 2420 33400 2780 33440
rect 2820 33400 3180 33440
rect 3220 33400 3580 33440
rect 3620 33400 3980 33440
rect 4020 33400 4380 33440
rect 4420 33400 4780 33440
rect 4820 33400 5180 33440
rect 5220 33400 5580 33440
rect 5620 33400 5980 33440
rect 6020 33400 6380 33440
rect 6420 33400 6780 33440
rect 6820 33400 7180 33440
rect 7220 33400 7580 33440
rect 7620 33400 7980 33440
rect 8020 33400 8380 33440
rect 8420 33400 8780 33440
rect 8820 33400 9180 33440
rect 9220 33400 9580 33440
rect 9620 33400 9980 33440
rect 10020 33400 10380 33440
rect 10420 33400 10780 33440
rect 10820 33400 11180 33440
rect 11220 33400 11580 33440
rect 11620 33400 11980 33440
rect 12020 33400 12380 33440
rect 12420 33400 12780 33440
rect 12820 33400 13180 33440
rect 13220 33400 13580 33440
rect 13620 33400 13980 33440
rect 14020 33400 14380 33440
rect 14420 33400 14780 33440
rect 14820 33400 15180 33440
rect 15220 33400 15580 33440
rect 15620 33400 16000 33440
rect 0 33040 16000 33400
rect 0 33000 380 33040
rect 420 33000 780 33040
rect 820 33000 1180 33040
rect 1220 33000 1580 33040
rect 1620 33000 1980 33040
rect 2020 33000 2380 33040
rect 2420 33000 2780 33040
rect 2820 33000 3180 33040
rect 3220 33000 3580 33040
rect 3620 33000 3980 33040
rect 4020 33000 4380 33040
rect 4420 33000 4780 33040
rect 4820 33000 5180 33040
rect 5220 33000 5580 33040
rect 5620 33000 5980 33040
rect 6020 33000 6380 33040
rect 6420 33000 6780 33040
rect 6820 33000 7180 33040
rect 7220 33000 7580 33040
rect 7620 33000 7980 33040
rect 8020 33000 8380 33040
rect 8420 33000 8780 33040
rect 8820 33000 9180 33040
rect 9220 33000 9580 33040
rect 9620 33000 9980 33040
rect 10020 33000 10380 33040
rect 10420 33000 10780 33040
rect 10820 33000 11180 33040
rect 11220 33000 11580 33040
rect 11620 33000 11980 33040
rect 12020 33000 12380 33040
rect 12420 33000 12780 33040
rect 12820 33000 13180 33040
rect 13220 33000 13580 33040
rect 13620 33000 13980 33040
rect 14020 33000 14380 33040
rect 14420 33000 14780 33040
rect 14820 33000 15180 33040
rect 15220 33000 15580 33040
rect 15620 33000 16000 33040
rect 0 32440 16000 33000
rect 200 32000 249 32040
rect 7751 32000 7800 32040
rect 200 31160 7800 32000
rect 8200 31600 15800 32440
rect 8200 31560 8249 31600
rect 15751 31560 15800 31600
rect 0 30600 16000 31160
rect 0 30560 380 30600
rect 420 30560 780 30600
rect 820 30560 1180 30600
rect 1220 30560 1580 30600
rect 1620 30560 1980 30600
rect 2020 30560 2380 30600
rect 2420 30560 2780 30600
rect 2820 30560 3180 30600
rect 3220 30560 3580 30600
rect 3620 30560 3980 30600
rect 4020 30560 4380 30600
rect 4420 30560 4780 30600
rect 4820 30560 5180 30600
rect 5220 30560 5580 30600
rect 5620 30560 5980 30600
rect 6020 30560 6380 30600
rect 6420 30560 6780 30600
rect 6820 30560 7180 30600
rect 7220 30560 7580 30600
rect 7620 30560 7980 30600
rect 8020 30560 8380 30600
rect 8420 30560 8780 30600
rect 8820 30560 9180 30600
rect 9220 30560 9580 30600
rect 9620 30560 9980 30600
rect 10020 30560 10380 30600
rect 10420 30560 10780 30600
rect 10820 30560 11180 30600
rect 11220 30560 11580 30600
rect 11620 30560 11980 30600
rect 12020 30560 12380 30600
rect 12420 30560 12780 30600
rect 12820 30560 13180 30600
rect 13220 30560 13580 30600
rect 13620 30560 13980 30600
rect 14020 30560 14380 30600
rect 14420 30560 14780 30600
rect 14820 30560 15180 30600
rect 15220 30560 15580 30600
rect 15620 30560 16000 30600
rect 0 30200 16000 30560
rect 0 30160 380 30200
rect 420 30160 780 30200
rect 820 30160 1180 30200
rect 1220 30160 1580 30200
rect 1620 30160 1980 30200
rect 2020 30160 2380 30200
rect 2420 30160 2780 30200
rect 2820 30160 3180 30200
rect 3220 30160 3580 30200
rect 3620 30160 3980 30200
rect 4020 30160 4380 30200
rect 4420 30160 4780 30200
rect 4820 30160 5180 30200
rect 5220 30160 5580 30200
rect 5620 30160 5980 30200
rect 6020 30160 6380 30200
rect 6420 30160 6780 30200
rect 6820 30160 7180 30200
rect 7220 30160 7580 30200
rect 7620 30160 7980 30200
rect 8020 30160 8380 30200
rect 8420 30160 8780 30200
rect 8820 30160 9180 30200
rect 9220 30160 9580 30200
rect 9620 30160 9980 30200
rect 10020 30160 10380 30200
rect 10420 30160 10780 30200
rect 10820 30160 11180 30200
rect 11220 30160 11580 30200
rect 11620 30160 11980 30200
rect 12020 30160 12380 30200
rect 12420 30160 12780 30200
rect 12820 30160 13180 30200
rect 13220 30160 13580 30200
rect 13620 30160 13980 30200
rect 14020 30160 14380 30200
rect 14420 30160 14780 30200
rect 14820 30160 15180 30200
rect 15220 30160 15580 30200
rect 15620 30160 16000 30200
rect 0 29800 16000 30160
rect 0 29760 380 29800
rect 420 29760 780 29800
rect 820 29760 1180 29800
rect 1220 29760 1580 29800
rect 1620 29760 1980 29800
rect 2020 29760 2380 29800
rect 2420 29760 2780 29800
rect 2820 29760 3180 29800
rect 3220 29760 3580 29800
rect 3620 29760 3980 29800
rect 4020 29760 4380 29800
rect 4420 29760 4780 29800
rect 4820 29760 5180 29800
rect 5220 29760 5580 29800
rect 5620 29760 5980 29800
rect 6020 29760 6380 29800
rect 6420 29760 6780 29800
rect 6820 29760 7180 29800
rect 7220 29760 7580 29800
rect 7620 29760 7980 29800
rect 8020 29760 8380 29800
rect 8420 29760 8780 29800
rect 8820 29760 9180 29800
rect 9220 29760 9580 29800
rect 9620 29760 9980 29800
rect 10020 29760 10380 29800
rect 10420 29760 10780 29800
rect 10820 29760 11180 29800
rect 11220 29760 11580 29800
rect 11620 29760 11980 29800
rect 12020 29760 12380 29800
rect 12420 29760 12780 29800
rect 12820 29760 13180 29800
rect 13220 29760 13580 29800
rect 13620 29760 13980 29800
rect 14020 29760 14380 29800
rect 14420 29760 14780 29800
rect 14820 29760 15180 29800
rect 15220 29760 15580 29800
rect 15620 29760 16000 29800
rect 0 29400 16000 29760
rect 0 29360 380 29400
rect 420 29360 780 29400
rect 820 29360 1180 29400
rect 1220 29360 1580 29400
rect 1620 29360 1980 29400
rect 2020 29360 2380 29400
rect 2420 29360 2780 29400
rect 2820 29360 3180 29400
rect 3220 29360 3580 29400
rect 3620 29360 3980 29400
rect 4020 29360 4380 29400
rect 4420 29360 4780 29400
rect 4820 29360 5180 29400
rect 5220 29360 5580 29400
rect 5620 29360 5980 29400
rect 6020 29360 6380 29400
rect 6420 29360 6780 29400
rect 6820 29360 7180 29400
rect 7220 29360 7580 29400
rect 7620 29360 7980 29400
rect 8020 29360 8380 29400
rect 8420 29360 8780 29400
rect 8820 29360 9180 29400
rect 9220 29360 9580 29400
rect 9620 29360 9980 29400
rect 10020 29360 10380 29400
rect 10420 29360 10780 29400
rect 10820 29360 11180 29400
rect 11220 29360 11580 29400
rect 11620 29360 11980 29400
rect 12020 29360 12380 29400
rect 12420 29360 12780 29400
rect 12820 29360 13180 29400
rect 13220 29360 13580 29400
rect 13620 29360 13980 29400
rect 14020 29360 14380 29400
rect 14420 29360 14780 29400
rect 14820 29360 15180 29400
rect 15220 29360 15580 29400
rect 15620 29360 16000 29400
rect 0 29000 16000 29360
rect 0 28960 380 29000
rect 420 28960 780 29000
rect 820 28960 1180 29000
rect 1220 28960 1580 29000
rect 1620 28960 1980 29000
rect 2020 28960 2380 29000
rect 2420 28960 2780 29000
rect 2820 28960 3180 29000
rect 3220 28960 3580 29000
rect 3620 28960 3980 29000
rect 4020 28960 4380 29000
rect 4420 28960 4780 29000
rect 4820 28960 5180 29000
rect 5220 28960 5580 29000
rect 5620 28960 5980 29000
rect 6020 28960 6380 29000
rect 6420 28960 6780 29000
rect 6820 28960 7180 29000
rect 7220 28960 7580 29000
rect 7620 28960 7980 29000
rect 8020 28960 8380 29000
rect 8420 28960 8780 29000
rect 8820 28960 9180 29000
rect 9220 28960 9580 29000
rect 9620 28960 9980 29000
rect 10020 28960 10380 29000
rect 10420 28960 10780 29000
rect 10820 28960 11180 29000
rect 11220 28960 11580 29000
rect 11620 28960 11980 29000
rect 12020 28960 12380 29000
rect 12420 28960 12780 29000
rect 12820 28960 13180 29000
rect 13220 28960 13580 29000
rect 13620 28960 13980 29000
rect 14020 28960 14380 29000
rect 14420 28960 14780 29000
rect 14820 28960 15180 29000
rect 15220 28960 15580 29000
rect 15620 28960 16000 29000
rect 0 28600 16000 28960
rect 0 28560 380 28600
rect 420 28560 780 28600
rect 820 28560 1180 28600
rect 1220 28560 1580 28600
rect 1620 28560 1980 28600
rect 2020 28560 2380 28600
rect 2420 28560 2780 28600
rect 2820 28560 3180 28600
rect 3220 28560 3580 28600
rect 3620 28560 3980 28600
rect 4020 28560 4380 28600
rect 4420 28560 4780 28600
rect 4820 28560 5180 28600
rect 5220 28560 5580 28600
rect 5620 28560 5980 28600
rect 6020 28560 6380 28600
rect 6420 28560 6780 28600
rect 6820 28560 7180 28600
rect 7220 28560 7580 28600
rect 7620 28560 7980 28600
rect 8020 28560 8380 28600
rect 8420 28560 8780 28600
rect 8820 28560 9180 28600
rect 9220 28560 9580 28600
rect 9620 28560 9980 28600
rect 10020 28560 10380 28600
rect 10420 28560 10780 28600
rect 10820 28560 11180 28600
rect 11220 28560 11580 28600
rect 11620 28560 11980 28600
rect 12020 28560 12380 28600
rect 12420 28560 12780 28600
rect 12820 28560 13180 28600
rect 13220 28560 13580 28600
rect 13620 28560 13980 28600
rect 14020 28560 14380 28600
rect 14420 28560 14780 28600
rect 14820 28560 15180 28600
rect 15220 28560 15580 28600
rect 15620 28560 16000 28600
rect 0 28000 16000 28560
rect 0 26420 16000 26800
rect 0 26380 380 26420
rect 420 26380 780 26420
rect 820 26380 1180 26420
rect 1220 26380 1580 26420
rect 1620 26380 1980 26420
rect 2020 26380 2380 26420
rect 2420 26380 2780 26420
rect 2820 26380 3180 26420
rect 3220 26380 3580 26420
rect 3620 26380 3980 26420
rect 4020 26380 4380 26420
rect 4420 26380 4780 26420
rect 4820 26380 5180 26420
rect 5220 26380 5580 26420
rect 5620 26380 5980 26420
rect 6020 26380 6380 26420
rect 6420 26380 6780 26420
rect 6820 26380 7180 26420
rect 7220 26380 7580 26420
rect 7620 26380 7980 26420
rect 8020 26380 8380 26420
rect 8420 26380 8780 26420
rect 8820 26380 9180 26420
rect 9220 26380 9580 26420
rect 9620 26380 9980 26420
rect 10020 26380 10380 26420
rect 10420 26380 10780 26420
rect 10820 26380 11180 26420
rect 11220 26380 11580 26420
rect 11620 26380 11980 26420
rect 12020 26380 12380 26420
rect 12420 26380 12780 26420
rect 12820 26380 13180 26420
rect 13220 26380 13580 26420
rect 13620 26380 13980 26420
rect 14020 26380 14380 26420
rect 14420 26380 14780 26420
rect 14820 26380 15180 26420
rect 15220 26380 15580 26420
rect 15620 26380 16000 26420
rect 0 26020 16000 26380
rect 0 25980 380 26020
rect 420 25980 780 26020
rect 820 25980 1180 26020
rect 1220 25980 1580 26020
rect 1620 25980 1980 26020
rect 2020 25980 2380 26020
rect 2420 25980 2780 26020
rect 2820 25980 3180 26020
rect 3220 25980 3580 26020
rect 3620 25980 3980 26020
rect 4020 25980 4380 26020
rect 4420 25980 4780 26020
rect 4820 25980 5180 26020
rect 5220 25980 5580 26020
rect 5620 25980 5980 26020
rect 6020 25980 6380 26020
rect 6420 25980 6780 26020
rect 6820 25980 7180 26020
rect 7220 25980 7580 26020
rect 7620 25980 7980 26020
rect 8020 25980 8380 26020
rect 8420 25980 8780 26020
rect 8820 25980 9180 26020
rect 9220 25980 9580 26020
rect 9620 25980 9980 26020
rect 10020 25980 10380 26020
rect 10420 25980 10780 26020
rect 10820 25980 11180 26020
rect 11220 25980 11580 26020
rect 11620 25980 11980 26020
rect 12020 25980 12380 26020
rect 12420 25980 12780 26020
rect 12820 25980 13180 26020
rect 13220 25980 13580 26020
rect 13620 25980 13980 26020
rect 14020 25980 14380 26020
rect 14420 25980 14780 26020
rect 14820 25980 15180 26020
rect 15220 25980 15580 26020
rect 15620 25980 16000 26020
rect 0 25620 16000 25980
rect 0 25580 380 25620
rect 420 25580 780 25620
rect 820 25580 1180 25620
rect 1220 25580 1580 25620
rect 1620 25580 1980 25620
rect 2020 25580 2380 25620
rect 2420 25580 2780 25620
rect 2820 25580 3180 25620
rect 3220 25580 3580 25620
rect 3620 25580 3980 25620
rect 4020 25580 4380 25620
rect 4420 25580 4780 25620
rect 4820 25580 5180 25620
rect 5220 25580 5580 25620
rect 5620 25580 5980 25620
rect 6020 25580 6380 25620
rect 6420 25580 6780 25620
rect 6820 25580 7180 25620
rect 7220 25580 7580 25620
rect 7620 25580 7980 25620
rect 8020 25580 8380 25620
rect 8420 25580 8780 25620
rect 8820 25580 9180 25620
rect 9220 25580 9580 25620
rect 9620 25580 9980 25620
rect 10020 25580 10380 25620
rect 10420 25580 10780 25620
rect 10820 25580 11180 25620
rect 11220 25580 11580 25620
rect 11620 25580 11980 25620
rect 12020 25580 12380 25620
rect 12420 25580 12780 25620
rect 12820 25580 13180 25620
rect 13220 25580 13580 25620
rect 13620 25580 13980 25620
rect 14020 25580 14380 25620
rect 14420 25580 14780 25620
rect 14820 25580 15180 25620
rect 15220 25580 15580 25620
rect 15620 25580 16000 25620
rect 0 25200 16000 25580
rect 0 23270 16000 23800
rect 0 23230 380 23270
rect 420 23230 780 23270
rect 820 23230 1180 23270
rect 1220 23230 1580 23270
rect 1620 23230 1980 23270
rect 2020 23230 2380 23270
rect 2420 23230 2780 23270
rect 2820 23230 3180 23270
rect 3220 23230 3580 23270
rect 3620 23230 3980 23270
rect 4020 23230 4380 23270
rect 4420 23230 4780 23270
rect 4820 23230 5180 23270
rect 5220 23230 5580 23270
rect 5620 23230 5980 23270
rect 6020 23230 6380 23270
rect 6420 23230 6780 23270
rect 6820 23230 7180 23270
rect 7220 23230 7580 23270
rect 7620 23230 7980 23270
rect 8020 23230 8380 23270
rect 8420 23230 8780 23270
rect 8820 23230 9180 23270
rect 9220 23230 9580 23270
rect 9620 23230 9980 23270
rect 10020 23230 10380 23270
rect 10420 23230 10780 23270
rect 10820 23230 11180 23270
rect 11220 23230 11580 23270
rect 11620 23230 11980 23270
rect 12020 23230 12380 23270
rect 12420 23230 12780 23270
rect 12820 23230 13180 23270
rect 13220 23230 13580 23270
rect 13620 23230 13980 23270
rect 14020 23230 14380 23270
rect 14420 23230 14780 23270
rect 14820 23230 15180 23270
rect 15220 23230 15580 23270
rect 15620 23230 16000 23270
rect 0 22870 16000 23230
rect 0 22830 380 22870
rect 420 22830 780 22870
rect 820 22830 1180 22870
rect 1220 22830 1580 22870
rect 1620 22830 1980 22870
rect 2020 22830 2380 22870
rect 2420 22830 2780 22870
rect 2820 22830 3180 22870
rect 3220 22830 3580 22870
rect 3620 22830 3980 22870
rect 4020 22830 4380 22870
rect 4420 22830 4780 22870
rect 4820 22830 5180 22870
rect 5220 22830 5580 22870
rect 5620 22830 5980 22870
rect 6020 22830 6380 22870
rect 6420 22830 6780 22870
rect 6820 22830 7180 22870
rect 7220 22830 7580 22870
rect 7620 22830 7980 22870
rect 8020 22830 8380 22870
rect 8420 22830 8780 22870
rect 8820 22830 9180 22870
rect 9220 22830 9580 22870
rect 9620 22830 9980 22870
rect 10020 22830 10380 22870
rect 10420 22830 10780 22870
rect 10820 22830 11180 22870
rect 11220 22830 11580 22870
rect 11620 22830 11980 22870
rect 12020 22830 12380 22870
rect 12420 22830 12780 22870
rect 12820 22830 13180 22870
rect 13220 22830 13580 22870
rect 13620 22830 13980 22870
rect 14020 22830 14380 22870
rect 14420 22830 14780 22870
rect 14820 22830 15180 22870
rect 15220 22830 15580 22870
rect 15620 22830 16000 22870
rect 0 22470 16000 22830
rect 0 22430 380 22470
rect 420 22430 780 22470
rect 820 22430 1180 22470
rect 1220 22430 1580 22470
rect 1620 22430 1980 22470
rect 2020 22430 2380 22470
rect 2420 22430 2780 22470
rect 2820 22430 3180 22470
rect 3220 22430 3580 22470
rect 3620 22430 3980 22470
rect 4020 22430 4380 22470
rect 4420 22430 4780 22470
rect 4820 22430 5180 22470
rect 5220 22430 5580 22470
rect 5620 22430 5980 22470
rect 6020 22430 6380 22470
rect 6420 22430 6780 22470
rect 6820 22430 7180 22470
rect 7220 22430 7580 22470
rect 7620 22430 7980 22470
rect 8020 22430 8380 22470
rect 8420 22430 8780 22470
rect 8820 22430 9180 22470
rect 9220 22430 9580 22470
rect 9620 22430 9980 22470
rect 10020 22430 10380 22470
rect 10420 22430 10780 22470
rect 10820 22430 11180 22470
rect 11220 22430 11580 22470
rect 11620 22430 11980 22470
rect 12020 22430 12380 22470
rect 12420 22430 12780 22470
rect 12820 22430 13180 22470
rect 13220 22430 13580 22470
rect 13620 22430 13980 22470
rect 14020 22430 14380 22470
rect 14420 22430 14780 22470
rect 14820 22430 15180 22470
rect 15220 22430 15580 22470
rect 15620 22430 16000 22470
rect 0 22070 16000 22430
rect 0 22030 380 22070
rect 420 22030 780 22070
rect 820 22030 1180 22070
rect 1220 22030 1580 22070
rect 1620 22030 1980 22070
rect 2020 22030 2380 22070
rect 2420 22030 2780 22070
rect 2820 22030 3180 22070
rect 3220 22030 3580 22070
rect 3620 22030 3980 22070
rect 4020 22030 4380 22070
rect 4420 22030 4780 22070
rect 4820 22030 5180 22070
rect 5220 22030 5580 22070
rect 5620 22030 5980 22070
rect 6020 22030 6380 22070
rect 6420 22030 6780 22070
rect 6820 22030 7180 22070
rect 7220 22030 7580 22070
rect 7620 22030 7980 22070
rect 8020 22030 8380 22070
rect 8420 22030 8780 22070
rect 8820 22030 9180 22070
rect 9220 22030 9580 22070
rect 9620 22030 9980 22070
rect 10020 22030 10380 22070
rect 10420 22030 10780 22070
rect 10820 22030 11180 22070
rect 11220 22030 11580 22070
rect 11620 22030 11980 22070
rect 12020 22030 12380 22070
rect 12420 22030 12780 22070
rect 12820 22030 13180 22070
rect 13220 22030 13580 22070
rect 13620 22030 13980 22070
rect 14020 22030 14380 22070
rect 14420 22030 14780 22070
rect 14820 22030 15180 22070
rect 15220 22030 15580 22070
rect 15620 22030 16000 22070
rect 0 21670 16000 22030
rect 0 21630 380 21670
rect 420 21630 780 21670
rect 820 21630 1180 21670
rect 1220 21630 1580 21670
rect 1620 21630 1980 21670
rect 2020 21630 2380 21670
rect 2420 21630 2780 21670
rect 2820 21630 3180 21670
rect 3220 21630 3580 21670
rect 3620 21630 3980 21670
rect 4020 21630 4380 21670
rect 4420 21630 4780 21670
rect 4820 21630 5180 21670
rect 5220 21630 5580 21670
rect 5620 21630 5980 21670
rect 6020 21630 6380 21670
rect 6420 21630 6780 21670
rect 6820 21630 7180 21670
rect 7220 21630 7580 21670
rect 7620 21630 7980 21670
rect 8020 21630 8380 21670
rect 8420 21630 8780 21670
rect 8820 21630 9180 21670
rect 9220 21630 9580 21670
rect 9620 21630 9980 21670
rect 10020 21630 10380 21670
rect 10420 21630 10780 21670
rect 10820 21630 11180 21670
rect 11220 21630 11580 21670
rect 11620 21630 11980 21670
rect 12020 21630 12380 21670
rect 12420 21630 12780 21670
rect 12820 21630 13180 21670
rect 13220 21630 13580 21670
rect 13620 21630 13980 21670
rect 14020 21630 14380 21670
rect 14420 21630 14780 21670
rect 14820 21630 15180 21670
rect 15220 21630 15580 21670
rect 15620 21630 16000 21670
rect 0 21270 16000 21630
rect 0 21230 380 21270
rect 420 21230 780 21270
rect 820 21230 1180 21270
rect 1220 21230 1580 21270
rect 1620 21230 1980 21270
rect 2020 21230 2380 21270
rect 2420 21230 2780 21270
rect 2820 21230 3180 21270
rect 3220 21230 3580 21270
rect 3620 21230 3980 21270
rect 4020 21230 4380 21270
rect 4420 21230 4780 21270
rect 4820 21230 5180 21270
rect 5220 21230 5580 21270
rect 5620 21230 5980 21270
rect 6020 21230 6380 21270
rect 6420 21230 6780 21270
rect 6820 21230 7180 21270
rect 7220 21230 7580 21270
rect 7620 21230 7980 21270
rect 8020 21230 8380 21270
rect 8420 21230 8780 21270
rect 8820 21230 9180 21270
rect 9220 21230 9580 21270
rect 9620 21230 9980 21270
rect 10020 21230 10380 21270
rect 10420 21230 10780 21270
rect 10820 21230 11180 21270
rect 11220 21230 11580 21270
rect 11620 21230 11980 21270
rect 12020 21230 12380 21270
rect 12420 21230 12780 21270
rect 12820 21230 13180 21270
rect 13220 21230 13580 21270
rect 13620 21230 13980 21270
rect 14020 21230 14380 21270
rect 14420 21230 14780 21270
rect 14820 21230 15180 21270
rect 15220 21230 15580 21270
rect 15620 21230 16000 21270
rect 0 20870 16000 21230
rect 0 20830 380 20870
rect 420 20830 780 20870
rect 820 20830 1180 20870
rect 1220 20830 1580 20870
rect 1620 20830 1980 20870
rect 2020 20830 2380 20870
rect 2420 20830 2780 20870
rect 2820 20830 3180 20870
rect 3220 20830 3580 20870
rect 3620 20830 3980 20870
rect 4020 20830 4380 20870
rect 4420 20830 4780 20870
rect 4820 20830 5180 20870
rect 5220 20830 5580 20870
rect 5620 20830 5980 20870
rect 6020 20830 6380 20870
rect 6420 20830 6780 20870
rect 6820 20830 7180 20870
rect 7220 20830 7580 20870
rect 7620 20830 7980 20870
rect 8020 20830 8380 20870
rect 8420 20830 8780 20870
rect 8820 20830 9180 20870
rect 9220 20830 9580 20870
rect 9620 20830 9980 20870
rect 10020 20830 10380 20870
rect 10420 20830 10780 20870
rect 10820 20830 11180 20870
rect 11220 20830 11580 20870
rect 11620 20830 11980 20870
rect 12020 20830 12380 20870
rect 12420 20830 12780 20870
rect 12820 20830 13180 20870
rect 13220 20830 13580 20870
rect 13620 20830 13980 20870
rect 14020 20830 14380 20870
rect 14420 20830 14780 20870
rect 14820 20830 15180 20870
rect 15220 20830 15580 20870
rect 15620 20830 16000 20870
rect 0 20470 16000 20830
rect 0 20430 380 20470
rect 420 20430 780 20470
rect 820 20430 1180 20470
rect 1220 20430 1580 20470
rect 1620 20430 1980 20470
rect 2020 20430 2380 20470
rect 2420 20430 2780 20470
rect 2820 20430 3180 20470
rect 3220 20430 3580 20470
rect 3620 20430 3980 20470
rect 4020 20430 4380 20470
rect 4420 20430 4780 20470
rect 4820 20430 5180 20470
rect 5220 20430 5580 20470
rect 5620 20430 5980 20470
rect 6020 20430 6380 20470
rect 6420 20430 6780 20470
rect 6820 20430 7180 20470
rect 7220 20430 7580 20470
rect 7620 20430 7980 20470
rect 8020 20430 8380 20470
rect 8420 20430 8780 20470
rect 8820 20430 9180 20470
rect 9220 20430 9580 20470
rect 9620 20430 9980 20470
rect 10020 20430 10380 20470
rect 10420 20430 10780 20470
rect 10820 20430 11180 20470
rect 11220 20430 11580 20470
rect 11620 20430 11980 20470
rect 12020 20430 12380 20470
rect 12420 20430 12780 20470
rect 12820 20430 13180 20470
rect 13220 20430 13580 20470
rect 13620 20430 13980 20470
rect 14020 20430 14380 20470
rect 14420 20430 14780 20470
rect 14820 20430 15180 20470
rect 15220 20430 15580 20470
rect 15620 20430 16000 20470
rect 0 20070 16000 20430
rect 0 20030 380 20070
rect 420 20030 780 20070
rect 820 20030 1180 20070
rect 1220 20030 1580 20070
rect 1620 20030 1980 20070
rect 2020 20030 2380 20070
rect 2420 20030 2780 20070
rect 2820 20030 3180 20070
rect 3220 20030 3580 20070
rect 3620 20030 3980 20070
rect 4020 20030 4380 20070
rect 4420 20030 4780 20070
rect 4820 20030 5180 20070
rect 5220 20030 5580 20070
rect 5620 20030 5980 20070
rect 6020 20030 6380 20070
rect 6420 20030 6780 20070
rect 6820 20030 7180 20070
rect 7220 20030 7580 20070
rect 7620 20030 7980 20070
rect 8020 20030 8380 20070
rect 8420 20030 8780 20070
rect 8820 20030 9180 20070
rect 9220 20030 9580 20070
rect 9620 20030 9980 20070
rect 10020 20030 10380 20070
rect 10420 20030 10780 20070
rect 10820 20030 11180 20070
rect 11220 20030 11580 20070
rect 11620 20030 11980 20070
rect 12020 20030 12380 20070
rect 12420 20030 12780 20070
rect 12820 20030 13180 20070
rect 13220 20030 13580 20070
rect 13620 20030 13980 20070
rect 14020 20030 14380 20070
rect 14420 20030 14780 20070
rect 14820 20030 15180 20070
rect 15220 20030 15580 20070
rect 15620 20030 16000 20070
rect 0 19670 16000 20030
rect 0 19630 380 19670
rect 420 19630 780 19670
rect 820 19630 1180 19670
rect 1220 19630 1580 19670
rect 1620 19630 1980 19670
rect 2020 19630 2380 19670
rect 2420 19630 2780 19670
rect 2820 19630 3180 19670
rect 3220 19630 3580 19670
rect 3620 19630 3980 19670
rect 4020 19630 4380 19670
rect 4420 19630 4780 19670
rect 4820 19630 5180 19670
rect 5220 19630 5580 19670
rect 5620 19630 5980 19670
rect 6020 19630 6380 19670
rect 6420 19630 6780 19670
rect 6820 19630 7180 19670
rect 7220 19630 7580 19670
rect 7620 19630 7980 19670
rect 8020 19630 8380 19670
rect 8420 19630 8780 19670
rect 8820 19630 9180 19670
rect 9220 19630 9580 19670
rect 9620 19630 9980 19670
rect 10020 19630 10380 19670
rect 10420 19630 10780 19670
rect 10820 19630 11180 19670
rect 11220 19630 11580 19670
rect 11620 19630 11980 19670
rect 12020 19630 12380 19670
rect 12420 19630 12780 19670
rect 12820 19630 13180 19670
rect 13220 19630 13580 19670
rect 13620 19630 13980 19670
rect 14020 19630 14380 19670
rect 14420 19630 14780 19670
rect 14820 19630 15180 19670
rect 15220 19630 15580 19670
rect 15620 19630 16000 19670
rect 0 19270 16000 19630
rect 0 19230 380 19270
rect 420 19230 780 19270
rect 820 19230 1180 19270
rect 1220 19230 1580 19270
rect 1620 19230 1980 19270
rect 2020 19230 2380 19270
rect 2420 19230 2780 19270
rect 2820 19230 3180 19270
rect 3220 19230 3580 19270
rect 3620 19230 3980 19270
rect 4020 19230 4380 19270
rect 4420 19230 4780 19270
rect 4820 19230 5180 19270
rect 5220 19230 5580 19270
rect 5620 19230 5980 19270
rect 6020 19230 6380 19270
rect 6420 19230 6780 19270
rect 6820 19230 7180 19270
rect 7220 19230 7580 19270
rect 7620 19230 7980 19270
rect 8020 19230 8380 19270
rect 8420 19230 8780 19270
rect 8820 19230 9180 19270
rect 9220 19230 9580 19270
rect 9620 19230 9980 19270
rect 10020 19230 10380 19270
rect 10420 19230 10780 19270
rect 10820 19230 11180 19270
rect 11220 19230 11580 19270
rect 11620 19230 11980 19270
rect 12020 19230 12380 19270
rect 12420 19230 12780 19270
rect 12820 19230 13180 19270
rect 13220 19230 13580 19270
rect 13620 19230 13980 19270
rect 14020 19230 14380 19270
rect 14420 19230 14780 19270
rect 14820 19230 15180 19270
rect 15220 19230 15580 19270
rect 15620 19230 16000 19270
rect 0 18700 16000 19230
rect 0 17770 16000 18300
rect 0 17730 380 17770
rect 420 17730 780 17770
rect 820 17730 1180 17770
rect 1220 17730 1580 17770
rect 1620 17730 1980 17770
rect 2020 17730 2380 17770
rect 2420 17730 2780 17770
rect 2820 17730 3180 17770
rect 3220 17730 3580 17770
rect 3620 17730 3980 17770
rect 4020 17730 4380 17770
rect 4420 17730 4780 17770
rect 4820 17730 5180 17770
rect 5220 17730 5580 17770
rect 5620 17730 5980 17770
rect 6020 17730 6380 17770
rect 6420 17730 6780 17770
rect 6820 17730 7180 17770
rect 7220 17730 7580 17770
rect 7620 17730 7980 17770
rect 8020 17730 8380 17770
rect 8420 17730 8780 17770
rect 8820 17730 9180 17770
rect 9220 17730 9580 17770
rect 9620 17730 9980 17770
rect 10020 17730 10380 17770
rect 10420 17730 10780 17770
rect 10820 17730 11180 17770
rect 11220 17730 11580 17770
rect 11620 17730 11980 17770
rect 12020 17730 12380 17770
rect 12420 17730 12780 17770
rect 12820 17730 13180 17770
rect 13220 17730 13580 17770
rect 13620 17730 13980 17770
rect 14020 17730 14380 17770
rect 14420 17730 14780 17770
rect 14820 17730 15180 17770
rect 15220 17730 15580 17770
rect 15620 17730 16000 17770
rect 0 17370 16000 17730
rect 0 17330 380 17370
rect 420 17330 780 17370
rect 820 17330 1180 17370
rect 1220 17330 1580 17370
rect 1620 17330 1980 17370
rect 2020 17330 2380 17370
rect 2420 17330 2780 17370
rect 2820 17330 3180 17370
rect 3220 17330 3580 17370
rect 3620 17330 3980 17370
rect 4020 17330 4380 17370
rect 4420 17330 4780 17370
rect 4820 17330 5180 17370
rect 5220 17330 5580 17370
rect 5620 17330 5980 17370
rect 6020 17330 6380 17370
rect 6420 17330 6780 17370
rect 6820 17330 7180 17370
rect 7220 17330 7580 17370
rect 7620 17330 7980 17370
rect 8020 17330 8380 17370
rect 8420 17330 8780 17370
rect 8820 17330 9180 17370
rect 9220 17330 9580 17370
rect 9620 17330 9980 17370
rect 10020 17330 10380 17370
rect 10420 17330 10780 17370
rect 10820 17330 11180 17370
rect 11220 17330 11580 17370
rect 11620 17330 11980 17370
rect 12020 17330 12380 17370
rect 12420 17330 12780 17370
rect 12820 17330 13180 17370
rect 13220 17330 13580 17370
rect 13620 17330 13980 17370
rect 14020 17330 14380 17370
rect 14420 17330 14780 17370
rect 14820 17330 15180 17370
rect 15220 17330 15580 17370
rect 15620 17330 16000 17370
rect 0 16970 16000 17330
rect 0 16930 380 16970
rect 420 16930 780 16970
rect 820 16930 1180 16970
rect 1220 16930 1580 16970
rect 1620 16930 1980 16970
rect 2020 16930 2380 16970
rect 2420 16930 2780 16970
rect 2820 16930 3180 16970
rect 3220 16930 3580 16970
rect 3620 16930 3980 16970
rect 4020 16930 4380 16970
rect 4420 16930 4780 16970
rect 4820 16930 5180 16970
rect 5220 16930 5580 16970
rect 5620 16930 5980 16970
rect 6020 16930 6380 16970
rect 6420 16930 6780 16970
rect 6820 16930 7180 16970
rect 7220 16930 7580 16970
rect 7620 16930 7980 16970
rect 8020 16930 8380 16970
rect 8420 16930 8780 16970
rect 8820 16930 9180 16970
rect 9220 16930 9580 16970
rect 9620 16930 9980 16970
rect 10020 16930 10380 16970
rect 10420 16930 10780 16970
rect 10820 16930 11180 16970
rect 11220 16930 11580 16970
rect 11620 16930 11980 16970
rect 12020 16930 12380 16970
rect 12420 16930 12780 16970
rect 12820 16930 13180 16970
rect 13220 16930 13580 16970
rect 13620 16930 13980 16970
rect 14020 16930 14380 16970
rect 14420 16930 14780 16970
rect 14820 16930 15180 16970
rect 15220 16930 15580 16970
rect 15620 16930 16000 16970
rect 0 16570 16000 16930
rect 0 16530 380 16570
rect 420 16530 780 16570
rect 820 16530 1180 16570
rect 1220 16530 1580 16570
rect 1620 16530 1980 16570
rect 2020 16530 2380 16570
rect 2420 16530 2780 16570
rect 2820 16530 3180 16570
rect 3220 16530 3580 16570
rect 3620 16530 3980 16570
rect 4020 16530 4380 16570
rect 4420 16530 4780 16570
rect 4820 16530 5180 16570
rect 5220 16530 5580 16570
rect 5620 16530 5980 16570
rect 6020 16530 6380 16570
rect 6420 16530 6780 16570
rect 6820 16530 7180 16570
rect 7220 16530 7580 16570
rect 7620 16530 7980 16570
rect 8020 16530 8380 16570
rect 8420 16530 8780 16570
rect 8820 16530 9180 16570
rect 9220 16530 9580 16570
rect 9620 16530 9980 16570
rect 10020 16530 10380 16570
rect 10420 16530 10780 16570
rect 10820 16530 11180 16570
rect 11220 16530 11580 16570
rect 11620 16530 11980 16570
rect 12020 16530 12380 16570
rect 12420 16530 12780 16570
rect 12820 16530 13180 16570
rect 13220 16530 13580 16570
rect 13620 16530 13980 16570
rect 14020 16530 14380 16570
rect 14420 16530 14780 16570
rect 14820 16530 15180 16570
rect 15220 16530 15580 16570
rect 15620 16530 16000 16570
rect 0 16170 16000 16530
rect 0 16130 380 16170
rect 420 16130 780 16170
rect 820 16130 1180 16170
rect 1220 16130 1580 16170
rect 1620 16130 1980 16170
rect 2020 16130 2380 16170
rect 2420 16130 2780 16170
rect 2820 16130 3180 16170
rect 3220 16130 3580 16170
rect 3620 16130 3980 16170
rect 4020 16130 4380 16170
rect 4420 16130 4780 16170
rect 4820 16130 5180 16170
rect 5220 16130 5580 16170
rect 5620 16130 5980 16170
rect 6020 16130 6380 16170
rect 6420 16130 6780 16170
rect 6820 16130 7180 16170
rect 7220 16130 7580 16170
rect 7620 16130 7980 16170
rect 8020 16130 8380 16170
rect 8420 16130 8780 16170
rect 8820 16130 9180 16170
rect 9220 16130 9580 16170
rect 9620 16130 9980 16170
rect 10020 16130 10380 16170
rect 10420 16130 10780 16170
rect 10820 16130 11180 16170
rect 11220 16130 11580 16170
rect 11620 16130 11980 16170
rect 12020 16130 12380 16170
rect 12420 16130 12780 16170
rect 12820 16130 13180 16170
rect 13220 16130 13580 16170
rect 13620 16130 13980 16170
rect 14020 16130 14380 16170
rect 14420 16130 14780 16170
rect 14820 16130 15180 16170
rect 15220 16130 15580 16170
rect 15620 16130 16000 16170
rect 0 15770 16000 16130
rect 0 15730 380 15770
rect 420 15730 780 15770
rect 820 15730 1180 15770
rect 1220 15730 1580 15770
rect 1620 15730 1980 15770
rect 2020 15730 2380 15770
rect 2420 15730 2780 15770
rect 2820 15730 3180 15770
rect 3220 15730 3580 15770
rect 3620 15730 3980 15770
rect 4020 15730 4380 15770
rect 4420 15730 4780 15770
rect 4820 15730 5180 15770
rect 5220 15730 5580 15770
rect 5620 15730 5980 15770
rect 6020 15730 6380 15770
rect 6420 15730 6780 15770
rect 6820 15730 7180 15770
rect 7220 15730 7580 15770
rect 7620 15730 7980 15770
rect 8020 15730 8380 15770
rect 8420 15730 8780 15770
rect 8820 15730 9180 15770
rect 9220 15730 9580 15770
rect 9620 15730 9980 15770
rect 10020 15730 10380 15770
rect 10420 15730 10780 15770
rect 10820 15730 11180 15770
rect 11220 15730 11580 15770
rect 11620 15730 11980 15770
rect 12020 15730 12380 15770
rect 12420 15730 12780 15770
rect 12820 15730 13180 15770
rect 13220 15730 13580 15770
rect 13620 15730 13980 15770
rect 14020 15730 14380 15770
rect 14420 15730 14780 15770
rect 14820 15730 15180 15770
rect 15220 15730 15580 15770
rect 15620 15730 16000 15770
rect 0 15370 16000 15730
rect 0 15330 380 15370
rect 420 15330 780 15370
rect 820 15330 1180 15370
rect 1220 15330 1580 15370
rect 1620 15330 1980 15370
rect 2020 15330 2380 15370
rect 2420 15330 2780 15370
rect 2820 15330 3180 15370
rect 3220 15330 3580 15370
rect 3620 15330 3980 15370
rect 4020 15330 4380 15370
rect 4420 15330 4780 15370
rect 4820 15330 5180 15370
rect 5220 15330 5580 15370
rect 5620 15330 5980 15370
rect 6020 15330 6380 15370
rect 6420 15330 6780 15370
rect 6820 15330 7180 15370
rect 7220 15330 7580 15370
rect 7620 15330 7980 15370
rect 8020 15330 8380 15370
rect 8420 15330 8780 15370
rect 8820 15330 9180 15370
rect 9220 15330 9580 15370
rect 9620 15330 9980 15370
rect 10020 15330 10380 15370
rect 10420 15330 10780 15370
rect 10820 15330 11180 15370
rect 11220 15330 11580 15370
rect 11620 15330 11980 15370
rect 12020 15330 12380 15370
rect 12420 15330 12780 15370
rect 12820 15330 13180 15370
rect 13220 15330 13580 15370
rect 13620 15330 13980 15370
rect 14020 15330 14380 15370
rect 14420 15330 14780 15370
rect 14820 15330 15180 15370
rect 15220 15330 15580 15370
rect 15620 15330 16000 15370
rect 0 14970 16000 15330
rect 0 14930 380 14970
rect 420 14930 780 14970
rect 820 14930 1180 14970
rect 1220 14930 1580 14970
rect 1620 14930 1980 14970
rect 2020 14930 2380 14970
rect 2420 14930 2780 14970
rect 2820 14930 3180 14970
rect 3220 14930 3580 14970
rect 3620 14930 3980 14970
rect 4020 14930 4380 14970
rect 4420 14930 4780 14970
rect 4820 14930 5180 14970
rect 5220 14930 5580 14970
rect 5620 14930 5980 14970
rect 6020 14930 6380 14970
rect 6420 14930 6780 14970
rect 6820 14930 7180 14970
rect 7220 14930 7580 14970
rect 7620 14930 7980 14970
rect 8020 14930 8380 14970
rect 8420 14930 8780 14970
rect 8820 14930 9180 14970
rect 9220 14930 9580 14970
rect 9620 14930 9980 14970
rect 10020 14930 10380 14970
rect 10420 14930 10780 14970
rect 10820 14930 11180 14970
rect 11220 14930 11580 14970
rect 11620 14930 11980 14970
rect 12020 14930 12380 14970
rect 12420 14930 12780 14970
rect 12820 14930 13180 14970
rect 13220 14930 13580 14970
rect 13620 14930 13980 14970
rect 14020 14930 14380 14970
rect 14420 14930 14780 14970
rect 14820 14930 15180 14970
rect 15220 14930 15580 14970
rect 15620 14930 16000 14970
rect 0 14570 16000 14930
rect 0 14530 380 14570
rect 420 14530 780 14570
rect 820 14530 1180 14570
rect 1220 14530 1580 14570
rect 1620 14530 1980 14570
rect 2020 14530 2380 14570
rect 2420 14530 2780 14570
rect 2820 14530 3180 14570
rect 3220 14530 3580 14570
rect 3620 14530 3980 14570
rect 4020 14530 4380 14570
rect 4420 14530 4780 14570
rect 4820 14530 5180 14570
rect 5220 14530 5580 14570
rect 5620 14530 5980 14570
rect 6020 14530 6380 14570
rect 6420 14530 6780 14570
rect 6820 14530 7180 14570
rect 7220 14530 7580 14570
rect 7620 14530 7980 14570
rect 8020 14530 8380 14570
rect 8420 14530 8780 14570
rect 8820 14530 9180 14570
rect 9220 14530 9580 14570
rect 9620 14530 9980 14570
rect 10020 14530 10380 14570
rect 10420 14530 10780 14570
rect 10820 14530 11180 14570
rect 11220 14530 11580 14570
rect 11620 14530 11980 14570
rect 12020 14530 12380 14570
rect 12420 14530 12780 14570
rect 12820 14530 13180 14570
rect 13220 14530 13580 14570
rect 13620 14530 13980 14570
rect 14020 14530 14380 14570
rect 14420 14530 14780 14570
rect 14820 14530 15180 14570
rect 15220 14530 15580 14570
rect 15620 14530 16000 14570
rect 0 14170 16000 14530
rect 0 14130 380 14170
rect 420 14130 780 14170
rect 820 14130 1180 14170
rect 1220 14130 1580 14170
rect 1620 14130 1980 14170
rect 2020 14130 2380 14170
rect 2420 14130 2780 14170
rect 2820 14130 3180 14170
rect 3220 14130 3580 14170
rect 3620 14130 3980 14170
rect 4020 14130 4380 14170
rect 4420 14130 4780 14170
rect 4820 14130 5180 14170
rect 5220 14130 5580 14170
rect 5620 14130 5980 14170
rect 6020 14130 6380 14170
rect 6420 14130 6780 14170
rect 6820 14130 7180 14170
rect 7220 14130 7580 14170
rect 7620 14130 7980 14170
rect 8020 14130 8380 14170
rect 8420 14130 8780 14170
rect 8820 14130 9180 14170
rect 9220 14130 9580 14170
rect 9620 14130 9980 14170
rect 10020 14130 10380 14170
rect 10420 14130 10780 14170
rect 10820 14130 11180 14170
rect 11220 14130 11580 14170
rect 11620 14130 11980 14170
rect 12020 14130 12380 14170
rect 12420 14130 12780 14170
rect 12820 14130 13180 14170
rect 13220 14130 13580 14170
rect 13620 14130 13980 14170
rect 14020 14130 14380 14170
rect 14420 14130 14780 14170
rect 14820 14130 15180 14170
rect 15220 14130 15580 14170
rect 15620 14130 16000 14170
rect 0 13770 16000 14130
rect 0 13730 380 13770
rect 420 13730 780 13770
rect 820 13730 1180 13770
rect 1220 13730 1580 13770
rect 1620 13730 1980 13770
rect 2020 13730 2380 13770
rect 2420 13730 2780 13770
rect 2820 13730 3180 13770
rect 3220 13730 3580 13770
rect 3620 13730 3980 13770
rect 4020 13730 4380 13770
rect 4420 13730 4780 13770
rect 4820 13730 5180 13770
rect 5220 13730 5580 13770
rect 5620 13730 5980 13770
rect 6020 13730 6380 13770
rect 6420 13730 6780 13770
rect 6820 13730 7180 13770
rect 7220 13730 7580 13770
rect 7620 13730 7980 13770
rect 8020 13730 8380 13770
rect 8420 13730 8780 13770
rect 8820 13730 9180 13770
rect 9220 13730 9580 13770
rect 9620 13730 9980 13770
rect 10020 13730 10380 13770
rect 10420 13730 10780 13770
rect 10820 13730 11180 13770
rect 11220 13730 11580 13770
rect 11620 13730 11980 13770
rect 12020 13730 12380 13770
rect 12420 13730 12780 13770
rect 12820 13730 13180 13770
rect 13220 13730 13580 13770
rect 13620 13730 13980 13770
rect 14020 13730 14380 13770
rect 14420 13730 14780 13770
rect 14820 13730 15180 13770
rect 15220 13730 15580 13770
rect 15620 13730 16000 13770
rect 0 13200 16000 13730
rect 0 11470 16000 12000
rect 0 11430 380 11470
rect 420 11430 780 11470
rect 820 11430 1180 11470
rect 1220 11430 1580 11470
rect 1620 11430 1980 11470
rect 2020 11430 2380 11470
rect 2420 11430 2780 11470
rect 2820 11430 3180 11470
rect 3220 11430 3580 11470
rect 3620 11430 3980 11470
rect 4020 11430 4380 11470
rect 4420 11430 4780 11470
rect 4820 11430 5180 11470
rect 5220 11430 5580 11470
rect 5620 11430 5980 11470
rect 6020 11430 6380 11470
rect 6420 11430 6780 11470
rect 6820 11430 7180 11470
rect 7220 11430 7580 11470
rect 7620 11430 7980 11470
rect 8020 11430 8380 11470
rect 8420 11430 8780 11470
rect 8820 11430 9180 11470
rect 9220 11430 9580 11470
rect 9620 11430 9980 11470
rect 10020 11430 10380 11470
rect 10420 11430 10780 11470
rect 10820 11430 11180 11470
rect 11220 11430 11580 11470
rect 11620 11430 11980 11470
rect 12020 11430 12380 11470
rect 12420 11430 12780 11470
rect 12820 11430 13180 11470
rect 13220 11430 13580 11470
rect 13620 11430 13980 11470
rect 14020 11430 14380 11470
rect 14420 11430 14780 11470
rect 14820 11430 15180 11470
rect 15220 11430 15580 11470
rect 15620 11430 16000 11470
rect 0 11070 16000 11430
rect 0 11030 380 11070
rect 420 11030 780 11070
rect 820 11030 1180 11070
rect 1220 11030 1580 11070
rect 1620 11030 1980 11070
rect 2020 11030 2380 11070
rect 2420 11030 2780 11070
rect 2820 11030 3180 11070
rect 3220 11030 3580 11070
rect 3620 11030 3980 11070
rect 4020 11030 4380 11070
rect 4420 11030 4780 11070
rect 4820 11030 5180 11070
rect 5220 11030 5580 11070
rect 5620 11030 5980 11070
rect 6020 11030 6380 11070
rect 6420 11030 6780 11070
rect 6820 11030 7180 11070
rect 7220 11030 7580 11070
rect 7620 11030 7980 11070
rect 8020 11030 8380 11070
rect 8420 11030 8780 11070
rect 8820 11030 9180 11070
rect 9220 11030 9580 11070
rect 9620 11030 9980 11070
rect 10020 11030 10380 11070
rect 10420 11030 10780 11070
rect 10820 11030 11180 11070
rect 11220 11030 11580 11070
rect 11620 11030 11980 11070
rect 12020 11030 12380 11070
rect 12420 11030 12780 11070
rect 12820 11030 13180 11070
rect 13220 11030 13580 11070
rect 13620 11030 13980 11070
rect 14020 11030 14380 11070
rect 14420 11030 14780 11070
rect 14820 11030 15180 11070
rect 15220 11030 15580 11070
rect 15620 11030 16000 11070
rect 0 10670 16000 11030
rect 0 10630 380 10670
rect 420 10630 780 10670
rect 820 10630 1180 10670
rect 1220 10630 1580 10670
rect 1620 10630 1980 10670
rect 2020 10630 2380 10670
rect 2420 10630 2780 10670
rect 2820 10630 3180 10670
rect 3220 10630 3580 10670
rect 3620 10630 3980 10670
rect 4020 10630 4380 10670
rect 4420 10630 4780 10670
rect 4820 10630 5180 10670
rect 5220 10630 5580 10670
rect 5620 10630 5980 10670
rect 6020 10630 6380 10670
rect 6420 10630 6780 10670
rect 6820 10630 7180 10670
rect 7220 10630 7580 10670
rect 7620 10630 7980 10670
rect 8020 10630 8380 10670
rect 8420 10630 8780 10670
rect 8820 10630 9180 10670
rect 9220 10630 9580 10670
rect 9620 10630 9980 10670
rect 10020 10630 10380 10670
rect 10420 10630 10780 10670
rect 10820 10630 11180 10670
rect 11220 10630 11580 10670
rect 11620 10630 11980 10670
rect 12020 10630 12380 10670
rect 12420 10630 12780 10670
rect 12820 10630 13180 10670
rect 13220 10630 13580 10670
rect 13620 10630 13980 10670
rect 14020 10630 14380 10670
rect 14420 10630 14780 10670
rect 14820 10630 15180 10670
rect 15220 10630 15580 10670
rect 15620 10630 16000 10670
rect 0 10270 16000 10630
rect 0 10230 380 10270
rect 420 10230 780 10270
rect 820 10230 1180 10270
rect 1220 10230 1580 10270
rect 1620 10230 1980 10270
rect 2020 10230 2380 10270
rect 2420 10230 2780 10270
rect 2820 10230 3180 10270
rect 3220 10230 3580 10270
rect 3620 10230 3980 10270
rect 4020 10230 4380 10270
rect 4420 10230 4780 10270
rect 4820 10230 5180 10270
rect 5220 10230 5580 10270
rect 5620 10230 5980 10270
rect 6020 10230 6380 10270
rect 6420 10230 6780 10270
rect 6820 10230 7180 10270
rect 7220 10230 7580 10270
rect 7620 10230 7980 10270
rect 8020 10230 8380 10270
rect 8420 10230 8780 10270
rect 8820 10230 9180 10270
rect 9220 10230 9580 10270
rect 9620 10230 9980 10270
rect 10020 10230 10380 10270
rect 10420 10230 10780 10270
rect 10820 10230 11180 10270
rect 11220 10230 11580 10270
rect 11620 10230 11980 10270
rect 12020 10230 12380 10270
rect 12420 10230 12780 10270
rect 12820 10230 13180 10270
rect 13220 10230 13580 10270
rect 13620 10230 13980 10270
rect 14020 10230 14380 10270
rect 14420 10230 14780 10270
rect 14820 10230 15180 10270
rect 15220 10230 15580 10270
rect 15620 10230 16000 10270
rect 0 9870 16000 10230
rect 0 9830 380 9870
rect 420 9830 780 9870
rect 820 9830 1180 9870
rect 1220 9830 1580 9870
rect 1620 9830 1980 9870
rect 2020 9830 2380 9870
rect 2420 9830 2780 9870
rect 2820 9830 3180 9870
rect 3220 9830 3580 9870
rect 3620 9830 3980 9870
rect 4020 9830 4380 9870
rect 4420 9830 4780 9870
rect 4820 9830 5180 9870
rect 5220 9830 5580 9870
rect 5620 9830 5980 9870
rect 6020 9830 6380 9870
rect 6420 9830 6780 9870
rect 6820 9830 7180 9870
rect 7220 9830 7580 9870
rect 7620 9830 7980 9870
rect 8020 9830 8380 9870
rect 8420 9830 8780 9870
rect 8820 9830 9180 9870
rect 9220 9830 9580 9870
rect 9620 9830 9980 9870
rect 10020 9830 10380 9870
rect 10420 9830 10780 9870
rect 10820 9830 11180 9870
rect 11220 9830 11580 9870
rect 11620 9830 11980 9870
rect 12020 9830 12380 9870
rect 12420 9830 12780 9870
rect 12820 9830 13180 9870
rect 13220 9830 13580 9870
rect 13620 9830 13980 9870
rect 14020 9830 14380 9870
rect 14420 9830 14780 9870
rect 14820 9830 15180 9870
rect 15220 9830 15580 9870
rect 15620 9830 16000 9870
rect 0 9470 16000 9830
rect 0 9430 380 9470
rect 420 9430 780 9470
rect 820 9430 1180 9470
rect 1220 9430 1580 9470
rect 1620 9430 1980 9470
rect 2020 9430 2380 9470
rect 2420 9430 2780 9470
rect 2820 9430 3180 9470
rect 3220 9430 3580 9470
rect 3620 9430 3980 9470
rect 4020 9430 4380 9470
rect 4420 9430 4780 9470
rect 4820 9430 5180 9470
rect 5220 9430 5580 9470
rect 5620 9430 5980 9470
rect 6020 9430 6380 9470
rect 6420 9430 6780 9470
rect 6820 9430 7180 9470
rect 7220 9430 7580 9470
rect 7620 9430 7980 9470
rect 8020 9430 8380 9470
rect 8420 9430 8780 9470
rect 8820 9430 9180 9470
rect 9220 9430 9580 9470
rect 9620 9430 9980 9470
rect 10020 9430 10380 9470
rect 10420 9430 10780 9470
rect 10820 9430 11180 9470
rect 11220 9430 11580 9470
rect 11620 9430 11980 9470
rect 12020 9430 12380 9470
rect 12420 9430 12780 9470
rect 12820 9430 13180 9470
rect 13220 9430 13580 9470
rect 13620 9430 13980 9470
rect 14020 9430 14380 9470
rect 14420 9430 14780 9470
rect 14820 9430 15180 9470
rect 15220 9430 15580 9470
rect 15620 9430 16000 9470
rect 0 9070 16000 9430
rect 0 9030 380 9070
rect 420 9030 780 9070
rect 820 9030 1180 9070
rect 1220 9030 1580 9070
rect 1620 9030 1980 9070
rect 2020 9030 2380 9070
rect 2420 9030 2780 9070
rect 2820 9030 3180 9070
rect 3220 9030 3580 9070
rect 3620 9030 3980 9070
rect 4020 9030 4380 9070
rect 4420 9030 4780 9070
rect 4820 9030 5180 9070
rect 5220 9030 5580 9070
rect 5620 9030 5980 9070
rect 6020 9030 6380 9070
rect 6420 9030 6780 9070
rect 6820 9030 7180 9070
rect 7220 9030 7580 9070
rect 7620 9030 7980 9070
rect 8020 9030 8380 9070
rect 8420 9030 8780 9070
rect 8820 9030 9180 9070
rect 9220 9030 9580 9070
rect 9620 9030 9980 9070
rect 10020 9030 10380 9070
rect 10420 9030 10780 9070
rect 10820 9030 11180 9070
rect 11220 9030 11580 9070
rect 11620 9030 11980 9070
rect 12020 9030 12380 9070
rect 12420 9030 12780 9070
rect 12820 9030 13180 9070
rect 13220 9030 13580 9070
rect 13620 9030 13980 9070
rect 14020 9030 14380 9070
rect 14420 9030 14780 9070
rect 14820 9030 15180 9070
rect 15220 9030 15580 9070
rect 15620 9030 16000 9070
rect 0 8670 16000 9030
rect 0 8630 380 8670
rect 420 8630 780 8670
rect 820 8630 1180 8670
rect 1220 8630 1580 8670
rect 1620 8630 1980 8670
rect 2020 8630 2380 8670
rect 2420 8630 2780 8670
rect 2820 8630 3180 8670
rect 3220 8630 3580 8670
rect 3620 8630 3980 8670
rect 4020 8630 4380 8670
rect 4420 8630 4780 8670
rect 4820 8630 5180 8670
rect 5220 8630 5580 8670
rect 5620 8630 5980 8670
rect 6020 8630 6380 8670
rect 6420 8630 6780 8670
rect 6820 8630 7180 8670
rect 7220 8630 7580 8670
rect 7620 8630 7980 8670
rect 8020 8630 8380 8670
rect 8420 8630 8780 8670
rect 8820 8630 9180 8670
rect 9220 8630 9580 8670
rect 9620 8630 9980 8670
rect 10020 8630 10380 8670
rect 10420 8630 10780 8670
rect 10820 8630 11180 8670
rect 11220 8630 11580 8670
rect 11620 8630 11980 8670
rect 12020 8630 12380 8670
rect 12420 8630 12780 8670
rect 12820 8630 13180 8670
rect 13220 8630 13580 8670
rect 13620 8630 13980 8670
rect 14020 8630 14380 8670
rect 14420 8630 14780 8670
rect 14820 8630 15180 8670
rect 15220 8630 15580 8670
rect 15620 8630 16000 8670
rect 0 8270 16000 8630
rect 0 8230 380 8270
rect 420 8230 780 8270
rect 820 8230 1180 8270
rect 1220 8230 1580 8270
rect 1620 8230 1980 8270
rect 2020 8230 2380 8270
rect 2420 8230 2780 8270
rect 2820 8230 3180 8270
rect 3220 8230 3580 8270
rect 3620 8230 3980 8270
rect 4020 8230 4380 8270
rect 4420 8230 4780 8270
rect 4820 8230 5180 8270
rect 5220 8230 5580 8270
rect 5620 8230 5980 8270
rect 6020 8230 6380 8270
rect 6420 8230 6780 8270
rect 6820 8230 7180 8270
rect 7220 8230 7580 8270
rect 7620 8230 7980 8270
rect 8020 8230 8380 8270
rect 8420 8230 8780 8270
rect 8820 8230 9180 8270
rect 9220 8230 9580 8270
rect 9620 8230 9980 8270
rect 10020 8230 10380 8270
rect 10420 8230 10780 8270
rect 10820 8230 11180 8270
rect 11220 8230 11580 8270
rect 11620 8230 11980 8270
rect 12020 8230 12380 8270
rect 12420 8230 12780 8270
rect 12820 8230 13180 8270
rect 13220 8230 13580 8270
rect 13620 8230 13980 8270
rect 14020 8230 14380 8270
rect 14420 8230 14780 8270
rect 14820 8230 15180 8270
rect 15220 8230 15580 8270
rect 15620 8230 16000 8270
rect 0 7870 16000 8230
rect 0 7830 380 7870
rect 420 7830 780 7870
rect 820 7830 1180 7870
rect 1220 7830 1580 7870
rect 1620 7830 1980 7870
rect 2020 7830 2380 7870
rect 2420 7830 2780 7870
rect 2820 7830 3180 7870
rect 3220 7830 3580 7870
rect 3620 7830 3980 7870
rect 4020 7830 4380 7870
rect 4420 7830 4780 7870
rect 4820 7830 5180 7870
rect 5220 7830 5580 7870
rect 5620 7830 5980 7870
rect 6020 7830 6380 7870
rect 6420 7830 6780 7870
rect 6820 7830 7180 7870
rect 7220 7830 7580 7870
rect 7620 7830 7980 7870
rect 8020 7830 8380 7870
rect 8420 7830 8780 7870
rect 8820 7830 9180 7870
rect 9220 7830 9580 7870
rect 9620 7830 9980 7870
rect 10020 7830 10380 7870
rect 10420 7830 10780 7870
rect 10820 7830 11180 7870
rect 11220 7830 11580 7870
rect 11620 7830 11980 7870
rect 12020 7830 12380 7870
rect 12420 7830 12780 7870
rect 12820 7830 13180 7870
rect 13220 7830 13580 7870
rect 13620 7830 13980 7870
rect 14020 7830 14380 7870
rect 14420 7830 14780 7870
rect 14820 7830 15180 7870
rect 15220 7830 15580 7870
rect 15620 7830 16000 7870
rect 0 7470 16000 7830
rect 0 7430 380 7470
rect 420 7430 780 7470
rect 820 7430 1180 7470
rect 1220 7430 1580 7470
rect 1620 7430 1980 7470
rect 2020 7430 2380 7470
rect 2420 7430 2780 7470
rect 2820 7430 3180 7470
rect 3220 7430 3580 7470
rect 3620 7430 3980 7470
rect 4020 7430 4380 7470
rect 4420 7430 4780 7470
rect 4820 7430 5180 7470
rect 5220 7430 5580 7470
rect 5620 7430 5980 7470
rect 6020 7430 6380 7470
rect 6420 7430 6780 7470
rect 6820 7430 7180 7470
rect 7220 7430 7580 7470
rect 7620 7430 7980 7470
rect 8020 7430 8380 7470
rect 8420 7430 8780 7470
rect 8820 7430 9180 7470
rect 9220 7430 9580 7470
rect 9620 7430 9980 7470
rect 10020 7430 10380 7470
rect 10420 7430 10780 7470
rect 10820 7430 11180 7470
rect 11220 7430 11580 7470
rect 11620 7430 11980 7470
rect 12020 7430 12380 7470
rect 12420 7430 12780 7470
rect 12820 7430 13180 7470
rect 13220 7430 13580 7470
rect 13620 7430 13980 7470
rect 14020 7430 14380 7470
rect 14420 7430 14780 7470
rect 14820 7430 15180 7470
rect 15220 7430 15580 7470
rect 15620 7430 16000 7470
rect 0 6900 16000 7430
rect 0 5970 16000 6500
rect 0 5930 380 5970
rect 420 5930 780 5970
rect 820 5930 1180 5970
rect 1220 5930 1580 5970
rect 1620 5930 1980 5970
rect 2020 5930 2380 5970
rect 2420 5930 2780 5970
rect 2820 5930 3180 5970
rect 3220 5930 3580 5970
rect 3620 5930 3980 5970
rect 4020 5930 4380 5970
rect 4420 5930 4780 5970
rect 4820 5930 5180 5970
rect 5220 5930 5580 5970
rect 5620 5930 5980 5970
rect 6020 5930 6380 5970
rect 6420 5930 6780 5970
rect 6820 5930 7180 5970
rect 7220 5930 7580 5970
rect 7620 5930 7980 5970
rect 8020 5930 8380 5970
rect 8420 5930 8780 5970
rect 8820 5930 9180 5970
rect 9220 5930 9580 5970
rect 9620 5930 9980 5970
rect 10020 5930 10380 5970
rect 10420 5930 10780 5970
rect 10820 5930 11180 5970
rect 11220 5930 11580 5970
rect 11620 5930 11980 5970
rect 12020 5930 12380 5970
rect 12420 5930 12780 5970
rect 12820 5930 13180 5970
rect 13220 5930 13580 5970
rect 13620 5930 13980 5970
rect 14020 5930 14380 5970
rect 14420 5930 14780 5970
rect 14820 5930 15180 5970
rect 15220 5930 15580 5970
rect 15620 5930 16000 5970
rect 0 5570 16000 5930
rect 0 5530 380 5570
rect 420 5530 780 5570
rect 820 5530 1180 5570
rect 1220 5530 1580 5570
rect 1620 5530 1980 5570
rect 2020 5530 2380 5570
rect 2420 5530 2780 5570
rect 2820 5530 3180 5570
rect 3220 5530 3580 5570
rect 3620 5530 3980 5570
rect 4020 5530 4380 5570
rect 4420 5530 4780 5570
rect 4820 5530 5180 5570
rect 5220 5530 5580 5570
rect 5620 5530 5980 5570
rect 6020 5530 6380 5570
rect 6420 5530 6780 5570
rect 6820 5530 7180 5570
rect 7220 5530 7580 5570
rect 7620 5530 7980 5570
rect 8020 5530 8380 5570
rect 8420 5530 8780 5570
rect 8820 5530 9180 5570
rect 9220 5530 9580 5570
rect 9620 5530 9980 5570
rect 10020 5530 10380 5570
rect 10420 5530 10780 5570
rect 10820 5530 11180 5570
rect 11220 5530 11580 5570
rect 11620 5530 11980 5570
rect 12020 5530 12380 5570
rect 12420 5530 12780 5570
rect 12820 5530 13180 5570
rect 13220 5530 13580 5570
rect 13620 5530 13980 5570
rect 14020 5530 14380 5570
rect 14420 5530 14780 5570
rect 14820 5530 15180 5570
rect 15220 5530 15580 5570
rect 15620 5530 16000 5570
rect 0 5170 16000 5530
rect 0 5130 380 5170
rect 420 5130 780 5170
rect 820 5130 1180 5170
rect 1220 5130 1580 5170
rect 1620 5130 1980 5170
rect 2020 5130 2380 5170
rect 2420 5130 2780 5170
rect 2820 5130 3180 5170
rect 3220 5130 3580 5170
rect 3620 5130 3980 5170
rect 4020 5130 4380 5170
rect 4420 5130 4780 5170
rect 4820 5130 5180 5170
rect 5220 5130 5580 5170
rect 5620 5130 5980 5170
rect 6020 5130 6380 5170
rect 6420 5130 6780 5170
rect 6820 5130 7180 5170
rect 7220 5130 7580 5170
rect 7620 5130 7980 5170
rect 8020 5130 8380 5170
rect 8420 5130 8780 5170
rect 8820 5130 9180 5170
rect 9220 5130 9580 5170
rect 9620 5130 9980 5170
rect 10020 5130 10380 5170
rect 10420 5130 10780 5170
rect 10820 5130 11180 5170
rect 11220 5130 11580 5170
rect 11620 5130 11980 5170
rect 12020 5130 12380 5170
rect 12420 5130 12780 5170
rect 12820 5130 13180 5170
rect 13220 5130 13580 5170
rect 13620 5130 13980 5170
rect 14020 5130 14380 5170
rect 14420 5130 14780 5170
rect 14820 5130 15180 5170
rect 15220 5130 15580 5170
rect 15620 5130 16000 5170
rect 0 4770 16000 5130
rect 0 4730 380 4770
rect 420 4730 780 4770
rect 820 4730 1180 4770
rect 1220 4730 1580 4770
rect 1620 4730 1980 4770
rect 2020 4730 2380 4770
rect 2420 4730 2780 4770
rect 2820 4730 3180 4770
rect 3220 4730 3580 4770
rect 3620 4730 3980 4770
rect 4020 4730 4380 4770
rect 4420 4730 4780 4770
rect 4820 4730 5180 4770
rect 5220 4730 5580 4770
rect 5620 4730 5980 4770
rect 6020 4730 6380 4770
rect 6420 4730 6780 4770
rect 6820 4730 7180 4770
rect 7220 4730 7580 4770
rect 7620 4730 7980 4770
rect 8020 4730 8380 4770
rect 8420 4730 8780 4770
rect 8820 4730 9180 4770
rect 9220 4730 9580 4770
rect 9620 4730 9980 4770
rect 10020 4730 10380 4770
rect 10420 4730 10780 4770
rect 10820 4730 11180 4770
rect 11220 4730 11580 4770
rect 11620 4730 11980 4770
rect 12020 4730 12380 4770
rect 12420 4730 12780 4770
rect 12820 4730 13180 4770
rect 13220 4730 13580 4770
rect 13620 4730 13980 4770
rect 14020 4730 14380 4770
rect 14420 4730 14780 4770
rect 14820 4730 15180 4770
rect 15220 4730 15580 4770
rect 15620 4730 16000 4770
rect 0 4370 16000 4730
rect 0 4330 380 4370
rect 420 4330 780 4370
rect 820 4330 1180 4370
rect 1220 4330 1580 4370
rect 1620 4330 1980 4370
rect 2020 4330 2380 4370
rect 2420 4330 2780 4370
rect 2820 4330 3180 4370
rect 3220 4330 3580 4370
rect 3620 4330 3980 4370
rect 4020 4330 4380 4370
rect 4420 4330 4780 4370
rect 4820 4330 5180 4370
rect 5220 4330 5580 4370
rect 5620 4330 5980 4370
rect 6020 4330 6380 4370
rect 6420 4330 6780 4370
rect 6820 4330 7180 4370
rect 7220 4330 7580 4370
rect 7620 4330 7980 4370
rect 8020 4330 8380 4370
rect 8420 4330 8780 4370
rect 8820 4330 9180 4370
rect 9220 4330 9580 4370
rect 9620 4330 9980 4370
rect 10020 4330 10380 4370
rect 10420 4330 10780 4370
rect 10820 4330 11180 4370
rect 11220 4330 11580 4370
rect 11620 4330 11980 4370
rect 12020 4330 12380 4370
rect 12420 4330 12780 4370
rect 12820 4330 13180 4370
rect 13220 4330 13580 4370
rect 13620 4330 13980 4370
rect 14020 4330 14380 4370
rect 14420 4330 14780 4370
rect 14820 4330 15180 4370
rect 15220 4330 15580 4370
rect 15620 4330 16000 4370
rect 0 3970 16000 4330
rect 0 3930 380 3970
rect 420 3930 780 3970
rect 820 3930 1180 3970
rect 1220 3930 1580 3970
rect 1620 3930 1980 3970
rect 2020 3930 2380 3970
rect 2420 3930 2780 3970
rect 2820 3930 3180 3970
rect 3220 3930 3580 3970
rect 3620 3930 3980 3970
rect 4020 3930 4380 3970
rect 4420 3930 4780 3970
rect 4820 3930 5180 3970
rect 5220 3930 5580 3970
rect 5620 3930 5980 3970
rect 6020 3930 6380 3970
rect 6420 3930 6780 3970
rect 6820 3930 7180 3970
rect 7220 3930 7580 3970
rect 7620 3930 7980 3970
rect 8020 3930 8380 3970
rect 8420 3930 8780 3970
rect 8820 3930 9180 3970
rect 9220 3930 9580 3970
rect 9620 3930 9980 3970
rect 10020 3930 10380 3970
rect 10420 3930 10780 3970
rect 10820 3930 11180 3970
rect 11220 3930 11580 3970
rect 11620 3930 11980 3970
rect 12020 3930 12380 3970
rect 12420 3930 12780 3970
rect 12820 3930 13180 3970
rect 13220 3930 13580 3970
rect 13620 3930 13980 3970
rect 14020 3930 14380 3970
rect 14420 3930 14780 3970
rect 14820 3930 15180 3970
rect 15220 3930 15580 3970
rect 15620 3930 16000 3970
rect 0 3570 16000 3930
rect 0 3530 380 3570
rect 420 3530 780 3570
rect 820 3530 1180 3570
rect 1220 3530 1580 3570
rect 1620 3530 1980 3570
rect 2020 3530 2380 3570
rect 2420 3530 2780 3570
rect 2820 3530 3180 3570
rect 3220 3530 3580 3570
rect 3620 3530 3980 3570
rect 4020 3530 4380 3570
rect 4420 3530 4780 3570
rect 4820 3530 5180 3570
rect 5220 3530 5580 3570
rect 5620 3530 5980 3570
rect 6020 3530 6380 3570
rect 6420 3530 6780 3570
rect 6820 3530 7180 3570
rect 7220 3530 7580 3570
rect 7620 3530 7980 3570
rect 8020 3530 8380 3570
rect 8420 3530 8780 3570
rect 8820 3530 9180 3570
rect 9220 3530 9580 3570
rect 9620 3530 9980 3570
rect 10020 3530 10380 3570
rect 10420 3530 10780 3570
rect 10820 3530 11180 3570
rect 11220 3530 11580 3570
rect 11620 3530 11980 3570
rect 12020 3530 12380 3570
rect 12420 3530 12780 3570
rect 12820 3530 13180 3570
rect 13220 3530 13580 3570
rect 13620 3530 13980 3570
rect 14020 3530 14380 3570
rect 14420 3530 14780 3570
rect 14820 3530 15180 3570
rect 15220 3530 15580 3570
rect 15620 3530 16000 3570
rect 0 3170 16000 3530
rect 0 3130 380 3170
rect 420 3130 780 3170
rect 820 3130 1180 3170
rect 1220 3130 1580 3170
rect 1620 3130 1980 3170
rect 2020 3130 2380 3170
rect 2420 3130 2780 3170
rect 2820 3130 3180 3170
rect 3220 3130 3580 3170
rect 3620 3130 3980 3170
rect 4020 3130 4380 3170
rect 4420 3130 4780 3170
rect 4820 3130 5180 3170
rect 5220 3130 5580 3170
rect 5620 3130 5980 3170
rect 6020 3130 6380 3170
rect 6420 3130 6780 3170
rect 6820 3130 7180 3170
rect 7220 3130 7580 3170
rect 7620 3130 7980 3170
rect 8020 3130 8380 3170
rect 8420 3130 8780 3170
rect 8820 3130 9180 3170
rect 9220 3130 9580 3170
rect 9620 3130 9980 3170
rect 10020 3130 10380 3170
rect 10420 3130 10780 3170
rect 10820 3130 11180 3170
rect 11220 3130 11580 3170
rect 11620 3130 11980 3170
rect 12020 3130 12380 3170
rect 12420 3130 12780 3170
rect 12820 3130 13180 3170
rect 13220 3130 13580 3170
rect 13620 3130 13980 3170
rect 14020 3130 14380 3170
rect 14420 3130 14780 3170
rect 14820 3130 15180 3170
rect 15220 3130 15580 3170
rect 15620 3130 16000 3170
rect 0 2770 16000 3130
rect 0 2730 380 2770
rect 420 2730 780 2770
rect 820 2730 1180 2770
rect 1220 2730 1580 2770
rect 1620 2730 1980 2770
rect 2020 2730 2380 2770
rect 2420 2730 2780 2770
rect 2820 2730 3180 2770
rect 3220 2730 3580 2770
rect 3620 2730 3980 2770
rect 4020 2730 4380 2770
rect 4420 2730 4780 2770
rect 4820 2730 5180 2770
rect 5220 2730 5580 2770
rect 5620 2730 5980 2770
rect 6020 2730 6380 2770
rect 6420 2730 6780 2770
rect 6820 2730 7180 2770
rect 7220 2730 7580 2770
rect 7620 2730 7980 2770
rect 8020 2730 8380 2770
rect 8420 2730 8780 2770
rect 8820 2730 9180 2770
rect 9220 2730 9580 2770
rect 9620 2730 9980 2770
rect 10020 2730 10380 2770
rect 10420 2730 10780 2770
rect 10820 2730 11180 2770
rect 11220 2730 11580 2770
rect 11620 2730 11980 2770
rect 12020 2730 12380 2770
rect 12420 2730 12780 2770
rect 12820 2730 13180 2770
rect 13220 2730 13580 2770
rect 13620 2730 13980 2770
rect 14020 2730 14380 2770
rect 14420 2730 14780 2770
rect 14820 2730 15180 2770
rect 15220 2730 15580 2770
rect 15620 2730 16000 2770
rect 0 2370 16000 2730
rect 0 2330 380 2370
rect 420 2330 780 2370
rect 820 2330 1180 2370
rect 1220 2330 1580 2370
rect 1620 2330 1980 2370
rect 2020 2330 2380 2370
rect 2420 2330 2780 2370
rect 2820 2330 3180 2370
rect 3220 2330 3580 2370
rect 3620 2330 3980 2370
rect 4020 2330 4380 2370
rect 4420 2330 4780 2370
rect 4820 2330 5180 2370
rect 5220 2330 5580 2370
rect 5620 2330 5980 2370
rect 6020 2330 6380 2370
rect 6420 2330 6780 2370
rect 6820 2330 7180 2370
rect 7220 2330 7580 2370
rect 7620 2330 7980 2370
rect 8020 2330 8380 2370
rect 8420 2330 8780 2370
rect 8820 2330 9180 2370
rect 9220 2330 9580 2370
rect 9620 2330 9980 2370
rect 10020 2330 10380 2370
rect 10420 2330 10780 2370
rect 10820 2330 11180 2370
rect 11220 2330 11580 2370
rect 11620 2330 11980 2370
rect 12020 2330 12380 2370
rect 12420 2330 12780 2370
rect 12820 2330 13180 2370
rect 13220 2330 13580 2370
rect 13620 2330 13980 2370
rect 14020 2330 14380 2370
rect 14420 2330 14780 2370
rect 14820 2330 15180 2370
rect 15220 2330 15580 2370
rect 15620 2330 16000 2370
rect 0 1970 16000 2330
rect 0 1930 380 1970
rect 420 1930 780 1970
rect 820 1930 1180 1970
rect 1220 1930 1580 1970
rect 1620 1930 1980 1970
rect 2020 1930 2380 1970
rect 2420 1930 2780 1970
rect 2820 1930 3180 1970
rect 3220 1930 3580 1970
rect 3620 1930 3980 1970
rect 4020 1930 4380 1970
rect 4420 1930 4780 1970
rect 4820 1930 5180 1970
rect 5220 1930 5580 1970
rect 5620 1930 5980 1970
rect 6020 1930 6380 1970
rect 6420 1930 6780 1970
rect 6820 1930 7180 1970
rect 7220 1930 7580 1970
rect 7620 1930 7980 1970
rect 8020 1930 8380 1970
rect 8420 1930 8780 1970
rect 8820 1930 9180 1970
rect 9220 1930 9580 1970
rect 9620 1930 9980 1970
rect 10020 1930 10380 1970
rect 10420 1930 10780 1970
rect 10820 1930 11180 1970
rect 11220 1930 11580 1970
rect 11620 1930 11980 1970
rect 12020 1930 12380 1970
rect 12420 1930 12780 1970
rect 12820 1930 13180 1970
rect 13220 1930 13580 1970
rect 13620 1930 13980 1970
rect 14020 1930 14380 1970
rect 14420 1930 14780 1970
rect 14820 1930 15180 1970
rect 15220 1930 15580 1970
rect 15620 1930 16000 1970
rect 0 1400 16000 1930
rect 1000 520 15000 600
rect 1000 480 1180 520
rect 1220 480 1580 520
rect 1620 480 1980 520
rect 2020 480 2380 520
rect 2420 480 2780 520
rect 2820 480 3180 520
rect 3220 480 3580 520
rect 3620 480 3980 520
rect 4020 480 4380 520
rect 4420 480 4780 520
rect 4820 480 5180 520
rect 5220 480 5580 520
rect 5620 480 5980 520
rect 6020 480 6380 520
rect 6420 480 6780 520
rect 6820 480 7180 520
rect 7220 480 7580 520
rect 7620 480 7980 520
rect 8020 480 8380 520
rect 8420 480 8780 520
rect 8820 480 9180 520
rect 9220 480 9580 520
rect 9620 480 9980 520
rect 10020 480 10380 520
rect 10420 480 10780 520
rect 10820 480 11180 520
rect 11220 480 11580 520
rect 11620 480 11980 520
rect 12020 480 12380 520
rect 12420 480 12780 520
rect 12820 480 13180 520
rect 13220 480 13580 520
rect 13620 480 13980 520
rect 14020 480 14380 520
rect 14420 480 14780 520
rect 14820 480 15000 520
rect 1000 120 15000 480
rect 1000 80 1180 120
rect 1220 80 1580 120
rect 1620 80 1980 120
rect 2020 80 2380 120
rect 2420 80 2780 120
rect 2820 80 3180 120
rect 3220 80 3580 120
rect 3620 80 3980 120
rect 4020 80 4380 120
rect 4420 80 4780 120
rect 4820 80 5180 120
rect 5220 80 5580 120
rect 5620 80 5980 120
rect 6020 80 6380 120
rect 6420 80 6780 120
rect 6820 80 7180 120
rect 7220 80 7580 120
rect 7620 80 7980 120
rect 8020 80 8380 120
rect 8420 80 8780 120
rect 8820 80 9180 120
rect 9220 80 9580 120
rect 9620 80 9980 120
rect 10020 80 10380 120
rect 10420 80 10780 120
rect 10820 80 11180 120
rect 11220 80 11580 120
rect 11620 80 11980 120
rect 12020 80 12380 120
rect 12420 80 12780 120
rect 12820 80 13180 120
rect 13220 80 13580 120
rect 13620 80 13980 120
rect 14020 80 14380 120
rect 14420 80 14780 120
rect 14820 80 15000 120
rect 1000 0 15000 80
<< via4 >>
rect 380 35000 420 35040
rect 780 35000 820 35040
rect 1180 35000 1220 35040
rect 1580 35000 1620 35040
rect 1980 35000 2020 35040
rect 2380 35000 2420 35040
rect 2780 35000 2820 35040
rect 3180 35000 3220 35040
rect 3580 35000 3620 35040
rect 3980 35000 4020 35040
rect 4380 35000 4420 35040
rect 4780 35000 4820 35040
rect 5180 35000 5220 35040
rect 5580 35000 5620 35040
rect 5980 35000 6020 35040
rect 6380 35000 6420 35040
rect 6780 35000 6820 35040
rect 7180 35000 7220 35040
rect 7580 35000 7620 35040
rect 7980 35000 8020 35040
rect 8380 35000 8420 35040
rect 8780 35000 8820 35040
rect 9180 35000 9220 35040
rect 9580 35000 9620 35040
rect 9980 35000 10020 35040
rect 10380 35000 10420 35040
rect 10780 35000 10820 35040
rect 11180 35000 11220 35040
rect 11580 35000 11620 35040
rect 11980 35000 12020 35040
rect 12380 35000 12420 35040
rect 12780 35000 12820 35040
rect 13180 35000 13220 35040
rect 13580 35000 13620 35040
rect 13980 35000 14020 35040
rect 14380 35000 14420 35040
rect 14780 35000 14820 35040
rect 15180 35000 15220 35040
rect 15580 35000 15620 35040
rect 380 34600 420 34640
rect 780 34600 820 34640
rect 1180 34600 1220 34640
rect 1580 34600 1620 34640
rect 1980 34600 2020 34640
rect 2380 34600 2420 34640
rect 2780 34600 2820 34640
rect 3180 34600 3220 34640
rect 3580 34600 3620 34640
rect 3980 34600 4020 34640
rect 4380 34600 4420 34640
rect 4780 34600 4820 34640
rect 5180 34600 5220 34640
rect 5580 34600 5620 34640
rect 5980 34600 6020 34640
rect 6380 34600 6420 34640
rect 6780 34600 6820 34640
rect 7180 34600 7220 34640
rect 7580 34600 7620 34640
rect 7980 34600 8020 34640
rect 8380 34600 8420 34640
rect 8780 34600 8820 34640
rect 9180 34600 9220 34640
rect 9580 34600 9620 34640
rect 9980 34600 10020 34640
rect 10380 34600 10420 34640
rect 10780 34600 10820 34640
rect 11180 34600 11220 34640
rect 11580 34600 11620 34640
rect 11980 34600 12020 34640
rect 12380 34600 12420 34640
rect 12780 34600 12820 34640
rect 13180 34600 13220 34640
rect 13580 34600 13620 34640
rect 13980 34600 14020 34640
rect 14380 34600 14420 34640
rect 14780 34600 14820 34640
rect 15180 34600 15220 34640
rect 15580 34600 15620 34640
rect 380 34200 420 34240
rect 780 34200 820 34240
rect 1180 34200 1220 34240
rect 1580 34200 1620 34240
rect 1980 34200 2020 34240
rect 2380 34200 2420 34240
rect 2780 34200 2820 34240
rect 3180 34200 3220 34240
rect 3580 34200 3620 34240
rect 3980 34200 4020 34240
rect 4380 34200 4420 34240
rect 4780 34200 4820 34240
rect 5180 34200 5220 34240
rect 5580 34200 5620 34240
rect 5980 34200 6020 34240
rect 6380 34200 6420 34240
rect 6780 34200 6820 34240
rect 7180 34200 7220 34240
rect 7580 34200 7620 34240
rect 7980 34200 8020 34240
rect 8380 34200 8420 34240
rect 8780 34200 8820 34240
rect 9180 34200 9220 34240
rect 9580 34200 9620 34240
rect 9980 34200 10020 34240
rect 10380 34200 10420 34240
rect 10780 34200 10820 34240
rect 11180 34200 11220 34240
rect 11580 34200 11620 34240
rect 11980 34200 12020 34240
rect 12380 34200 12420 34240
rect 12780 34200 12820 34240
rect 13180 34200 13220 34240
rect 13580 34200 13620 34240
rect 13980 34200 14020 34240
rect 14380 34200 14420 34240
rect 14780 34200 14820 34240
rect 15180 34200 15220 34240
rect 15580 34200 15620 34240
rect 380 33800 420 33840
rect 780 33800 820 33840
rect 1180 33800 1220 33840
rect 1580 33800 1620 33840
rect 1980 33800 2020 33840
rect 2380 33800 2420 33840
rect 2780 33800 2820 33840
rect 3180 33800 3220 33840
rect 3580 33800 3620 33840
rect 3980 33800 4020 33840
rect 4380 33800 4420 33840
rect 4780 33800 4820 33840
rect 5180 33800 5220 33840
rect 5580 33800 5620 33840
rect 5980 33800 6020 33840
rect 6380 33800 6420 33840
rect 6780 33800 6820 33840
rect 7180 33800 7220 33840
rect 7580 33800 7620 33840
rect 7980 33800 8020 33840
rect 8380 33800 8420 33840
rect 8780 33800 8820 33840
rect 9180 33800 9220 33840
rect 9580 33800 9620 33840
rect 9980 33800 10020 33840
rect 10380 33800 10420 33840
rect 10780 33800 10820 33840
rect 11180 33800 11220 33840
rect 11580 33800 11620 33840
rect 11980 33800 12020 33840
rect 12380 33800 12420 33840
rect 12780 33800 12820 33840
rect 13180 33800 13220 33840
rect 13580 33800 13620 33840
rect 13980 33800 14020 33840
rect 14380 33800 14420 33840
rect 14780 33800 14820 33840
rect 15180 33800 15220 33840
rect 15580 33800 15620 33840
rect 380 33400 420 33440
rect 780 33400 820 33440
rect 1180 33400 1220 33440
rect 1580 33400 1620 33440
rect 1980 33400 2020 33440
rect 2380 33400 2420 33440
rect 2780 33400 2820 33440
rect 3180 33400 3220 33440
rect 3580 33400 3620 33440
rect 3980 33400 4020 33440
rect 4380 33400 4420 33440
rect 4780 33400 4820 33440
rect 5180 33400 5220 33440
rect 5580 33400 5620 33440
rect 5980 33400 6020 33440
rect 6380 33400 6420 33440
rect 6780 33400 6820 33440
rect 7180 33400 7220 33440
rect 7580 33400 7620 33440
rect 7980 33400 8020 33440
rect 8380 33400 8420 33440
rect 8780 33400 8820 33440
rect 9180 33400 9220 33440
rect 9580 33400 9620 33440
rect 9980 33400 10020 33440
rect 10380 33400 10420 33440
rect 10780 33400 10820 33440
rect 11180 33400 11220 33440
rect 11580 33400 11620 33440
rect 11980 33400 12020 33440
rect 12380 33400 12420 33440
rect 12780 33400 12820 33440
rect 13180 33400 13220 33440
rect 13580 33400 13620 33440
rect 13980 33400 14020 33440
rect 14380 33400 14420 33440
rect 14780 33400 14820 33440
rect 15180 33400 15220 33440
rect 15580 33400 15620 33440
rect 380 33000 420 33040
rect 780 33000 820 33040
rect 1180 33000 1220 33040
rect 1580 33000 1620 33040
rect 1980 33000 2020 33040
rect 2380 33000 2420 33040
rect 2780 33000 2820 33040
rect 3180 33000 3220 33040
rect 3580 33000 3620 33040
rect 3980 33000 4020 33040
rect 4380 33000 4420 33040
rect 4780 33000 4820 33040
rect 5180 33000 5220 33040
rect 5580 33000 5620 33040
rect 5980 33000 6020 33040
rect 6380 33000 6420 33040
rect 6780 33000 6820 33040
rect 7180 33000 7220 33040
rect 7580 33000 7620 33040
rect 7980 33000 8020 33040
rect 8380 33000 8420 33040
rect 8780 33000 8820 33040
rect 9180 33000 9220 33040
rect 9580 33000 9620 33040
rect 9980 33000 10020 33040
rect 10380 33000 10420 33040
rect 10780 33000 10820 33040
rect 11180 33000 11220 33040
rect 11580 33000 11620 33040
rect 11980 33000 12020 33040
rect 12380 33000 12420 33040
rect 12780 33000 12820 33040
rect 13180 33000 13220 33040
rect 13580 33000 13620 33040
rect 13980 33000 14020 33040
rect 14380 33000 14420 33040
rect 14780 33000 14820 33040
rect 15180 33000 15220 33040
rect 15580 33000 15620 33040
rect 380 30560 420 30600
rect 780 30560 820 30600
rect 1180 30560 1220 30600
rect 1580 30560 1620 30600
rect 1980 30560 2020 30600
rect 2380 30560 2420 30600
rect 2780 30560 2820 30600
rect 3180 30560 3220 30600
rect 3580 30560 3620 30600
rect 3980 30560 4020 30600
rect 4380 30560 4420 30600
rect 4780 30560 4820 30600
rect 5180 30560 5220 30600
rect 5580 30560 5620 30600
rect 5980 30560 6020 30600
rect 6380 30560 6420 30600
rect 6780 30560 6820 30600
rect 7180 30560 7220 30600
rect 7580 30560 7620 30600
rect 7980 30560 8020 30600
rect 8380 30560 8420 30600
rect 8780 30560 8820 30600
rect 9180 30560 9220 30600
rect 9580 30560 9620 30600
rect 9980 30560 10020 30600
rect 10380 30560 10420 30600
rect 10780 30560 10820 30600
rect 11180 30560 11220 30600
rect 11580 30560 11620 30600
rect 11980 30560 12020 30600
rect 12380 30560 12420 30600
rect 12780 30560 12820 30600
rect 13180 30560 13220 30600
rect 13580 30560 13620 30600
rect 13980 30560 14020 30600
rect 14380 30560 14420 30600
rect 14780 30560 14820 30600
rect 15180 30560 15220 30600
rect 15580 30560 15620 30600
rect 380 30160 420 30200
rect 780 30160 820 30200
rect 1180 30160 1220 30200
rect 1580 30160 1620 30200
rect 1980 30160 2020 30200
rect 2380 30160 2420 30200
rect 2780 30160 2820 30200
rect 3180 30160 3220 30200
rect 3580 30160 3620 30200
rect 3980 30160 4020 30200
rect 4380 30160 4420 30200
rect 4780 30160 4820 30200
rect 5180 30160 5220 30200
rect 5580 30160 5620 30200
rect 5980 30160 6020 30200
rect 6380 30160 6420 30200
rect 6780 30160 6820 30200
rect 7180 30160 7220 30200
rect 7580 30160 7620 30200
rect 7980 30160 8020 30200
rect 8380 30160 8420 30200
rect 8780 30160 8820 30200
rect 9180 30160 9220 30200
rect 9580 30160 9620 30200
rect 9980 30160 10020 30200
rect 10380 30160 10420 30200
rect 10780 30160 10820 30200
rect 11180 30160 11220 30200
rect 11580 30160 11620 30200
rect 11980 30160 12020 30200
rect 12380 30160 12420 30200
rect 12780 30160 12820 30200
rect 13180 30160 13220 30200
rect 13580 30160 13620 30200
rect 13980 30160 14020 30200
rect 14380 30160 14420 30200
rect 14780 30160 14820 30200
rect 15180 30160 15220 30200
rect 15580 30160 15620 30200
rect 380 29760 420 29800
rect 780 29760 820 29800
rect 1180 29760 1220 29800
rect 1580 29760 1620 29800
rect 1980 29760 2020 29800
rect 2380 29760 2420 29800
rect 2780 29760 2820 29800
rect 3180 29760 3220 29800
rect 3580 29760 3620 29800
rect 3980 29760 4020 29800
rect 4380 29760 4420 29800
rect 4780 29760 4820 29800
rect 5180 29760 5220 29800
rect 5580 29760 5620 29800
rect 5980 29760 6020 29800
rect 6380 29760 6420 29800
rect 6780 29760 6820 29800
rect 7180 29760 7220 29800
rect 7580 29760 7620 29800
rect 7980 29760 8020 29800
rect 8380 29760 8420 29800
rect 8780 29760 8820 29800
rect 9180 29760 9220 29800
rect 9580 29760 9620 29800
rect 9980 29760 10020 29800
rect 10380 29760 10420 29800
rect 10780 29760 10820 29800
rect 11180 29760 11220 29800
rect 11580 29760 11620 29800
rect 11980 29760 12020 29800
rect 12380 29760 12420 29800
rect 12780 29760 12820 29800
rect 13180 29760 13220 29800
rect 13580 29760 13620 29800
rect 13980 29760 14020 29800
rect 14380 29760 14420 29800
rect 14780 29760 14820 29800
rect 15180 29760 15220 29800
rect 15580 29760 15620 29800
rect 380 29360 420 29400
rect 780 29360 820 29400
rect 1180 29360 1220 29400
rect 1580 29360 1620 29400
rect 1980 29360 2020 29400
rect 2380 29360 2420 29400
rect 2780 29360 2820 29400
rect 3180 29360 3220 29400
rect 3580 29360 3620 29400
rect 3980 29360 4020 29400
rect 4380 29360 4420 29400
rect 4780 29360 4820 29400
rect 5180 29360 5220 29400
rect 5580 29360 5620 29400
rect 5980 29360 6020 29400
rect 6380 29360 6420 29400
rect 6780 29360 6820 29400
rect 7180 29360 7220 29400
rect 7580 29360 7620 29400
rect 7980 29360 8020 29400
rect 8380 29360 8420 29400
rect 8780 29360 8820 29400
rect 9180 29360 9220 29400
rect 9580 29360 9620 29400
rect 9980 29360 10020 29400
rect 10380 29360 10420 29400
rect 10780 29360 10820 29400
rect 11180 29360 11220 29400
rect 11580 29360 11620 29400
rect 11980 29360 12020 29400
rect 12380 29360 12420 29400
rect 12780 29360 12820 29400
rect 13180 29360 13220 29400
rect 13580 29360 13620 29400
rect 13980 29360 14020 29400
rect 14380 29360 14420 29400
rect 14780 29360 14820 29400
rect 15180 29360 15220 29400
rect 15580 29360 15620 29400
rect 380 28960 420 29000
rect 780 28960 820 29000
rect 1180 28960 1220 29000
rect 1580 28960 1620 29000
rect 1980 28960 2020 29000
rect 2380 28960 2420 29000
rect 2780 28960 2820 29000
rect 3180 28960 3220 29000
rect 3580 28960 3620 29000
rect 3980 28960 4020 29000
rect 4380 28960 4420 29000
rect 4780 28960 4820 29000
rect 5180 28960 5220 29000
rect 5580 28960 5620 29000
rect 5980 28960 6020 29000
rect 6380 28960 6420 29000
rect 6780 28960 6820 29000
rect 7180 28960 7220 29000
rect 7580 28960 7620 29000
rect 7980 28960 8020 29000
rect 8380 28960 8420 29000
rect 8780 28960 8820 29000
rect 9180 28960 9220 29000
rect 9580 28960 9620 29000
rect 9980 28960 10020 29000
rect 10380 28960 10420 29000
rect 10780 28960 10820 29000
rect 11180 28960 11220 29000
rect 11580 28960 11620 29000
rect 11980 28960 12020 29000
rect 12380 28960 12420 29000
rect 12780 28960 12820 29000
rect 13180 28960 13220 29000
rect 13580 28960 13620 29000
rect 13980 28960 14020 29000
rect 14380 28960 14420 29000
rect 14780 28960 14820 29000
rect 15180 28960 15220 29000
rect 15580 28960 15620 29000
rect 380 28560 420 28600
rect 780 28560 820 28600
rect 1180 28560 1220 28600
rect 1580 28560 1620 28600
rect 1980 28560 2020 28600
rect 2380 28560 2420 28600
rect 2780 28560 2820 28600
rect 3180 28560 3220 28600
rect 3580 28560 3620 28600
rect 3980 28560 4020 28600
rect 4380 28560 4420 28600
rect 4780 28560 4820 28600
rect 5180 28560 5220 28600
rect 5580 28560 5620 28600
rect 5980 28560 6020 28600
rect 6380 28560 6420 28600
rect 6780 28560 6820 28600
rect 7180 28560 7220 28600
rect 7580 28560 7620 28600
rect 7980 28560 8020 28600
rect 8380 28560 8420 28600
rect 8780 28560 8820 28600
rect 9180 28560 9220 28600
rect 9580 28560 9620 28600
rect 9980 28560 10020 28600
rect 10380 28560 10420 28600
rect 10780 28560 10820 28600
rect 11180 28560 11220 28600
rect 11580 28560 11620 28600
rect 11980 28560 12020 28600
rect 12380 28560 12420 28600
rect 12780 28560 12820 28600
rect 13180 28560 13220 28600
rect 13580 28560 13620 28600
rect 13980 28560 14020 28600
rect 14380 28560 14420 28600
rect 14780 28560 14820 28600
rect 15180 28560 15220 28600
rect 15580 28560 15620 28600
rect 380 26380 420 26420
rect 780 26380 820 26420
rect 1180 26380 1220 26420
rect 1580 26380 1620 26420
rect 1980 26380 2020 26420
rect 2380 26380 2420 26420
rect 2780 26380 2820 26420
rect 3180 26380 3220 26420
rect 3580 26380 3620 26420
rect 3980 26380 4020 26420
rect 4380 26380 4420 26420
rect 4780 26380 4820 26420
rect 5180 26380 5220 26420
rect 5580 26380 5620 26420
rect 5980 26380 6020 26420
rect 6380 26380 6420 26420
rect 6780 26380 6820 26420
rect 7180 26380 7220 26420
rect 7580 26380 7620 26420
rect 7980 26380 8020 26420
rect 8380 26380 8420 26420
rect 8780 26380 8820 26420
rect 9180 26380 9220 26420
rect 9580 26380 9620 26420
rect 9980 26380 10020 26420
rect 10380 26380 10420 26420
rect 10780 26380 10820 26420
rect 11180 26380 11220 26420
rect 11580 26380 11620 26420
rect 11980 26380 12020 26420
rect 12380 26380 12420 26420
rect 12780 26380 12820 26420
rect 13180 26380 13220 26420
rect 13580 26380 13620 26420
rect 13980 26380 14020 26420
rect 14380 26380 14420 26420
rect 14780 26380 14820 26420
rect 15180 26380 15220 26420
rect 15580 26380 15620 26420
rect 380 25980 420 26020
rect 780 25980 820 26020
rect 1180 25980 1220 26020
rect 1580 25980 1620 26020
rect 1980 25980 2020 26020
rect 2380 25980 2420 26020
rect 2780 25980 2820 26020
rect 3180 25980 3220 26020
rect 3580 25980 3620 26020
rect 3980 25980 4020 26020
rect 4380 25980 4420 26020
rect 4780 25980 4820 26020
rect 5180 25980 5220 26020
rect 5580 25980 5620 26020
rect 5980 25980 6020 26020
rect 6380 25980 6420 26020
rect 6780 25980 6820 26020
rect 7180 25980 7220 26020
rect 7580 25980 7620 26020
rect 7980 25980 8020 26020
rect 8380 25980 8420 26020
rect 8780 25980 8820 26020
rect 9180 25980 9220 26020
rect 9580 25980 9620 26020
rect 9980 25980 10020 26020
rect 10380 25980 10420 26020
rect 10780 25980 10820 26020
rect 11180 25980 11220 26020
rect 11580 25980 11620 26020
rect 11980 25980 12020 26020
rect 12380 25980 12420 26020
rect 12780 25980 12820 26020
rect 13180 25980 13220 26020
rect 13580 25980 13620 26020
rect 13980 25980 14020 26020
rect 14380 25980 14420 26020
rect 14780 25980 14820 26020
rect 15180 25980 15220 26020
rect 15580 25980 15620 26020
rect 380 25580 420 25620
rect 780 25580 820 25620
rect 1180 25580 1220 25620
rect 1580 25580 1620 25620
rect 1980 25580 2020 25620
rect 2380 25580 2420 25620
rect 2780 25580 2820 25620
rect 3180 25580 3220 25620
rect 3580 25580 3620 25620
rect 3980 25580 4020 25620
rect 4380 25580 4420 25620
rect 4780 25580 4820 25620
rect 5180 25580 5220 25620
rect 5580 25580 5620 25620
rect 5980 25580 6020 25620
rect 6380 25580 6420 25620
rect 6780 25580 6820 25620
rect 7180 25580 7220 25620
rect 7580 25580 7620 25620
rect 7980 25580 8020 25620
rect 8380 25580 8420 25620
rect 8780 25580 8820 25620
rect 9180 25580 9220 25620
rect 9580 25580 9620 25620
rect 9980 25580 10020 25620
rect 10380 25580 10420 25620
rect 10780 25580 10820 25620
rect 11180 25580 11220 25620
rect 11580 25580 11620 25620
rect 11980 25580 12020 25620
rect 12380 25580 12420 25620
rect 12780 25580 12820 25620
rect 13180 25580 13220 25620
rect 13580 25580 13620 25620
rect 13980 25580 14020 25620
rect 14380 25580 14420 25620
rect 14780 25580 14820 25620
rect 15180 25580 15220 25620
rect 15580 25580 15620 25620
rect 380 23230 420 23270
rect 780 23230 820 23270
rect 1180 23230 1220 23270
rect 1580 23230 1620 23270
rect 1980 23230 2020 23270
rect 2380 23230 2420 23270
rect 2780 23230 2820 23270
rect 3180 23230 3220 23270
rect 3580 23230 3620 23270
rect 3980 23230 4020 23270
rect 4380 23230 4420 23270
rect 4780 23230 4820 23270
rect 5180 23230 5220 23270
rect 5580 23230 5620 23270
rect 5980 23230 6020 23270
rect 6380 23230 6420 23270
rect 6780 23230 6820 23270
rect 7180 23230 7220 23270
rect 7580 23230 7620 23270
rect 7980 23230 8020 23270
rect 8380 23230 8420 23270
rect 8780 23230 8820 23270
rect 9180 23230 9220 23270
rect 9580 23230 9620 23270
rect 9980 23230 10020 23270
rect 10380 23230 10420 23270
rect 10780 23230 10820 23270
rect 11180 23230 11220 23270
rect 11580 23230 11620 23270
rect 11980 23230 12020 23270
rect 12380 23230 12420 23270
rect 12780 23230 12820 23270
rect 13180 23230 13220 23270
rect 13580 23230 13620 23270
rect 13980 23230 14020 23270
rect 14380 23230 14420 23270
rect 14780 23230 14820 23270
rect 15180 23230 15220 23270
rect 15580 23230 15620 23270
rect 380 22830 420 22870
rect 780 22830 820 22870
rect 1180 22830 1220 22870
rect 1580 22830 1620 22870
rect 1980 22830 2020 22870
rect 2380 22830 2420 22870
rect 2780 22830 2820 22870
rect 3180 22830 3220 22870
rect 3580 22830 3620 22870
rect 3980 22830 4020 22870
rect 4380 22830 4420 22870
rect 4780 22830 4820 22870
rect 5180 22830 5220 22870
rect 5580 22830 5620 22870
rect 5980 22830 6020 22870
rect 6380 22830 6420 22870
rect 6780 22830 6820 22870
rect 7180 22830 7220 22870
rect 7580 22830 7620 22870
rect 7980 22830 8020 22870
rect 8380 22830 8420 22870
rect 8780 22830 8820 22870
rect 9180 22830 9220 22870
rect 9580 22830 9620 22870
rect 9980 22830 10020 22870
rect 10380 22830 10420 22870
rect 10780 22830 10820 22870
rect 11180 22830 11220 22870
rect 11580 22830 11620 22870
rect 11980 22830 12020 22870
rect 12380 22830 12420 22870
rect 12780 22830 12820 22870
rect 13180 22830 13220 22870
rect 13580 22830 13620 22870
rect 13980 22830 14020 22870
rect 14380 22830 14420 22870
rect 14780 22830 14820 22870
rect 15180 22830 15220 22870
rect 15580 22830 15620 22870
rect 380 22430 420 22470
rect 780 22430 820 22470
rect 1180 22430 1220 22470
rect 1580 22430 1620 22470
rect 1980 22430 2020 22470
rect 2380 22430 2420 22470
rect 2780 22430 2820 22470
rect 3180 22430 3220 22470
rect 3580 22430 3620 22470
rect 3980 22430 4020 22470
rect 4380 22430 4420 22470
rect 4780 22430 4820 22470
rect 5180 22430 5220 22470
rect 5580 22430 5620 22470
rect 5980 22430 6020 22470
rect 6380 22430 6420 22470
rect 6780 22430 6820 22470
rect 7180 22430 7220 22470
rect 7580 22430 7620 22470
rect 7980 22430 8020 22470
rect 8380 22430 8420 22470
rect 8780 22430 8820 22470
rect 9180 22430 9220 22470
rect 9580 22430 9620 22470
rect 9980 22430 10020 22470
rect 10380 22430 10420 22470
rect 10780 22430 10820 22470
rect 11180 22430 11220 22470
rect 11580 22430 11620 22470
rect 11980 22430 12020 22470
rect 12380 22430 12420 22470
rect 12780 22430 12820 22470
rect 13180 22430 13220 22470
rect 13580 22430 13620 22470
rect 13980 22430 14020 22470
rect 14380 22430 14420 22470
rect 14780 22430 14820 22470
rect 15180 22430 15220 22470
rect 15580 22430 15620 22470
rect 380 22030 420 22070
rect 780 22030 820 22070
rect 1180 22030 1220 22070
rect 1580 22030 1620 22070
rect 1980 22030 2020 22070
rect 2380 22030 2420 22070
rect 2780 22030 2820 22070
rect 3180 22030 3220 22070
rect 3580 22030 3620 22070
rect 3980 22030 4020 22070
rect 4380 22030 4420 22070
rect 4780 22030 4820 22070
rect 5180 22030 5220 22070
rect 5580 22030 5620 22070
rect 5980 22030 6020 22070
rect 6380 22030 6420 22070
rect 6780 22030 6820 22070
rect 7180 22030 7220 22070
rect 7580 22030 7620 22070
rect 7980 22030 8020 22070
rect 8380 22030 8420 22070
rect 8780 22030 8820 22070
rect 9180 22030 9220 22070
rect 9580 22030 9620 22070
rect 9980 22030 10020 22070
rect 10380 22030 10420 22070
rect 10780 22030 10820 22070
rect 11180 22030 11220 22070
rect 11580 22030 11620 22070
rect 11980 22030 12020 22070
rect 12380 22030 12420 22070
rect 12780 22030 12820 22070
rect 13180 22030 13220 22070
rect 13580 22030 13620 22070
rect 13980 22030 14020 22070
rect 14380 22030 14420 22070
rect 14780 22030 14820 22070
rect 15180 22030 15220 22070
rect 15580 22030 15620 22070
rect 380 21630 420 21670
rect 780 21630 820 21670
rect 1180 21630 1220 21670
rect 1580 21630 1620 21670
rect 1980 21630 2020 21670
rect 2380 21630 2420 21670
rect 2780 21630 2820 21670
rect 3180 21630 3220 21670
rect 3580 21630 3620 21670
rect 3980 21630 4020 21670
rect 4380 21630 4420 21670
rect 4780 21630 4820 21670
rect 5180 21630 5220 21670
rect 5580 21630 5620 21670
rect 5980 21630 6020 21670
rect 6380 21630 6420 21670
rect 6780 21630 6820 21670
rect 7180 21630 7220 21670
rect 7580 21630 7620 21670
rect 7980 21630 8020 21670
rect 8380 21630 8420 21670
rect 8780 21630 8820 21670
rect 9180 21630 9220 21670
rect 9580 21630 9620 21670
rect 9980 21630 10020 21670
rect 10380 21630 10420 21670
rect 10780 21630 10820 21670
rect 11180 21630 11220 21670
rect 11580 21630 11620 21670
rect 11980 21630 12020 21670
rect 12380 21630 12420 21670
rect 12780 21630 12820 21670
rect 13180 21630 13220 21670
rect 13580 21630 13620 21670
rect 13980 21630 14020 21670
rect 14380 21630 14420 21670
rect 14780 21630 14820 21670
rect 15180 21630 15220 21670
rect 15580 21630 15620 21670
rect 380 21230 420 21270
rect 780 21230 820 21270
rect 1180 21230 1220 21270
rect 1580 21230 1620 21270
rect 1980 21230 2020 21270
rect 2380 21230 2420 21270
rect 2780 21230 2820 21270
rect 3180 21230 3220 21270
rect 3580 21230 3620 21270
rect 3980 21230 4020 21270
rect 4380 21230 4420 21270
rect 4780 21230 4820 21270
rect 5180 21230 5220 21270
rect 5580 21230 5620 21270
rect 5980 21230 6020 21270
rect 6380 21230 6420 21270
rect 6780 21230 6820 21270
rect 7180 21230 7220 21270
rect 7580 21230 7620 21270
rect 7980 21230 8020 21270
rect 8380 21230 8420 21270
rect 8780 21230 8820 21270
rect 9180 21230 9220 21270
rect 9580 21230 9620 21270
rect 9980 21230 10020 21270
rect 10380 21230 10420 21270
rect 10780 21230 10820 21270
rect 11180 21230 11220 21270
rect 11580 21230 11620 21270
rect 11980 21230 12020 21270
rect 12380 21230 12420 21270
rect 12780 21230 12820 21270
rect 13180 21230 13220 21270
rect 13580 21230 13620 21270
rect 13980 21230 14020 21270
rect 14380 21230 14420 21270
rect 14780 21230 14820 21270
rect 15180 21230 15220 21270
rect 15580 21230 15620 21270
rect 380 20830 420 20870
rect 780 20830 820 20870
rect 1180 20830 1220 20870
rect 1580 20830 1620 20870
rect 1980 20830 2020 20870
rect 2380 20830 2420 20870
rect 2780 20830 2820 20870
rect 3180 20830 3220 20870
rect 3580 20830 3620 20870
rect 3980 20830 4020 20870
rect 4380 20830 4420 20870
rect 4780 20830 4820 20870
rect 5180 20830 5220 20870
rect 5580 20830 5620 20870
rect 5980 20830 6020 20870
rect 6380 20830 6420 20870
rect 6780 20830 6820 20870
rect 7180 20830 7220 20870
rect 7580 20830 7620 20870
rect 7980 20830 8020 20870
rect 8380 20830 8420 20870
rect 8780 20830 8820 20870
rect 9180 20830 9220 20870
rect 9580 20830 9620 20870
rect 9980 20830 10020 20870
rect 10380 20830 10420 20870
rect 10780 20830 10820 20870
rect 11180 20830 11220 20870
rect 11580 20830 11620 20870
rect 11980 20830 12020 20870
rect 12380 20830 12420 20870
rect 12780 20830 12820 20870
rect 13180 20830 13220 20870
rect 13580 20830 13620 20870
rect 13980 20830 14020 20870
rect 14380 20830 14420 20870
rect 14780 20830 14820 20870
rect 15180 20830 15220 20870
rect 15580 20830 15620 20870
rect 380 20430 420 20470
rect 780 20430 820 20470
rect 1180 20430 1220 20470
rect 1580 20430 1620 20470
rect 1980 20430 2020 20470
rect 2380 20430 2420 20470
rect 2780 20430 2820 20470
rect 3180 20430 3220 20470
rect 3580 20430 3620 20470
rect 3980 20430 4020 20470
rect 4380 20430 4420 20470
rect 4780 20430 4820 20470
rect 5180 20430 5220 20470
rect 5580 20430 5620 20470
rect 5980 20430 6020 20470
rect 6380 20430 6420 20470
rect 6780 20430 6820 20470
rect 7180 20430 7220 20470
rect 7580 20430 7620 20470
rect 7980 20430 8020 20470
rect 8380 20430 8420 20470
rect 8780 20430 8820 20470
rect 9180 20430 9220 20470
rect 9580 20430 9620 20470
rect 9980 20430 10020 20470
rect 10380 20430 10420 20470
rect 10780 20430 10820 20470
rect 11180 20430 11220 20470
rect 11580 20430 11620 20470
rect 11980 20430 12020 20470
rect 12380 20430 12420 20470
rect 12780 20430 12820 20470
rect 13180 20430 13220 20470
rect 13580 20430 13620 20470
rect 13980 20430 14020 20470
rect 14380 20430 14420 20470
rect 14780 20430 14820 20470
rect 15180 20430 15220 20470
rect 15580 20430 15620 20470
rect 380 20030 420 20070
rect 780 20030 820 20070
rect 1180 20030 1220 20070
rect 1580 20030 1620 20070
rect 1980 20030 2020 20070
rect 2380 20030 2420 20070
rect 2780 20030 2820 20070
rect 3180 20030 3220 20070
rect 3580 20030 3620 20070
rect 3980 20030 4020 20070
rect 4380 20030 4420 20070
rect 4780 20030 4820 20070
rect 5180 20030 5220 20070
rect 5580 20030 5620 20070
rect 5980 20030 6020 20070
rect 6380 20030 6420 20070
rect 6780 20030 6820 20070
rect 7180 20030 7220 20070
rect 7580 20030 7620 20070
rect 7980 20030 8020 20070
rect 8380 20030 8420 20070
rect 8780 20030 8820 20070
rect 9180 20030 9220 20070
rect 9580 20030 9620 20070
rect 9980 20030 10020 20070
rect 10380 20030 10420 20070
rect 10780 20030 10820 20070
rect 11180 20030 11220 20070
rect 11580 20030 11620 20070
rect 11980 20030 12020 20070
rect 12380 20030 12420 20070
rect 12780 20030 12820 20070
rect 13180 20030 13220 20070
rect 13580 20030 13620 20070
rect 13980 20030 14020 20070
rect 14380 20030 14420 20070
rect 14780 20030 14820 20070
rect 15180 20030 15220 20070
rect 15580 20030 15620 20070
rect 380 19630 420 19670
rect 780 19630 820 19670
rect 1180 19630 1220 19670
rect 1580 19630 1620 19670
rect 1980 19630 2020 19670
rect 2380 19630 2420 19670
rect 2780 19630 2820 19670
rect 3180 19630 3220 19670
rect 3580 19630 3620 19670
rect 3980 19630 4020 19670
rect 4380 19630 4420 19670
rect 4780 19630 4820 19670
rect 5180 19630 5220 19670
rect 5580 19630 5620 19670
rect 5980 19630 6020 19670
rect 6380 19630 6420 19670
rect 6780 19630 6820 19670
rect 7180 19630 7220 19670
rect 7580 19630 7620 19670
rect 7980 19630 8020 19670
rect 8380 19630 8420 19670
rect 8780 19630 8820 19670
rect 9180 19630 9220 19670
rect 9580 19630 9620 19670
rect 9980 19630 10020 19670
rect 10380 19630 10420 19670
rect 10780 19630 10820 19670
rect 11180 19630 11220 19670
rect 11580 19630 11620 19670
rect 11980 19630 12020 19670
rect 12380 19630 12420 19670
rect 12780 19630 12820 19670
rect 13180 19630 13220 19670
rect 13580 19630 13620 19670
rect 13980 19630 14020 19670
rect 14380 19630 14420 19670
rect 14780 19630 14820 19670
rect 15180 19630 15220 19670
rect 15580 19630 15620 19670
rect 380 19230 420 19270
rect 780 19230 820 19270
rect 1180 19230 1220 19270
rect 1580 19230 1620 19270
rect 1980 19230 2020 19270
rect 2380 19230 2420 19270
rect 2780 19230 2820 19270
rect 3180 19230 3220 19270
rect 3580 19230 3620 19270
rect 3980 19230 4020 19270
rect 4380 19230 4420 19270
rect 4780 19230 4820 19270
rect 5180 19230 5220 19270
rect 5580 19230 5620 19270
rect 5980 19230 6020 19270
rect 6380 19230 6420 19270
rect 6780 19230 6820 19270
rect 7180 19230 7220 19270
rect 7580 19230 7620 19270
rect 7980 19230 8020 19270
rect 8380 19230 8420 19270
rect 8780 19230 8820 19270
rect 9180 19230 9220 19270
rect 9580 19230 9620 19270
rect 9980 19230 10020 19270
rect 10380 19230 10420 19270
rect 10780 19230 10820 19270
rect 11180 19230 11220 19270
rect 11580 19230 11620 19270
rect 11980 19230 12020 19270
rect 12380 19230 12420 19270
rect 12780 19230 12820 19270
rect 13180 19230 13220 19270
rect 13580 19230 13620 19270
rect 13980 19230 14020 19270
rect 14380 19230 14420 19270
rect 14780 19230 14820 19270
rect 15180 19230 15220 19270
rect 15580 19230 15620 19270
rect 380 17730 420 17770
rect 780 17730 820 17770
rect 1180 17730 1220 17770
rect 1580 17730 1620 17770
rect 1980 17730 2020 17770
rect 2380 17730 2420 17770
rect 2780 17730 2820 17770
rect 3180 17730 3220 17770
rect 3580 17730 3620 17770
rect 3980 17730 4020 17770
rect 4380 17730 4420 17770
rect 4780 17730 4820 17770
rect 5180 17730 5220 17770
rect 5580 17730 5620 17770
rect 5980 17730 6020 17770
rect 6380 17730 6420 17770
rect 6780 17730 6820 17770
rect 7180 17730 7220 17770
rect 7580 17730 7620 17770
rect 7980 17730 8020 17770
rect 8380 17730 8420 17770
rect 8780 17730 8820 17770
rect 9180 17730 9220 17770
rect 9580 17730 9620 17770
rect 9980 17730 10020 17770
rect 10380 17730 10420 17770
rect 10780 17730 10820 17770
rect 11180 17730 11220 17770
rect 11580 17730 11620 17770
rect 11980 17730 12020 17770
rect 12380 17730 12420 17770
rect 12780 17730 12820 17770
rect 13180 17730 13220 17770
rect 13580 17730 13620 17770
rect 13980 17730 14020 17770
rect 14380 17730 14420 17770
rect 14780 17730 14820 17770
rect 15180 17730 15220 17770
rect 15580 17730 15620 17770
rect 380 17330 420 17370
rect 780 17330 820 17370
rect 1180 17330 1220 17370
rect 1580 17330 1620 17370
rect 1980 17330 2020 17370
rect 2380 17330 2420 17370
rect 2780 17330 2820 17370
rect 3180 17330 3220 17370
rect 3580 17330 3620 17370
rect 3980 17330 4020 17370
rect 4380 17330 4420 17370
rect 4780 17330 4820 17370
rect 5180 17330 5220 17370
rect 5580 17330 5620 17370
rect 5980 17330 6020 17370
rect 6380 17330 6420 17370
rect 6780 17330 6820 17370
rect 7180 17330 7220 17370
rect 7580 17330 7620 17370
rect 7980 17330 8020 17370
rect 8380 17330 8420 17370
rect 8780 17330 8820 17370
rect 9180 17330 9220 17370
rect 9580 17330 9620 17370
rect 9980 17330 10020 17370
rect 10380 17330 10420 17370
rect 10780 17330 10820 17370
rect 11180 17330 11220 17370
rect 11580 17330 11620 17370
rect 11980 17330 12020 17370
rect 12380 17330 12420 17370
rect 12780 17330 12820 17370
rect 13180 17330 13220 17370
rect 13580 17330 13620 17370
rect 13980 17330 14020 17370
rect 14380 17330 14420 17370
rect 14780 17330 14820 17370
rect 15180 17330 15220 17370
rect 15580 17330 15620 17370
rect 380 16930 420 16970
rect 780 16930 820 16970
rect 1180 16930 1220 16970
rect 1580 16930 1620 16970
rect 1980 16930 2020 16970
rect 2380 16930 2420 16970
rect 2780 16930 2820 16970
rect 3180 16930 3220 16970
rect 3580 16930 3620 16970
rect 3980 16930 4020 16970
rect 4380 16930 4420 16970
rect 4780 16930 4820 16970
rect 5180 16930 5220 16970
rect 5580 16930 5620 16970
rect 5980 16930 6020 16970
rect 6380 16930 6420 16970
rect 6780 16930 6820 16970
rect 7180 16930 7220 16970
rect 7580 16930 7620 16970
rect 7980 16930 8020 16970
rect 8380 16930 8420 16970
rect 8780 16930 8820 16970
rect 9180 16930 9220 16970
rect 9580 16930 9620 16970
rect 9980 16930 10020 16970
rect 10380 16930 10420 16970
rect 10780 16930 10820 16970
rect 11180 16930 11220 16970
rect 11580 16930 11620 16970
rect 11980 16930 12020 16970
rect 12380 16930 12420 16970
rect 12780 16930 12820 16970
rect 13180 16930 13220 16970
rect 13580 16930 13620 16970
rect 13980 16930 14020 16970
rect 14380 16930 14420 16970
rect 14780 16930 14820 16970
rect 15180 16930 15220 16970
rect 15580 16930 15620 16970
rect 380 16530 420 16570
rect 780 16530 820 16570
rect 1180 16530 1220 16570
rect 1580 16530 1620 16570
rect 1980 16530 2020 16570
rect 2380 16530 2420 16570
rect 2780 16530 2820 16570
rect 3180 16530 3220 16570
rect 3580 16530 3620 16570
rect 3980 16530 4020 16570
rect 4380 16530 4420 16570
rect 4780 16530 4820 16570
rect 5180 16530 5220 16570
rect 5580 16530 5620 16570
rect 5980 16530 6020 16570
rect 6380 16530 6420 16570
rect 6780 16530 6820 16570
rect 7180 16530 7220 16570
rect 7580 16530 7620 16570
rect 7980 16530 8020 16570
rect 8380 16530 8420 16570
rect 8780 16530 8820 16570
rect 9180 16530 9220 16570
rect 9580 16530 9620 16570
rect 9980 16530 10020 16570
rect 10380 16530 10420 16570
rect 10780 16530 10820 16570
rect 11180 16530 11220 16570
rect 11580 16530 11620 16570
rect 11980 16530 12020 16570
rect 12380 16530 12420 16570
rect 12780 16530 12820 16570
rect 13180 16530 13220 16570
rect 13580 16530 13620 16570
rect 13980 16530 14020 16570
rect 14380 16530 14420 16570
rect 14780 16530 14820 16570
rect 15180 16530 15220 16570
rect 15580 16530 15620 16570
rect 380 16130 420 16170
rect 780 16130 820 16170
rect 1180 16130 1220 16170
rect 1580 16130 1620 16170
rect 1980 16130 2020 16170
rect 2380 16130 2420 16170
rect 2780 16130 2820 16170
rect 3180 16130 3220 16170
rect 3580 16130 3620 16170
rect 3980 16130 4020 16170
rect 4380 16130 4420 16170
rect 4780 16130 4820 16170
rect 5180 16130 5220 16170
rect 5580 16130 5620 16170
rect 5980 16130 6020 16170
rect 6380 16130 6420 16170
rect 6780 16130 6820 16170
rect 7180 16130 7220 16170
rect 7580 16130 7620 16170
rect 7980 16130 8020 16170
rect 8380 16130 8420 16170
rect 8780 16130 8820 16170
rect 9180 16130 9220 16170
rect 9580 16130 9620 16170
rect 9980 16130 10020 16170
rect 10380 16130 10420 16170
rect 10780 16130 10820 16170
rect 11180 16130 11220 16170
rect 11580 16130 11620 16170
rect 11980 16130 12020 16170
rect 12380 16130 12420 16170
rect 12780 16130 12820 16170
rect 13180 16130 13220 16170
rect 13580 16130 13620 16170
rect 13980 16130 14020 16170
rect 14380 16130 14420 16170
rect 14780 16130 14820 16170
rect 15180 16130 15220 16170
rect 15580 16130 15620 16170
rect 380 15730 420 15770
rect 780 15730 820 15770
rect 1180 15730 1220 15770
rect 1580 15730 1620 15770
rect 1980 15730 2020 15770
rect 2380 15730 2420 15770
rect 2780 15730 2820 15770
rect 3180 15730 3220 15770
rect 3580 15730 3620 15770
rect 3980 15730 4020 15770
rect 4380 15730 4420 15770
rect 4780 15730 4820 15770
rect 5180 15730 5220 15770
rect 5580 15730 5620 15770
rect 5980 15730 6020 15770
rect 6380 15730 6420 15770
rect 6780 15730 6820 15770
rect 7180 15730 7220 15770
rect 7580 15730 7620 15770
rect 7980 15730 8020 15770
rect 8380 15730 8420 15770
rect 8780 15730 8820 15770
rect 9180 15730 9220 15770
rect 9580 15730 9620 15770
rect 9980 15730 10020 15770
rect 10380 15730 10420 15770
rect 10780 15730 10820 15770
rect 11180 15730 11220 15770
rect 11580 15730 11620 15770
rect 11980 15730 12020 15770
rect 12380 15730 12420 15770
rect 12780 15730 12820 15770
rect 13180 15730 13220 15770
rect 13580 15730 13620 15770
rect 13980 15730 14020 15770
rect 14380 15730 14420 15770
rect 14780 15730 14820 15770
rect 15180 15730 15220 15770
rect 15580 15730 15620 15770
rect 380 15330 420 15370
rect 780 15330 820 15370
rect 1180 15330 1220 15370
rect 1580 15330 1620 15370
rect 1980 15330 2020 15370
rect 2380 15330 2420 15370
rect 2780 15330 2820 15370
rect 3180 15330 3220 15370
rect 3580 15330 3620 15370
rect 3980 15330 4020 15370
rect 4380 15330 4420 15370
rect 4780 15330 4820 15370
rect 5180 15330 5220 15370
rect 5580 15330 5620 15370
rect 5980 15330 6020 15370
rect 6380 15330 6420 15370
rect 6780 15330 6820 15370
rect 7180 15330 7220 15370
rect 7580 15330 7620 15370
rect 7980 15330 8020 15370
rect 8380 15330 8420 15370
rect 8780 15330 8820 15370
rect 9180 15330 9220 15370
rect 9580 15330 9620 15370
rect 9980 15330 10020 15370
rect 10380 15330 10420 15370
rect 10780 15330 10820 15370
rect 11180 15330 11220 15370
rect 11580 15330 11620 15370
rect 11980 15330 12020 15370
rect 12380 15330 12420 15370
rect 12780 15330 12820 15370
rect 13180 15330 13220 15370
rect 13580 15330 13620 15370
rect 13980 15330 14020 15370
rect 14380 15330 14420 15370
rect 14780 15330 14820 15370
rect 15180 15330 15220 15370
rect 15580 15330 15620 15370
rect 380 14930 420 14970
rect 780 14930 820 14970
rect 1180 14930 1220 14970
rect 1580 14930 1620 14970
rect 1980 14930 2020 14970
rect 2380 14930 2420 14970
rect 2780 14930 2820 14970
rect 3180 14930 3220 14970
rect 3580 14930 3620 14970
rect 3980 14930 4020 14970
rect 4380 14930 4420 14970
rect 4780 14930 4820 14970
rect 5180 14930 5220 14970
rect 5580 14930 5620 14970
rect 5980 14930 6020 14970
rect 6380 14930 6420 14970
rect 6780 14930 6820 14970
rect 7180 14930 7220 14970
rect 7580 14930 7620 14970
rect 7980 14930 8020 14970
rect 8380 14930 8420 14970
rect 8780 14930 8820 14970
rect 9180 14930 9220 14970
rect 9580 14930 9620 14970
rect 9980 14930 10020 14970
rect 10380 14930 10420 14970
rect 10780 14930 10820 14970
rect 11180 14930 11220 14970
rect 11580 14930 11620 14970
rect 11980 14930 12020 14970
rect 12380 14930 12420 14970
rect 12780 14930 12820 14970
rect 13180 14930 13220 14970
rect 13580 14930 13620 14970
rect 13980 14930 14020 14970
rect 14380 14930 14420 14970
rect 14780 14930 14820 14970
rect 15180 14930 15220 14970
rect 15580 14930 15620 14970
rect 380 14530 420 14570
rect 780 14530 820 14570
rect 1180 14530 1220 14570
rect 1580 14530 1620 14570
rect 1980 14530 2020 14570
rect 2380 14530 2420 14570
rect 2780 14530 2820 14570
rect 3180 14530 3220 14570
rect 3580 14530 3620 14570
rect 3980 14530 4020 14570
rect 4380 14530 4420 14570
rect 4780 14530 4820 14570
rect 5180 14530 5220 14570
rect 5580 14530 5620 14570
rect 5980 14530 6020 14570
rect 6380 14530 6420 14570
rect 6780 14530 6820 14570
rect 7180 14530 7220 14570
rect 7580 14530 7620 14570
rect 7980 14530 8020 14570
rect 8380 14530 8420 14570
rect 8780 14530 8820 14570
rect 9180 14530 9220 14570
rect 9580 14530 9620 14570
rect 9980 14530 10020 14570
rect 10380 14530 10420 14570
rect 10780 14530 10820 14570
rect 11180 14530 11220 14570
rect 11580 14530 11620 14570
rect 11980 14530 12020 14570
rect 12380 14530 12420 14570
rect 12780 14530 12820 14570
rect 13180 14530 13220 14570
rect 13580 14530 13620 14570
rect 13980 14530 14020 14570
rect 14380 14530 14420 14570
rect 14780 14530 14820 14570
rect 15180 14530 15220 14570
rect 15580 14530 15620 14570
rect 380 14130 420 14170
rect 780 14130 820 14170
rect 1180 14130 1220 14170
rect 1580 14130 1620 14170
rect 1980 14130 2020 14170
rect 2380 14130 2420 14170
rect 2780 14130 2820 14170
rect 3180 14130 3220 14170
rect 3580 14130 3620 14170
rect 3980 14130 4020 14170
rect 4380 14130 4420 14170
rect 4780 14130 4820 14170
rect 5180 14130 5220 14170
rect 5580 14130 5620 14170
rect 5980 14130 6020 14170
rect 6380 14130 6420 14170
rect 6780 14130 6820 14170
rect 7180 14130 7220 14170
rect 7580 14130 7620 14170
rect 7980 14130 8020 14170
rect 8380 14130 8420 14170
rect 8780 14130 8820 14170
rect 9180 14130 9220 14170
rect 9580 14130 9620 14170
rect 9980 14130 10020 14170
rect 10380 14130 10420 14170
rect 10780 14130 10820 14170
rect 11180 14130 11220 14170
rect 11580 14130 11620 14170
rect 11980 14130 12020 14170
rect 12380 14130 12420 14170
rect 12780 14130 12820 14170
rect 13180 14130 13220 14170
rect 13580 14130 13620 14170
rect 13980 14130 14020 14170
rect 14380 14130 14420 14170
rect 14780 14130 14820 14170
rect 15180 14130 15220 14170
rect 15580 14130 15620 14170
rect 380 13730 420 13770
rect 780 13730 820 13770
rect 1180 13730 1220 13770
rect 1580 13730 1620 13770
rect 1980 13730 2020 13770
rect 2380 13730 2420 13770
rect 2780 13730 2820 13770
rect 3180 13730 3220 13770
rect 3580 13730 3620 13770
rect 3980 13730 4020 13770
rect 4380 13730 4420 13770
rect 4780 13730 4820 13770
rect 5180 13730 5220 13770
rect 5580 13730 5620 13770
rect 5980 13730 6020 13770
rect 6380 13730 6420 13770
rect 6780 13730 6820 13770
rect 7180 13730 7220 13770
rect 7580 13730 7620 13770
rect 7980 13730 8020 13770
rect 8380 13730 8420 13770
rect 8780 13730 8820 13770
rect 9180 13730 9220 13770
rect 9580 13730 9620 13770
rect 9980 13730 10020 13770
rect 10380 13730 10420 13770
rect 10780 13730 10820 13770
rect 11180 13730 11220 13770
rect 11580 13730 11620 13770
rect 11980 13730 12020 13770
rect 12380 13730 12420 13770
rect 12780 13730 12820 13770
rect 13180 13730 13220 13770
rect 13580 13730 13620 13770
rect 13980 13730 14020 13770
rect 14380 13730 14420 13770
rect 14780 13730 14820 13770
rect 15180 13730 15220 13770
rect 15580 13730 15620 13770
rect 380 11430 420 11470
rect 780 11430 820 11470
rect 1180 11430 1220 11470
rect 1580 11430 1620 11470
rect 1980 11430 2020 11470
rect 2380 11430 2420 11470
rect 2780 11430 2820 11470
rect 3180 11430 3220 11470
rect 3580 11430 3620 11470
rect 3980 11430 4020 11470
rect 4380 11430 4420 11470
rect 4780 11430 4820 11470
rect 5180 11430 5220 11470
rect 5580 11430 5620 11470
rect 5980 11430 6020 11470
rect 6380 11430 6420 11470
rect 6780 11430 6820 11470
rect 7180 11430 7220 11470
rect 7580 11430 7620 11470
rect 7980 11430 8020 11470
rect 8380 11430 8420 11470
rect 8780 11430 8820 11470
rect 9180 11430 9220 11470
rect 9580 11430 9620 11470
rect 9980 11430 10020 11470
rect 10380 11430 10420 11470
rect 10780 11430 10820 11470
rect 11180 11430 11220 11470
rect 11580 11430 11620 11470
rect 11980 11430 12020 11470
rect 12380 11430 12420 11470
rect 12780 11430 12820 11470
rect 13180 11430 13220 11470
rect 13580 11430 13620 11470
rect 13980 11430 14020 11470
rect 14380 11430 14420 11470
rect 14780 11430 14820 11470
rect 15180 11430 15220 11470
rect 15580 11430 15620 11470
rect 380 11030 420 11070
rect 780 11030 820 11070
rect 1180 11030 1220 11070
rect 1580 11030 1620 11070
rect 1980 11030 2020 11070
rect 2380 11030 2420 11070
rect 2780 11030 2820 11070
rect 3180 11030 3220 11070
rect 3580 11030 3620 11070
rect 3980 11030 4020 11070
rect 4380 11030 4420 11070
rect 4780 11030 4820 11070
rect 5180 11030 5220 11070
rect 5580 11030 5620 11070
rect 5980 11030 6020 11070
rect 6380 11030 6420 11070
rect 6780 11030 6820 11070
rect 7180 11030 7220 11070
rect 7580 11030 7620 11070
rect 7980 11030 8020 11070
rect 8380 11030 8420 11070
rect 8780 11030 8820 11070
rect 9180 11030 9220 11070
rect 9580 11030 9620 11070
rect 9980 11030 10020 11070
rect 10380 11030 10420 11070
rect 10780 11030 10820 11070
rect 11180 11030 11220 11070
rect 11580 11030 11620 11070
rect 11980 11030 12020 11070
rect 12380 11030 12420 11070
rect 12780 11030 12820 11070
rect 13180 11030 13220 11070
rect 13580 11030 13620 11070
rect 13980 11030 14020 11070
rect 14380 11030 14420 11070
rect 14780 11030 14820 11070
rect 15180 11030 15220 11070
rect 15580 11030 15620 11070
rect 380 10630 420 10670
rect 780 10630 820 10670
rect 1180 10630 1220 10670
rect 1580 10630 1620 10670
rect 1980 10630 2020 10670
rect 2380 10630 2420 10670
rect 2780 10630 2820 10670
rect 3180 10630 3220 10670
rect 3580 10630 3620 10670
rect 3980 10630 4020 10670
rect 4380 10630 4420 10670
rect 4780 10630 4820 10670
rect 5180 10630 5220 10670
rect 5580 10630 5620 10670
rect 5980 10630 6020 10670
rect 6380 10630 6420 10670
rect 6780 10630 6820 10670
rect 7180 10630 7220 10670
rect 7580 10630 7620 10670
rect 7980 10630 8020 10670
rect 8380 10630 8420 10670
rect 8780 10630 8820 10670
rect 9180 10630 9220 10670
rect 9580 10630 9620 10670
rect 9980 10630 10020 10670
rect 10380 10630 10420 10670
rect 10780 10630 10820 10670
rect 11180 10630 11220 10670
rect 11580 10630 11620 10670
rect 11980 10630 12020 10670
rect 12380 10630 12420 10670
rect 12780 10630 12820 10670
rect 13180 10630 13220 10670
rect 13580 10630 13620 10670
rect 13980 10630 14020 10670
rect 14380 10630 14420 10670
rect 14780 10630 14820 10670
rect 15180 10630 15220 10670
rect 15580 10630 15620 10670
rect 380 10230 420 10270
rect 780 10230 820 10270
rect 1180 10230 1220 10270
rect 1580 10230 1620 10270
rect 1980 10230 2020 10270
rect 2380 10230 2420 10270
rect 2780 10230 2820 10270
rect 3180 10230 3220 10270
rect 3580 10230 3620 10270
rect 3980 10230 4020 10270
rect 4380 10230 4420 10270
rect 4780 10230 4820 10270
rect 5180 10230 5220 10270
rect 5580 10230 5620 10270
rect 5980 10230 6020 10270
rect 6380 10230 6420 10270
rect 6780 10230 6820 10270
rect 7180 10230 7220 10270
rect 7580 10230 7620 10270
rect 7980 10230 8020 10270
rect 8380 10230 8420 10270
rect 8780 10230 8820 10270
rect 9180 10230 9220 10270
rect 9580 10230 9620 10270
rect 9980 10230 10020 10270
rect 10380 10230 10420 10270
rect 10780 10230 10820 10270
rect 11180 10230 11220 10270
rect 11580 10230 11620 10270
rect 11980 10230 12020 10270
rect 12380 10230 12420 10270
rect 12780 10230 12820 10270
rect 13180 10230 13220 10270
rect 13580 10230 13620 10270
rect 13980 10230 14020 10270
rect 14380 10230 14420 10270
rect 14780 10230 14820 10270
rect 15180 10230 15220 10270
rect 15580 10230 15620 10270
rect 380 9830 420 9870
rect 780 9830 820 9870
rect 1180 9830 1220 9870
rect 1580 9830 1620 9870
rect 1980 9830 2020 9870
rect 2380 9830 2420 9870
rect 2780 9830 2820 9870
rect 3180 9830 3220 9870
rect 3580 9830 3620 9870
rect 3980 9830 4020 9870
rect 4380 9830 4420 9870
rect 4780 9830 4820 9870
rect 5180 9830 5220 9870
rect 5580 9830 5620 9870
rect 5980 9830 6020 9870
rect 6380 9830 6420 9870
rect 6780 9830 6820 9870
rect 7180 9830 7220 9870
rect 7580 9830 7620 9870
rect 7980 9830 8020 9870
rect 8380 9830 8420 9870
rect 8780 9830 8820 9870
rect 9180 9830 9220 9870
rect 9580 9830 9620 9870
rect 9980 9830 10020 9870
rect 10380 9830 10420 9870
rect 10780 9830 10820 9870
rect 11180 9830 11220 9870
rect 11580 9830 11620 9870
rect 11980 9830 12020 9870
rect 12380 9830 12420 9870
rect 12780 9830 12820 9870
rect 13180 9830 13220 9870
rect 13580 9830 13620 9870
rect 13980 9830 14020 9870
rect 14380 9830 14420 9870
rect 14780 9830 14820 9870
rect 15180 9830 15220 9870
rect 15580 9830 15620 9870
rect 380 9430 420 9470
rect 780 9430 820 9470
rect 1180 9430 1220 9470
rect 1580 9430 1620 9470
rect 1980 9430 2020 9470
rect 2380 9430 2420 9470
rect 2780 9430 2820 9470
rect 3180 9430 3220 9470
rect 3580 9430 3620 9470
rect 3980 9430 4020 9470
rect 4380 9430 4420 9470
rect 4780 9430 4820 9470
rect 5180 9430 5220 9470
rect 5580 9430 5620 9470
rect 5980 9430 6020 9470
rect 6380 9430 6420 9470
rect 6780 9430 6820 9470
rect 7180 9430 7220 9470
rect 7580 9430 7620 9470
rect 7980 9430 8020 9470
rect 8380 9430 8420 9470
rect 8780 9430 8820 9470
rect 9180 9430 9220 9470
rect 9580 9430 9620 9470
rect 9980 9430 10020 9470
rect 10380 9430 10420 9470
rect 10780 9430 10820 9470
rect 11180 9430 11220 9470
rect 11580 9430 11620 9470
rect 11980 9430 12020 9470
rect 12380 9430 12420 9470
rect 12780 9430 12820 9470
rect 13180 9430 13220 9470
rect 13580 9430 13620 9470
rect 13980 9430 14020 9470
rect 14380 9430 14420 9470
rect 14780 9430 14820 9470
rect 15180 9430 15220 9470
rect 15580 9430 15620 9470
rect 380 9030 420 9070
rect 780 9030 820 9070
rect 1180 9030 1220 9070
rect 1580 9030 1620 9070
rect 1980 9030 2020 9070
rect 2380 9030 2420 9070
rect 2780 9030 2820 9070
rect 3180 9030 3220 9070
rect 3580 9030 3620 9070
rect 3980 9030 4020 9070
rect 4380 9030 4420 9070
rect 4780 9030 4820 9070
rect 5180 9030 5220 9070
rect 5580 9030 5620 9070
rect 5980 9030 6020 9070
rect 6380 9030 6420 9070
rect 6780 9030 6820 9070
rect 7180 9030 7220 9070
rect 7580 9030 7620 9070
rect 7980 9030 8020 9070
rect 8380 9030 8420 9070
rect 8780 9030 8820 9070
rect 9180 9030 9220 9070
rect 9580 9030 9620 9070
rect 9980 9030 10020 9070
rect 10380 9030 10420 9070
rect 10780 9030 10820 9070
rect 11180 9030 11220 9070
rect 11580 9030 11620 9070
rect 11980 9030 12020 9070
rect 12380 9030 12420 9070
rect 12780 9030 12820 9070
rect 13180 9030 13220 9070
rect 13580 9030 13620 9070
rect 13980 9030 14020 9070
rect 14380 9030 14420 9070
rect 14780 9030 14820 9070
rect 15180 9030 15220 9070
rect 15580 9030 15620 9070
rect 380 8630 420 8670
rect 780 8630 820 8670
rect 1180 8630 1220 8670
rect 1580 8630 1620 8670
rect 1980 8630 2020 8670
rect 2380 8630 2420 8670
rect 2780 8630 2820 8670
rect 3180 8630 3220 8670
rect 3580 8630 3620 8670
rect 3980 8630 4020 8670
rect 4380 8630 4420 8670
rect 4780 8630 4820 8670
rect 5180 8630 5220 8670
rect 5580 8630 5620 8670
rect 5980 8630 6020 8670
rect 6380 8630 6420 8670
rect 6780 8630 6820 8670
rect 7180 8630 7220 8670
rect 7580 8630 7620 8670
rect 7980 8630 8020 8670
rect 8380 8630 8420 8670
rect 8780 8630 8820 8670
rect 9180 8630 9220 8670
rect 9580 8630 9620 8670
rect 9980 8630 10020 8670
rect 10380 8630 10420 8670
rect 10780 8630 10820 8670
rect 11180 8630 11220 8670
rect 11580 8630 11620 8670
rect 11980 8630 12020 8670
rect 12380 8630 12420 8670
rect 12780 8630 12820 8670
rect 13180 8630 13220 8670
rect 13580 8630 13620 8670
rect 13980 8630 14020 8670
rect 14380 8630 14420 8670
rect 14780 8630 14820 8670
rect 15180 8630 15220 8670
rect 15580 8630 15620 8670
rect 380 8230 420 8270
rect 780 8230 820 8270
rect 1180 8230 1220 8270
rect 1580 8230 1620 8270
rect 1980 8230 2020 8270
rect 2380 8230 2420 8270
rect 2780 8230 2820 8270
rect 3180 8230 3220 8270
rect 3580 8230 3620 8270
rect 3980 8230 4020 8270
rect 4380 8230 4420 8270
rect 4780 8230 4820 8270
rect 5180 8230 5220 8270
rect 5580 8230 5620 8270
rect 5980 8230 6020 8270
rect 6380 8230 6420 8270
rect 6780 8230 6820 8270
rect 7180 8230 7220 8270
rect 7580 8230 7620 8270
rect 7980 8230 8020 8270
rect 8380 8230 8420 8270
rect 8780 8230 8820 8270
rect 9180 8230 9220 8270
rect 9580 8230 9620 8270
rect 9980 8230 10020 8270
rect 10380 8230 10420 8270
rect 10780 8230 10820 8270
rect 11180 8230 11220 8270
rect 11580 8230 11620 8270
rect 11980 8230 12020 8270
rect 12380 8230 12420 8270
rect 12780 8230 12820 8270
rect 13180 8230 13220 8270
rect 13580 8230 13620 8270
rect 13980 8230 14020 8270
rect 14380 8230 14420 8270
rect 14780 8230 14820 8270
rect 15180 8230 15220 8270
rect 15580 8230 15620 8270
rect 380 7830 420 7870
rect 780 7830 820 7870
rect 1180 7830 1220 7870
rect 1580 7830 1620 7870
rect 1980 7830 2020 7870
rect 2380 7830 2420 7870
rect 2780 7830 2820 7870
rect 3180 7830 3220 7870
rect 3580 7830 3620 7870
rect 3980 7830 4020 7870
rect 4380 7830 4420 7870
rect 4780 7830 4820 7870
rect 5180 7830 5220 7870
rect 5580 7830 5620 7870
rect 5980 7830 6020 7870
rect 6380 7830 6420 7870
rect 6780 7830 6820 7870
rect 7180 7830 7220 7870
rect 7580 7830 7620 7870
rect 7980 7830 8020 7870
rect 8380 7830 8420 7870
rect 8780 7830 8820 7870
rect 9180 7830 9220 7870
rect 9580 7830 9620 7870
rect 9980 7830 10020 7870
rect 10380 7830 10420 7870
rect 10780 7830 10820 7870
rect 11180 7830 11220 7870
rect 11580 7830 11620 7870
rect 11980 7830 12020 7870
rect 12380 7830 12420 7870
rect 12780 7830 12820 7870
rect 13180 7830 13220 7870
rect 13580 7830 13620 7870
rect 13980 7830 14020 7870
rect 14380 7830 14420 7870
rect 14780 7830 14820 7870
rect 15180 7830 15220 7870
rect 15580 7830 15620 7870
rect 380 7430 420 7470
rect 780 7430 820 7470
rect 1180 7430 1220 7470
rect 1580 7430 1620 7470
rect 1980 7430 2020 7470
rect 2380 7430 2420 7470
rect 2780 7430 2820 7470
rect 3180 7430 3220 7470
rect 3580 7430 3620 7470
rect 3980 7430 4020 7470
rect 4380 7430 4420 7470
rect 4780 7430 4820 7470
rect 5180 7430 5220 7470
rect 5580 7430 5620 7470
rect 5980 7430 6020 7470
rect 6380 7430 6420 7470
rect 6780 7430 6820 7470
rect 7180 7430 7220 7470
rect 7580 7430 7620 7470
rect 7980 7430 8020 7470
rect 8380 7430 8420 7470
rect 8780 7430 8820 7470
rect 9180 7430 9220 7470
rect 9580 7430 9620 7470
rect 9980 7430 10020 7470
rect 10380 7430 10420 7470
rect 10780 7430 10820 7470
rect 11180 7430 11220 7470
rect 11580 7430 11620 7470
rect 11980 7430 12020 7470
rect 12380 7430 12420 7470
rect 12780 7430 12820 7470
rect 13180 7430 13220 7470
rect 13580 7430 13620 7470
rect 13980 7430 14020 7470
rect 14380 7430 14420 7470
rect 14780 7430 14820 7470
rect 15180 7430 15220 7470
rect 15580 7430 15620 7470
rect 380 5930 420 5970
rect 780 5930 820 5970
rect 1180 5930 1220 5970
rect 1580 5930 1620 5970
rect 1980 5930 2020 5970
rect 2380 5930 2420 5970
rect 2780 5930 2820 5970
rect 3180 5930 3220 5970
rect 3580 5930 3620 5970
rect 3980 5930 4020 5970
rect 4380 5930 4420 5970
rect 4780 5930 4820 5970
rect 5180 5930 5220 5970
rect 5580 5930 5620 5970
rect 5980 5930 6020 5970
rect 6380 5930 6420 5970
rect 6780 5930 6820 5970
rect 7180 5930 7220 5970
rect 7580 5930 7620 5970
rect 7980 5930 8020 5970
rect 8380 5930 8420 5970
rect 8780 5930 8820 5970
rect 9180 5930 9220 5970
rect 9580 5930 9620 5970
rect 9980 5930 10020 5970
rect 10380 5930 10420 5970
rect 10780 5930 10820 5970
rect 11180 5930 11220 5970
rect 11580 5930 11620 5970
rect 11980 5930 12020 5970
rect 12380 5930 12420 5970
rect 12780 5930 12820 5970
rect 13180 5930 13220 5970
rect 13580 5930 13620 5970
rect 13980 5930 14020 5970
rect 14380 5930 14420 5970
rect 14780 5930 14820 5970
rect 15180 5930 15220 5970
rect 15580 5930 15620 5970
rect 380 5530 420 5570
rect 780 5530 820 5570
rect 1180 5530 1220 5570
rect 1580 5530 1620 5570
rect 1980 5530 2020 5570
rect 2380 5530 2420 5570
rect 2780 5530 2820 5570
rect 3180 5530 3220 5570
rect 3580 5530 3620 5570
rect 3980 5530 4020 5570
rect 4380 5530 4420 5570
rect 4780 5530 4820 5570
rect 5180 5530 5220 5570
rect 5580 5530 5620 5570
rect 5980 5530 6020 5570
rect 6380 5530 6420 5570
rect 6780 5530 6820 5570
rect 7180 5530 7220 5570
rect 7580 5530 7620 5570
rect 7980 5530 8020 5570
rect 8380 5530 8420 5570
rect 8780 5530 8820 5570
rect 9180 5530 9220 5570
rect 9580 5530 9620 5570
rect 9980 5530 10020 5570
rect 10380 5530 10420 5570
rect 10780 5530 10820 5570
rect 11180 5530 11220 5570
rect 11580 5530 11620 5570
rect 11980 5530 12020 5570
rect 12380 5530 12420 5570
rect 12780 5530 12820 5570
rect 13180 5530 13220 5570
rect 13580 5530 13620 5570
rect 13980 5530 14020 5570
rect 14380 5530 14420 5570
rect 14780 5530 14820 5570
rect 15180 5530 15220 5570
rect 15580 5530 15620 5570
rect 380 5130 420 5170
rect 780 5130 820 5170
rect 1180 5130 1220 5170
rect 1580 5130 1620 5170
rect 1980 5130 2020 5170
rect 2380 5130 2420 5170
rect 2780 5130 2820 5170
rect 3180 5130 3220 5170
rect 3580 5130 3620 5170
rect 3980 5130 4020 5170
rect 4380 5130 4420 5170
rect 4780 5130 4820 5170
rect 5180 5130 5220 5170
rect 5580 5130 5620 5170
rect 5980 5130 6020 5170
rect 6380 5130 6420 5170
rect 6780 5130 6820 5170
rect 7180 5130 7220 5170
rect 7580 5130 7620 5170
rect 7980 5130 8020 5170
rect 8380 5130 8420 5170
rect 8780 5130 8820 5170
rect 9180 5130 9220 5170
rect 9580 5130 9620 5170
rect 9980 5130 10020 5170
rect 10380 5130 10420 5170
rect 10780 5130 10820 5170
rect 11180 5130 11220 5170
rect 11580 5130 11620 5170
rect 11980 5130 12020 5170
rect 12380 5130 12420 5170
rect 12780 5130 12820 5170
rect 13180 5130 13220 5170
rect 13580 5130 13620 5170
rect 13980 5130 14020 5170
rect 14380 5130 14420 5170
rect 14780 5130 14820 5170
rect 15180 5130 15220 5170
rect 15580 5130 15620 5170
rect 380 4730 420 4770
rect 780 4730 820 4770
rect 1180 4730 1220 4770
rect 1580 4730 1620 4770
rect 1980 4730 2020 4770
rect 2380 4730 2420 4770
rect 2780 4730 2820 4770
rect 3180 4730 3220 4770
rect 3580 4730 3620 4770
rect 3980 4730 4020 4770
rect 4380 4730 4420 4770
rect 4780 4730 4820 4770
rect 5180 4730 5220 4770
rect 5580 4730 5620 4770
rect 5980 4730 6020 4770
rect 6380 4730 6420 4770
rect 6780 4730 6820 4770
rect 7180 4730 7220 4770
rect 7580 4730 7620 4770
rect 7980 4730 8020 4770
rect 8380 4730 8420 4770
rect 8780 4730 8820 4770
rect 9180 4730 9220 4770
rect 9580 4730 9620 4770
rect 9980 4730 10020 4770
rect 10380 4730 10420 4770
rect 10780 4730 10820 4770
rect 11180 4730 11220 4770
rect 11580 4730 11620 4770
rect 11980 4730 12020 4770
rect 12380 4730 12420 4770
rect 12780 4730 12820 4770
rect 13180 4730 13220 4770
rect 13580 4730 13620 4770
rect 13980 4730 14020 4770
rect 14380 4730 14420 4770
rect 14780 4730 14820 4770
rect 15180 4730 15220 4770
rect 15580 4730 15620 4770
rect 380 4330 420 4370
rect 780 4330 820 4370
rect 1180 4330 1220 4370
rect 1580 4330 1620 4370
rect 1980 4330 2020 4370
rect 2380 4330 2420 4370
rect 2780 4330 2820 4370
rect 3180 4330 3220 4370
rect 3580 4330 3620 4370
rect 3980 4330 4020 4370
rect 4380 4330 4420 4370
rect 4780 4330 4820 4370
rect 5180 4330 5220 4370
rect 5580 4330 5620 4370
rect 5980 4330 6020 4370
rect 6380 4330 6420 4370
rect 6780 4330 6820 4370
rect 7180 4330 7220 4370
rect 7580 4330 7620 4370
rect 7980 4330 8020 4370
rect 8380 4330 8420 4370
rect 8780 4330 8820 4370
rect 9180 4330 9220 4370
rect 9580 4330 9620 4370
rect 9980 4330 10020 4370
rect 10380 4330 10420 4370
rect 10780 4330 10820 4370
rect 11180 4330 11220 4370
rect 11580 4330 11620 4370
rect 11980 4330 12020 4370
rect 12380 4330 12420 4370
rect 12780 4330 12820 4370
rect 13180 4330 13220 4370
rect 13580 4330 13620 4370
rect 13980 4330 14020 4370
rect 14380 4330 14420 4370
rect 14780 4330 14820 4370
rect 15180 4330 15220 4370
rect 15580 4330 15620 4370
rect 380 3930 420 3970
rect 780 3930 820 3970
rect 1180 3930 1220 3970
rect 1580 3930 1620 3970
rect 1980 3930 2020 3970
rect 2380 3930 2420 3970
rect 2780 3930 2820 3970
rect 3180 3930 3220 3970
rect 3580 3930 3620 3970
rect 3980 3930 4020 3970
rect 4380 3930 4420 3970
rect 4780 3930 4820 3970
rect 5180 3930 5220 3970
rect 5580 3930 5620 3970
rect 5980 3930 6020 3970
rect 6380 3930 6420 3970
rect 6780 3930 6820 3970
rect 7180 3930 7220 3970
rect 7580 3930 7620 3970
rect 7980 3930 8020 3970
rect 8380 3930 8420 3970
rect 8780 3930 8820 3970
rect 9180 3930 9220 3970
rect 9580 3930 9620 3970
rect 9980 3930 10020 3970
rect 10380 3930 10420 3970
rect 10780 3930 10820 3970
rect 11180 3930 11220 3970
rect 11580 3930 11620 3970
rect 11980 3930 12020 3970
rect 12380 3930 12420 3970
rect 12780 3930 12820 3970
rect 13180 3930 13220 3970
rect 13580 3930 13620 3970
rect 13980 3930 14020 3970
rect 14380 3930 14420 3970
rect 14780 3930 14820 3970
rect 15180 3930 15220 3970
rect 15580 3930 15620 3970
rect 380 3530 420 3570
rect 780 3530 820 3570
rect 1180 3530 1220 3570
rect 1580 3530 1620 3570
rect 1980 3530 2020 3570
rect 2380 3530 2420 3570
rect 2780 3530 2820 3570
rect 3180 3530 3220 3570
rect 3580 3530 3620 3570
rect 3980 3530 4020 3570
rect 4380 3530 4420 3570
rect 4780 3530 4820 3570
rect 5180 3530 5220 3570
rect 5580 3530 5620 3570
rect 5980 3530 6020 3570
rect 6380 3530 6420 3570
rect 6780 3530 6820 3570
rect 7180 3530 7220 3570
rect 7580 3530 7620 3570
rect 7980 3530 8020 3570
rect 8380 3530 8420 3570
rect 8780 3530 8820 3570
rect 9180 3530 9220 3570
rect 9580 3530 9620 3570
rect 9980 3530 10020 3570
rect 10380 3530 10420 3570
rect 10780 3530 10820 3570
rect 11180 3530 11220 3570
rect 11580 3530 11620 3570
rect 11980 3530 12020 3570
rect 12380 3530 12420 3570
rect 12780 3530 12820 3570
rect 13180 3530 13220 3570
rect 13580 3530 13620 3570
rect 13980 3530 14020 3570
rect 14380 3530 14420 3570
rect 14780 3530 14820 3570
rect 15180 3530 15220 3570
rect 15580 3530 15620 3570
rect 380 3130 420 3170
rect 780 3130 820 3170
rect 1180 3130 1220 3170
rect 1580 3130 1620 3170
rect 1980 3130 2020 3170
rect 2380 3130 2420 3170
rect 2780 3130 2820 3170
rect 3180 3130 3220 3170
rect 3580 3130 3620 3170
rect 3980 3130 4020 3170
rect 4380 3130 4420 3170
rect 4780 3130 4820 3170
rect 5180 3130 5220 3170
rect 5580 3130 5620 3170
rect 5980 3130 6020 3170
rect 6380 3130 6420 3170
rect 6780 3130 6820 3170
rect 7180 3130 7220 3170
rect 7580 3130 7620 3170
rect 7980 3130 8020 3170
rect 8380 3130 8420 3170
rect 8780 3130 8820 3170
rect 9180 3130 9220 3170
rect 9580 3130 9620 3170
rect 9980 3130 10020 3170
rect 10380 3130 10420 3170
rect 10780 3130 10820 3170
rect 11180 3130 11220 3170
rect 11580 3130 11620 3170
rect 11980 3130 12020 3170
rect 12380 3130 12420 3170
rect 12780 3130 12820 3170
rect 13180 3130 13220 3170
rect 13580 3130 13620 3170
rect 13980 3130 14020 3170
rect 14380 3130 14420 3170
rect 14780 3130 14820 3170
rect 15180 3130 15220 3170
rect 15580 3130 15620 3170
rect 380 2730 420 2770
rect 780 2730 820 2770
rect 1180 2730 1220 2770
rect 1580 2730 1620 2770
rect 1980 2730 2020 2770
rect 2380 2730 2420 2770
rect 2780 2730 2820 2770
rect 3180 2730 3220 2770
rect 3580 2730 3620 2770
rect 3980 2730 4020 2770
rect 4380 2730 4420 2770
rect 4780 2730 4820 2770
rect 5180 2730 5220 2770
rect 5580 2730 5620 2770
rect 5980 2730 6020 2770
rect 6380 2730 6420 2770
rect 6780 2730 6820 2770
rect 7180 2730 7220 2770
rect 7580 2730 7620 2770
rect 7980 2730 8020 2770
rect 8380 2730 8420 2770
rect 8780 2730 8820 2770
rect 9180 2730 9220 2770
rect 9580 2730 9620 2770
rect 9980 2730 10020 2770
rect 10380 2730 10420 2770
rect 10780 2730 10820 2770
rect 11180 2730 11220 2770
rect 11580 2730 11620 2770
rect 11980 2730 12020 2770
rect 12380 2730 12420 2770
rect 12780 2730 12820 2770
rect 13180 2730 13220 2770
rect 13580 2730 13620 2770
rect 13980 2730 14020 2770
rect 14380 2730 14420 2770
rect 14780 2730 14820 2770
rect 15180 2730 15220 2770
rect 15580 2730 15620 2770
rect 380 2330 420 2370
rect 780 2330 820 2370
rect 1180 2330 1220 2370
rect 1580 2330 1620 2370
rect 1980 2330 2020 2370
rect 2380 2330 2420 2370
rect 2780 2330 2820 2370
rect 3180 2330 3220 2370
rect 3580 2330 3620 2370
rect 3980 2330 4020 2370
rect 4380 2330 4420 2370
rect 4780 2330 4820 2370
rect 5180 2330 5220 2370
rect 5580 2330 5620 2370
rect 5980 2330 6020 2370
rect 6380 2330 6420 2370
rect 6780 2330 6820 2370
rect 7180 2330 7220 2370
rect 7580 2330 7620 2370
rect 7980 2330 8020 2370
rect 8380 2330 8420 2370
rect 8780 2330 8820 2370
rect 9180 2330 9220 2370
rect 9580 2330 9620 2370
rect 9980 2330 10020 2370
rect 10380 2330 10420 2370
rect 10780 2330 10820 2370
rect 11180 2330 11220 2370
rect 11580 2330 11620 2370
rect 11980 2330 12020 2370
rect 12380 2330 12420 2370
rect 12780 2330 12820 2370
rect 13180 2330 13220 2370
rect 13580 2330 13620 2370
rect 13980 2330 14020 2370
rect 14380 2330 14420 2370
rect 14780 2330 14820 2370
rect 15180 2330 15220 2370
rect 15580 2330 15620 2370
rect 380 1930 420 1970
rect 780 1930 820 1970
rect 1180 1930 1220 1970
rect 1580 1930 1620 1970
rect 1980 1930 2020 1970
rect 2380 1930 2420 1970
rect 2780 1930 2820 1970
rect 3180 1930 3220 1970
rect 3580 1930 3620 1970
rect 3980 1930 4020 1970
rect 4380 1930 4420 1970
rect 4780 1930 4820 1970
rect 5180 1930 5220 1970
rect 5580 1930 5620 1970
rect 5980 1930 6020 1970
rect 6380 1930 6420 1970
rect 6780 1930 6820 1970
rect 7180 1930 7220 1970
rect 7580 1930 7620 1970
rect 7980 1930 8020 1970
rect 8380 1930 8420 1970
rect 8780 1930 8820 1970
rect 9180 1930 9220 1970
rect 9580 1930 9620 1970
rect 9980 1930 10020 1970
rect 10380 1930 10420 1970
rect 10780 1930 10820 1970
rect 11180 1930 11220 1970
rect 11580 1930 11620 1970
rect 11980 1930 12020 1970
rect 12380 1930 12420 1970
rect 12780 1930 12820 1970
rect 13180 1930 13220 1970
rect 13580 1930 13620 1970
rect 13980 1930 14020 1970
rect 14380 1930 14420 1970
rect 14780 1930 14820 1970
rect 15180 1930 15220 1970
rect 15580 1930 15620 1970
rect 1180 480 1220 520
rect 1580 480 1620 520
rect 1980 480 2020 520
rect 2380 480 2420 520
rect 2780 480 2820 520
rect 3180 480 3220 520
rect 3580 480 3620 520
rect 3980 480 4020 520
rect 4380 480 4420 520
rect 4780 480 4820 520
rect 5180 480 5220 520
rect 5580 480 5620 520
rect 5980 480 6020 520
rect 6380 480 6420 520
rect 6780 480 6820 520
rect 7180 480 7220 520
rect 7580 480 7620 520
rect 7980 480 8020 520
rect 8380 480 8420 520
rect 8780 480 8820 520
rect 9180 480 9220 520
rect 9580 480 9620 520
rect 9980 480 10020 520
rect 10380 480 10420 520
rect 10780 480 10820 520
rect 11180 480 11220 520
rect 11580 480 11620 520
rect 11980 480 12020 520
rect 12380 480 12420 520
rect 12780 480 12820 520
rect 13180 480 13220 520
rect 13580 480 13620 520
rect 13980 480 14020 520
rect 14380 480 14420 520
rect 14780 480 14820 520
rect 1180 80 1220 120
rect 1580 80 1620 120
rect 1980 80 2020 120
rect 2380 80 2420 120
rect 2780 80 2820 120
rect 3180 80 3220 120
rect 3580 80 3620 120
rect 3980 80 4020 120
rect 4380 80 4420 120
rect 4780 80 4820 120
rect 5180 80 5220 120
rect 5580 80 5620 120
rect 5980 80 6020 120
rect 6380 80 6420 120
rect 6780 80 6820 120
rect 7180 80 7220 120
rect 7580 80 7620 120
rect 7980 80 8020 120
rect 8380 80 8420 120
rect 8780 80 8820 120
rect 9180 80 9220 120
rect 9580 80 9620 120
rect 9980 80 10020 120
rect 10380 80 10420 120
rect 10780 80 10820 120
rect 11180 80 11220 120
rect 11580 80 11620 120
rect 11980 80 12020 120
rect 12380 80 12420 120
rect 12780 80 12820 120
rect 13180 80 13220 120
rect 13580 80 13620 120
rect 13980 80 14020 120
rect 14380 80 14420 120
rect 14780 80 14820 120
<< metal5 >>
rect 0 35062 16000 35600
rect 0 35040 538 35062
rect 0 35000 380 35040
rect 420 35000 538 35040
rect 0 34938 538 35000
rect 662 35040 938 35062
rect 662 35000 780 35040
rect 820 35000 938 35040
rect 662 34938 938 35000
rect 1062 35040 1338 35062
rect 1062 35000 1180 35040
rect 1220 35000 1338 35040
rect 1062 34938 1338 35000
rect 1462 35040 1738 35062
rect 1462 35000 1580 35040
rect 1620 35000 1738 35040
rect 1462 34938 1738 35000
rect 1862 35040 2138 35062
rect 1862 35000 1980 35040
rect 2020 35000 2138 35040
rect 1862 34938 2138 35000
rect 2262 35040 2538 35062
rect 2262 35000 2380 35040
rect 2420 35000 2538 35040
rect 2262 34938 2538 35000
rect 2662 35040 2938 35062
rect 2662 35000 2780 35040
rect 2820 35000 2938 35040
rect 2662 34938 2938 35000
rect 3062 35040 3338 35062
rect 3062 35000 3180 35040
rect 3220 35000 3338 35040
rect 3062 34938 3338 35000
rect 3462 35040 3738 35062
rect 3462 35000 3580 35040
rect 3620 35000 3738 35040
rect 3462 34938 3738 35000
rect 3862 35040 4138 35062
rect 3862 35000 3980 35040
rect 4020 35000 4138 35040
rect 3862 34938 4138 35000
rect 4262 35040 4538 35062
rect 4262 35000 4380 35040
rect 4420 35000 4538 35040
rect 4262 34938 4538 35000
rect 4662 35040 4938 35062
rect 4662 35000 4780 35040
rect 4820 35000 4938 35040
rect 4662 34938 4938 35000
rect 5062 35040 5338 35062
rect 5062 35000 5180 35040
rect 5220 35000 5338 35040
rect 5062 34938 5338 35000
rect 5462 35040 5738 35062
rect 5462 35000 5580 35040
rect 5620 35000 5738 35040
rect 5462 34938 5738 35000
rect 5862 35040 6138 35062
rect 5862 35000 5980 35040
rect 6020 35000 6138 35040
rect 5862 34938 6138 35000
rect 6262 35040 6538 35062
rect 6262 35000 6380 35040
rect 6420 35000 6538 35040
rect 6262 34938 6538 35000
rect 6662 35040 6938 35062
rect 6662 35000 6780 35040
rect 6820 35000 6938 35040
rect 6662 34938 6938 35000
rect 7062 35040 7338 35062
rect 7062 35000 7180 35040
rect 7220 35000 7338 35040
rect 7062 34938 7338 35000
rect 7462 35040 7738 35062
rect 7462 35000 7580 35040
rect 7620 35000 7738 35040
rect 7462 34938 7738 35000
rect 7862 35040 8138 35062
rect 7862 35000 7980 35040
rect 8020 35000 8138 35040
rect 7862 34938 8138 35000
rect 8262 35040 8538 35062
rect 8262 35000 8380 35040
rect 8420 35000 8538 35040
rect 8262 34938 8538 35000
rect 8662 35040 8938 35062
rect 8662 35000 8780 35040
rect 8820 35000 8938 35040
rect 8662 34938 8938 35000
rect 9062 35040 9338 35062
rect 9062 35000 9180 35040
rect 9220 35000 9338 35040
rect 9062 34938 9338 35000
rect 9462 35040 9738 35062
rect 9462 35000 9580 35040
rect 9620 35000 9738 35040
rect 9462 34938 9738 35000
rect 9862 35040 10138 35062
rect 9862 35000 9980 35040
rect 10020 35000 10138 35040
rect 9862 34938 10138 35000
rect 10262 35040 10538 35062
rect 10262 35000 10380 35040
rect 10420 35000 10538 35040
rect 10262 34938 10538 35000
rect 10662 35040 10938 35062
rect 10662 35000 10780 35040
rect 10820 35000 10938 35040
rect 10662 34938 10938 35000
rect 11062 35040 11338 35062
rect 11062 35000 11180 35040
rect 11220 35000 11338 35040
rect 11062 34938 11338 35000
rect 11462 35040 11738 35062
rect 11462 35000 11580 35040
rect 11620 35000 11738 35040
rect 11462 34938 11738 35000
rect 11862 35040 12138 35062
rect 11862 35000 11980 35040
rect 12020 35000 12138 35040
rect 11862 34938 12138 35000
rect 12262 35040 12538 35062
rect 12262 35000 12380 35040
rect 12420 35000 12538 35040
rect 12262 34938 12538 35000
rect 12662 35040 12938 35062
rect 12662 35000 12780 35040
rect 12820 35000 12938 35040
rect 12662 34938 12938 35000
rect 13062 35040 13338 35062
rect 13062 35000 13180 35040
rect 13220 35000 13338 35040
rect 13062 34938 13338 35000
rect 13462 35040 13738 35062
rect 13462 35000 13580 35040
rect 13620 35000 13738 35040
rect 13462 34938 13738 35000
rect 13862 35040 14138 35062
rect 13862 35000 13980 35040
rect 14020 35000 14138 35040
rect 13862 34938 14138 35000
rect 14262 35040 14538 35062
rect 14262 35000 14380 35040
rect 14420 35000 14538 35040
rect 14262 34938 14538 35000
rect 14662 35040 14938 35062
rect 14662 35000 14780 35040
rect 14820 35000 14938 35040
rect 14662 34938 14938 35000
rect 15062 35040 15338 35062
rect 15062 35000 15180 35040
rect 15220 35000 15338 35040
rect 15062 34938 15338 35000
rect 15462 35040 16000 35062
rect 15462 35000 15580 35040
rect 15620 35000 16000 35040
rect 15462 34938 16000 35000
rect 0 34662 16000 34938
rect 0 34640 538 34662
rect 0 34600 380 34640
rect 420 34600 538 34640
rect 0 34538 538 34600
rect 662 34640 938 34662
rect 662 34600 780 34640
rect 820 34600 938 34640
rect 662 34538 938 34600
rect 1062 34640 1338 34662
rect 1062 34600 1180 34640
rect 1220 34600 1338 34640
rect 1062 34538 1338 34600
rect 1462 34640 1738 34662
rect 1462 34600 1580 34640
rect 1620 34600 1738 34640
rect 1462 34538 1738 34600
rect 1862 34640 2138 34662
rect 1862 34600 1980 34640
rect 2020 34600 2138 34640
rect 1862 34538 2138 34600
rect 2262 34640 2538 34662
rect 2262 34600 2380 34640
rect 2420 34600 2538 34640
rect 2262 34538 2538 34600
rect 2662 34640 2938 34662
rect 2662 34600 2780 34640
rect 2820 34600 2938 34640
rect 2662 34538 2938 34600
rect 3062 34640 3338 34662
rect 3062 34600 3180 34640
rect 3220 34600 3338 34640
rect 3062 34538 3338 34600
rect 3462 34640 3738 34662
rect 3462 34600 3580 34640
rect 3620 34600 3738 34640
rect 3462 34538 3738 34600
rect 3862 34640 4138 34662
rect 3862 34600 3980 34640
rect 4020 34600 4138 34640
rect 3862 34538 4138 34600
rect 4262 34640 4538 34662
rect 4262 34600 4380 34640
rect 4420 34600 4538 34640
rect 4262 34538 4538 34600
rect 4662 34640 4938 34662
rect 4662 34600 4780 34640
rect 4820 34600 4938 34640
rect 4662 34538 4938 34600
rect 5062 34640 5338 34662
rect 5062 34600 5180 34640
rect 5220 34600 5338 34640
rect 5062 34538 5338 34600
rect 5462 34640 5738 34662
rect 5462 34600 5580 34640
rect 5620 34600 5738 34640
rect 5462 34538 5738 34600
rect 5862 34640 6138 34662
rect 5862 34600 5980 34640
rect 6020 34600 6138 34640
rect 5862 34538 6138 34600
rect 6262 34640 6538 34662
rect 6262 34600 6380 34640
rect 6420 34600 6538 34640
rect 6262 34538 6538 34600
rect 6662 34640 6938 34662
rect 6662 34600 6780 34640
rect 6820 34600 6938 34640
rect 6662 34538 6938 34600
rect 7062 34640 7338 34662
rect 7062 34600 7180 34640
rect 7220 34600 7338 34640
rect 7062 34538 7338 34600
rect 7462 34640 7738 34662
rect 7462 34600 7580 34640
rect 7620 34600 7738 34640
rect 7462 34538 7738 34600
rect 7862 34640 8138 34662
rect 7862 34600 7980 34640
rect 8020 34600 8138 34640
rect 7862 34538 8138 34600
rect 8262 34640 8538 34662
rect 8262 34600 8380 34640
rect 8420 34600 8538 34640
rect 8262 34538 8538 34600
rect 8662 34640 8938 34662
rect 8662 34600 8780 34640
rect 8820 34600 8938 34640
rect 8662 34538 8938 34600
rect 9062 34640 9338 34662
rect 9062 34600 9180 34640
rect 9220 34600 9338 34640
rect 9062 34538 9338 34600
rect 9462 34640 9738 34662
rect 9462 34600 9580 34640
rect 9620 34600 9738 34640
rect 9462 34538 9738 34600
rect 9862 34640 10138 34662
rect 9862 34600 9980 34640
rect 10020 34600 10138 34640
rect 9862 34538 10138 34600
rect 10262 34640 10538 34662
rect 10262 34600 10380 34640
rect 10420 34600 10538 34640
rect 10262 34538 10538 34600
rect 10662 34640 10938 34662
rect 10662 34600 10780 34640
rect 10820 34600 10938 34640
rect 10662 34538 10938 34600
rect 11062 34640 11338 34662
rect 11062 34600 11180 34640
rect 11220 34600 11338 34640
rect 11062 34538 11338 34600
rect 11462 34640 11738 34662
rect 11462 34600 11580 34640
rect 11620 34600 11738 34640
rect 11462 34538 11738 34600
rect 11862 34640 12138 34662
rect 11862 34600 11980 34640
rect 12020 34600 12138 34640
rect 11862 34538 12138 34600
rect 12262 34640 12538 34662
rect 12262 34600 12380 34640
rect 12420 34600 12538 34640
rect 12262 34538 12538 34600
rect 12662 34640 12938 34662
rect 12662 34600 12780 34640
rect 12820 34600 12938 34640
rect 12662 34538 12938 34600
rect 13062 34640 13338 34662
rect 13062 34600 13180 34640
rect 13220 34600 13338 34640
rect 13062 34538 13338 34600
rect 13462 34640 13738 34662
rect 13462 34600 13580 34640
rect 13620 34600 13738 34640
rect 13462 34538 13738 34600
rect 13862 34640 14138 34662
rect 13862 34600 13980 34640
rect 14020 34600 14138 34640
rect 13862 34538 14138 34600
rect 14262 34640 14538 34662
rect 14262 34600 14380 34640
rect 14420 34600 14538 34640
rect 14262 34538 14538 34600
rect 14662 34640 14938 34662
rect 14662 34600 14780 34640
rect 14820 34600 14938 34640
rect 14662 34538 14938 34600
rect 15062 34640 15338 34662
rect 15062 34600 15180 34640
rect 15220 34600 15338 34640
rect 15062 34538 15338 34600
rect 15462 34640 16000 34662
rect 15462 34600 15580 34640
rect 15620 34600 16000 34640
rect 15462 34538 16000 34600
rect 0 34262 16000 34538
rect 0 34240 538 34262
rect 0 34200 380 34240
rect 420 34200 538 34240
rect 0 34138 538 34200
rect 662 34240 938 34262
rect 662 34200 780 34240
rect 820 34200 938 34240
rect 662 34138 938 34200
rect 1062 34240 1338 34262
rect 1062 34200 1180 34240
rect 1220 34200 1338 34240
rect 1062 34138 1338 34200
rect 1462 34240 1738 34262
rect 1462 34200 1580 34240
rect 1620 34200 1738 34240
rect 1462 34138 1738 34200
rect 1862 34240 2138 34262
rect 1862 34200 1980 34240
rect 2020 34200 2138 34240
rect 1862 34138 2138 34200
rect 2262 34240 2538 34262
rect 2262 34200 2380 34240
rect 2420 34200 2538 34240
rect 2262 34138 2538 34200
rect 2662 34240 2938 34262
rect 2662 34200 2780 34240
rect 2820 34200 2938 34240
rect 2662 34138 2938 34200
rect 3062 34240 3338 34262
rect 3062 34200 3180 34240
rect 3220 34200 3338 34240
rect 3062 34138 3338 34200
rect 3462 34240 3738 34262
rect 3462 34200 3580 34240
rect 3620 34200 3738 34240
rect 3462 34138 3738 34200
rect 3862 34240 4138 34262
rect 3862 34200 3980 34240
rect 4020 34200 4138 34240
rect 3862 34138 4138 34200
rect 4262 34240 4538 34262
rect 4262 34200 4380 34240
rect 4420 34200 4538 34240
rect 4262 34138 4538 34200
rect 4662 34240 4938 34262
rect 4662 34200 4780 34240
rect 4820 34200 4938 34240
rect 4662 34138 4938 34200
rect 5062 34240 5338 34262
rect 5062 34200 5180 34240
rect 5220 34200 5338 34240
rect 5062 34138 5338 34200
rect 5462 34240 5738 34262
rect 5462 34200 5580 34240
rect 5620 34200 5738 34240
rect 5462 34138 5738 34200
rect 5862 34240 6138 34262
rect 5862 34200 5980 34240
rect 6020 34200 6138 34240
rect 5862 34138 6138 34200
rect 6262 34240 6538 34262
rect 6262 34200 6380 34240
rect 6420 34200 6538 34240
rect 6262 34138 6538 34200
rect 6662 34240 6938 34262
rect 6662 34200 6780 34240
rect 6820 34200 6938 34240
rect 6662 34138 6938 34200
rect 7062 34240 7338 34262
rect 7062 34200 7180 34240
rect 7220 34200 7338 34240
rect 7062 34138 7338 34200
rect 7462 34240 7738 34262
rect 7462 34200 7580 34240
rect 7620 34200 7738 34240
rect 7462 34138 7738 34200
rect 7862 34240 8138 34262
rect 7862 34200 7980 34240
rect 8020 34200 8138 34240
rect 7862 34138 8138 34200
rect 8262 34240 8538 34262
rect 8262 34200 8380 34240
rect 8420 34200 8538 34240
rect 8262 34138 8538 34200
rect 8662 34240 8938 34262
rect 8662 34200 8780 34240
rect 8820 34200 8938 34240
rect 8662 34138 8938 34200
rect 9062 34240 9338 34262
rect 9062 34200 9180 34240
rect 9220 34200 9338 34240
rect 9062 34138 9338 34200
rect 9462 34240 9738 34262
rect 9462 34200 9580 34240
rect 9620 34200 9738 34240
rect 9462 34138 9738 34200
rect 9862 34240 10138 34262
rect 9862 34200 9980 34240
rect 10020 34200 10138 34240
rect 9862 34138 10138 34200
rect 10262 34240 10538 34262
rect 10262 34200 10380 34240
rect 10420 34200 10538 34240
rect 10262 34138 10538 34200
rect 10662 34240 10938 34262
rect 10662 34200 10780 34240
rect 10820 34200 10938 34240
rect 10662 34138 10938 34200
rect 11062 34240 11338 34262
rect 11062 34200 11180 34240
rect 11220 34200 11338 34240
rect 11062 34138 11338 34200
rect 11462 34240 11738 34262
rect 11462 34200 11580 34240
rect 11620 34200 11738 34240
rect 11462 34138 11738 34200
rect 11862 34240 12138 34262
rect 11862 34200 11980 34240
rect 12020 34200 12138 34240
rect 11862 34138 12138 34200
rect 12262 34240 12538 34262
rect 12262 34200 12380 34240
rect 12420 34200 12538 34240
rect 12262 34138 12538 34200
rect 12662 34240 12938 34262
rect 12662 34200 12780 34240
rect 12820 34200 12938 34240
rect 12662 34138 12938 34200
rect 13062 34240 13338 34262
rect 13062 34200 13180 34240
rect 13220 34200 13338 34240
rect 13062 34138 13338 34200
rect 13462 34240 13738 34262
rect 13462 34200 13580 34240
rect 13620 34200 13738 34240
rect 13462 34138 13738 34200
rect 13862 34240 14138 34262
rect 13862 34200 13980 34240
rect 14020 34200 14138 34240
rect 13862 34138 14138 34200
rect 14262 34240 14538 34262
rect 14262 34200 14380 34240
rect 14420 34200 14538 34240
rect 14262 34138 14538 34200
rect 14662 34240 14938 34262
rect 14662 34200 14780 34240
rect 14820 34200 14938 34240
rect 14662 34138 14938 34200
rect 15062 34240 15338 34262
rect 15062 34200 15180 34240
rect 15220 34200 15338 34240
rect 15062 34138 15338 34200
rect 15462 34240 16000 34262
rect 15462 34200 15580 34240
rect 15620 34200 16000 34240
rect 15462 34138 16000 34200
rect 0 33862 16000 34138
rect 0 33840 538 33862
rect 0 33800 380 33840
rect 420 33800 538 33840
rect 0 33738 538 33800
rect 662 33840 938 33862
rect 662 33800 780 33840
rect 820 33800 938 33840
rect 662 33738 938 33800
rect 1062 33840 1338 33862
rect 1062 33800 1180 33840
rect 1220 33800 1338 33840
rect 1062 33738 1338 33800
rect 1462 33840 1738 33862
rect 1462 33800 1580 33840
rect 1620 33800 1738 33840
rect 1462 33738 1738 33800
rect 1862 33840 2138 33862
rect 1862 33800 1980 33840
rect 2020 33800 2138 33840
rect 1862 33738 2138 33800
rect 2262 33840 2538 33862
rect 2262 33800 2380 33840
rect 2420 33800 2538 33840
rect 2262 33738 2538 33800
rect 2662 33840 2938 33862
rect 2662 33800 2780 33840
rect 2820 33800 2938 33840
rect 2662 33738 2938 33800
rect 3062 33840 3338 33862
rect 3062 33800 3180 33840
rect 3220 33800 3338 33840
rect 3062 33738 3338 33800
rect 3462 33840 3738 33862
rect 3462 33800 3580 33840
rect 3620 33800 3738 33840
rect 3462 33738 3738 33800
rect 3862 33840 4138 33862
rect 3862 33800 3980 33840
rect 4020 33800 4138 33840
rect 3862 33738 4138 33800
rect 4262 33840 4538 33862
rect 4262 33800 4380 33840
rect 4420 33800 4538 33840
rect 4262 33738 4538 33800
rect 4662 33840 4938 33862
rect 4662 33800 4780 33840
rect 4820 33800 4938 33840
rect 4662 33738 4938 33800
rect 5062 33840 5338 33862
rect 5062 33800 5180 33840
rect 5220 33800 5338 33840
rect 5062 33738 5338 33800
rect 5462 33840 5738 33862
rect 5462 33800 5580 33840
rect 5620 33800 5738 33840
rect 5462 33738 5738 33800
rect 5862 33840 6138 33862
rect 5862 33800 5980 33840
rect 6020 33800 6138 33840
rect 5862 33738 6138 33800
rect 6262 33840 6538 33862
rect 6262 33800 6380 33840
rect 6420 33800 6538 33840
rect 6262 33738 6538 33800
rect 6662 33840 6938 33862
rect 6662 33800 6780 33840
rect 6820 33800 6938 33840
rect 6662 33738 6938 33800
rect 7062 33840 7338 33862
rect 7062 33800 7180 33840
rect 7220 33800 7338 33840
rect 7062 33738 7338 33800
rect 7462 33840 7738 33862
rect 7462 33800 7580 33840
rect 7620 33800 7738 33840
rect 7462 33738 7738 33800
rect 7862 33840 8138 33862
rect 7862 33800 7980 33840
rect 8020 33800 8138 33840
rect 7862 33738 8138 33800
rect 8262 33840 8538 33862
rect 8262 33800 8380 33840
rect 8420 33800 8538 33840
rect 8262 33738 8538 33800
rect 8662 33840 8938 33862
rect 8662 33800 8780 33840
rect 8820 33800 8938 33840
rect 8662 33738 8938 33800
rect 9062 33840 9338 33862
rect 9062 33800 9180 33840
rect 9220 33800 9338 33840
rect 9062 33738 9338 33800
rect 9462 33840 9738 33862
rect 9462 33800 9580 33840
rect 9620 33800 9738 33840
rect 9462 33738 9738 33800
rect 9862 33840 10138 33862
rect 9862 33800 9980 33840
rect 10020 33800 10138 33840
rect 9862 33738 10138 33800
rect 10262 33840 10538 33862
rect 10262 33800 10380 33840
rect 10420 33800 10538 33840
rect 10262 33738 10538 33800
rect 10662 33840 10938 33862
rect 10662 33800 10780 33840
rect 10820 33800 10938 33840
rect 10662 33738 10938 33800
rect 11062 33840 11338 33862
rect 11062 33800 11180 33840
rect 11220 33800 11338 33840
rect 11062 33738 11338 33800
rect 11462 33840 11738 33862
rect 11462 33800 11580 33840
rect 11620 33800 11738 33840
rect 11462 33738 11738 33800
rect 11862 33840 12138 33862
rect 11862 33800 11980 33840
rect 12020 33800 12138 33840
rect 11862 33738 12138 33800
rect 12262 33840 12538 33862
rect 12262 33800 12380 33840
rect 12420 33800 12538 33840
rect 12262 33738 12538 33800
rect 12662 33840 12938 33862
rect 12662 33800 12780 33840
rect 12820 33800 12938 33840
rect 12662 33738 12938 33800
rect 13062 33840 13338 33862
rect 13062 33800 13180 33840
rect 13220 33800 13338 33840
rect 13062 33738 13338 33800
rect 13462 33840 13738 33862
rect 13462 33800 13580 33840
rect 13620 33800 13738 33840
rect 13462 33738 13738 33800
rect 13862 33840 14138 33862
rect 13862 33800 13980 33840
rect 14020 33800 14138 33840
rect 13862 33738 14138 33800
rect 14262 33840 14538 33862
rect 14262 33800 14380 33840
rect 14420 33800 14538 33840
rect 14262 33738 14538 33800
rect 14662 33840 14938 33862
rect 14662 33800 14780 33840
rect 14820 33800 14938 33840
rect 14662 33738 14938 33800
rect 15062 33840 15338 33862
rect 15062 33800 15180 33840
rect 15220 33800 15338 33840
rect 15062 33738 15338 33800
rect 15462 33840 16000 33862
rect 15462 33800 15580 33840
rect 15620 33800 16000 33840
rect 15462 33738 16000 33800
rect 0 33462 16000 33738
rect 0 33440 538 33462
rect 0 33400 380 33440
rect 420 33400 538 33440
rect 0 33338 538 33400
rect 662 33440 938 33462
rect 662 33400 780 33440
rect 820 33400 938 33440
rect 662 33338 938 33400
rect 1062 33440 1338 33462
rect 1062 33400 1180 33440
rect 1220 33400 1338 33440
rect 1062 33338 1338 33400
rect 1462 33440 1738 33462
rect 1462 33400 1580 33440
rect 1620 33400 1738 33440
rect 1462 33338 1738 33400
rect 1862 33440 2138 33462
rect 1862 33400 1980 33440
rect 2020 33400 2138 33440
rect 1862 33338 2138 33400
rect 2262 33440 2538 33462
rect 2262 33400 2380 33440
rect 2420 33400 2538 33440
rect 2262 33338 2538 33400
rect 2662 33440 2938 33462
rect 2662 33400 2780 33440
rect 2820 33400 2938 33440
rect 2662 33338 2938 33400
rect 3062 33440 3338 33462
rect 3062 33400 3180 33440
rect 3220 33400 3338 33440
rect 3062 33338 3338 33400
rect 3462 33440 3738 33462
rect 3462 33400 3580 33440
rect 3620 33400 3738 33440
rect 3462 33338 3738 33400
rect 3862 33440 4138 33462
rect 3862 33400 3980 33440
rect 4020 33400 4138 33440
rect 3862 33338 4138 33400
rect 4262 33440 4538 33462
rect 4262 33400 4380 33440
rect 4420 33400 4538 33440
rect 4262 33338 4538 33400
rect 4662 33440 4938 33462
rect 4662 33400 4780 33440
rect 4820 33400 4938 33440
rect 4662 33338 4938 33400
rect 5062 33440 5338 33462
rect 5062 33400 5180 33440
rect 5220 33400 5338 33440
rect 5062 33338 5338 33400
rect 5462 33440 5738 33462
rect 5462 33400 5580 33440
rect 5620 33400 5738 33440
rect 5462 33338 5738 33400
rect 5862 33440 6138 33462
rect 5862 33400 5980 33440
rect 6020 33400 6138 33440
rect 5862 33338 6138 33400
rect 6262 33440 6538 33462
rect 6262 33400 6380 33440
rect 6420 33400 6538 33440
rect 6262 33338 6538 33400
rect 6662 33440 6938 33462
rect 6662 33400 6780 33440
rect 6820 33400 6938 33440
rect 6662 33338 6938 33400
rect 7062 33440 7338 33462
rect 7062 33400 7180 33440
rect 7220 33400 7338 33440
rect 7062 33338 7338 33400
rect 7462 33440 7738 33462
rect 7462 33400 7580 33440
rect 7620 33400 7738 33440
rect 7462 33338 7738 33400
rect 7862 33440 8138 33462
rect 7862 33400 7980 33440
rect 8020 33400 8138 33440
rect 7862 33338 8138 33400
rect 8262 33440 8538 33462
rect 8262 33400 8380 33440
rect 8420 33400 8538 33440
rect 8262 33338 8538 33400
rect 8662 33440 8938 33462
rect 8662 33400 8780 33440
rect 8820 33400 8938 33440
rect 8662 33338 8938 33400
rect 9062 33440 9338 33462
rect 9062 33400 9180 33440
rect 9220 33400 9338 33440
rect 9062 33338 9338 33400
rect 9462 33440 9738 33462
rect 9462 33400 9580 33440
rect 9620 33400 9738 33440
rect 9462 33338 9738 33400
rect 9862 33440 10138 33462
rect 9862 33400 9980 33440
rect 10020 33400 10138 33440
rect 9862 33338 10138 33400
rect 10262 33440 10538 33462
rect 10262 33400 10380 33440
rect 10420 33400 10538 33440
rect 10262 33338 10538 33400
rect 10662 33440 10938 33462
rect 10662 33400 10780 33440
rect 10820 33400 10938 33440
rect 10662 33338 10938 33400
rect 11062 33440 11338 33462
rect 11062 33400 11180 33440
rect 11220 33400 11338 33440
rect 11062 33338 11338 33400
rect 11462 33440 11738 33462
rect 11462 33400 11580 33440
rect 11620 33400 11738 33440
rect 11462 33338 11738 33400
rect 11862 33440 12138 33462
rect 11862 33400 11980 33440
rect 12020 33400 12138 33440
rect 11862 33338 12138 33400
rect 12262 33440 12538 33462
rect 12262 33400 12380 33440
rect 12420 33400 12538 33440
rect 12262 33338 12538 33400
rect 12662 33440 12938 33462
rect 12662 33400 12780 33440
rect 12820 33400 12938 33440
rect 12662 33338 12938 33400
rect 13062 33440 13338 33462
rect 13062 33400 13180 33440
rect 13220 33400 13338 33440
rect 13062 33338 13338 33400
rect 13462 33440 13738 33462
rect 13462 33400 13580 33440
rect 13620 33400 13738 33440
rect 13462 33338 13738 33400
rect 13862 33440 14138 33462
rect 13862 33400 13980 33440
rect 14020 33400 14138 33440
rect 13862 33338 14138 33400
rect 14262 33440 14538 33462
rect 14262 33400 14380 33440
rect 14420 33400 14538 33440
rect 14262 33338 14538 33400
rect 14662 33440 14938 33462
rect 14662 33400 14780 33440
rect 14820 33400 14938 33440
rect 14662 33338 14938 33400
rect 15062 33440 15338 33462
rect 15062 33400 15180 33440
rect 15220 33400 15338 33440
rect 15062 33338 15338 33400
rect 15462 33440 16000 33462
rect 15462 33400 15580 33440
rect 15620 33400 16000 33440
rect 15462 33338 16000 33400
rect 0 33062 16000 33338
rect 0 33040 538 33062
rect 0 33000 380 33040
rect 420 33000 538 33040
rect 0 32938 538 33000
rect 662 33040 938 33062
rect 662 33000 780 33040
rect 820 33000 938 33040
rect 662 32938 938 33000
rect 1062 33040 1338 33062
rect 1062 33000 1180 33040
rect 1220 33000 1338 33040
rect 1062 32938 1338 33000
rect 1462 33040 1738 33062
rect 1462 33000 1580 33040
rect 1620 33000 1738 33040
rect 1462 32938 1738 33000
rect 1862 33040 2138 33062
rect 1862 33000 1980 33040
rect 2020 33000 2138 33040
rect 1862 32938 2138 33000
rect 2262 33040 2538 33062
rect 2262 33000 2380 33040
rect 2420 33000 2538 33040
rect 2262 32938 2538 33000
rect 2662 33040 2938 33062
rect 2662 33000 2780 33040
rect 2820 33000 2938 33040
rect 2662 32938 2938 33000
rect 3062 33040 3338 33062
rect 3062 33000 3180 33040
rect 3220 33000 3338 33040
rect 3062 32938 3338 33000
rect 3462 33040 3738 33062
rect 3462 33000 3580 33040
rect 3620 33000 3738 33040
rect 3462 32938 3738 33000
rect 3862 33040 4138 33062
rect 3862 33000 3980 33040
rect 4020 33000 4138 33040
rect 3862 32938 4138 33000
rect 4262 33040 4538 33062
rect 4262 33000 4380 33040
rect 4420 33000 4538 33040
rect 4262 32938 4538 33000
rect 4662 33040 4938 33062
rect 4662 33000 4780 33040
rect 4820 33000 4938 33040
rect 4662 32938 4938 33000
rect 5062 33040 5338 33062
rect 5062 33000 5180 33040
rect 5220 33000 5338 33040
rect 5062 32938 5338 33000
rect 5462 33040 5738 33062
rect 5462 33000 5580 33040
rect 5620 33000 5738 33040
rect 5462 32938 5738 33000
rect 5862 33040 6138 33062
rect 5862 33000 5980 33040
rect 6020 33000 6138 33040
rect 5862 32938 6138 33000
rect 6262 33040 6538 33062
rect 6262 33000 6380 33040
rect 6420 33000 6538 33040
rect 6262 32938 6538 33000
rect 6662 33040 6938 33062
rect 6662 33000 6780 33040
rect 6820 33000 6938 33040
rect 6662 32938 6938 33000
rect 7062 33040 7338 33062
rect 7062 33000 7180 33040
rect 7220 33000 7338 33040
rect 7062 32938 7338 33000
rect 7462 33040 7738 33062
rect 7462 33000 7580 33040
rect 7620 33000 7738 33040
rect 7462 32938 7738 33000
rect 7862 33040 8138 33062
rect 7862 33000 7980 33040
rect 8020 33000 8138 33040
rect 7862 32938 8138 33000
rect 8262 33040 8538 33062
rect 8262 33000 8380 33040
rect 8420 33000 8538 33040
rect 8262 32938 8538 33000
rect 8662 33040 8938 33062
rect 8662 33000 8780 33040
rect 8820 33000 8938 33040
rect 8662 32938 8938 33000
rect 9062 33040 9338 33062
rect 9062 33000 9180 33040
rect 9220 33000 9338 33040
rect 9062 32938 9338 33000
rect 9462 33040 9738 33062
rect 9462 33000 9580 33040
rect 9620 33000 9738 33040
rect 9462 32938 9738 33000
rect 9862 33040 10138 33062
rect 9862 33000 9980 33040
rect 10020 33000 10138 33040
rect 9862 32938 10138 33000
rect 10262 33040 10538 33062
rect 10262 33000 10380 33040
rect 10420 33000 10538 33040
rect 10262 32938 10538 33000
rect 10662 33040 10938 33062
rect 10662 33000 10780 33040
rect 10820 33000 10938 33040
rect 10662 32938 10938 33000
rect 11062 33040 11338 33062
rect 11062 33000 11180 33040
rect 11220 33000 11338 33040
rect 11062 32938 11338 33000
rect 11462 33040 11738 33062
rect 11462 33000 11580 33040
rect 11620 33000 11738 33040
rect 11462 32938 11738 33000
rect 11862 33040 12138 33062
rect 11862 33000 11980 33040
rect 12020 33000 12138 33040
rect 11862 32938 12138 33000
rect 12262 33040 12538 33062
rect 12262 33000 12380 33040
rect 12420 33000 12538 33040
rect 12262 32938 12538 33000
rect 12662 33040 12938 33062
rect 12662 33000 12780 33040
rect 12820 33000 12938 33040
rect 12662 32938 12938 33000
rect 13062 33040 13338 33062
rect 13062 33000 13180 33040
rect 13220 33000 13338 33040
rect 13062 32938 13338 33000
rect 13462 33040 13738 33062
rect 13462 33000 13580 33040
rect 13620 33000 13738 33040
rect 13462 32938 13738 33000
rect 13862 33040 14138 33062
rect 13862 33000 13980 33040
rect 14020 33000 14138 33040
rect 13862 32938 14138 33000
rect 14262 33040 14538 33062
rect 14262 33000 14380 33040
rect 14420 33000 14538 33040
rect 14262 32938 14538 33000
rect 14662 33040 14938 33062
rect 14662 33000 14780 33040
rect 14820 33000 14938 33040
rect 14662 32938 14938 33000
rect 15062 33040 15338 33062
rect 15062 33000 15180 33040
rect 15220 33000 15338 33040
rect 15062 32938 15338 33000
rect 15462 33040 16000 33062
rect 15462 33000 15580 33040
rect 15620 33000 16000 33040
rect 15462 32938 16000 33000
rect 0 32662 16000 32938
rect 0 32538 538 32662
rect 662 32538 938 32662
rect 1062 32538 1338 32662
rect 1462 32538 1738 32662
rect 1862 32538 2138 32662
rect 2262 32538 2538 32662
rect 2662 32538 2938 32662
rect 3062 32538 3338 32662
rect 3462 32538 3738 32662
rect 3862 32538 4138 32662
rect 4262 32538 4538 32662
rect 4662 32538 4938 32662
rect 5062 32538 5338 32662
rect 5462 32538 5738 32662
rect 5862 32538 6138 32662
rect 6262 32538 6538 32662
rect 6662 32538 6938 32662
rect 7062 32538 7338 32662
rect 7462 32538 7738 32662
rect 7862 32538 8138 32662
rect 8262 32538 8538 32662
rect 8662 32538 8938 32662
rect 9062 32538 9338 32662
rect 9462 32538 9738 32662
rect 9862 32538 10138 32662
rect 10262 32538 10538 32662
rect 10662 32538 10938 32662
rect 11062 32538 11338 32662
rect 11462 32538 11738 32662
rect 11862 32538 12138 32662
rect 12262 32538 12538 32662
rect 12662 32538 12938 32662
rect 13062 32538 13338 32662
rect 13462 32538 13738 32662
rect 13862 32538 14138 32662
rect 14262 32538 14538 32662
rect 14662 32538 14938 32662
rect 15062 32538 15338 32662
rect 15462 32538 16000 32662
rect 0 32000 16000 32538
rect 0 31062 16000 31600
rect 0 30938 538 31062
rect 662 30938 938 31062
rect 1062 30938 1338 31062
rect 1462 30938 1738 31062
rect 1862 30938 2138 31062
rect 2262 30938 2538 31062
rect 2662 30938 2938 31062
rect 3062 30938 3338 31062
rect 3462 30938 3738 31062
rect 3862 30938 4138 31062
rect 4262 30938 4538 31062
rect 4662 30938 4938 31062
rect 5062 30938 5338 31062
rect 5462 30938 5738 31062
rect 5862 30938 6138 31062
rect 6262 30938 6538 31062
rect 6662 30938 6938 31062
rect 7062 30938 7338 31062
rect 7462 30938 7738 31062
rect 7862 30938 8138 31062
rect 8262 30938 8538 31062
rect 8662 30938 8938 31062
rect 9062 30938 9338 31062
rect 9462 30938 9738 31062
rect 9862 30938 10138 31062
rect 10262 30938 10538 31062
rect 10662 30938 10938 31062
rect 11062 30938 11338 31062
rect 11462 30938 11738 31062
rect 11862 30938 12138 31062
rect 12262 30938 12538 31062
rect 12662 30938 12938 31062
rect 13062 30938 13338 31062
rect 13462 30938 13738 31062
rect 13862 30938 14138 31062
rect 14262 30938 14538 31062
rect 14662 30938 14938 31062
rect 15062 30938 15338 31062
rect 15462 30938 16000 31062
rect 0 30662 16000 30938
rect 0 30600 538 30662
rect 0 30560 380 30600
rect 420 30560 538 30600
rect 0 30538 538 30560
rect 662 30600 938 30662
rect 662 30560 780 30600
rect 820 30560 938 30600
rect 662 30538 938 30560
rect 1062 30600 1338 30662
rect 1062 30560 1180 30600
rect 1220 30560 1338 30600
rect 1062 30538 1338 30560
rect 1462 30600 1738 30662
rect 1462 30560 1580 30600
rect 1620 30560 1738 30600
rect 1462 30538 1738 30560
rect 1862 30600 2138 30662
rect 1862 30560 1980 30600
rect 2020 30560 2138 30600
rect 1862 30538 2138 30560
rect 2262 30600 2538 30662
rect 2262 30560 2380 30600
rect 2420 30560 2538 30600
rect 2262 30538 2538 30560
rect 2662 30600 2938 30662
rect 2662 30560 2780 30600
rect 2820 30560 2938 30600
rect 2662 30538 2938 30560
rect 3062 30600 3338 30662
rect 3062 30560 3180 30600
rect 3220 30560 3338 30600
rect 3062 30538 3338 30560
rect 3462 30600 3738 30662
rect 3462 30560 3580 30600
rect 3620 30560 3738 30600
rect 3462 30538 3738 30560
rect 3862 30600 4138 30662
rect 3862 30560 3980 30600
rect 4020 30560 4138 30600
rect 3862 30538 4138 30560
rect 4262 30600 4538 30662
rect 4262 30560 4380 30600
rect 4420 30560 4538 30600
rect 4262 30538 4538 30560
rect 4662 30600 4938 30662
rect 4662 30560 4780 30600
rect 4820 30560 4938 30600
rect 4662 30538 4938 30560
rect 5062 30600 5338 30662
rect 5062 30560 5180 30600
rect 5220 30560 5338 30600
rect 5062 30538 5338 30560
rect 5462 30600 5738 30662
rect 5462 30560 5580 30600
rect 5620 30560 5738 30600
rect 5462 30538 5738 30560
rect 5862 30600 6138 30662
rect 5862 30560 5980 30600
rect 6020 30560 6138 30600
rect 5862 30538 6138 30560
rect 6262 30600 6538 30662
rect 6262 30560 6380 30600
rect 6420 30560 6538 30600
rect 6262 30538 6538 30560
rect 6662 30600 6938 30662
rect 6662 30560 6780 30600
rect 6820 30560 6938 30600
rect 6662 30538 6938 30560
rect 7062 30600 7338 30662
rect 7062 30560 7180 30600
rect 7220 30560 7338 30600
rect 7062 30538 7338 30560
rect 7462 30600 7738 30662
rect 7462 30560 7580 30600
rect 7620 30560 7738 30600
rect 7462 30538 7738 30560
rect 7862 30600 8138 30662
rect 7862 30560 7980 30600
rect 8020 30560 8138 30600
rect 7862 30538 8138 30560
rect 8262 30600 8538 30662
rect 8262 30560 8380 30600
rect 8420 30560 8538 30600
rect 8262 30538 8538 30560
rect 8662 30600 8938 30662
rect 8662 30560 8780 30600
rect 8820 30560 8938 30600
rect 8662 30538 8938 30560
rect 9062 30600 9338 30662
rect 9062 30560 9180 30600
rect 9220 30560 9338 30600
rect 9062 30538 9338 30560
rect 9462 30600 9738 30662
rect 9462 30560 9580 30600
rect 9620 30560 9738 30600
rect 9462 30538 9738 30560
rect 9862 30600 10138 30662
rect 9862 30560 9980 30600
rect 10020 30560 10138 30600
rect 9862 30538 10138 30560
rect 10262 30600 10538 30662
rect 10262 30560 10380 30600
rect 10420 30560 10538 30600
rect 10262 30538 10538 30560
rect 10662 30600 10938 30662
rect 10662 30560 10780 30600
rect 10820 30560 10938 30600
rect 10662 30538 10938 30560
rect 11062 30600 11338 30662
rect 11062 30560 11180 30600
rect 11220 30560 11338 30600
rect 11062 30538 11338 30560
rect 11462 30600 11738 30662
rect 11462 30560 11580 30600
rect 11620 30560 11738 30600
rect 11462 30538 11738 30560
rect 11862 30600 12138 30662
rect 11862 30560 11980 30600
rect 12020 30560 12138 30600
rect 11862 30538 12138 30560
rect 12262 30600 12538 30662
rect 12262 30560 12380 30600
rect 12420 30560 12538 30600
rect 12262 30538 12538 30560
rect 12662 30600 12938 30662
rect 12662 30560 12780 30600
rect 12820 30560 12938 30600
rect 12662 30538 12938 30560
rect 13062 30600 13338 30662
rect 13062 30560 13180 30600
rect 13220 30560 13338 30600
rect 13062 30538 13338 30560
rect 13462 30600 13738 30662
rect 13462 30560 13580 30600
rect 13620 30560 13738 30600
rect 13462 30538 13738 30560
rect 13862 30600 14138 30662
rect 13862 30560 13980 30600
rect 14020 30560 14138 30600
rect 13862 30538 14138 30560
rect 14262 30600 14538 30662
rect 14262 30560 14380 30600
rect 14420 30560 14538 30600
rect 14262 30538 14538 30560
rect 14662 30600 14938 30662
rect 14662 30560 14780 30600
rect 14820 30560 14938 30600
rect 14662 30538 14938 30560
rect 15062 30600 15338 30662
rect 15062 30560 15180 30600
rect 15220 30560 15338 30600
rect 15062 30538 15338 30560
rect 15462 30600 16000 30662
rect 15462 30560 15580 30600
rect 15620 30560 16000 30600
rect 15462 30538 16000 30560
rect 0 30262 16000 30538
rect 0 30200 538 30262
rect 0 30160 380 30200
rect 420 30160 538 30200
rect 0 30138 538 30160
rect 662 30200 938 30262
rect 662 30160 780 30200
rect 820 30160 938 30200
rect 662 30138 938 30160
rect 1062 30200 1338 30262
rect 1062 30160 1180 30200
rect 1220 30160 1338 30200
rect 1062 30138 1338 30160
rect 1462 30200 1738 30262
rect 1462 30160 1580 30200
rect 1620 30160 1738 30200
rect 1462 30138 1738 30160
rect 1862 30200 2138 30262
rect 1862 30160 1980 30200
rect 2020 30160 2138 30200
rect 1862 30138 2138 30160
rect 2262 30200 2538 30262
rect 2262 30160 2380 30200
rect 2420 30160 2538 30200
rect 2262 30138 2538 30160
rect 2662 30200 2938 30262
rect 2662 30160 2780 30200
rect 2820 30160 2938 30200
rect 2662 30138 2938 30160
rect 3062 30200 3338 30262
rect 3062 30160 3180 30200
rect 3220 30160 3338 30200
rect 3062 30138 3338 30160
rect 3462 30200 3738 30262
rect 3462 30160 3580 30200
rect 3620 30160 3738 30200
rect 3462 30138 3738 30160
rect 3862 30200 4138 30262
rect 3862 30160 3980 30200
rect 4020 30160 4138 30200
rect 3862 30138 4138 30160
rect 4262 30200 4538 30262
rect 4262 30160 4380 30200
rect 4420 30160 4538 30200
rect 4262 30138 4538 30160
rect 4662 30200 4938 30262
rect 4662 30160 4780 30200
rect 4820 30160 4938 30200
rect 4662 30138 4938 30160
rect 5062 30200 5338 30262
rect 5062 30160 5180 30200
rect 5220 30160 5338 30200
rect 5062 30138 5338 30160
rect 5462 30200 5738 30262
rect 5462 30160 5580 30200
rect 5620 30160 5738 30200
rect 5462 30138 5738 30160
rect 5862 30200 6138 30262
rect 5862 30160 5980 30200
rect 6020 30160 6138 30200
rect 5862 30138 6138 30160
rect 6262 30200 6538 30262
rect 6262 30160 6380 30200
rect 6420 30160 6538 30200
rect 6262 30138 6538 30160
rect 6662 30200 6938 30262
rect 6662 30160 6780 30200
rect 6820 30160 6938 30200
rect 6662 30138 6938 30160
rect 7062 30200 7338 30262
rect 7062 30160 7180 30200
rect 7220 30160 7338 30200
rect 7062 30138 7338 30160
rect 7462 30200 7738 30262
rect 7462 30160 7580 30200
rect 7620 30160 7738 30200
rect 7462 30138 7738 30160
rect 7862 30200 8138 30262
rect 7862 30160 7980 30200
rect 8020 30160 8138 30200
rect 7862 30138 8138 30160
rect 8262 30200 8538 30262
rect 8262 30160 8380 30200
rect 8420 30160 8538 30200
rect 8262 30138 8538 30160
rect 8662 30200 8938 30262
rect 8662 30160 8780 30200
rect 8820 30160 8938 30200
rect 8662 30138 8938 30160
rect 9062 30200 9338 30262
rect 9062 30160 9180 30200
rect 9220 30160 9338 30200
rect 9062 30138 9338 30160
rect 9462 30200 9738 30262
rect 9462 30160 9580 30200
rect 9620 30160 9738 30200
rect 9462 30138 9738 30160
rect 9862 30200 10138 30262
rect 9862 30160 9980 30200
rect 10020 30160 10138 30200
rect 9862 30138 10138 30160
rect 10262 30200 10538 30262
rect 10262 30160 10380 30200
rect 10420 30160 10538 30200
rect 10262 30138 10538 30160
rect 10662 30200 10938 30262
rect 10662 30160 10780 30200
rect 10820 30160 10938 30200
rect 10662 30138 10938 30160
rect 11062 30200 11338 30262
rect 11062 30160 11180 30200
rect 11220 30160 11338 30200
rect 11062 30138 11338 30160
rect 11462 30200 11738 30262
rect 11462 30160 11580 30200
rect 11620 30160 11738 30200
rect 11462 30138 11738 30160
rect 11862 30200 12138 30262
rect 11862 30160 11980 30200
rect 12020 30160 12138 30200
rect 11862 30138 12138 30160
rect 12262 30200 12538 30262
rect 12262 30160 12380 30200
rect 12420 30160 12538 30200
rect 12262 30138 12538 30160
rect 12662 30200 12938 30262
rect 12662 30160 12780 30200
rect 12820 30160 12938 30200
rect 12662 30138 12938 30160
rect 13062 30200 13338 30262
rect 13062 30160 13180 30200
rect 13220 30160 13338 30200
rect 13062 30138 13338 30160
rect 13462 30200 13738 30262
rect 13462 30160 13580 30200
rect 13620 30160 13738 30200
rect 13462 30138 13738 30160
rect 13862 30200 14138 30262
rect 13862 30160 13980 30200
rect 14020 30160 14138 30200
rect 13862 30138 14138 30160
rect 14262 30200 14538 30262
rect 14262 30160 14380 30200
rect 14420 30160 14538 30200
rect 14262 30138 14538 30160
rect 14662 30200 14938 30262
rect 14662 30160 14780 30200
rect 14820 30160 14938 30200
rect 14662 30138 14938 30160
rect 15062 30200 15338 30262
rect 15062 30160 15180 30200
rect 15220 30160 15338 30200
rect 15062 30138 15338 30160
rect 15462 30200 16000 30262
rect 15462 30160 15580 30200
rect 15620 30160 16000 30200
rect 15462 30138 16000 30160
rect 0 29862 16000 30138
rect 0 29800 538 29862
rect 0 29760 380 29800
rect 420 29760 538 29800
rect 0 29738 538 29760
rect 662 29800 938 29862
rect 662 29760 780 29800
rect 820 29760 938 29800
rect 662 29738 938 29760
rect 1062 29800 1338 29862
rect 1062 29760 1180 29800
rect 1220 29760 1338 29800
rect 1062 29738 1338 29760
rect 1462 29800 1738 29862
rect 1462 29760 1580 29800
rect 1620 29760 1738 29800
rect 1462 29738 1738 29760
rect 1862 29800 2138 29862
rect 1862 29760 1980 29800
rect 2020 29760 2138 29800
rect 1862 29738 2138 29760
rect 2262 29800 2538 29862
rect 2262 29760 2380 29800
rect 2420 29760 2538 29800
rect 2262 29738 2538 29760
rect 2662 29800 2938 29862
rect 2662 29760 2780 29800
rect 2820 29760 2938 29800
rect 2662 29738 2938 29760
rect 3062 29800 3338 29862
rect 3062 29760 3180 29800
rect 3220 29760 3338 29800
rect 3062 29738 3338 29760
rect 3462 29800 3738 29862
rect 3462 29760 3580 29800
rect 3620 29760 3738 29800
rect 3462 29738 3738 29760
rect 3862 29800 4138 29862
rect 3862 29760 3980 29800
rect 4020 29760 4138 29800
rect 3862 29738 4138 29760
rect 4262 29800 4538 29862
rect 4262 29760 4380 29800
rect 4420 29760 4538 29800
rect 4262 29738 4538 29760
rect 4662 29800 4938 29862
rect 4662 29760 4780 29800
rect 4820 29760 4938 29800
rect 4662 29738 4938 29760
rect 5062 29800 5338 29862
rect 5062 29760 5180 29800
rect 5220 29760 5338 29800
rect 5062 29738 5338 29760
rect 5462 29800 5738 29862
rect 5462 29760 5580 29800
rect 5620 29760 5738 29800
rect 5462 29738 5738 29760
rect 5862 29800 6138 29862
rect 5862 29760 5980 29800
rect 6020 29760 6138 29800
rect 5862 29738 6138 29760
rect 6262 29800 6538 29862
rect 6262 29760 6380 29800
rect 6420 29760 6538 29800
rect 6262 29738 6538 29760
rect 6662 29800 6938 29862
rect 6662 29760 6780 29800
rect 6820 29760 6938 29800
rect 6662 29738 6938 29760
rect 7062 29800 7338 29862
rect 7062 29760 7180 29800
rect 7220 29760 7338 29800
rect 7062 29738 7338 29760
rect 7462 29800 7738 29862
rect 7462 29760 7580 29800
rect 7620 29760 7738 29800
rect 7462 29738 7738 29760
rect 7862 29800 8138 29862
rect 7862 29760 7980 29800
rect 8020 29760 8138 29800
rect 7862 29738 8138 29760
rect 8262 29800 8538 29862
rect 8262 29760 8380 29800
rect 8420 29760 8538 29800
rect 8262 29738 8538 29760
rect 8662 29800 8938 29862
rect 8662 29760 8780 29800
rect 8820 29760 8938 29800
rect 8662 29738 8938 29760
rect 9062 29800 9338 29862
rect 9062 29760 9180 29800
rect 9220 29760 9338 29800
rect 9062 29738 9338 29760
rect 9462 29800 9738 29862
rect 9462 29760 9580 29800
rect 9620 29760 9738 29800
rect 9462 29738 9738 29760
rect 9862 29800 10138 29862
rect 9862 29760 9980 29800
rect 10020 29760 10138 29800
rect 9862 29738 10138 29760
rect 10262 29800 10538 29862
rect 10262 29760 10380 29800
rect 10420 29760 10538 29800
rect 10262 29738 10538 29760
rect 10662 29800 10938 29862
rect 10662 29760 10780 29800
rect 10820 29760 10938 29800
rect 10662 29738 10938 29760
rect 11062 29800 11338 29862
rect 11062 29760 11180 29800
rect 11220 29760 11338 29800
rect 11062 29738 11338 29760
rect 11462 29800 11738 29862
rect 11462 29760 11580 29800
rect 11620 29760 11738 29800
rect 11462 29738 11738 29760
rect 11862 29800 12138 29862
rect 11862 29760 11980 29800
rect 12020 29760 12138 29800
rect 11862 29738 12138 29760
rect 12262 29800 12538 29862
rect 12262 29760 12380 29800
rect 12420 29760 12538 29800
rect 12262 29738 12538 29760
rect 12662 29800 12938 29862
rect 12662 29760 12780 29800
rect 12820 29760 12938 29800
rect 12662 29738 12938 29760
rect 13062 29800 13338 29862
rect 13062 29760 13180 29800
rect 13220 29760 13338 29800
rect 13062 29738 13338 29760
rect 13462 29800 13738 29862
rect 13462 29760 13580 29800
rect 13620 29760 13738 29800
rect 13462 29738 13738 29760
rect 13862 29800 14138 29862
rect 13862 29760 13980 29800
rect 14020 29760 14138 29800
rect 13862 29738 14138 29760
rect 14262 29800 14538 29862
rect 14262 29760 14380 29800
rect 14420 29760 14538 29800
rect 14262 29738 14538 29760
rect 14662 29800 14938 29862
rect 14662 29760 14780 29800
rect 14820 29760 14938 29800
rect 14662 29738 14938 29760
rect 15062 29800 15338 29862
rect 15062 29760 15180 29800
rect 15220 29760 15338 29800
rect 15062 29738 15338 29760
rect 15462 29800 16000 29862
rect 15462 29760 15580 29800
rect 15620 29760 16000 29800
rect 15462 29738 16000 29760
rect 0 29462 16000 29738
rect 0 29400 538 29462
rect 0 29360 380 29400
rect 420 29360 538 29400
rect 0 29338 538 29360
rect 662 29400 938 29462
rect 662 29360 780 29400
rect 820 29360 938 29400
rect 662 29338 938 29360
rect 1062 29400 1338 29462
rect 1062 29360 1180 29400
rect 1220 29360 1338 29400
rect 1062 29338 1338 29360
rect 1462 29400 1738 29462
rect 1462 29360 1580 29400
rect 1620 29360 1738 29400
rect 1462 29338 1738 29360
rect 1862 29400 2138 29462
rect 1862 29360 1980 29400
rect 2020 29360 2138 29400
rect 1862 29338 2138 29360
rect 2262 29400 2538 29462
rect 2262 29360 2380 29400
rect 2420 29360 2538 29400
rect 2262 29338 2538 29360
rect 2662 29400 2938 29462
rect 2662 29360 2780 29400
rect 2820 29360 2938 29400
rect 2662 29338 2938 29360
rect 3062 29400 3338 29462
rect 3062 29360 3180 29400
rect 3220 29360 3338 29400
rect 3062 29338 3338 29360
rect 3462 29400 3738 29462
rect 3462 29360 3580 29400
rect 3620 29360 3738 29400
rect 3462 29338 3738 29360
rect 3862 29400 4138 29462
rect 3862 29360 3980 29400
rect 4020 29360 4138 29400
rect 3862 29338 4138 29360
rect 4262 29400 4538 29462
rect 4262 29360 4380 29400
rect 4420 29360 4538 29400
rect 4262 29338 4538 29360
rect 4662 29400 4938 29462
rect 4662 29360 4780 29400
rect 4820 29360 4938 29400
rect 4662 29338 4938 29360
rect 5062 29400 5338 29462
rect 5062 29360 5180 29400
rect 5220 29360 5338 29400
rect 5062 29338 5338 29360
rect 5462 29400 5738 29462
rect 5462 29360 5580 29400
rect 5620 29360 5738 29400
rect 5462 29338 5738 29360
rect 5862 29400 6138 29462
rect 5862 29360 5980 29400
rect 6020 29360 6138 29400
rect 5862 29338 6138 29360
rect 6262 29400 6538 29462
rect 6262 29360 6380 29400
rect 6420 29360 6538 29400
rect 6262 29338 6538 29360
rect 6662 29400 6938 29462
rect 6662 29360 6780 29400
rect 6820 29360 6938 29400
rect 6662 29338 6938 29360
rect 7062 29400 7338 29462
rect 7062 29360 7180 29400
rect 7220 29360 7338 29400
rect 7062 29338 7338 29360
rect 7462 29400 7738 29462
rect 7462 29360 7580 29400
rect 7620 29360 7738 29400
rect 7462 29338 7738 29360
rect 7862 29400 8138 29462
rect 7862 29360 7980 29400
rect 8020 29360 8138 29400
rect 7862 29338 8138 29360
rect 8262 29400 8538 29462
rect 8262 29360 8380 29400
rect 8420 29360 8538 29400
rect 8262 29338 8538 29360
rect 8662 29400 8938 29462
rect 8662 29360 8780 29400
rect 8820 29360 8938 29400
rect 8662 29338 8938 29360
rect 9062 29400 9338 29462
rect 9062 29360 9180 29400
rect 9220 29360 9338 29400
rect 9062 29338 9338 29360
rect 9462 29400 9738 29462
rect 9462 29360 9580 29400
rect 9620 29360 9738 29400
rect 9462 29338 9738 29360
rect 9862 29400 10138 29462
rect 9862 29360 9980 29400
rect 10020 29360 10138 29400
rect 9862 29338 10138 29360
rect 10262 29400 10538 29462
rect 10262 29360 10380 29400
rect 10420 29360 10538 29400
rect 10262 29338 10538 29360
rect 10662 29400 10938 29462
rect 10662 29360 10780 29400
rect 10820 29360 10938 29400
rect 10662 29338 10938 29360
rect 11062 29400 11338 29462
rect 11062 29360 11180 29400
rect 11220 29360 11338 29400
rect 11062 29338 11338 29360
rect 11462 29400 11738 29462
rect 11462 29360 11580 29400
rect 11620 29360 11738 29400
rect 11462 29338 11738 29360
rect 11862 29400 12138 29462
rect 11862 29360 11980 29400
rect 12020 29360 12138 29400
rect 11862 29338 12138 29360
rect 12262 29400 12538 29462
rect 12262 29360 12380 29400
rect 12420 29360 12538 29400
rect 12262 29338 12538 29360
rect 12662 29400 12938 29462
rect 12662 29360 12780 29400
rect 12820 29360 12938 29400
rect 12662 29338 12938 29360
rect 13062 29400 13338 29462
rect 13062 29360 13180 29400
rect 13220 29360 13338 29400
rect 13062 29338 13338 29360
rect 13462 29400 13738 29462
rect 13462 29360 13580 29400
rect 13620 29360 13738 29400
rect 13462 29338 13738 29360
rect 13862 29400 14138 29462
rect 13862 29360 13980 29400
rect 14020 29360 14138 29400
rect 13862 29338 14138 29360
rect 14262 29400 14538 29462
rect 14262 29360 14380 29400
rect 14420 29360 14538 29400
rect 14262 29338 14538 29360
rect 14662 29400 14938 29462
rect 14662 29360 14780 29400
rect 14820 29360 14938 29400
rect 14662 29338 14938 29360
rect 15062 29400 15338 29462
rect 15062 29360 15180 29400
rect 15220 29360 15338 29400
rect 15062 29338 15338 29360
rect 15462 29400 16000 29462
rect 15462 29360 15580 29400
rect 15620 29360 16000 29400
rect 15462 29338 16000 29360
rect 0 29062 16000 29338
rect 0 29000 538 29062
rect 0 28960 380 29000
rect 420 28960 538 29000
rect 0 28938 538 28960
rect 662 29000 938 29062
rect 662 28960 780 29000
rect 820 28960 938 29000
rect 662 28938 938 28960
rect 1062 29000 1338 29062
rect 1062 28960 1180 29000
rect 1220 28960 1338 29000
rect 1062 28938 1338 28960
rect 1462 29000 1738 29062
rect 1462 28960 1580 29000
rect 1620 28960 1738 29000
rect 1462 28938 1738 28960
rect 1862 29000 2138 29062
rect 1862 28960 1980 29000
rect 2020 28960 2138 29000
rect 1862 28938 2138 28960
rect 2262 29000 2538 29062
rect 2262 28960 2380 29000
rect 2420 28960 2538 29000
rect 2262 28938 2538 28960
rect 2662 29000 2938 29062
rect 2662 28960 2780 29000
rect 2820 28960 2938 29000
rect 2662 28938 2938 28960
rect 3062 29000 3338 29062
rect 3062 28960 3180 29000
rect 3220 28960 3338 29000
rect 3062 28938 3338 28960
rect 3462 29000 3738 29062
rect 3462 28960 3580 29000
rect 3620 28960 3738 29000
rect 3462 28938 3738 28960
rect 3862 29000 4138 29062
rect 3862 28960 3980 29000
rect 4020 28960 4138 29000
rect 3862 28938 4138 28960
rect 4262 29000 4538 29062
rect 4262 28960 4380 29000
rect 4420 28960 4538 29000
rect 4262 28938 4538 28960
rect 4662 29000 4938 29062
rect 4662 28960 4780 29000
rect 4820 28960 4938 29000
rect 4662 28938 4938 28960
rect 5062 29000 5338 29062
rect 5062 28960 5180 29000
rect 5220 28960 5338 29000
rect 5062 28938 5338 28960
rect 5462 29000 5738 29062
rect 5462 28960 5580 29000
rect 5620 28960 5738 29000
rect 5462 28938 5738 28960
rect 5862 29000 6138 29062
rect 5862 28960 5980 29000
rect 6020 28960 6138 29000
rect 5862 28938 6138 28960
rect 6262 29000 6538 29062
rect 6262 28960 6380 29000
rect 6420 28960 6538 29000
rect 6262 28938 6538 28960
rect 6662 29000 6938 29062
rect 6662 28960 6780 29000
rect 6820 28960 6938 29000
rect 6662 28938 6938 28960
rect 7062 29000 7338 29062
rect 7062 28960 7180 29000
rect 7220 28960 7338 29000
rect 7062 28938 7338 28960
rect 7462 29000 7738 29062
rect 7462 28960 7580 29000
rect 7620 28960 7738 29000
rect 7462 28938 7738 28960
rect 7862 29000 8138 29062
rect 7862 28960 7980 29000
rect 8020 28960 8138 29000
rect 7862 28938 8138 28960
rect 8262 29000 8538 29062
rect 8262 28960 8380 29000
rect 8420 28960 8538 29000
rect 8262 28938 8538 28960
rect 8662 29000 8938 29062
rect 8662 28960 8780 29000
rect 8820 28960 8938 29000
rect 8662 28938 8938 28960
rect 9062 29000 9338 29062
rect 9062 28960 9180 29000
rect 9220 28960 9338 29000
rect 9062 28938 9338 28960
rect 9462 29000 9738 29062
rect 9462 28960 9580 29000
rect 9620 28960 9738 29000
rect 9462 28938 9738 28960
rect 9862 29000 10138 29062
rect 9862 28960 9980 29000
rect 10020 28960 10138 29000
rect 9862 28938 10138 28960
rect 10262 29000 10538 29062
rect 10262 28960 10380 29000
rect 10420 28960 10538 29000
rect 10262 28938 10538 28960
rect 10662 29000 10938 29062
rect 10662 28960 10780 29000
rect 10820 28960 10938 29000
rect 10662 28938 10938 28960
rect 11062 29000 11338 29062
rect 11062 28960 11180 29000
rect 11220 28960 11338 29000
rect 11062 28938 11338 28960
rect 11462 29000 11738 29062
rect 11462 28960 11580 29000
rect 11620 28960 11738 29000
rect 11462 28938 11738 28960
rect 11862 29000 12138 29062
rect 11862 28960 11980 29000
rect 12020 28960 12138 29000
rect 11862 28938 12138 28960
rect 12262 29000 12538 29062
rect 12262 28960 12380 29000
rect 12420 28960 12538 29000
rect 12262 28938 12538 28960
rect 12662 29000 12938 29062
rect 12662 28960 12780 29000
rect 12820 28960 12938 29000
rect 12662 28938 12938 28960
rect 13062 29000 13338 29062
rect 13062 28960 13180 29000
rect 13220 28960 13338 29000
rect 13062 28938 13338 28960
rect 13462 29000 13738 29062
rect 13462 28960 13580 29000
rect 13620 28960 13738 29000
rect 13462 28938 13738 28960
rect 13862 29000 14138 29062
rect 13862 28960 13980 29000
rect 14020 28960 14138 29000
rect 13862 28938 14138 28960
rect 14262 29000 14538 29062
rect 14262 28960 14380 29000
rect 14420 28960 14538 29000
rect 14262 28938 14538 28960
rect 14662 29000 14938 29062
rect 14662 28960 14780 29000
rect 14820 28960 14938 29000
rect 14662 28938 14938 28960
rect 15062 29000 15338 29062
rect 15062 28960 15180 29000
rect 15220 28960 15338 29000
rect 15062 28938 15338 28960
rect 15462 29000 16000 29062
rect 15462 28960 15580 29000
rect 15620 28960 16000 29000
rect 15462 28938 16000 28960
rect 0 28662 16000 28938
rect 0 28600 538 28662
rect 0 28560 380 28600
rect 420 28560 538 28600
rect 0 28538 538 28560
rect 662 28600 938 28662
rect 662 28560 780 28600
rect 820 28560 938 28600
rect 662 28538 938 28560
rect 1062 28600 1338 28662
rect 1062 28560 1180 28600
rect 1220 28560 1338 28600
rect 1062 28538 1338 28560
rect 1462 28600 1738 28662
rect 1462 28560 1580 28600
rect 1620 28560 1738 28600
rect 1462 28538 1738 28560
rect 1862 28600 2138 28662
rect 1862 28560 1980 28600
rect 2020 28560 2138 28600
rect 1862 28538 2138 28560
rect 2262 28600 2538 28662
rect 2262 28560 2380 28600
rect 2420 28560 2538 28600
rect 2262 28538 2538 28560
rect 2662 28600 2938 28662
rect 2662 28560 2780 28600
rect 2820 28560 2938 28600
rect 2662 28538 2938 28560
rect 3062 28600 3338 28662
rect 3062 28560 3180 28600
rect 3220 28560 3338 28600
rect 3062 28538 3338 28560
rect 3462 28600 3738 28662
rect 3462 28560 3580 28600
rect 3620 28560 3738 28600
rect 3462 28538 3738 28560
rect 3862 28600 4138 28662
rect 3862 28560 3980 28600
rect 4020 28560 4138 28600
rect 3862 28538 4138 28560
rect 4262 28600 4538 28662
rect 4262 28560 4380 28600
rect 4420 28560 4538 28600
rect 4262 28538 4538 28560
rect 4662 28600 4938 28662
rect 4662 28560 4780 28600
rect 4820 28560 4938 28600
rect 4662 28538 4938 28560
rect 5062 28600 5338 28662
rect 5062 28560 5180 28600
rect 5220 28560 5338 28600
rect 5062 28538 5338 28560
rect 5462 28600 5738 28662
rect 5462 28560 5580 28600
rect 5620 28560 5738 28600
rect 5462 28538 5738 28560
rect 5862 28600 6138 28662
rect 5862 28560 5980 28600
rect 6020 28560 6138 28600
rect 5862 28538 6138 28560
rect 6262 28600 6538 28662
rect 6262 28560 6380 28600
rect 6420 28560 6538 28600
rect 6262 28538 6538 28560
rect 6662 28600 6938 28662
rect 6662 28560 6780 28600
rect 6820 28560 6938 28600
rect 6662 28538 6938 28560
rect 7062 28600 7338 28662
rect 7062 28560 7180 28600
rect 7220 28560 7338 28600
rect 7062 28538 7338 28560
rect 7462 28600 7738 28662
rect 7462 28560 7580 28600
rect 7620 28560 7738 28600
rect 7462 28538 7738 28560
rect 7862 28600 8138 28662
rect 7862 28560 7980 28600
rect 8020 28560 8138 28600
rect 7862 28538 8138 28560
rect 8262 28600 8538 28662
rect 8262 28560 8380 28600
rect 8420 28560 8538 28600
rect 8262 28538 8538 28560
rect 8662 28600 8938 28662
rect 8662 28560 8780 28600
rect 8820 28560 8938 28600
rect 8662 28538 8938 28560
rect 9062 28600 9338 28662
rect 9062 28560 9180 28600
rect 9220 28560 9338 28600
rect 9062 28538 9338 28560
rect 9462 28600 9738 28662
rect 9462 28560 9580 28600
rect 9620 28560 9738 28600
rect 9462 28538 9738 28560
rect 9862 28600 10138 28662
rect 9862 28560 9980 28600
rect 10020 28560 10138 28600
rect 9862 28538 10138 28560
rect 10262 28600 10538 28662
rect 10262 28560 10380 28600
rect 10420 28560 10538 28600
rect 10262 28538 10538 28560
rect 10662 28600 10938 28662
rect 10662 28560 10780 28600
rect 10820 28560 10938 28600
rect 10662 28538 10938 28560
rect 11062 28600 11338 28662
rect 11062 28560 11180 28600
rect 11220 28560 11338 28600
rect 11062 28538 11338 28560
rect 11462 28600 11738 28662
rect 11462 28560 11580 28600
rect 11620 28560 11738 28600
rect 11462 28538 11738 28560
rect 11862 28600 12138 28662
rect 11862 28560 11980 28600
rect 12020 28560 12138 28600
rect 11862 28538 12138 28560
rect 12262 28600 12538 28662
rect 12262 28560 12380 28600
rect 12420 28560 12538 28600
rect 12262 28538 12538 28560
rect 12662 28600 12938 28662
rect 12662 28560 12780 28600
rect 12820 28560 12938 28600
rect 12662 28538 12938 28560
rect 13062 28600 13338 28662
rect 13062 28560 13180 28600
rect 13220 28560 13338 28600
rect 13062 28538 13338 28560
rect 13462 28600 13738 28662
rect 13462 28560 13580 28600
rect 13620 28560 13738 28600
rect 13462 28538 13738 28560
rect 13862 28600 14138 28662
rect 13862 28560 13980 28600
rect 14020 28560 14138 28600
rect 13862 28538 14138 28560
rect 14262 28600 14538 28662
rect 14262 28560 14380 28600
rect 14420 28560 14538 28600
rect 14262 28538 14538 28560
rect 14662 28600 14938 28662
rect 14662 28560 14780 28600
rect 14820 28560 14938 28600
rect 14662 28538 14938 28560
rect 15062 28600 15338 28662
rect 15062 28560 15180 28600
rect 15220 28560 15338 28600
rect 15062 28538 15338 28560
rect 15462 28600 16000 28662
rect 15462 28560 15580 28600
rect 15620 28560 16000 28600
rect 15462 28538 16000 28560
rect 0 28000 16000 28538
rect 0 26420 16000 26800
rect 0 26380 380 26420
rect 420 26380 780 26420
rect 820 26380 1180 26420
rect 1220 26380 1580 26420
rect 1620 26380 1980 26420
rect 2020 26380 2380 26420
rect 2420 26380 2780 26420
rect 2820 26380 3180 26420
rect 3220 26380 3580 26420
rect 3620 26380 3980 26420
rect 4020 26380 4380 26420
rect 4420 26380 4780 26420
rect 4820 26380 5180 26420
rect 5220 26380 5580 26420
rect 5620 26380 5980 26420
rect 6020 26380 6380 26420
rect 6420 26380 6780 26420
rect 6820 26380 7180 26420
rect 7220 26380 7580 26420
rect 7620 26380 7980 26420
rect 8020 26380 8380 26420
rect 8420 26380 8780 26420
rect 8820 26380 9180 26420
rect 9220 26380 9580 26420
rect 9620 26380 9980 26420
rect 10020 26380 10380 26420
rect 10420 26380 10780 26420
rect 10820 26380 11180 26420
rect 11220 26380 11580 26420
rect 11620 26380 11980 26420
rect 12020 26380 12380 26420
rect 12420 26380 12780 26420
rect 12820 26380 13180 26420
rect 13220 26380 13580 26420
rect 13620 26380 13980 26420
rect 14020 26380 14380 26420
rect 14420 26380 14780 26420
rect 14820 26380 15180 26420
rect 15220 26380 15580 26420
rect 15620 26380 16000 26420
rect 0 26262 16000 26380
rect 0 26138 538 26262
rect 662 26138 938 26262
rect 1062 26138 1338 26262
rect 1462 26138 1738 26262
rect 1862 26138 2138 26262
rect 2262 26138 2538 26262
rect 2662 26138 2938 26262
rect 3062 26138 3338 26262
rect 3462 26138 3738 26262
rect 3862 26138 4138 26262
rect 4262 26138 4538 26262
rect 4662 26138 4938 26262
rect 5062 26138 5338 26262
rect 5462 26138 5738 26262
rect 5862 26138 6138 26262
rect 6262 26138 6538 26262
rect 6662 26138 6938 26262
rect 7062 26138 7338 26262
rect 7462 26138 7738 26262
rect 7862 26138 8138 26262
rect 8262 26138 8538 26262
rect 8662 26138 8938 26262
rect 9062 26138 9338 26262
rect 9462 26138 9738 26262
rect 9862 26138 10138 26262
rect 10262 26138 10538 26262
rect 10662 26138 10938 26262
rect 11062 26138 11338 26262
rect 11462 26138 11738 26262
rect 11862 26138 12138 26262
rect 12262 26138 12538 26262
rect 12662 26138 12938 26262
rect 13062 26138 13338 26262
rect 13462 26138 13738 26262
rect 13862 26138 14138 26262
rect 14262 26138 14538 26262
rect 14662 26138 14938 26262
rect 15062 26138 15338 26262
rect 15462 26138 16000 26262
rect 0 26020 16000 26138
rect 0 25980 380 26020
rect 420 25980 780 26020
rect 820 25980 1180 26020
rect 1220 25980 1580 26020
rect 1620 25980 1980 26020
rect 2020 25980 2380 26020
rect 2420 25980 2780 26020
rect 2820 25980 3180 26020
rect 3220 25980 3580 26020
rect 3620 25980 3980 26020
rect 4020 25980 4380 26020
rect 4420 25980 4780 26020
rect 4820 25980 5180 26020
rect 5220 25980 5580 26020
rect 5620 25980 5980 26020
rect 6020 25980 6380 26020
rect 6420 25980 6780 26020
rect 6820 25980 7180 26020
rect 7220 25980 7580 26020
rect 7620 25980 7980 26020
rect 8020 25980 8380 26020
rect 8420 25980 8780 26020
rect 8820 25980 9180 26020
rect 9220 25980 9580 26020
rect 9620 25980 9980 26020
rect 10020 25980 10380 26020
rect 10420 25980 10780 26020
rect 10820 25980 11180 26020
rect 11220 25980 11580 26020
rect 11620 25980 11980 26020
rect 12020 25980 12380 26020
rect 12420 25980 12780 26020
rect 12820 25980 13180 26020
rect 13220 25980 13580 26020
rect 13620 25980 13980 26020
rect 14020 25980 14380 26020
rect 14420 25980 14780 26020
rect 14820 25980 15180 26020
rect 15220 25980 15580 26020
rect 15620 25980 16000 26020
rect 0 25862 16000 25980
rect 0 25738 538 25862
rect 662 25738 938 25862
rect 1062 25738 1338 25862
rect 1462 25738 1738 25862
rect 1862 25738 2138 25862
rect 2262 25738 2538 25862
rect 2662 25738 2938 25862
rect 3062 25738 3338 25862
rect 3462 25738 3738 25862
rect 3862 25738 4138 25862
rect 4262 25738 4538 25862
rect 4662 25738 4938 25862
rect 5062 25738 5338 25862
rect 5462 25738 5738 25862
rect 5862 25738 6138 25862
rect 6262 25738 6538 25862
rect 6662 25738 6938 25862
rect 7062 25738 7338 25862
rect 7462 25738 7738 25862
rect 7862 25738 8138 25862
rect 8262 25738 8538 25862
rect 8662 25738 8938 25862
rect 9062 25738 9338 25862
rect 9462 25738 9738 25862
rect 9862 25738 10138 25862
rect 10262 25738 10538 25862
rect 10662 25738 10938 25862
rect 11062 25738 11338 25862
rect 11462 25738 11738 25862
rect 11862 25738 12138 25862
rect 12262 25738 12538 25862
rect 12662 25738 12938 25862
rect 13062 25738 13338 25862
rect 13462 25738 13738 25862
rect 13862 25738 14138 25862
rect 14262 25738 14538 25862
rect 14662 25738 14938 25862
rect 15062 25738 15338 25862
rect 15462 25738 16000 25862
rect 0 25620 16000 25738
rect 0 25580 380 25620
rect 420 25580 780 25620
rect 820 25580 1180 25620
rect 1220 25580 1580 25620
rect 1620 25580 1980 25620
rect 2020 25580 2380 25620
rect 2420 25580 2780 25620
rect 2820 25580 3180 25620
rect 3220 25580 3580 25620
rect 3620 25580 3980 25620
rect 4020 25580 4380 25620
rect 4420 25580 4780 25620
rect 4820 25580 5180 25620
rect 5220 25580 5580 25620
rect 5620 25580 5980 25620
rect 6020 25580 6380 25620
rect 6420 25580 6780 25620
rect 6820 25580 7180 25620
rect 7220 25580 7580 25620
rect 7620 25580 7980 25620
rect 8020 25580 8380 25620
rect 8420 25580 8780 25620
rect 8820 25580 9180 25620
rect 9220 25580 9580 25620
rect 9620 25580 9980 25620
rect 10020 25580 10380 25620
rect 10420 25580 10780 25620
rect 10820 25580 11180 25620
rect 11220 25580 11580 25620
rect 11620 25580 11980 25620
rect 12020 25580 12380 25620
rect 12420 25580 12780 25620
rect 12820 25580 13180 25620
rect 13220 25580 13580 25620
rect 13620 25580 13980 25620
rect 14020 25580 14380 25620
rect 14420 25580 14780 25620
rect 14820 25580 15180 25620
rect 15220 25580 15580 25620
rect 15620 25580 16000 25620
rect 0 25200 16000 25580
rect 0 23312 16000 23800
rect 0 23270 538 23312
rect 0 23230 380 23270
rect 420 23230 538 23270
rect 0 23188 538 23230
rect 662 23270 938 23312
rect 662 23230 780 23270
rect 820 23230 938 23270
rect 662 23188 938 23230
rect 1062 23270 1338 23312
rect 1062 23230 1180 23270
rect 1220 23230 1338 23270
rect 1062 23188 1338 23230
rect 1462 23270 1738 23312
rect 1462 23230 1580 23270
rect 1620 23230 1738 23270
rect 1462 23188 1738 23230
rect 1862 23270 2138 23312
rect 1862 23230 1980 23270
rect 2020 23230 2138 23270
rect 1862 23188 2138 23230
rect 2262 23270 2538 23312
rect 2262 23230 2380 23270
rect 2420 23230 2538 23270
rect 2262 23188 2538 23230
rect 2662 23270 2938 23312
rect 2662 23230 2780 23270
rect 2820 23230 2938 23270
rect 2662 23188 2938 23230
rect 3062 23270 3338 23312
rect 3062 23230 3180 23270
rect 3220 23230 3338 23270
rect 3062 23188 3338 23230
rect 3462 23270 3738 23312
rect 3462 23230 3580 23270
rect 3620 23230 3738 23270
rect 3462 23188 3738 23230
rect 3862 23270 4138 23312
rect 3862 23230 3980 23270
rect 4020 23230 4138 23270
rect 3862 23188 4138 23230
rect 4262 23270 4538 23312
rect 4262 23230 4380 23270
rect 4420 23230 4538 23270
rect 4262 23188 4538 23230
rect 4662 23270 4938 23312
rect 4662 23230 4780 23270
rect 4820 23230 4938 23270
rect 4662 23188 4938 23230
rect 5062 23270 5338 23312
rect 5062 23230 5180 23270
rect 5220 23230 5338 23270
rect 5062 23188 5338 23230
rect 5462 23270 5738 23312
rect 5462 23230 5580 23270
rect 5620 23230 5738 23270
rect 5462 23188 5738 23230
rect 5862 23270 6138 23312
rect 5862 23230 5980 23270
rect 6020 23230 6138 23270
rect 5862 23188 6138 23230
rect 6262 23270 6538 23312
rect 6262 23230 6380 23270
rect 6420 23230 6538 23270
rect 6262 23188 6538 23230
rect 6662 23270 6938 23312
rect 6662 23230 6780 23270
rect 6820 23230 6938 23270
rect 6662 23188 6938 23230
rect 7062 23270 7338 23312
rect 7062 23230 7180 23270
rect 7220 23230 7338 23270
rect 7062 23188 7338 23230
rect 7462 23270 7738 23312
rect 7462 23230 7580 23270
rect 7620 23230 7738 23270
rect 7462 23188 7738 23230
rect 7862 23270 8138 23312
rect 7862 23230 7980 23270
rect 8020 23230 8138 23270
rect 7862 23188 8138 23230
rect 8262 23270 8538 23312
rect 8262 23230 8380 23270
rect 8420 23230 8538 23270
rect 8262 23188 8538 23230
rect 8662 23270 8938 23312
rect 8662 23230 8780 23270
rect 8820 23230 8938 23270
rect 8662 23188 8938 23230
rect 9062 23270 9338 23312
rect 9062 23230 9180 23270
rect 9220 23230 9338 23270
rect 9062 23188 9338 23230
rect 9462 23270 9738 23312
rect 9462 23230 9580 23270
rect 9620 23230 9738 23270
rect 9462 23188 9738 23230
rect 9862 23270 10138 23312
rect 9862 23230 9980 23270
rect 10020 23230 10138 23270
rect 9862 23188 10138 23230
rect 10262 23270 10538 23312
rect 10262 23230 10380 23270
rect 10420 23230 10538 23270
rect 10262 23188 10538 23230
rect 10662 23270 10938 23312
rect 10662 23230 10780 23270
rect 10820 23230 10938 23270
rect 10662 23188 10938 23230
rect 11062 23270 11338 23312
rect 11062 23230 11180 23270
rect 11220 23230 11338 23270
rect 11062 23188 11338 23230
rect 11462 23270 11738 23312
rect 11462 23230 11580 23270
rect 11620 23230 11738 23270
rect 11462 23188 11738 23230
rect 11862 23270 12138 23312
rect 11862 23230 11980 23270
rect 12020 23230 12138 23270
rect 11862 23188 12138 23230
rect 12262 23270 12538 23312
rect 12262 23230 12380 23270
rect 12420 23230 12538 23270
rect 12262 23188 12538 23230
rect 12662 23270 12938 23312
rect 12662 23230 12780 23270
rect 12820 23230 12938 23270
rect 12662 23188 12938 23230
rect 13062 23270 13338 23312
rect 13062 23230 13180 23270
rect 13220 23230 13338 23270
rect 13062 23188 13338 23230
rect 13462 23270 13738 23312
rect 13462 23230 13580 23270
rect 13620 23230 13738 23270
rect 13462 23188 13738 23230
rect 13862 23270 14138 23312
rect 13862 23230 13980 23270
rect 14020 23230 14138 23270
rect 13862 23188 14138 23230
rect 14262 23270 14538 23312
rect 14262 23230 14380 23270
rect 14420 23230 14538 23270
rect 14262 23188 14538 23230
rect 14662 23270 14938 23312
rect 14662 23230 14780 23270
rect 14820 23230 14938 23270
rect 14662 23188 14938 23230
rect 15062 23270 15338 23312
rect 15062 23230 15180 23270
rect 15220 23230 15338 23270
rect 15062 23188 15338 23230
rect 15462 23270 16000 23312
rect 15462 23230 15580 23270
rect 15620 23230 16000 23270
rect 15462 23188 16000 23230
rect 0 22912 16000 23188
rect 0 22870 538 22912
rect 0 22830 380 22870
rect 420 22830 538 22870
rect 0 22788 538 22830
rect 662 22870 938 22912
rect 662 22830 780 22870
rect 820 22830 938 22870
rect 662 22788 938 22830
rect 1062 22870 1338 22912
rect 1062 22830 1180 22870
rect 1220 22830 1338 22870
rect 1062 22788 1338 22830
rect 1462 22870 1738 22912
rect 1462 22830 1580 22870
rect 1620 22830 1738 22870
rect 1462 22788 1738 22830
rect 1862 22870 2138 22912
rect 1862 22830 1980 22870
rect 2020 22830 2138 22870
rect 1862 22788 2138 22830
rect 2262 22870 2538 22912
rect 2262 22830 2380 22870
rect 2420 22830 2538 22870
rect 2262 22788 2538 22830
rect 2662 22870 2938 22912
rect 2662 22830 2780 22870
rect 2820 22830 2938 22870
rect 2662 22788 2938 22830
rect 3062 22870 3338 22912
rect 3062 22830 3180 22870
rect 3220 22830 3338 22870
rect 3062 22788 3338 22830
rect 3462 22870 3738 22912
rect 3462 22830 3580 22870
rect 3620 22830 3738 22870
rect 3462 22788 3738 22830
rect 3862 22870 4138 22912
rect 3862 22830 3980 22870
rect 4020 22830 4138 22870
rect 3862 22788 4138 22830
rect 4262 22870 4538 22912
rect 4262 22830 4380 22870
rect 4420 22830 4538 22870
rect 4262 22788 4538 22830
rect 4662 22870 4938 22912
rect 4662 22830 4780 22870
rect 4820 22830 4938 22870
rect 4662 22788 4938 22830
rect 5062 22870 5338 22912
rect 5062 22830 5180 22870
rect 5220 22830 5338 22870
rect 5062 22788 5338 22830
rect 5462 22870 5738 22912
rect 5462 22830 5580 22870
rect 5620 22830 5738 22870
rect 5462 22788 5738 22830
rect 5862 22870 6138 22912
rect 5862 22830 5980 22870
rect 6020 22830 6138 22870
rect 5862 22788 6138 22830
rect 6262 22870 6538 22912
rect 6262 22830 6380 22870
rect 6420 22830 6538 22870
rect 6262 22788 6538 22830
rect 6662 22870 6938 22912
rect 6662 22830 6780 22870
rect 6820 22830 6938 22870
rect 6662 22788 6938 22830
rect 7062 22870 7338 22912
rect 7062 22830 7180 22870
rect 7220 22830 7338 22870
rect 7062 22788 7338 22830
rect 7462 22870 7738 22912
rect 7462 22830 7580 22870
rect 7620 22830 7738 22870
rect 7462 22788 7738 22830
rect 7862 22870 8138 22912
rect 7862 22830 7980 22870
rect 8020 22830 8138 22870
rect 7862 22788 8138 22830
rect 8262 22870 8538 22912
rect 8262 22830 8380 22870
rect 8420 22830 8538 22870
rect 8262 22788 8538 22830
rect 8662 22870 8938 22912
rect 8662 22830 8780 22870
rect 8820 22830 8938 22870
rect 8662 22788 8938 22830
rect 9062 22870 9338 22912
rect 9062 22830 9180 22870
rect 9220 22830 9338 22870
rect 9062 22788 9338 22830
rect 9462 22870 9738 22912
rect 9462 22830 9580 22870
rect 9620 22830 9738 22870
rect 9462 22788 9738 22830
rect 9862 22870 10138 22912
rect 9862 22830 9980 22870
rect 10020 22830 10138 22870
rect 9862 22788 10138 22830
rect 10262 22870 10538 22912
rect 10262 22830 10380 22870
rect 10420 22830 10538 22870
rect 10262 22788 10538 22830
rect 10662 22870 10938 22912
rect 10662 22830 10780 22870
rect 10820 22830 10938 22870
rect 10662 22788 10938 22830
rect 11062 22870 11338 22912
rect 11062 22830 11180 22870
rect 11220 22830 11338 22870
rect 11062 22788 11338 22830
rect 11462 22870 11738 22912
rect 11462 22830 11580 22870
rect 11620 22830 11738 22870
rect 11462 22788 11738 22830
rect 11862 22870 12138 22912
rect 11862 22830 11980 22870
rect 12020 22830 12138 22870
rect 11862 22788 12138 22830
rect 12262 22870 12538 22912
rect 12262 22830 12380 22870
rect 12420 22830 12538 22870
rect 12262 22788 12538 22830
rect 12662 22870 12938 22912
rect 12662 22830 12780 22870
rect 12820 22830 12938 22870
rect 12662 22788 12938 22830
rect 13062 22870 13338 22912
rect 13062 22830 13180 22870
rect 13220 22830 13338 22870
rect 13062 22788 13338 22830
rect 13462 22870 13738 22912
rect 13462 22830 13580 22870
rect 13620 22830 13738 22870
rect 13462 22788 13738 22830
rect 13862 22870 14138 22912
rect 13862 22830 13980 22870
rect 14020 22830 14138 22870
rect 13862 22788 14138 22830
rect 14262 22870 14538 22912
rect 14262 22830 14380 22870
rect 14420 22830 14538 22870
rect 14262 22788 14538 22830
rect 14662 22870 14938 22912
rect 14662 22830 14780 22870
rect 14820 22830 14938 22870
rect 14662 22788 14938 22830
rect 15062 22870 15338 22912
rect 15062 22830 15180 22870
rect 15220 22830 15338 22870
rect 15062 22788 15338 22830
rect 15462 22870 16000 22912
rect 15462 22830 15580 22870
rect 15620 22830 16000 22870
rect 15462 22788 16000 22830
rect 0 22512 16000 22788
rect 0 22470 538 22512
rect 0 22430 380 22470
rect 420 22430 538 22470
rect 0 22388 538 22430
rect 662 22470 938 22512
rect 662 22430 780 22470
rect 820 22430 938 22470
rect 662 22388 938 22430
rect 1062 22470 1338 22512
rect 1062 22430 1180 22470
rect 1220 22430 1338 22470
rect 1062 22388 1338 22430
rect 1462 22470 1738 22512
rect 1462 22430 1580 22470
rect 1620 22430 1738 22470
rect 1462 22388 1738 22430
rect 1862 22470 2138 22512
rect 1862 22430 1980 22470
rect 2020 22430 2138 22470
rect 1862 22388 2138 22430
rect 2262 22470 2538 22512
rect 2262 22430 2380 22470
rect 2420 22430 2538 22470
rect 2262 22388 2538 22430
rect 2662 22470 2938 22512
rect 2662 22430 2780 22470
rect 2820 22430 2938 22470
rect 2662 22388 2938 22430
rect 3062 22470 3338 22512
rect 3062 22430 3180 22470
rect 3220 22430 3338 22470
rect 3062 22388 3338 22430
rect 3462 22470 3738 22512
rect 3462 22430 3580 22470
rect 3620 22430 3738 22470
rect 3462 22388 3738 22430
rect 3862 22470 4138 22512
rect 3862 22430 3980 22470
rect 4020 22430 4138 22470
rect 3862 22388 4138 22430
rect 4262 22470 4538 22512
rect 4262 22430 4380 22470
rect 4420 22430 4538 22470
rect 4262 22388 4538 22430
rect 4662 22470 4938 22512
rect 4662 22430 4780 22470
rect 4820 22430 4938 22470
rect 4662 22388 4938 22430
rect 5062 22470 5338 22512
rect 5062 22430 5180 22470
rect 5220 22430 5338 22470
rect 5062 22388 5338 22430
rect 5462 22470 5738 22512
rect 5462 22430 5580 22470
rect 5620 22430 5738 22470
rect 5462 22388 5738 22430
rect 5862 22470 6138 22512
rect 5862 22430 5980 22470
rect 6020 22430 6138 22470
rect 5862 22388 6138 22430
rect 6262 22470 6538 22512
rect 6262 22430 6380 22470
rect 6420 22430 6538 22470
rect 6262 22388 6538 22430
rect 6662 22470 6938 22512
rect 6662 22430 6780 22470
rect 6820 22430 6938 22470
rect 6662 22388 6938 22430
rect 7062 22470 7338 22512
rect 7062 22430 7180 22470
rect 7220 22430 7338 22470
rect 7062 22388 7338 22430
rect 7462 22470 7738 22512
rect 7462 22430 7580 22470
rect 7620 22430 7738 22470
rect 7462 22388 7738 22430
rect 7862 22470 8138 22512
rect 7862 22430 7980 22470
rect 8020 22430 8138 22470
rect 7862 22388 8138 22430
rect 8262 22470 8538 22512
rect 8262 22430 8380 22470
rect 8420 22430 8538 22470
rect 8262 22388 8538 22430
rect 8662 22470 8938 22512
rect 8662 22430 8780 22470
rect 8820 22430 8938 22470
rect 8662 22388 8938 22430
rect 9062 22470 9338 22512
rect 9062 22430 9180 22470
rect 9220 22430 9338 22470
rect 9062 22388 9338 22430
rect 9462 22470 9738 22512
rect 9462 22430 9580 22470
rect 9620 22430 9738 22470
rect 9462 22388 9738 22430
rect 9862 22470 10138 22512
rect 9862 22430 9980 22470
rect 10020 22430 10138 22470
rect 9862 22388 10138 22430
rect 10262 22470 10538 22512
rect 10262 22430 10380 22470
rect 10420 22430 10538 22470
rect 10262 22388 10538 22430
rect 10662 22470 10938 22512
rect 10662 22430 10780 22470
rect 10820 22430 10938 22470
rect 10662 22388 10938 22430
rect 11062 22470 11338 22512
rect 11062 22430 11180 22470
rect 11220 22430 11338 22470
rect 11062 22388 11338 22430
rect 11462 22470 11738 22512
rect 11462 22430 11580 22470
rect 11620 22430 11738 22470
rect 11462 22388 11738 22430
rect 11862 22470 12138 22512
rect 11862 22430 11980 22470
rect 12020 22430 12138 22470
rect 11862 22388 12138 22430
rect 12262 22470 12538 22512
rect 12262 22430 12380 22470
rect 12420 22430 12538 22470
rect 12262 22388 12538 22430
rect 12662 22470 12938 22512
rect 12662 22430 12780 22470
rect 12820 22430 12938 22470
rect 12662 22388 12938 22430
rect 13062 22470 13338 22512
rect 13062 22430 13180 22470
rect 13220 22430 13338 22470
rect 13062 22388 13338 22430
rect 13462 22470 13738 22512
rect 13462 22430 13580 22470
rect 13620 22430 13738 22470
rect 13462 22388 13738 22430
rect 13862 22470 14138 22512
rect 13862 22430 13980 22470
rect 14020 22430 14138 22470
rect 13862 22388 14138 22430
rect 14262 22470 14538 22512
rect 14262 22430 14380 22470
rect 14420 22430 14538 22470
rect 14262 22388 14538 22430
rect 14662 22470 14938 22512
rect 14662 22430 14780 22470
rect 14820 22430 14938 22470
rect 14662 22388 14938 22430
rect 15062 22470 15338 22512
rect 15062 22430 15180 22470
rect 15220 22430 15338 22470
rect 15062 22388 15338 22430
rect 15462 22470 16000 22512
rect 15462 22430 15580 22470
rect 15620 22430 16000 22470
rect 15462 22388 16000 22430
rect 0 22112 16000 22388
rect 0 22070 538 22112
rect 0 22030 380 22070
rect 420 22030 538 22070
rect 0 21988 538 22030
rect 662 22070 938 22112
rect 662 22030 780 22070
rect 820 22030 938 22070
rect 662 21988 938 22030
rect 1062 22070 1338 22112
rect 1062 22030 1180 22070
rect 1220 22030 1338 22070
rect 1062 21988 1338 22030
rect 1462 22070 1738 22112
rect 1462 22030 1580 22070
rect 1620 22030 1738 22070
rect 1462 21988 1738 22030
rect 1862 22070 2138 22112
rect 1862 22030 1980 22070
rect 2020 22030 2138 22070
rect 1862 21988 2138 22030
rect 2262 22070 2538 22112
rect 2262 22030 2380 22070
rect 2420 22030 2538 22070
rect 2262 21988 2538 22030
rect 2662 22070 2938 22112
rect 2662 22030 2780 22070
rect 2820 22030 2938 22070
rect 2662 21988 2938 22030
rect 3062 22070 3338 22112
rect 3062 22030 3180 22070
rect 3220 22030 3338 22070
rect 3062 21988 3338 22030
rect 3462 22070 3738 22112
rect 3462 22030 3580 22070
rect 3620 22030 3738 22070
rect 3462 21988 3738 22030
rect 3862 22070 4138 22112
rect 3862 22030 3980 22070
rect 4020 22030 4138 22070
rect 3862 21988 4138 22030
rect 4262 22070 4538 22112
rect 4262 22030 4380 22070
rect 4420 22030 4538 22070
rect 4262 21988 4538 22030
rect 4662 22070 4938 22112
rect 4662 22030 4780 22070
rect 4820 22030 4938 22070
rect 4662 21988 4938 22030
rect 5062 22070 5338 22112
rect 5062 22030 5180 22070
rect 5220 22030 5338 22070
rect 5062 21988 5338 22030
rect 5462 22070 5738 22112
rect 5462 22030 5580 22070
rect 5620 22030 5738 22070
rect 5462 21988 5738 22030
rect 5862 22070 6138 22112
rect 5862 22030 5980 22070
rect 6020 22030 6138 22070
rect 5862 21988 6138 22030
rect 6262 22070 6538 22112
rect 6262 22030 6380 22070
rect 6420 22030 6538 22070
rect 6262 21988 6538 22030
rect 6662 22070 6938 22112
rect 6662 22030 6780 22070
rect 6820 22030 6938 22070
rect 6662 21988 6938 22030
rect 7062 22070 7338 22112
rect 7062 22030 7180 22070
rect 7220 22030 7338 22070
rect 7062 21988 7338 22030
rect 7462 22070 7738 22112
rect 7462 22030 7580 22070
rect 7620 22030 7738 22070
rect 7462 21988 7738 22030
rect 7862 22070 8138 22112
rect 7862 22030 7980 22070
rect 8020 22030 8138 22070
rect 7862 21988 8138 22030
rect 8262 22070 8538 22112
rect 8262 22030 8380 22070
rect 8420 22030 8538 22070
rect 8262 21988 8538 22030
rect 8662 22070 8938 22112
rect 8662 22030 8780 22070
rect 8820 22030 8938 22070
rect 8662 21988 8938 22030
rect 9062 22070 9338 22112
rect 9062 22030 9180 22070
rect 9220 22030 9338 22070
rect 9062 21988 9338 22030
rect 9462 22070 9738 22112
rect 9462 22030 9580 22070
rect 9620 22030 9738 22070
rect 9462 21988 9738 22030
rect 9862 22070 10138 22112
rect 9862 22030 9980 22070
rect 10020 22030 10138 22070
rect 9862 21988 10138 22030
rect 10262 22070 10538 22112
rect 10262 22030 10380 22070
rect 10420 22030 10538 22070
rect 10262 21988 10538 22030
rect 10662 22070 10938 22112
rect 10662 22030 10780 22070
rect 10820 22030 10938 22070
rect 10662 21988 10938 22030
rect 11062 22070 11338 22112
rect 11062 22030 11180 22070
rect 11220 22030 11338 22070
rect 11062 21988 11338 22030
rect 11462 22070 11738 22112
rect 11462 22030 11580 22070
rect 11620 22030 11738 22070
rect 11462 21988 11738 22030
rect 11862 22070 12138 22112
rect 11862 22030 11980 22070
rect 12020 22030 12138 22070
rect 11862 21988 12138 22030
rect 12262 22070 12538 22112
rect 12262 22030 12380 22070
rect 12420 22030 12538 22070
rect 12262 21988 12538 22030
rect 12662 22070 12938 22112
rect 12662 22030 12780 22070
rect 12820 22030 12938 22070
rect 12662 21988 12938 22030
rect 13062 22070 13338 22112
rect 13062 22030 13180 22070
rect 13220 22030 13338 22070
rect 13062 21988 13338 22030
rect 13462 22070 13738 22112
rect 13462 22030 13580 22070
rect 13620 22030 13738 22070
rect 13462 21988 13738 22030
rect 13862 22070 14138 22112
rect 13862 22030 13980 22070
rect 14020 22030 14138 22070
rect 13862 21988 14138 22030
rect 14262 22070 14538 22112
rect 14262 22030 14380 22070
rect 14420 22030 14538 22070
rect 14262 21988 14538 22030
rect 14662 22070 14938 22112
rect 14662 22030 14780 22070
rect 14820 22030 14938 22070
rect 14662 21988 14938 22030
rect 15062 22070 15338 22112
rect 15062 22030 15180 22070
rect 15220 22030 15338 22070
rect 15062 21988 15338 22030
rect 15462 22070 16000 22112
rect 15462 22030 15580 22070
rect 15620 22030 16000 22070
rect 15462 21988 16000 22030
rect 0 21712 16000 21988
rect 0 21670 538 21712
rect 0 21630 380 21670
rect 420 21630 538 21670
rect 0 21588 538 21630
rect 662 21670 938 21712
rect 662 21630 780 21670
rect 820 21630 938 21670
rect 662 21588 938 21630
rect 1062 21670 1338 21712
rect 1062 21630 1180 21670
rect 1220 21630 1338 21670
rect 1062 21588 1338 21630
rect 1462 21670 1738 21712
rect 1462 21630 1580 21670
rect 1620 21630 1738 21670
rect 1462 21588 1738 21630
rect 1862 21670 2138 21712
rect 1862 21630 1980 21670
rect 2020 21630 2138 21670
rect 1862 21588 2138 21630
rect 2262 21670 2538 21712
rect 2262 21630 2380 21670
rect 2420 21630 2538 21670
rect 2262 21588 2538 21630
rect 2662 21670 2938 21712
rect 2662 21630 2780 21670
rect 2820 21630 2938 21670
rect 2662 21588 2938 21630
rect 3062 21670 3338 21712
rect 3062 21630 3180 21670
rect 3220 21630 3338 21670
rect 3062 21588 3338 21630
rect 3462 21670 3738 21712
rect 3462 21630 3580 21670
rect 3620 21630 3738 21670
rect 3462 21588 3738 21630
rect 3862 21670 4138 21712
rect 3862 21630 3980 21670
rect 4020 21630 4138 21670
rect 3862 21588 4138 21630
rect 4262 21670 4538 21712
rect 4262 21630 4380 21670
rect 4420 21630 4538 21670
rect 4262 21588 4538 21630
rect 4662 21670 4938 21712
rect 4662 21630 4780 21670
rect 4820 21630 4938 21670
rect 4662 21588 4938 21630
rect 5062 21670 5338 21712
rect 5062 21630 5180 21670
rect 5220 21630 5338 21670
rect 5062 21588 5338 21630
rect 5462 21670 5738 21712
rect 5462 21630 5580 21670
rect 5620 21630 5738 21670
rect 5462 21588 5738 21630
rect 5862 21670 6138 21712
rect 5862 21630 5980 21670
rect 6020 21630 6138 21670
rect 5862 21588 6138 21630
rect 6262 21670 6538 21712
rect 6262 21630 6380 21670
rect 6420 21630 6538 21670
rect 6262 21588 6538 21630
rect 6662 21670 6938 21712
rect 6662 21630 6780 21670
rect 6820 21630 6938 21670
rect 6662 21588 6938 21630
rect 7062 21670 7338 21712
rect 7062 21630 7180 21670
rect 7220 21630 7338 21670
rect 7062 21588 7338 21630
rect 7462 21670 7738 21712
rect 7462 21630 7580 21670
rect 7620 21630 7738 21670
rect 7462 21588 7738 21630
rect 7862 21670 8138 21712
rect 7862 21630 7980 21670
rect 8020 21630 8138 21670
rect 7862 21588 8138 21630
rect 8262 21670 8538 21712
rect 8262 21630 8380 21670
rect 8420 21630 8538 21670
rect 8262 21588 8538 21630
rect 8662 21670 8938 21712
rect 8662 21630 8780 21670
rect 8820 21630 8938 21670
rect 8662 21588 8938 21630
rect 9062 21670 9338 21712
rect 9062 21630 9180 21670
rect 9220 21630 9338 21670
rect 9062 21588 9338 21630
rect 9462 21670 9738 21712
rect 9462 21630 9580 21670
rect 9620 21630 9738 21670
rect 9462 21588 9738 21630
rect 9862 21670 10138 21712
rect 9862 21630 9980 21670
rect 10020 21630 10138 21670
rect 9862 21588 10138 21630
rect 10262 21670 10538 21712
rect 10262 21630 10380 21670
rect 10420 21630 10538 21670
rect 10262 21588 10538 21630
rect 10662 21670 10938 21712
rect 10662 21630 10780 21670
rect 10820 21630 10938 21670
rect 10662 21588 10938 21630
rect 11062 21670 11338 21712
rect 11062 21630 11180 21670
rect 11220 21630 11338 21670
rect 11062 21588 11338 21630
rect 11462 21670 11738 21712
rect 11462 21630 11580 21670
rect 11620 21630 11738 21670
rect 11462 21588 11738 21630
rect 11862 21670 12138 21712
rect 11862 21630 11980 21670
rect 12020 21630 12138 21670
rect 11862 21588 12138 21630
rect 12262 21670 12538 21712
rect 12262 21630 12380 21670
rect 12420 21630 12538 21670
rect 12262 21588 12538 21630
rect 12662 21670 12938 21712
rect 12662 21630 12780 21670
rect 12820 21630 12938 21670
rect 12662 21588 12938 21630
rect 13062 21670 13338 21712
rect 13062 21630 13180 21670
rect 13220 21630 13338 21670
rect 13062 21588 13338 21630
rect 13462 21670 13738 21712
rect 13462 21630 13580 21670
rect 13620 21630 13738 21670
rect 13462 21588 13738 21630
rect 13862 21670 14138 21712
rect 13862 21630 13980 21670
rect 14020 21630 14138 21670
rect 13862 21588 14138 21630
rect 14262 21670 14538 21712
rect 14262 21630 14380 21670
rect 14420 21630 14538 21670
rect 14262 21588 14538 21630
rect 14662 21670 14938 21712
rect 14662 21630 14780 21670
rect 14820 21630 14938 21670
rect 14662 21588 14938 21630
rect 15062 21670 15338 21712
rect 15062 21630 15180 21670
rect 15220 21630 15338 21670
rect 15062 21588 15338 21630
rect 15462 21670 16000 21712
rect 15462 21630 15580 21670
rect 15620 21630 16000 21670
rect 15462 21588 16000 21630
rect 0 21312 16000 21588
rect 0 21270 538 21312
rect 0 21230 380 21270
rect 420 21230 538 21270
rect 0 21188 538 21230
rect 662 21270 938 21312
rect 662 21230 780 21270
rect 820 21230 938 21270
rect 662 21188 938 21230
rect 1062 21270 1338 21312
rect 1062 21230 1180 21270
rect 1220 21230 1338 21270
rect 1062 21188 1338 21230
rect 1462 21270 1738 21312
rect 1462 21230 1580 21270
rect 1620 21230 1738 21270
rect 1462 21188 1738 21230
rect 1862 21270 2138 21312
rect 1862 21230 1980 21270
rect 2020 21230 2138 21270
rect 1862 21188 2138 21230
rect 2262 21270 2538 21312
rect 2262 21230 2380 21270
rect 2420 21230 2538 21270
rect 2262 21188 2538 21230
rect 2662 21270 2938 21312
rect 2662 21230 2780 21270
rect 2820 21230 2938 21270
rect 2662 21188 2938 21230
rect 3062 21270 3338 21312
rect 3062 21230 3180 21270
rect 3220 21230 3338 21270
rect 3062 21188 3338 21230
rect 3462 21270 3738 21312
rect 3462 21230 3580 21270
rect 3620 21230 3738 21270
rect 3462 21188 3738 21230
rect 3862 21270 4138 21312
rect 3862 21230 3980 21270
rect 4020 21230 4138 21270
rect 3862 21188 4138 21230
rect 4262 21270 4538 21312
rect 4262 21230 4380 21270
rect 4420 21230 4538 21270
rect 4262 21188 4538 21230
rect 4662 21270 4938 21312
rect 4662 21230 4780 21270
rect 4820 21230 4938 21270
rect 4662 21188 4938 21230
rect 5062 21270 5338 21312
rect 5062 21230 5180 21270
rect 5220 21230 5338 21270
rect 5062 21188 5338 21230
rect 5462 21270 5738 21312
rect 5462 21230 5580 21270
rect 5620 21230 5738 21270
rect 5462 21188 5738 21230
rect 5862 21270 6138 21312
rect 5862 21230 5980 21270
rect 6020 21230 6138 21270
rect 5862 21188 6138 21230
rect 6262 21270 6538 21312
rect 6262 21230 6380 21270
rect 6420 21230 6538 21270
rect 6262 21188 6538 21230
rect 6662 21270 6938 21312
rect 6662 21230 6780 21270
rect 6820 21230 6938 21270
rect 6662 21188 6938 21230
rect 7062 21270 7338 21312
rect 7062 21230 7180 21270
rect 7220 21230 7338 21270
rect 7062 21188 7338 21230
rect 7462 21270 7738 21312
rect 7462 21230 7580 21270
rect 7620 21230 7738 21270
rect 7462 21188 7738 21230
rect 7862 21270 8138 21312
rect 7862 21230 7980 21270
rect 8020 21230 8138 21270
rect 7862 21188 8138 21230
rect 8262 21270 8538 21312
rect 8262 21230 8380 21270
rect 8420 21230 8538 21270
rect 8262 21188 8538 21230
rect 8662 21270 8938 21312
rect 8662 21230 8780 21270
rect 8820 21230 8938 21270
rect 8662 21188 8938 21230
rect 9062 21270 9338 21312
rect 9062 21230 9180 21270
rect 9220 21230 9338 21270
rect 9062 21188 9338 21230
rect 9462 21270 9738 21312
rect 9462 21230 9580 21270
rect 9620 21230 9738 21270
rect 9462 21188 9738 21230
rect 9862 21270 10138 21312
rect 9862 21230 9980 21270
rect 10020 21230 10138 21270
rect 9862 21188 10138 21230
rect 10262 21270 10538 21312
rect 10262 21230 10380 21270
rect 10420 21230 10538 21270
rect 10262 21188 10538 21230
rect 10662 21270 10938 21312
rect 10662 21230 10780 21270
rect 10820 21230 10938 21270
rect 10662 21188 10938 21230
rect 11062 21270 11338 21312
rect 11062 21230 11180 21270
rect 11220 21230 11338 21270
rect 11062 21188 11338 21230
rect 11462 21270 11738 21312
rect 11462 21230 11580 21270
rect 11620 21230 11738 21270
rect 11462 21188 11738 21230
rect 11862 21270 12138 21312
rect 11862 21230 11980 21270
rect 12020 21230 12138 21270
rect 11862 21188 12138 21230
rect 12262 21270 12538 21312
rect 12262 21230 12380 21270
rect 12420 21230 12538 21270
rect 12262 21188 12538 21230
rect 12662 21270 12938 21312
rect 12662 21230 12780 21270
rect 12820 21230 12938 21270
rect 12662 21188 12938 21230
rect 13062 21270 13338 21312
rect 13062 21230 13180 21270
rect 13220 21230 13338 21270
rect 13062 21188 13338 21230
rect 13462 21270 13738 21312
rect 13462 21230 13580 21270
rect 13620 21230 13738 21270
rect 13462 21188 13738 21230
rect 13862 21270 14138 21312
rect 13862 21230 13980 21270
rect 14020 21230 14138 21270
rect 13862 21188 14138 21230
rect 14262 21270 14538 21312
rect 14262 21230 14380 21270
rect 14420 21230 14538 21270
rect 14262 21188 14538 21230
rect 14662 21270 14938 21312
rect 14662 21230 14780 21270
rect 14820 21230 14938 21270
rect 14662 21188 14938 21230
rect 15062 21270 15338 21312
rect 15062 21230 15180 21270
rect 15220 21230 15338 21270
rect 15062 21188 15338 21230
rect 15462 21270 16000 21312
rect 15462 21230 15580 21270
rect 15620 21230 16000 21270
rect 15462 21188 16000 21230
rect 0 20912 16000 21188
rect 0 20870 538 20912
rect 0 20830 380 20870
rect 420 20830 538 20870
rect 0 20788 538 20830
rect 662 20870 938 20912
rect 662 20830 780 20870
rect 820 20830 938 20870
rect 662 20788 938 20830
rect 1062 20870 1338 20912
rect 1062 20830 1180 20870
rect 1220 20830 1338 20870
rect 1062 20788 1338 20830
rect 1462 20870 1738 20912
rect 1462 20830 1580 20870
rect 1620 20830 1738 20870
rect 1462 20788 1738 20830
rect 1862 20870 2138 20912
rect 1862 20830 1980 20870
rect 2020 20830 2138 20870
rect 1862 20788 2138 20830
rect 2262 20870 2538 20912
rect 2262 20830 2380 20870
rect 2420 20830 2538 20870
rect 2262 20788 2538 20830
rect 2662 20870 2938 20912
rect 2662 20830 2780 20870
rect 2820 20830 2938 20870
rect 2662 20788 2938 20830
rect 3062 20870 3338 20912
rect 3062 20830 3180 20870
rect 3220 20830 3338 20870
rect 3062 20788 3338 20830
rect 3462 20870 3738 20912
rect 3462 20830 3580 20870
rect 3620 20830 3738 20870
rect 3462 20788 3738 20830
rect 3862 20870 4138 20912
rect 3862 20830 3980 20870
rect 4020 20830 4138 20870
rect 3862 20788 4138 20830
rect 4262 20870 4538 20912
rect 4262 20830 4380 20870
rect 4420 20830 4538 20870
rect 4262 20788 4538 20830
rect 4662 20870 4938 20912
rect 4662 20830 4780 20870
rect 4820 20830 4938 20870
rect 4662 20788 4938 20830
rect 5062 20870 5338 20912
rect 5062 20830 5180 20870
rect 5220 20830 5338 20870
rect 5062 20788 5338 20830
rect 5462 20870 5738 20912
rect 5462 20830 5580 20870
rect 5620 20830 5738 20870
rect 5462 20788 5738 20830
rect 5862 20870 6138 20912
rect 5862 20830 5980 20870
rect 6020 20830 6138 20870
rect 5862 20788 6138 20830
rect 6262 20870 6538 20912
rect 6262 20830 6380 20870
rect 6420 20830 6538 20870
rect 6262 20788 6538 20830
rect 6662 20870 6938 20912
rect 6662 20830 6780 20870
rect 6820 20830 6938 20870
rect 6662 20788 6938 20830
rect 7062 20870 7338 20912
rect 7062 20830 7180 20870
rect 7220 20830 7338 20870
rect 7062 20788 7338 20830
rect 7462 20870 7738 20912
rect 7462 20830 7580 20870
rect 7620 20830 7738 20870
rect 7462 20788 7738 20830
rect 7862 20870 8138 20912
rect 7862 20830 7980 20870
rect 8020 20830 8138 20870
rect 7862 20788 8138 20830
rect 8262 20870 8538 20912
rect 8262 20830 8380 20870
rect 8420 20830 8538 20870
rect 8262 20788 8538 20830
rect 8662 20870 8938 20912
rect 8662 20830 8780 20870
rect 8820 20830 8938 20870
rect 8662 20788 8938 20830
rect 9062 20870 9338 20912
rect 9062 20830 9180 20870
rect 9220 20830 9338 20870
rect 9062 20788 9338 20830
rect 9462 20870 9738 20912
rect 9462 20830 9580 20870
rect 9620 20830 9738 20870
rect 9462 20788 9738 20830
rect 9862 20870 10138 20912
rect 9862 20830 9980 20870
rect 10020 20830 10138 20870
rect 9862 20788 10138 20830
rect 10262 20870 10538 20912
rect 10262 20830 10380 20870
rect 10420 20830 10538 20870
rect 10262 20788 10538 20830
rect 10662 20870 10938 20912
rect 10662 20830 10780 20870
rect 10820 20830 10938 20870
rect 10662 20788 10938 20830
rect 11062 20870 11338 20912
rect 11062 20830 11180 20870
rect 11220 20830 11338 20870
rect 11062 20788 11338 20830
rect 11462 20870 11738 20912
rect 11462 20830 11580 20870
rect 11620 20830 11738 20870
rect 11462 20788 11738 20830
rect 11862 20870 12138 20912
rect 11862 20830 11980 20870
rect 12020 20830 12138 20870
rect 11862 20788 12138 20830
rect 12262 20870 12538 20912
rect 12262 20830 12380 20870
rect 12420 20830 12538 20870
rect 12262 20788 12538 20830
rect 12662 20870 12938 20912
rect 12662 20830 12780 20870
rect 12820 20830 12938 20870
rect 12662 20788 12938 20830
rect 13062 20870 13338 20912
rect 13062 20830 13180 20870
rect 13220 20830 13338 20870
rect 13062 20788 13338 20830
rect 13462 20870 13738 20912
rect 13462 20830 13580 20870
rect 13620 20830 13738 20870
rect 13462 20788 13738 20830
rect 13862 20870 14138 20912
rect 13862 20830 13980 20870
rect 14020 20830 14138 20870
rect 13862 20788 14138 20830
rect 14262 20870 14538 20912
rect 14262 20830 14380 20870
rect 14420 20830 14538 20870
rect 14262 20788 14538 20830
rect 14662 20870 14938 20912
rect 14662 20830 14780 20870
rect 14820 20830 14938 20870
rect 14662 20788 14938 20830
rect 15062 20870 15338 20912
rect 15062 20830 15180 20870
rect 15220 20830 15338 20870
rect 15062 20788 15338 20830
rect 15462 20870 16000 20912
rect 15462 20830 15580 20870
rect 15620 20830 16000 20870
rect 15462 20788 16000 20830
rect 0 20512 16000 20788
rect 0 20470 538 20512
rect 0 20430 380 20470
rect 420 20430 538 20470
rect 0 20388 538 20430
rect 662 20470 938 20512
rect 662 20430 780 20470
rect 820 20430 938 20470
rect 662 20388 938 20430
rect 1062 20470 1338 20512
rect 1062 20430 1180 20470
rect 1220 20430 1338 20470
rect 1062 20388 1338 20430
rect 1462 20470 1738 20512
rect 1462 20430 1580 20470
rect 1620 20430 1738 20470
rect 1462 20388 1738 20430
rect 1862 20470 2138 20512
rect 1862 20430 1980 20470
rect 2020 20430 2138 20470
rect 1862 20388 2138 20430
rect 2262 20470 2538 20512
rect 2262 20430 2380 20470
rect 2420 20430 2538 20470
rect 2262 20388 2538 20430
rect 2662 20470 2938 20512
rect 2662 20430 2780 20470
rect 2820 20430 2938 20470
rect 2662 20388 2938 20430
rect 3062 20470 3338 20512
rect 3062 20430 3180 20470
rect 3220 20430 3338 20470
rect 3062 20388 3338 20430
rect 3462 20470 3738 20512
rect 3462 20430 3580 20470
rect 3620 20430 3738 20470
rect 3462 20388 3738 20430
rect 3862 20470 4138 20512
rect 3862 20430 3980 20470
rect 4020 20430 4138 20470
rect 3862 20388 4138 20430
rect 4262 20470 4538 20512
rect 4262 20430 4380 20470
rect 4420 20430 4538 20470
rect 4262 20388 4538 20430
rect 4662 20470 4938 20512
rect 4662 20430 4780 20470
rect 4820 20430 4938 20470
rect 4662 20388 4938 20430
rect 5062 20470 5338 20512
rect 5062 20430 5180 20470
rect 5220 20430 5338 20470
rect 5062 20388 5338 20430
rect 5462 20470 5738 20512
rect 5462 20430 5580 20470
rect 5620 20430 5738 20470
rect 5462 20388 5738 20430
rect 5862 20470 6138 20512
rect 5862 20430 5980 20470
rect 6020 20430 6138 20470
rect 5862 20388 6138 20430
rect 6262 20470 6538 20512
rect 6262 20430 6380 20470
rect 6420 20430 6538 20470
rect 6262 20388 6538 20430
rect 6662 20470 6938 20512
rect 6662 20430 6780 20470
rect 6820 20430 6938 20470
rect 6662 20388 6938 20430
rect 7062 20470 7338 20512
rect 7062 20430 7180 20470
rect 7220 20430 7338 20470
rect 7062 20388 7338 20430
rect 7462 20470 7738 20512
rect 7462 20430 7580 20470
rect 7620 20430 7738 20470
rect 7462 20388 7738 20430
rect 7862 20470 8138 20512
rect 7862 20430 7980 20470
rect 8020 20430 8138 20470
rect 7862 20388 8138 20430
rect 8262 20470 8538 20512
rect 8262 20430 8380 20470
rect 8420 20430 8538 20470
rect 8262 20388 8538 20430
rect 8662 20470 8938 20512
rect 8662 20430 8780 20470
rect 8820 20430 8938 20470
rect 8662 20388 8938 20430
rect 9062 20470 9338 20512
rect 9062 20430 9180 20470
rect 9220 20430 9338 20470
rect 9062 20388 9338 20430
rect 9462 20470 9738 20512
rect 9462 20430 9580 20470
rect 9620 20430 9738 20470
rect 9462 20388 9738 20430
rect 9862 20470 10138 20512
rect 9862 20430 9980 20470
rect 10020 20430 10138 20470
rect 9862 20388 10138 20430
rect 10262 20470 10538 20512
rect 10262 20430 10380 20470
rect 10420 20430 10538 20470
rect 10262 20388 10538 20430
rect 10662 20470 10938 20512
rect 10662 20430 10780 20470
rect 10820 20430 10938 20470
rect 10662 20388 10938 20430
rect 11062 20470 11338 20512
rect 11062 20430 11180 20470
rect 11220 20430 11338 20470
rect 11062 20388 11338 20430
rect 11462 20470 11738 20512
rect 11462 20430 11580 20470
rect 11620 20430 11738 20470
rect 11462 20388 11738 20430
rect 11862 20470 12138 20512
rect 11862 20430 11980 20470
rect 12020 20430 12138 20470
rect 11862 20388 12138 20430
rect 12262 20470 12538 20512
rect 12262 20430 12380 20470
rect 12420 20430 12538 20470
rect 12262 20388 12538 20430
rect 12662 20470 12938 20512
rect 12662 20430 12780 20470
rect 12820 20430 12938 20470
rect 12662 20388 12938 20430
rect 13062 20470 13338 20512
rect 13062 20430 13180 20470
rect 13220 20430 13338 20470
rect 13062 20388 13338 20430
rect 13462 20470 13738 20512
rect 13462 20430 13580 20470
rect 13620 20430 13738 20470
rect 13462 20388 13738 20430
rect 13862 20470 14138 20512
rect 13862 20430 13980 20470
rect 14020 20430 14138 20470
rect 13862 20388 14138 20430
rect 14262 20470 14538 20512
rect 14262 20430 14380 20470
rect 14420 20430 14538 20470
rect 14262 20388 14538 20430
rect 14662 20470 14938 20512
rect 14662 20430 14780 20470
rect 14820 20430 14938 20470
rect 14662 20388 14938 20430
rect 15062 20470 15338 20512
rect 15062 20430 15180 20470
rect 15220 20430 15338 20470
rect 15062 20388 15338 20430
rect 15462 20470 16000 20512
rect 15462 20430 15580 20470
rect 15620 20430 16000 20470
rect 15462 20388 16000 20430
rect 0 20112 16000 20388
rect 0 20070 538 20112
rect 0 20030 380 20070
rect 420 20030 538 20070
rect 0 19988 538 20030
rect 662 20070 938 20112
rect 662 20030 780 20070
rect 820 20030 938 20070
rect 662 19988 938 20030
rect 1062 20070 1338 20112
rect 1062 20030 1180 20070
rect 1220 20030 1338 20070
rect 1062 19988 1338 20030
rect 1462 20070 1738 20112
rect 1462 20030 1580 20070
rect 1620 20030 1738 20070
rect 1462 19988 1738 20030
rect 1862 20070 2138 20112
rect 1862 20030 1980 20070
rect 2020 20030 2138 20070
rect 1862 19988 2138 20030
rect 2262 20070 2538 20112
rect 2262 20030 2380 20070
rect 2420 20030 2538 20070
rect 2262 19988 2538 20030
rect 2662 20070 2938 20112
rect 2662 20030 2780 20070
rect 2820 20030 2938 20070
rect 2662 19988 2938 20030
rect 3062 20070 3338 20112
rect 3062 20030 3180 20070
rect 3220 20030 3338 20070
rect 3062 19988 3338 20030
rect 3462 20070 3738 20112
rect 3462 20030 3580 20070
rect 3620 20030 3738 20070
rect 3462 19988 3738 20030
rect 3862 20070 4138 20112
rect 3862 20030 3980 20070
rect 4020 20030 4138 20070
rect 3862 19988 4138 20030
rect 4262 20070 4538 20112
rect 4262 20030 4380 20070
rect 4420 20030 4538 20070
rect 4262 19988 4538 20030
rect 4662 20070 4938 20112
rect 4662 20030 4780 20070
rect 4820 20030 4938 20070
rect 4662 19988 4938 20030
rect 5062 20070 5338 20112
rect 5062 20030 5180 20070
rect 5220 20030 5338 20070
rect 5062 19988 5338 20030
rect 5462 20070 5738 20112
rect 5462 20030 5580 20070
rect 5620 20030 5738 20070
rect 5462 19988 5738 20030
rect 5862 20070 6138 20112
rect 5862 20030 5980 20070
rect 6020 20030 6138 20070
rect 5862 19988 6138 20030
rect 6262 20070 6538 20112
rect 6262 20030 6380 20070
rect 6420 20030 6538 20070
rect 6262 19988 6538 20030
rect 6662 20070 6938 20112
rect 6662 20030 6780 20070
rect 6820 20030 6938 20070
rect 6662 19988 6938 20030
rect 7062 20070 7338 20112
rect 7062 20030 7180 20070
rect 7220 20030 7338 20070
rect 7062 19988 7338 20030
rect 7462 20070 7738 20112
rect 7462 20030 7580 20070
rect 7620 20030 7738 20070
rect 7462 19988 7738 20030
rect 7862 20070 8138 20112
rect 7862 20030 7980 20070
rect 8020 20030 8138 20070
rect 7862 19988 8138 20030
rect 8262 20070 8538 20112
rect 8262 20030 8380 20070
rect 8420 20030 8538 20070
rect 8262 19988 8538 20030
rect 8662 20070 8938 20112
rect 8662 20030 8780 20070
rect 8820 20030 8938 20070
rect 8662 19988 8938 20030
rect 9062 20070 9338 20112
rect 9062 20030 9180 20070
rect 9220 20030 9338 20070
rect 9062 19988 9338 20030
rect 9462 20070 9738 20112
rect 9462 20030 9580 20070
rect 9620 20030 9738 20070
rect 9462 19988 9738 20030
rect 9862 20070 10138 20112
rect 9862 20030 9980 20070
rect 10020 20030 10138 20070
rect 9862 19988 10138 20030
rect 10262 20070 10538 20112
rect 10262 20030 10380 20070
rect 10420 20030 10538 20070
rect 10262 19988 10538 20030
rect 10662 20070 10938 20112
rect 10662 20030 10780 20070
rect 10820 20030 10938 20070
rect 10662 19988 10938 20030
rect 11062 20070 11338 20112
rect 11062 20030 11180 20070
rect 11220 20030 11338 20070
rect 11062 19988 11338 20030
rect 11462 20070 11738 20112
rect 11462 20030 11580 20070
rect 11620 20030 11738 20070
rect 11462 19988 11738 20030
rect 11862 20070 12138 20112
rect 11862 20030 11980 20070
rect 12020 20030 12138 20070
rect 11862 19988 12138 20030
rect 12262 20070 12538 20112
rect 12262 20030 12380 20070
rect 12420 20030 12538 20070
rect 12262 19988 12538 20030
rect 12662 20070 12938 20112
rect 12662 20030 12780 20070
rect 12820 20030 12938 20070
rect 12662 19988 12938 20030
rect 13062 20070 13338 20112
rect 13062 20030 13180 20070
rect 13220 20030 13338 20070
rect 13062 19988 13338 20030
rect 13462 20070 13738 20112
rect 13462 20030 13580 20070
rect 13620 20030 13738 20070
rect 13462 19988 13738 20030
rect 13862 20070 14138 20112
rect 13862 20030 13980 20070
rect 14020 20030 14138 20070
rect 13862 19988 14138 20030
rect 14262 20070 14538 20112
rect 14262 20030 14380 20070
rect 14420 20030 14538 20070
rect 14262 19988 14538 20030
rect 14662 20070 14938 20112
rect 14662 20030 14780 20070
rect 14820 20030 14938 20070
rect 14662 19988 14938 20030
rect 15062 20070 15338 20112
rect 15062 20030 15180 20070
rect 15220 20030 15338 20070
rect 15062 19988 15338 20030
rect 15462 20070 16000 20112
rect 15462 20030 15580 20070
rect 15620 20030 16000 20070
rect 15462 19988 16000 20030
rect 0 19712 16000 19988
rect 0 19670 538 19712
rect 0 19630 380 19670
rect 420 19630 538 19670
rect 0 19588 538 19630
rect 662 19670 938 19712
rect 662 19630 780 19670
rect 820 19630 938 19670
rect 662 19588 938 19630
rect 1062 19670 1338 19712
rect 1062 19630 1180 19670
rect 1220 19630 1338 19670
rect 1062 19588 1338 19630
rect 1462 19670 1738 19712
rect 1462 19630 1580 19670
rect 1620 19630 1738 19670
rect 1462 19588 1738 19630
rect 1862 19670 2138 19712
rect 1862 19630 1980 19670
rect 2020 19630 2138 19670
rect 1862 19588 2138 19630
rect 2262 19670 2538 19712
rect 2262 19630 2380 19670
rect 2420 19630 2538 19670
rect 2262 19588 2538 19630
rect 2662 19670 2938 19712
rect 2662 19630 2780 19670
rect 2820 19630 2938 19670
rect 2662 19588 2938 19630
rect 3062 19670 3338 19712
rect 3062 19630 3180 19670
rect 3220 19630 3338 19670
rect 3062 19588 3338 19630
rect 3462 19670 3738 19712
rect 3462 19630 3580 19670
rect 3620 19630 3738 19670
rect 3462 19588 3738 19630
rect 3862 19670 4138 19712
rect 3862 19630 3980 19670
rect 4020 19630 4138 19670
rect 3862 19588 4138 19630
rect 4262 19670 4538 19712
rect 4262 19630 4380 19670
rect 4420 19630 4538 19670
rect 4262 19588 4538 19630
rect 4662 19670 4938 19712
rect 4662 19630 4780 19670
rect 4820 19630 4938 19670
rect 4662 19588 4938 19630
rect 5062 19670 5338 19712
rect 5062 19630 5180 19670
rect 5220 19630 5338 19670
rect 5062 19588 5338 19630
rect 5462 19670 5738 19712
rect 5462 19630 5580 19670
rect 5620 19630 5738 19670
rect 5462 19588 5738 19630
rect 5862 19670 6138 19712
rect 5862 19630 5980 19670
rect 6020 19630 6138 19670
rect 5862 19588 6138 19630
rect 6262 19670 6538 19712
rect 6262 19630 6380 19670
rect 6420 19630 6538 19670
rect 6262 19588 6538 19630
rect 6662 19670 6938 19712
rect 6662 19630 6780 19670
rect 6820 19630 6938 19670
rect 6662 19588 6938 19630
rect 7062 19670 7338 19712
rect 7062 19630 7180 19670
rect 7220 19630 7338 19670
rect 7062 19588 7338 19630
rect 7462 19670 7738 19712
rect 7462 19630 7580 19670
rect 7620 19630 7738 19670
rect 7462 19588 7738 19630
rect 7862 19670 8138 19712
rect 7862 19630 7980 19670
rect 8020 19630 8138 19670
rect 7862 19588 8138 19630
rect 8262 19670 8538 19712
rect 8262 19630 8380 19670
rect 8420 19630 8538 19670
rect 8262 19588 8538 19630
rect 8662 19670 8938 19712
rect 8662 19630 8780 19670
rect 8820 19630 8938 19670
rect 8662 19588 8938 19630
rect 9062 19670 9338 19712
rect 9062 19630 9180 19670
rect 9220 19630 9338 19670
rect 9062 19588 9338 19630
rect 9462 19670 9738 19712
rect 9462 19630 9580 19670
rect 9620 19630 9738 19670
rect 9462 19588 9738 19630
rect 9862 19670 10138 19712
rect 9862 19630 9980 19670
rect 10020 19630 10138 19670
rect 9862 19588 10138 19630
rect 10262 19670 10538 19712
rect 10262 19630 10380 19670
rect 10420 19630 10538 19670
rect 10262 19588 10538 19630
rect 10662 19670 10938 19712
rect 10662 19630 10780 19670
rect 10820 19630 10938 19670
rect 10662 19588 10938 19630
rect 11062 19670 11338 19712
rect 11062 19630 11180 19670
rect 11220 19630 11338 19670
rect 11062 19588 11338 19630
rect 11462 19670 11738 19712
rect 11462 19630 11580 19670
rect 11620 19630 11738 19670
rect 11462 19588 11738 19630
rect 11862 19670 12138 19712
rect 11862 19630 11980 19670
rect 12020 19630 12138 19670
rect 11862 19588 12138 19630
rect 12262 19670 12538 19712
rect 12262 19630 12380 19670
rect 12420 19630 12538 19670
rect 12262 19588 12538 19630
rect 12662 19670 12938 19712
rect 12662 19630 12780 19670
rect 12820 19630 12938 19670
rect 12662 19588 12938 19630
rect 13062 19670 13338 19712
rect 13062 19630 13180 19670
rect 13220 19630 13338 19670
rect 13062 19588 13338 19630
rect 13462 19670 13738 19712
rect 13462 19630 13580 19670
rect 13620 19630 13738 19670
rect 13462 19588 13738 19630
rect 13862 19670 14138 19712
rect 13862 19630 13980 19670
rect 14020 19630 14138 19670
rect 13862 19588 14138 19630
rect 14262 19670 14538 19712
rect 14262 19630 14380 19670
rect 14420 19630 14538 19670
rect 14262 19588 14538 19630
rect 14662 19670 14938 19712
rect 14662 19630 14780 19670
rect 14820 19630 14938 19670
rect 14662 19588 14938 19630
rect 15062 19670 15338 19712
rect 15062 19630 15180 19670
rect 15220 19630 15338 19670
rect 15062 19588 15338 19630
rect 15462 19670 16000 19712
rect 15462 19630 15580 19670
rect 15620 19630 16000 19670
rect 15462 19588 16000 19630
rect 0 19312 16000 19588
rect 0 19270 538 19312
rect 0 19230 380 19270
rect 420 19230 538 19270
rect 0 19188 538 19230
rect 662 19270 938 19312
rect 662 19230 780 19270
rect 820 19230 938 19270
rect 662 19188 938 19230
rect 1062 19270 1338 19312
rect 1062 19230 1180 19270
rect 1220 19230 1338 19270
rect 1062 19188 1338 19230
rect 1462 19270 1738 19312
rect 1462 19230 1580 19270
rect 1620 19230 1738 19270
rect 1462 19188 1738 19230
rect 1862 19270 2138 19312
rect 1862 19230 1980 19270
rect 2020 19230 2138 19270
rect 1862 19188 2138 19230
rect 2262 19270 2538 19312
rect 2262 19230 2380 19270
rect 2420 19230 2538 19270
rect 2262 19188 2538 19230
rect 2662 19270 2938 19312
rect 2662 19230 2780 19270
rect 2820 19230 2938 19270
rect 2662 19188 2938 19230
rect 3062 19270 3338 19312
rect 3062 19230 3180 19270
rect 3220 19230 3338 19270
rect 3062 19188 3338 19230
rect 3462 19270 3738 19312
rect 3462 19230 3580 19270
rect 3620 19230 3738 19270
rect 3462 19188 3738 19230
rect 3862 19270 4138 19312
rect 3862 19230 3980 19270
rect 4020 19230 4138 19270
rect 3862 19188 4138 19230
rect 4262 19270 4538 19312
rect 4262 19230 4380 19270
rect 4420 19230 4538 19270
rect 4262 19188 4538 19230
rect 4662 19270 4938 19312
rect 4662 19230 4780 19270
rect 4820 19230 4938 19270
rect 4662 19188 4938 19230
rect 5062 19270 5338 19312
rect 5062 19230 5180 19270
rect 5220 19230 5338 19270
rect 5062 19188 5338 19230
rect 5462 19270 5738 19312
rect 5462 19230 5580 19270
rect 5620 19230 5738 19270
rect 5462 19188 5738 19230
rect 5862 19270 6138 19312
rect 5862 19230 5980 19270
rect 6020 19230 6138 19270
rect 5862 19188 6138 19230
rect 6262 19270 6538 19312
rect 6262 19230 6380 19270
rect 6420 19230 6538 19270
rect 6262 19188 6538 19230
rect 6662 19270 6938 19312
rect 6662 19230 6780 19270
rect 6820 19230 6938 19270
rect 6662 19188 6938 19230
rect 7062 19270 7338 19312
rect 7062 19230 7180 19270
rect 7220 19230 7338 19270
rect 7062 19188 7338 19230
rect 7462 19270 7738 19312
rect 7462 19230 7580 19270
rect 7620 19230 7738 19270
rect 7462 19188 7738 19230
rect 7862 19270 8138 19312
rect 7862 19230 7980 19270
rect 8020 19230 8138 19270
rect 7862 19188 8138 19230
rect 8262 19270 8538 19312
rect 8262 19230 8380 19270
rect 8420 19230 8538 19270
rect 8262 19188 8538 19230
rect 8662 19270 8938 19312
rect 8662 19230 8780 19270
rect 8820 19230 8938 19270
rect 8662 19188 8938 19230
rect 9062 19270 9338 19312
rect 9062 19230 9180 19270
rect 9220 19230 9338 19270
rect 9062 19188 9338 19230
rect 9462 19270 9738 19312
rect 9462 19230 9580 19270
rect 9620 19230 9738 19270
rect 9462 19188 9738 19230
rect 9862 19270 10138 19312
rect 9862 19230 9980 19270
rect 10020 19230 10138 19270
rect 9862 19188 10138 19230
rect 10262 19270 10538 19312
rect 10262 19230 10380 19270
rect 10420 19230 10538 19270
rect 10262 19188 10538 19230
rect 10662 19270 10938 19312
rect 10662 19230 10780 19270
rect 10820 19230 10938 19270
rect 10662 19188 10938 19230
rect 11062 19270 11338 19312
rect 11062 19230 11180 19270
rect 11220 19230 11338 19270
rect 11062 19188 11338 19230
rect 11462 19270 11738 19312
rect 11462 19230 11580 19270
rect 11620 19230 11738 19270
rect 11462 19188 11738 19230
rect 11862 19270 12138 19312
rect 11862 19230 11980 19270
rect 12020 19230 12138 19270
rect 11862 19188 12138 19230
rect 12262 19270 12538 19312
rect 12262 19230 12380 19270
rect 12420 19230 12538 19270
rect 12262 19188 12538 19230
rect 12662 19270 12938 19312
rect 12662 19230 12780 19270
rect 12820 19230 12938 19270
rect 12662 19188 12938 19230
rect 13062 19270 13338 19312
rect 13062 19230 13180 19270
rect 13220 19230 13338 19270
rect 13062 19188 13338 19230
rect 13462 19270 13738 19312
rect 13462 19230 13580 19270
rect 13620 19230 13738 19270
rect 13462 19188 13738 19230
rect 13862 19270 14138 19312
rect 13862 19230 13980 19270
rect 14020 19230 14138 19270
rect 13862 19188 14138 19230
rect 14262 19270 14538 19312
rect 14262 19230 14380 19270
rect 14420 19230 14538 19270
rect 14262 19188 14538 19230
rect 14662 19270 14938 19312
rect 14662 19230 14780 19270
rect 14820 19230 14938 19270
rect 14662 19188 14938 19230
rect 15062 19270 15338 19312
rect 15062 19230 15180 19270
rect 15220 19230 15338 19270
rect 15062 19188 15338 19230
rect 15462 19270 16000 19312
rect 15462 19230 15580 19270
rect 15620 19230 16000 19270
rect 15462 19188 16000 19230
rect 0 18700 16000 19188
rect 0 17812 16000 18300
rect 0 17770 538 17812
rect 0 17730 380 17770
rect 420 17730 538 17770
rect 0 17688 538 17730
rect 662 17770 938 17812
rect 662 17730 780 17770
rect 820 17730 938 17770
rect 662 17688 938 17730
rect 1062 17770 1338 17812
rect 1062 17730 1180 17770
rect 1220 17730 1338 17770
rect 1062 17688 1338 17730
rect 1462 17770 1738 17812
rect 1462 17730 1580 17770
rect 1620 17730 1738 17770
rect 1462 17688 1738 17730
rect 1862 17770 2138 17812
rect 1862 17730 1980 17770
rect 2020 17730 2138 17770
rect 1862 17688 2138 17730
rect 2262 17770 2538 17812
rect 2262 17730 2380 17770
rect 2420 17730 2538 17770
rect 2262 17688 2538 17730
rect 2662 17770 2938 17812
rect 2662 17730 2780 17770
rect 2820 17730 2938 17770
rect 2662 17688 2938 17730
rect 3062 17770 3338 17812
rect 3062 17730 3180 17770
rect 3220 17730 3338 17770
rect 3062 17688 3338 17730
rect 3462 17770 3738 17812
rect 3462 17730 3580 17770
rect 3620 17730 3738 17770
rect 3462 17688 3738 17730
rect 3862 17770 4138 17812
rect 3862 17730 3980 17770
rect 4020 17730 4138 17770
rect 3862 17688 4138 17730
rect 4262 17770 4538 17812
rect 4262 17730 4380 17770
rect 4420 17730 4538 17770
rect 4262 17688 4538 17730
rect 4662 17770 4938 17812
rect 4662 17730 4780 17770
rect 4820 17730 4938 17770
rect 4662 17688 4938 17730
rect 5062 17770 5338 17812
rect 5062 17730 5180 17770
rect 5220 17730 5338 17770
rect 5062 17688 5338 17730
rect 5462 17770 5738 17812
rect 5462 17730 5580 17770
rect 5620 17730 5738 17770
rect 5462 17688 5738 17730
rect 5862 17770 6138 17812
rect 5862 17730 5980 17770
rect 6020 17730 6138 17770
rect 5862 17688 6138 17730
rect 6262 17770 6538 17812
rect 6262 17730 6380 17770
rect 6420 17730 6538 17770
rect 6262 17688 6538 17730
rect 6662 17770 6938 17812
rect 6662 17730 6780 17770
rect 6820 17730 6938 17770
rect 6662 17688 6938 17730
rect 7062 17770 7338 17812
rect 7062 17730 7180 17770
rect 7220 17730 7338 17770
rect 7062 17688 7338 17730
rect 7462 17770 7738 17812
rect 7462 17730 7580 17770
rect 7620 17730 7738 17770
rect 7462 17688 7738 17730
rect 7862 17770 8138 17812
rect 7862 17730 7980 17770
rect 8020 17730 8138 17770
rect 7862 17688 8138 17730
rect 8262 17770 8538 17812
rect 8262 17730 8380 17770
rect 8420 17730 8538 17770
rect 8262 17688 8538 17730
rect 8662 17770 8938 17812
rect 8662 17730 8780 17770
rect 8820 17730 8938 17770
rect 8662 17688 8938 17730
rect 9062 17770 9338 17812
rect 9062 17730 9180 17770
rect 9220 17730 9338 17770
rect 9062 17688 9338 17730
rect 9462 17770 9738 17812
rect 9462 17730 9580 17770
rect 9620 17730 9738 17770
rect 9462 17688 9738 17730
rect 9862 17770 10138 17812
rect 9862 17730 9980 17770
rect 10020 17730 10138 17770
rect 9862 17688 10138 17730
rect 10262 17770 10538 17812
rect 10262 17730 10380 17770
rect 10420 17730 10538 17770
rect 10262 17688 10538 17730
rect 10662 17770 10938 17812
rect 10662 17730 10780 17770
rect 10820 17730 10938 17770
rect 10662 17688 10938 17730
rect 11062 17770 11338 17812
rect 11062 17730 11180 17770
rect 11220 17730 11338 17770
rect 11062 17688 11338 17730
rect 11462 17770 11738 17812
rect 11462 17730 11580 17770
rect 11620 17730 11738 17770
rect 11462 17688 11738 17730
rect 11862 17770 12138 17812
rect 11862 17730 11980 17770
rect 12020 17730 12138 17770
rect 11862 17688 12138 17730
rect 12262 17770 12538 17812
rect 12262 17730 12380 17770
rect 12420 17730 12538 17770
rect 12262 17688 12538 17730
rect 12662 17770 12938 17812
rect 12662 17730 12780 17770
rect 12820 17730 12938 17770
rect 12662 17688 12938 17730
rect 13062 17770 13338 17812
rect 13062 17730 13180 17770
rect 13220 17730 13338 17770
rect 13062 17688 13338 17730
rect 13462 17770 13738 17812
rect 13462 17730 13580 17770
rect 13620 17730 13738 17770
rect 13462 17688 13738 17730
rect 13862 17770 14138 17812
rect 13862 17730 13980 17770
rect 14020 17730 14138 17770
rect 13862 17688 14138 17730
rect 14262 17770 14538 17812
rect 14262 17730 14380 17770
rect 14420 17730 14538 17770
rect 14262 17688 14538 17730
rect 14662 17770 14938 17812
rect 14662 17730 14780 17770
rect 14820 17730 14938 17770
rect 14662 17688 14938 17730
rect 15062 17770 15338 17812
rect 15062 17730 15180 17770
rect 15220 17730 15338 17770
rect 15062 17688 15338 17730
rect 15462 17770 16000 17812
rect 15462 17730 15580 17770
rect 15620 17730 16000 17770
rect 15462 17688 16000 17730
rect 0 17412 16000 17688
rect 0 17370 538 17412
rect 0 17330 380 17370
rect 420 17330 538 17370
rect 0 17288 538 17330
rect 662 17370 938 17412
rect 662 17330 780 17370
rect 820 17330 938 17370
rect 662 17288 938 17330
rect 1062 17370 1338 17412
rect 1062 17330 1180 17370
rect 1220 17330 1338 17370
rect 1062 17288 1338 17330
rect 1462 17370 1738 17412
rect 1462 17330 1580 17370
rect 1620 17330 1738 17370
rect 1462 17288 1738 17330
rect 1862 17370 2138 17412
rect 1862 17330 1980 17370
rect 2020 17330 2138 17370
rect 1862 17288 2138 17330
rect 2262 17370 2538 17412
rect 2262 17330 2380 17370
rect 2420 17330 2538 17370
rect 2262 17288 2538 17330
rect 2662 17370 2938 17412
rect 2662 17330 2780 17370
rect 2820 17330 2938 17370
rect 2662 17288 2938 17330
rect 3062 17370 3338 17412
rect 3062 17330 3180 17370
rect 3220 17330 3338 17370
rect 3062 17288 3338 17330
rect 3462 17370 3738 17412
rect 3462 17330 3580 17370
rect 3620 17330 3738 17370
rect 3462 17288 3738 17330
rect 3862 17370 4138 17412
rect 3862 17330 3980 17370
rect 4020 17330 4138 17370
rect 3862 17288 4138 17330
rect 4262 17370 4538 17412
rect 4262 17330 4380 17370
rect 4420 17330 4538 17370
rect 4262 17288 4538 17330
rect 4662 17370 4938 17412
rect 4662 17330 4780 17370
rect 4820 17330 4938 17370
rect 4662 17288 4938 17330
rect 5062 17370 5338 17412
rect 5062 17330 5180 17370
rect 5220 17330 5338 17370
rect 5062 17288 5338 17330
rect 5462 17370 5738 17412
rect 5462 17330 5580 17370
rect 5620 17330 5738 17370
rect 5462 17288 5738 17330
rect 5862 17370 6138 17412
rect 5862 17330 5980 17370
rect 6020 17330 6138 17370
rect 5862 17288 6138 17330
rect 6262 17370 6538 17412
rect 6262 17330 6380 17370
rect 6420 17330 6538 17370
rect 6262 17288 6538 17330
rect 6662 17370 6938 17412
rect 6662 17330 6780 17370
rect 6820 17330 6938 17370
rect 6662 17288 6938 17330
rect 7062 17370 7338 17412
rect 7062 17330 7180 17370
rect 7220 17330 7338 17370
rect 7062 17288 7338 17330
rect 7462 17370 7738 17412
rect 7462 17330 7580 17370
rect 7620 17330 7738 17370
rect 7462 17288 7738 17330
rect 7862 17370 8138 17412
rect 7862 17330 7980 17370
rect 8020 17330 8138 17370
rect 7862 17288 8138 17330
rect 8262 17370 8538 17412
rect 8262 17330 8380 17370
rect 8420 17330 8538 17370
rect 8262 17288 8538 17330
rect 8662 17370 8938 17412
rect 8662 17330 8780 17370
rect 8820 17330 8938 17370
rect 8662 17288 8938 17330
rect 9062 17370 9338 17412
rect 9062 17330 9180 17370
rect 9220 17330 9338 17370
rect 9062 17288 9338 17330
rect 9462 17370 9738 17412
rect 9462 17330 9580 17370
rect 9620 17330 9738 17370
rect 9462 17288 9738 17330
rect 9862 17370 10138 17412
rect 9862 17330 9980 17370
rect 10020 17330 10138 17370
rect 9862 17288 10138 17330
rect 10262 17370 10538 17412
rect 10262 17330 10380 17370
rect 10420 17330 10538 17370
rect 10262 17288 10538 17330
rect 10662 17370 10938 17412
rect 10662 17330 10780 17370
rect 10820 17330 10938 17370
rect 10662 17288 10938 17330
rect 11062 17370 11338 17412
rect 11062 17330 11180 17370
rect 11220 17330 11338 17370
rect 11062 17288 11338 17330
rect 11462 17370 11738 17412
rect 11462 17330 11580 17370
rect 11620 17330 11738 17370
rect 11462 17288 11738 17330
rect 11862 17370 12138 17412
rect 11862 17330 11980 17370
rect 12020 17330 12138 17370
rect 11862 17288 12138 17330
rect 12262 17370 12538 17412
rect 12262 17330 12380 17370
rect 12420 17330 12538 17370
rect 12262 17288 12538 17330
rect 12662 17370 12938 17412
rect 12662 17330 12780 17370
rect 12820 17330 12938 17370
rect 12662 17288 12938 17330
rect 13062 17370 13338 17412
rect 13062 17330 13180 17370
rect 13220 17330 13338 17370
rect 13062 17288 13338 17330
rect 13462 17370 13738 17412
rect 13462 17330 13580 17370
rect 13620 17330 13738 17370
rect 13462 17288 13738 17330
rect 13862 17370 14138 17412
rect 13862 17330 13980 17370
rect 14020 17330 14138 17370
rect 13862 17288 14138 17330
rect 14262 17370 14538 17412
rect 14262 17330 14380 17370
rect 14420 17330 14538 17370
rect 14262 17288 14538 17330
rect 14662 17370 14938 17412
rect 14662 17330 14780 17370
rect 14820 17330 14938 17370
rect 14662 17288 14938 17330
rect 15062 17370 15338 17412
rect 15062 17330 15180 17370
rect 15220 17330 15338 17370
rect 15062 17288 15338 17330
rect 15462 17370 16000 17412
rect 15462 17330 15580 17370
rect 15620 17330 16000 17370
rect 15462 17288 16000 17330
rect 0 17012 16000 17288
rect 0 16970 538 17012
rect 0 16930 380 16970
rect 420 16930 538 16970
rect 0 16888 538 16930
rect 662 16970 938 17012
rect 662 16930 780 16970
rect 820 16930 938 16970
rect 662 16888 938 16930
rect 1062 16970 1338 17012
rect 1062 16930 1180 16970
rect 1220 16930 1338 16970
rect 1062 16888 1338 16930
rect 1462 16970 1738 17012
rect 1462 16930 1580 16970
rect 1620 16930 1738 16970
rect 1462 16888 1738 16930
rect 1862 16970 2138 17012
rect 1862 16930 1980 16970
rect 2020 16930 2138 16970
rect 1862 16888 2138 16930
rect 2262 16970 2538 17012
rect 2262 16930 2380 16970
rect 2420 16930 2538 16970
rect 2262 16888 2538 16930
rect 2662 16970 2938 17012
rect 2662 16930 2780 16970
rect 2820 16930 2938 16970
rect 2662 16888 2938 16930
rect 3062 16970 3338 17012
rect 3062 16930 3180 16970
rect 3220 16930 3338 16970
rect 3062 16888 3338 16930
rect 3462 16970 3738 17012
rect 3462 16930 3580 16970
rect 3620 16930 3738 16970
rect 3462 16888 3738 16930
rect 3862 16970 4138 17012
rect 3862 16930 3980 16970
rect 4020 16930 4138 16970
rect 3862 16888 4138 16930
rect 4262 16970 4538 17012
rect 4262 16930 4380 16970
rect 4420 16930 4538 16970
rect 4262 16888 4538 16930
rect 4662 16970 4938 17012
rect 4662 16930 4780 16970
rect 4820 16930 4938 16970
rect 4662 16888 4938 16930
rect 5062 16970 5338 17012
rect 5062 16930 5180 16970
rect 5220 16930 5338 16970
rect 5062 16888 5338 16930
rect 5462 16970 5738 17012
rect 5462 16930 5580 16970
rect 5620 16930 5738 16970
rect 5462 16888 5738 16930
rect 5862 16970 6138 17012
rect 5862 16930 5980 16970
rect 6020 16930 6138 16970
rect 5862 16888 6138 16930
rect 6262 16970 6538 17012
rect 6262 16930 6380 16970
rect 6420 16930 6538 16970
rect 6262 16888 6538 16930
rect 6662 16970 6938 17012
rect 6662 16930 6780 16970
rect 6820 16930 6938 16970
rect 6662 16888 6938 16930
rect 7062 16970 7338 17012
rect 7062 16930 7180 16970
rect 7220 16930 7338 16970
rect 7062 16888 7338 16930
rect 7462 16970 7738 17012
rect 7462 16930 7580 16970
rect 7620 16930 7738 16970
rect 7462 16888 7738 16930
rect 7862 16970 8138 17012
rect 7862 16930 7980 16970
rect 8020 16930 8138 16970
rect 7862 16888 8138 16930
rect 8262 16970 8538 17012
rect 8262 16930 8380 16970
rect 8420 16930 8538 16970
rect 8262 16888 8538 16930
rect 8662 16970 8938 17012
rect 8662 16930 8780 16970
rect 8820 16930 8938 16970
rect 8662 16888 8938 16930
rect 9062 16970 9338 17012
rect 9062 16930 9180 16970
rect 9220 16930 9338 16970
rect 9062 16888 9338 16930
rect 9462 16970 9738 17012
rect 9462 16930 9580 16970
rect 9620 16930 9738 16970
rect 9462 16888 9738 16930
rect 9862 16970 10138 17012
rect 9862 16930 9980 16970
rect 10020 16930 10138 16970
rect 9862 16888 10138 16930
rect 10262 16970 10538 17012
rect 10262 16930 10380 16970
rect 10420 16930 10538 16970
rect 10262 16888 10538 16930
rect 10662 16970 10938 17012
rect 10662 16930 10780 16970
rect 10820 16930 10938 16970
rect 10662 16888 10938 16930
rect 11062 16970 11338 17012
rect 11062 16930 11180 16970
rect 11220 16930 11338 16970
rect 11062 16888 11338 16930
rect 11462 16970 11738 17012
rect 11462 16930 11580 16970
rect 11620 16930 11738 16970
rect 11462 16888 11738 16930
rect 11862 16970 12138 17012
rect 11862 16930 11980 16970
rect 12020 16930 12138 16970
rect 11862 16888 12138 16930
rect 12262 16970 12538 17012
rect 12262 16930 12380 16970
rect 12420 16930 12538 16970
rect 12262 16888 12538 16930
rect 12662 16970 12938 17012
rect 12662 16930 12780 16970
rect 12820 16930 12938 16970
rect 12662 16888 12938 16930
rect 13062 16970 13338 17012
rect 13062 16930 13180 16970
rect 13220 16930 13338 16970
rect 13062 16888 13338 16930
rect 13462 16970 13738 17012
rect 13462 16930 13580 16970
rect 13620 16930 13738 16970
rect 13462 16888 13738 16930
rect 13862 16970 14138 17012
rect 13862 16930 13980 16970
rect 14020 16930 14138 16970
rect 13862 16888 14138 16930
rect 14262 16970 14538 17012
rect 14262 16930 14380 16970
rect 14420 16930 14538 16970
rect 14262 16888 14538 16930
rect 14662 16970 14938 17012
rect 14662 16930 14780 16970
rect 14820 16930 14938 16970
rect 14662 16888 14938 16930
rect 15062 16970 15338 17012
rect 15062 16930 15180 16970
rect 15220 16930 15338 16970
rect 15062 16888 15338 16930
rect 15462 16970 16000 17012
rect 15462 16930 15580 16970
rect 15620 16930 16000 16970
rect 15462 16888 16000 16930
rect 0 16612 16000 16888
rect 0 16570 538 16612
rect 0 16530 380 16570
rect 420 16530 538 16570
rect 0 16488 538 16530
rect 662 16570 938 16612
rect 662 16530 780 16570
rect 820 16530 938 16570
rect 662 16488 938 16530
rect 1062 16570 1338 16612
rect 1062 16530 1180 16570
rect 1220 16530 1338 16570
rect 1062 16488 1338 16530
rect 1462 16570 1738 16612
rect 1462 16530 1580 16570
rect 1620 16530 1738 16570
rect 1462 16488 1738 16530
rect 1862 16570 2138 16612
rect 1862 16530 1980 16570
rect 2020 16530 2138 16570
rect 1862 16488 2138 16530
rect 2262 16570 2538 16612
rect 2262 16530 2380 16570
rect 2420 16530 2538 16570
rect 2262 16488 2538 16530
rect 2662 16570 2938 16612
rect 2662 16530 2780 16570
rect 2820 16530 2938 16570
rect 2662 16488 2938 16530
rect 3062 16570 3338 16612
rect 3062 16530 3180 16570
rect 3220 16530 3338 16570
rect 3062 16488 3338 16530
rect 3462 16570 3738 16612
rect 3462 16530 3580 16570
rect 3620 16530 3738 16570
rect 3462 16488 3738 16530
rect 3862 16570 4138 16612
rect 3862 16530 3980 16570
rect 4020 16530 4138 16570
rect 3862 16488 4138 16530
rect 4262 16570 4538 16612
rect 4262 16530 4380 16570
rect 4420 16530 4538 16570
rect 4262 16488 4538 16530
rect 4662 16570 4938 16612
rect 4662 16530 4780 16570
rect 4820 16530 4938 16570
rect 4662 16488 4938 16530
rect 5062 16570 5338 16612
rect 5062 16530 5180 16570
rect 5220 16530 5338 16570
rect 5062 16488 5338 16530
rect 5462 16570 5738 16612
rect 5462 16530 5580 16570
rect 5620 16530 5738 16570
rect 5462 16488 5738 16530
rect 5862 16570 6138 16612
rect 5862 16530 5980 16570
rect 6020 16530 6138 16570
rect 5862 16488 6138 16530
rect 6262 16570 6538 16612
rect 6262 16530 6380 16570
rect 6420 16530 6538 16570
rect 6262 16488 6538 16530
rect 6662 16570 6938 16612
rect 6662 16530 6780 16570
rect 6820 16530 6938 16570
rect 6662 16488 6938 16530
rect 7062 16570 7338 16612
rect 7062 16530 7180 16570
rect 7220 16530 7338 16570
rect 7062 16488 7338 16530
rect 7462 16570 7738 16612
rect 7462 16530 7580 16570
rect 7620 16530 7738 16570
rect 7462 16488 7738 16530
rect 7862 16570 8138 16612
rect 7862 16530 7980 16570
rect 8020 16530 8138 16570
rect 7862 16488 8138 16530
rect 8262 16570 8538 16612
rect 8262 16530 8380 16570
rect 8420 16530 8538 16570
rect 8262 16488 8538 16530
rect 8662 16570 8938 16612
rect 8662 16530 8780 16570
rect 8820 16530 8938 16570
rect 8662 16488 8938 16530
rect 9062 16570 9338 16612
rect 9062 16530 9180 16570
rect 9220 16530 9338 16570
rect 9062 16488 9338 16530
rect 9462 16570 9738 16612
rect 9462 16530 9580 16570
rect 9620 16530 9738 16570
rect 9462 16488 9738 16530
rect 9862 16570 10138 16612
rect 9862 16530 9980 16570
rect 10020 16530 10138 16570
rect 9862 16488 10138 16530
rect 10262 16570 10538 16612
rect 10262 16530 10380 16570
rect 10420 16530 10538 16570
rect 10262 16488 10538 16530
rect 10662 16570 10938 16612
rect 10662 16530 10780 16570
rect 10820 16530 10938 16570
rect 10662 16488 10938 16530
rect 11062 16570 11338 16612
rect 11062 16530 11180 16570
rect 11220 16530 11338 16570
rect 11062 16488 11338 16530
rect 11462 16570 11738 16612
rect 11462 16530 11580 16570
rect 11620 16530 11738 16570
rect 11462 16488 11738 16530
rect 11862 16570 12138 16612
rect 11862 16530 11980 16570
rect 12020 16530 12138 16570
rect 11862 16488 12138 16530
rect 12262 16570 12538 16612
rect 12262 16530 12380 16570
rect 12420 16530 12538 16570
rect 12262 16488 12538 16530
rect 12662 16570 12938 16612
rect 12662 16530 12780 16570
rect 12820 16530 12938 16570
rect 12662 16488 12938 16530
rect 13062 16570 13338 16612
rect 13062 16530 13180 16570
rect 13220 16530 13338 16570
rect 13062 16488 13338 16530
rect 13462 16570 13738 16612
rect 13462 16530 13580 16570
rect 13620 16530 13738 16570
rect 13462 16488 13738 16530
rect 13862 16570 14138 16612
rect 13862 16530 13980 16570
rect 14020 16530 14138 16570
rect 13862 16488 14138 16530
rect 14262 16570 14538 16612
rect 14262 16530 14380 16570
rect 14420 16530 14538 16570
rect 14262 16488 14538 16530
rect 14662 16570 14938 16612
rect 14662 16530 14780 16570
rect 14820 16530 14938 16570
rect 14662 16488 14938 16530
rect 15062 16570 15338 16612
rect 15062 16530 15180 16570
rect 15220 16530 15338 16570
rect 15062 16488 15338 16530
rect 15462 16570 16000 16612
rect 15462 16530 15580 16570
rect 15620 16530 16000 16570
rect 15462 16488 16000 16530
rect 0 16212 16000 16488
rect 0 16170 538 16212
rect 0 16130 380 16170
rect 420 16130 538 16170
rect 0 16088 538 16130
rect 662 16170 938 16212
rect 662 16130 780 16170
rect 820 16130 938 16170
rect 662 16088 938 16130
rect 1062 16170 1338 16212
rect 1062 16130 1180 16170
rect 1220 16130 1338 16170
rect 1062 16088 1338 16130
rect 1462 16170 1738 16212
rect 1462 16130 1580 16170
rect 1620 16130 1738 16170
rect 1462 16088 1738 16130
rect 1862 16170 2138 16212
rect 1862 16130 1980 16170
rect 2020 16130 2138 16170
rect 1862 16088 2138 16130
rect 2262 16170 2538 16212
rect 2262 16130 2380 16170
rect 2420 16130 2538 16170
rect 2262 16088 2538 16130
rect 2662 16170 2938 16212
rect 2662 16130 2780 16170
rect 2820 16130 2938 16170
rect 2662 16088 2938 16130
rect 3062 16170 3338 16212
rect 3062 16130 3180 16170
rect 3220 16130 3338 16170
rect 3062 16088 3338 16130
rect 3462 16170 3738 16212
rect 3462 16130 3580 16170
rect 3620 16130 3738 16170
rect 3462 16088 3738 16130
rect 3862 16170 4138 16212
rect 3862 16130 3980 16170
rect 4020 16130 4138 16170
rect 3862 16088 4138 16130
rect 4262 16170 4538 16212
rect 4262 16130 4380 16170
rect 4420 16130 4538 16170
rect 4262 16088 4538 16130
rect 4662 16170 4938 16212
rect 4662 16130 4780 16170
rect 4820 16130 4938 16170
rect 4662 16088 4938 16130
rect 5062 16170 5338 16212
rect 5062 16130 5180 16170
rect 5220 16130 5338 16170
rect 5062 16088 5338 16130
rect 5462 16170 5738 16212
rect 5462 16130 5580 16170
rect 5620 16130 5738 16170
rect 5462 16088 5738 16130
rect 5862 16170 6138 16212
rect 5862 16130 5980 16170
rect 6020 16130 6138 16170
rect 5862 16088 6138 16130
rect 6262 16170 6538 16212
rect 6262 16130 6380 16170
rect 6420 16130 6538 16170
rect 6262 16088 6538 16130
rect 6662 16170 6938 16212
rect 6662 16130 6780 16170
rect 6820 16130 6938 16170
rect 6662 16088 6938 16130
rect 7062 16170 7338 16212
rect 7062 16130 7180 16170
rect 7220 16130 7338 16170
rect 7062 16088 7338 16130
rect 7462 16170 7738 16212
rect 7462 16130 7580 16170
rect 7620 16130 7738 16170
rect 7462 16088 7738 16130
rect 7862 16170 8138 16212
rect 7862 16130 7980 16170
rect 8020 16130 8138 16170
rect 7862 16088 8138 16130
rect 8262 16170 8538 16212
rect 8262 16130 8380 16170
rect 8420 16130 8538 16170
rect 8262 16088 8538 16130
rect 8662 16170 8938 16212
rect 8662 16130 8780 16170
rect 8820 16130 8938 16170
rect 8662 16088 8938 16130
rect 9062 16170 9338 16212
rect 9062 16130 9180 16170
rect 9220 16130 9338 16170
rect 9062 16088 9338 16130
rect 9462 16170 9738 16212
rect 9462 16130 9580 16170
rect 9620 16130 9738 16170
rect 9462 16088 9738 16130
rect 9862 16170 10138 16212
rect 9862 16130 9980 16170
rect 10020 16130 10138 16170
rect 9862 16088 10138 16130
rect 10262 16170 10538 16212
rect 10262 16130 10380 16170
rect 10420 16130 10538 16170
rect 10262 16088 10538 16130
rect 10662 16170 10938 16212
rect 10662 16130 10780 16170
rect 10820 16130 10938 16170
rect 10662 16088 10938 16130
rect 11062 16170 11338 16212
rect 11062 16130 11180 16170
rect 11220 16130 11338 16170
rect 11062 16088 11338 16130
rect 11462 16170 11738 16212
rect 11462 16130 11580 16170
rect 11620 16130 11738 16170
rect 11462 16088 11738 16130
rect 11862 16170 12138 16212
rect 11862 16130 11980 16170
rect 12020 16130 12138 16170
rect 11862 16088 12138 16130
rect 12262 16170 12538 16212
rect 12262 16130 12380 16170
rect 12420 16130 12538 16170
rect 12262 16088 12538 16130
rect 12662 16170 12938 16212
rect 12662 16130 12780 16170
rect 12820 16130 12938 16170
rect 12662 16088 12938 16130
rect 13062 16170 13338 16212
rect 13062 16130 13180 16170
rect 13220 16130 13338 16170
rect 13062 16088 13338 16130
rect 13462 16170 13738 16212
rect 13462 16130 13580 16170
rect 13620 16130 13738 16170
rect 13462 16088 13738 16130
rect 13862 16170 14138 16212
rect 13862 16130 13980 16170
rect 14020 16130 14138 16170
rect 13862 16088 14138 16130
rect 14262 16170 14538 16212
rect 14262 16130 14380 16170
rect 14420 16130 14538 16170
rect 14262 16088 14538 16130
rect 14662 16170 14938 16212
rect 14662 16130 14780 16170
rect 14820 16130 14938 16170
rect 14662 16088 14938 16130
rect 15062 16170 15338 16212
rect 15062 16130 15180 16170
rect 15220 16130 15338 16170
rect 15062 16088 15338 16130
rect 15462 16170 16000 16212
rect 15462 16130 15580 16170
rect 15620 16130 16000 16170
rect 15462 16088 16000 16130
rect 0 15812 16000 16088
rect 0 15770 538 15812
rect 0 15730 380 15770
rect 420 15730 538 15770
rect 0 15688 538 15730
rect 662 15770 938 15812
rect 662 15730 780 15770
rect 820 15730 938 15770
rect 662 15688 938 15730
rect 1062 15770 1338 15812
rect 1062 15730 1180 15770
rect 1220 15730 1338 15770
rect 1062 15688 1338 15730
rect 1462 15770 1738 15812
rect 1462 15730 1580 15770
rect 1620 15730 1738 15770
rect 1462 15688 1738 15730
rect 1862 15770 2138 15812
rect 1862 15730 1980 15770
rect 2020 15730 2138 15770
rect 1862 15688 2138 15730
rect 2262 15770 2538 15812
rect 2262 15730 2380 15770
rect 2420 15730 2538 15770
rect 2262 15688 2538 15730
rect 2662 15770 2938 15812
rect 2662 15730 2780 15770
rect 2820 15730 2938 15770
rect 2662 15688 2938 15730
rect 3062 15770 3338 15812
rect 3062 15730 3180 15770
rect 3220 15730 3338 15770
rect 3062 15688 3338 15730
rect 3462 15770 3738 15812
rect 3462 15730 3580 15770
rect 3620 15730 3738 15770
rect 3462 15688 3738 15730
rect 3862 15770 4138 15812
rect 3862 15730 3980 15770
rect 4020 15730 4138 15770
rect 3862 15688 4138 15730
rect 4262 15770 4538 15812
rect 4262 15730 4380 15770
rect 4420 15730 4538 15770
rect 4262 15688 4538 15730
rect 4662 15770 4938 15812
rect 4662 15730 4780 15770
rect 4820 15730 4938 15770
rect 4662 15688 4938 15730
rect 5062 15770 5338 15812
rect 5062 15730 5180 15770
rect 5220 15730 5338 15770
rect 5062 15688 5338 15730
rect 5462 15770 5738 15812
rect 5462 15730 5580 15770
rect 5620 15730 5738 15770
rect 5462 15688 5738 15730
rect 5862 15770 6138 15812
rect 5862 15730 5980 15770
rect 6020 15730 6138 15770
rect 5862 15688 6138 15730
rect 6262 15770 6538 15812
rect 6262 15730 6380 15770
rect 6420 15730 6538 15770
rect 6262 15688 6538 15730
rect 6662 15770 6938 15812
rect 6662 15730 6780 15770
rect 6820 15730 6938 15770
rect 6662 15688 6938 15730
rect 7062 15770 7338 15812
rect 7062 15730 7180 15770
rect 7220 15730 7338 15770
rect 7062 15688 7338 15730
rect 7462 15770 7738 15812
rect 7462 15730 7580 15770
rect 7620 15730 7738 15770
rect 7462 15688 7738 15730
rect 7862 15770 8138 15812
rect 7862 15730 7980 15770
rect 8020 15730 8138 15770
rect 7862 15688 8138 15730
rect 8262 15770 8538 15812
rect 8262 15730 8380 15770
rect 8420 15730 8538 15770
rect 8262 15688 8538 15730
rect 8662 15770 8938 15812
rect 8662 15730 8780 15770
rect 8820 15730 8938 15770
rect 8662 15688 8938 15730
rect 9062 15770 9338 15812
rect 9062 15730 9180 15770
rect 9220 15730 9338 15770
rect 9062 15688 9338 15730
rect 9462 15770 9738 15812
rect 9462 15730 9580 15770
rect 9620 15730 9738 15770
rect 9462 15688 9738 15730
rect 9862 15770 10138 15812
rect 9862 15730 9980 15770
rect 10020 15730 10138 15770
rect 9862 15688 10138 15730
rect 10262 15770 10538 15812
rect 10262 15730 10380 15770
rect 10420 15730 10538 15770
rect 10262 15688 10538 15730
rect 10662 15770 10938 15812
rect 10662 15730 10780 15770
rect 10820 15730 10938 15770
rect 10662 15688 10938 15730
rect 11062 15770 11338 15812
rect 11062 15730 11180 15770
rect 11220 15730 11338 15770
rect 11062 15688 11338 15730
rect 11462 15770 11738 15812
rect 11462 15730 11580 15770
rect 11620 15730 11738 15770
rect 11462 15688 11738 15730
rect 11862 15770 12138 15812
rect 11862 15730 11980 15770
rect 12020 15730 12138 15770
rect 11862 15688 12138 15730
rect 12262 15770 12538 15812
rect 12262 15730 12380 15770
rect 12420 15730 12538 15770
rect 12262 15688 12538 15730
rect 12662 15770 12938 15812
rect 12662 15730 12780 15770
rect 12820 15730 12938 15770
rect 12662 15688 12938 15730
rect 13062 15770 13338 15812
rect 13062 15730 13180 15770
rect 13220 15730 13338 15770
rect 13062 15688 13338 15730
rect 13462 15770 13738 15812
rect 13462 15730 13580 15770
rect 13620 15730 13738 15770
rect 13462 15688 13738 15730
rect 13862 15770 14138 15812
rect 13862 15730 13980 15770
rect 14020 15730 14138 15770
rect 13862 15688 14138 15730
rect 14262 15770 14538 15812
rect 14262 15730 14380 15770
rect 14420 15730 14538 15770
rect 14262 15688 14538 15730
rect 14662 15770 14938 15812
rect 14662 15730 14780 15770
rect 14820 15730 14938 15770
rect 14662 15688 14938 15730
rect 15062 15770 15338 15812
rect 15062 15730 15180 15770
rect 15220 15730 15338 15770
rect 15062 15688 15338 15730
rect 15462 15770 16000 15812
rect 15462 15730 15580 15770
rect 15620 15730 16000 15770
rect 15462 15688 16000 15730
rect 0 15412 16000 15688
rect 0 15370 538 15412
rect 0 15330 380 15370
rect 420 15330 538 15370
rect 0 15288 538 15330
rect 662 15370 938 15412
rect 662 15330 780 15370
rect 820 15330 938 15370
rect 662 15288 938 15330
rect 1062 15370 1338 15412
rect 1062 15330 1180 15370
rect 1220 15330 1338 15370
rect 1062 15288 1338 15330
rect 1462 15370 1738 15412
rect 1462 15330 1580 15370
rect 1620 15330 1738 15370
rect 1462 15288 1738 15330
rect 1862 15370 2138 15412
rect 1862 15330 1980 15370
rect 2020 15330 2138 15370
rect 1862 15288 2138 15330
rect 2262 15370 2538 15412
rect 2262 15330 2380 15370
rect 2420 15330 2538 15370
rect 2262 15288 2538 15330
rect 2662 15370 2938 15412
rect 2662 15330 2780 15370
rect 2820 15330 2938 15370
rect 2662 15288 2938 15330
rect 3062 15370 3338 15412
rect 3062 15330 3180 15370
rect 3220 15330 3338 15370
rect 3062 15288 3338 15330
rect 3462 15370 3738 15412
rect 3462 15330 3580 15370
rect 3620 15330 3738 15370
rect 3462 15288 3738 15330
rect 3862 15370 4138 15412
rect 3862 15330 3980 15370
rect 4020 15330 4138 15370
rect 3862 15288 4138 15330
rect 4262 15370 4538 15412
rect 4262 15330 4380 15370
rect 4420 15330 4538 15370
rect 4262 15288 4538 15330
rect 4662 15370 4938 15412
rect 4662 15330 4780 15370
rect 4820 15330 4938 15370
rect 4662 15288 4938 15330
rect 5062 15370 5338 15412
rect 5062 15330 5180 15370
rect 5220 15330 5338 15370
rect 5062 15288 5338 15330
rect 5462 15370 5738 15412
rect 5462 15330 5580 15370
rect 5620 15330 5738 15370
rect 5462 15288 5738 15330
rect 5862 15370 6138 15412
rect 5862 15330 5980 15370
rect 6020 15330 6138 15370
rect 5862 15288 6138 15330
rect 6262 15370 6538 15412
rect 6262 15330 6380 15370
rect 6420 15330 6538 15370
rect 6262 15288 6538 15330
rect 6662 15370 6938 15412
rect 6662 15330 6780 15370
rect 6820 15330 6938 15370
rect 6662 15288 6938 15330
rect 7062 15370 7338 15412
rect 7062 15330 7180 15370
rect 7220 15330 7338 15370
rect 7062 15288 7338 15330
rect 7462 15370 7738 15412
rect 7462 15330 7580 15370
rect 7620 15330 7738 15370
rect 7462 15288 7738 15330
rect 7862 15370 8138 15412
rect 7862 15330 7980 15370
rect 8020 15330 8138 15370
rect 7862 15288 8138 15330
rect 8262 15370 8538 15412
rect 8262 15330 8380 15370
rect 8420 15330 8538 15370
rect 8262 15288 8538 15330
rect 8662 15370 8938 15412
rect 8662 15330 8780 15370
rect 8820 15330 8938 15370
rect 8662 15288 8938 15330
rect 9062 15370 9338 15412
rect 9062 15330 9180 15370
rect 9220 15330 9338 15370
rect 9062 15288 9338 15330
rect 9462 15370 9738 15412
rect 9462 15330 9580 15370
rect 9620 15330 9738 15370
rect 9462 15288 9738 15330
rect 9862 15370 10138 15412
rect 9862 15330 9980 15370
rect 10020 15330 10138 15370
rect 9862 15288 10138 15330
rect 10262 15370 10538 15412
rect 10262 15330 10380 15370
rect 10420 15330 10538 15370
rect 10262 15288 10538 15330
rect 10662 15370 10938 15412
rect 10662 15330 10780 15370
rect 10820 15330 10938 15370
rect 10662 15288 10938 15330
rect 11062 15370 11338 15412
rect 11062 15330 11180 15370
rect 11220 15330 11338 15370
rect 11062 15288 11338 15330
rect 11462 15370 11738 15412
rect 11462 15330 11580 15370
rect 11620 15330 11738 15370
rect 11462 15288 11738 15330
rect 11862 15370 12138 15412
rect 11862 15330 11980 15370
rect 12020 15330 12138 15370
rect 11862 15288 12138 15330
rect 12262 15370 12538 15412
rect 12262 15330 12380 15370
rect 12420 15330 12538 15370
rect 12262 15288 12538 15330
rect 12662 15370 12938 15412
rect 12662 15330 12780 15370
rect 12820 15330 12938 15370
rect 12662 15288 12938 15330
rect 13062 15370 13338 15412
rect 13062 15330 13180 15370
rect 13220 15330 13338 15370
rect 13062 15288 13338 15330
rect 13462 15370 13738 15412
rect 13462 15330 13580 15370
rect 13620 15330 13738 15370
rect 13462 15288 13738 15330
rect 13862 15370 14138 15412
rect 13862 15330 13980 15370
rect 14020 15330 14138 15370
rect 13862 15288 14138 15330
rect 14262 15370 14538 15412
rect 14262 15330 14380 15370
rect 14420 15330 14538 15370
rect 14262 15288 14538 15330
rect 14662 15370 14938 15412
rect 14662 15330 14780 15370
rect 14820 15330 14938 15370
rect 14662 15288 14938 15330
rect 15062 15370 15338 15412
rect 15062 15330 15180 15370
rect 15220 15330 15338 15370
rect 15062 15288 15338 15330
rect 15462 15370 16000 15412
rect 15462 15330 15580 15370
rect 15620 15330 16000 15370
rect 15462 15288 16000 15330
rect 0 15012 16000 15288
rect 0 14970 538 15012
rect 0 14930 380 14970
rect 420 14930 538 14970
rect 0 14888 538 14930
rect 662 14970 938 15012
rect 662 14930 780 14970
rect 820 14930 938 14970
rect 662 14888 938 14930
rect 1062 14970 1338 15012
rect 1062 14930 1180 14970
rect 1220 14930 1338 14970
rect 1062 14888 1338 14930
rect 1462 14970 1738 15012
rect 1462 14930 1580 14970
rect 1620 14930 1738 14970
rect 1462 14888 1738 14930
rect 1862 14970 2138 15012
rect 1862 14930 1980 14970
rect 2020 14930 2138 14970
rect 1862 14888 2138 14930
rect 2262 14970 2538 15012
rect 2262 14930 2380 14970
rect 2420 14930 2538 14970
rect 2262 14888 2538 14930
rect 2662 14970 2938 15012
rect 2662 14930 2780 14970
rect 2820 14930 2938 14970
rect 2662 14888 2938 14930
rect 3062 14970 3338 15012
rect 3062 14930 3180 14970
rect 3220 14930 3338 14970
rect 3062 14888 3338 14930
rect 3462 14970 3738 15012
rect 3462 14930 3580 14970
rect 3620 14930 3738 14970
rect 3462 14888 3738 14930
rect 3862 14970 4138 15012
rect 3862 14930 3980 14970
rect 4020 14930 4138 14970
rect 3862 14888 4138 14930
rect 4262 14970 4538 15012
rect 4262 14930 4380 14970
rect 4420 14930 4538 14970
rect 4262 14888 4538 14930
rect 4662 14970 4938 15012
rect 4662 14930 4780 14970
rect 4820 14930 4938 14970
rect 4662 14888 4938 14930
rect 5062 14970 5338 15012
rect 5062 14930 5180 14970
rect 5220 14930 5338 14970
rect 5062 14888 5338 14930
rect 5462 14970 5738 15012
rect 5462 14930 5580 14970
rect 5620 14930 5738 14970
rect 5462 14888 5738 14930
rect 5862 14970 6138 15012
rect 5862 14930 5980 14970
rect 6020 14930 6138 14970
rect 5862 14888 6138 14930
rect 6262 14970 6538 15012
rect 6262 14930 6380 14970
rect 6420 14930 6538 14970
rect 6262 14888 6538 14930
rect 6662 14970 6938 15012
rect 6662 14930 6780 14970
rect 6820 14930 6938 14970
rect 6662 14888 6938 14930
rect 7062 14970 7338 15012
rect 7062 14930 7180 14970
rect 7220 14930 7338 14970
rect 7062 14888 7338 14930
rect 7462 14970 7738 15012
rect 7462 14930 7580 14970
rect 7620 14930 7738 14970
rect 7462 14888 7738 14930
rect 7862 14970 8138 15012
rect 7862 14930 7980 14970
rect 8020 14930 8138 14970
rect 7862 14888 8138 14930
rect 8262 14970 8538 15012
rect 8262 14930 8380 14970
rect 8420 14930 8538 14970
rect 8262 14888 8538 14930
rect 8662 14970 8938 15012
rect 8662 14930 8780 14970
rect 8820 14930 8938 14970
rect 8662 14888 8938 14930
rect 9062 14970 9338 15012
rect 9062 14930 9180 14970
rect 9220 14930 9338 14970
rect 9062 14888 9338 14930
rect 9462 14970 9738 15012
rect 9462 14930 9580 14970
rect 9620 14930 9738 14970
rect 9462 14888 9738 14930
rect 9862 14970 10138 15012
rect 9862 14930 9980 14970
rect 10020 14930 10138 14970
rect 9862 14888 10138 14930
rect 10262 14970 10538 15012
rect 10262 14930 10380 14970
rect 10420 14930 10538 14970
rect 10262 14888 10538 14930
rect 10662 14970 10938 15012
rect 10662 14930 10780 14970
rect 10820 14930 10938 14970
rect 10662 14888 10938 14930
rect 11062 14970 11338 15012
rect 11062 14930 11180 14970
rect 11220 14930 11338 14970
rect 11062 14888 11338 14930
rect 11462 14970 11738 15012
rect 11462 14930 11580 14970
rect 11620 14930 11738 14970
rect 11462 14888 11738 14930
rect 11862 14970 12138 15012
rect 11862 14930 11980 14970
rect 12020 14930 12138 14970
rect 11862 14888 12138 14930
rect 12262 14970 12538 15012
rect 12262 14930 12380 14970
rect 12420 14930 12538 14970
rect 12262 14888 12538 14930
rect 12662 14970 12938 15012
rect 12662 14930 12780 14970
rect 12820 14930 12938 14970
rect 12662 14888 12938 14930
rect 13062 14970 13338 15012
rect 13062 14930 13180 14970
rect 13220 14930 13338 14970
rect 13062 14888 13338 14930
rect 13462 14970 13738 15012
rect 13462 14930 13580 14970
rect 13620 14930 13738 14970
rect 13462 14888 13738 14930
rect 13862 14970 14138 15012
rect 13862 14930 13980 14970
rect 14020 14930 14138 14970
rect 13862 14888 14138 14930
rect 14262 14970 14538 15012
rect 14262 14930 14380 14970
rect 14420 14930 14538 14970
rect 14262 14888 14538 14930
rect 14662 14970 14938 15012
rect 14662 14930 14780 14970
rect 14820 14930 14938 14970
rect 14662 14888 14938 14930
rect 15062 14970 15338 15012
rect 15062 14930 15180 14970
rect 15220 14930 15338 14970
rect 15062 14888 15338 14930
rect 15462 14970 16000 15012
rect 15462 14930 15580 14970
rect 15620 14930 16000 14970
rect 15462 14888 16000 14930
rect 0 14612 16000 14888
rect 0 14570 538 14612
rect 0 14530 380 14570
rect 420 14530 538 14570
rect 0 14488 538 14530
rect 662 14570 938 14612
rect 662 14530 780 14570
rect 820 14530 938 14570
rect 662 14488 938 14530
rect 1062 14570 1338 14612
rect 1062 14530 1180 14570
rect 1220 14530 1338 14570
rect 1062 14488 1338 14530
rect 1462 14570 1738 14612
rect 1462 14530 1580 14570
rect 1620 14530 1738 14570
rect 1462 14488 1738 14530
rect 1862 14570 2138 14612
rect 1862 14530 1980 14570
rect 2020 14530 2138 14570
rect 1862 14488 2138 14530
rect 2262 14570 2538 14612
rect 2262 14530 2380 14570
rect 2420 14530 2538 14570
rect 2262 14488 2538 14530
rect 2662 14570 2938 14612
rect 2662 14530 2780 14570
rect 2820 14530 2938 14570
rect 2662 14488 2938 14530
rect 3062 14570 3338 14612
rect 3062 14530 3180 14570
rect 3220 14530 3338 14570
rect 3062 14488 3338 14530
rect 3462 14570 3738 14612
rect 3462 14530 3580 14570
rect 3620 14530 3738 14570
rect 3462 14488 3738 14530
rect 3862 14570 4138 14612
rect 3862 14530 3980 14570
rect 4020 14530 4138 14570
rect 3862 14488 4138 14530
rect 4262 14570 4538 14612
rect 4262 14530 4380 14570
rect 4420 14530 4538 14570
rect 4262 14488 4538 14530
rect 4662 14570 4938 14612
rect 4662 14530 4780 14570
rect 4820 14530 4938 14570
rect 4662 14488 4938 14530
rect 5062 14570 5338 14612
rect 5062 14530 5180 14570
rect 5220 14530 5338 14570
rect 5062 14488 5338 14530
rect 5462 14570 5738 14612
rect 5462 14530 5580 14570
rect 5620 14530 5738 14570
rect 5462 14488 5738 14530
rect 5862 14570 6138 14612
rect 5862 14530 5980 14570
rect 6020 14530 6138 14570
rect 5862 14488 6138 14530
rect 6262 14570 6538 14612
rect 6262 14530 6380 14570
rect 6420 14530 6538 14570
rect 6262 14488 6538 14530
rect 6662 14570 6938 14612
rect 6662 14530 6780 14570
rect 6820 14530 6938 14570
rect 6662 14488 6938 14530
rect 7062 14570 7338 14612
rect 7062 14530 7180 14570
rect 7220 14530 7338 14570
rect 7062 14488 7338 14530
rect 7462 14570 7738 14612
rect 7462 14530 7580 14570
rect 7620 14530 7738 14570
rect 7462 14488 7738 14530
rect 7862 14570 8138 14612
rect 7862 14530 7980 14570
rect 8020 14530 8138 14570
rect 7862 14488 8138 14530
rect 8262 14570 8538 14612
rect 8262 14530 8380 14570
rect 8420 14530 8538 14570
rect 8262 14488 8538 14530
rect 8662 14570 8938 14612
rect 8662 14530 8780 14570
rect 8820 14530 8938 14570
rect 8662 14488 8938 14530
rect 9062 14570 9338 14612
rect 9062 14530 9180 14570
rect 9220 14530 9338 14570
rect 9062 14488 9338 14530
rect 9462 14570 9738 14612
rect 9462 14530 9580 14570
rect 9620 14530 9738 14570
rect 9462 14488 9738 14530
rect 9862 14570 10138 14612
rect 9862 14530 9980 14570
rect 10020 14530 10138 14570
rect 9862 14488 10138 14530
rect 10262 14570 10538 14612
rect 10262 14530 10380 14570
rect 10420 14530 10538 14570
rect 10262 14488 10538 14530
rect 10662 14570 10938 14612
rect 10662 14530 10780 14570
rect 10820 14530 10938 14570
rect 10662 14488 10938 14530
rect 11062 14570 11338 14612
rect 11062 14530 11180 14570
rect 11220 14530 11338 14570
rect 11062 14488 11338 14530
rect 11462 14570 11738 14612
rect 11462 14530 11580 14570
rect 11620 14530 11738 14570
rect 11462 14488 11738 14530
rect 11862 14570 12138 14612
rect 11862 14530 11980 14570
rect 12020 14530 12138 14570
rect 11862 14488 12138 14530
rect 12262 14570 12538 14612
rect 12262 14530 12380 14570
rect 12420 14530 12538 14570
rect 12262 14488 12538 14530
rect 12662 14570 12938 14612
rect 12662 14530 12780 14570
rect 12820 14530 12938 14570
rect 12662 14488 12938 14530
rect 13062 14570 13338 14612
rect 13062 14530 13180 14570
rect 13220 14530 13338 14570
rect 13062 14488 13338 14530
rect 13462 14570 13738 14612
rect 13462 14530 13580 14570
rect 13620 14530 13738 14570
rect 13462 14488 13738 14530
rect 13862 14570 14138 14612
rect 13862 14530 13980 14570
rect 14020 14530 14138 14570
rect 13862 14488 14138 14530
rect 14262 14570 14538 14612
rect 14262 14530 14380 14570
rect 14420 14530 14538 14570
rect 14262 14488 14538 14530
rect 14662 14570 14938 14612
rect 14662 14530 14780 14570
rect 14820 14530 14938 14570
rect 14662 14488 14938 14530
rect 15062 14570 15338 14612
rect 15062 14530 15180 14570
rect 15220 14530 15338 14570
rect 15062 14488 15338 14530
rect 15462 14570 16000 14612
rect 15462 14530 15580 14570
rect 15620 14530 16000 14570
rect 15462 14488 16000 14530
rect 0 14212 16000 14488
rect 0 14170 538 14212
rect 0 14130 380 14170
rect 420 14130 538 14170
rect 0 14088 538 14130
rect 662 14170 938 14212
rect 662 14130 780 14170
rect 820 14130 938 14170
rect 662 14088 938 14130
rect 1062 14170 1338 14212
rect 1062 14130 1180 14170
rect 1220 14130 1338 14170
rect 1062 14088 1338 14130
rect 1462 14170 1738 14212
rect 1462 14130 1580 14170
rect 1620 14130 1738 14170
rect 1462 14088 1738 14130
rect 1862 14170 2138 14212
rect 1862 14130 1980 14170
rect 2020 14130 2138 14170
rect 1862 14088 2138 14130
rect 2262 14170 2538 14212
rect 2262 14130 2380 14170
rect 2420 14130 2538 14170
rect 2262 14088 2538 14130
rect 2662 14170 2938 14212
rect 2662 14130 2780 14170
rect 2820 14130 2938 14170
rect 2662 14088 2938 14130
rect 3062 14170 3338 14212
rect 3062 14130 3180 14170
rect 3220 14130 3338 14170
rect 3062 14088 3338 14130
rect 3462 14170 3738 14212
rect 3462 14130 3580 14170
rect 3620 14130 3738 14170
rect 3462 14088 3738 14130
rect 3862 14170 4138 14212
rect 3862 14130 3980 14170
rect 4020 14130 4138 14170
rect 3862 14088 4138 14130
rect 4262 14170 4538 14212
rect 4262 14130 4380 14170
rect 4420 14130 4538 14170
rect 4262 14088 4538 14130
rect 4662 14170 4938 14212
rect 4662 14130 4780 14170
rect 4820 14130 4938 14170
rect 4662 14088 4938 14130
rect 5062 14170 5338 14212
rect 5062 14130 5180 14170
rect 5220 14130 5338 14170
rect 5062 14088 5338 14130
rect 5462 14170 5738 14212
rect 5462 14130 5580 14170
rect 5620 14130 5738 14170
rect 5462 14088 5738 14130
rect 5862 14170 6138 14212
rect 5862 14130 5980 14170
rect 6020 14130 6138 14170
rect 5862 14088 6138 14130
rect 6262 14170 6538 14212
rect 6262 14130 6380 14170
rect 6420 14130 6538 14170
rect 6262 14088 6538 14130
rect 6662 14170 6938 14212
rect 6662 14130 6780 14170
rect 6820 14130 6938 14170
rect 6662 14088 6938 14130
rect 7062 14170 7338 14212
rect 7062 14130 7180 14170
rect 7220 14130 7338 14170
rect 7062 14088 7338 14130
rect 7462 14170 7738 14212
rect 7462 14130 7580 14170
rect 7620 14130 7738 14170
rect 7462 14088 7738 14130
rect 7862 14170 8138 14212
rect 7862 14130 7980 14170
rect 8020 14130 8138 14170
rect 7862 14088 8138 14130
rect 8262 14170 8538 14212
rect 8262 14130 8380 14170
rect 8420 14130 8538 14170
rect 8262 14088 8538 14130
rect 8662 14170 8938 14212
rect 8662 14130 8780 14170
rect 8820 14130 8938 14170
rect 8662 14088 8938 14130
rect 9062 14170 9338 14212
rect 9062 14130 9180 14170
rect 9220 14130 9338 14170
rect 9062 14088 9338 14130
rect 9462 14170 9738 14212
rect 9462 14130 9580 14170
rect 9620 14130 9738 14170
rect 9462 14088 9738 14130
rect 9862 14170 10138 14212
rect 9862 14130 9980 14170
rect 10020 14130 10138 14170
rect 9862 14088 10138 14130
rect 10262 14170 10538 14212
rect 10262 14130 10380 14170
rect 10420 14130 10538 14170
rect 10262 14088 10538 14130
rect 10662 14170 10938 14212
rect 10662 14130 10780 14170
rect 10820 14130 10938 14170
rect 10662 14088 10938 14130
rect 11062 14170 11338 14212
rect 11062 14130 11180 14170
rect 11220 14130 11338 14170
rect 11062 14088 11338 14130
rect 11462 14170 11738 14212
rect 11462 14130 11580 14170
rect 11620 14130 11738 14170
rect 11462 14088 11738 14130
rect 11862 14170 12138 14212
rect 11862 14130 11980 14170
rect 12020 14130 12138 14170
rect 11862 14088 12138 14130
rect 12262 14170 12538 14212
rect 12262 14130 12380 14170
rect 12420 14130 12538 14170
rect 12262 14088 12538 14130
rect 12662 14170 12938 14212
rect 12662 14130 12780 14170
rect 12820 14130 12938 14170
rect 12662 14088 12938 14130
rect 13062 14170 13338 14212
rect 13062 14130 13180 14170
rect 13220 14130 13338 14170
rect 13062 14088 13338 14130
rect 13462 14170 13738 14212
rect 13462 14130 13580 14170
rect 13620 14130 13738 14170
rect 13462 14088 13738 14130
rect 13862 14170 14138 14212
rect 13862 14130 13980 14170
rect 14020 14130 14138 14170
rect 13862 14088 14138 14130
rect 14262 14170 14538 14212
rect 14262 14130 14380 14170
rect 14420 14130 14538 14170
rect 14262 14088 14538 14130
rect 14662 14170 14938 14212
rect 14662 14130 14780 14170
rect 14820 14130 14938 14170
rect 14662 14088 14938 14130
rect 15062 14170 15338 14212
rect 15062 14130 15180 14170
rect 15220 14130 15338 14170
rect 15062 14088 15338 14130
rect 15462 14170 16000 14212
rect 15462 14130 15580 14170
rect 15620 14130 16000 14170
rect 15462 14088 16000 14130
rect 0 13812 16000 14088
rect 0 13770 538 13812
rect 0 13730 380 13770
rect 420 13730 538 13770
rect 0 13688 538 13730
rect 662 13770 938 13812
rect 662 13730 780 13770
rect 820 13730 938 13770
rect 662 13688 938 13730
rect 1062 13770 1338 13812
rect 1062 13730 1180 13770
rect 1220 13730 1338 13770
rect 1062 13688 1338 13730
rect 1462 13770 1738 13812
rect 1462 13730 1580 13770
rect 1620 13730 1738 13770
rect 1462 13688 1738 13730
rect 1862 13770 2138 13812
rect 1862 13730 1980 13770
rect 2020 13730 2138 13770
rect 1862 13688 2138 13730
rect 2262 13770 2538 13812
rect 2262 13730 2380 13770
rect 2420 13730 2538 13770
rect 2262 13688 2538 13730
rect 2662 13770 2938 13812
rect 2662 13730 2780 13770
rect 2820 13730 2938 13770
rect 2662 13688 2938 13730
rect 3062 13770 3338 13812
rect 3062 13730 3180 13770
rect 3220 13730 3338 13770
rect 3062 13688 3338 13730
rect 3462 13770 3738 13812
rect 3462 13730 3580 13770
rect 3620 13730 3738 13770
rect 3462 13688 3738 13730
rect 3862 13770 4138 13812
rect 3862 13730 3980 13770
rect 4020 13730 4138 13770
rect 3862 13688 4138 13730
rect 4262 13770 4538 13812
rect 4262 13730 4380 13770
rect 4420 13730 4538 13770
rect 4262 13688 4538 13730
rect 4662 13770 4938 13812
rect 4662 13730 4780 13770
rect 4820 13730 4938 13770
rect 4662 13688 4938 13730
rect 5062 13770 5338 13812
rect 5062 13730 5180 13770
rect 5220 13730 5338 13770
rect 5062 13688 5338 13730
rect 5462 13770 5738 13812
rect 5462 13730 5580 13770
rect 5620 13730 5738 13770
rect 5462 13688 5738 13730
rect 5862 13770 6138 13812
rect 5862 13730 5980 13770
rect 6020 13730 6138 13770
rect 5862 13688 6138 13730
rect 6262 13770 6538 13812
rect 6262 13730 6380 13770
rect 6420 13730 6538 13770
rect 6262 13688 6538 13730
rect 6662 13770 6938 13812
rect 6662 13730 6780 13770
rect 6820 13730 6938 13770
rect 6662 13688 6938 13730
rect 7062 13770 7338 13812
rect 7062 13730 7180 13770
rect 7220 13730 7338 13770
rect 7062 13688 7338 13730
rect 7462 13770 7738 13812
rect 7462 13730 7580 13770
rect 7620 13730 7738 13770
rect 7462 13688 7738 13730
rect 7862 13770 8138 13812
rect 7862 13730 7980 13770
rect 8020 13730 8138 13770
rect 7862 13688 8138 13730
rect 8262 13770 8538 13812
rect 8262 13730 8380 13770
rect 8420 13730 8538 13770
rect 8262 13688 8538 13730
rect 8662 13770 8938 13812
rect 8662 13730 8780 13770
rect 8820 13730 8938 13770
rect 8662 13688 8938 13730
rect 9062 13770 9338 13812
rect 9062 13730 9180 13770
rect 9220 13730 9338 13770
rect 9062 13688 9338 13730
rect 9462 13770 9738 13812
rect 9462 13730 9580 13770
rect 9620 13730 9738 13770
rect 9462 13688 9738 13730
rect 9862 13770 10138 13812
rect 9862 13730 9980 13770
rect 10020 13730 10138 13770
rect 9862 13688 10138 13730
rect 10262 13770 10538 13812
rect 10262 13730 10380 13770
rect 10420 13730 10538 13770
rect 10262 13688 10538 13730
rect 10662 13770 10938 13812
rect 10662 13730 10780 13770
rect 10820 13730 10938 13770
rect 10662 13688 10938 13730
rect 11062 13770 11338 13812
rect 11062 13730 11180 13770
rect 11220 13730 11338 13770
rect 11062 13688 11338 13730
rect 11462 13770 11738 13812
rect 11462 13730 11580 13770
rect 11620 13730 11738 13770
rect 11462 13688 11738 13730
rect 11862 13770 12138 13812
rect 11862 13730 11980 13770
rect 12020 13730 12138 13770
rect 11862 13688 12138 13730
rect 12262 13770 12538 13812
rect 12262 13730 12380 13770
rect 12420 13730 12538 13770
rect 12262 13688 12538 13730
rect 12662 13770 12938 13812
rect 12662 13730 12780 13770
rect 12820 13730 12938 13770
rect 12662 13688 12938 13730
rect 13062 13770 13338 13812
rect 13062 13730 13180 13770
rect 13220 13730 13338 13770
rect 13062 13688 13338 13730
rect 13462 13770 13738 13812
rect 13462 13730 13580 13770
rect 13620 13730 13738 13770
rect 13462 13688 13738 13730
rect 13862 13770 14138 13812
rect 13862 13730 13980 13770
rect 14020 13730 14138 13770
rect 13862 13688 14138 13730
rect 14262 13770 14538 13812
rect 14262 13730 14380 13770
rect 14420 13730 14538 13770
rect 14262 13688 14538 13730
rect 14662 13770 14938 13812
rect 14662 13730 14780 13770
rect 14820 13730 14938 13770
rect 14662 13688 14938 13730
rect 15062 13770 15338 13812
rect 15062 13730 15180 13770
rect 15220 13730 15338 13770
rect 15062 13688 15338 13730
rect 15462 13770 16000 13812
rect 15462 13730 15580 13770
rect 15620 13730 16000 13770
rect 15462 13688 16000 13730
rect 0 13200 16000 13688
rect 0 11512 16000 12000
rect 0 11470 538 11512
rect 0 11430 380 11470
rect 420 11430 538 11470
rect 0 11388 538 11430
rect 662 11470 938 11512
rect 662 11430 780 11470
rect 820 11430 938 11470
rect 662 11388 938 11430
rect 1062 11470 1338 11512
rect 1062 11430 1180 11470
rect 1220 11430 1338 11470
rect 1062 11388 1338 11430
rect 1462 11470 1738 11512
rect 1462 11430 1580 11470
rect 1620 11430 1738 11470
rect 1462 11388 1738 11430
rect 1862 11470 2138 11512
rect 1862 11430 1980 11470
rect 2020 11430 2138 11470
rect 1862 11388 2138 11430
rect 2262 11470 2538 11512
rect 2262 11430 2380 11470
rect 2420 11430 2538 11470
rect 2262 11388 2538 11430
rect 2662 11470 2938 11512
rect 2662 11430 2780 11470
rect 2820 11430 2938 11470
rect 2662 11388 2938 11430
rect 3062 11470 3338 11512
rect 3062 11430 3180 11470
rect 3220 11430 3338 11470
rect 3062 11388 3338 11430
rect 3462 11470 3738 11512
rect 3462 11430 3580 11470
rect 3620 11430 3738 11470
rect 3462 11388 3738 11430
rect 3862 11470 4138 11512
rect 3862 11430 3980 11470
rect 4020 11430 4138 11470
rect 3862 11388 4138 11430
rect 4262 11470 4538 11512
rect 4262 11430 4380 11470
rect 4420 11430 4538 11470
rect 4262 11388 4538 11430
rect 4662 11470 4938 11512
rect 4662 11430 4780 11470
rect 4820 11430 4938 11470
rect 4662 11388 4938 11430
rect 5062 11470 5338 11512
rect 5062 11430 5180 11470
rect 5220 11430 5338 11470
rect 5062 11388 5338 11430
rect 5462 11470 5738 11512
rect 5462 11430 5580 11470
rect 5620 11430 5738 11470
rect 5462 11388 5738 11430
rect 5862 11470 6138 11512
rect 5862 11430 5980 11470
rect 6020 11430 6138 11470
rect 5862 11388 6138 11430
rect 6262 11470 6538 11512
rect 6262 11430 6380 11470
rect 6420 11430 6538 11470
rect 6262 11388 6538 11430
rect 6662 11470 6938 11512
rect 6662 11430 6780 11470
rect 6820 11430 6938 11470
rect 6662 11388 6938 11430
rect 7062 11470 7338 11512
rect 7062 11430 7180 11470
rect 7220 11430 7338 11470
rect 7062 11388 7338 11430
rect 7462 11470 7738 11512
rect 7462 11430 7580 11470
rect 7620 11430 7738 11470
rect 7462 11388 7738 11430
rect 7862 11470 8138 11512
rect 7862 11430 7980 11470
rect 8020 11430 8138 11470
rect 7862 11388 8138 11430
rect 8262 11470 8538 11512
rect 8262 11430 8380 11470
rect 8420 11430 8538 11470
rect 8262 11388 8538 11430
rect 8662 11470 8938 11512
rect 8662 11430 8780 11470
rect 8820 11430 8938 11470
rect 8662 11388 8938 11430
rect 9062 11470 9338 11512
rect 9062 11430 9180 11470
rect 9220 11430 9338 11470
rect 9062 11388 9338 11430
rect 9462 11470 9738 11512
rect 9462 11430 9580 11470
rect 9620 11430 9738 11470
rect 9462 11388 9738 11430
rect 9862 11470 10138 11512
rect 9862 11430 9980 11470
rect 10020 11430 10138 11470
rect 9862 11388 10138 11430
rect 10262 11470 10538 11512
rect 10262 11430 10380 11470
rect 10420 11430 10538 11470
rect 10262 11388 10538 11430
rect 10662 11470 10938 11512
rect 10662 11430 10780 11470
rect 10820 11430 10938 11470
rect 10662 11388 10938 11430
rect 11062 11470 11338 11512
rect 11062 11430 11180 11470
rect 11220 11430 11338 11470
rect 11062 11388 11338 11430
rect 11462 11470 11738 11512
rect 11462 11430 11580 11470
rect 11620 11430 11738 11470
rect 11462 11388 11738 11430
rect 11862 11470 12138 11512
rect 11862 11430 11980 11470
rect 12020 11430 12138 11470
rect 11862 11388 12138 11430
rect 12262 11470 12538 11512
rect 12262 11430 12380 11470
rect 12420 11430 12538 11470
rect 12262 11388 12538 11430
rect 12662 11470 12938 11512
rect 12662 11430 12780 11470
rect 12820 11430 12938 11470
rect 12662 11388 12938 11430
rect 13062 11470 13338 11512
rect 13062 11430 13180 11470
rect 13220 11430 13338 11470
rect 13062 11388 13338 11430
rect 13462 11470 13738 11512
rect 13462 11430 13580 11470
rect 13620 11430 13738 11470
rect 13462 11388 13738 11430
rect 13862 11470 14138 11512
rect 13862 11430 13980 11470
rect 14020 11430 14138 11470
rect 13862 11388 14138 11430
rect 14262 11470 14538 11512
rect 14262 11430 14380 11470
rect 14420 11430 14538 11470
rect 14262 11388 14538 11430
rect 14662 11470 14938 11512
rect 14662 11430 14780 11470
rect 14820 11430 14938 11470
rect 14662 11388 14938 11430
rect 15062 11470 15338 11512
rect 15062 11430 15180 11470
rect 15220 11430 15338 11470
rect 15062 11388 15338 11430
rect 15462 11470 16000 11512
rect 15462 11430 15580 11470
rect 15620 11430 16000 11470
rect 15462 11388 16000 11430
rect 0 11112 16000 11388
rect 0 11070 538 11112
rect 0 11030 380 11070
rect 420 11030 538 11070
rect 0 10988 538 11030
rect 662 11070 938 11112
rect 662 11030 780 11070
rect 820 11030 938 11070
rect 662 10988 938 11030
rect 1062 11070 1338 11112
rect 1062 11030 1180 11070
rect 1220 11030 1338 11070
rect 1062 10988 1338 11030
rect 1462 11070 1738 11112
rect 1462 11030 1580 11070
rect 1620 11030 1738 11070
rect 1462 10988 1738 11030
rect 1862 11070 2138 11112
rect 1862 11030 1980 11070
rect 2020 11030 2138 11070
rect 1862 10988 2138 11030
rect 2262 11070 2538 11112
rect 2262 11030 2380 11070
rect 2420 11030 2538 11070
rect 2262 10988 2538 11030
rect 2662 11070 2938 11112
rect 2662 11030 2780 11070
rect 2820 11030 2938 11070
rect 2662 10988 2938 11030
rect 3062 11070 3338 11112
rect 3062 11030 3180 11070
rect 3220 11030 3338 11070
rect 3062 10988 3338 11030
rect 3462 11070 3738 11112
rect 3462 11030 3580 11070
rect 3620 11030 3738 11070
rect 3462 10988 3738 11030
rect 3862 11070 4138 11112
rect 3862 11030 3980 11070
rect 4020 11030 4138 11070
rect 3862 10988 4138 11030
rect 4262 11070 4538 11112
rect 4262 11030 4380 11070
rect 4420 11030 4538 11070
rect 4262 10988 4538 11030
rect 4662 11070 4938 11112
rect 4662 11030 4780 11070
rect 4820 11030 4938 11070
rect 4662 10988 4938 11030
rect 5062 11070 5338 11112
rect 5062 11030 5180 11070
rect 5220 11030 5338 11070
rect 5062 10988 5338 11030
rect 5462 11070 5738 11112
rect 5462 11030 5580 11070
rect 5620 11030 5738 11070
rect 5462 10988 5738 11030
rect 5862 11070 6138 11112
rect 5862 11030 5980 11070
rect 6020 11030 6138 11070
rect 5862 10988 6138 11030
rect 6262 11070 6538 11112
rect 6262 11030 6380 11070
rect 6420 11030 6538 11070
rect 6262 10988 6538 11030
rect 6662 11070 6938 11112
rect 6662 11030 6780 11070
rect 6820 11030 6938 11070
rect 6662 10988 6938 11030
rect 7062 11070 7338 11112
rect 7062 11030 7180 11070
rect 7220 11030 7338 11070
rect 7062 10988 7338 11030
rect 7462 11070 7738 11112
rect 7462 11030 7580 11070
rect 7620 11030 7738 11070
rect 7462 10988 7738 11030
rect 7862 11070 8138 11112
rect 7862 11030 7980 11070
rect 8020 11030 8138 11070
rect 7862 10988 8138 11030
rect 8262 11070 8538 11112
rect 8262 11030 8380 11070
rect 8420 11030 8538 11070
rect 8262 10988 8538 11030
rect 8662 11070 8938 11112
rect 8662 11030 8780 11070
rect 8820 11030 8938 11070
rect 8662 10988 8938 11030
rect 9062 11070 9338 11112
rect 9062 11030 9180 11070
rect 9220 11030 9338 11070
rect 9062 10988 9338 11030
rect 9462 11070 9738 11112
rect 9462 11030 9580 11070
rect 9620 11030 9738 11070
rect 9462 10988 9738 11030
rect 9862 11070 10138 11112
rect 9862 11030 9980 11070
rect 10020 11030 10138 11070
rect 9862 10988 10138 11030
rect 10262 11070 10538 11112
rect 10262 11030 10380 11070
rect 10420 11030 10538 11070
rect 10262 10988 10538 11030
rect 10662 11070 10938 11112
rect 10662 11030 10780 11070
rect 10820 11030 10938 11070
rect 10662 10988 10938 11030
rect 11062 11070 11338 11112
rect 11062 11030 11180 11070
rect 11220 11030 11338 11070
rect 11062 10988 11338 11030
rect 11462 11070 11738 11112
rect 11462 11030 11580 11070
rect 11620 11030 11738 11070
rect 11462 10988 11738 11030
rect 11862 11070 12138 11112
rect 11862 11030 11980 11070
rect 12020 11030 12138 11070
rect 11862 10988 12138 11030
rect 12262 11070 12538 11112
rect 12262 11030 12380 11070
rect 12420 11030 12538 11070
rect 12262 10988 12538 11030
rect 12662 11070 12938 11112
rect 12662 11030 12780 11070
rect 12820 11030 12938 11070
rect 12662 10988 12938 11030
rect 13062 11070 13338 11112
rect 13062 11030 13180 11070
rect 13220 11030 13338 11070
rect 13062 10988 13338 11030
rect 13462 11070 13738 11112
rect 13462 11030 13580 11070
rect 13620 11030 13738 11070
rect 13462 10988 13738 11030
rect 13862 11070 14138 11112
rect 13862 11030 13980 11070
rect 14020 11030 14138 11070
rect 13862 10988 14138 11030
rect 14262 11070 14538 11112
rect 14262 11030 14380 11070
rect 14420 11030 14538 11070
rect 14262 10988 14538 11030
rect 14662 11070 14938 11112
rect 14662 11030 14780 11070
rect 14820 11030 14938 11070
rect 14662 10988 14938 11030
rect 15062 11070 15338 11112
rect 15062 11030 15180 11070
rect 15220 11030 15338 11070
rect 15062 10988 15338 11030
rect 15462 11070 16000 11112
rect 15462 11030 15580 11070
rect 15620 11030 16000 11070
rect 15462 10988 16000 11030
rect 0 10712 16000 10988
rect 0 10670 538 10712
rect 0 10630 380 10670
rect 420 10630 538 10670
rect 0 10588 538 10630
rect 662 10670 938 10712
rect 662 10630 780 10670
rect 820 10630 938 10670
rect 662 10588 938 10630
rect 1062 10670 1338 10712
rect 1062 10630 1180 10670
rect 1220 10630 1338 10670
rect 1062 10588 1338 10630
rect 1462 10670 1738 10712
rect 1462 10630 1580 10670
rect 1620 10630 1738 10670
rect 1462 10588 1738 10630
rect 1862 10670 2138 10712
rect 1862 10630 1980 10670
rect 2020 10630 2138 10670
rect 1862 10588 2138 10630
rect 2262 10670 2538 10712
rect 2262 10630 2380 10670
rect 2420 10630 2538 10670
rect 2262 10588 2538 10630
rect 2662 10670 2938 10712
rect 2662 10630 2780 10670
rect 2820 10630 2938 10670
rect 2662 10588 2938 10630
rect 3062 10670 3338 10712
rect 3062 10630 3180 10670
rect 3220 10630 3338 10670
rect 3062 10588 3338 10630
rect 3462 10670 3738 10712
rect 3462 10630 3580 10670
rect 3620 10630 3738 10670
rect 3462 10588 3738 10630
rect 3862 10670 4138 10712
rect 3862 10630 3980 10670
rect 4020 10630 4138 10670
rect 3862 10588 4138 10630
rect 4262 10670 4538 10712
rect 4262 10630 4380 10670
rect 4420 10630 4538 10670
rect 4262 10588 4538 10630
rect 4662 10670 4938 10712
rect 4662 10630 4780 10670
rect 4820 10630 4938 10670
rect 4662 10588 4938 10630
rect 5062 10670 5338 10712
rect 5062 10630 5180 10670
rect 5220 10630 5338 10670
rect 5062 10588 5338 10630
rect 5462 10670 5738 10712
rect 5462 10630 5580 10670
rect 5620 10630 5738 10670
rect 5462 10588 5738 10630
rect 5862 10670 6138 10712
rect 5862 10630 5980 10670
rect 6020 10630 6138 10670
rect 5862 10588 6138 10630
rect 6262 10670 6538 10712
rect 6262 10630 6380 10670
rect 6420 10630 6538 10670
rect 6262 10588 6538 10630
rect 6662 10670 6938 10712
rect 6662 10630 6780 10670
rect 6820 10630 6938 10670
rect 6662 10588 6938 10630
rect 7062 10670 7338 10712
rect 7062 10630 7180 10670
rect 7220 10630 7338 10670
rect 7062 10588 7338 10630
rect 7462 10670 7738 10712
rect 7462 10630 7580 10670
rect 7620 10630 7738 10670
rect 7462 10588 7738 10630
rect 7862 10670 8138 10712
rect 7862 10630 7980 10670
rect 8020 10630 8138 10670
rect 7862 10588 8138 10630
rect 8262 10670 8538 10712
rect 8262 10630 8380 10670
rect 8420 10630 8538 10670
rect 8262 10588 8538 10630
rect 8662 10670 8938 10712
rect 8662 10630 8780 10670
rect 8820 10630 8938 10670
rect 8662 10588 8938 10630
rect 9062 10670 9338 10712
rect 9062 10630 9180 10670
rect 9220 10630 9338 10670
rect 9062 10588 9338 10630
rect 9462 10670 9738 10712
rect 9462 10630 9580 10670
rect 9620 10630 9738 10670
rect 9462 10588 9738 10630
rect 9862 10670 10138 10712
rect 9862 10630 9980 10670
rect 10020 10630 10138 10670
rect 9862 10588 10138 10630
rect 10262 10670 10538 10712
rect 10262 10630 10380 10670
rect 10420 10630 10538 10670
rect 10262 10588 10538 10630
rect 10662 10670 10938 10712
rect 10662 10630 10780 10670
rect 10820 10630 10938 10670
rect 10662 10588 10938 10630
rect 11062 10670 11338 10712
rect 11062 10630 11180 10670
rect 11220 10630 11338 10670
rect 11062 10588 11338 10630
rect 11462 10670 11738 10712
rect 11462 10630 11580 10670
rect 11620 10630 11738 10670
rect 11462 10588 11738 10630
rect 11862 10670 12138 10712
rect 11862 10630 11980 10670
rect 12020 10630 12138 10670
rect 11862 10588 12138 10630
rect 12262 10670 12538 10712
rect 12262 10630 12380 10670
rect 12420 10630 12538 10670
rect 12262 10588 12538 10630
rect 12662 10670 12938 10712
rect 12662 10630 12780 10670
rect 12820 10630 12938 10670
rect 12662 10588 12938 10630
rect 13062 10670 13338 10712
rect 13062 10630 13180 10670
rect 13220 10630 13338 10670
rect 13062 10588 13338 10630
rect 13462 10670 13738 10712
rect 13462 10630 13580 10670
rect 13620 10630 13738 10670
rect 13462 10588 13738 10630
rect 13862 10670 14138 10712
rect 13862 10630 13980 10670
rect 14020 10630 14138 10670
rect 13862 10588 14138 10630
rect 14262 10670 14538 10712
rect 14262 10630 14380 10670
rect 14420 10630 14538 10670
rect 14262 10588 14538 10630
rect 14662 10670 14938 10712
rect 14662 10630 14780 10670
rect 14820 10630 14938 10670
rect 14662 10588 14938 10630
rect 15062 10670 15338 10712
rect 15062 10630 15180 10670
rect 15220 10630 15338 10670
rect 15062 10588 15338 10630
rect 15462 10670 16000 10712
rect 15462 10630 15580 10670
rect 15620 10630 16000 10670
rect 15462 10588 16000 10630
rect 0 10312 16000 10588
rect 0 10270 538 10312
rect 0 10230 380 10270
rect 420 10230 538 10270
rect 0 10188 538 10230
rect 662 10270 938 10312
rect 662 10230 780 10270
rect 820 10230 938 10270
rect 662 10188 938 10230
rect 1062 10270 1338 10312
rect 1062 10230 1180 10270
rect 1220 10230 1338 10270
rect 1062 10188 1338 10230
rect 1462 10270 1738 10312
rect 1462 10230 1580 10270
rect 1620 10230 1738 10270
rect 1462 10188 1738 10230
rect 1862 10270 2138 10312
rect 1862 10230 1980 10270
rect 2020 10230 2138 10270
rect 1862 10188 2138 10230
rect 2262 10270 2538 10312
rect 2262 10230 2380 10270
rect 2420 10230 2538 10270
rect 2262 10188 2538 10230
rect 2662 10270 2938 10312
rect 2662 10230 2780 10270
rect 2820 10230 2938 10270
rect 2662 10188 2938 10230
rect 3062 10270 3338 10312
rect 3062 10230 3180 10270
rect 3220 10230 3338 10270
rect 3062 10188 3338 10230
rect 3462 10270 3738 10312
rect 3462 10230 3580 10270
rect 3620 10230 3738 10270
rect 3462 10188 3738 10230
rect 3862 10270 4138 10312
rect 3862 10230 3980 10270
rect 4020 10230 4138 10270
rect 3862 10188 4138 10230
rect 4262 10270 4538 10312
rect 4262 10230 4380 10270
rect 4420 10230 4538 10270
rect 4262 10188 4538 10230
rect 4662 10270 4938 10312
rect 4662 10230 4780 10270
rect 4820 10230 4938 10270
rect 4662 10188 4938 10230
rect 5062 10270 5338 10312
rect 5062 10230 5180 10270
rect 5220 10230 5338 10270
rect 5062 10188 5338 10230
rect 5462 10270 5738 10312
rect 5462 10230 5580 10270
rect 5620 10230 5738 10270
rect 5462 10188 5738 10230
rect 5862 10270 6138 10312
rect 5862 10230 5980 10270
rect 6020 10230 6138 10270
rect 5862 10188 6138 10230
rect 6262 10270 6538 10312
rect 6262 10230 6380 10270
rect 6420 10230 6538 10270
rect 6262 10188 6538 10230
rect 6662 10270 6938 10312
rect 6662 10230 6780 10270
rect 6820 10230 6938 10270
rect 6662 10188 6938 10230
rect 7062 10270 7338 10312
rect 7062 10230 7180 10270
rect 7220 10230 7338 10270
rect 7062 10188 7338 10230
rect 7462 10270 7738 10312
rect 7462 10230 7580 10270
rect 7620 10230 7738 10270
rect 7462 10188 7738 10230
rect 7862 10270 8138 10312
rect 7862 10230 7980 10270
rect 8020 10230 8138 10270
rect 7862 10188 8138 10230
rect 8262 10270 8538 10312
rect 8262 10230 8380 10270
rect 8420 10230 8538 10270
rect 8262 10188 8538 10230
rect 8662 10270 8938 10312
rect 8662 10230 8780 10270
rect 8820 10230 8938 10270
rect 8662 10188 8938 10230
rect 9062 10270 9338 10312
rect 9062 10230 9180 10270
rect 9220 10230 9338 10270
rect 9062 10188 9338 10230
rect 9462 10270 9738 10312
rect 9462 10230 9580 10270
rect 9620 10230 9738 10270
rect 9462 10188 9738 10230
rect 9862 10270 10138 10312
rect 9862 10230 9980 10270
rect 10020 10230 10138 10270
rect 9862 10188 10138 10230
rect 10262 10270 10538 10312
rect 10262 10230 10380 10270
rect 10420 10230 10538 10270
rect 10262 10188 10538 10230
rect 10662 10270 10938 10312
rect 10662 10230 10780 10270
rect 10820 10230 10938 10270
rect 10662 10188 10938 10230
rect 11062 10270 11338 10312
rect 11062 10230 11180 10270
rect 11220 10230 11338 10270
rect 11062 10188 11338 10230
rect 11462 10270 11738 10312
rect 11462 10230 11580 10270
rect 11620 10230 11738 10270
rect 11462 10188 11738 10230
rect 11862 10270 12138 10312
rect 11862 10230 11980 10270
rect 12020 10230 12138 10270
rect 11862 10188 12138 10230
rect 12262 10270 12538 10312
rect 12262 10230 12380 10270
rect 12420 10230 12538 10270
rect 12262 10188 12538 10230
rect 12662 10270 12938 10312
rect 12662 10230 12780 10270
rect 12820 10230 12938 10270
rect 12662 10188 12938 10230
rect 13062 10270 13338 10312
rect 13062 10230 13180 10270
rect 13220 10230 13338 10270
rect 13062 10188 13338 10230
rect 13462 10270 13738 10312
rect 13462 10230 13580 10270
rect 13620 10230 13738 10270
rect 13462 10188 13738 10230
rect 13862 10270 14138 10312
rect 13862 10230 13980 10270
rect 14020 10230 14138 10270
rect 13862 10188 14138 10230
rect 14262 10270 14538 10312
rect 14262 10230 14380 10270
rect 14420 10230 14538 10270
rect 14262 10188 14538 10230
rect 14662 10270 14938 10312
rect 14662 10230 14780 10270
rect 14820 10230 14938 10270
rect 14662 10188 14938 10230
rect 15062 10270 15338 10312
rect 15062 10230 15180 10270
rect 15220 10230 15338 10270
rect 15062 10188 15338 10230
rect 15462 10270 16000 10312
rect 15462 10230 15580 10270
rect 15620 10230 16000 10270
rect 15462 10188 16000 10230
rect 0 9912 16000 10188
rect 0 9870 538 9912
rect 0 9830 380 9870
rect 420 9830 538 9870
rect 0 9788 538 9830
rect 662 9870 938 9912
rect 662 9830 780 9870
rect 820 9830 938 9870
rect 662 9788 938 9830
rect 1062 9870 1338 9912
rect 1062 9830 1180 9870
rect 1220 9830 1338 9870
rect 1062 9788 1338 9830
rect 1462 9870 1738 9912
rect 1462 9830 1580 9870
rect 1620 9830 1738 9870
rect 1462 9788 1738 9830
rect 1862 9870 2138 9912
rect 1862 9830 1980 9870
rect 2020 9830 2138 9870
rect 1862 9788 2138 9830
rect 2262 9870 2538 9912
rect 2262 9830 2380 9870
rect 2420 9830 2538 9870
rect 2262 9788 2538 9830
rect 2662 9870 2938 9912
rect 2662 9830 2780 9870
rect 2820 9830 2938 9870
rect 2662 9788 2938 9830
rect 3062 9870 3338 9912
rect 3062 9830 3180 9870
rect 3220 9830 3338 9870
rect 3062 9788 3338 9830
rect 3462 9870 3738 9912
rect 3462 9830 3580 9870
rect 3620 9830 3738 9870
rect 3462 9788 3738 9830
rect 3862 9870 4138 9912
rect 3862 9830 3980 9870
rect 4020 9830 4138 9870
rect 3862 9788 4138 9830
rect 4262 9870 4538 9912
rect 4262 9830 4380 9870
rect 4420 9830 4538 9870
rect 4262 9788 4538 9830
rect 4662 9870 4938 9912
rect 4662 9830 4780 9870
rect 4820 9830 4938 9870
rect 4662 9788 4938 9830
rect 5062 9870 5338 9912
rect 5062 9830 5180 9870
rect 5220 9830 5338 9870
rect 5062 9788 5338 9830
rect 5462 9870 5738 9912
rect 5462 9830 5580 9870
rect 5620 9830 5738 9870
rect 5462 9788 5738 9830
rect 5862 9870 6138 9912
rect 5862 9830 5980 9870
rect 6020 9830 6138 9870
rect 5862 9788 6138 9830
rect 6262 9870 6538 9912
rect 6262 9830 6380 9870
rect 6420 9830 6538 9870
rect 6262 9788 6538 9830
rect 6662 9870 6938 9912
rect 6662 9830 6780 9870
rect 6820 9830 6938 9870
rect 6662 9788 6938 9830
rect 7062 9870 7338 9912
rect 7062 9830 7180 9870
rect 7220 9830 7338 9870
rect 7062 9788 7338 9830
rect 7462 9870 7738 9912
rect 7462 9830 7580 9870
rect 7620 9830 7738 9870
rect 7462 9788 7738 9830
rect 7862 9870 8138 9912
rect 7862 9830 7980 9870
rect 8020 9830 8138 9870
rect 7862 9788 8138 9830
rect 8262 9870 8538 9912
rect 8262 9830 8380 9870
rect 8420 9830 8538 9870
rect 8262 9788 8538 9830
rect 8662 9870 8938 9912
rect 8662 9830 8780 9870
rect 8820 9830 8938 9870
rect 8662 9788 8938 9830
rect 9062 9870 9338 9912
rect 9062 9830 9180 9870
rect 9220 9830 9338 9870
rect 9062 9788 9338 9830
rect 9462 9870 9738 9912
rect 9462 9830 9580 9870
rect 9620 9830 9738 9870
rect 9462 9788 9738 9830
rect 9862 9870 10138 9912
rect 9862 9830 9980 9870
rect 10020 9830 10138 9870
rect 9862 9788 10138 9830
rect 10262 9870 10538 9912
rect 10262 9830 10380 9870
rect 10420 9830 10538 9870
rect 10262 9788 10538 9830
rect 10662 9870 10938 9912
rect 10662 9830 10780 9870
rect 10820 9830 10938 9870
rect 10662 9788 10938 9830
rect 11062 9870 11338 9912
rect 11062 9830 11180 9870
rect 11220 9830 11338 9870
rect 11062 9788 11338 9830
rect 11462 9870 11738 9912
rect 11462 9830 11580 9870
rect 11620 9830 11738 9870
rect 11462 9788 11738 9830
rect 11862 9870 12138 9912
rect 11862 9830 11980 9870
rect 12020 9830 12138 9870
rect 11862 9788 12138 9830
rect 12262 9870 12538 9912
rect 12262 9830 12380 9870
rect 12420 9830 12538 9870
rect 12262 9788 12538 9830
rect 12662 9870 12938 9912
rect 12662 9830 12780 9870
rect 12820 9830 12938 9870
rect 12662 9788 12938 9830
rect 13062 9870 13338 9912
rect 13062 9830 13180 9870
rect 13220 9830 13338 9870
rect 13062 9788 13338 9830
rect 13462 9870 13738 9912
rect 13462 9830 13580 9870
rect 13620 9830 13738 9870
rect 13462 9788 13738 9830
rect 13862 9870 14138 9912
rect 13862 9830 13980 9870
rect 14020 9830 14138 9870
rect 13862 9788 14138 9830
rect 14262 9870 14538 9912
rect 14262 9830 14380 9870
rect 14420 9830 14538 9870
rect 14262 9788 14538 9830
rect 14662 9870 14938 9912
rect 14662 9830 14780 9870
rect 14820 9830 14938 9870
rect 14662 9788 14938 9830
rect 15062 9870 15338 9912
rect 15062 9830 15180 9870
rect 15220 9830 15338 9870
rect 15062 9788 15338 9830
rect 15462 9870 16000 9912
rect 15462 9830 15580 9870
rect 15620 9830 16000 9870
rect 15462 9788 16000 9830
rect 0 9512 16000 9788
rect 0 9470 538 9512
rect 0 9430 380 9470
rect 420 9430 538 9470
rect 0 9388 538 9430
rect 662 9470 938 9512
rect 662 9430 780 9470
rect 820 9430 938 9470
rect 662 9388 938 9430
rect 1062 9470 1338 9512
rect 1062 9430 1180 9470
rect 1220 9430 1338 9470
rect 1062 9388 1338 9430
rect 1462 9470 1738 9512
rect 1462 9430 1580 9470
rect 1620 9430 1738 9470
rect 1462 9388 1738 9430
rect 1862 9470 2138 9512
rect 1862 9430 1980 9470
rect 2020 9430 2138 9470
rect 1862 9388 2138 9430
rect 2262 9470 2538 9512
rect 2262 9430 2380 9470
rect 2420 9430 2538 9470
rect 2262 9388 2538 9430
rect 2662 9470 2938 9512
rect 2662 9430 2780 9470
rect 2820 9430 2938 9470
rect 2662 9388 2938 9430
rect 3062 9470 3338 9512
rect 3062 9430 3180 9470
rect 3220 9430 3338 9470
rect 3062 9388 3338 9430
rect 3462 9470 3738 9512
rect 3462 9430 3580 9470
rect 3620 9430 3738 9470
rect 3462 9388 3738 9430
rect 3862 9470 4138 9512
rect 3862 9430 3980 9470
rect 4020 9430 4138 9470
rect 3862 9388 4138 9430
rect 4262 9470 4538 9512
rect 4262 9430 4380 9470
rect 4420 9430 4538 9470
rect 4262 9388 4538 9430
rect 4662 9470 4938 9512
rect 4662 9430 4780 9470
rect 4820 9430 4938 9470
rect 4662 9388 4938 9430
rect 5062 9470 5338 9512
rect 5062 9430 5180 9470
rect 5220 9430 5338 9470
rect 5062 9388 5338 9430
rect 5462 9470 5738 9512
rect 5462 9430 5580 9470
rect 5620 9430 5738 9470
rect 5462 9388 5738 9430
rect 5862 9470 6138 9512
rect 5862 9430 5980 9470
rect 6020 9430 6138 9470
rect 5862 9388 6138 9430
rect 6262 9470 6538 9512
rect 6262 9430 6380 9470
rect 6420 9430 6538 9470
rect 6262 9388 6538 9430
rect 6662 9470 6938 9512
rect 6662 9430 6780 9470
rect 6820 9430 6938 9470
rect 6662 9388 6938 9430
rect 7062 9470 7338 9512
rect 7062 9430 7180 9470
rect 7220 9430 7338 9470
rect 7062 9388 7338 9430
rect 7462 9470 7738 9512
rect 7462 9430 7580 9470
rect 7620 9430 7738 9470
rect 7462 9388 7738 9430
rect 7862 9470 8138 9512
rect 7862 9430 7980 9470
rect 8020 9430 8138 9470
rect 7862 9388 8138 9430
rect 8262 9470 8538 9512
rect 8262 9430 8380 9470
rect 8420 9430 8538 9470
rect 8262 9388 8538 9430
rect 8662 9470 8938 9512
rect 8662 9430 8780 9470
rect 8820 9430 8938 9470
rect 8662 9388 8938 9430
rect 9062 9470 9338 9512
rect 9062 9430 9180 9470
rect 9220 9430 9338 9470
rect 9062 9388 9338 9430
rect 9462 9470 9738 9512
rect 9462 9430 9580 9470
rect 9620 9430 9738 9470
rect 9462 9388 9738 9430
rect 9862 9470 10138 9512
rect 9862 9430 9980 9470
rect 10020 9430 10138 9470
rect 9862 9388 10138 9430
rect 10262 9470 10538 9512
rect 10262 9430 10380 9470
rect 10420 9430 10538 9470
rect 10262 9388 10538 9430
rect 10662 9470 10938 9512
rect 10662 9430 10780 9470
rect 10820 9430 10938 9470
rect 10662 9388 10938 9430
rect 11062 9470 11338 9512
rect 11062 9430 11180 9470
rect 11220 9430 11338 9470
rect 11062 9388 11338 9430
rect 11462 9470 11738 9512
rect 11462 9430 11580 9470
rect 11620 9430 11738 9470
rect 11462 9388 11738 9430
rect 11862 9470 12138 9512
rect 11862 9430 11980 9470
rect 12020 9430 12138 9470
rect 11862 9388 12138 9430
rect 12262 9470 12538 9512
rect 12262 9430 12380 9470
rect 12420 9430 12538 9470
rect 12262 9388 12538 9430
rect 12662 9470 12938 9512
rect 12662 9430 12780 9470
rect 12820 9430 12938 9470
rect 12662 9388 12938 9430
rect 13062 9470 13338 9512
rect 13062 9430 13180 9470
rect 13220 9430 13338 9470
rect 13062 9388 13338 9430
rect 13462 9470 13738 9512
rect 13462 9430 13580 9470
rect 13620 9430 13738 9470
rect 13462 9388 13738 9430
rect 13862 9470 14138 9512
rect 13862 9430 13980 9470
rect 14020 9430 14138 9470
rect 13862 9388 14138 9430
rect 14262 9470 14538 9512
rect 14262 9430 14380 9470
rect 14420 9430 14538 9470
rect 14262 9388 14538 9430
rect 14662 9470 14938 9512
rect 14662 9430 14780 9470
rect 14820 9430 14938 9470
rect 14662 9388 14938 9430
rect 15062 9470 15338 9512
rect 15062 9430 15180 9470
rect 15220 9430 15338 9470
rect 15062 9388 15338 9430
rect 15462 9470 16000 9512
rect 15462 9430 15580 9470
rect 15620 9430 16000 9470
rect 15462 9388 16000 9430
rect 0 9112 16000 9388
rect 0 9070 538 9112
rect 0 9030 380 9070
rect 420 9030 538 9070
rect 0 8988 538 9030
rect 662 9070 938 9112
rect 662 9030 780 9070
rect 820 9030 938 9070
rect 662 8988 938 9030
rect 1062 9070 1338 9112
rect 1062 9030 1180 9070
rect 1220 9030 1338 9070
rect 1062 8988 1338 9030
rect 1462 9070 1738 9112
rect 1462 9030 1580 9070
rect 1620 9030 1738 9070
rect 1462 8988 1738 9030
rect 1862 9070 2138 9112
rect 1862 9030 1980 9070
rect 2020 9030 2138 9070
rect 1862 8988 2138 9030
rect 2262 9070 2538 9112
rect 2262 9030 2380 9070
rect 2420 9030 2538 9070
rect 2262 8988 2538 9030
rect 2662 9070 2938 9112
rect 2662 9030 2780 9070
rect 2820 9030 2938 9070
rect 2662 8988 2938 9030
rect 3062 9070 3338 9112
rect 3062 9030 3180 9070
rect 3220 9030 3338 9070
rect 3062 8988 3338 9030
rect 3462 9070 3738 9112
rect 3462 9030 3580 9070
rect 3620 9030 3738 9070
rect 3462 8988 3738 9030
rect 3862 9070 4138 9112
rect 3862 9030 3980 9070
rect 4020 9030 4138 9070
rect 3862 8988 4138 9030
rect 4262 9070 4538 9112
rect 4262 9030 4380 9070
rect 4420 9030 4538 9070
rect 4262 8988 4538 9030
rect 4662 9070 4938 9112
rect 4662 9030 4780 9070
rect 4820 9030 4938 9070
rect 4662 8988 4938 9030
rect 5062 9070 5338 9112
rect 5062 9030 5180 9070
rect 5220 9030 5338 9070
rect 5062 8988 5338 9030
rect 5462 9070 5738 9112
rect 5462 9030 5580 9070
rect 5620 9030 5738 9070
rect 5462 8988 5738 9030
rect 5862 9070 6138 9112
rect 5862 9030 5980 9070
rect 6020 9030 6138 9070
rect 5862 8988 6138 9030
rect 6262 9070 6538 9112
rect 6262 9030 6380 9070
rect 6420 9030 6538 9070
rect 6262 8988 6538 9030
rect 6662 9070 6938 9112
rect 6662 9030 6780 9070
rect 6820 9030 6938 9070
rect 6662 8988 6938 9030
rect 7062 9070 7338 9112
rect 7062 9030 7180 9070
rect 7220 9030 7338 9070
rect 7062 8988 7338 9030
rect 7462 9070 7738 9112
rect 7462 9030 7580 9070
rect 7620 9030 7738 9070
rect 7462 8988 7738 9030
rect 7862 9070 8138 9112
rect 7862 9030 7980 9070
rect 8020 9030 8138 9070
rect 7862 8988 8138 9030
rect 8262 9070 8538 9112
rect 8262 9030 8380 9070
rect 8420 9030 8538 9070
rect 8262 8988 8538 9030
rect 8662 9070 8938 9112
rect 8662 9030 8780 9070
rect 8820 9030 8938 9070
rect 8662 8988 8938 9030
rect 9062 9070 9338 9112
rect 9062 9030 9180 9070
rect 9220 9030 9338 9070
rect 9062 8988 9338 9030
rect 9462 9070 9738 9112
rect 9462 9030 9580 9070
rect 9620 9030 9738 9070
rect 9462 8988 9738 9030
rect 9862 9070 10138 9112
rect 9862 9030 9980 9070
rect 10020 9030 10138 9070
rect 9862 8988 10138 9030
rect 10262 9070 10538 9112
rect 10262 9030 10380 9070
rect 10420 9030 10538 9070
rect 10262 8988 10538 9030
rect 10662 9070 10938 9112
rect 10662 9030 10780 9070
rect 10820 9030 10938 9070
rect 10662 8988 10938 9030
rect 11062 9070 11338 9112
rect 11062 9030 11180 9070
rect 11220 9030 11338 9070
rect 11062 8988 11338 9030
rect 11462 9070 11738 9112
rect 11462 9030 11580 9070
rect 11620 9030 11738 9070
rect 11462 8988 11738 9030
rect 11862 9070 12138 9112
rect 11862 9030 11980 9070
rect 12020 9030 12138 9070
rect 11862 8988 12138 9030
rect 12262 9070 12538 9112
rect 12262 9030 12380 9070
rect 12420 9030 12538 9070
rect 12262 8988 12538 9030
rect 12662 9070 12938 9112
rect 12662 9030 12780 9070
rect 12820 9030 12938 9070
rect 12662 8988 12938 9030
rect 13062 9070 13338 9112
rect 13062 9030 13180 9070
rect 13220 9030 13338 9070
rect 13062 8988 13338 9030
rect 13462 9070 13738 9112
rect 13462 9030 13580 9070
rect 13620 9030 13738 9070
rect 13462 8988 13738 9030
rect 13862 9070 14138 9112
rect 13862 9030 13980 9070
rect 14020 9030 14138 9070
rect 13862 8988 14138 9030
rect 14262 9070 14538 9112
rect 14262 9030 14380 9070
rect 14420 9030 14538 9070
rect 14262 8988 14538 9030
rect 14662 9070 14938 9112
rect 14662 9030 14780 9070
rect 14820 9030 14938 9070
rect 14662 8988 14938 9030
rect 15062 9070 15338 9112
rect 15062 9030 15180 9070
rect 15220 9030 15338 9070
rect 15062 8988 15338 9030
rect 15462 9070 16000 9112
rect 15462 9030 15580 9070
rect 15620 9030 16000 9070
rect 15462 8988 16000 9030
rect 0 8712 16000 8988
rect 0 8670 538 8712
rect 0 8630 380 8670
rect 420 8630 538 8670
rect 0 8588 538 8630
rect 662 8670 938 8712
rect 662 8630 780 8670
rect 820 8630 938 8670
rect 662 8588 938 8630
rect 1062 8670 1338 8712
rect 1062 8630 1180 8670
rect 1220 8630 1338 8670
rect 1062 8588 1338 8630
rect 1462 8670 1738 8712
rect 1462 8630 1580 8670
rect 1620 8630 1738 8670
rect 1462 8588 1738 8630
rect 1862 8670 2138 8712
rect 1862 8630 1980 8670
rect 2020 8630 2138 8670
rect 1862 8588 2138 8630
rect 2262 8670 2538 8712
rect 2262 8630 2380 8670
rect 2420 8630 2538 8670
rect 2262 8588 2538 8630
rect 2662 8670 2938 8712
rect 2662 8630 2780 8670
rect 2820 8630 2938 8670
rect 2662 8588 2938 8630
rect 3062 8670 3338 8712
rect 3062 8630 3180 8670
rect 3220 8630 3338 8670
rect 3062 8588 3338 8630
rect 3462 8670 3738 8712
rect 3462 8630 3580 8670
rect 3620 8630 3738 8670
rect 3462 8588 3738 8630
rect 3862 8670 4138 8712
rect 3862 8630 3980 8670
rect 4020 8630 4138 8670
rect 3862 8588 4138 8630
rect 4262 8670 4538 8712
rect 4262 8630 4380 8670
rect 4420 8630 4538 8670
rect 4262 8588 4538 8630
rect 4662 8670 4938 8712
rect 4662 8630 4780 8670
rect 4820 8630 4938 8670
rect 4662 8588 4938 8630
rect 5062 8670 5338 8712
rect 5062 8630 5180 8670
rect 5220 8630 5338 8670
rect 5062 8588 5338 8630
rect 5462 8670 5738 8712
rect 5462 8630 5580 8670
rect 5620 8630 5738 8670
rect 5462 8588 5738 8630
rect 5862 8670 6138 8712
rect 5862 8630 5980 8670
rect 6020 8630 6138 8670
rect 5862 8588 6138 8630
rect 6262 8670 6538 8712
rect 6262 8630 6380 8670
rect 6420 8630 6538 8670
rect 6262 8588 6538 8630
rect 6662 8670 6938 8712
rect 6662 8630 6780 8670
rect 6820 8630 6938 8670
rect 6662 8588 6938 8630
rect 7062 8670 7338 8712
rect 7062 8630 7180 8670
rect 7220 8630 7338 8670
rect 7062 8588 7338 8630
rect 7462 8670 7738 8712
rect 7462 8630 7580 8670
rect 7620 8630 7738 8670
rect 7462 8588 7738 8630
rect 7862 8670 8138 8712
rect 7862 8630 7980 8670
rect 8020 8630 8138 8670
rect 7862 8588 8138 8630
rect 8262 8670 8538 8712
rect 8262 8630 8380 8670
rect 8420 8630 8538 8670
rect 8262 8588 8538 8630
rect 8662 8670 8938 8712
rect 8662 8630 8780 8670
rect 8820 8630 8938 8670
rect 8662 8588 8938 8630
rect 9062 8670 9338 8712
rect 9062 8630 9180 8670
rect 9220 8630 9338 8670
rect 9062 8588 9338 8630
rect 9462 8670 9738 8712
rect 9462 8630 9580 8670
rect 9620 8630 9738 8670
rect 9462 8588 9738 8630
rect 9862 8670 10138 8712
rect 9862 8630 9980 8670
rect 10020 8630 10138 8670
rect 9862 8588 10138 8630
rect 10262 8670 10538 8712
rect 10262 8630 10380 8670
rect 10420 8630 10538 8670
rect 10262 8588 10538 8630
rect 10662 8670 10938 8712
rect 10662 8630 10780 8670
rect 10820 8630 10938 8670
rect 10662 8588 10938 8630
rect 11062 8670 11338 8712
rect 11062 8630 11180 8670
rect 11220 8630 11338 8670
rect 11062 8588 11338 8630
rect 11462 8670 11738 8712
rect 11462 8630 11580 8670
rect 11620 8630 11738 8670
rect 11462 8588 11738 8630
rect 11862 8670 12138 8712
rect 11862 8630 11980 8670
rect 12020 8630 12138 8670
rect 11862 8588 12138 8630
rect 12262 8670 12538 8712
rect 12262 8630 12380 8670
rect 12420 8630 12538 8670
rect 12262 8588 12538 8630
rect 12662 8670 12938 8712
rect 12662 8630 12780 8670
rect 12820 8630 12938 8670
rect 12662 8588 12938 8630
rect 13062 8670 13338 8712
rect 13062 8630 13180 8670
rect 13220 8630 13338 8670
rect 13062 8588 13338 8630
rect 13462 8670 13738 8712
rect 13462 8630 13580 8670
rect 13620 8630 13738 8670
rect 13462 8588 13738 8630
rect 13862 8670 14138 8712
rect 13862 8630 13980 8670
rect 14020 8630 14138 8670
rect 13862 8588 14138 8630
rect 14262 8670 14538 8712
rect 14262 8630 14380 8670
rect 14420 8630 14538 8670
rect 14262 8588 14538 8630
rect 14662 8670 14938 8712
rect 14662 8630 14780 8670
rect 14820 8630 14938 8670
rect 14662 8588 14938 8630
rect 15062 8670 15338 8712
rect 15062 8630 15180 8670
rect 15220 8630 15338 8670
rect 15062 8588 15338 8630
rect 15462 8670 16000 8712
rect 15462 8630 15580 8670
rect 15620 8630 16000 8670
rect 15462 8588 16000 8630
rect 0 8312 16000 8588
rect 0 8270 538 8312
rect 0 8230 380 8270
rect 420 8230 538 8270
rect 0 8188 538 8230
rect 662 8270 938 8312
rect 662 8230 780 8270
rect 820 8230 938 8270
rect 662 8188 938 8230
rect 1062 8270 1338 8312
rect 1062 8230 1180 8270
rect 1220 8230 1338 8270
rect 1062 8188 1338 8230
rect 1462 8270 1738 8312
rect 1462 8230 1580 8270
rect 1620 8230 1738 8270
rect 1462 8188 1738 8230
rect 1862 8270 2138 8312
rect 1862 8230 1980 8270
rect 2020 8230 2138 8270
rect 1862 8188 2138 8230
rect 2262 8270 2538 8312
rect 2262 8230 2380 8270
rect 2420 8230 2538 8270
rect 2262 8188 2538 8230
rect 2662 8270 2938 8312
rect 2662 8230 2780 8270
rect 2820 8230 2938 8270
rect 2662 8188 2938 8230
rect 3062 8270 3338 8312
rect 3062 8230 3180 8270
rect 3220 8230 3338 8270
rect 3062 8188 3338 8230
rect 3462 8270 3738 8312
rect 3462 8230 3580 8270
rect 3620 8230 3738 8270
rect 3462 8188 3738 8230
rect 3862 8270 4138 8312
rect 3862 8230 3980 8270
rect 4020 8230 4138 8270
rect 3862 8188 4138 8230
rect 4262 8270 4538 8312
rect 4262 8230 4380 8270
rect 4420 8230 4538 8270
rect 4262 8188 4538 8230
rect 4662 8270 4938 8312
rect 4662 8230 4780 8270
rect 4820 8230 4938 8270
rect 4662 8188 4938 8230
rect 5062 8270 5338 8312
rect 5062 8230 5180 8270
rect 5220 8230 5338 8270
rect 5062 8188 5338 8230
rect 5462 8270 5738 8312
rect 5462 8230 5580 8270
rect 5620 8230 5738 8270
rect 5462 8188 5738 8230
rect 5862 8270 6138 8312
rect 5862 8230 5980 8270
rect 6020 8230 6138 8270
rect 5862 8188 6138 8230
rect 6262 8270 6538 8312
rect 6262 8230 6380 8270
rect 6420 8230 6538 8270
rect 6262 8188 6538 8230
rect 6662 8270 6938 8312
rect 6662 8230 6780 8270
rect 6820 8230 6938 8270
rect 6662 8188 6938 8230
rect 7062 8270 7338 8312
rect 7062 8230 7180 8270
rect 7220 8230 7338 8270
rect 7062 8188 7338 8230
rect 7462 8270 7738 8312
rect 7462 8230 7580 8270
rect 7620 8230 7738 8270
rect 7462 8188 7738 8230
rect 7862 8270 8138 8312
rect 7862 8230 7980 8270
rect 8020 8230 8138 8270
rect 7862 8188 8138 8230
rect 8262 8270 8538 8312
rect 8262 8230 8380 8270
rect 8420 8230 8538 8270
rect 8262 8188 8538 8230
rect 8662 8270 8938 8312
rect 8662 8230 8780 8270
rect 8820 8230 8938 8270
rect 8662 8188 8938 8230
rect 9062 8270 9338 8312
rect 9062 8230 9180 8270
rect 9220 8230 9338 8270
rect 9062 8188 9338 8230
rect 9462 8270 9738 8312
rect 9462 8230 9580 8270
rect 9620 8230 9738 8270
rect 9462 8188 9738 8230
rect 9862 8270 10138 8312
rect 9862 8230 9980 8270
rect 10020 8230 10138 8270
rect 9862 8188 10138 8230
rect 10262 8270 10538 8312
rect 10262 8230 10380 8270
rect 10420 8230 10538 8270
rect 10262 8188 10538 8230
rect 10662 8270 10938 8312
rect 10662 8230 10780 8270
rect 10820 8230 10938 8270
rect 10662 8188 10938 8230
rect 11062 8270 11338 8312
rect 11062 8230 11180 8270
rect 11220 8230 11338 8270
rect 11062 8188 11338 8230
rect 11462 8270 11738 8312
rect 11462 8230 11580 8270
rect 11620 8230 11738 8270
rect 11462 8188 11738 8230
rect 11862 8270 12138 8312
rect 11862 8230 11980 8270
rect 12020 8230 12138 8270
rect 11862 8188 12138 8230
rect 12262 8270 12538 8312
rect 12262 8230 12380 8270
rect 12420 8230 12538 8270
rect 12262 8188 12538 8230
rect 12662 8270 12938 8312
rect 12662 8230 12780 8270
rect 12820 8230 12938 8270
rect 12662 8188 12938 8230
rect 13062 8270 13338 8312
rect 13062 8230 13180 8270
rect 13220 8230 13338 8270
rect 13062 8188 13338 8230
rect 13462 8270 13738 8312
rect 13462 8230 13580 8270
rect 13620 8230 13738 8270
rect 13462 8188 13738 8230
rect 13862 8270 14138 8312
rect 13862 8230 13980 8270
rect 14020 8230 14138 8270
rect 13862 8188 14138 8230
rect 14262 8270 14538 8312
rect 14262 8230 14380 8270
rect 14420 8230 14538 8270
rect 14262 8188 14538 8230
rect 14662 8270 14938 8312
rect 14662 8230 14780 8270
rect 14820 8230 14938 8270
rect 14662 8188 14938 8230
rect 15062 8270 15338 8312
rect 15062 8230 15180 8270
rect 15220 8230 15338 8270
rect 15062 8188 15338 8230
rect 15462 8270 16000 8312
rect 15462 8230 15580 8270
rect 15620 8230 16000 8270
rect 15462 8188 16000 8230
rect 0 7912 16000 8188
rect 0 7870 538 7912
rect 0 7830 380 7870
rect 420 7830 538 7870
rect 0 7788 538 7830
rect 662 7870 938 7912
rect 662 7830 780 7870
rect 820 7830 938 7870
rect 662 7788 938 7830
rect 1062 7870 1338 7912
rect 1062 7830 1180 7870
rect 1220 7830 1338 7870
rect 1062 7788 1338 7830
rect 1462 7870 1738 7912
rect 1462 7830 1580 7870
rect 1620 7830 1738 7870
rect 1462 7788 1738 7830
rect 1862 7870 2138 7912
rect 1862 7830 1980 7870
rect 2020 7830 2138 7870
rect 1862 7788 2138 7830
rect 2262 7870 2538 7912
rect 2262 7830 2380 7870
rect 2420 7830 2538 7870
rect 2262 7788 2538 7830
rect 2662 7870 2938 7912
rect 2662 7830 2780 7870
rect 2820 7830 2938 7870
rect 2662 7788 2938 7830
rect 3062 7870 3338 7912
rect 3062 7830 3180 7870
rect 3220 7830 3338 7870
rect 3062 7788 3338 7830
rect 3462 7870 3738 7912
rect 3462 7830 3580 7870
rect 3620 7830 3738 7870
rect 3462 7788 3738 7830
rect 3862 7870 4138 7912
rect 3862 7830 3980 7870
rect 4020 7830 4138 7870
rect 3862 7788 4138 7830
rect 4262 7870 4538 7912
rect 4262 7830 4380 7870
rect 4420 7830 4538 7870
rect 4262 7788 4538 7830
rect 4662 7870 4938 7912
rect 4662 7830 4780 7870
rect 4820 7830 4938 7870
rect 4662 7788 4938 7830
rect 5062 7870 5338 7912
rect 5062 7830 5180 7870
rect 5220 7830 5338 7870
rect 5062 7788 5338 7830
rect 5462 7870 5738 7912
rect 5462 7830 5580 7870
rect 5620 7830 5738 7870
rect 5462 7788 5738 7830
rect 5862 7870 6138 7912
rect 5862 7830 5980 7870
rect 6020 7830 6138 7870
rect 5862 7788 6138 7830
rect 6262 7870 6538 7912
rect 6262 7830 6380 7870
rect 6420 7830 6538 7870
rect 6262 7788 6538 7830
rect 6662 7870 6938 7912
rect 6662 7830 6780 7870
rect 6820 7830 6938 7870
rect 6662 7788 6938 7830
rect 7062 7870 7338 7912
rect 7062 7830 7180 7870
rect 7220 7830 7338 7870
rect 7062 7788 7338 7830
rect 7462 7870 7738 7912
rect 7462 7830 7580 7870
rect 7620 7830 7738 7870
rect 7462 7788 7738 7830
rect 7862 7870 8138 7912
rect 7862 7830 7980 7870
rect 8020 7830 8138 7870
rect 7862 7788 8138 7830
rect 8262 7870 8538 7912
rect 8262 7830 8380 7870
rect 8420 7830 8538 7870
rect 8262 7788 8538 7830
rect 8662 7870 8938 7912
rect 8662 7830 8780 7870
rect 8820 7830 8938 7870
rect 8662 7788 8938 7830
rect 9062 7870 9338 7912
rect 9062 7830 9180 7870
rect 9220 7830 9338 7870
rect 9062 7788 9338 7830
rect 9462 7870 9738 7912
rect 9462 7830 9580 7870
rect 9620 7830 9738 7870
rect 9462 7788 9738 7830
rect 9862 7870 10138 7912
rect 9862 7830 9980 7870
rect 10020 7830 10138 7870
rect 9862 7788 10138 7830
rect 10262 7870 10538 7912
rect 10262 7830 10380 7870
rect 10420 7830 10538 7870
rect 10262 7788 10538 7830
rect 10662 7870 10938 7912
rect 10662 7830 10780 7870
rect 10820 7830 10938 7870
rect 10662 7788 10938 7830
rect 11062 7870 11338 7912
rect 11062 7830 11180 7870
rect 11220 7830 11338 7870
rect 11062 7788 11338 7830
rect 11462 7870 11738 7912
rect 11462 7830 11580 7870
rect 11620 7830 11738 7870
rect 11462 7788 11738 7830
rect 11862 7870 12138 7912
rect 11862 7830 11980 7870
rect 12020 7830 12138 7870
rect 11862 7788 12138 7830
rect 12262 7870 12538 7912
rect 12262 7830 12380 7870
rect 12420 7830 12538 7870
rect 12262 7788 12538 7830
rect 12662 7870 12938 7912
rect 12662 7830 12780 7870
rect 12820 7830 12938 7870
rect 12662 7788 12938 7830
rect 13062 7870 13338 7912
rect 13062 7830 13180 7870
rect 13220 7830 13338 7870
rect 13062 7788 13338 7830
rect 13462 7870 13738 7912
rect 13462 7830 13580 7870
rect 13620 7830 13738 7870
rect 13462 7788 13738 7830
rect 13862 7870 14138 7912
rect 13862 7830 13980 7870
rect 14020 7830 14138 7870
rect 13862 7788 14138 7830
rect 14262 7870 14538 7912
rect 14262 7830 14380 7870
rect 14420 7830 14538 7870
rect 14262 7788 14538 7830
rect 14662 7870 14938 7912
rect 14662 7830 14780 7870
rect 14820 7830 14938 7870
rect 14662 7788 14938 7830
rect 15062 7870 15338 7912
rect 15062 7830 15180 7870
rect 15220 7830 15338 7870
rect 15062 7788 15338 7830
rect 15462 7870 16000 7912
rect 15462 7830 15580 7870
rect 15620 7830 16000 7870
rect 15462 7788 16000 7830
rect 0 7512 16000 7788
rect 0 7470 538 7512
rect 0 7430 380 7470
rect 420 7430 538 7470
rect 0 7388 538 7430
rect 662 7470 938 7512
rect 662 7430 780 7470
rect 820 7430 938 7470
rect 662 7388 938 7430
rect 1062 7470 1338 7512
rect 1062 7430 1180 7470
rect 1220 7430 1338 7470
rect 1062 7388 1338 7430
rect 1462 7470 1738 7512
rect 1462 7430 1580 7470
rect 1620 7430 1738 7470
rect 1462 7388 1738 7430
rect 1862 7470 2138 7512
rect 1862 7430 1980 7470
rect 2020 7430 2138 7470
rect 1862 7388 2138 7430
rect 2262 7470 2538 7512
rect 2262 7430 2380 7470
rect 2420 7430 2538 7470
rect 2262 7388 2538 7430
rect 2662 7470 2938 7512
rect 2662 7430 2780 7470
rect 2820 7430 2938 7470
rect 2662 7388 2938 7430
rect 3062 7470 3338 7512
rect 3062 7430 3180 7470
rect 3220 7430 3338 7470
rect 3062 7388 3338 7430
rect 3462 7470 3738 7512
rect 3462 7430 3580 7470
rect 3620 7430 3738 7470
rect 3462 7388 3738 7430
rect 3862 7470 4138 7512
rect 3862 7430 3980 7470
rect 4020 7430 4138 7470
rect 3862 7388 4138 7430
rect 4262 7470 4538 7512
rect 4262 7430 4380 7470
rect 4420 7430 4538 7470
rect 4262 7388 4538 7430
rect 4662 7470 4938 7512
rect 4662 7430 4780 7470
rect 4820 7430 4938 7470
rect 4662 7388 4938 7430
rect 5062 7470 5338 7512
rect 5062 7430 5180 7470
rect 5220 7430 5338 7470
rect 5062 7388 5338 7430
rect 5462 7470 5738 7512
rect 5462 7430 5580 7470
rect 5620 7430 5738 7470
rect 5462 7388 5738 7430
rect 5862 7470 6138 7512
rect 5862 7430 5980 7470
rect 6020 7430 6138 7470
rect 5862 7388 6138 7430
rect 6262 7470 6538 7512
rect 6262 7430 6380 7470
rect 6420 7430 6538 7470
rect 6262 7388 6538 7430
rect 6662 7470 6938 7512
rect 6662 7430 6780 7470
rect 6820 7430 6938 7470
rect 6662 7388 6938 7430
rect 7062 7470 7338 7512
rect 7062 7430 7180 7470
rect 7220 7430 7338 7470
rect 7062 7388 7338 7430
rect 7462 7470 7738 7512
rect 7462 7430 7580 7470
rect 7620 7430 7738 7470
rect 7462 7388 7738 7430
rect 7862 7470 8138 7512
rect 7862 7430 7980 7470
rect 8020 7430 8138 7470
rect 7862 7388 8138 7430
rect 8262 7470 8538 7512
rect 8262 7430 8380 7470
rect 8420 7430 8538 7470
rect 8262 7388 8538 7430
rect 8662 7470 8938 7512
rect 8662 7430 8780 7470
rect 8820 7430 8938 7470
rect 8662 7388 8938 7430
rect 9062 7470 9338 7512
rect 9062 7430 9180 7470
rect 9220 7430 9338 7470
rect 9062 7388 9338 7430
rect 9462 7470 9738 7512
rect 9462 7430 9580 7470
rect 9620 7430 9738 7470
rect 9462 7388 9738 7430
rect 9862 7470 10138 7512
rect 9862 7430 9980 7470
rect 10020 7430 10138 7470
rect 9862 7388 10138 7430
rect 10262 7470 10538 7512
rect 10262 7430 10380 7470
rect 10420 7430 10538 7470
rect 10262 7388 10538 7430
rect 10662 7470 10938 7512
rect 10662 7430 10780 7470
rect 10820 7430 10938 7470
rect 10662 7388 10938 7430
rect 11062 7470 11338 7512
rect 11062 7430 11180 7470
rect 11220 7430 11338 7470
rect 11062 7388 11338 7430
rect 11462 7470 11738 7512
rect 11462 7430 11580 7470
rect 11620 7430 11738 7470
rect 11462 7388 11738 7430
rect 11862 7470 12138 7512
rect 11862 7430 11980 7470
rect 12020 7430 12138 7470
rect 11862 7388 12138 7430
rect 12262 7470 12538 7512
rect 12262 7430 12380 7470
rect 12420 7430 12538 7470
rect 12262 7388 12538 7430
rect 12662 7470 12938 7512
rect 12662 7430 12780 7470
rect 12820 7430 12938 7470
rect 12662 7388 12938 7430
rect 13062 7470 13338 7512
rect 13062 7430 13180 7470
rect 13220 7430 13338 7470
rect 13062 7388 13338 7430
rect 13462 7470 13738 7512
rect 13462 7430 13580 7470
rect 13620 7430 13738 7470
rect 13462 7388 13738 7430
rect 13862 7470 14138 7512
rect 13862 7430 13980 7470
rect 14020 7430 14138 7470
rect 13862 7388 14138 7430
rect 14262 7470 14538 7512
rect 14262 7430 14380 7470
rect 14420 7430 14538 7470
rect 14262 7388 14538 7430
rect 14662 7470 14938 7512
rect 14662 7430 14780 7470
rect 14820 7430 14938 7470
rect 14662 7388 14938 7430
rect 15062 7470 15338 7512
rect 15062 7430 15180 7470
rect 15220 7430 15338 7470
rect 15062 7388 15338 7430
rect 15462 7470 16000 7512
rect 15462 7430 15580 7470
rect 15620 7430 16000 7470
rect 15462 7388 16000 7430
rect 0 6900 16000 7388
rect 0 6012 16000 6500
rect 0 5970 538 6012
rect 0 5930 380 5970
rect 420 5930 538 5970
rect 0 5888 538 5930
rect 662 5970 938 6012
rect 662 5930 780 5970
rect 820 5930 938 5970
rect 662 5888 938 5930
rect 1062 5970 1338 6012
rect 1062 5930 1180 5970
rect 1220 5930 1338 5970
rect 1062 5888 1338 5930
rect 1462 5970 1738 6012
rect 1462 5930 1580 5970
rect 1620 5930 1738 5970
rect 1462 5888 1738 5930
rect 1862 5970 2138 6012
rect 1862 5930 1980 5970
rect 2020 5930 2138 5970
rect 1862 5888 2138 5930
rect 2262 5970 2538 6012
rect 2262 5930 2380 5970
rect 2420 5930 2538 5970
rect 2262 5888 2538 5930
rect 2662 5970 2938 6012
rect 2662 5930 2780 5970
rect 2820 5930 2938 5970
rect 2662 5888 2938 5930
rect 3062 5970 3338 6012
rect 3062 5930 3180 5970
rect 3220 5930 3338 5970
rect 3062 5888 3338 5930
rect 3462 5970 3738 6012
rect 3462 5930 3580 5970
rect 3620 5930 3738 5970
rect 3462 5888 3738 5930
rect 3862 5970 4138 6012
rect 3862 5930 3980 5970
rect 4020 5930 4138 5970
rect 3862 5888 4138 5930
rect 4262 5970 4538 6012
rect 4262 5930 4380 5970
rect 4420 5930 4538 5970
rect 4262 5888 4538 5930
rect 4662 5970 4938 6012
rect 4662 5930 4780 5970
rect 4820 5930 4938 5970
rect 4662 5888 4938 5930
rect 5062 5970 5338 6012
rect 5062 5930 5180 5970
rect 5220 5930 5338 5970
rect 5062 5888 5338 5930
rect 5462 5970 5738 6012
rect 5462 5930 5580 5970
rect 5620 5930 5738 5970
rect 5462 5888 5738 5930
rect 5862 5970 6138 6012
rect 5862 5930 5980 5970
rect 6020 5930 6138 5970
rect 5862 5888 6138 5930
rect 6262 5970 6538 6012
rect 6262 5930 6380 5970
rect 6420 5930 6538 5970
rect 6262 5888 6538 5930
rect 6662 5970 6938 6012
rect 6662 5930 6780 5970
rect 6820 5930 6938 5970
rect 6662 5888 6938 5930
rect 7062 5970 7338 6012
rect 7062 5930 7180 5970
rect 7220 5930 7338 5970
rect 7062 5888 7338 5930
rect 7462 5970 7738 6012
rect 7462 5930 7580 5970
rect 7620 5930 7738 5970
rect 7462 5888 7738 5930
rect 7862 5970 8138 6012
rect 7862 5930 7980 5970
rect 8020 5930 8138 5970
rect 7862 5888 8138 5930
rect 8262 5970 8538 6012
rect 8262 5930 8380 5970
rect 8420 5930 8538 5970
rect 8262 5888 8538 5930
rect 8662 5970 8938 6012
rect 8662 5930 8780 5970
rect 8820 5930 8938 5970
rect 8662 5888 8938 5930
rect 9062 5970 9338 6012
rect 9062 5930 9180 5970
rect 9220 5930 9338 5970
rect 9062 5888 9338 5930
rect 9462 5970 9738 6012
rect 9462 5930 9580 5970
rect 9620 5930 9738 5970
rect 9462 5888 9738 5930
rect 9862 5970 10138 6012
rect 9862 5930 9980 5970
rect 10020 5930 10138 5970
rect 9862 5888 10138 5930
rect 10262 5970 10538 6012
rect 10262 5930 10380 5970
rect 10420 5930 10538 5970
rect 10262 5888 10538 5930
rect 10662 5970 10938 6012
rect 10662 5930 10780 5970
rect 10820 5930 10938 5970
rect 10662 5888 10938 5930
rect 11062 5970 11338 6012
rect 11062 5930 11180 5970
rect 11220 5930 11338 5970
rect 11062 5888 11338 5930
rect 11462 5970 11738 6012
rect 11462 5930 11580 5970
rect 11620 5930 11738 5970
rect 11462 5888 11738 5930
rect 11862 5970 12138 6012
rect 11862 5930 11980 5970
rect 12020 5930 12138 5970
rect 11862 5888 12138 5930
rect 12262 5970 12538 6012
rect 12262 5930 12380 5970
rect 12420 5930 12538 5970
rect 12262 5888 12538 5930
rect 12662 5970 12938 6012
rect 12662 5930 12780 5970
rect 12820 5930 12938 5970
rect 12662 5888 12938 5930
rect 13062 5970 13338 6012
rect 13062 5930 13180 5970
rect 13220 5930 13338 5970
rect 13062 5888 13338 5930
rect 13462 5970 13738 6012
rect 13462 5930 13580 5970
rect 13620 5930 13738 5970
rect 13462 5888 13738 5930
rect 13862 5970 14138 6012
rect 13862 5930 13980 5970
rect 14020 5930 14138 5970
rect 13862 5888 14138 5930
rect 14262 5970 14538 6012
rect 14262 5930 14380 5970
rect 14420 5930 14538 5970
rect 14262 5888 14538 5930
rect 14662 5970 14938 6012
rect 14662 5930 14780 5970
rect 14820 5930 14938 5970
rect 14662 5888 14938 5930
rect 15062 5970 15338 6012
rect 15062 5930 15180 5970
rect 15220 5930 15338 5970
rect 15062 5888 15338 5930
rect 15462 5970 16000 6012
rect 15462 5930 15580 5970
rect 15620 5930 16000 5970
rect 15462 5888 16000 5930
rect 0 5612 16000 5888
rect 0 5570 538 5612
rect 0 5530 380 5570
rect 420 5530 538 5570
rect 0 5488 538 5530
rect 662 5570 938 5612
rect 662 5530 780 5570
rect 820 5530 938 5570
rect 662 5488 938 5530
rect 1062 5570 1338 5612
rect 1062 5530 1180 5570
rect 1220 5530 1338 5570
rect 1062 5488 1338 5530
rect 1462 5570 1738 5612
rect 1462 5530 1580 5570
rect 1620 5530 1738 5570
rect 1462 5488 1738 5530
rect 1862 5570 2138 5612
rect 1862 5530 1980 5570
rect 2020 5530 2138 5570
rect 1862 5488 2138 5530
rect 2262 5570 2538 5612
rect 2262 5530 2380 5570
rect 2420 5530 2538 5570
rect 2262 5488 2538 5530
rect 2662 5570 2938 5612
rect 2662 5530 2780 5570
rect 2820 5530 2938 5570
rect 2662 5488 2938 5530
rect 3062 5570 3338 5612
rect 3062 5530 3180 5570
rect 3220 5530 3338 5570
rect 3062 5488 3338 5530
rect 3462 5570 3738 5612
rect 3462 5530 3580 5570
rect 3620 5530 3738 5570
rect 3462 5488 3738 5530
rect 3862 5570 4138 5612
rect 3862 5530 3980 5570
rect 4020 5530 4138 5570
rect 3862 5488 4138 5530
rect 4262 5570 4538 5612
rect 4262 5530 4380 5570
rect 4420 5530 4538 5570
rect 4262 5488 4538 5530
rect 4662 5570 4938 5612
rect 4662 5530 4780 5570
rect 4820 5530 4938 5570
rect 4662 5488 4938 5530
rect 5062 5570 5338 5612
rect 5062 5530 5180 5570
rect 5220 5530 5338 5570
rect 5062 5488 5338 5530
rect 5462 5570 5738 5612
rect 5462 5530 5580 5570
rect 5620 5530 5738 5570
rect 5462 5488 5738 5530
rect 5862 5570 6138 5612
rect 5862 5530 5980 5570
rect 6020 5530 6138 5570
rect 5862 5488 6138 5530
rect 6262 5570 6538 5612
rect 6262 5530 6380 5570
rect 6420 5530 6538 5570
rect 6262 5488 6538 5530
rect 6662 5570 6938 5612
rect 6662 5530 6780 5570
rect 6820 5530 6938 5570
rect 6662 5488 6938 5530
rect 7062 5570 7338 5612
rect 7062 5530 7180 5570
rect 7220 5530 7338 5570
rect 7062 5488 7338 5530
rect 7462 5570 7738 5612
rect 7462 5530 7580 5570
rect 7620 5530 7738 5570
rect 7462 5488 7738 5530
rect 7862 5570 8138 5612
rect 7862 5530 7980 5570
rect 8020 5530 8138 5570
rect 7862 5488 8138 5530
rect 8262 5570 8538 5612
rect 8262 5530 8380 5570
rect 8420 5530 8538 5570
rect 8262 5488 8538 5530
rect 8662 5570 8938 5612
rect 8662 5530 8780 5570
rect 8820 5530 8938 5570
rect 8662 5488 8938 5530
rect 9062 5570 9338 5612
rect 9062 5530 9180 5570
rect 9220 5530 9338 5570
rect 9062 5488 9338 5530
rect 9462 5570 9738 5612
rect 9462 5530 9580 5570
rect 9620 5530 9738 5570
rect 9462 5488 9738 5530
rect 9862 5570 10138 5612
rect 9862 5530 9980 5570
rect 10020 5530 10138 5570
rect 9862 5488 10138 5530
rect 10262 5570 10538 5612
rect 10262 5530 10380 5570
rect 10420 5530 10538 5570
rect 10262 5488 10538 5530
rect 10662 5570 10938 5612
rect 10662 5530 10780 5570
rect 10820 5530 10938 5570
rect 10662 5488 10938 5530
rect 11062 5570 11338 5612
rect 11062 5530 11180 5570
rect 11220 5530 11338 5570
rect 11062 5488 11338 5530
rect 11462 5570 11738 5612
rect 11462 5530 11580 5570
rect 11620 5530 11738 5570
rect 11462 5488 11738 5530
rect 11862 5570 12138 5612
rect 11862 5530 11980 5570
rect 12020 5530 12138 5570
rect 11862 5488 12138 5530
rect 12262 5570 12538 5612
rect 12262 5530 12380 5570
rect 12420 5530 12538 5570
rect 12262 5488 12538 5530
rect 12662 5570 12938 5612
rect 12662 5530 12780 5570
rect 12820 5530 12938 5570
rect 12662 5488 12938 5530
rect 13062 5570 13338 5612
rect 13062 5530 13180 5570
rect 13220 5530 13338 5570
rect 13062 5488 13338 5530
rect 13462 5570 13738 5612
rect 13462 5530 13580 5570
rect 13620 5530 13738 5570
rect 13462 5488 13738 5530
rect 13862 5570 14138 5612
rect 13862 5530 13980 5570
rect 14020 5530 14138 5570
rect 13862 5488 14138 5530
rect 14262 5570 14538 5612
rect 14262 5530 14380 5570
rect 14420 5530 14538 5570
rect 14262 5488 14538 5530
rect 14662 5570 14938 5612
rect 14662 5530 14780 5570
rect 14820 5530 14938 5570
rect 14662 5488 14938 5530
rect 15062 5570 15338 5612
rect 15062 5530 15180 5570
rect 15220 5530 15338 5570
rect 15062 5488 15338 5530
rect 15462 5570 16000 5612
rect 15462 5530 15580 5570
rect 15620 5530 16000 5570
rect 15462 5488 16000 5530
rect 0 5212 16000 5488
rect 0 5170 538 5212
rect 0 5130 380 5170
rect 420 5130 538 5170
rect 0 5088 538 5130
rect 662 5170 938 5212
rect 662 5130 780 5170
rect 820 5130 938 5170
rect 662 5088 938 5130
rect 1062 5170 1338 5212
rect 1062 5130 1180 5170
rect 1220 5130 1338 5170
rect 1062 5088 1338 5130
rect 1462 5170 1738 5212
rect 1462 5130 1580 5170
rect 1620 5130 1738 5170
rect 1462 5088 1738 5130
rect 1862 5170 2138 5212
rect 1862 5130 1980 5170
rect 2020 5130 2138 5170
rect 1862 5088 2138 5130
rect 2262 5170 2538 5212
rect 2262 5130 2380 5170
rect 2420 5130 2538 5170
rect 2262 5088 2538 5130
rect 2662 5170 2938 5212
rect 2662 5130 2780 5170
rect 2820 5130 2938 5170
rect 2662 5088 2938 5130
rect 3062 5170 3338 5212
rect 3062 5130 3180 5170
rect 3220 5130 3338 5170
rect 3062 5088 3338 5130
rect 3462 5170 3738 5212
rect 3462 5130 3580 5170
rect 3620 5130 3738 5170
rect 3462 5088 3738 5130
rect 3862 5170 4138 5212
rect 3862 5130 3980 5170
rect 4020 5130 4138 5170
rect 3862 5088 4138 5130
rect 4262 5170 4538 5212
rect 4262 5130 4380 5170
rect 4420 5130 4538 5170
rect 4262 5088 4538 5130
rect 4662 5170 4938 5212
rect 4662 5130 4780 5170
rect 4820 5130 4938 5170
rect 4662 5088 4938 5130
rect 5062 5170 5338 5212
rect 5062 5130 5180 5170
rect 5220 5130 5338 5170
rect 5062 5088 5338 5130
rect 5462 5170 5738 5212
rect 5462 5130 5580 5170
rect 5620 5130 5738 5170
rect 5462 5088 5738 5130
rect 5862 5170 6138 5212
rect 5862 5130 5980 5170
rect 6020 5130 6138 5170
rect 5862 5088 6138 5130
rect 6262 5170 6538 5212
rect 6262 5130 6380 5170
rect 6420 5130 6538 5170
rect 6262 5088 6538 5130
rect 6662 5170 6938 5212
rect 6662 5130 6780 5170
rect 6820 5130 6938 5170
rect 6662 5088 6938 5130
rect 7062 5170 7338 5212
rect 7062 5130 7180 5170
rect 7220 5130 7338 5170
rect 7062 5088 7338 5130
rect 7462 5170 7738 5212
rect 7462 5130 7580 5170
rect 7620 5130 7738 5170
rect 7462 5088 7738 5130
rect 7862 5170 8138 5212
rect 7862 5130 7980 5170
rect 8020 5130 8138 5170
rect 7862 5088 8138 5130
rect 8262 5170 8538 5212
rect 8262 5130 8380 5170
rect 8420 5130 8538 5170
rect 8262 5088 8538 5130
rect 8662 5170 8938 5212
rect 8662 5130 8780 5170
rect 8820 5130 8938 5170
rect 8662 5088 8938 5130
rect 9062 5170 9338 5212
rect 9062 5130 9180 5170
rect 9220 5130 9338 5170
rect 9062 5088 9338 5130
rect 9462 5170 9738 5212
rect 9462 5130 9580 5170
rect 9620 5130 9738 5170
rect 9462 5088 9738 5130
rect 9862 5170 10138 5212
rect 9862 5130 9980 5170
rect 10020 5130 10138 5170
rect 9862 5088 10138 5130
rect 10262 5170 10538 5212
rect 10262 5130 10380 5170
rect 10420 5130 10538 5170
rect 10262 5088 10538 5130
rect 10662 5170 10938 5212
rect 10662 5130 10780 5170
rect 10820 5130 10938 5170
rect 10662 5088 10938 5130
rect 11062 5170 11338 5212
rect 11062 5130 11180 5170
rect 11220 5130 11338 5170
rect 11062 5088 11338 5130
rect 11462 5170 11738 5212
rect 11462 5130 11580 5170
rect 11620 5130 11738 5170
rect 11462 5088 11738 5130
rect 11862 5170 12138 5212
rect 11862 5130 11980 5170
rect 12020 5130 12138 5170
rect 11862 5088 12138 5130
rect 12262 5170 12538 5212
rect 12262 5130 12380 5170
rect 12420 5130 12538 5170
rect 12262 5088 12538 5130
rect 12662 5170 12938 5212
rect 12662 5130 12780 5170
rect 12820 5130 12938 5170
rect 12662 5088 12938 5130
rect 13062 5170 13338 5212
rect 13062 5130 13180 5170
rect 13220 5130 13338 5170
rect 13062 5088 13338 5130
rect 13462 5170 13738 5212
rect 13462 5130 13580 5170
rect 13620 5130 13738 5170
rect 13462 5088 13738 5130
rect 13862 5170 14138 5212
rect 13862 5130 13980 5170
rect 14020 5130 14138 5170
rect 13862 5088 14138 5130
rect 14262 5170 14538 5212
rect 14262 5130 14380 5170
rect 14420 5130 14538 5170
rect 14262 5088 14538 5130
rect 14662 5170 14938 5212
rect 14662 5130 14780 5170
rect 14820 5130 14938 5170
rect 14662 5088 14938 5130
rect 15062 5170 15338 5212
rect 15062 5130 15180 5170
rect 15220 5130 15338 5170
rect 15062 5088 15338 5130
rect 15462 5170 16000 5212
rect 15462 5130 15580 5170
rect 15620 5130 16000 5170
rect 15462 5088 16000 5130
rect 0 4812 16000 5088
rect 0 4770 538 4812
rect 0 4730 380 4770
rect 420 4730 538 4770
rect 0 4688 538 4730
rect 662 4770 938 4812
rect 662 4730 780 4770
rect 820 4730 938 4770
rect 662 4688 938 4730
rect 1062 4770 1338 4812
rect 1062 4730 1180 4770
rect 1220 4730 1338 4770
rect 1062 4688 1338 4730
rect 1462 4770 1738 4812
rect 1462 4730 1580 4770
rect 1620 4730 1738 4770
rect 1462 4688 1738 4730
rect 1862 4770 2138 4812
rect 1862 4730 1980 4770
rect 2020 4730 2138 4770
rect 1862 4688 2138 4730
rect 2262 4770 2538 4812
rect 2262 4730 2380 4770
rect 2420 4730 2538 4770
rect 2262 4688 2538 4730
rect 2662 4770 2938 4812
rect 2662 4730 2780 4770
rect 2820 4730 2938 4770
rect 2662 4688 2938 4730
rect 3062 4770 3338 4812
rect 3062 4730 3180 4770
rect 3220 4730 3338 4770
rect 3062 4688 3338 4730
rect 3462 4770 3738 4812
rect 3462 4730 3580 4770
rect 3620 4730 3738 4770
rect 3462 4688 3738 4730
rect 3862 4770 4138 4812
rect 3862 4730 3980 4770
rect 4020 4730 4138 4770
rect 3862 4688 4138 4730
rect 4262 4770 4538 4812
rect 4262 4730 4380 4770
rect 4420 4730 4538 4770
rect 4262 4688 4538 4730
rect 4662 4770 4938 4812
rect 4662 4730 4780 4770
rect 4820 4730 4938 4770
rect 4662 4688 4938 4730
rect 5062 4770 5338 4812
rect 5062 4730 5180 4770
rect 5220 4730 5338 4770
rect 5062 4688 5338 4730
rect 5462 4770 5738 4812
rect 5462 4730 5580 4770
rect 5620 4730 5738 4770
rect 5462 4688 5738 4730
rect 5862 4770 6138 4812
rect 5862 4730 5980 4770
rect 6020 4730 6138 4770
rect 5862 4688 6138 4730
rect 6262 4770 6538 4812
rect 6262 4730 6380 4770
rect 6420 4730 6538 4770
rect 6262 4688 6538 4730
rect 6662 4770 6938 4812
rect 6662 4730 6780 4770
rect 6820 4730 6938 4770
rect 6662 4688 6938 4730
rect 7062 4770 7338 4812
rect 7062 4730 7180 4770
rect 7220 4730 7338 4770
rect 7062 4688 7338 4730
rect 7462 4770 7738 4812
rect 7462 4730 7580 4770
rect 7620 4730 7738 4770
rect 7462 4688 7738 4730
rect 7862 4770 8138 4812
rect 7862 4730 7980 4770
rect 8020 4730 8138 4770
rect 7862 4688 8138 4730
rect 8262 4770 8538 4812
rect 8262 4730 8380 4770
rect 8420 4730 8538 4770
rect 8262 4688 8538 4730
rect 8662 4770 8938 4812
rect 8662 4730 8780 4770
rect 8820 4730 8938 4770
rect 8662 4688 8938 4730
rect 9062 4770 9338 4812
rect 9062 4730 9180 4770
rect 9220 4730 9338 4770
rect 9062 4688 9338 4730
rect 9462 4770 9738 4812
rect 9462 4730 9580 4770
rect 9620 4730 9738 4770
rect 9462 4688 9738 4730
rect 9862 4770 10138 4812
rect 9862 4730 9980 4770
rect 10020 4730 10138 4770
rect 9862 4688 10138 4730
rect 10262 4770 10538 4812
rect 10262 4730 10380 4770
rect 10420 4730 10538 4770
rect 10262 4688 10538 4730
rect 10662 4770 10938 4812
rect 10662 4730 10780 4770
rect 10820 4730 10938 4770
rect 10662 4688 10938 4730
rect 11062 4770 11338 4812
rect 11062 4730 11180 4770
rect 11220 4730 11338 4770
rect 11062 4688 11338 4730
rect 11462 4770 11738 4812
rect 11462 4730 11580 4770
rect 11620 4730 11738 4770
rect 11462 4688 11738 4730
rect 11862 4770 12138 4812
rect 11862 4730 11980 4770
rect 12020 4730 12138 4770
rect 11862 4688 12138 4730
rect 12262 4770 12538 4812
rect 12262 4730 12380 4770
rect 12420 4730 12538 4770
rect 12262 4688 12538 4730
rect 12662 4770 12938 4812
rect 12662 4730 12780 4770
rect 12820 4730 12938 4770
rect 12662 4688 12938 4730
rect 13062 4770 13338 4812
rect 13062 4730 13180 4770
rect 13220 4730 13338 4770
rect 13062 4688 13338 4730
rect 13462 4770 13738 4812
rect 13462 4730 13580 4770
rect 13620 4730 13738 4770
rect 13462 4688 13738 4730
rect 13862 4770 14138 4812
rect 13862 4730 13980 4770
rect 14020 4730 14138 4770
rect 13862 4688 14138 4730
rect 14262 4770 14538 4812
rect 14262 4730 14380 4770
rect 14420 4730 14538 4770
rect 14262 4688 14538 4730
rect 14662 4770 14938 4812
rect 14662 4730 14780 4770
rect 14820 4730 14938 4770
rect 14662 4688 14938 4730
rect 15062 4770 15338 4812
rect 15062 4730 15180 4770
rect 15220 4730 15338 4770
rect 15062 4688 15338 4730
rect 15462 4770 16000 4812
rect 15462 4730 15580 4770
rect 15620 4730 16000 4770
rect 15462 4688 16000 4730
rect 0 4412 16000 4688
rect 0 4370 538 4412
rect 0 4330 380 4370
rect 420 4330 538 4370
rect 0 4288 538 4330
rect 662 4370 938 4412
rect 662 4330 780 4370
rect 820 4330 938 4370
rect 662 4288 938 4330
rect 1062 4370 1338 4412
rect 1062 4330 1180 4370
rect 1220 4330 1338 4370
rect 1062 4288 1338 4330
rect 1462 4370 1738 4412
rect 1462 4330 1580 4370
rect 1620 4330 1738 4370
rect 1462 4288 1738 4330
rect 1862 4370 2138 4412
rect 1862 4330 1980 4370
rect 2020 4330 2138 4370
rect 1862 4288 2138 4330
rect 2262 4370 2538 4412
rect 2262 4330 2380 4370
rect 2420 4330 2538 4370
rect 2262 4288 2538 4330
rect 2662 4370 2938 4412
rect 2662 4330 2780 4370
rect 2820 4330 2938 4370
rect 2662 4288 2938 4330
rect 3062 4370 3338 4412
rect 3062 4330 3180 4370
rect 3220 4330 3338 4370
rect 3062 4288 3338 4330
rect 3462 4370 3738 4412
rect 3462 4330 3580 4370
rect 3620 4330 3738 4370
rect 3462 4288 3738 4330
rect 3862 4370 4138 4412
rect 3862 4330 3980 4370
rect 4020 4330 4138 4370
rect 3862 4288 4138 4330
rect 4262 4370 4538 4412
rect 4262 4330 4380 4370
rect 4420 4330 4538 4370
rect 4262 4288 4538 4330
rect 4662 4370 4938 4412
rect 4662 4330 4780 4370
rect 4820 4330 4938 4370
rect 4662 4288 4938 4330
rect 5062 4370 5338 4412
rect 5062 4330 5180 4370
rect 5220 4330 5338 4370
rect 5062 4288 5338 4330
rect 5462 4370 5738 4412
rect 5462 4330 5580 4370
rect 5620 4330 5738 4370
rect 5462 4288 5738 4330
rect 5862 4370 6138 4412
rect 5862 4330 5980 4370
rect 6020 4330 6138 4370
rect 5862 4288 6138 4330
rect 6262 4370 6538 4412
rect 6262 4330 6380 4370
rect 6420 4330 6538 4370
rect 6262 4288 6538 4330
rect 6662 4370 6938 4412
rect 6662 4330 6780 4370
rect 6820 4330 6938 4370
rect 6662 4288 6938 4330
rect 7062 4370 7338 4412
rect 7062 4330 7180 4370
rect 7220 4330 7338 4370
rect 7062 4288 7338 4330
rect 7462 4370 7738 4412
rect 7462 4330 7580 4370
rect 7620 4330 7738 4370
rect 7462 4288 7738 4330
rect 7862 4370 8138 4412
rect 7862 4330 7980 4370
rect 8020 4330 8138 4370
rect 7862 4288 8138 4330
rect 8262 4370 8538 4412
rect 8262 4330 8380 4370
rect 8420 4330 8538 4370
rect 8262 4288 8538 4330
rect 8662 4370 8938 4412
rect 8662 4330 8780 4370
rect 8820 4330 8938 4370
rect 8662 4288 8938 4330
rect 9062 4370 9338 4412
rect 9062 4330 9180 4370
rect 9220 4330 9338 4370
rect 9062 4288 9338 4330
rect 9462 4370 9738 4412
rect 9462 4330 9580 4370
rect 9620 4330 9738 4370
rect 9462 4288 9738 4330
rect 9862 4370 10138 4412
rect 9862 4330 9980 4370
rect 10020 4330 10138 4370
rect 9862 4288 10138 4330
rect 10262 4370 10538 4412
rect 10262 4330 10380 4370
rect 10420 4330 10538 4370
rect 10262 4288 10538 4330
rect 10662 4370 10938 4412
rect 10662 4330 10780 4370
rect 10820 4330 10938 4370
rect 10662 4288 10938 4330
rect 11062 4370 11338 4412
rect 11062 4330 11180 4370
rect 11220 4330 11338 4370
rect 11062 4288 11338 4330
rect 11462 4370 11738 4412
rect 11462 4330 11580 4370
rect 11620 4330 11738 4370
rect 11462 4288 11738 4330
rect 11862 4370 12138 4412
rect 11862 4330 11980 4370
rect 12020 4330 12138 4370
rect 11862 4288 12138 4330
rect 12262 4370 12538 4412
rect 12262 4330 12380 4370
rect 12420 4330 12538 4370
rect 12262 4288 12538 4330
rect 12662 4370 12938 4412
rect 12662 4330 12780 4370
rect 12820 4330 12938 4370
rect 12662 4288 12938 4330
rect 13062 4370 13338 4412
rect 13062 4330 13180 4370
rect 13220 4330 13338 4370
rect 13062 4288 13338 4330
rect 13462 4370 13738 4412
rect 13462 4330 13580 4370
rect 13620 4330 13738 4370
rect 13462 4288 13738 4330
rect 13862 4370 14138 4412
rect 13862 4330 13980 4370
rect 14020 4330 14138 4370
rect 13862 4288 14138 4330
rect 14262 4370 14538 4412
rect 14262 4330 14380 4370
rect 14420 4330 14538 4370
rect 14262 4288 14538 4330
rect 14662 4370 14938 4412
rect 14662 4330 14780 4370
rect 14820 4330 14938 4370
rect 14662 4288 14938 4330
rect 15062 4370 15338 4412
rect 15062 4330 15180 4370
rect 15220 4330 15338 4370
rect 15062 4288 15338 4330
rect 15462 4370 16000 4412
rect 15462 4330 15580 4370
rect 15620 4330 16000 4370
rect 15462 4288 16000 4330
rect 0 4012 16000 4288
rect 0 3970 538 4012
rect 0 3930 380 3970
rect 420 3930 538 3970
rect 0 3888 538 3930
rect 662 3970 938 4012
rect 662 3930 780 3970
rect 820 3930 938 3970
rect 662 3888 938 3930
rect 1062 3970 1338 4012
rect 1062 3930 1180 3970
rect 1220 3930 1338 3970
rect 1062 3888 1338 3930
rect 1462 3970 1738 4012
rect 1462 3930 1580 3970
rect 1620 3930 1738 3970
rect 1462 3888 1738 3930
rect 1862 3970 2138 4012
rect 1862 3930 1980 3970
rect 2020 3930 2138 3970
rect 1862 3888 2138 3930
rect 2262 3970 2538 4012
rect 2262 3930 2380 3970
rect 2420 3930 2538 3970
rect 2262 3888 2538 3930
rect 2662 3970 2938 4012
rect 2662 3930 2780 3970
rect 2820 3930 2938 3970
rect 2662 3888 2938 3930
rect 3062 3970 3338 4012
rect 3062 3930 3180 3970
rect 3220 3930 3338 3970
rect 3062 3888 3338 3930
rect 3462 3970 3738 4012
rect 3462 3930 3580 3970
rect 3620 3930 3738 3970
rect 3462 3888 3738 3930
rect 3862 3970 4138 4012
rect 3862 3930 3980 3970
rect 4020 3930 4138 3970
rect 3862 3888 4138 3930
rect 4262 3970 4538 4012
rect 4262 3930 4380 3970
rect 4420 3930 4538 3970
rect 4262 3888 4538 3930
rect 4662 3970 4938 4012
rect 4662 3930 4780 3970
rect 4820 3930 4938 3970
rect 4662 3888 4938 3930
rect 5062 3970 5338 4012
rect 5062 3930 5180 3970
rect 5220 3930 5338 3970
rect 5062 3888 5338 3930
rect 5462 3970 5738 4012
rect 5462 3930 5580 3970
rect 5620 3930 5738 3970
rect 5462 3888 5738 3930
rect 5862 3970 6138 4012
rect 5862 3930 5980 3970
rect 6020 3930 6138 3970
rect 5862 3888 6138 3930
rect 6262 3970 6538 4012
rect 6262 3930 6380 3970
rect 6420 3930 6538 3970
rect 6262 3888 6538 3930
rect 6662 3970 6938 4012
rect 6662 3930 6780 3970
rect 6820 3930 6938 3970
rect 6662 3888 6938 3930
rect 7062 3970 7338 4012
rect 7062 3930 7180 3970
rect 7220 3930 7338 3970
rect 7062 3888 7338 3930
rect 7462 3970 7738 4012
rect 7462 3930 7580 3970
rect 7620 3930 7738 3970
rect 7462 3888 7738 3930
rect 7862 3970 8138 4012
rect 7862 3930 7980 3970
rect 8020 3930 8138 3970
rect 7862 3888 8138 3930
rect 8262 3970 8538 4012
rect 8262 3930 8380 3970
rect 8420 3930 8538 3970
rect 8262 3888 8538 3930
rect 8662 3970 8938 4012
rect 8662 3930 8780 3970
rect 8820 3930 8938 3970
rect 8662 3888 8938 3930
rect 9062 3970 9338 4012
rect 9062 3930 9180 3970
rect 9220 3930 9338 3970
rect 9062 3888 9338 3930
rect 9462 3970 9738 4012
rect 9462 3930 9580 3970
rect 9620 3930 9738 3970
rect 9462 3888 9738 3930
rect 9862 3970 10138 4012
rect 9862 3930 9980 3970
rect 10020 3930 10138 3970
rect 9862 3888 10138 3930
rect 10262 3970 10538 4012
rect 10262 3930 10380 3970
rect 10420 3930 10538 3970
rect 10262 3888 10538 3930
rect 10662 3970 10938 4012
rect 10662 3930 10780 3970
rect 10820 3930 10938 3970
rect 10662 3888 10938 3930
rect 11062 3970 11338 4012
rect 11062 3930 11180 3970
rect 11220 3930 11338 3970
rect 11062 3888 11338 3930
rect 11462 3970 11738 4012
rect 11462 3930 11580 3970
rect 11620 3930 11738 3970
rect 11462 3888 11738 3930
rect 11862 3970 12138 4012
rect 11862 3930 11980 3970
rect 12020 3930 12138 3970
rect 11862 3888 12138 3930
rect 12262 3970 12538 4012
rect 12262 3930 12380 3970
rect 12420 3930 12538 3970
rect 12262 3888 12538 3930
rect 12662 3970 12938 4012
rect 12662 3930 12780 3970
rect 12820 3930 12938 3970
rect 12662 3888 12938 3930
rect 13062 3970 13338 4012
rect 13062 3930 13180 3970
rect 13220 3930 13338 3970
rect 13062 3888 13338 3930
rect 13462 3970 13738 4012
rect 13462 3930 13580 3970
rect 13620 3930 13738 3970
rect 13462 3888 13738 3930
rect 13862 3970 14138 4012
rect 13862 3930 13980 3970
rect 14020 3930 14138 3970
rect 13862 3888 14138 3930
rect 14262 3970 14538 4012
rect 14262 3930 14380 3970
rect 14420 3930 14538 3970
rect 14262 3888 14538 3930
rect 14662 3970 14938 4012
rect 14662 3930 14780 3970
rect 14820 3930 14938 3970
rect 14662 3888 14938 3930
rect 15062 3970 15338 4012
rect 15062 3930 15180 3970
rect 15220 3930 15338 3970
rect 15062 3888 15338 3930
rect 15462 3970 16000 4012
rect 15462 3930 15580 3970
rect 15620 3930 16000 3970
rect 15462 3888 16000 3930
rect 0 3612 16000 3888
rect 0 3570 538 3612
rect 0 3530 380 3570
rect 420 3530 538 3570
rect 0 3488 538 3530
rect 662 3570 938 3612
rect 662 3530 780 3570
rect 820 3530 938 3570
rect 662 3488 938 3530
rect 1062 3570 1338 3612
rect 1062 3530 1180 3570
rect 1220 3530 1338 3570
rect 1062 3488 1338 3530
rect 1462 3570 1738 3612
rect 1462 3530 1580 3570
rect 1620 3530 1738 3570
rect 1462 3488 1738 3530
rect 1862 3570 2138 3612
rect 1862 3530 1980 3570
rect 2020 3530 2138 3570
rect 1862 3488 2138 3530
rect 2262 3570 2538 3612
rect 2262 3530 2380 3570
rect 2420 3530 2538 3570
rect 2262 3488 2538 3530
rect 2662 3570 2938 3612
rect 2662 3530 2780 3570
rect 2820 3530 2938 3570
rect 2662 3488 2938 3530
rect 3062 3570 3338 3612
rect 3062 3530 3180 3570
rect 3220 3530 3338 3570
rect 3062 3488 3338 3530
rect 3462 3570 3738 3612
rect 3462 3530 3580 3570
rect 3620 3530 3738 3570
rect 3462 3488 3738 3530
rect 3862 3570 4138 3612
rect 3862 3530 3980 3570
rect 4020 3530 4138 3570
rect 3862 3488 4138 3530
rect 4262 3570 4538 3612
rect 4262 3530 4380 3570
rect 4420 3530 4538 3570
rect 4262 3488 4538 3530
rect 4662 3570 4938 3612
rect 4662 3530 4780 3570
rect 4820 3530 4938 3570
rect 4662 3488 4938 3530
rect 5062 3570 5338 3612
rect 5062 3530 5180 3570
rect 5220 3530 5338 3570
rect 5062 3488 5338 3530
rect 5462 3570 5738 3612
rect 5462 3530 5580 3570
rect 5620 3530 5738 3570
rect 5462 3488 5738 3530
rect 5862 3570 6138 3612
rect 5862 3530 5980 3570
rect 6020 3530 6138 3570
rect 5862 3488 6138 3530
rect 6262 3570 6538 3612
rect 6262 3530 6380 3570
rect 6420 3530 6538 3570
rect 6262 3488 6538 3530
rect 6662 3570 6938 3612
rect 6662 3530 6780 3570
rect 6820 3530 6938 3570
rect 6662 3488 6938 3530
rect 7062 3570 7338 3612
rect 7062 3530 7180 3570
rect 7220 3530 7338 3570
rect 7062 3488 7338 3530
rect 7462 3570 7738 3612
rect 7462 3530 7580 3570
rect 7620 3530 7738 3570
rect 7462 3488 7738 3530
rect 7862 3570 8138 3612
rect 7862 3530 7980 3570
rect 8020 3530 8138 3570
rect 7862 3488 8138 3530
rect 8262 3570 8538 3612
rect 8262 3530 8380 3570
rect 8420 3530 8538 3570
rect 8262 3488 8538 3530
rect 8662 3570 8938 3612
rect 8662 3530 8780 3570
rect 8820 3530 8938 3570
rect 8662 3488 8938 3530
rect 9062 3570 9338 3612
rect 9062 3530 9180 3570
rect 9220 3530 9338 3570
rect 9062 3488 9338 3530
rect 9462 3570 9738 3612
rect 9462 3530 9580 3570
rect 9620 3530 9738 3570
rect 9462 3488 9738 3530
rect 9862 3570 10138 3612
rect 9862 3530 9980 3570
rect 10020 3530 10138 3570
rect 9862 3488 10138 3530
rect 10262 3570 10538 3612
rect 10262 3530 10380 3570
rect 10420 3530 10538 3570
rect 10262 3488 10538 3530
rect 10662 3570 10938 3612
rect 10662 3530 10780 3570
rect 10820 3530 10938 3570
rect 10662 3488 10938 3530
rect 11062 3570 11338 3612
rect 11062 3530 11180 3570
rect 11220 3530 11338 3570
rect 11062 3488 11338 3530
rect 11462 3570 11738 3612
rect 11462 3530 11580 3570
rect 11620 3530 11738 3570
rect 11462 3488 11738 3530
rect 11862 3570 12138 3612
rect 11862 3530 11980 3570
rect 12020 3530 12138 3570
rect 11862 3488 12138 3530
rect 12262 3570 12538 3612
rect 12262 3530 12380 3570
rect 12420 3530 12538 3570
rect 12262 3488 12538 3530
rect 12662 3570 12938 3612
rect 12662 3530 12780 3570
rect 12820 3530 12938 3570
rect 12662 3488 12938 3530
rect 13062 3570 13338 3612
rect 13062 3530 13180 3570
rect 13220 3530 13338 3570
rect 13062 3488 13338 3530
rect 13462 3570 13738 3612
rect 13462 3530 13580 3570
rect 13620 3530 13738 3570
rect 13462 3488 13738 3530
rect 13862 3570 14138 3612
rect 13862 3530 13980 3570
rect 14020 3530 14138 3570
rect 13862 3488 14138 3530
rect 14262 3570 14538 3612
rect 14262 3530 14380 3570
rect 14420 3530 14538 3570
rect 14262 3488 14538 3530
rect 14662 3570 14938 3612
rect 14662 3530 14780 3570
rect 14820 3530 14938 3570
rect 14662 3488 14938 3530
rect 15062 3570 15338 3612
rect 15062 3530 15180 3570
rect 15220 3530 15338 3570
rect 15062 3488 15338 3530
rect 15462 3570 16000 3612
rect 15462 3530 15580 3570
rect 15620 3530 16000 3570
rect 15462 3488 16000 3530
rect 0 3212 16000 3488
rect 0 3170 538 3212
rect 0 3130 380 3170
rect 420 3130 538 3170
rect 0 3088 538 3130
rect 662 3170 938 3212
rect 662 3130 780 3170
rect 820 3130 938 3170
rect 662 3088 938 3130
rect 1062 3170 1338 3212
rect 1062 3130 1180 3170
rect 1220 3130 1338 3170
rect 1062 3088 1338 3130
rect 1462 3170 1738 3212
rect 1462 3130 1580 3170
rect 1620 3130 1738 3170
rect 1462 3088 1738 3130
rect 1862 3170 2138 3212
rect 1862 3130 1980 3170
rect 2020 3130 2138 3170
rect 1862 3088 2138 3130
rect 2262 3170 2538 3212
rect 2262 3130 2380 3170
rect 2420 3130 2538 3170
rect 2262 3088 2538 3130
rect 2662 3170 2938 3212
rect 2662 3130 2780 3170
rect 2820 3130 2938 3170
rect 2662 3088 2938 3130
rect 3062 3170 3338 3212
rect 3062 3130 3180 3170
rect 3220 3130 3338 3170
rect 3062 3088 3338 3130
rect 3462 3170 3738 3212
rect 3462 3130 3580 3170
rect 3620 3130 3738 3170
rect 3462 3088 3738 3130
rect 3862 3170 4138 3212
rect 3862 3130 3980 3170
rect 4020 3130 4138 3170
rect 3862 3088 4138 3130
rect 4262 3170 4538 3212
rect 4262 3130 4380 3170
rect 4420 3130 4538 3170
rect 4262 3088 4538 3130
rect 4662 3170 4938 3212
rect 4662 3130 4780 3170
rect 4820 3130 4938 3170
rect 4662 3088 4938 3130
rect 5062 3170 5338 3212
rect 5062 3130 5180 3170
rect 5220 3130 5338 3170
rect 5062 3088 5338 3130
rect 5462 3170 5738 3212
rect 5462 3130 5580 3170
rect 5620 3130 5738 3170
rect 5462 3088 5738 3130
rect 5862 3170 6138 3212
rect 5862 3130 5980 3170
rect 6020 3130 6138 3170
rect 5862 3088 6138 3130
rect 6262 3170 6538 3212
rect 6262 3130 6380 3170
rect 6420 3130 6538 3170
rect 6262 3088 6538 3130
rect 6662 3170 6938 3212
rect 6662 3130 6780 3170
rect 6820 3130 6938 3170
rect 6662 3088 6938 3130
rect 7062 3170 7338 3212
rect 7062 3130 7180 3170
rect 7220 3130 7338 3170
rect 7062 3088 7338 3130
rect 7462 3170 7738 3212
rect 7462 3130 7580 3170
rect 7620 3130 7738 3170
rect 7462 3088 7738 3130
rect 7862 3170 8138 3212
rect 7862 3130 7980 3170
rect 8020 3130 8138 3170
rect 7862 3088 8138 3130
rect 8262 3170 8538 3212
rect 8262 3130 8380 3170
rect 8420 3130 8538 3170
rect 8262 3088 8538 3130
rect 8662 3170 8938 3212
rect 8662 3130 8780 3170
rect 8820 3130 8938 3170
rect 8662 3088 8938 3130
rect 9062 3170 9338 3212
rect 9062 3130 9180 3170
rect 9220 3130 9338 3170
rect 9062 3088 9338 3130
rect 9462 3170 9738 3212
rect 9462 3130 9580 3170
rect 9620 3130 9738 3170
rect 9462 3088 9738 3130
rect 9862 3170 10138 3212
rect 9862 3130 9980 3170
rect 10020 3130 10138 3170
rect 9862 3088 10138 3130
rect 10262 3170 10538 3212
rect 10262 3130 10380 3170
rect 10420 3130 10538 3170
rect 10262 3088 10538 3130
rect 10662 3170 10938 3212
rect 10662 3130 10780 3170
rect 10820 3130 10938 3170
rect 10662 3088 10938 3130
rect 11062 3170 11338 3212
rect 11062 3130 11180 3170
rect 11220 3130 11338 3170
rect 11062 3088 11338 3130
rect 11462 3170 11738 3212
rect 11462 3130 11580 3170
rect 11620 3130 11738 3170
rect 11462 3088 11738 3130
rect 11862 3170 12138 3212
rect 11862 3130 11980 3170
rect 12020 3130 12138 3170
rect 11862 3088 12138 3130
rect 12262 3170 12538 3212
rect 12262 3130 12380 3170
rect 12420 3130 12538 3170
rect 12262 3088 12538 3130
rect 12662 3170 12938 3212
rect 12662 3130 12780 3170
rect 12820 3130 12938 3170
rect 12662 3088 12938 3130
rect 13062 3170 13338 3212
rect 13062 3130 13180 3170
rect 13220 3130 13338 3170
rect 13062 3088 13338 3130
rect 13462 3170 13738 3212
rect 13462 3130 13580 3170
rect 13620 3130 13738 3170
rect 13462 3088 13738 3130
rect 13862 3170 14138 3212
rect 13862 3130 13980 3170
rect 14020 3130 14138 3170
rect 13862 3088 14138 3130
rect 14262 3170 14538 3212
rect 14262 3130 14380 3170
rect 14420 3130 14538 3170
rect 14262 3088 14538 3130
rect 14662 3170 14938 3212
rect 14662 3130 14780 3170
rect 14820 3130 14938 3170
rect 14662 3088 14938 3130
rect 15062 3170 15338 3212
rect 15062 3130 15180 3170
rect 15220 3130 15338 3170
rect 15062 3088 15338 3130
rect 15462 3170 16000 3212
rect 15462 3130 15580 3170
rect 15620 3130 16000 3170
rect 15462 3088 16000 3130
rect 0 2812 16000 3088
rect 0 2770 538 2812
rect 0 2730 380 2770
rect 420 2730 538 2770
rect 0 2688 538 2730
rect 662 2770 938 2812
rect 662 2730 780 2770
rect 820 2730 938 2770
rect 662 2688 938 2730
rect 1062 2770 1338 2812
rect 1062 2730 1180 2770
rect 1220 2730 1338 2770
rect 1062 2688 1338 2730
rect 1462 2770 1738 2812
rect 1462 2730 1580 2770
rect 1620 2730 1738 2770
rect 1462 2688 1738 2730
rect 1862 2770 2138 2812
rect 1862 2730 1980 2770
rect 2020 2730 2138 2770
rect 1862 2688 2138 2730
rect 2262 2770 2538 2812
rect 2262 2730 2380 2770
rect 2420 2730 2538 2770
rect 2262 2688 2538 2730
rect 2662 2770 2938 2812
rect 2662 2730 2780 2770
rect 2820 2730 2938 2770
rect 2662 2688 2938 2730
rect 3062 2770 3338 2812
rect 3062 2730 3180 2770
rect 3220 2730 3338 2770
rect 3062 2688 3338 2730
rect 3462 2770 3738 2812
rect 3462 2730 3580 2770
rect 3620 2730 3738 2770
rect 3462 2688 3738 2730
rect 3862 2770 4138 2812
rect 3862 2730 3980 2770
rect 4020 2730 4138 2770
rect 3862 2688 4138 2730
rect 4262 2770 4538 2812
rect 4262 2730 4380 2770
rect 4420 2730 4538 2770
rect 4262 2688 4538 2730
rect 4662 2770 4938 2812
rect 4662 2730 4780 2770
rect 4820 2730 4938 2770
rect 4662 2688 4938 2730
rect 5062 2770 5338 2812
rect 5062 2730 5180 2770
rect 5220 2730 5338 2770
rect 5062 2688 5338 2730
rect 5462 2770 5738 2812
rect 5462 2730 5580 2770
rect 5620 2730 5738 2770
rect 5462 2688 5738 2730
rect 5862 2770 6138 2812
rect 5862 2730 5980 2770
rect 6020 2730 6138 2770
rect 5862 2688 6138 2730
rect 6262 2770 6538 2812
rect 6262 2730 6380 2770
rect 6420 2730 6538 2770
rect 6262 2688 6538 2730
rect 6662 2770 6938 2812
rect 6662 2730 6780 2770
rect 6820 2730 6938 2770
rect 6662 2688 6938 2730
rect 7062 2770 7338 2812
rect 7062 2730 7180 2770
rect 7220 2730 7338 2770
rect 7062 2688 7338 2730
rect 7462 2770 7738 2812
rect 7462 2730 7580 2770
rect 7620 2730 7738 2770
rect 7462 2688 7738 2730
rect 7862 2770 8138 2812
rect 7862 2730 7980 2770
rect 8020 2730 8138 2770
rect 7862 2688 8138 2730
rect 8262 2770 8538 2812
rect 8262 2730 8380 2770
rect 8420 2730 8538 2770
rect 8262 2688 8538 2730
rect 8662 2770 8938 2812
rect 8662 2730 8780 2770
rect 8820 2730 8938 2770
rect 8662 2688 8938 2730
rect 9062 2770 9338 2812
rect 9062 2730 9180 2770
rect 9220 2730 9338 2770
rect 9062 2688 9338 2730
rect 9462 2770 9738 2812
rect 9462 2730 9580 2770
rect 9620 2730 9738 2770
rect 9462 2688 9738 2730
rect 9862 2770 10138 2812
rect 9862 2730 9980 2770
rect 10020 2730 10138 2770
rect 9862 2688 10138 2730
rect 10262 2770 10538 2812
rect 10262 2730 10380 2770
rect 10420 2730 10538 2770
rect 10262 2688 10538 2730
rect 10662 2770 10938 2812
rect 10662 2730 10780 2770
rect 10820 2730 10938 2770
rect 10662 2688 10938 2730
rect 11062 2770 11338 2812
rect 11062 2730 11180 2770
rect 11220 2730 11338 2770
rect 11062 2688 11338 2730
rect 11462 2770 11738 2812
rect 11462 2730 11580 2770
rect 11620 2730 11738 2770
rect 11462 2688 11738 2730
rect 11862 2770 12138 2812
rect 11862 2730 11980 2770
rect 12020 2730 12138 2770
rect 11862 2688 12138 2730
rect 12262 2770 12538 2812
rect 12262 2730 12380 2770
rect 12420 2730 12538 2770
rect 12262 2688 12538 2730
rect 12662 2770 12938 2812
rect 12662 2730 12780 2770
rect 12820 2730 12938 2770
rect 12662 2688 12938 2730
rect 13062 2770 13338 2812
rect 13062 2730 13180 2770
rect 13220 2730 13338 2770
rect 13062 2688 13338 2730
rect 13462 2770 13738 2812
rect 13462 2730 13580 2770
rect 13620 2730 13738 2770
rect 13462 2688 13738 2730
rect 13862 2770 14138 2812
rect 13862 2730 13980 2770
rect 14020 2730 14138 2770
rect 13862 2688 14138 2730
rect 14262 2770 14538 2812
rect 14262 2730 14380 2770
rect 14420 2730 14538 2770
rect 14262 2688 14538 2730
rect 14662 2770 14938 2812
rect 14662 2730 14780 2770
rect 14820 2730 14938 2770
rect 14662 2688 14938 2730
rect 15062 2770 15338 2812
rect 15062 2730 15180 2770
rect 15220 2730 15338 2770
rect 15062 2688 15338 2730
rect 15462 2770 16000 2812
rect 15462 2730 15580 2770
rect 15620 2730 16000 2770
rect 15462 2688 16000 2730
rect 0 2412 16000 2688
rect 0 2370 538 2412
rect 0 2330 380 2370
rect 420 2330 538 2370
rect 0 2288 538 2330
rect 662 2370 938 2412
rect 662 2330 780 2370
rect 820 2330 938 2370
rect 662 2288 938 2330
rect 1062 2370 1338 2412
rect 1062 2330 1180 2370
rect 1220 2330 1338 2370
rect 1062 2288 1338 2330
rect 1462 2370 1738 2412
rect 1462 2330 1580 2370
rect 1620 2330 1738 2370
rect 1462 2288 1738 2330
rect 1862 2370 2138 2412
rect 1862 2330 1980 2370
rect 2020 2330 2138 2370
rect 1862 2288 2138 2330
rect 2262 2370 2538 2412
rect 2262 2330 2380 2370
rect 2420 2330 2538 2370
rect 2262 2288 2538 2330
rect 2662 2370 2938 2412
rect 2662 2330 2780 2370
rect 2820 2330 2938 2370
rect 2662 2288 2938 2330
rect 3062 2370 3338 2412
rect 3062 2330 3180 2370
rect 3220 2330 3338 2370
rect 3062 2288 3338 2330
rect 3462 2370 3738 2412
rect 3462 2330 3580 2370
rect 3620 2330 3738 2370
rect 3462 2288 3738 2330
rect 3862 2370 4138 2412
rect 3862 2330 3980 2370
rect 4020 2330 4138 2370
rect 3862 2288 4138 2330
rect 4262 2370 4538 2412
rect 4262 2330 4380 2370
rect 4420 2330 4538 2370
rect 4262 2288 4538 2330
rect 4662 2370 4938 2412
rect 4662 2330 4780 2370
rect 4820 2330 4938 2370
rect 4662 2288 4938 2330
rect 5062 2370 5338 2412
rect 5062 2330 5180 2370
rect 5220 2330 5338 2370
rect 5062 2288 5338 2330
rect 5462 2370 5738 2412
rect 5462 2330 5580 2370
rect 5620 2330 5738 2370
rect 5462 2288 5738 2330
rect 5862 2370 6138 2412
rect 5862 2330 5980 2370
rect 6020 2330 6138 2370
rect 5862 2288 6138 2330
rect 6262 2370 6538 2412
rect 6262 2330 6380 2370
rect 6420 2330 6538 2370
rect 6262 2288 6538 2330
rect 6662 2370 6938 2412
rect 6662 2330 6780 2370
rect 6820 2330 6938 2370
rect 6662 2288 6938 2330
rect 7062 2370 7338 2412
rect 7062 2330 7180 2370
rect 7220 2330 7338 2370
rect 7062 2288 7338 2330
rect 7462 2370 7738 2412
rect 7462 2330 7580 2370
rect 7620 2330 7738 2370
rect 7462 2288 7738 2330
rect 7862 2370 8138 2412
rect 7862 2330 7980 2370
rect 8020 2330 8138 2370
rect 7862 2288 8138 2330
rect 8262 2370 8538 2412
rect 8262 2330 8380 2370
rect 8420 2330 8538 2370
rect 8262 2288 8538 2330
rect 8662 2370 8938 2412
rect 8662 2330 8780 2370
rect 8820 2330 8938 2370
rect 8662 2288 8938 2330
rect 9062 2370 9338 2412
rect 9062 2330 9180 2370
rect 9220 2330 9338 2370
rect 9062 2288 9338 2330
rect 9462 2370 9738 2412
rect 9462 2330 9580 2370
rect 9620 2330 9738 2370
rect 9462 2288 9738 2330
rect 9862 2370 10138 2412
rect 9862 2330 9980 2370
rect 10020 2330 10138 2370
rect 9862 2288 10138 2330
rect 10262 2370 10538 2412
rect 10262 2330 10380 2370
rect 10420 2330 10538 2370
rect 10262 2288 10538 2330
rect 10662 2370 10938 2412
rect 10662 2330 10780 2370
rect 10820 2330 10938 2370
rect 10662 2288 10938 2330
rect 11062 2370 11338 2412
rect 11062 2330 11180 2370
rect 11220 2330 11338 2370
rect 11062 2288 11338 2330
rect 11462 2370 11738 2412
rect 11462 2330 11580 2370
rect 11620 2330 11738 2370
rect 11462 2288 11738 2330
rect 11862 2370 12138 2412
rect 11862 2330 11980 2370
rect 12020 2330 12138 2370
rect 11862 2288 12138 2330
rect 12262 2370 12538 2412
rect 12262 2330 12380 2370
rect 12420 2330 12538 2370
rect 12262 2288 12538 2330
rect 12662 2370 12938 2412
rect 12662 2330 12780 2370
rect 12820 2330 12938 2370
rect 12662 2288 12938 2330
rect 13062 2370 13338 2412
rect 13062 2330 13180 2370
rect 13220 2330 13338 2370
rect 13062 2288 13338 2330
rect 13462 2370 13738 2412
rect 13462 2330 13580 2370
rect 13620 2330 13738 2370
rect 13462 2288 13738 2330
rect 13862 2370 14138 2412
rect 13862 2330 13980 2370
rect 14020 2330 14138 2370
rect 13862 2288 14138 2330
rect 14262 2370 14538 2412
rect 14262 2330 14380 2370
rect 14420 2330 14538 2370
rect 14262 2288 14538 2330
rect 14662 2370 14938 2412
rect 14662 2330 14780 2370
rect 14820 2330 14938 2370
rect 14662 2288 14938 2330
rect 15062 2370 15338 2412
rect 15062 2330 15180 2370
rect 15220 2330 15338 2370
rect 15062 2288 15338 2330
rect 15462 2370 16000 2412
rect 15462 2330 15580 2370
rect 15620 2330 16000 2370
rect 15462 2288 16000 2330
rect 0 2012 16000 2288
rect 0 1970 538 2012
rect 0 1930 380 1970
rect 420 1930 538 1970
rect 0 1888 538 1930
rect 662 1970 938 2012
rect 662 1930 780 1970
rect 820 1930 938 1970
rect 662 1888 938 1930
rect 1062 1970 1338 2012
rect 1062 1930 1180 1970
rect 1220 1930 1338 1970
rect 1062 1888 1338 1930
rect 1462 1970 1738 2012
rect 1462 1930 1580 1970
rect 1620 1930 1738 1970
rect 1462 1888 1738 1930
rect 1862 1970 2138 2012
rect 1862 1930 1980 1970
rect 2020 1930 2138 1970
rect 1862 1888 2138 1930
rect 2262 1970 2538 2012
rect 2262 1930 2380 1970
rect 2420 1930 2538 1970
rect 2262 1888 2538 1930
rect 2662 1970 2938 2012
rect 2662 1930 2780 1970
rect 2820 1930 2938 1970
rect 2662 1888 2938 1930
rect 3062 1970 3338 2012
rect 3062 1930 3180 1970
rect 3220 1930 3338 1970
rect 3062 1888 3338 1930
rect 3462 1970 3738 2012
rect 3462 1930 3580 1970
rect 3620 1930 3738 1970
rect 3462 1888 3738 1930
rect 3862 1970 4138 2012
rect 3862 1930 3980 1970
rect 4020 1930 4138 1970
rect 3862 1888 4138 1930
rect 4262 1970 4538 2012
rect 4262 1930 4380 1970
rect 4420 1930 4538 1970
rect 4262 1888 4538 1930
rect 4662 1970 4938 2012
rect 4662 1930 4780 1970
rect 4820 1930 4938 1970
rect 4662 1888 4938 1930
rect 5062 1970 5338 2012
rect 5062 1930 5180 1970
rect 5220 1930 5338 1970
rect 5062 1888 5338 1930
rect 5462 1970 5738 2012
rect 5462 1930 5580 1970
rect 5620 1930 5738 1970
rect 5462 1888 5738 1930
rect 5862 1970 6138 2012
rect 5862 1930 5980 1970
rect 6020 1930 6138 1970
rect 5862 1888 6138 1930
rect 6262 1970 6538 2012
rect 6262 1930 6380 1970
rect 6420 1930 6538 1970
rect 6262 1888 6538 1930
rect 6662 1970 6938 2012
rect 6662 1930 6780 1970
rect 6820 1930 6938 1970
rect 6662 1888 6938 1930
rect 7062 1970 7338 2012
rect 7062 1930 7180 1970
rect 7220 1930 7338 1970
rect 7062 1888 7338 1930
rect 7462 1970 7738 2012
rect 7462 1930 7580 1970
rect 7620 1930 7738 1970
rect 7462 1888 7738 1930
rect 7862 1970 8138 2012
rect 7862 1930 7980 1970
rect 8020 1930 8138 1970
rect 7862 1888 8138 1930
rect 8262 1970 8538 2012
rect 8262 1930 8380 1970
rect 8420 1930 8538 1970
rect 8262 1888 8538 1930
rect 8662 1970 8938 2012
rect 8662 1930 8780 1970
rect 8820 1930 8938 1970
rect 8662 1888 8938 1930
rect 9062 1970 9338 2012
rect 9062 1930 9180 1970
rect 9220 1930 9338 1970
rect 9062 1888 9338 1930
rect 9462 1970 9738 2012
rect 9462 1930 9580 1970
rect 9620 1930 9738 1970
rect 9462 1888 9738 1930
rect 9862 1970 10138 2012
rect 9862 1930 9980 1970
rect 10020 1930 10138 1970
rect 9862 1888 10138 1930
rect 10262 1970 10538 2012
rect 10262 1930 10380 1970
rect 10420 1930 10538 1970
rect 10262 1888 10538 1930
rect 10662 1970 10938 2012
rect 10662 1930 10780 1970
rect 10820 1930 10938 1970
rect 10662 1888 10938 1930
rect 11062 1970 11338 2012
rect 11062 1930 11180 1970
rect 11220 1930 11338 1970
rect 11062 1888 11338 1930
rect 11462 1970 11738 2012
rect 11462 1930 11580 1970
rect 11620 1930 11738 1970
rect 11462 1888 11738 1930
rect 11862 1970 12138 2012
rect 11862 1930 11980 1970
rect 12020 1930 12138 1970
rect 11862 1888 12138 1930
rect 12262 1970 12538 2012
rect 12262 1930 12380 1970
rect 12420 1930 12538 1970
rect 12262 1888 12538 1930
rect 12662 1970 12938 2012
rect 12662 1930 12780 1970
rect 12820 1930 12938 1970
rect 12662 1888 12938 1930
rect 13062 1970 13338 2012
rect 13062 1930 13180 1970
rect 13220 1930 13338 1970
rect 13062 1888 13338 1930
rect 13462 1970 13738 2012
rect 13462 1930 13580 1970
rect 13620 1930 13738 1970
rect 13462 1888 13738 1930
rect 13862 1970 14138 2012
rect 13862 1930 13980 1970
rect 14020 1930 14138 1970
rect 13862 1888 14138 1930
rect 14262 1970 14538 2012
rect 14262 1930 14380 1970
rect 14420 1930 14538 1970
rect 14262 1888 14538 1930
rect 14662 1970 14938 2012
rect 14662 1930 14780 1970
rect 14820 1930 14938 1970
rect 14662 1888 14938 1930
rect 15062 1970 15338 2012
rect 15062 1930 15180 1970
rect 15220 1930 15338 1970
rect 15062 1888 15338 1930
rect 15462 1970 16000 2012
rect 15462 1930 15580 1970
rect 15620 1930 16000 1970
rect 15462 1888 16000 1930
rect 0 1400 16000 1888
rect 1000 520 15000 600
rect 1000 480 1180 520
rect 1220 480 1580 520
rect 1620 480 1980 520
rect 2020 480 2380 520
rect 2420 480 2780 520
rect 2820 480 3180 520
rect 3220 480 3580 520
rect 3620 480 3980 520
rect 4020 480 4380 520
rect 4420 480 4780 520
rect 4820 480 5180 520
rect 5220 480 5580 520
rect 5620 480 5980 520
rect 6020 480 6380 520
rect 6420 480 6780 520
rect 6820 480 7180 520
rect 7220 480 7580 520
rect 7620 480 7980 520
rect 8020 480 8380 520
rect 8420 480 8780 520
rect 8820 480 9180 520
rect 9220 480 9580 520
rect 9620 480 9980 520
rect 10020 480 10380 520
rect 10420 480 10780 520
rect 10820 480 11180 520
rect 11220 480 11580 520
rect 11620 480 11980 520
rect 12020 480 12380 520
rect 12420 480 12780 520
rect 12820 480 13180 520
rect 13220 480 13580 520
rect 13620 480 13980 520
rect 14020 480 14380 520
rect 14420 480 14780 520
rect 14820 480 15000 520
rect 1000 362 15000 480
rect 1000 238 1138 362
rect 1262 238 1538 362
rect 1662 238 1938 362
rect 2062 238 2338 362
rect 2462 238 2738 362
rect 2862 238 3138 362
rect 3262 238 3538 362
rect 3662 238 3938 362
rect 4062 238 4338 362
rect 4462 238 4738 362
rect 4862 238 5138 362
rect 5262 238 5538 362
rect 5662 238 5938 362
rect 6062 238 6338 362
rect 6462 238 6738 362
rect 6862 238 7138 362
rect 7262 238 7538 362
rect 7662 238 7938 362
rect 8062 238 8338 362
rect 8462 238 8738 362
rect 8862 238 9138 362
rect 9262 238 9538 362
rect 9662 238 9938 362
rect 10062 238 10338 362
rect 10462 238 10738 362
rect 10862 238 11138 362
rect 11262 238 11538 362
rect 11662 238 11938 362
rect 12062 238 12338 362
rect 12462 238 12738 362
rect 12862 238 13138 362
rect 13262 238 13538 362
rect 13662 238 13938 362
rect 14062 238 14338 362
rect 14462 238 14738 362
rect 14862 238 15000 362
rect 1000 120 15000 238
rect 1000 80 1180 120
rect 1220 80 1580 120
rect 1620 80 1980 120
rect 2020 80 2380 120
rect 2420 80 2780 120
rect 2820 80 3180 120
rect 3220 80 3580 120
rect 3620 80 3980 120
rect 4020 80 4380 120
rect 4420 80 4780 120
rect 4820 80 5180 120
rect 5220 80 5580 120
rect 5620 80 5980 120
rect 6020 80 6380 120
rect 6420 80 6780 120
rect 6820 80 7180 120
rect 7220 80 7580 120
rect 7620 80 7980 120
rect 8020 80 8380 120
rect 8420 80 8780 120
rect 8820 80 9180 120
rect 9220 80 9580 120
rect 9620 80 9980 120
rect 10020 80 10380 120
rect 10420 80 10780 120
rect 10820 80 11180 120
rect 11220 80 11580 120
rect 11620 80 11980 120
rect 12020 80 12380 120
rect 12420 80 12780 120
rect 12820 80 13180 120
rect 13220 80 13580 120
rect 13620 80 13980 120
rect 14020 80 14380 120
rect 14420 80 14780 120
rect 14820 80 15000 120
rect 1000 0 15000 80
<< via5 >>
rect 538 34938 662 35062
rect 938 34938 1062 35062
rect 1338 34938 1462 35062
rect 1738 34938 1862 35062
rect 2138 34938 2262 35062
rect 2538 34938 2662 35062
rect 2938 34938 3062 35062
rect 3338 34938 3462 35062
rect 3738 34938 3862 35062
rect 4138 34938 4262 35062
rect 4538 34938 4662 35062
rect 4938 34938 5062 35062
rect 5338 34938 5462 35062
rect 5738 34938 5862 35062
rect 6138 34938 6262 35062
rect 6538 34938 6662 35062
rect 6938 34938 7062 35062
rect 7338 34938 7462 35062
rect 7738 34938 7862 35062
rect 8138 34938 8262 35062
rect 8538 34938 8662 35062
rect 8938 34938 9062 35062
rect 9338 34938 9462 35062
rect 9738 34938 9862 35062
rect 10138 34938 10262 35062
rect 10538 34938 10662 35062
rect 10938 34938 11062 35062
rect 11338 34938 11462 35062
rect 11738 34938 11862 35062
rect 12138 34938 12262 35062
rect 12538 34938 12662 35062
rect 12938 34938 13062 35062
rect 13338 34938 13462 35062
rect 13738 34938 13862 35062
rect 14138 34938 14262 35062
rect 14538 34938 14662 35062
rect 14938 34938 15062 35062
rect 15338 34938 15462 35062
rect 538 34538 662 34662
rect 938 34538 1062 34662
rect 1338 34538 1462 34662
rect 1738 34538 1862 34662
rect 2138 34538 2262 34662
rect 2538 34538 2662 34662
rect 2938 34538 3062 34662
rect 3338 34538 3462 34662
rect 3738 34538 3862 34662
rect 4138 34538 4262 34662
rect 4538 34538 4662 34662
rect 4938 34538 5062 34662
rect 5338 34538 5462 34662
rect 5738 34538 5862 34662
rect 6138 34538 6262 34662
rect 6538 34538 6662 34662
rect 6938 34538 7062 34662
rect 7338 34538 7462 34662
rect 7738 34538 7862 34662
rect 8138 34538 8262 34662
rect 8538 34538 8662 34662
rect 8938 34538 9062 34662
rect 9338 34538 9462 34662
rect 9738 34538 9862 34662
rect 10138 34538 10262 34662
rect 10538 34538 10662 34662
rect 10938 34538 11062 34662
rect 11338 34538 11462 34662
rect 11738 34538 11862 34662
rect 12138 34538 12262 34662
rect 12538 34538 12662 34662
rect 12938 34538 13062 34662
rect 13338 34538 13462 34662
rect 13738 34538 13862 34662
rect 14138 34538 14262 34662
rect 14538 34538 14662 34662
rect 14938 34538 15062 34662
rect 15338 34538 15462 34662
rect 538 34138 662 34262
rect 938 34138 1062 34262
rect 1338 34138 1462 34262
rect 1738 34138 1862 34262
rect 2138 34138 2262 34262
rect 2538 34138 2662 34262
rect 2938 34138 3062 34262
rect 3338 34138 3462 34262
rect 3738 34138 3862 34262
rect 4138 34138 4262 34262
rect 4538 34138 4662 34262
rect 4938 34138 5062 34262
rect 5338 34138 5462 34262
rect 5738 34138 5862 34262
rect 6138 34138 6262 34262
rect 6538 34138 6662 34262
rect 6938 34138 7062 34262
rect 7338 34138 7462 34262
rect 7738 34138 7862 34262
rect 8138 34138 8262 34262
rect 8538 34138 8662 34262
rect 8938 34138 9062 34262
rect 9338 34138 9462 34262
rect 9738 34138 9862 34262
rect 10138 34138 10262 34262
rect 10538 34138 10662 34262
rect 10938 34138 11062 34262
rect 11338 34138 11462 34262
rect 11738 34138 11862 34262
rect 12138 34138 12262 34262
rect 12538 34138 12662 34262
rect 12938 34138 13062 34262
rect 13338 34138 13462 34262
rect 13738 34138 13862 34262
rect 14138 34138 14262 34262
rect 14538 34138 14662 34262
rect 14938 34138 15062 34262
rect 15338 34138 15462 34262
rect 538 33738 662 33862
rect 938 33738 1062 33862
rect 1338 33738 1462 33862
rect 1738 33738 1862 33862
rect 2138 33738 2262 33862
rect 2538 33738 2662 33862
rect 2938 33738 3062 33862
rect 3338 33738 3462 33862
rect 3738 33738 3862 33862
rect 4138 33738 4262 33862
rect 4538 33738 4662 33862
rect 4938 33738 5062 33862
rect 5338 33738 5462 33862
rect 5738 33738 5862 33862
rect 6138 33738 6262 33862
rect 6538 33738 6662 33862
rect 6938 33738 7062 33862
rect 7338 33738 7462 33862
rect 7738 33738 7862 33862
rect 8138 33738 8262 33862
rect 8538 33738 8662 33862
rect 8938 33738 9062 33862
rect 9338 33738 9462 33862
rect 9738 33738 9862 33862
rect 10138 33738 10262 33862
rect 10538 33738 10662 33862
rect 10938 33738 11062 33862
rect 11338 33738 11462 33862
rect 11738 33738 11862 33862
rect 12138 33738 12262 33862
rect 12538 33738 12662 33862
rect 12938 33738 13062 33862
rect 13338 33738 13462 33862
rect 13738 33738 13862 33862
rect 14138 33738 14262 33862
rect 14538 33738 14662 33862
rect 14938 33738 15062 33862
rect 15338 33738 15462 33862
rect 538 33338 662 33462
rect 938 33338 1062 33462
rect 1338 33338 1462 33462
rect 1738 33338 1862 33462
rect 2138 33338 2262 33462
rect 2538 33338 2662 33462
rect 2938 33338 3062 33462
rect 3338 33338 3462 33462
rect 3738 33338 3862 33462
rect 4138 33338 4262 33462
rect 4538 33338 4662 33462
rect 4938 33338 5062 33462
rect 5338 33338 5462 33462
rect 5738 33338 5862 33462
rect 6138 33338 6262 33462
rect 6538 33338 6662 33462
rect 6938 33338 7062 33462
rect 7338 33338 7462 33462
rect 7738 33338 7862 33462
rect 8138 33338 8262 33462
rect 8538 33338 8662 33462
rect 8938 33338 9062 33462
rect 9338 33338 9462 33462
rect 9738 33338 9862 33462
rect 10138 33338 10262 33462
rect 10538 33338 10662 33462
rect 10938 33338 11062 33462
rect 11338 33338 11462 33462
rect 11738 33338 11862 33462
rect 12138 33338 12262 33462
rect 12538 33338 12662 33462
rect 12938 33338 13062 33462
rect 13338 33338 13462 33462
rect 13738 33338 13862 33462
rect 14138 33338 14262 33462
rect 14538 33338 14662 33462
rect 14938 33338 15062 33462
rect 15338 33338 15462 33462
rect 538 32938 662 33062
rect 938 32938 1062 33062
rect 1338 32938 1462 33062
rect 1738 32938 1862 33062
rect 2138 32938 2262 33062
rect 2538 32938 2662 33062
rect 2938 32938 3062 33062
rect 3338 32938 3462 33062
rect 3738 32938 3862 33062
rect 4138 32938 4262 33062
rect 4538 32938 4662 33062
rect 4938 32938 5062 33062
rect 5338 32938 5462 33062
rect 5738 32938 5862 33062
rect 6138 32938 6262 33062
rect 6538 32938 6662 33062
rect 6938 32938 7062 33062
rect 7338 32938 7462 33062
rect 7738 32938 7862 33062
rect 8138 32938 8262 33062
rect 8538 32938 8662 33062
rect 8938 32938 9062 33062
rect 9338 32938 9462 33062
rect 9738 32938 9862 33062
rect 10138 32938 10262 33062
rect 10538 32938 10662 33062
rect 10938 32938 11062 33062
rect 11338 32938 11462 33062
rect 11738 32938 11862 33062
rect 12138 32938 12262 33062
rect 12538 32938 12662 33062
rect 12938 32938 13062 33062
rect 13338 32938 13462 33062
rect 13738 32938 13862 33062
rect 14138 32938 14262 33062
rect 14538 32938 14662 33062
rect 14938 32938 15062 33062
rect 15338 32938 15462 33062
rect 538 32538 662 32662
rect 938 32538 1062 32662
rect 1338 32538 1462 32662
rect 1738 32538 1862 32662
rect 2138 32538 2262 32662
rect 2538 32538 2662 32662
rect 2938 32538 3062 32662
rect 3338 32538 3462 32662
rect 3738 32538 3862 32662
rect 4138 32538 4262 32662
rect 4538 32538 4662 32662
rect 4938 32538 5062 32662
rect 5338 32538 5462 32662
rect 5738 32538 5862 32662
rect 6138 32538 6262 32662
rect 6538 32538 6662 32662
rect 6938 32538 7062 32662
rect 7338 32538 7462 32662
rect 7738 32538 7862 32662
rect 8138 32538 8262 32662
rect 8538 32538 8662 32662
rect 8938 32538 9062 32662
rect 9338 32538 9462 32662
rect 9738 32538 9862 32662
rect 10138 32538 10262 32662
rect 10538 32538 10662 32662
rect 10938 32538 11062 32662
rect 11338 32538 11462 32662
rect 11738 32538 11862 32662
rect 12138 32538 12262 32662
rect 12538 32538 12662 32662
rect 12938 32538 13062 32662
rect 13338 32538 13462 32662
rect 13738 32538 13862 32662
rect 14138 32538 14262 32662
rect 14538 32538 14662 32662
rect 14938 32538 15062 32662
rect 15338 32538 15462 32662
rect 538 30938 662 31062
rect 938 30938 1062 31062
rect 1338 30938 1462 31062
rect 1738 30938 1862 31062
rect 2138 30938 2262 31062
rect 2538 30938 2662 31062
rect 2938 30938 3062 31062
rect 3338 30938 3462 31062
rect 3738 30938 3862 31062
rect 4138 30938 4262 31062
rect 4538 30938 4662 31062
rect 4938 30938 5062 31062
rect 5338 30938 5462 31062
rect 5738 30938 5862 31062
rect 6138 30938 6262 31062
rect 6538 30938 6662 31062
rect 6938 30938 7062 31062
rect 7338 30938 7462 31062
rect 7738 30938 7862 31062
rect 8138 30938 8262 31062
rect 8538 30938 8662 31062
rect 8938 30938 9062 31062
rect 9338 30938 9462 31062
rect 9738 30938 9862 31062
rect 10138 30938 10262 31062
rect 10538 30938 10662 31062
rect 10938 30938 11062 31062
rect 11338 30938 11462 31062
rect 11738 30938 11862 31062
rect 12138 30938 12262 31062
rect 12538 30938 12662 31062
rect 12938 30938 13062 31062
rect 13338 30938 13462 31062
rect 13738 30938 13862 31062
rect 14138 30938 14262 31062
rect 14538 30938 14662 31062
rect 14938 30938 15062 31062
rect 15338 30938 15462 31062
rect 538 30538 662 30662
rect 938 30538 1062 30662
rect 1338 30538 1462 30662
rect 1738 30538 1862 30662
rect 2138 30538 2262 30662
rect 2538 30538 2662 30662
rect 2938 30538 3062 30662
rect 3338 30538 3462 30662
rect 3738 30538 3862 30662
rect 4138 30538 4262 30662
rect 4538 30538 4662 30662
rect 4938 30538 5062 30662
rect 5338 30538 5462 30662
rect 5738 30538 5862 30662
rect 6138 30538 6262 30662
rect 6538 30538 6662 30662
rect 6938 30538 7062 30662
rect 7338 30538 7462 30662
rect 7738 30538 7862 30662
rect 8138 30538 8262 30662
rect 8538 30538 8662 30662
rect 8938 30538 9062 30662
rect 9338 30538 9462 30662
rect 9738 30538 9862 30662
rect 10138 30538 10262 30662
rect 10538 30538 10662 30662
rect 10938 30538 11062 30662
rect 11338 30538 11462 30662
rect 11738 30538 11862 30662
rect 12138 30538 12262 30662
rect 12538 30538 12662 30662
rect 12938 30538 13062 30662
rect 13338 30538 13462 30662
rect 13738 30538 13862 30662
rect 14138 30538 14262 30662
rect 14538 30538 14662 30662
rect 14938 30538 15062 30662
rect 15338 30538 15462 30662
rect 538 30138 662 30262
rect 938 30138 1062 30262
rect 1338 30138 1462 30262
rect 1738 30138 1862 30262
rect 2138 30138 2262 30262
rect 2538 30138 2662 30262
rect 2938 30138 3062 30262
rect 3338 30138 3462 30262
rect 3738 30138 3862 30262
rect 4138 30138 4262 30262
rect 4538 30138 4662 30262
rect 4938 30138 5062 30262
rect 5338 30138 5462 30262
rect 5738 30138 5862 30262
rect 6138 30138 6262 30262
rect 6538 30138 6662 30262
rect 6938 30138 7062 30262
rect 7338 30138 7462 30262
rect 7738 30138 7862 30262
rect 8138 30138 8262 30262
rect 8538 30138 8662 30262
rect 8938 30138 9062 30262
rect 9338 30138 9462 30262
rect 9738 30138 9862 30262
rect 10138 30138 10262 30262
rect 10538 30138 10662 30262
rect 10938 30138 11062 30262
rect 11338 30138 11462 30262
rect 11738 30138 11862 30262
rect 12138 30138 12262 30262
rect 12538 30138 12662 30262
rect 12938 30138 13062 30262
rect 13338 30138 13462 30262
rect 13738 30138 13862 30262
rect 14138 30138 14262 30262
rect 14538 30138 14662 30262
rect 14938 30138 15062 30262
rect 15338 30138 15462 30262
rect 538 29738 662 29862
rect 938 29738 1062 29862
rect 1338 29738 1462 29862
rect 1738 29738 1862 29862
rect 2138 29738 2262 29862
rect 2538 29738 2662 29862
rect 2938 29738 3062 29862
rect 3338 29738 3462 29862
rect 3738 29738 3862 29862
rect 4138 29738 4262 29862
rect 4538 29738 4662 29862
rect 4938 29738 5062 29862
rect 5338 29738 5462 29862
rect 5738 29738 5862 29862
rect 6138 29738 6262 29862
rect 6538 29738 6662 29862
rect 6938 29738 7062 29862
rect 7338 29738 7462 29862
rect 7738 29738 7862 29862
rect 8138 29738 8262 29862
rect 8538 29738 8662 29862
rect 8938 29738 9062 29862
rect 9338 29738 9462 29862
rect 9738 29738 9862 29862
rect 10138 29738 10262 29862
rect 10538 29738 10662 29862
rect 10938 29738 11062 29862
rect 11338 29738 11462 29862
rect 11738 29738 11862 29862
rect 12138 29738 12262 29862
rect 12538 29738 12662 29862
rect 12938 29738 13062 29862
rect 13338 29738 13462 29862
rect 13738 29738 13862 29862
rect 14138 29738 14262 29862
rect 14538 29738 14662 29862
rect 14938 29738 15062 29862
rect 15338 29738 15462 29862
rect 538 29338 662 29462
rect 938 29338 1062 29462
rect 1338 29338 1462 29462
rect 1738 29338 1862 29462
rect 2138 29338 2262 29462
rect 2538 29338 2662 29462
rect 2938 29338 3062 29462
rect 3338 29338 3462 29462
rect 3738 29338 3862 29462
rect 4138 29338 4262 29462
rect 4538 29338 4662 29462
rect 4938 29338 5062 29462
rect 5338 29338 5462 29462
rect 5738 29338 5862 29462
rect 6138 29338 6262 29462
rect 6538 29338 6662 29462
rect 6938 29338 7062 29462
rect 7338 29338 7462 29462
rect 7738 29338 7862 29462
rect 8138 29338 8262 29462
rect 8538 29338 8662 29462
rect 8938 29338 9062 29462
rect 9338 29338 9462 29462
rect 9738 29338 9862 29462
rect 10138 29338 10262 29462
rect 10538 29338 10662 29462
rect 10938 29338 11062 29462
rect 11338 29338 11462 29462
rect 11738 29338 11862 29462
rect 12138 29338 12262 29462
rect 12538 29338 12662 29462
rect 12938 29338 13062 29462
rect 13338 29338 13462 29462
rect 13738 29338 13862 29462
rect 14138 29338 14262 29462
rect 14538 29338 14662 29462
rect 14938 29338 15062 29462
rect 15338 29338 15462 29462
rect 538 28938 662 29062
rect 938 28938 1062 29062
rect 1338 28938 1462 29062
rect 1738 28938 1862 29062
rect 2138 28938 2262 29062
rect 2538 28938 2662 29062
rect 2938 28938 3062 29062
rect 3338 28938 3462 29062
rect 3738 28938 3862 29062
rect 4138 28938 4262 29062
rect 4538 28938 4662 29062
rect 4938 28938 5062 29062
rect 5338 28938 5462 29062
rect 5738 28938 5862 29062
rect 6138 28938 6262 29062
rect 6538 28938 6662 29062
rect 6938 28938 7062 29062
rect 7338 28938 7462 29062
rect 7738 28938 7862 29062
rect 8138 28938 8262 29062
rect 8538 28938 8662 29062
rect 8938 28938 9062 29062
rect 9338 28938 9462 29062
rect 9738 28938 9862 29062
rect 10138 28938 10262 29062
rect 10538 28938 10662 29062
rect 10938 28938 11062 29062
rect 11338 28938 11462 29062
rect 11738 28938 11862 29062
rect 12138 28938 12262 29062
rect 12538 28938 12662 29062
rect 12938 28938 13062 29062
rect 13338 28938 13462 29062
rect 13738 28938 13862 29062
rect 14138 28938 14262 29062
rect 14538 28938 14662 29062
rect 14938 28938 15062 29062
rect 15338 28938 15462 29062
rect 538 28538 662 28662
rect 938 28538 1062 28662
rect 1338 28538 1462 28662
rect 1738 28538 1862 28662
rect 2138 28538 2262 28662
rect 2538 28538 2662 28662
rect 2938 28538 3062 28662
rect 3338 28538 3462 28662
rect 3738 28538 3862 28662
rect 4138 28538 4262 28662
rect 4538 28538 4662 28662
rect 4938 28538 5062 28662
rect 5338 28538 5462 28662
rect 5738 28538 5862 28662
rect 6138 28538 6262 28662
rect 6538 28538 6662 28662
rect 6938 28538 7062 28662
rect 7338 28538 7462 28662
rect 7738 28538 7862 28662
rect 8138 28538 8262 28662
rect 8538 28538 8662 28662
rect 8938 28538 9062 28662
rect 9338 28538 9462 28662
rect 9738 28538 9862 28662
rect 10138 28538 10262 28662
rect 10538 28538 10662 28662
rect 10938 28538 11062 28662
rect 11338 28538 11462 28662
rect 11738 28538 11862 28662
rect 12138 28538 12262 28662
rect 12538 28538 12662 28662
rect 12938 28538 13062 28662
rect 13338 28538 13462 28662
rect 13738 28538 13862 28662
rect 14138 28538 14262 28662
rect 14538 28538 14662 28662
rect 14938 28538 15062 28662
rect 15338 28538 15462 28662
rect 538 26138 662 26262
rect 938 26138 1062 26262
rect 1338 26138 1462 26262
rect 1738 26138 1862 26262
rect 2138 26138 2262 26262
rect 2538 26138 2662 26262
rect 2938 26138 3062 26262
rect 3338 26138 3462 26262
rect 3738 26138 3862 26262
rect 4138 26138 4262 26262
rect 4538 26138 4662 26262
rect 4938 26138 5062 26262
rect 5338 26138 5462 26262
rect 5738 26138 5862 26262
rect 6138 26138 6262 26262
rect 6538 26138 6662 26262
rect 6938 26138 7062 26262
rect 7338 26138 7462 26262
rect 7738 26138 7862 26262
rect 8138 26138 8262 26262
rect 8538 26138 8662 26262
rect 8938 26138 9062 26262
rect 9338 26138 9462 26262
rect 9738 26138 9862 26262
rect 10138 26138 10262 26262
rect 10538 26138 10662 26262
rect 10938 26138 11062 26262
rect 11338 26138 11462 26262
rect 11738 26138 11862 26262
rect 12138 26138 12262 26262
rect 12538 26138 12662 26262
rect 12938 26138 13062 26262
rect 13338 26138 13462 26262
rect 13738 26138 13862 26262
rect 14138 26138 14262 26262
rect 14538 26138 14662 26262
rect 14938 26138 15062 26262
rect 15338 26138 15462 26262
rect 538 25738 662 25862
rect 938 25738 1062 25862
rect 1338 25738 1462 25862
rect 1738 25738 1862 25862
rect 2138 25738 2262 25862
rect 2538 25738 2662 25862
rect 2938 25738 3062 25862
rect 3338 25738 3462 25862
rect 3738 25738 3862 25862
rect 4138 25738 4262 25862
rect 4538 25738 4662 25862
rect 4938 25738 5062 25862
rect 5338 25738 5462 25862
rect 5738 25738 5862 25862
rect 6138 25738 6262 25862
rect 6538 25738 6662 25862
rect 6938 25738 7062 25862
rect 7338 25738 7462 25862
rect 7738 25738 7862 25862
rect 8138 25738 8262 25862
rect 8538 25738 8662 25862
rect 8938 25738 9062 25862
rect 9338 25738 9462 25862
rect 9738 25738 9862 25862
rect 10138 25738 10262 25862
rect 10538 25738 10662 25862
rect 10938 25738 11062 25862
rect 11338 25738 11462 25862
rect 11738 25738 11862 25862
rect 12138 25738 12262 25862
rect 12538 25738 12662 25862
rect 12938 25738 13062 25862
rect 13338 25738 13462 25862
rect 13738 25738 13862 25862
rect 14138 25738 14262 25862
rect 14538 25738 14662 25862
rect 14938 25738 15062 25862
rect 15338 25738 15462 25862
rect 538 23188 662 23312
rect 938 23188 1062 23312
rect 1338 23188 1462 23312
rect 1738 23188 1862 23312
rect 2138 23188 2262 23312
rect 2538 23188 2662 23312
rect 2938 23188 3062 23312
rect 3338 23188 3462 23312
rect 3738 23188 3862 23312
rect 4138 23188 4262 23312
rect 4538 23188 4662 23312
rect 4938 23188 5062 23312
rect 5338 23188 5462 23312
rect 5738 23188 5862 23312
rect 6138 23188 6262 23312
rect 6538 23188 6662 23312
rect 6938 23188 7062 23312
rect 7338 23188 7462 23312
rect 7738 23188 7862 23312
rect 8138 23188 8262 23312
rect 8538 23188 8662 23312
rect 8938 23188 9062 23312
rect 9338 23188 9462 23312
rect 9738 23188 9862 23312
rect 10138 23188 10262 23312
rect 10538 23188 10662 23312
rect 10938 23188 11062 23312
rect 11338 23188 11462 23312
rect 11738 23188 11862 23312
rect 12138 23188 12262 23312
rect 12538 23188 12662 23312
rect 12938 23188 13062 23312
rect 13338 23188 13462 23312
rect 13738 23188 13862 23312
rect 14138 23188 14262 23312
rect 14538 23188 14662 23312
rect 14938 23188 15062 23312
rect 15338 23188 15462 23312
rect 538 22788 662 22912
rect 938 22788 1062 22912
rect 1338 22788 1462 22912
rect 1738 22788 1862 22912
rect 2138 22788 2262 22912
rect 2538 22788 2662 22912
rect 2938 22788 3062 22912
rect 3338 22788 3462 22912
rect 3738 22788 3862 22912
rect 4138 22788 4262 22912
rect 4538 22788 4662 22912
rect 4938 22788 5062 22912
rect 5338 22788 5462 22912
rect 5738 22788 5862 22912
rect 6138 22788 6262 22912
rect 6538 22788 6662 22912
rect 6938 22788 7062 22912
rect 7338 22788 7462 22912
rect 7738 22788 7862 22912
rect 8138 22788 8262 22912
rect 8538 22788 8662 22912
rect 8938 22788 9062 22912
rect 9338 22788 9462 22912
rect 9738 22788 9862 22912
rect 10138 22788 10262 22912
rect 10538 22788 10662 22912
rect 10938 22788 11062 22912
rect 11338 22788 11462 22912
rect 11738 22788 11862 22912
rect 12138 22788 12262 22912
rect 12538 22788 12662 22912
rect 12938 22788 13062 22912
rect 13338 22788 13462 22912
rect 13738 22788 13862 22912
rect 14138 22788 14262 22912
rect 14538 22788 14662 22912
rect 14938 22788 15062 22912
rect 15338 22788 15462 22912
rect 538 22388 662 22512
rect 938 22388 1062 22512
rect 1338 22388 1462 22512
rect 1738 22388 1862 22512
rect 2138 22388 2262 22512
rect 2538 22388 2662 22512
rect 2938 22388 3062 22512
rect 3338 22388 3462 22512
rect 3738 22388 3862 22512
rect 4138 22388 4262 22512
rect 4538 22388 4662 22512
rect 4938 22388 5062 22512
rect 5338 22388 5462 22512
rect 5738 22388 5862 22512
rect 6138 22388 6262 22512
rect 6538 22388 6662 22512
rect 6938 22388 7062 22512
rect 7338 22388 7462 22512
rect 7738 22388 7862 22512
rect 8138 22388 8262 22512
rect 8538 22388 8662 22512
rect 8938 22388 9062 22512
rect 9338 22388 9462 22512
rect 9738 22388 9862 22512
rect 10138 22388 10262 22512
rect 10538 22388 10662 22512
rect 10938 22388 11062 22512
rect 11338 22388 11462 22512
rect 11738 22388 11862 22512
rect 12138 22388 12262 22512
rect 12538 22388 12662 22512
rect 12938 22388 13062 22512
rect 13338 22388 13462 22512
rect 13738 22388 13862 22512
rect 14138 22388 14262 22512
rect 14538 22388 14662 22512
rect 14938 22388 15062 22512
rect 15338 22388 15462 22512
rect 538 21988 662 22112
rect 938 21988 1062 22112
rect 1338 21988 1462 22112
rect 1738 21988 1862 22112
rect 2138 21988 2262 22112
rect 2538 21988 2662 22112
rect 2938 21988 3062 22112
rect 3338 21988 3462 22112
rect 3738 21988 3862 22112
rect 4138 21988 4262 22112
rect 4538 21988 4662 22112
rect 4938 21988 5062 22112
rect 5338 21988 5462 22112
rect 5738 21988 5862 22112
rect 6138 21988 6262 22112
rect 6538 21988 6662 22112
rect 6938 21988 7062 22112
rect 7338 21988 7462 22112
rect 7738 21988 7862 22112
rect 8138 21988 8262 22112
rect 8538 21988 8662 22112
rect 8938 21988 9062 22112
rect 9338 21988 9462 22112
rect 9738 21988 9862 22112
rect 10138 21988 10262 22112
rect 10538 21988 10662 22112
rect 10938 21988 11062 22112
rect 11338 21988 11462 22112
rect 11738 21988 11862 22112
rect 12138 21988 12262 22112
rect 12538 21988 12662 22112
rect 12938 21988 13062 22112
rect 13338 21988 13462 22112
rect 13738 21988 13862 22112
rect 14138 21988 14262 22112
rect 14538 21988 14662 22112
rect 14938 21988 15062 22112
rect 15338 21988 15462 22112
rect 538 21588 662 21712
rect 938 21588 1062 21712
rect 1338 21588 1462 21712
rect 1738 21588 1862 21712
rect 2138 21588 2262 21712
rect 2538 21588 2662 21712
rect 2938 21588 3062 21712
rect 3338 21588 3462 21712
rect 3738 21588 3862 21712
rect 4138 21588 4262 21712
rect 4538 21588 4662 21712
rect 4938 21588 5062 21712
rect 5338 21588 5462 21712
rect 5738 21588 5862 21712
rect 6138 21588 6262 21712
rect 6538 21588 6662 21712
rect 6938 21588 7062 21712
rect 7338 21588 7462 21712
rect 7738 21588 7862 21712
rect 8138 21588 8262 21712
rect 8538 21588 8662 21712
rect 8938 21588 9062 21712
rect 9338 21588 9462 21712
rect 9738 21588 9862 21712
rect 10138 21588 10262 21712
rect 10538 21588 10662 21712
rect 10938 21588 11062 21712
rect 11338 21588 11462 21712
rect 11738 21588 11862 21712
rect 12138 21588 12262 21712
rect 12538 21588 12662 21712
rect 12938 21588 13062 21712
rect 13338 21588 13462 21712
rect 13738 21588 13862 21712
rect 14138 21588 14262 21712
rect 14538 21588 14662 21712
rect 14938 21588 15062 21712
rect 15338 21588 15462 21712
rect 538 21188 662 21312
rect 938 21188 1062 21312
rect 1338 21188 1462 21312
rect 1738 21188 1862 21312
rect 2138 21188 2262 21312
rect 2538 21188 2662 21312
rect 2938 21188 3062 21312
rect 3338 21188 3462 21312
rect 3738 21188 3862 21312
rect 4138 21188 4262 21312
rect 4538 21188 4662 21312
rect 4938 21188 5062 21312
rect 5338 21188 5462 21312
rect 5738 21188 5862 21312
rect 6138 21188 6262 21312
rect 6538 21188 6662 21312
rect 6938 21188 7062 21312
rect 7338 21188 7462 21312
rect 7738 21188 7862 21312
rect 8138 21188 8262 21312
rect 8538 21188 8662 21312
rect 8938 21188 9062 21312
rect 9338 21188 9462 21312
rect 9738 21188 9862 21312
rect 10138 21188 10262 21312
rect 10538 21188 10662 21312
rect 10938 21188 11062 21312
rect 11338 21188 11462 21312
rect 11738 21188 11862 21312
rect 12138 21188 12262 21312
rect 12538 21188 12662 21312
rect 12938 21188 13062 21312
rect 13338 21188 13462 21312
rect 13738 21188 13862 21312
rect 14138 21188 14262 21312
rect 14538 21188 14662 21312
rect 14938 21188 15062 21312
rect 15338 21188 15462 21312
rect 538 20788 662 20912
rect 938 20788 1062 20912
rect 1338 20788 1462 20912
rect 1738 20788 1862 20912
rect 2138 20788 2262 20912
rect 2538 20788 2662 20912
rect 2938 20788 3062 20912
rect 3338 20788 3462 20912
rect 3738 20788 3862 20912
rect 4138 20788 4262 20912
rect 4538 20788 4662 20912
rect 4938 20788 5062 20912
rect 5338 20788 5462 20912
rect 5738 20788 5862 20912
rect 6138 20788 6262 20912
rect 6538 20788 6662 20912
rect 6938 20788 7062 20912
rect 7338 20788 7462 20912
rect 7738 20788 7862 20912
rect 8138 20788 8262 20912
rect 8538 20788 8662 20912
rect 8938 20788 9062 20912
rect 9338 20788 9462 20912
rect 9738 20788 9862 20912
rect 10138 20788 10262 20912
rect 10538 20788 10662 20912
rect 10938 20788 11062 20912
rect 11338 20788 11462 20912
rect 11738 20788 11862 20912
rect 12138 20788 12262 20912
rect 12538 20788 12662 20912
rect 12938 20788 13062 20912
rect 13338 20788 13462 20912
rect 13738 20788 13862 20912
rect 14138 20788 14262 20912
rect 14538 20788 14662 20912
rect 14938 20788 15062 20912
rect 15338 20788 15462 20912
rect 538 20388 662 20512
rect 938 20388 1062 20512
rect 1338 20388 1462 20512
rect 1738 20388 1862 20512
rect 2138 20388 2262 20512
rect 2538 20388 2662 20512
rect 2938 20388 3062 20512
rect 3338 20388 3462 20512
rect 3738 20388 3862 20512
rect 4138 20388 4262 20512
rect 4538 20388 4662 20512
rect 4938 20388 5062 20512
rect 5338 20388 5462 20512
rect 5738 20388 5862 20512
rect 6138 20388 6262 20512
rect 6538 20388 6662 20512
rect 6938 20388 7062 20512
rect 7338 20388 7462 20512
rect 7738 20388 7862 20512
rect 8138 20388 8262 20512
rect 8538 20388 8662 20512
rect 8938 20388 9062 20512
rect 9338 20388 9462 20512
rect 9738 20388 9862 20512
rect 10138 20388 10262 20512
rect 10538 20388 10662 20512
rect 10938 20388 11062 20512
rect 11338 20388 11462 20512
rect 11738 20388 11862 20512
rect 12138 20388 12262 20512
rect 12538 20388 12662 20512
rect 12938 20388 13062 20512
rect 13338 20388 13462 20512
rect 13738 20388 13862 20512
rect 14138 20388 14262 20512
rect 14538 20388 14662 20512
rect 14938 20388 15062 20512
rect 15338 20388 15462 20512
rect 538 19988 662 20112
rect 938 19988 1062 20112
rect 1338 19988 1462 20112
rect 1738 19988 1862 20112
rect 2138 19988 2262 20112
rect 2538 19988 2662 20112
rect 2938 19988 3062 20112
rect 3338 19988 3462 20112
rect 3738 19988 3862 20112
rect 4138 19988 4262 20112
rect 4538 19988 4662 20112
rect 4938 19988 5062 20112
rect 5338 19988 5462 20112
rect 5738 19988 5862 20112
rect 6138 19988 6262 20112
rect 6538 19988 6662 20112
rect 6938 19988 7062 20112
rect 7338 19988 7462 20112
rect 7738 19988 7862 20112
rect 8138 19988 8262 20112
rect 8538 19988 8662 20112
rect 8938 19988 9062 20112
rect 9338 19988 9462 20112
rect 9738 19988 9862 20112
rect 10138 19988 10262 20112
rect 10538 19988 10662 20112
rect 10938 19988 11062 20112
rect 11338 19988 11462 20112
rect 11738 19988 11862 20112
rect 12138 19988 12262 20112
rect 12538 19988 12662 20112
rect 12938 19988 13062 20112
rect 13338 19988 13462 20112
rect 13738 19988 13862 20112
rect 14138 19988 14262 20112
rect 14538 19988 14662 20112
rect 14938 19988 15062 20112
rect 15338 19988 15462 20112
rect 538 19588 662 19712
rect 938 19588 1062 19712
rect 1338 19588 1462 19712
rect 1738 19588 1862 19712
rect 2138 19588 2262 19712
rect 2538 19588 2662 19712
rect 2938 19588 3062 19712
rect 3338 19588 3462 19712
rect 3738 19588 3862 19712
rect 4138 19588 4262 19712
rect 4538 19588 4662 19712
rect 4938 19588 5062 19712
rect 5338 19588 5462 19712
rect 5738 19588 5862 19712
rect 6138 19588 6262 19712
rect 6538 19588 6662 19712
rect 6938 19588 7062 19712
rect 7338 19588 7462 19712
rect 7738 19588 7862 19712
rect 8138 19588 8262 19712
rect 8538 19588 8662 19712
rect 8938 19588 9062 19712
rect 9338 19588 9462 19712
rect 9738 19588 9862 19712
rect 10138 19588 10262 19712
rect 10538 19588 10662 19712
rect 10938 19588 11062 19712
rect 11338 19588 11462 19712
rect 11738 19588 11862 19712
rect 12138 19588 12262 19712
rect 12538 19588 12662 19712
rect 12938 19588 13062 19712
rect 13338 19588 13462 19712
rect 13738 19588 13862 19712
rect 14138 19588 14262 19712
rect 14538 19588 14662 19712
rect 14938 19588 15062 19712
rect 15338 19588 15462 19712
rect 538 19188 662 19312
rect 938 19188 1062 19312
rect 1338 19188 1462 19312
rect 1738 19188 1862 19312
rect 2138 19188 2262 19312
rect 2538 19188 2662 19312
rect 2938 19188 3062 19312
rect 3338 19188 3462 19312
rect 3738 19188 3862 19312
rect 4138 19188 4262 19312
rect 4538 19188 4662 19312
rect 4938 19188 5062 19312
rect 5338 19188 5462 19312
rect 5738 19188 5862 19312
rect 6138 19188 6262 19312
rect 6538 19188 6662 19312
rect 6938 19188 7062 19312
rect 7338 19188 7462 19312
rect 7738 19188 7862 19312
rect 8138 19188 8262 19312
rect 8538 19188 8662 19312
rect 8938 19188 9062 19312
rect 9338 19188 9462 19312
rect 9738 19188 9862 19312
rect 10138 19188 10262 19312
rect 10538 19188 10662 19312
rect 10938 19188 11062 19312
rect 11338 19188 11462 19312
rect 11738 19188 11862 19312
rect 12138 19188 12262 19312
rect 12538 19188 12662 19312
rect 12938 19188 13062 19312
rect 13338 19188 13462 19312
rect 13738 19188 13862 19312
rect 14138 19188 14262 19312
rect 14538 19188 14662 19312
rect 14938 19188 15062 19312
rect 15338 19188 15462 19312
rect 538 17688 662 17812
rect 938 17688 1062 17812
rect 1338 17688 1462 17812
rect 1738 17688 1862 17812
rect 2138 17688 2262 17812
rect 2538 17688 2662 17812
rect 2938 17688 3062 17812
rect 3338 17688 3462 17812
rect 3738 17688 3862 17812
rect 4138 17688 4262 17812
rect 4538 17688 4662 17812
rect 4938 17688 5062 17812
rect 5338 17688 5462 17812
rect 5738 17688 5862 17812
rect 6138 17688 6262 17812
rect 6538 17688 6662 17812
rect 6938 17688 7062 17812
rect 7338 17688 7462 17812
rect 7738 17688 7862 17812
rect 8138 17688 8262 17812
rect 8538 17688 8662 17812
rect 8938 17688 9062 17812
rect 9338 17688 9462 17812
rect 9738 17688 9862 17812
rect 10138 17688 10262 17812
rect 10538 17688 10662 17812
rect 10938 17688 11062 17812
rect 11338 17688 11462 17812
rect 11738 17688 11862 17812
rect 12138 17688 12262 17812
rect 12538 17688 12662 17812
rect 12938 17688 13062 17812
rect 13338 17688 13462 17812
rect 13738 17688 13862 17812
rect 14138 17688 14262 17812
rect 14538 17688 14662 17812
rect 14938 17688 15062 17812
rect 15338 17688 15462 17812
rect 538 17288 662 17412
rect 938 17288 1062 17412
rect 1338 17288 1462 17412
rect 1738 17288 1862 17412
rect 2138 17288 2262 17412
rect 2538 17288 2662 17412
rect 2938 17288 3062 17412
rect 3338 17288 3462 17412
rect 3738 17288 3862 17412
rect 4138 17288 4262 17412
rect 4538 17288 4662 17412
rect 4938 17288 5062 17412
rect 5338 17288 5462 17412
rect 5738 17288 5862 17412
rect 6138 17288 6262 17412
rect 6538 17288 6662 17412
rect 6938 17288 7062 17412
rect 7338 17288 7462 17412
rect 7738 17288 7862 17412
rect 8138 17288 8262 17412
rect 8538 17288 8662 17412
rect 8938 17288 9062 17412
rect 9338 17288 9462 17412
rect 9738 17288 9862 17412
rect 10138 17288 10262 17412
rect 10538 17288 10662 17412
rect 10938 17288 11062 17412
rect 11338 17288 11462 17412
rect 11738 17288 11862 17412
rect 12138 17288 12262 17412
rect 12538 17288 12662 17412
rect 12938 17288 13062 17412
rect 13338 17288 13462 17412
rect 13738 17288 13862 17412
rect 14138 17288 14262 17412
rect 14538 17288 14662 17412
rect 14938 17288 15062 17412
rect 15338 17288 15462 17412
rect 538 16888 662 17012
rect 938 16888 1062 17012
rect 1338 16888 1462 17012
rect 1738 16888 1862 17012
rect 2138 16888 2262 17012
rect 2538 16888 2662 17012
rect 2938 16888 3062 17012
rect 3338 16888 3462 17012
rect 3738 16888 3862 17012
rect 4138 16888 4262 17012
rect 4538 16888 4662 17012
rect 4938 16888 5062 17012
rect 5338 16888 5462 17012
rect 5738 16888 5862 17012
rect 6138 16888 6262 17012
rect 6538 16888 6662 17012
rect 6938 16888 7062 17012
rect 7338 16888 7462 17012
rect 7738 16888 7862 17012
rect 8138 16888 8262 17012
rect 8538 16888 8662 17012
rect 8938 16888 9062 17012
rect 9338 16888 9462 17012
rect 9738 16888 9862 17012
rect 10138 16888 10262 17012
rect 10538 16888 10662 17012
rect 10938 16888 11062 17012
rect 11338 16888 11462 17012
rect 11738 16888 11862 17012
rect 12138 16888 12262 17012
rect 12538 16888 12662 17012
rect 12938 16888 13062 17012
rect 13338 16888 13462 17012
rect 13738 16888 13862 17012
rect 14138 16888 14262 17012
rect 14538 16888 14662 17012
rect 14938 16888 15062 17012
rect 15338 16888 15462 17012
rect 538 16488 662 16612
rect 938 16488 1062 16612
rect 1338 16488 1462 16612
rect 1738 16488 1862 16612
rect 2138 16488 2262 16612
rect 2538 16488 2662 16612
rect 2938 16488 3062 16612
rect 3338 16488 3462 16612
rect 3738 16488 3862 16612
rect 4138 16488 4262 16612
rect 4538 16488 4662 16612
rect 4938 16488 5062 16612
rect 5338 16488 5462 16612
rect 5738 16488 5862 16612
rect 6138 16488 6262 16612
rect 6538 16488 6662 16612
rect 6938 16488 7062 16612
rect 7338 16488 7462 16612
rect 7738 16488 7862 16612
rect 8138 16488 8262 16612
rect 8538 16488 8662 16612
rect 8938 16488 9062 16612
rect 9338 16488 9462 16612
rect 9738 16488 9862 16612
rect 10138 16488 10262 16612
rect 10538 16488 10662 16612
rect 10938 16488 11062 16612
rect 11338 16488 11462 16612
rect 11738 16488 11862 16612
rect 12138 16488 12262 16612
rect 12538 16488 12662 16612
rect 12938 16488 13062 16612
rect 13338 16488 13462 16612
rect 13738 16488 13862 16612
rect 14138 16488 14262 16612
rect 14538 16488 14662 16612
rect 14938 16488 15062 16612
rect 15338 16488 15462 16612
rect 538 16088 662 16212
rect 938 16088 1062 16212
rect 1338 16088 1462 16212
rect 1738 16088 1862 16212
rect 2138 16088 2262 16212
rect 2538 16088 2662 16212
rect 2938 16088 3062 16212
rect 3338 16088 3462 16212
rect 3738 16088 3862 16212
rect 4138 16088 4262 16212
rect 4538 16088 4662 16212
rect 4938 16088 5062 16212
rect 5338 16088 5462 16212
rect 5738 16088 5862 16212
rect 6138 16088 6262 16212
rect 6538 16088 6662 16212
rect 6938 16088 7062 16212
rect 7338 16088 7462 16212
rect 7738 16088 7862 16212
rect 8138 16088 8262 16212
rect 8538 16088 8662 16212
rect 8938 16088 9062 16212
rect 9338 16088 9462 16212
rect 9738 16088 9862 16212
rect 10138 16088 10262 16212
rect 10538 16088 10662 16212
rect 10938 16088 11062 16212
rect 11338 16088 11462 16212
rect 11738 16088 11862 16212
rect 12138 16088 12262 16212
rect 12538 16088 12662 16212
rect 12938 16088 13062 16212
rect 13338 16088 13462 16212
rect 13738 16088 13862 16212
rect 14138 16088 14262 16212
rect 14538 16088 14662 16212
rect 14938 16088 15062 16212
rect 15338 16088 15462 16212
rect 538 15688 662 15812
rect 938 15688 1062 15812
rect 1338 15688 1462 15812
rect 1738 15688 1862 15812
rect 2138 15688 2262 15812
rect 2538 15688 2662 15812
rect 2938 15688 3062 15812
rect 3338 15688 3462 15812
rect 3738 15688 3862 15812
rect 4138 15688 4262 15812
rect 4538 15688 4662 15812
rect 4938 15688 5062 15812
rect 5338 15688 5462 15812
rect 5738 15688 5862 15812
rect 6138 15688 6262 15812
rect 6538 15688 6662 15812
rect 6938 15688 7062 15812
rect 7338 15688 7462 15812
rect 7738 15688 7862 15812
rect 8138 15688 8262 15812
rect 8538 15688 8662 15812
rect 8938 15688 9062 15812
rect 9338 15688 9462 15812
rect 9738 15688 9862 15812
rect 10138 15688 10262 15812
rect 10538 15688 10662 15812
rect 10938 15688 11062 15812
rect 11338 15688 11462 15812
rect 11738 15688 11862 15812
rect 12138 15688 12262 15812
rect 12538 15688 12662 15812
rect 12938 15688 13062 15812
rect 13338 15688 13462 15812
rect 13738 15688 13862 15812
rect 14138 15688 14262 15812
rect 14538 15688 14662 15812
rect 14938 15688 15062 15812
rect 15338 15688 15462 15812
rect 538 15288 662 15412
rect 938 15288 1062 15412
rect 1338 15288 1462 15412
rect 1738 15288 1862 15412
rect 2138 15288 2262 15412
rect 2538 15288 2662 15412
rect 2938 15288 3062 15412
rect 3338 15288 3462 15412
rect 3738 15288 3862 15412
rect 4138 15288 4262 15412
rect 4538 15288 4662 15412
rect 4938 15288 5062 15412
rect 5338 15288 5462 15412
rect 5738 15288 5862 15412
rect 6138 15288 6262 15412
rect 6538 15288 6662 15412
rect 6938 15288 7062 15412
rect 7338 15288 7462 15412
rect 7738 15288 7862 15412
rect 8138 15288 8262 15412
rect 8538 15288 8662 15412
rect 8938 15288 9062 15412
rect 9338 15288 9462 15412
rect 9738 15288 9862 15412
rect 10138 15288 10262 15412
rect 10538 15288 10662 15412
rect 10938 15288 11062 15412
rect 11338 15288 11462 15412
rect 11738 15288 11862 15412
rect 12138 15288 12262 15412
rect 12538 15288 12662 15412
rect 12938 15288 13062 15412
rect 13338 15288 13462 15412
rect 13738 15288 13862 15412
rect 14138 15288 14262 15412
rect 14538 15288 14662 15412
rect 14938 15288 15062 15412
rect 15338 15288 15462 15412
rect 538 14888 662 15012
rect 938 14888 1062 15012
rect 1338 14888 1462 15012
rect 1738 14888 1862 15012
rect 2138 14888 2262 15012
rect 2538 14888 2662 15012
rect 2938 14888 3062 15012
rect 3338 14888 3462 15012
rect 3738 14888 3862 15012
rect 4138 14888 4262 15012
rect 4538 14888 4662 15012
rect 4938 14888 5062 15012
rect 5338 14888 5462 15012
rect 5738 14888 5862 15012
rect 6138 14888 6262 15012
rect 6538 14888 6662 15012
rect 6938 14888 7062 15012
rect 7338 14888 7462 15012
rect 7738 14888 7862 15012
rect 8138 14888 8262 15012
rect 8538 14888 8662 15012
rect 8938 14888 9062 15012
rect 9338 14888 9462 15012
rect 9738 14888 9862 15012
rect 10138 14888 10262 15012
rect 10538 14888 10662 15012
rect 10938 14888 11062 15012
rect 11338 14888 11462 15012
rect 11738 14888 11862 15012
rect 12138 14888 12262 15012
rect 12538 14888 12662 15012
rect 12938 14888 13062 15012
rect 13338 14888 13462 15012
rect 13738 14888 13862 15012
rect 14138 14888 14262 15012
rect 14538 14888 14662 15012
rect 14938 14888 15062 15012
rect 15338 14888 15462 15012
rect 538 14488 662 14612
rect 938 14488 1062 14612
rect 1338 14488 1462 14612
rect 1738 14488 1862 14612
rect 2138 14488 2262 14612
rect 2538 14488 2662 14612
rect 2938 14488 3062 14612
rect 3338 14488 3462 14612
rect 3738 14488 3862 14612
rect 4138 14488 4262 14612
rect 4538 14488 4662 14612
rect 4938 14488 5062 14612
rect 5338 14488 5462 14612
rect 5738 14488 5862 14612
rect 6138 14488 6262 14612
rect 6538 14488 6662 14612
rect 6938 14488 7062 14612
rect 7338 14488 7462 14612
rect 7738 14488 7862 14612
rect 8138 14488 8262 14612
rect 8538 14488 8662 14612
rect 8938 14488 9062 14612
rect 9338 14488 9462 14612
rect 9738 14488 9862 14612
rect 10138 14488 10262 14612
rect 10538 14488 10662 14612
rect 10938 14488 11062 14612
rect 11338 14488 11462 14612
rect 11738 14488 11862 14612
rect 12138 14488 12262 14612
rect 12538 14488 12662 14612
rect 12938 14488 13062 14612
rect 13338 14488 13462 14612
rect 13738 14488 13862 14612
rect 14138 14488 14262 14612
rect 14538 14488 14662 14612
rect 14938 14488 15062 14612
rect 15338 14488 15462 14612
rect 538 14088 662 14212
rect 938 14088 1062 14212
rect 1338 14088 1462 14212
rect 1738 14088 1862 14212
rect 2138 14088 2262 14212
rect 2538 14088 2662 14212
rect 2938 14088 3062 14212
rect 3338 14088 3462 14212
rect 3738 14088 3862 14212
rect 4138 14088 4262 14212
rect 4538 14088 4662 14212
rect 4938 14088 5062 14212
rect 5338 14088 5462 14212
rect 5738 14088 5862 14212
rect 6138 14088 6262 14212
rect 6538 14088 6662 14212
rect 6938 14088 7062 14212
rect 7338 14088 7462 14212
rect 7738 14088 7862 14212
rect 8138 14088 8262 14212
rect 8538 14088 8662 14212
rect 8938 14088 9062 14212
rect 9338 14088 9462 14212
rect 9738 14088 9862 14212
rect 10138 14088 10262 14212
rect 10538 14088 10662 14212
rect 10938 14088 11062 14212
rect 11338 14088 11462 14212
rect 11738 14088 11862 14212
rect 12138 14088 12262 14212
rect 12538 14088 12662 14212
rect 12938 14088 13062 14212
rect 13338 14088 13462 14212
rect 13738 14088 13862 14212
rect 14138 14088 14262 14212
rect 14538 14088 14662 14212
rect 14938 14088 15062 14212
rect 15338 14088 15462 14212
rect 538 13688 662 13812
rect 938 13688 1062 13812
rect 1338 13688 1462 13812
rect 1738 13688 1862 13812
rect 2138 13688 2262 13812
rect 2538 13688 2662 13812
rect 2938 13688 3062 13812
rect 3338 13688 3462 13812
rect 3738 13688 3862 13812
rect 4138 13688 4262 13812
rect 4538 13688 4662 13812
rect 4938 13688 5062 13812
rect 5338 13688 5462 13812
rect 5738 13688 5862 13812
rect 6138 13688 6262 13812
rect 6538 13688 6662 13812
rect 6938 13688 7062 13812
rect 7338 13688 7462 13812
rect 7738 13688 7862 13812
rect 8138 13688 8262 13812
rect 8538 13688 8662 13812
rect 8938 13688 9062 13812
rect 9338 13688 9462 13812
rect 9738 13688 9862 13812
rect 10138 13688 10262 13812
rect 10538 13688 10662 13812
rect 10938 13688 11062 13812
rect 11338 13688 11462 13812
rect 11738 13688 11862 13812
rect 12138 13688 12262 13812
rect 12538 13688 12662 13812
rect 12938 13688 13062 13812
rect 13338 13688 13462 13812
rect 13738 13688 13862 13812
rect 14138 13688 14262 13812
rect 14538 13688 14662 13812
rect 14938 13688 15062 13812
rect 15338 13688 15462 13812
rect 538 11388 662 11512
rect 938 11388 1062 11512
rect 1338 11388 1462 11512
rect 1738 11388 1862 11512
rect 2138 11388 2262 11512
rect 2538 11388 2662 11512
rect 2938 11388 3062 11512
rect 3338 11388 3462 11512
rect 3738 11388 3862 11512
rect 4138 11388 4262 11512
rect 4538 11388 4662 11512
rect 4938 11388 5062 11512
rect 5338 11388 5462 11512
rect 5738 11388 5862 11512
rect 6138 11388 6262 11512
rect 6538 11388 6662 11512
rect 6938 11388 7062 11512
rect 7338 11388 7462 11512
rect 7738 11388 7862 11512
rect 8138 11388 8262 11512
rect 8538 11388 8662 11512
rect 8938 11388 9062 11512
rect 9338 11388 9462 11512
rect 9738 11388 9862 11512
rect 10138 11388 10262 11512
rect 10538 11388 10662 11512
rect 10938 11388 11062 11512
rect 11338 11388 11462 11512
rect 11738 11388 11862 11512
rect 12138 11388 12262 11512
rect 12538 11388 12662 11512
rect 12938 11388 13062 11512
rect 13338 11388 13462 11512
rect 13738 11388 13862 11512
rect 14138 11388 14262 11512
rect 14538 11388 14662 11512
rect 14938 11388 15062 11512
rect 15338 11388 15462 11512
rect 538 10988 662 11112
rect 938 10988 1062 11112
rect 1338 10988 1462 11112
rect 1738 10988 1862 11112
rect 2138 10988 2262 11112
rect 2538 10988 2662 11112
rect 2938 10988 3062 11112
rect 3338 10988 3462 11112
rect 3738 10988 3862 11112
rect 4138 10988 4262 11112
rect 4538 10988 4662 11112
rect 4938 10988 5062 11112
rect 5338 10988 5462 11112
rect 5738 10988 5862 11112
rect 6138 10988 6262 11112
rect 6538 10988 6662 11112
rect 6938 10988 7062 11112
rect 7338 10988 7462 11112
rect 7738 10988 7862 11112
rect 8138 10988 8262 11112
rect 8538 10988 8662 11112
rect 8938 10988 9062 11112
rect 9338 10988 9462 11112
rect 9738 10988 9862 11112
rect 10138 10988 10262 11112
rect 10538 10988 10662 11112
rect 10938 10988 11062 11112
rect 11338 10988 11462 11112
rect 11738 10988 11862 11112
rect 12138 10988 12262 11112
rect 12538 10988 12662 11112
rect 12938 10988 13062 11112
rect 13338 10988 13462 11112
rect 13738 10988 13862 11112
rect 14138 10988 14262 11112
rect 14538 10988 14662 11112
rect 14938 10988 15062 11112
rect 15338 10988 15462 11112
rect 538 10588 662 10712
rect 938 10588 1062 10712
rect 1338 10588 1462 10712
rect 1738 10588 1862 10712
rect 2138 10588 2262 10712
rect 2538 10588 2662 10712
rect 2938 10588 3062 10712
rect 3338 10588 3462 10712
rect 3738 10588 3862 10712
rect 4138 10588 4262 10712
rect 4538 10588 4662 10712
rect 4938 10588 5062 10712
rect 5338 10588 5462 10712
rect 5738 10588 5862 10712
rect 6138 10588 6262 10712
rect 6538 10588 6662 10712
rect 6938 10588 7062 10712
rect 7338 10588 7462 10712
rect 7738 10588 7862 10712
rect 8138 10588 8262 10712
rect 8538 10588 8662 10712
rect 8938 10588 9062 10712
rect 9338 10588 9462 10712
rect 9738 10588 9862 10712
rect 10138 10588 10262 10712
rect 10538 10588 10662 10712
rect 10938 10588 11062 10712
rect 11338 10588 11462 10712
rect 11738 10588 11862 10712
rect 12138 10588 12262 10712
rect 12538 10588 12662 10712
rect 12938 10588 13062 10712
rect 13338 10588 13462 10712
rect 13738 10588 13862 10712
rect 14138 10588 14262 10712
rect 14538 10588 14662 10712
rect 14938 10588 15062 10712
rect 15338 10588 15462 10712
rect 538 10188 662 10312
rect 938 10188 1062 10312
rect 1338 10188 1462 10312
rect 1738 10188 1862 10312
rect 2138 10188 2262 10312
rect 2538 10188 2662 10312
rect 2938 10188 3062 10312
rect 3338 10188 3462 10312
rect 3738 10188 3862 10312
rect 4138 10188 4262 10312
rect 4538 10188 4662 10312
rect 4938 10188 5062 10312
rect 5338 10188 5462 10312
rect 5738 10188 5862 10312
rect 6138 10188 6262 10312
rect 6538 10188 6662 10312
rect 6938 10188 7062 10312
rect 7338 10188 7462 10312
rect 7738 10188 7862 10312
rect 8138 10188 8262 10312
rect 8538 10188 8662 10312
rect 8938 10188 9062 10312
rect 9338 10188 9462 10312
rect 9738 10188 9862 10312
rect 10138 10188 10262 10312
rect 10538 10188 10662 10312
rect 10938 10188 11062 10312
rect 11338 10188 11462 10312
rect 11738 10188 11862 10312
rect 12138 10188 12262 10312
rect 12538 10188 12662 10312
rect 12938 10188 13062 10312
rect 13338 10188 13462 10312
rect 13738 10188 13862 10312
rect 14138 10188 14262 10312
rect 14538 10188 14662 10312
rect 14938 10188 15062 10312
rect 15338 10188 15462 10312
rect 538 9788 662 9912
rect 938 9788 1062 9912
rect 1338 9788 1462 9912
rect 1738 9788 1862 9912
rect 2138 9788 2262 9912
rect 2538 9788 2662 9912
rect 2938 9788 3062 9912
rect 3338 9788 3462 9912
rect 3738 9788 3862 9912
rect 4138 9788 4262 9912
rect 4538 9788 4662 9912
rect 4938 9788 5062 9912
rect 5338 9788 5462 9912
rect 5738 9788 5862 9912
rect 6138 9788 6262 9912
rect 6538 9788 6662 9912
rect 6938 9788 7062 9912
rect 7338 9788 7462 9912
rect 7738 9788 7862 9912
rect 8138 9788 8262 9912
rect 8538 9788 8662 9912
rect 8938 9788 9062 9912
rect 9338 9788 9462 9912
rect 9738 9788 9862 9912
rect 10138 9788 10262 9912
rect 10538 9788 10662 9912
rect 10938 9788 11062 9912
rect 11338 9788 11462 9912
rect 11738 9788 11862 9912
rect 12138 9788 12262 9912
rect 12538 9788 12662 9912
rect 12938 9788 13062 9912
rect 13338 9788 13462 9912
rect 13738 9788 13862 9912
rect 14138 9788 14262 9912
rect 14538 9788 14662 9912
rect 14938 9788 15062 9912
rect 15338 9788 15462 9912
rect 538 9388 662 9512
rect 938 9388 1062 9512
rect 1338 9388 1462 9512
rect 1738 9388 1862 9512
rect 2138 9388 2262 9512
rect 2538 9388 2662 9512
rect 2938 9388 3062 9512
rect 3338 9388 3462 9512
rect 3738 9388 3862 9512
rect 4138 9388 4262 9512
rect 4538 9388 4662 9512
rect 4938 9388 5062 9512
rect 5338 9388 5462 9512
rect 5738 9388 5862 9512
rect 6138 9388 6262 9512
rect 6538 9388 6662 9512
rect 6938 9388 7062 9512
rect 7338 9388 7462 9512
rect 7738 9388 7862 9512
rect 8138 9388 8262 9512
rect 8538 9388 8662 9512
rect 8938 9388 9062 9512
rect 9338 9388 9462 9512
rect 9738 9388 9862 9512
rect 10138 9388 10262 9512
rect 10538 9388 10662 9512
rect 10938 9388 11062 9512
rect 11338 9388 11462 9512
rect 11738 9388 11862 9512
rect 12138 9388 12262 9512
rect 12538 9388 12662 9512
rect 12938 9388 13062 9512
rect 13338 9388 13462 9512
rect 13738 9388 13862 9512
rect 14138 9388 14262 9512
rect 14538 9388 14662 9512
rect 14938 9388 15062 9512
rect 15338 9388 15462 9512
rect 538 8988 662 9112
rect 938 8988 1062 9112
rect 1338 8988 1462 9112
rect 1738 8988 1862 9112
rect 2138 8988 2262 9112
rect 2538 8988 2662 9112
rect 2938 8988 3062 9112
rect 3338 8988 3462 9112
rect 3738 8988 3862 9112
rect 4138 8988 4262 9112
rect 4538 8988 4662 9112
rect 4938 8988 5062 9112
rect 5338 8988 5462 9112
rect 5738 8988 5862 9112
rect 6138 8988 6262 9112
rect 6538 8988 6662 9112
rect 6938 8988 7062 9112
rect 7338 8988 7462 9112
rect 7738 8988 7862 9112
rect 8138 8988 8262 9112
rect 8538 8988 8662 9112
rect 8938 8988 9062 9112
rect 9338 8988 9462 9112
rect 9738 8988 9862 9112
rect 10138 8988 10262 9112
rect 10538 8988 10662 9112
rect 10938 8988 11062 9112
rect 11338 8988 11462 9112
rect 11738 8988 11862 9112
rect 12138 8988 12262 9112
rect 12538 8988 12662 9112
rect 12938 8988 13062 9112
rect 13338 8988 13462 9112
rect 13738 8988 13862 9112
rect 14138 8988 14262 9112
rect 14538 8988 14662 9112
rect 14938 8988 15062 9112
rect 15338 8988 15462 9112
rect 538 8588 662 8712
rect 938 8588 1062 8712
rect 1338 8588 1462 8712
rect 1738 8588 1862 8712
rect 2138 8588 2262 8712
rect 2538 8588 2662 8712
rect 2938 8588 3062 8712
rect 3338 8588 3462 8712
rect 3738 8588 3862 8712
rect 4138 8588 4262 8712
rect 4538 8588 4662 8712
rect 4938 8588 5062 8712
rect 5338 8588 5462 8712
rect 5738 8588 5862 8712
rect 6138 8588 6262 8712
rect 6538 8588 6662 8712
rect 6938 8588 7062 8712
rect 7338 8588 7462 8712
rect 7738 8588 7862 8712
rect 8138 8588 8262 8712
rect 8538 8588 8662 8712
rect 8938 8588 9062 8712
rect 9338 8588 9462 8712
rect 9738 8588 9862 8712
rect 10138 8588 10262 8712
rect 10538 8588 10662 8712
rect 10938 8588 11062 8712
rect 11338 8588 11462 8712
rect 11738 8588 11862 8712
rect 12138 8588 12262 8712
rect 12538 8588 12662 8712
rect 12938 8588 13062 8712
rect 13338 8588 13462 8712
rect 13738 8588 13862 8712
rect 14138 8588 14262 8712
rect 14538 8588 14662 8712
rect 14938 8588 15062 8712
rect 15338 8588 15462 8712
rect 538 8188 662 8312
rect 938 8188 1062 8312
rect 1338 8188 1462 8312
rect 1738 8188 1862 8312
rect 2138 8188 2262 8312
rect 2538 8188 2662 8312
rect 2938 8188 3062 8312
rect 3338 8188 3462 8312
rect 3738 8188 3862 8312
rect 4138 8188 4262 8312
rect 4538 8188 4662 8312
rect 4938 8188 5062 8312
rect 5338 8188 5462 8312
rect 5738 8188 5862 8312
rect 6138 8188 6262 8312
rect 6538 8188 6662 8312
rect 6938 8188 7062 8312
rect 7338 8188 7462 8312
rect 7738 8188 7862 8312
rect 8138 8188 8262 8312
rect 8538 8188 8662 8312
rect 8938 8188 9062 8312
rect 9338 8188 9462 8312
rect 9738 8188 9862 8312
rect 10138 8188 10262 8312
rect 10538 8188 10662 8312
rect 10938 8188 11062 8312
rect 11338 8188 11462 8312
rect 11738 8188 11862 8312
rect 12138 8188 12262 8312
rect 12538 8188 12662 8312
rect 12938 8188 13062 8312
rect 13338 8188 13462 8312
rect 13738 8188 13862 8312
rect 14138 8188 14262 8312
rect 14538 8188 14662 8312
rect 14938 8188 15062 8312
rect 15338 8188 15462 8312
rect 538 7788 662 7912
rect 938 7788 1062 7912
rect 1338 7788 1462 7912
rect 1738 7788 1862 7912
rect 2138 7788 2262 7912
rect 2538 7788 2662 7912
rect 2938 7788 3062 7912
rect 3338 7788 3462 7912
rect 3738 7788 3862 7912
rect 4138 7788 4262 7912
rect 4538 7788 4662 7912
rect 4938 7788 5062 7912
rect 5338 7788 5462 7912
rect 5738 7788 5862 7912
rect 6138 7788 6262 7912
rect 6538 7788 6662 7912
rect 6938 7788 7062 7912
rect 7338 7788 7462 7912
rect 7738 7788 7862 7912
rect 8138 7788 8262 7912
rect 8538 7788 8662 7912
rect 8938 7788 9062 7912
rect 9338 7788 9462 7912
rect 9738 7788 9862 7912
rect 10138 7788 10262 7912
rect 10538 7788 10662 7912
rect 10938 7788 11062 7912
rect 11338 7788 11462 7912
rect 11738 7788 11862 7912
rect 12138 7788 12262 7912
rect 12538 7788 12662 7912
rect 12938 7788 13062 7912
rect 13338 7788 13462 7912
rect 13738 7788 13862 7912
rect 14138 7788 14262 7912
rect 14538 7788 14662 7912
rect 14938 7788 15062 7912
rect 15338 7788 15462 7912
rect 538 7388 662 7512
rect 938 7388 1062 7512
rect 1338 7388 1462 7512
rect 1738 7388 1862 7512
rect 2138 7388 2262 7512
rect 2538 7388 2662 7512
rect 2938 7388 3062 7512
rect 3338 7388 3462 7512
rect 3738 7388 3862 7512
rect 4138 7388 4262 7512
rect 4538 7388 4662 7512
rect 4938 7388 5062 7512
rect 5338 7388 5462 7512
rect 5738 7388 5862 7512
rect 6138 7388 6262 7512
rect 6538 7388 6662 7512
rect 6938 7388 7062 7512
rect 7338 7388 7462 7512
rect 7738 7388 7862 7512
rect 8138 7388 8262 7512
rect 8538 7388 8662 7512
rect 8938 7388 9062 7512
rect 9338 7388 9462 7512
rect 9738 7388 9862 7512
rect 10138 7388 10262 7512
rect 10538 7388 10662 7512
rect 10938 7388 11062 7512
rect 11338 7388 11462 7512
rect 11738 7388 11862 7512
rect 12138 7388 12262 7512
rect 12538 7388 12662 7512
rect 12938 7388 13062 7512
rect 13338 7388 13462 7512
rect 13738 7388 13862 7512
rect 14138 7388 14262 7512
rect 14538 7388 14662 7512
rect 14938 7388 15062 7512
rect 15338 7388 15462 7512
rect 538 5888 662 6012
rect 938 5888 1062 6012
rect 1338 5888 1462 6012
rect 1738 5888 1862 6012
rect 2138 5888 2262 6012
rect 2538 5888 2662 6012
rect 2938 5888 3062 6012
rect 3338 5888 3462 6012
rect 3738 5888 3862 6012
rect 4138 5888 4262 6012
rect 4538 5888 4662 6012
rect 4938 5888 5062 6012
rect 5338 5888 5462 6012
rect 5738 5888 5862 6012
rect 6138 5888 6262 6012
rect 6538 5888 6662 6012
rect 6938 5888 7062 6012
rect 7338 5888 7462 6012
rect 7738 5888 7862 6012
rect 8138 5888 8262 6012
rect 8538 5888 8662 6012
rect 8938 5888 9062 6012
rect 9338 5888 9462 6012
rect 9738 5888 9862 6012
rect 10138 5888 10262 6012
rect 10538 5888 10662 6012
rect 10938 5888 11062 6012
rect 11338 5888 11462 6012
rect 11738 5888 11862 6012
rect 12138 5888 12262 6012
rect 12538 5888 12662 6012
rect 12938 5888 13062 6012
rect 13338 5888 13462 6012
rect 13738 5888 13862 6012
rect 14138 5888 14262 6012
rect 14538 5888 14662 6012
rect 14938 5888 15062 6012
rect 15338 5888 15462 6012
rect 538 5488 662 5612
rect 938 5488 1062 5612
rect 1338 5488 1462 5612
rect 1738 5488 1862 5612
rect 2138 5488 2262 5612
rect 2538 5488 2662 5612
rect 2938 5488 3062 5612
rect 3338 5488 3462 5612
rect 3738 5488 3862 5612
rect 4138 5488 4262 5612
rect 4538 5488 4662 5612
rect 4938 5488 5062 5612
rect 5338 5488 5462 5612
rect 5738 5488 5862 5612
rect 6138 5488 6262 5612
rect 6538 5488 6662 5612
rect 6938 5488 7062 5612
rect 7338 5488 7462 5612
rect 7738 5488 7862 5612
rect 8138 5488 8262 5612
rect 8538 5488 8662 5612
rect 8938 5488 9062 5612
rect 9338 5488 9462 5612
rect 9738 5488 9862 5612
rect 10138 5488 10262 5612
rect 10538 5488 10662 5612
rect 10938 5488 11062 5612
rect 11338 5488 11462 5612
rect 11738 5488 11862 5612
rect 12138 5488 12262 5612
rect 12538 5488 12662 5612
rect 12938 5488 13062 5612
rect 13338 5488 13462 5612
rect 13738 5488 13862 5612
rect 14138 5488 14262 5612
rect 14538 5488 14662 5612
rect 14938 5488 15062 5612
rect 15338 5488 15462 5612
rect 538 5088 662 5212
rect 938 5088 1062 5212
rect 1338 5088 1462 5212
rect 1738 5088 1862 5212
rect 2138 5088 2262 5212
rect 2538 5088 2662 5212
rect 2938 5088 3062 5212
rect 3338 5088 3462 5212
rect 3738 5088 3862 5212
rect 4138 5088 4262 5212
rect 4538 5088 4662 5212
rect 4938 5088 5062 5212
rect 5338 5088 5462 5212
rect 5738 5088 5862 5212
rect 6138 5088 6262 5212
rect 6538 5088 6662 5212
rect 6938 5088 7062 5212
rect 7338 5088 7462 5212
rect 7738 5088 7862 5212
rect 8138 5088 8262 5212
rect 8538 5088 8662 5212
rect 8938 5088 9062 5212
rect 9338 5088 9462 5212
rect 9738 5088 9862 5212
rect 10138 5088 10262 5212
rect 10538 5088 10662 5212
rect 10938 5088 11062 5212
rect 11338 5088 11462 5212
rect 11738 5088 11862 5212
rect 12138 5088 12262 5212
rect 12538 5088 12662 5212
rect 12938 5088 13062 5212
rect 13338 5088 13462 5212
rect 13738 5088 13862 5212
rect 14138 5088 14262 5212
rect 14538 5088 14662 5212
rect 14938 5088 15062 5212
rect 15338 5088 15462 5212
rect 538 4688 662 4812
rect 938 4688 1062 4812
rect 1338 4688 1462 4812
rect 1738 4688 1862 4812
rect 2138 4688 2262 4812
rect 2538 4688 2662 4812
rect 2938 4688 3062 4812
rect 3338 4688 3462 4812
rect 3738 4688 3862 4812
rect 4138 4688 4262 4812
rect 4538 4688 4662 4812
rect 4938 4688 5062 4812
rect 5338 4688 5462 4812
rect 5738 4688 5862 4812
rect 6138 4688 6262 4812
rect 6538 4688 6662 4812
rect 6938 4688 7062 4812
rect 7338 4688 7462 4812
rect 7738 4688 7862 4812
rect 8138 4688 8262 4812
rect 8538 4688 8662 4812
rect 8938 4688 9062 4812
rect 9338 4688 9462 4812
rect 9738 4688 9862 4812
rect 10138 4688 10262 4812
rect 10538 4688 10662 4812
rect 10938 4688 11062 4812
rect 11338 4688 11462 4812
rect 11738 4688 11862 4812
rect 12138 4688 12262 4812
rect 12538 4688 12662 4812
rect 12938 4688 13062 4812
rect 13338 4688 13462 4812
rect 13738 4688 13862 4812
rect 14138 4688 14262 4812
rect 14538 4688 14662 4812
rect 14938 4688 15062 4812
rect 15338 4688 15462 4812
rect 538 4288 662 4412
rect 938 4288 1062 4412
rect 1338 4288 1462 4412
rect 1738 4288 1862 4412
rect 2138 4288 2262 4412
rect 2538 4288 2662 4412
rect 2938 4288 3062 4412
rect 3338 4288 3462 4412
rect 3738 4288 3862 4412
rect 4138 4288 4262 4412
rect 4538 4288 4662 4412
rect 4938 4288 5062 4412
rect 5338 4288 5462 4412
rect 5738 4288 5862 4412
rect 6138 4288 6262 4412
rect 6538 4288 6662 4412
rect 6938 4288 7062 4412
rect 7338 4288 7462 4412
rect 7738 4288 7862 4412
rect 8138 4288 8262 4412
rect 8538 4288 8662 4412
rect 8938 4288 9062 4412
rect 9338 4288 9462 4412
rect 9738 4288 9862 4412
rect 10138 4288 10262 4412
rect 10538 4288 10662 4412
rect 10938 4288 11062 4412
rect 11338 4288 11462 4412
rect 11738 4288 11862 4412
rect 12138 4288 12262 4412
rect 12538 4288 12662 4412
rect 12938 4288 13062 4412
rect 13338 4288 13462 4412
rect 13738 4288 13862 4412
rect 14138 4288 14262 4412
rect 14538 4288 14662 4412
rect 14938 4288 15062 4412
rect 15338 4288 15462 4412
rect 538 3888 662 4012
rect 938 3888 1062 4012
rect 1338 3888 1462 4012
rect 1738 3888 1862 4012
rect 2138 3888 2262 4012
rect 2538 3888 2662 4012
rect 2938 3888 3062 4012
rect 3338 3888 3462 4012
rect 3738 3888 3862 4012
rect 4138 3888 4262 4012
rect 4538 3888 4662 4012
rect 4938 3888 5062 4012
rect 5338 3888 5462 4012
rect 5738 3888 5862 4012
rect 6138 3888 6262 4012
rect 6538 3888 6662 4012
rect 6938 3888 7062 4012
rect 7338 3888 7462 4012
rect 7738 3888 7862 4012
rect 8138 3888 8262 4012
rect 8538 3888 8662 4012
rect 8938 3888 9062 4012
rect 9338 3888 9462 4012
rect 9738 3888 9862 4012
rect 10138 3888 10262 4012
rect 10538 3888 10662 4012
rect 10938 3888 11062 4012
rect 11338 3888 11462 4012
rect 11738 3888 11862 4012
rect 12138 3888 12262 4012
rect 12538 3888 12662 4012
rect 12938 3888 13062 4012
rect 13338 3888 13462 4012
rect 13738 3888 13862 4012
rect 14138 3888 14262 4012
rect 14538 3888 14662 4012
rect 14938 3888 15062 4012
rect 15338 3888 15462 4012
rect 538 3488 662 3612
rect 938 3488 1062 3612
rect 1338 3488 1462 3612
rect 1738 3488 1862 3612
rect 2138 3488 2262 3612
rect 2538 3488 2662 3612
rect 2938 3488 3062 3612
rect 3338 3488 3462 3612
rect 3738 3488 3862 3612
rect 4138 3488 4262 3612
rect 4538 3488 4662 3612
rect 4938 3488 5062 3612
rect 5338 3488 5462 3612
rect 5738 3488 5862 3612
rect 6138 3488 6262 3612
rect 6538 3488 6662 3612
rect 6938 3488 7062 3612
rect 7338 3488 7462 3612
rect 7738 3488 7862 3612
rect 8138 3488 8262 3612
rect 8538 3488 8662 3612
rect 8938 3488 9062 3612
rect 9338 3488 9462 3612
rect 9738 3488 9862 3612
rect 10138 3488 10262 3612
rect 10538 3488 10662 3612
rect 10938 3488 11062 3612
rect 11338 3488 11462 3612
rect 11738 3488 11862 3612
rect 12138 3488 12262 3612
rect 12538 3488 12662 3612
rect 12938 3488 13062 3612
rect 13338 3488 13462 3612
rect 13738 3488 13862 3612
rect 14138 3488 14262 3612
rect 14538 3488 14662 3612
rect 14938 3488 15062 3612
rect 15338 3488 15462 3612
rect 538 3088 662 3212
rect 938 3088 1062 3212
rect 1338 3088 1462 3212
rect 1738 3088 1862 3212
rect 2138 3088 2262 3212
rect 2538 3088 2662 3212
rect 2938 3088 3062 3212
rect 3338 3088 3462 3212
rect 3738 3088 3862 3212
rect 4138 3088 4262 3212
rect 4538 3088 4662 3212
rect 4938 3088 5062 3212
rect 5338 3088 5462 3212
rect 5738 3088 5862 3212
rect 6138 3088 6262 3212
rect 6538 3088 6662 3212
rect 6938 3088 7062 3212
rect 7338 3088 7462 3212
rect 7738 3088 7862 3212
rect 8138 3088 8262 3212
rect 8538 3088 8662 3212
rect 8938 3088 9062 3212
rect 9338 3088 9462 3212
rect 9738 3088 9862 3212
rect 10138 3088 10262 3212
rect 10538 3088 10662 3212
rect 10938 3088 11062 3212
rect 11338 3088 11462 3212
rect 11738 3088 11862 3212
rect 12138 3088 12262 3212
rect 12538 3088 12662 3212
rect 12938 3088 13062 3212
rect 13338 3088 13462 3212
rect 13738 3088 13862 3212
rect 14138 3088 14262 3212
rect 14538 3088 14662 3212
rect 14938 3088 15062 3212
rect 15338 3088 15462 3212
rect 538 2688 662 2812
rect 938 2688 1062 2812
rect 1338 2688 1462 2812
rect 1738 2688 1862 2812
rect 2138 2688 2262 2812
rect 2538 2688 2662 2812
rect 2938 2688 3062 2812
rect 3338 2688 3462 2812
rect 3738 2688 3862 2812
rect 4138 2688 4262 2812
rect 4538 2688 4662 2812
rect 4938 2688 5062 2812
rect 5338 2688 5462 2812
rect 5738 2688 5862 2812
rect 6138 2688 6262 2812
rect 6538 2688 6662 2812
rect 6938 2688 7062 2812
rect 7338 2688 7462 2812
rect 7738 2688 7862 2812
rect 8138 2688 8262 2812
rect 8538 2688 8662 2812
rect 8938 2688 9062 2812
rect 9338 2688 9462 2812
rect 9738 2688 9862 2812
rect 10138 2688 10262 2812
rect 10538 2688 10662 2812
rect 10938 2688 11062 2812
rect 11338 2688 11462 2812
rect 11738 2688 11862 2812
rect 12138 2688 12262 2812
rect 12538 2688 12662 2812
rect 12938 2688 13062 2812
rect 13338 2688 13462 2812
rect 13738 2688 13862 2812
rect 14138 2688 14262 2812
rect 14538 2688 14662 2812
rect 14938 2688 15062 2812
rect 15338 2688 15462 2812
rect 538 2288 662 2412
rect 938 2288 1062 2412
rect 1338 2288 1462 2412
rect 1738 2288 1862 2412
rect 2138 2288 2262 2412
rect 2538 2288 2662 2412
rect 2938 2288 3062 2412
rect 3338 2288 3462 2412
rect 3738 2288 3862 2412
rect 4138 2288 4262 2412
rect 4538 2288 4662 2412
rect 4938 2288 5062 2412
rect 5338 2288 5462 2412
rect 5738 2288 5862 2412
rect 6138 2288 6262 2412
rect 6538 2288 6662 2412
rect 6938 2288 7062 2412
rect 7338 2288 7462 2412
rect 7738 2288 7862 2412
rect 8138 2288 8262 2412
rect 8538 2288 8662 2412
rect 8938 2288 9062 2412
rect 9338 2288 9462 2412
rect 9738 2288 9862 2412
rect 10138 2288 10262 2412
rect 10538 2288 10662 2412
rect 10938 2288 11062 2412
rect 11338 2288 11462 2412
rect 11738 2288 11862 2412
rect 12138 2288 12262 2412
rect 12538 2288 12662 2412
rect 12938 2288 13062 2412
rect 13338 2288 13462 2412
rect 13738 2288 13862 2412
rect 14138 2288 14262 2412
rect 14538 2288 14662 2412
rect 14938 2288 15062 2412
rect 15338 2288 15462 2412
rect 538 1888 662 2012
rect 938 1888 1062 2012
rect 1338 1888 1462 2012
rect 1738 1888 1862 2012
rect 2138 1888 2262 2012
rect 2538 1888 2662 2012
rect 2938 1888 3062 2012
rect 3338 1888 3462 2012
rect 3738 1888 3862 2012
rect 4138 1888 4262 2012
rect 4538 1888 4662 2012
rect 4938 1888 5062 2012
rect 5338 1888 5462 2012
rect 5738 1888 5862 2012
rect 6138 1888 6262 2012
rect 6538 1888 6662 2012
rect 6938 1888 7062 2012
rect 7338 1888 7462 2012
rect 7738 1888 7862 2012
rect 8138 1888 8262 2012
rect 8538 1888 8662 2012
rect 8938 1888 9062 2012
rect 9338 1888 9462 2012
rect 9738 1888 9862 2012
rect 10138 1888 10262 2012
rect 10538 1888 10662 2012
rect 10938 1888 11062 2012
rect 11338 1888 11462 2012
rect 11738 1888 11862 2012
rect 12138 1888 12262 2012
rect 12538 1888 12662 2012
rect 12938 1888 13062 2012
rect 13338 1888 13462 2012
rect 13738 1888 13862 2012
rect 14138 1888 14262 2012
rect 14538 1888 14662 2012
rect 14938 1888 15062 2012
rect 15338 1888 15462 2012
rect 1138 238 1262 362
rect 1538 238 1662 362
rect 1938 238 2062 362
rect 2338 238 2462 362
rect 2738 238 2862 362
rect 3138 238 3262 362
rect 3538 238 3662 362
rect 3938 238 4062 362
rect 4338 238 4462 362
rect 4738 238 4862 362
rect 5138 238 5262 362
rect 5538 238 5662 362
rect 5938 238 6062 362
rect 6338 238 6462 362
rect 6738 238 6862 362
rect 7138 238 7262 362
rect 7538 238 7662 362
rect 7938 238 8062 362
rect 8338 238 8462 362
rect 8738 238 8862 362
rect 9138 238 9262 362
rect 9538 238 9662 362
rect 9938 238 10062 362
rect 10338 238 10462 362
rect 10738 238 10862 362
rect 11138 238 11262 362
rect 11538 238 11662 362
rect 11938 238 12062 362
rect 12338 238 12462 362
rect 12738 238 12862 362
rect 13138 238 13262 362
rect 13538 238 13662 362
rect 13938 238 14062 362
rect 14338 238 14462 362
rect 14738 238 14862 362
<< metal6 >>
rect 0 35062 16000 35600
rect 0 34938 538 35062
rect 662 34938 938 35062
rect 1062 34938 1338 35062
rect 1462 34938 1738 35062
rect 1862 34938 2138 35062
rect 2262 34938 2538 35062
rect 2662 34938 2938 35062
rect 3062 34938 3338 35062
rect 3462 34938 3738 35062
rect 3862 34938 4138 35062
rect 4262 34938 4538 35062
rect 4662 34938 4938 35062
rect 5062 34938 5338 35062
rect 5462 34938 5738 35062
rect 5862 34938 6138 35062
rect 6262 34938 6538 35062
rect 6662 34938 6938 35062
rect 7062 34938 7338 35062
rect 7462 34938 7738 35062
rect 7862 34938 8138 35062
rect 8262 34938 8538 35062
rect 8662 34938 8938 35062
rect 9062 34938 9338 35062
rect 9462 34938 9738 35062
rect 9862 34938 10138 35062
rect 10262 34938 10538 35062
rect 10662 34938 10938 35062
rect 11062 34938 11338 35062
rect 11462 34938 11738 35062
rect 11862 34938 12138 35062
rect 12262 34938 12538 35062
rect 12662 34938 12938 35062
rect 13062 34938 13338 35062
rect 13462 34938 13738 35062
rect 13862 34938 14138 35062
rect 14262 34938 14538 35062
rect 14662 34938 14938 35062
rect 15062 34938 15338 35062
rect 15462 34938 16000 35062
rect 0 34662 16000 34938
rect 0 34538 538 34662
rect 662 34538 938 34662
rect 1062 34538 1338 34662
rect 1462 34538 1738 34662
rect 1862 34538 2138 34662
rect 2262 34538 2538 34662
rect 2662 34538 2938 34662
rect 3062 34538 3338 34662
rect 3462 34538 3738 34662
rect 3862 34538 4138 34662
rect 4262 34538 4538 34662
rect 4662 34538 4938 34662
rect 5062 34538 5338 34662
rect 5462 34538 5738 34662
rect 5862 34538 6138 34662
rect 6262 34538 6538 34662
rect 6662 34538 6938 34662
rect 7062 34538 7338 34662
rect 7462 34538 7738 34662
rect 7862 34538 8138 34662
rect 8262 34538 8538 34662
rect 8662 34538 8938 34662
rect 9062 34538 9338 34662
rect 9462 34538 9738 34662
rect 9862 34538 10138 34662
rect 10262 34538 10538 34662
rect 10662 34538 10938 34662
rect 11062 34538 11338 34662
rect 11462 34538 11738 34662
rect 11862 34538 12138 34662
rect 12262 34538 12538 34662
rect 12662 34538 12938 34662
rect 13062 34538 13338 34662
rect 13462 34538 13738 34662
rect 13862 34538 14138 34662
rect 14262 34538 14538 34662
rect 14662 34538 14938 34662
rect 15062 34538 15338 34662
rect 15462 34538 16000 34662
rect 0 34262 16000 34538
rect 0 34138 538 34262
rect 662 34138 938 34262
rect 1062 34138 1338 34262
rect 1462 34138 1738 34262
rect 1862 34138 2138 34262
rect 2262 34138 2538 34262
rect 2662 34138 2938 34262
rect 3062 34138 3338 34262
rect 3462 34138 3738 34262
rect 3862 34138 4138 34262
rect 4262 34138 4538 34262
rect 4662 34138 4938 34262
rect 5062 34138 5338 34262
rect 5462 34138 5738 34262
rect 5862 34138 6138 34262
rect 6262 34138 6538 34262
rect 6662 34138 6938 34262
rect 7062 34138 7338 34262
rect 7462 34138 7738 34262
rect 7862 34138 8138 34262
rect 8262 34138 8538 34262
rect 8662 34138 8938 34262
rect 9062 34138 9338 34262
rect 9462 34138 9738 34262
rect 9862 34138 10138 34262
rect 10262 34138 10538 34262
rect 10662 34138 10938 34262
rect 11062 34138 11338 34262
rect 11462 34138 11738 34262
rect 11862 34138 12138 34262
rect 12262 34138 12538 34262
rect 12662 34138 12938 34262
rect 13062 34138 13338 34262
rect 13462 34138 13738 34262
rect 13862 34138 14138 34262
rect 14262 34138 14538 34262
rect 14662 34138 14938 34262
rect 15062 34138 15338 34262
rect 15462 34138 16000 34262
rect 0 33862 16000 34138
rect 0 33738 538 33862
rect 662 33738 938 33862
rect 1062 33738 1338 33862
rect 1462 33738 1738 33862
rect 1862 33738 2138 33862
rect 2262 33738 2538 33862
rect 2662 33738 2938 33862
rect 3062 33738 3338 33862
rect 3462 33738 3738 33862
rect 3862 33738 4138 33862
rect 4262 33738 4538 33862
rect 4662 33738 4938 33862
rect 5062 33738 5338 33862
rect 5462 33738 5738 33862
rect 5862 33738 6138 33862
rect 6262 33738 6538 33862
rect 6662 33738 6938 33862
rect 7062 33738 7338 33862
rect 7462 33738 7738 33862
rect 7862 33738 8138 33862
rect 8262 33738 8538 33862
rect 8662 33738 8938 33862
rect 9062 33738 9338 33862
rect 9462 33738 9738 33862
rect 9862 33738 10138 33862
rect 10262 33738 10538 33862
rect 10662 33738 10938 33862
rect 11062 33738 11338 33862
rect 11462 33738 11738 33862
rect 11862 33738 12138 33862
rect 12262 33738 12538 33862
rect 12662 33738 12938 33862
rect 13062 33738 13338 33862
rect 13462 33738 13738 33862
rect 13862 33738 14138 33862
rect 14262 33738 14538 33862
rect 14662 33738 14938 33862
rect 15062 33738 15338 33862
rect 15462 33738 16000 33862
rect 0 33462 16000 33738
rect 0 33338 538 33462
rect 662 33338 938 33462
rect 1062 33338 1338 33462
rect 1462 33338 1738 33462
rect 1862 33338 2138 33462
rect 2262 33338 2538 33462
rect 2662 33338 2938 33462
rect 3062 33338 3338 33462
rect 3462 33338 3738 33462
rect 3862 33338 4138 33462
rect 4262 33338 4538 33462
rect 4662 33338 4938 33462
rect 5062 33338 5338 33462
rect 5462 33338 5738 33462
rect 5862 33338 6138 33462
rect 6262 33338 6538 33462
rect 6662 33338 6938 33462
rect 7062 33338 7338 33462
rect 7462 33338 7738 33462
rect 7862 33338 8138 33462
rect 8262 33338 8538 33462
rect 8662 33338 8938 33462
rect 9062 33338 9338 33462
rect 9462 33338 9738 33462
rect 9862 33338 10138 33462
rect 10262 33338 10538 33462
rect 10662 33338 10938 33462
rect 11062 33338 11338 33462
rect 11462 33338 11738 33462
rect 11862 33338 12138 33462
rect 12262 33338 12538 33462
rect 12662 33338 12938 33462
rect 13062 33338 13338 33462
rect 13462 33338 13738 33462
rect 13862 33338 14138 33462
rect 14262 33338 14538 33462
rect 14662 33338 14938 33462
rect 15062 33338 15338 33462
rect 15462 33338 16000 33462
rect 0 33062 16000 33338
rect 0 32938 538 33062
rect 662 32938 938 33062
rect 1062 32938 1338 33062
rect 1462 32938 1738 33062
rect 1862 32938 2138 33062
rect 2262 32938 2538 33062
rect 2662 32938 2938 33062
rect 3062 32938 3338 33062
rect 3462 32938 3738 33062
rect 3862 32938 4138 33062
rect 4262 32938 4538 33062
rect 4662 32938 4938 33062
rect 5062 32938 5338 33062
rect 5462 32938 5738 33062
rect 5862 32938 6138 33062
rect 6262 32938 6538 33062
rect 6662 32938 6938 33062
rect 7062 32938 7338 33062
rect 7462 32938 7738 33062
rect 7862 32938 8138 33062
rect 8262 32938 8538 33062
rect 8662 32938 8938 33062
rect 9062 32938 9338 33062
rect 9462 32938 9738 33062
rect 9862 32938 10138 33062
rect 10262 32938 10538 33062
rect 10662 32938 10938 33062
rect 11062 32938 11338 33062
rect 11462 32938 11738 33062
rect 11862 32938 12138 33062
rect 12262 32938 12538 33062
rect 12662 32938 12938 33062
rect 13062 32938 13338 33062
rect 13462 32938 13738 33062
rect 13862 32938 14138 33062
rect 14262 32938 14538 33062
rect 14662 32938 14938 33062
rect 15062 32938 15338 33062
rect 15462 32938 16000 33062
rect 0 32662 16000 32938
rect 0 32538 538 32662
rect 662 32538 938 32662
rect 1062 32538 1338 32662
rect 1462 32538 1738 32662
rect 1862 32538 2138 32662
rect 2262 32538 2538 32662
rect 2662 32538 2938 32662
rect 3062 32538 3338 32662
rect 3462 32538 3738 32662
rect 3862 32538 4138 32662
rect 4262 32538 4538 32662
rect 4662 32538 4938 32662
rect 5062 32538 5338 32662
rect 5462 32538 5738 32662
rect 5862 32538 6138 32662
rect 6262 32538 6538 32662
rect 6662 32538 6938 32662
rect 7062 32538 7338 32662
rect 7462 32538 7738 32662
rect 7862 32538 8138 32662
rect 8262 32538 8538 32662
rect 8662 32538 8938 32662
rect 9062 32538 9338 32662
rect 9462 32538 9738 32662
rect 9862 32538 10138 32662
rect 10262 32538 10538 32662
rect 10662 32538 10938 32662
rect 11062 32538 11338 32662
rect 11462 32538 11738 32662
rect 11862 32538 12138 32662
rect 12262 32538 12538 32662
rect 12662 32538 12938 32662
rect 13062 32538 13338 32662
rect 13462 32538 13738 32662
rect 13862 32538 14138 32662
rect 14262 32538 14538 32662
rect 14662 32538 14938 32662
rect 15062 32538 15338 32662
rect 15462 32538 16000 32662
rect 0 32000 16000 32538
rect 0 31062 16000 31600
rect 0 30938 538 31062
rect 662 30938 938 31062
rect 1062 30938 1338 31062
rect 1462 30938 1738 31062
rect 1862 30938 2138 31062
rect 2262 30938 2538 31062
rect 2662 30938 2938 31062
rect 3062 30938 3338 31062
rect 3462 30938 3738 31062
rect 3862 30938 4138 31062
rect 4262 30938 4538 31062
rect 4662 30938 4938 31062
rect 5062 30938 5338 31062
rect 5462 30938 5738 31062
rect 5862 30938 6138 31062
rect 6262 30938 6538 31062
rect 6662 30938 6938 31062
rect 7062 30938 7338 31062
rect 7462 30938 7738 31062
rect 7862 30938 8138 31062
rect 8262 30938 8538 31062
rect 8662 30938 8938 31062
rect 9062 30938 9338 31062
rect 9462 30938 9738 31062
rect 9862 30938 10138 31062
rect 10262 30938 10538 31062
rect 10662 30938 10938 31062
rect 11062 30938 11338 31062
rect 11462 30938 11738 31062
rect 11862 30938 12138 31062
rect 12262 30938 12538 31062
rect 12662 30938 12938 31062
rect 13062 30938 13338 31062
rect 13462 30938 13738 31062
rect 13862 30938 14138 31062
rect 14262 30938 14538 31062
rect 14662 30938 14938 31062
rect 15062 30938 15338 31062
rect 15462 30938 16000 31062
rect 0 30662 16000 30938
rect 0 30538 538 30662
rect 662 30538 938 30662
rect 1062 30538 1338 30662
rect 1462 30538 1738 30662
rect 1862 30538 2138 30662
rect 2262 30538 2538 30662
rect 2662 30538 2938 30662
rect 3062 30538 3338 30662
rect 3462 30538 3738 30662
rect 3862 30538 4138 30662
rect 4262 30538 4538 30662
rect 4662 30538 4938 30662
rect 5062 30538 5338 30662
rect 5462 30538 5738 30662
rect 5862 30538 6138 30662
rect 6262 30538 6538 30662
rect 6662 30538 6938 30662
rect 7062 30538 7338 30662
rect 7462 30538 7738 30662
rect 7862 30538 8138 30662
rect 8262 30538 8538 30662
rect 8662 30538 8938 30662
rect 9062 30538 9338 30662
rect 9462 30538 9738 30662
rect 9862 30538 10138 30662
rect 10262 30538 10538 30662
rect 10662 30538 10938 30662
rect 11062 30538 11338 30662
rect 11462 30538 11738 30662
rect 11862 30538 12138 30662
rect 12262 30538 12538 30662
rect 12662 30538 12938 30662
rect 13062 30538 13338 30662
rect 13462 30538 13738 30662
rect 13862 30538 14138 30662
rect 14262 30538 14538 30662
rect 14662 30538 14938 30662
rect 15062 30538 15338 30662
rect 15462 30538 16000 30662
rect 0 30262 16000 30538
rect 0 30138 538 30262
rect 662 30138 938 30262
rect 1062 30138 1338 30262
rect 1462 30138 1738 30262
rect 1862 30138 2138 30262
rect 2262 30138 2538 30262
rect 2662 30138 2938 30262
rect 3062 30138 3338 30262
rect 3462 30138 3738 30262
rect 3862 30138 4138 30262
rect 4262 30138 4538 30262
rect 4662 30138 4938 30262
rect 5062 30138 5338 30262
rect 5462 30138 5738 30262
rect 5862 30138 6138 30262
rect 6262 30138 6538 30262
rect 6662 30138 6938 30262
rect 7062 30138 7338 30262
rect 7462 30138 7738 30262
rect 7862 30138 8138 30262
rect 8262 30138 8538 30262
rect 8662 30138 8938 30262
rect 9062 30138 9338 30262
rect 9462 30138 9738 30262
rect 9862 30138 10138 30262
rect 10262 30138 10538 30262
rect 10662 30138 10938 30262
rect 11062 30138 11338 30262
rect 11462 30138 11738 30262
rect 11862 30138 12138 30262
rect 12262 30138 12538 30262
rect 12662 30138 12938 30262
rect 13062 30138 13338 30262
rect 13462 30138 13738 30262
rect 13862 30138 14138 30262
rect 14262 30138 14538 30262
rect 14662 30138 14938 30262
rect 15062 30138 15338 30262
rect 15462 30138 16000 30262
rect 0 29862 16000 30138
rect 0 29738 538 29862
rect 662 29738 938 29862
rect 1062 29738 1338 29862
rect 1462 29738 1738 29862
rect 1862 29738 2138 29862
rect 2262 29738 2538 29862
rect 2662 29738 2938 29862
rect 3062 29738 3338 29862
rect 3462 29738 3738 29862
rect 3862 29738 4138 29862
rect 4262 29738 4538 29862
rect 4662 29738 4938 29862
rect 5062 29738 5338 29862
rect 5462 29738 5738 29862
rect 5862 29738 6138 29862
rect 6262 29738 6538 29862
rect 6662 29738 6938 29862
rect 7062 29738 7338 29862
rect 7462 29738 7738 29862
rect 7862 29738 8138 29862
rect 8262 29738 8538 29862
rect 8662 29738 8938 29862
rect 9062 29738 9338 29862
rect 9462 29738 9738 29862
rect 9862 29738 10138 29862
rect 10262 29738 10538 29862
rect 10662 29738 10938 29862
rect 11062 29738 11338 29862
rect 11462 29738 11738 29862
rect 11862 29738 12138 29862
rect 12262 29738 12538 29862
rect 12662 29738 12938 29862
rect 13062 29738 13338 29862
rect 13462 29738 13738 29862
rect 13862 29738 14138 29862
rect 14262 29738 14538 29862
rect 14662 29738 14938 29862
rect 15062 29738 15338 29862
rect 15462 29738 16000 29862
rect 0 29462 16000 29738
rect 0 29338 538 29462
rect 662 29338 938 29462
rect 1062 29338 1338 29462
rect 1462 29338 1738 29462
rect 1862 29338 2138 29462
rect 2262 29338 2538 29462
rect 2662 29338 2938 29462
rect 3062 29338 3338 29462
rect 3462 29338 3738 29462
rect 3862 29338 4138 29462
rect 4262 29338 4538 29462
rect 4662 29338 4938 29462
rect 5062 29338 5338 29462
rect 5462 29338 5738 29462
rect 5862 29338 6138 29462
rect 6262 29338 6538 29462
rect 6662 29338 6938 29462
rect 7062 29338 7338 29462
rect 7462 29338 7738 29462
rect 7862 29338 8138 29462
rect 8262 29338 8538 29462
rect 8662 29338 8938 29462
rect 9062 29338 9338 29462
rect 9462 29338 9738 29462
rect 9862 29338 10138 29462
rect 10262 29338 10538 29462
rect 10662 29338 10938 29462
rect 11062 29338 11338 29462
rect 11462 29338 11738 29462
rect 11862 29338 12138 29462
rect 12262 29338 12538 29462
rect 12662 29338 12938 29462
rect 13062 29338 13338 29462
rect 13462 29338 13738 29462
rect 13862 29338 14138 29462
rect 14262 29338 14538 29462
rect 14662 29338 14938 29462
rect 15062 29338 15338 29462
rect 15462 29338 16000 29462
rect 0 29062 16000 29338
rect 0 28938 538 29062
rect 662 28938 938 29062
rect 1062 28938 1338 29062
rect 1462 28938 1738 29062
rect 1862 28938 2138 29062
rect 2262 28938 2538 29062
rect 2662 28938 2938 29062
rect 3062 28938 3338 29062
rect 3462 28938 3738 29062
rect 3862 28938 4138 29062
rect 4262 28938 4538 29062
rect 4662 28938 4938 29062
rect 5062 28938 5338 29062
rect 5462 28938 5738 29062
rect 5862 28938 6138 29062
rect 6262 28938 6538 29062
rect 6662 28938 6938 29062
rect 7062 28938 7338 29062
rect 7462 28938 7738 29062
rect 7862 28938 8138 29062
rect 8262 28938 8538 29062
rect 8662 28938 8938 29062
rect 9062 28938 9338 29062
rect 9462 28938 9738 29062
rect 9862 28938 10138 29062
rect 10262 28938 10538 29062
rect 10662 28938 10938 29062
rect 11062 28938 11338 29062
rect 11462 28938 11738 29062
rect 11862 28938 12138 29062
rect 12262 28938 12538 29062
rect 12662 28938 12938 29062
rect 13062 28938 13338 29062
rect 13462 28938 13738 29062
rect 13862 28938 14138 29062
rect 14262 28938 14538 29062
rect 14662 28938 14938 29062
rect 15062 28938 15338 29062
rect 15462 28938 16000 29062
rect 0 28662 16000 28938
rect 0 28538 538 28662
rect 662 28538 938 28662
rect 1062 28538 1338 28662
rect 1462 28538 1738 28662
rect 1862 28538 2138 28662
rect 2262 28538 2538 28662
rect 2662 28538 2938 28662
rect 3062 28538 3338 28662
rect 3462 28538 3738 28662
rect 3862 28538 4138 28662
rect 4262 28538 4538 28662
rect 4662 28538 4938 28662
rect 5062 28538 5338 28662
rect 5462 28538 5738 28662
rect 5862 28538 6138 28662
rect 6262 28538 6538 28662
rect 6662 28538 6938 28662
rect 7062 28538 7338 28662
rect 7462 28538 7738 28662
rect 7862 28538 8138 28662
rect 8262 28538 8538 28662
rect 8662 28538 8938 28662
rect 9062 28538 9338 28662
rect 9462 28538 9738 28662
rect 9862 28538 10138 28662
rect 10262 28538 10538 28662
rect 10662 28538 10938 28662
rect 11062 28538 11338 28662
rect 11462 28538 11738 28662
rect 11862 28538 12138 28662
rect 12262 28538 12538 28662
rect 12662 28538 12938 28662
rect 13062 28538 13338 28662
rect 13462 28538 13738 28662
rect 13862 28538 14138 28662
rect 14262 28538 14538 28662
rect 14662 28538 14938 28662
rect 15062 28538 15338 28662
rect 15462 28538 16000 28662
rect 0 28000 16000 28538
rect 0 26262 16000 26800
rect 0 26190 538 26262
rect 662 26190 938 26262
rect 1062 26190 1338 26262
rect 1462 26190 1738 26262
rect 1862 26190 2138 26262
rect 2262 26190 2538 26262
rect 2662 26190 2938 26262
rect 3062 26190 3338 26262
rect 3462 26190 3738 26262
rect 3862 26190 4138 26262
rect 4262 26190 4538 26262
rect 4662 26190 4938 26262
rect 5062 26190 5338 26262
rect 5462 26190 5738 26262
rect 5862 26190 6138 26262
rect 6262 26190 6538 26262
rect 6662 26190 6938 26262
rect 7062 26190 7338 26262
rect 7462 26190 7738 26262
rect 7862 26190 8138 26262
rect 8262 26190 8538 26262
rect 8662 26190 8938 26262
rect 9062 26190 9338 26262
rect 9462 26190 9738 26262
rect 9862 26190 10138 26262
rect 10262 26190 10538 26262
rect 10662 26190 10938 26262
rect 11062 26190 11338 26262
rect 11462 26190 11738 26262
rect 11862 26190 12138 26262
rect 12262 26190 12538 26262
rect 12662 26190 12938 26262
rect 13062 26190 13338 26262
rect 13462 26190 13738 26262
rect 13862 26190 14138 26262
rect 14262 26190 14538 26262
rect 14662 26190 14938 26262
rect 15062 26190 15338 26262
rect 15462 26190 16000 26262
rect 0 25810 410 26190
rect 790 25810 810 26190
rect 1190 25810 1210 26190
rect 1590 25810 1610 26190
rect 1990 25810 2010 26190
rect 2390 25810 2410 26190
rect 2790 25810 2810 26190
rect 3190 25810 3210 26190
rect 3590 25810 3610 26190
rect 3990 25810 4010 26190
rect 4390 25810 4410 26190
rect 4790 25810 4810 26190
rect 5190 25810 5210 26190
rect 5590 25810 5610 26190
rect 5990 25810 6010 26190
rect 6390 25810 6410 26190
rect 6790 25810 6810 26190
rect 7190 25810 7210 26190
rect 7590 25810 7610 26190
rect 7990 25810 8010 26190
rect 8390 25810 8410 26190
rect 8790 25810 8810 26190
rect 9190 25810 9210 26190
rect 9590 25810 9610 26190
rect 9990 25810 10010 26190
rect 10390 25810 10410 26190
rect 10790 25810 10810 26190
rect 11190 25810 11210 26190
rect 11590 25810 11610 26190
rect 11990 25810 12010 26190
rect 12390 25810 12410 26190
rect 12790 25810 12810 26190
rect 13190 25810 13210 26190
rect 13590 25810 13610 26190
rect 13990 25810 14010 26190
rect 14390 25810 14410 26190
rect 14790 25810 14810 26190
rect 15190 25810 15210 26190
rect 15590 25810 16000 26190
rect 0 25738 538 25810
rect 662 25738 938 25810
rect 1062 25738 1338 25810
rect 1462 25738 1738 25810
rect 1862 25738 2138 25810
rect 2262 25738 2538 25810
rect 2662 25738 2938 25810
rect 3062 25738 3338 25810
rect 3462 25738 3738 25810
rect 3862 25738 4138 25810
rect 4262 25738 4538 25810
rect 4662 25738 4938 25810
rect 5062 25738 5338 25810
rect 5462 25738 5738 25810
rect 5862 25738 6138 25810
rect 6262 25738 6538 25810
rect 6662 25738 6938 25810
rect 7062 25738 7338 25810
rect 7462 25738 7738 25810
rect 7862 25738 8138 25810
rect 8262 25738 8538 25810
rect 8662 25738 8938 25810
rect 9062 25738 9338 25810
rect 9462 25738 9738 25810
rect 9862 25738 10138 25810
rect 10262 25738 10538 25810
rect 10662 25738 10938 25810
rect 11062 25738 11338 25810
rect 11462 25738 11738 25810
rect 11862 25738 12138 25810
rect 12262 25738 12538 25810
rect 12662 25738 12938 25810
rect 13062 25738 13338 25810
rect 13462 25738 13738 25810
rect 13862 25738 14138 25810
rect 14262 25738 14538 25810
rect 14662 25738 14938 25810
rect 15062 25738 15338 25810
rect 15462 25738 16000 25810
rect 0 25200 16000 25738
rect 0 23312 16000 23800
rect 0 23240 538 23312
rect 662 23240 938 23312
rect 1062 23240 1338 23312
rect 1462 23240 1738 23312
rect 1862 23240 2138 23312
rect 2262 23240 2538 23312
rect 2662 23240 2938 23312
rect 3062 23240 3338 23312
rect 3462 23240 3738 23312
rect 3862 23240 4138 23312
rect 4262 23240 4538 23312
rect 4662 23240 4938 23312
rect 5062 23240 5338 23312
rect 5462 23240 5738 23312
rect 5862 23240 6138 23312
rect 6262 23240 6538 23312
rect 6662 23240 6938 23312
rect 7062 23240 7338 23312
rect 7462 23240 7738 23312
rect 7862 23240 8138 23312
rect 8262 23240 8538 23312
rect 8662 23240 8938 23312
rect 9062 23240 9338 23312
rect 9462 23240 9738 23312
rect 9862 23240 10138 23312
rect 10262 23240 10538 23312
rect 10662 23240 10938 23312
rect 11062 23240 11338 23312
rect 11462 23240 11738 23312
rect 11862 23240 12138 23312
rect 12262 23240 12538 23312
rect 12662 23240 12938 23312
rect 13062 23240 13338 23312
rect 13462 23240 13738 23312
rect 13862 23240 14138 23312
rect 14262 23240 14538 23312
rect 14662 23240 14938 23312
rect 15062 23240 15338 23312
rect 15462 23240 16000 23312
rect 0 22860 410 23240
rect 790 22860 810 23240
rect 1190 22860 1210 23240
rect 1590 22860 1610 23240
rect 1990 22860 2010 23240
rect 2390 22860 2410 23240
rect 2790 22860 2810 23240
rect 3190 22860 3210 23240
rect 3590 22860 3610 23240
rect 3990 22860 4010 23240
rect 4390 22860 4410 23240
rect 4790 22860 4810 23240
rect 5190 22860 5210 23240
rect 5590 22860 5610 23240
rect 5990 22860 6010 23240
rect 6390 22860 6410 23240
rect 6790 22860 6810 23240
rect 7190 22860 7210 23240
rect 7590 22860 7610 23240
rect 7990 22860 8010 23240
rect 8390 22860 8410 23240
rect 8790 22860 8810 23240
rect 9190 22860 9210 23240
rect 9590 22860 9610 23240
rect 9990 22860 10010 23240
rect 10390 22860 10410 23240
rect 10790 22860 10810 23240
rect 11190 22860 11210 23240
rect 11590 22860 11610 23240
rect 11990 22860 12010 23240
rect 12390 22860 12410 23240
rect 12790 22860 12810 23240
rect 13190 22860 13210 23240
rect 13590 22860 13610 23240
rect 13990 22860 14010 23240
rect 14390 22860 14410 23240
rect 14790 22860 14810 23240
rect 15190 22860 15210 23240
rect 15590 22860 16000 23240
rect 0 22840 538 22860
rect 662 22840 938 22860
rect 1062 22840 1338 22860
rect 1462 22840 1738 22860
rect 1862 22840 2138 22860
rect 2262 22840 2538 22860
rect 2662 22840 2938 22860
rect 3062 22840 3338 22860
rect 3462 22840 3738 22860
rect 3862 22840 4138 22860
rect 4262 22840 4538 22860
rect 4662 22840 4938 22860
rect 5062 22840 5338 22860
rect 5462 22840 5738 22860
rect 5862 22840 6138 22860
rect 6262 22840 6538 22860
rect 6662 22840 6938 22860
rect 7062 22840 7338 22860
rect 7462 22840 7738 22860
rect 7862 22840 8138 22860
rect 8262 22840 8538 22860
rect 8662 22840 8938 22860
rect 9062 22840 9338 22860
rect 9462 22840 9738 22860
rect 9862 22840 10138 22860
rect 10262 22840 10538 22860
rect 10662 22840 10938 22860
rect 11062 22840 11338 22860
rect 11462 22840 11738 22860
rect 11862 22840 12138 22860
rect 12262 22840 12538 22860
rect 12662 22840 12938 22860
rect 13062 22840 13338 22860
rect 13462 22840 13738 22860
rect 13862 22840 14138 22860
rect 14262 22840 14538 22860
rect 14662 22840 14938 22860
rect 15062 22840 15338 22860
rect 15462 22840 16000 22860
rect 0 22460 410 22840
rect 790 22460 810 22840
rect 1190 22460 1210 22840
rect 1590 22460 1610 22840
rect 1990 22460 2010 22840
rect 2390 22460 2410 22840
rect 2790 22460 2810 22840
rect 3190 22460 3210 22840
rect 3590 22460 3610 22840
rect 3990 22460 4010 22840
rect 4390 22460 4410 22840
rect 4790 22460 4810 22840
rect 5190 22460 5210 22840
rect 5590 22460 5610 22840
rect 5990 22460 6010 22840
rect 6390 22460 6410 22840
rect 6790 22460 6810 22840
rect 7190 22460 7210 22840
rect 7590 22460 7610 22840
rect 7990 22460 8010 22840
rect 8390 22460 8410 22840
rect 8790 22460 8810 22840
rect 9190 22460 9210 22840
rect 9590 22460 9610 22840
rect 9990 22460 10010 22840
rect 10390 22460 10410 22840
rect 10790 22460 10810 22840
rect 11190 22460 11210 22840
rect 11590 22460 11610 22840
rect 11990 22460 12010 22840
rect 12390 22460 12410 22840
rect 12790 22460 12810 22840
rect 13190 22460 13210 22840
rect 13590 22460 13610 22840
rect 13990 22460 14010 22840
rect 14390 22460 14410 22840
rect 14790 22460 14810 22840
rect 15190 22460 15210 22840
rect 15590 22460 16000 22840
rect 0 22440 538 22460
rect 662 22440 938 22460
rect 1062 22440 1338 22460
rect 1462 22440 1738 22460
rect 1862 22440 2138 22460
rect 2262 22440 2538 22460
rect 2662 22440 2938 22460
rect 3062 22440 3338 22460
rect 3462 22440 3738 22460
rect 3862 22440 4138 22460
rect 4262 22440 4538 22460
rect 4662 22440 4938 22460
rect 5062 22440 5338 22460
rect 5462 22440 5738 22460
rect 5862 22440 6138 22460
rect 6262 22440 6538 22460
rect 6662 22440 6938 22460
rect 7062 22440 7338 22460
rect 7462 22440 7738 22460
rect 7862 22440 8138 22460
rect 8262 22440 8538 22460
rect 8662 22440 8938 22460
rect 9062 22440 9338 22460
rect 9462 22440 9738 22460
rect 9862 22440 10138 22460
rect 10262 22440 10538 22460
rect 10662 22440 10938 22460
rect 11062 22440 11338 22460
rect 11462 22440 11738 22460
rect 11862 22440 12138 22460
rect 12262 22440 12538 22460
rect 12662 22440 12938 22460
rect 13062 22440 13338 22460
rect 13462 22440 13738 22460
rect 13862 22440 14138 22460
rect 14262 22440 14538 22460
rect 14662 22440 14938 22460
rect 15062 22440 15338 22460
rect 15462 22440 16000 22460
rect 0 22060 410 22440
rect 790 22060 810 22440
rect 1190 22060 1210 22440
rect 1590 22060 1610 22440
rect 1990 22060 2010 22440
rect 2390 22060 2410 22440
rect 2790 22060 2810 22440
rect 3190 22060 3210 22440
rect 3590 22060 3610 22440
rect 3990 22060 4010 22440
rect 4390 22060 4410 22440
rect 4790 22060 4810 22440
rect 5190 22060 5210 22440
rect 5590 22060 5610 22440
rect 5990 22060 6010 22440
rect 6390 22060 6410 22440
rect 6790 22060 6810 22440
rect 7190 22060 7210 22440
rect 7590 22060 7610 22440
rect 7990 22060 8010 22440
rect 8390 22060 8410 22440
rect 8790 22060 8810 22440
rect 9190 22060 9210 22440
rect 9590 22060 9610 22440
rect 9990 22060 10010 22440
rect 10390 22060 10410 22440
rect 10790 22060 10810 22440
rect 11190 22060 11210 22440
rect 11590 22060 11610 22440
rect 11990 22060 12010 22440
rect 12390 22060 12410 22440
rect 12790 22060 12810 22440
rect 13190 22060 13210 22440
rect 13590 22060 13610 22440
rect 13990 22060 14010 22440
rect 14390 22060 14410 22440
rect 14790 22060 14810 22440
rect 15190 22060 15210 22440
rect 15590 22060 16000 22440
rect 0 22040 538 22060
rect 662 22040 938 22060
rect 1062 22040 1338 22060
rect 1462 22040 1738 22060
rect 1862 22040 2138 22060
rect 2262 22040 2538 22060
rect 2662 22040 2938 22060
rect 3062 22040 3338 22060
rect 3462 22040 3738 22060
rect 3862 22040 4138 22060
rect 4262 22040 4538 22060
rect 4662 22040 4938 22060
rect 5062 22040 5338 22060
rect 5462 22040 5738 22060
rect 5862 22040 6138 22060
rect 6262 22040 6538 22060
rect 6662 22040 6938 22060
rect 7062 22040 7338 22060
rect 7462 22040 7738 22060
rect 7862 22040 8138 22060
rect 8262 22040 8538 22060
rect 8662 22040 8938 22060
rect 9062 22040 9338 22060
rect 9462 22040 9738 22060
rect 9862 22040 10138 22060
rect 10262 22040 10538 22060
rect 10662 22040 10938 22060
rect 11062 22040 11338 22060
rect 11462 22040 11738 22060
rect 11862 22040 12138 22060
rect 12262 22040 12538 22060
rect 12662 22040 12938 22060
rect 13062 22040 13338 22060
rect 13462 22040 13738 22060
rect 13862 22040 14138 22060
rect 14262 22040 14538 22060
rect 14662 22040 14938 22060
rect 15062 22040 15338 22060
rect 15462 22040 16000 22060
rect 0 21660 410 22040
rect 790 21660 810 22040
rect 1190 21660 1210 22040
rect 1590 21660 1610 22040
rect 1990 21660 2010 22040
rect 2390 21660 2410 22040
rect 2790 21660 2810 22040
rect 3190 21660 3210 22040
rect 3590 21660 3610 22040
rect 3990 21660 4010 22040
rect 4390 21660 4410 22040
rect 4790 21660 4810 22040
rect 5190 21660 5210 22040
rect 5590 21660 5610 22040
rect 5990 21660 6010 22040
rect 6390 21660 6410 22040
rect 6790 21660 6810 22040
rect 7190 21660 7210 22040
rect 7590 21660 7610 22040
rect 7990 21660 8010 22040
rect 8390 21660 8410 22040
rect 8790 21660 8810 22040
rect 9190 21660 9210 22040
rect 9590 21660 9610 22040
rect 9990 21660 10010 22040
rect 10390 21660 10410 22040
rect 10790 21660 10810 22040
rect 11190 21660 11210 22040
rect 11590 21660 11610 22040
rect 11990 21660 12010 22040
rect 12390 21660 12410 22040
rect 12790 21660 12810 22040
rect 13190 21660 13210 22040
rect 13590 21660 13610 22040
rect 13990 21660 14010 22040
rect 14390 21660 14410 22040
rect 14790 21660 14810 22040
rect 15190 21660 15210 22040
rect 15590 21660 16000 22040
rect 0 21640 538 21660
rect 662 21640 938 21660
rect 1062 21640 1338 21660
rect 1462 21640 1738 21660
rect 1862 21640 2138 21660
rect 2262 21640 2538 21660
rect 2662 21640 2938 21660
rect 3062 21640 3338 21660
rect 3462 21640 3738 21660
rect 3862 21640 4138 21660
rect 4262 21640 4538 21660
rect 4662 21640 4938 21660
rect 5062 21640 5338 21660
rect 5462 21640 5738 21660
rect 5862 21640 6138 21660
rect 6262 21640 6538 21660
rect 6662 21640 6938 21660
rect 7062 21640 7338 21660
rect 7462 21640 7738 21660
rect 7862 21640 8138 21660
rect 8262 21640 8538 21660
rect 8662 21640 8938 21660
rect 9062 21640 9338 21660
rect 9462 21640 9738 21660
rect 9862 21640 10138 21660
rect 10262 21640 10538 21660
rect 10662 21640 10938 21660
rect 11062 21640 11338 21660
rect 11462 21640 11738 21660
rect 11862 21640 12138 21660
rect 12262 21640 12538 21660
rect 12662 21640 12938 21660
rect 13062 21640 13338 21660
rect 13462 21640 13738 21660
rect 13862 21640 14138 21660
rect 14262 21640 14538 21660
rect 14662 21640 14938 21660
rect 15062 21640 15338 21660
rect 15462 21640 16000 21660
rect 0 21260 410 21640
rect 790 21260 810 21640
rect 1190 21260 1210 21640
rect 1590 21260 1610 21640
rect 1990 21260 2010 21640
rect 2390 21260 2410 21640
rect 2790 21260 2810 21640
rect 3190 21260 3210 21640
rect 3590 21260 3610 21640
rect 3990 21260 4010 21640
rect 4390 21260 4410 21640
rect 4790 21260 4810 21640
rect 5190 21260 5210 21640
rect 5590 21260 5610 21640
rect 5990 21260 6010 21640
rect 6390 21260 6410 21640
rect 6790 21260 6810 21640
rect 7190 21260 7210 21640
rect 7590 21260 7610 21640
rect 7990 21260 8010 21640
rect 8390 21260 8410 21640
rect 8790 21260 8810 21640
rect 9190 21260 9210 21640
rect 9590 21260 9610 21640
rect 9990 21260 10010 21640
rect 10390 21260 10410 21640
rect 10790 21260 10810 21640
rect 11190 21260 11210 21640
rect 11590 21260 11610 21640
rect 11990 21260 12010 21640
rect 12390 21260 12410 21640
rect 12790 21260 12810 21640
rect 13190 21260 13210 21640
rect 13590 21260 13610 21640
rect 13990 21260 14010 21640
rect 14390 21260 14410 21640
rect 14790 21260 14810 21640
rect 15190 21260 15210 21640
rect 15590 21260 16000 21640
rect 0 21240 538 21260
rect 662 21240 938 21260
rect 1062 21240 1338 21260
rect 1462 21240 1738 21260
rect 1862 21240 2138 21260
rect 2262 21240 2538 21260
rect 2662 21240 2938 21260
rect 3062 21240 3338 21260
rect 3462 21240 3738 21260
rect 3862 21240 4138 21260
rect 4262 21240 4538 21260
rect 4662 21240 4938 21260
rect 5062 21240 5338 21260
rect 5462 21240 5738 21260
rect 5862 21240 6138 21260
rect 6262 21240 6538 21260
rect 6662 21240 6938 21260
rect 7062 21240 7338 21260
rect 7462 21240 7738 21260
rect 7862 21240 8138 21260
rect 8262 21240 8538 21260
rect 8662 21240 8938 21260
rect 9062 21240 9338 21260
rect 9462 21240 9738 21260
rect 9862 21240 10138 21260
rect 10262 21240 10538 21260
rect 10662 21240 10938 21260
rect 11062 21240 11338 21260
rect 11462 21240 11738 21260
rect 11862 21240 12138 21260
rect 12262 21240 12538 21260
rect 12662 21240 12938 21260
rect 13062 21240 13338 21260
rect 13462 21240 13738 21260
rect 13862 21240 14138 21260
rect 14262 21240 14538 21260
rect 14662 21240 14938 21260
rect 15062 21240 15338 21260
rect 15462 21240 16000 21260
rect 0 20860 410 21240
rect 790 20860 810 21240
rect 1190 20860 1210 21240
rect 1590 20860 1610 21240
rect 1990 20860 2010 21240
rect 2390 20860 2410 21240
rect 2790 20860 2810 21240
rect 3190 20860 3210 21240
rect 3590 20860 3610 21240
rect 3990 20860 4010 21240
rect 4390 20860 4410 21240
rect 4790 20860 4810 21240
rect 5190 20860 5210 21240
rect 5590 20860 5610 21240
rect 5990 20860 6010 21240
rect 6390 20860 6410 21240
rect 6790 20860 6810 21240
rect 7190 20860 7210 21240
rect 7590 20860 7610 21240
rect 7990 20860 8010 21240
rect 8390 20860 8410 21240
rect 8790 20860 8810 21240
rect 9190 20860 9210 21240
rect 9590 20860 9610 21240
rect 9990 20860 10010 21240
rect 10390 20860 10410 21240
rect 10790 20860 10810 21240
rect 11190 20860 11210 21240
rect 11590 20860 11610 21240
rect 11990 20860 12010 21240
rect 12390 20860 12410 21240
rect 12790 20860 12810 21240
rect 13190 20860 13210 21240
rect 13590 20860 13610 21240
rect 13990 20860 14010 21240
rect 14390 20860 14410 21240
rect 14790 20860 14810 21240
rect 15190 20860 15210 21240
rect 15590 20860 16000 21240
rect 0 20840 538 20860
rect 662 20840 938 20860
rect 1062 20840 1338 20860
rect 1462 20840 1738 20860
rect 1862 20840 2138 20860
rect 2262 20840 2538 20860
rect 2662 20840 2938 20860
rect 3062 20840 3338 20860
rect 3462 20840 3738 20860
rect 3862 20840 4138 20860
rect 4262 20840 4538 20860
rect 4662 20840 4938 20860
rect 5062 20840 5338 20860
rect 5462 20840 5738 20860
rect 5862 20840 6138 20860
rect 6262 20840 6538 20860
rect 6662 20840 6938 20860
rect 7062 20840 7338 20860
rect 7462 20840 7738 20860
rect 7862 20840 8138 20860
rect 8262 20840 8538 20860
rect 8662 20840 8938 20860
rect 9062 20840 9338 20860
rect 9462 20840 9738 20860
rect 9862 20840 10138 20860
rect 10262 20840 10538 20860
rect 10662 20840 10938 20860
rect 11062 20840 11338 20860
rect 11462 20840 11738 20860
rect 11862 20840 12138 20860
rect 12262 20840 12538 20860
rect 12662 20840 12938 20860
rect 13062 20840 13338 20860
rect 13462 20840 13738 20860
rect 13862 20840 14138 20860
rect 14262 20840 14538 20860
rect 14662 20840 14938 20860
rect 15062 20840 15338 20860
rect 15462 20840 16000 20860
rect 0 20460 410 20840
rect 790 20460 810 20840
rect 1190 20460 1210 20840
rect 1590 20460 1610 20840
rect 1990 20460 2010 20840
rect 2390 20460 2410 20840
rect 2790 20460 2810 20840
rect 3190 20460 3210 20840
rect 3590 20460 3610 20840
rect 3990 20460 4010 20840
rect 4390 20460 4410 20840
rect 4790 20460 4810 20840
rect 5190 20460 5210 20840
rect 5590 20460 5610 20840
rect 5990 20460 6010 20840
rect 6390 20460 6410 20840
rect 6790 20460 6810 20840
rect 7190 20460 7210 20840
rect 7590 20460 7610 20840
rect 7990 20460 8010 20840
rect 8390 20460 8410 20840
rect 8790 20460 8810 20840
rect 9190 20460 9210 20840
rect 9590 20460 9610 20840
rect 9990 20460 10010 20840
rect 10390 20460 10410 20840
rect 10790 20460 10810 20840
rect 11190 20460 11210 20840
rect 11590 20460 11610 20840
rect 11990 20460 12010 20840
rect 12390 20460 12410 20840
rect 12790 20460 12810 20840
rect 13190 20460 13210 20840
rect 13590 20460 13610 20840
rect 13990 20460 14010 20840
rect 14390 20460 14410 20840
rect 14790 20460 14810 20840
rect 15190 20460 15210 20840
rect 15590 20460 16000 20840
rect 0 20440 538 20460
rect 662 20440 938 20460
rect 1062 20440 1338 20460
rect 1462 20440 1738 20460
rect 1862 20440 2138 20460
rect 2262 20440 2538 20460
rect 2662 20440 2938 20460
rect 3062 20440 3338 20460
rect 3462 20440 3738 20460
rect 3862 20440 4138 20460
rect 4262 20440 4538 20460
rect 4662 20440 4938 20460
rect 5062 20440 5338 20460
rect 5462 20440 5738 20460
rect 5862 20440 6138 20460
rect 6262 20440 6538 20460
rect 6662 20440 6938 20460
rect 7062 20440 7338 20460
rect 7462 20440 7738 20460
rect 7862 20440 8138 20460
rect 8262 20440 8538 20460
rect 8662 20440 8938 20460
rect 9062 20440 9338 20460
rect 9462 20440 9738 20460
rect 9862 20440 10138 20460
rect 10262 20440 10538 20460
rect 10662 20440 10938 20460
rect 11062 20440 11338 20460
rect 11462 20440 11738 20460
rect 11862 20440 12138 20460
rect 12262 20440 12538 20460
rect 12662 20440 12938 20460
rect 13062 20440 13338 20460
rect 13462 20440 13738 20460
rect 13862 20440 14138 20460
rect 14262 20440 14538 20460
rect 14662 20440 14938 20460
rect 15062 20440 15338 20460
rect 15462 20440 16000 20460
rect 0 20060 410 20440
rect 790 20060 810 20440
rect 1190 20060 1210 20440
rect 1590 20060 1610 20440
rect 1990 20060 2010 20440
rect 2390 20060 2410 20440
rect 2790 20060 2810 20440
rect 3190 20060 3210 20440
rect 3590 20060 3610 20440
rect 3990 20060 4010 20440
rect 4390 20060 4410 20440
rect 4790 20060 4810 20440
rect 5190 20060 5210 20440
rect 5590 20060 5610 20440
rect 5990 20060 6010 20440
rect 6390 20060 6410 20440
rect 6790 20060 6810 20440
rect 7190 20060 7210 20440
rect 7590 20060 7610 20440
rect 7990 20060 8010 20440
rect 8390 20060 8410 20440
rect 8790 20060 8810 20440
rect 9190 20060 9210 20440
rect 9590 20060 9610 20440
rect 9990 20060 10010 20440
rect 10390 20060 10410 20440
rect 10790 20060 10810 20440
rect 11190 20060 11210 20440
rect 11590 20060 11610 20440
rect 11990 20060 12010 20440
rect 12390 20060 12410 20440
rect 12790 20060 12810 20440
rect 13190 20060 13210 20440
rect 13590 20060 13610 20440
rect 13990 20060 14010 20440
rect 14390 20060 14410 20440
rect 14790 20060 14810 20440
rect 15190 20060 15210 20440
rect 15590 20060 16000 20440
rect 0 20040 538 20060
rect 662 20040 938 20060
rect 1062 20040 1338 20060
rect 1462 20040 1738 20060
rect 1862 20040 2138 20060
rect 2262 20040 2538 20060
rect 2662 20040 2938 20060
rect 3062 20040 3338 20060
rect 3462 20040 3738 20060
rect 3862 20040 4138 20060
rect 4262 20040 4538 20060
rect 4662 20040 4938 20060
rect 5062 20040 5338 20060
rect 5462 20040 5738 20060
rect 5862 20040 6138 20060
rect 6262 20040 6538 20060
rect 6662 20040 6938 20060
rect 7062 20040 7338 20060
rect 7462 20040 7738 20060
rect 7862 20040 8138 20060
rect 8262 20040 8538 20060
rect 8662 20040 8938 20060
rect 9062 20040 9338 20060
rect 9462 20040 9738 20060
rect 9862 20040 10138 20060
rect 10262 20040 10538 20060
rect 10662 20040 10938 20060
rect 11062 20040 11338 20060
rect 11462 20040 11738 20060
rect 11862 20040 12138 20060
rect 12262 20040 12538 20060
rect 12662 20040 12938 20060
rect 13062 20040 13338 20060
rect 13462 20040 13738 20060
rect 13862 20040 14138 20060
rect 14262 20040 14538 20060
rect 14662 20040 14938 20060
rect 15062 20040 15338 20060
rect 15462 20040 16000 20060
rect 0 19660 410 20040
rect 790 19660 810 20040
rect 1190 19660 1210 20040
rect 1590 19660 1610 20040
rect 1990 19660 2010 20040
rect 2390 19660 2410 20040
rect 2790 19660 2810 20040
rect 3190 19660 3210 20040
rect 3590 19660 3610 20040
rect 3990 19660 4010 20040
rect 4390 19660 4410 20040
rect 4790 19660 4810 20040
rect 5190 19660 5210 20040
rect 5590 19660 5610 20040
rect 5990 19660 6010 20040
rect 6390 19660 6410 20040
rect 6790 19660 6810 20040
rect 7190 19660 7210 20040
rect 7590 19660 7610 20040
rect 7990 19660 8010 20040
rect 8390 19660 8410 20040
rect 8790 19660 8810 20040
rect 9190 19660 9210 20040
rect 9590 19660 9610 20040
rect 9990 19660 10010 20040
rect 10390 19660 10410 20040
rect 10790 19660 10810 20040
rect 11190 19660 11210 20040
rect 11590 19660 11610 20040
rect 11990 19660 12010 20040
rect 12390 19660 12410 20040
rect 12790 19660 12810 20040
rect 13190 19660 13210 20040
rect 13590 19660 13610 20040
rect 13990 19660 14010 20040
rect 14390 19660 14410 20040
rect 14790 19660 14810 20040
rect 15190 19660 15210 20040
rect 15590 19660 16000 20040
rect 0 19640 538 19660
rect 662 19640 938 19660
rect 1062 19640 1338 19660
rect 1462 19640 1738 19660
rect 1862 19640 2138 19660
rect 2262 19640 2538 19660
rect 2662 19640 2938 19660
rect 3062 19640 3338 19660
rect 3462 19640 3738 19660
rect 3862 19640 4138 19660
rect 4262 19640 4538 19660
rect 4662 19640 4938 19660
rect 5062 19640 5338 19660
rect 5462 19640 5738 19660
rect 5862 19640 6138 19660
rect 6262 19640 6538 19660
rect 6662 19640 6938 19660
rect 7062 19640 7338 19660
rect 7462 19640 7738 19660
rect 7862 19640 8138 19660
rect 8262 19640 8538 19660
rect 8662 19640 8938 19660
rect 9062 19640 9338 19660
rect 9462 19640 9738 19660
rect 9862 19640 10138 19660
rect 10262 19640 10538 19660
rect 10662 19640 10938 19660
rect 11062 19640 11338 19660
rect 11462 19640 11738 19660
rect 11862 19640 12138 19660
rect 12262 19640 12538 19660
rect 12662 19640 12938 19660
rect 13062 19640 13338 19660
rect 13462 19640 13738 19660
rect 13862 19640 14138 19660
rect 14262 19640 14538 19660
rect 14662 19640 14938 19660
rect 15062 19640 15338 19660
rect 15462 19640 16000 19660
rect 0 19260 410 19640
rect 790 19260 810 19640
rect 1190 19260 1210 19640
rect 1590 19260 1610 19640
rect 1990 19260 2010 19640
rect 2390 19260 2410 19640
rect 2790 19260 2810 19640
rect 3190 19260 3210 19640
rect 3590 19260 3610 19640
rect 3990 19260 4010 19640
rect 4390 19260 4410 19640
rect 4790 19260 4810 19640
rect 5190 19260 5210 19640
rect 5590 19260 5610 19640
rect 5990 19260 6010 19640
rect 6390 19260 6410 19640
rect 6790 19260 6810 19640
rect 7190 19260 7210 19640
rect 7590 19260 7610 19640
rect 7990 19260 8010 19640
rect 8390 19260 8410 19640
rect 8790 19260 8810 19640
rect 9190 19260 9210 19640
rect 9590 19260 9610 19640
rect 9990 19260 10010 19640
rect 10390 19260 10410 19640
rect 10790 19260 10810 19640
rect 11190 19260 11210 19640
rect 11590 19260 11610 19640
rect 11990 19260 12010 19640
rect 12390 19260 12410 19640
rect 12790 19260 12810 19640
rect 13190 19260 13210 19640
rect 13590 19260 13610 19640
rect 13990 19260 14010 19640
rect 14390 19260 14410 19640
rect 14790 19260 14810 19640
rect 15190 19260 15210 19640
rect 15590 19260 16000 19640
rect 0 19188 538 19260
rect 662 19188 938 19260
rect 1062 19188 1338 19260
rect 1462 19188 1738 19260
rect 1862 19188 2138 19260
rect 2262 19188 2538 19260
rect 2662 19188 2938 19260
rect 3062 19188 3338 19260
rect 3462 19188 3738 19260
rect 3862 19188 4138 19260
rect 4262 19188 4538 19260
rect 4662 19188 4938 19260
rect 5062 19188 5338 19260
rect 5462 19188 5738 19260
rect 5862 19188 6138 19260
rect 6262 19188 6538 19260
rect 6662 19188 6938 19260
rect 7062 19188 7338 19260
rect 7462 19188 7738 19260
rect 7862 19188 8138 19260
rect 8262 19188 8538 19260
rect 8662 19188 8938 19260
rect 9062 19188 9338 19260
rect 9462 19188 9738 19260
rect 9862 19188 10138 19260
rect 10262 19188 10538 19260
rect 10662 19188 10938 19260
rect 11062 19188 11338 19260
rect 11462 19188 11738 19260
rect 11862 19188 12138 19260
rect 12262 19188 12538 19260
rect 12662 19188 12938 19260
rect 13062 19188 13338 19260
rect 13462 19188 13738 19260
rect 13862 19188 14138 19260
rect 14262 19188 14538 19260
rect 14662 19188 14938 19260
rect 15062 19188 15338 19260
rect 15462 19188 16000 19260
rect 0 18700 16000 19188
rect 0 17812 16000 18300
rect 0 17740 538 17812
rect 662 17740 938 17812
rect 1062 17740 1338 17812
rect 1462 17740 1738 17812
rect 1862 17740 2138 17812
rect 2262 17740 2538 17812
rect 2662 17740 2938 17812
rect 3062 17740 3338 17812
rect 3462 17740 3738 17812
rect 3862 17740 4138 17812
rect 4262 17740 4538 17812
rect 4662 17740 4938 17812
rect 5062 17740 5338 17812
rect 5462 17740 5738 17812
rect 5862 17740 6138 17812
rect 6262 17740 6538 17812
rect 6662 17740 6938 17812
rect 7062 17740 7338 17812
rect 7462 17740 7738 17812
rect 7862 17740 8138 17812
rect 8262 17740 8538 17812
rect 8662 17740 8938 17812
rect 9062 17740 9338 17812
rect 9462 17740 9738 17812
rect 9862 17740 10138 17812
rect 10262 17740 10538 17812
rect 10662 17740 10938 17812
rect 11062 17740 11338 17812
rect 11462 17740 11738 17812
rect 11862 17740 12138 17812
rect 12262 17740 12538 17812
rect 12662 17740 12938 17812
rect 13062 17740 13338 17812
rect 13462 17740 13738 17812
rect 13862 17740 14138 17812
rect 14262 17740 14538 17812
rect 14662 17740 14938 17812
rect 15062 17740 15338 17812
rect 15462 17740 16000 17812
rect 0 17360 410 17740
rect 790 17360 810 17740
rect 1190 17360 1210 17740
rect 1590 17360 1610 17740
rect 1990 17360 2010 17740
rect 2390 17360 2410 17740
rect 2790 17360 2810 17740
rect 3190 17360 3210 17740
rect 3590 17360 3610 17740
rect 3990 17360 4010 17740
rect 4390 17360 4410 17740
rect 4790 17360 4810 17740
rect 5190 17360 5210 17740
rect 5590 17360 5610 17740
rect 5990 17360 6010 17740
rect 6390 17360 6410 17740
rect 6790 17360 6810 17740
rect 7190 17360 7210 17740
rect 7590 17360 7610 17740
rect 7990 17360 8010 17740
rect 8390 17360 8410 17740
rect 8790 17360 8810 17740
rect 9190 17360 9210 17740
rect 9590 17360 9610 17740
rect 9990 17360 10010 17740
rect 10390 17360 10410 17740
rect 10790 17360 10810 17740
rect 11190 17360 11210 17740
rect 11590 17360 11610 17740
rect 11990 17360 12010 17740
rect 12390 17360 12410 17740
rect 12790 17360 12810 17740
rect 13190 17360 13210 17740
rect 13590 17360 13610 17740
rect 13990 17360 14010 17740
rect 14390 17360 14410 17740
rect 14790 17360 14810 17740
rect 15190 17360 15210 17740
rect 15590 17360 16000 17740
rect 0 17340 538 17360
rect 662 17340 938 17360
rect 1062 17340 1338 17360
rect 1462 17340 1738 17360
rect 1862 17340 2138 17360
rect 2262 17340 2538 17360
rect 2662 17340 2938 17360
rect 3062 17340 3338 17360
rect 3462 17340 3738 17360
rect 3862 17340 4138 17360
rect 4262 17340 4538 17360
rect 4662 17340 4938 17360
rect 5062 17340 5338 17360
rect 5462 17340 5738 17360
rect 5862 17340 6138 17360
rect 6262 17340 6538 17360
rect 6662 17340 6938 17360
rect 7062 17340 7338 17360
rect 7462 17340 7738 17360
rect 7862 17340 8138 17360
rect 8262 17340 8538 17360
rect 8662 17340 8938 17360
rect 9062 17340 9338 17360
rect 9462 17340 9738 17360
rect 9862 17340 10138 17360
rect 10262 17340 10538 17360
rect 10662 17340 10938 17360
rect 11062 17340 11338 17360
rect 11462 17340 11738 17360
rect 11862 17340 12138 17360
rect 12262 17340 12538 17360
rect 12662 17340 12938 17360
rect 13062 17340 13338 17360
rect 13462 17340 13738 17360
rect 13862 17340 14138 17360
rect 14262 17340 14538 17360
rect 14662 17340 14938 17360
rect 15062 17340 15338 17360
rect 15462 17340 16000 17360
rect 0 16960 410 17340
rect 790 16960 810 17340
rect 1190 16960 1210 17340
rect 1590 16960 1610 17340
rect 1990 16960 2010 17340
rect 2390 16960 2410 17340
rect 2790 16960 2810 17340
rect 3190 16960 3210 17340
rect 3590 16960 3610 17340
rect 3990 16960 4010 17340
rect 4390 16960 4410 17340
rect 4790 16960 4810 17340
rect 5190 16960 5210 17340
rect 5590 16960 5610 17340
rect 5990 16960 6010 17340
rect 6390 16960 6410 17340
rect 6790 16960 6810 17340
rect 7190 16960 7210 17340
rect 7590 16960 7610 17340
rect 7990 16960 8010 17340
rect 8390 16960 8410 17340
rect 8790 16960 8810 17340
rect 9190 16960 9210 17340
rect 9590 16960 9610 17340
rect 9990 16960 10010 17340
rect 10390 16960 10410 17340
rect 10790 16960 10810 17340
rect 11190 16960 11210 17340
rect 11590 16960 11610 17340
rect 11990 16960 12010 17340
rect 12390 16960 12410 17340
rect 12790 16960 12810 17340
rect 13190 16960 13210 17340
rect 13590 16960 13610 17340
rect 13990 16960 14010 17340
rect 14390 16960 14410 17340
rect 14790 16960 14810 17340
rect 15190 16960 15210 17340
rect 15590 16960 16000 17340
rect 0 16940 538 16960
rect 662 16940 938 16960
rect 1062 16940 1338 16960
rect 1462 16940 1738 16960
rect 1862 16940 2138 16960
rect 2262 16940 2538 16960
rect 2662 16940 2938 16960
rect 3062 16940 3338 16960
rect 3462 16940 3738 16960
rect 3862 16940 4138 16960
rect 4262 16940 4538 16960
rect 4662 16940 4938 16960
rect 5062 16940 5338 16960
rect 5462 16940 5738 16960
rect 5862 16940 6138 16960
rect 6262 16940 6538 16960
rect 6662 16940 6938 16960
rect 7062 16940 7338 16960
rect 7462 16940 7738 16960
rect 7862 16940 8138 16960
rect 8262 16940 8538 16960
rect 8662 16940 8938 16960
rect 9062 16940 9338 16960
rect 9462 16940 9738 16960
rect 9862 16940 10138 16960
rect 10262 16940 10538 16960
rect 10662 16940 10938 16960
rect 11062 16940 11338 16960
rect 11462 16940 11738 16960
rect 11862 16940 12138 16960
rect 12262 16940 12538 16960
rect 12662 16940 12938 16960
rect 13062 16940 13338 16960
rect 13462 16940 13738 16960
rect 13862 16940 14138 16960
rect 14262 16940 14538 16960
rect 14662 16940 14938 16960
rect 15062 16940 15338 16960
rect 15462 16940 16000 16960
rect 0 16560 410 16940
rect 790 16560 810 16940
rect 1190 16560 1210 16940
rect 1590 16560 1610 16940
rect 1990 16560 2010 16940
rect 2390 16560 2410 16940
rect 2790 16560 2810 16940
rect 3190 16560 3210 16940
rect 3590 16560 3610 16940
rect 3990 16560 4010 16940
rect 4390 16560 4410 16940
rect 4790 16560 4810 16940
rect 5190 16560 5210 16940
rect 5590 16560 5610 16940
rect 5990 16560 6010 16940
rect 6390 16560 6410 16940
rect 6790 16560 6810 16940
rect 7190 16560 7210 16940
rect 7590 16560 7610 16940
rect 7990 16560 8010 16940
rect 8390 16560 8410 16940
rect 8790 16560 8810 16940
rect 9190 16560 9210 16940
rect 9590 16560 9610 16940
rect 9990 16560 10010 16940
rect 10390 16560 10410 16940
rect 10790 16560 10810 16940
rect 11190 16560 11210 16940
rect 11590 16560 11610 16940
rect 11990 16560 12010 16940
rect 12390 16560 12410 16940
rect 12790 16560 12810 16940
rect 13190 16560 13210 16940
rect 13590 16560 13610 16940
rect 13990 16560 14010 16940
rect 14390 16560 14410 16940
rect 14790 16560 14810 16940
rect 15190 16560 15210 16940
rect 15590 16560 16000 16940
rect 0 16540 538 16560
rect 662 16540 938 16560
rect 1062 16540 1338 16560
rect 1462 16540 1738 16560
rect 1862 16540 2138 16560
rect 2262 16540 2538 16560
rect 2662 16540 2938 16560
rect 3062 16540 3338 16560
rect 3462 16540 3738 16560
rect 3862 16540 4138 16560
rect 4262 16540 4538 16560
rect 4662 16540 4938 16560
rect 5062 16540 5338 16560
rect 5462 16540 5738 16560
rect 5862 16540 6138 16560
rect 6262 16540 6538 16560
rect 6662 16540 6938 16560
rect 7062 16540 7338 16560
rect 7462 16540 7738 16560
rect 7862 16540 8138 16560
rect 8262 16540 8538 16560
rect 8662 16540 8938 16560
rect 9062 16540 9338 16560
rect 9462 16540 9738 16560
rect 9862 16540 10138 16560
rect 10262 16540 10538 16560
rect 10662 16540 10938 16560
rect 11062 16540 11338 16560
rect 11462 16540 11738 16560
rect 11862 16540 12138 16560
rect 12262 16540 12538 16560
rect 12662 16540 12938 16560
rect 13062 16540 13338 16560
rect 13462 16540 13738 16560
rect 13862 16540 14138 16560
rect 14262 16540 14538 16560
rect 14662 16540 14938 16560
rect 15062 16540 15338 16560
rect 15462 16540 16000 16560
rect 0 16160 410 16540
rect 790 16160 810 16540
rect 1190 16160 1210 16540
rect 1590 16160 1610 16540
rect 1990 16160 2010 16540
rect 2390 16160 2410 16540
rect 2790 16160 2810 16540
rect 3190 16160 3210 16540
rect 3590 16160 3610 16540
rect 3990 16160 4010 16540
rect 4390 16160 4410 16540
rect 4790 16160 4810 16540
rect 5190 16160 5210 16540
rect 5590 16160 5610 16540
rect 5990 16160 6010 16540
rect 6390 16160 6410 16540
rect 6790 16160 6810 16540
rect 7190 16160 7210 16540
rect 7590 16160 7610 16540
rect 7990 16160 8010 16540
rect 8390 16160 8410 16540
rect 8790 16160 8810 16540
rect 9190 16160 9210 16540
rect 9590 16160 9610 16540
rect 9990 16160 10010 16540
rect 10390 16160 10410 16540
rect 10790 16160 10810 16540
rect 11190 16160 11210 16540
rect 11590 16160 11610 16540
rect 11990 16160 12010 16540
rect 12390 16160 12410 16540
rect 12790 16160 12810 16540
rect 13190 16160 13210 16540
rect 13590 16160 13610 16540
rect 13990 16160 14010 16540
rect 14390 16160 14410 16540
rect 14790 16160 14810 16540
rect 15190 16160 15210 16540
rect 15590 16160 16000 16540
rect 0 16140 538 16160
rect 662 16140 938 16160
rect 1062 16140 1338 16160
rect 1462 16140 1738 16160
rect 1862 16140 2138 16160
rect 2262 16140 2538 16160
rect 2662 16140 2938 16160
rect 3062 16140 3338 16160
rect 3462 16140 3738 16160
rect 3862 16140 4138 16160
rect 4262 16140 4538 16160
rect 4662 16140 4938 16160
rect 5062 16140 5338 16160
rect 5462 16140 5738 16160
rect 5862 16140 6138 16160
rect 6262 16140 6538 16160
rect 6662 16140 6938 16160
rect 7062 16140 7338 16160
rect 7462 16140 7738 16160
rect 7862 16140 8138 16160
rect 8262 16140 8538 16160
rect 8662 16140 8938 16160
rect 9062 16140 9338 16160
rect 9462 16140 9738 16160
rect 9862 16140 10138 16160
rect 10262 16140 10538 16160
rect 10662 16140 10938 16160
rect 11062 16140 11338 16160
rect 11462 16140 11738 16160
rect 11862 16140 12138 16160
rect 12262 16140 12538 16160
rect 12662 16140 12938 16160
rect 13062 16140 13338 16160
rect 13462 16140 13738 16160
rect 13862 16140 14138 16160
rect 14262 16140 14538 16160
rect 14662 16140 14938 16160
rect 15062 16140 15338 16160
rect 15462 16140 16000 16160
rect 0 15760 410 16140
rect 790 15760 810 16140
rect 1190 15760 1210 16140
rect 1590 15760 1610 16140
rect 1990 15760 2010 16140
rect 2390 15760 2410 16140
rect 2790 15760 2810 16140
rect 3190 15760 3210 16140
rect 3590 15760 3610 16140
rect 3990 15760 4010 16140
rect 4390 15760 4410 16140
rect 4790 15760 4810 16140
rect 5190 15760 5210 16140
rect 5590 15760 5610 16140
rect 5990 15760 6010 16140
rect 6390 15760 6410 16140
rect 6790 15760 6810 16140
rect 7190 15760 7210 16140
rect 7590 15760 7610 16140
rect 7990 15760 8010 16140
rect 8390 15760 8410 16140
rect 8790 15760 8810 16140
rect 9190 15760 9210 16140
rect 9590 15760 9610 16140
rect 9990 15760 10010 16140
rect 10390 15760 10410 16140
rect 10790 15760 10810 16140
rect 11190 15760 11210 16140
rect 11590 15760 11610 16140
rect 11990 15760 12010 16140
rect 12390 15760 12410 16140
rect 12790 15760 12810 16140
rect 13190 15760 13210 16140
rect 13590 15760 13610 16140
rect 13990 15760 14010 16140
rect 14390 15760 14410 16140
rect 14790 15760 14810 16140
rect 15190 15760 15210 16140
rect 15590 15760 16000 16140
rect 0 15740 538 15760
rect 662 15740 938 15760
rect 1062 15740 1338 15760
rect 1462 15740 1738 15760
rect 1862 15740 2138 15760
rect 2262 15740 2538 15760
rect 2662 15740 2938 15760
rect 3062 15740 3338 15760
rect 3462 15740 3738 15760
rect 3862 15740 4138 15760
rect 4262 15740 4538 15760
rect 4662 15740 4938 15760
rect 5062 15740 5338 15760
rect 5462 15740 5738 15760
rect 5862 15740 6138 15760
rect 6262 15740 6538 15760
rect 6662 15740 6938 15760
rect 7062 15740 7338 15760
rect 7462 15740 7738 15760
rect 7862 15740 8138 15760
rect 8262 15740 8538 15760
rect 8662 15740 8938 15760
rect 9062 15740 9338 15760
rect 9462 15740 9738 15760
rect 9862 15740 10138 15760
rect 10262 15740 10538 15760
rect 10662 15740 10938 15760
rect 11062 15740 11338 15760
rect 11462 15740 11738 15760
rect 11862 15740 12138 15760
rect 12262 15740 12538 15760
rect 12662 15740 12938 15760
rect 13062 15740 13338 15760
rect 13462 15740 13738 15760
rect 13862 15740 14138 15760
rect 14262 15740 14538 15760
rect 14662 15740 14938 15760
rect 15062 15740 15338 15760
rect 15462 15740 16000 15760
rect 0 15360 410 15740
rect 790 15360 810 15740
rect 1190 15360 1210 15740
rect 1590 15360 1610 15740
rect 1990 15360 2010 15740
rect 2390 15360 2410 15740
rect 2790 15360 2810 15740
rect 3190 15360 3210 15740
rect 3590 15360 3610 15740
rect 3990 15360 4010 15740
rect 4390 15360 4410 15740
rect 4790 15360 4810 15740
rect 5190 15360 5210 15740
rect 5590 15360 5610 15740
rect 5990 15360 6010 15740
rect 6390 15360 6410 15740
rect 6790 15360 6810 15740
rect 7190 15360 7210 15740
rect 7590 15360 7610 15740
rect 7990 15360 8010 15740
rect 8390 15360 8410 15740
rect 8790 15360 8810 15740
rect 9190 15360 9210 15740
rect 9590 15360 9610 15740
rect 9990 15360 10010 15740
rect 10390 15360 10410 15740
rect 10790 15360 10810 15740
rect 11190 15360 11210 15740
rect 11590 15360 11610 15740
rect 11990 15360 12010 15740
rect 12390 15360 12410 15740
rect 12790 15360 12810 15740
rect 13190 15360 13210 15740
rect 13590 15360 13610 15740
rect 13990 15360 14010 15740
rect 14390 15360 14410 15740
rect 14790 15360 14810 15740
rect 15190 15360 15210 15740
rect 15590 15360 16000 15740
rect 0 15340 538 15360
rect 662 15340 938 15360
rect 1062 15340 1338 15360
rect 1462 15340 1738 15360
rect 1862 15340 2138 15360
rect 2262 15340 2538 15360
rect 2662 15340 2938 15360
rect 3062 15340 3338 15360
rect 3462 15340 3738 15360
rect 3862 15340 4138 15360
rect 4262 15340 4538 15360
rect 4662 15340 4938 15360
rect 5062 15340 5338 15360
rect 5462 15340 5738 15360
rect 5862 15340 6138 15360
rect 6262 15340 6538 15360
rect 6662 15340 6938 15360
rect 7062 15340 7338 15360
rect 7462 15340 7738 15360
rect 7862 15340 8138 15360
rect 8262 15340 8538 15360
rect 8662 15340 8938 15360
rect 9062 15340 9338 15360
rect 9462 15340 9738 15360
rect 9862 15340 10138 15360
rect 10262 15340 10538 15360
rect 10662 15340 10938 15360
rect 11062 15340 11338 15360
rect 11462 15340 11738 15360
rect 11862 15340 12138 15360
rect 12262 15340 12538 15360
rect 12662 15340 12938 15360
rect 13062 15340 13338 15360
rect 13462 15340 13738 15360
rect 13862 15340 14138 15360
rect 14262 15340 14538 15360
rect 14662 15340 14938 15360
rect 15062 15340 15338 15360
rect 15462 15340 16000 15360
rect 0 14960 410 15340
rect 790 14960 810 15340
rect 1190 14960 1210 15340
rect 1590 14960 1610 15340
rect 1990 14960 2010 15340
rect 2390 14960 2410 15340
rect 2790 14960 2810 15340
rect 3190 14960 3210 15340
rect 3590 14960 3610 15340
rect 3990 14960 4010 15340
rect 4390 14960 4410 15340
rect 4790 14960 4810 15340
rect 5190 14960 5210 15340
rect 5590 14960 5610 15340
rect 5990 14960 6010 15340
rect 6390 14960 6410 15340
rect 6790 14960 6810 15340
rect 7190 14960 7210 15340
rect 7590 14960 7610 15340
rect 7990 14960 8010 15340
rect 8390 14960 8410 15340
rect 8790 14960 8810 15340
rect 9190 14960 9210 15340
rect 9590 14960 9610 15340
rect 9990 14960 10010 15340
rect 10390 14960 10410 15340
rect 10790 14960 10810 15340
rect 11190 14960 11210 15340
rect 11590 14960 11610 15340
rect 11990 14960 12010 15340
rect 12390 14960 12410 15340
rect 12790 14960 12810 15340
rect 13190 14960 13210 15340
rect 13590 14960 13610 15340
rect 13990 14960 14010 15340
rect 14390 14960 14410 15340
rect 14790 14960 14810 15340
rect 15190 14960 15210 15340
rect 15590 14960 16000 15340
rect 0 14940 538 14960
rect 662 14940 938 14960
rect 1062 14940 1338 14960
rect 1462 14940 1738 14960
rect 1862 14940 2138 14960
rect 2262 14940 2538 14960
rect 2662 14940 2938 14960
rect 3062 14940 3338 14960
rect 3462 14940 3738 14960
rect 3862 14940 4138 14960
rect 4262 14940 4538 14960
rect 4662 14940 4938 14960
rect 5062 14940 5338 14960
rect 5462 14940 5738 14960
rect 5862 14940 6138 14960
rect 6262 14940 6538 14960
rect 6662 14940 6938 14960
rect 7062 14940 7338 14960
rect 7462 14940 7738 14960
rect 7862 14940 8138 14960
rect 8262 14940 8538 14960
rect 8662 14940 8938 14960
rect 9062 14940 9338 14960
rect 9462 14940 9738 14960
rect 9862 14940 10138 14960
rect 10262 14940 10538 14960
rect 10662 14940 10938 14960
rect 11062 14940 11338 14960
rect 11462 14940 11738 14960
rect 11862 14940 12138 14960
rect 12262 14940 12538 14960
rect 12662 14940 12938 14960
rect 13062 14940 13338 14960
rect 13462 14940 13738 14960
rect 13862 14940 14138 14960
rect 14262 14940 14538 14960
rect 14662 14940 14938 14960
rect 15062 14940 15338 14960
rect 15462 14940 16000 14960
rect 0 14560 410 14940
rect 790 14560 810 14940
rect 1190 14560 1210 14940
rect 1590 14560 1610 14940
rect 1990 14560 2010 14940
rect 2390 14560 2410 14940
rect 2790 14560 2810 14940
rect 3190 14560 3210 14940
rect 3590 14560 3610 14940
rect 3990 14560 4010 14940
rect 4390 14560 4410 14940
rect 4790 14560 4810 14940
rect 5190 14560 5210 14940
rect 5590 14560 5610 14940
rect 5990 14560 6010 14940
rect 6390 14560 6410 14940
rect 6790 14560 6810 14940
rect 7190 14560 7210 14940
rect 7590 14560 7610 14940
rect 7990 14560 8010 14940
rect 8390 14560 8410 14940
rect 8790 14560 8810 14940
rect 9190 14560 9210 14940
rect 9590 14560 9610 14940
rect 9990 14560 10010 14940
rect 10390 14560 10410 14940
rect 10790 14560 10810 14940
rect 11190 14560 11210 14940
rect 11590 14560 11610 14940
rect 11990 14560 12010 14940
rect 12390 14560 12410 14940
rect 12790 14560 12810 14940
rect 13190 14560 13210 14940
rect 13590 14560 13610 14940
rect 13990 14560 14010 14940
rect 14390 14560 14410 14940
rect 14790 14560 14810 14940
rect 15190 14560 15210 14940
rect 15590 14560 16000 14940
rect 0 14540 538 14560
rect 662 14540 938 14560
rect 1062 14540 1338 14560
rect 1462 14540 1738 14560
rect 1862 14540 2138 14560
rect 2262 14540 2538 14560
rect 2662 14540 2938 14560
rect 3062 14540 3338 14560
rect 3462 14540 3738 14560
rect 3862 14540 4138 14560
rect 4262 14540 4538 14560
rect 4662 14540 4938 14560
rect 5062 14540 5338 14560
rect 5462 14540 5738 14560
rect 5862 14540 6138 14560
rect 6262 14540 6538 14560
rect 6662 14540 6938 14560
rect 7062 14540 7338 14560
rect 7462 14540 7738 14560
rect 7862 14540 8138 14560
rect 8262 14540 8538 14560
rect 8662 14540 8938 14560
rect 9062 14540 9338 14560
rect 9462 14540 9738 14560
rect 9862 14540 10138 14560
rect 10262 14540 10538 14560
rect 10662 14540 10938 14560
rect 11062 14540 11338 14560
rect 11462 14540 11738 14560
rect 11862 14540 12138 14560
rect 12262 14540 12538 14560
rect 12662 14540 12938 14560
rect 13062 14540 13338 14560
rect 13462 14540 13738 14560
rect 13862 14540 14138 14560
rect 14262 14540 14538 14560
rect 14662 14540 14938 14560
rect 15062 14540 15338 14560
rect 15462 14540 16000 14560
rect 0 14160 410 14540
rect 790 14160 810 14540
rect 1190 14160 1210 14540
rect 1590 14160 1610 14540
rect 1990 14160 2010 14540
rect 2390 14160 2410 14540
rect 2790 14160 2810 14540
rect 3190 14160 3210 14540
rect 3590 14160 3610 14540
rect 3990 14160 4010 14540
rect 4390 14160 4410 14540
rect 4790 14160 4810 14540
rect 5190 14160 5210 14540
rect 5590 14160 5610 14540
rect 5990 14160 6010 14540
rect 6390 14160 6410 14540
rect 6790 14160 6810 14540
rect 7190 14160 7210 14540
rect 7590 14160 7610 14540
rect 7990 14160 8010 14540
rect 8390 14160 8410 14540
rect 8790 14160 8810 14540
rect 9190 14160 9210 14540
rect 9590 14160 9610 14540
rect 9990 14160 10010 14540
rect 10390 14160 10410 14540
rect 10790 14160 10810 14540
rect 11190 14160 11210 14540
rect 11590 14160 11610 14540
rect 11990 14160 12010 14540
rect 12390 14160 12410 14540
rect 12790 14160 12810 14540
rect 13190 14160 13210 14540
rect 13590 14160 13610 14540
rect 13990 14160 14010 14540
rect 14390 14160 14410 14540
rect 14790 14160 14810 14540
rect 15190 14160 15210 14540
rect 15590 14160 16000 14540
rect 0 14140 538 14160
rect 662 14140 938 14160
rect 1062 14140 1338 14160
rect 1462 14140 1738 14160
rect 1862 14140 2138 14160
rect 2262 14140 2538 14160
rect 2662 14140 2938 14160
rect 3062 14140 3338 14160
rect 3462 14140 3738 14160
rect 3862 14140 4138 14160
rect 4262 14140 4538 14160
rect 4662 14140 4938 14160
rect 5062 14140 5338 14160
rect 5462 14140 5738 14160
rect 5862 14140 6138 14160
rect 6262 14140 6538 14160
rect 6662 14140 6938 14160
rect 7062 14140 7338 14160
rect 7462 14140 7738 14160
rect 7862 14140 8138 14160
rect 8262 14140 8538 14160
rect 8662 14140 8938 14160
rect 9062 14140 9338 14160
rect 9462 14140 9738 14160
rect 9862 14140 10138 14160
rect 10262 14140 10538 14160
rect 10662 14140 10938 14160
rect 11062 14140 11338 14160
rect 11462 14140 11738 14160
rect 11862 14140 12138 14160
rect 12262 14140 12538 14160
rect 12662 14140 12938 14160
rect 13062 14140 13338 14160
rect 13462 14140 13738 14160
rect 13862 14140 14138 14160
rect 14262 14140 14538 14160
rect 14662 14140 14938 14160
rect 15062 14140 15338 14160
rect 15462 14140 16000 14160
rect 0 13760 410 14140
rect 790 13760 810 14140
rect 1190 13760 1210 14140
rect 1590 13760 1610 14140
rect 1990 13760 2010 14140
rect 2390 13760 2410 14140
rect 2790 13760 2810 14140
rect 3190 13760 3210 14140
rect 3590 13760 3610 14140
rect 3990 13760 4010 14140
rect 4390 13760 4410 14140
rect 4790 13760 4810 14140
rect 5190 13760 5210 14140
rect 5590 13760 5610 14140
rect 5990 13760 6010 14140
rect 6390 13760 6410 14140
rect 6790 13760 6810 14140
rect 7190 13760 7210 14140
rect 7590 13760 7610 14140
rect 7990 13760 8010 14140
rect 8390 13760 8410 14140
rect 8790 13760 8810 14140
rect 9190 13760 9210 14140
rect 9590 13760 9610 14140
rect 9990 13760 10010 14140
rect 10390 13760 10410 14140
rect 10790 13760 10810 14140
rect 11190 13760 11210 14140
rect 11590 13760 11610 14140
rect 11990 13760 12010 14140
rect 12390 13760 12410 14140
rect 12790 13760 12810 14140
rect 13190 13760 13210 14140
rect 13590 13760 13610 14140
rect 13990 13760 14010 14140
rect 14390 13760 14410 14140
rect 14790 13760 14810 14140
rect 15190 13760 15210 14140
rect 15590 13760 16000 14140
rect 0 13688 538 13760
rect 662 13688 938 13760
rect 1062 13688 1338 13760
rect 1462 13688 1738 13760
rect 1862 13688 2138 13760
rect 2262 13688 2538 13760
rect 2662 13688 2938 13760
rect 3062 13688 3338 13760
rect 3462 13688 3738 13760
rect 3862 13688 4138 13760
rect 4262 13688 4538 13760
rect 4662 13688 4938 13760
rect 5062 13688 5338 13760
rect 5462 13688 5738 13760
rect 5862 13688 6138 13760
rect 6262 13688 6538 13760
rect 6662 13688 6938 13760
rect 7062 13688 7338 13760
rect 7462 13688 7738 13760
rect 7862 13688 8138 13760
rect 8262 13688 8538 13760
rect 8662 13688 8938 13760
rect 9062 13688 9338 13760
rect 9462 13688 9738 13760
rect 9862 13688 10138 13760
rect 10262 13688 10538 13760
rect 10662 13688 10938 13760
rect 11062 13688 11338 13760
rect 11462 13688 11738 13760
rect 11862 13688 12138 13760
rect 12262 13688 12538 13760
rect 12662 13688 12938 13760
rect 13062 13688 13338 13760
rect 13462 13688 13738 13760
rect 13862 13688 14138 13760
rect 14262 13688 14538 13760
rect 14662 13688 14938 13760
rect 15062 13688 15338 13760
rect 15462 13688 16000 13760
rect 0 13200 16000 13688
rect 0 11640 16000 12000
rect 380 11260 400 11640
rect 780 11512 15220 11640
rect 780 11388 938 11512
rect 1062 11388 1338 11512
rect 1462 11388 1738 11512
rect 1862 11388 2138 11512
rect 2262 11388 2538 11512
rect 2662 11388 2938 11512
rect 3062 11388 3338 11512
rect 3462 11388 3738 11512
rect 3862 11388 4138 11512
rect 4262 11388 4538 11512
rect 4662 11388 4938 11512
rect 5062 11388 5338 11512
rect 5462 11388 5738 11512
rect 5862 11388 6138 11512
rect 6262 11388 6538 11512
rect 6662 11388 6938 11512
rect 7062 11388 7338 11512
rect 7462 11388 7738 11512
rect 7862 11388 8138 11512
rect 8262 11388 8538 11512
rect 8662 11388 8938 11512
rect 9062 11388 9338 11512
rect 9462 11388 9738 11512
rect 9862 11388 10138 11512
rect 10262 11388 10538 11512
rect 10662 11388 10938 11512
rect 11062 11388 11338 11512
rect 11462 11388 11738 11512
rect 11862 11388 12138 11512
rect 12262 11388 12538 11512
rect 12662 11388 12938 11512
rect 13062 11388 13338 11512
rect 13462 11388 13738 11512
rect 13862 11388 14138 11512
rect 14262 11388 14538 11512
rect 14662 11388 14938 11512
rect 15062 11388 15220 11512
rect 780 11260 15220 11388
rect 15600 11260 15620 11640
rect 0 11240 16000 11260
rect 380 10860 400 11240
rect 780 11112 15220 11240
rect 780 10988 938 11112
rect 1062 10988 1338 11112
rect 1462 10988 1738 11112
rect 1862 10988 2138 11112
rect 2262 10988 2538 11112
rect 2662 10988 2938 11112
rect 3062 10988 3338 11112
rect 3462 10988 3738 11112
rect 3862 10988 4138 11112
rect 4262 10988 4538 11112
rect 4662 10988 4938 11112
rect 5062 10988 5338 11112
rect 5462 10988 5738 11112
rect 5862 10988 6138 11112
rect 6262 10988 6538 11112
rect 6662 10988 6938 11112
rect 7062 10988 7338 11112
rect 7462 10988 7738 11112
rect 7862 10988 8138 11112
rect 8262 10988 8538 11112
rect 8662 10988 8938 11112
rect 9062 10988 9338 11112
rect 9462 10988 9738 11112
rect 9862 10988 10138 11112
rect 10262 10988 10538 11112
rect 10662 10988 10938 11112
rect 11062 10988 11338 11112
rect 11462 10988 11738 11112
rect 11862 10988 12138 11112
rect 12262 10988 12538 11112
rect 12662 10988 12938 11112
rect 13062 10988 13338 11112
rect 13462 10988 13738 11112
rect 13862 10988 14138 11112
rect 14262 10988 14538 11112
rect 14662 10988 14938 11112
rect 15062 10988 15220 11112
rect 780 10860 15220 10988
rect 15600 10860 15620 11240
rect 0 10840 16000 10860
rect 380 10460 400 10840
rect 780 10712 15220 10840
rect 780 10588 938 10712
rect 1062 10588 1338 10712
rect 1462 10588 1738 10712
rect 1862 10588 2138 10712
rect 2262 10588 2538 10712
rect 2662 10588 2938 10712
rect 3062 10588 3338 10712
rect 3462 10588 3738 10712
rect 3862 10588 4138 10712
rect 4262 10588 4538 10712
rect 4662 10588 4938 10712
rect 5062 10588 5338 10712
rect 5462 10588 5738 10712
rect 5862 10588 6138 10712
rect 6262 10588 6538 10712
rect 6662 10588 6938 10712
rect 7062 10588 7338 10712
rect 7462 10588 7738 10712
rect 7862 10588 8138 10712
rect 8262 10588 8538 10712
rect 8662 10588 8938 10712
rect 9062 10588 9338 10712
rect 9462 10588 9738 10712
rect 9862 10588 10138 10712
rect 10262 10588 10538 10712
rect 10662 10588 10938 10712
rect 11062 10588 11338 10712
rect 11462 10588 11738 10712
rect 11862 10588 12138 10712
rect 12262 10588 12538 10712
rect 12662 10588 12938 10712
rect 13062 10588 13338 10712
rect 13462 10588 13738 10712
rect 13862 10588 14138 10712
rect 14262 10588 14538 10712
rect 14662 10588 14938 10712
rect 15062 10588 15220 10712
rect 780 10460 15220 10588
rect 15600 10460 15620 10840
rect 0 10440 16000 10460
rect 380 10060 400 10440
rect 780 10312 15220 10440
rect 780 10188 938 10312
rect 1062 10188 1338 10312
rect 1462 10188 1738 10312
rect 1862 10188 2138 10312
rect 2262 10188 2538 10312
rect 2662 10188 2938 10312
rect 3062 10188 3338 10312
rect 3462 10188 3738 10312
rect 3862 10188 4138 10312
rect 4262 10188 4538 10312
rect 4662 10188 4938 10312
rect 5062 10188 5338 10312
rect 5462 10188 5738 10312
rect 5862 10188 6138 10312
rect 6262 10188 6538 10312
rect 6662 10188 6938 10312
rect 7062 10188 7338 10312
rect 7462 10188 7738 10312
rect 7862 10188 8138 10312
rect 8262 10188 8538 10312
rect 8662 10188 8938 10312
rect 9062 10188 9338 10312
rect 9462 10188 9738 10312
rect 9862 10188 10138 10312
rect 10262 10188 10538 10312
rect 10662 10188 10938 10312
rect 11062 10188 11338 10312
rect 11462 10188 11738 10312
rect 11862 10188 12138 10312
rect 12262 10188 12538 10312
rect 12662 10188 12938 10312
rect 13062 10188 13338 10312
rect 13462 10188 13738 10312
rect 13862 10188 14138 10312
rect 14262 10188 14538 10312
rect 14662 10188 14938 10312
rect 15062 10188 15220 10312
rect 780 10060 15220 10188
rect 15600 10060 15620 10440
rect 0 10040 16000 10060
rect 380 9660 400 10040
rect 780 9912 15220 10040
rect 780 9788 938 9912
rect 1062 9788 1338 9912
rect 1462 9788 1738 9912
rect 1862 9788 2138 9912
rect 2262 9788 2538 9912
rect 2662 9788 2938 9912
rect 3062 9788 3338 9912
rect 3462 9788 3738 9912
rect 3862 9788 4138 9912
rect 4262 9788 4538 9912
rect 4662 9788 4938 9912
rect 5062 9788 5338 9912
rect 5462 9788 5738 9912
rect 5862 9788 6138 9912
rect 6262 9788 6538 9912
rect 6662 9788 6938 9912
rect 7062 9788 7338 9912
rect 7462 9788 7738 9912
rect 7862 9788 8138 9912
rect 8262 9788 8538 9912
rect 8662 9788 8938 9912
rect 9062 9788 9338 9912
rect 9462 9788 9738 9912
rect 9862 9788 10138 9912
rect 10262 9788 10538 9912
rect 10662 9788 10938 9912
rect 11062 9788 11338 9912
rect 11462 9788 11738 9912
rect 11862 9788 12138 9912
rect 12262 9788 12538 9912
rect 12662 9788 12938 9912
rect 13062 9788 13338 9912
rect 13462 9788 13738 9912
rect 13862 9788 14138 9912
rect 14262 9788 14538 9912
rect 14662 9788 14938 9912
rect 15062 9788 15220 9912
rect 780 9660 15220 9788
rect 15600 9660 15620 10040
rect 0 9640 16000 9660
rect 380 9260 400 9640
rect 780 9512 15220 9640
rect 780 9388 938 9512
rect 1062 9388 1338 9512
rect 1462 9388 1738 9512
rect 1862 9388 2138 9512
rect 2262 9388 2538 9512
rect 2662 9388 2938 9512
rect 3062 9388 3338 9512
rect 3462 9388 3738 9512
rect 3862 9388 4138 9512
rect 4262 9388 4538 9512
rect 4662 9388 4938 9512
rect 5062 9388 5338 9512
rect 5462 9388 5738 9512
rect 5862 9388 6138 9512
rect 6262 9388 6538 9512
rect 6662 9388 6938 9512
rect 7062 9388 7338 9512
rect 7462 9388 7738 9512
rect 7862 9388 8138 9512
rect 8262 9388 8538 9512
rect 8662 9388 8938 9512
rect 9062 9388 9338 9512
rect 9462 9388 9738 9512
rect 9862 9388 10138 9512
rect 10262 9388 10538 9512
rect 10662 9388 10938 9512
rect 11062 9388 11338 9512
rect 11462 9388 11738 9512
rect 11862 9388 12138 9512
rect 12262 9388 12538 9512
rect 12662 9388 12938 9512
rect 13062 9388 13338 9512
rect 13462 9388 13738 9512
rect 13862 9388 14138 9512
rect 14262 9388 14538 9512
rect 14662 9388 14938 9512
rect 15062 9388 15220 9512
rect 780 9260 15220 9388
rect 15600 9260 15620 9640
rect 0 9240 16000 9260
rect 380 8860 400 9240
rect 780 9112 15220 9240
rect 780 8988 938 9112
rect 1062 8988 1338 9112
rect 1462 8988 1738 9112
rect 1862 8988 2138 9112
rect 2262 8988 2538 9112
rect 2662 8988 2938 9112
rect 3062 8988 3338 9112
rect 3462 8988 3738 9112
rect 3862 8988 4138 9112
rect 4262 8988 4538 9112
rect 4662 8988 4938 9112
rect 5062 8988 5338 9112
rect 5462 8988 5738 9112
rect 5862 8988 6138 9112
rect 6262 8988 6538 9112
rect 6662 8988 6938 9112
rect 7062 8988 7338 9112
rect 7462 8988 7738 9112
rect 7862 8988 8138 9112
rect 8262 8988 8538 9112
rect 8662 8988 8938 9112
rect 9062 8988 9338 9112
rect 9462 8988 9738 9112
rect 9862 8988 10138 9112
rect 10262 8988 10538 9112
rect 10662 8988 10938 9112
rect 11062 8988 11338 9112
rect 11462 8988 11738 9112
rect 11862 8988 12138 9112
rect 12262 8988 12538 9112
rect 12662 8988 12938 9112
rect 13062 8988 13338 9112
rect 13462 8988 13738 9112
rect 13862 8988 14138 9112
rect 14262 8988 14538 9112
rect 14662 8988 14938 9112
rect 15062 8988 15220 9112
rect 780 8860 15220 8988
rect 15600 8860 15620 9240
rect 0 8840 16000 8860
rect 380 8460 400 8840
rect 780 8712 15220 8840
rect 780 8588 938 8712
rect 1062 8588 1338 8712
rect 1462 8588 1738 8712
rect 1862 8588 2138 8712
rect 2262 8588 2538 8712
rect 2662 8588 2938 8712
rect 3062 8588 3338 8712
rect 3462 8588 3738 8712
rect 3862 8588 4138 8712
rect 4262 8588 4538 8712
rect 4662 8588 4938 8712
rect 5062 8588 5338 8712
rect 5462 8588 5738 8712
rect 5862 8588 6138 8712
rect 6262 8588 6538 8712
rect 6662 8588 6938 8712
rect 7062 8588 7338 8712
rect 7462 8588 7738 8712
rect 7862 8588 8138 8712
rect 8262 8588 8538 8712
rect 8662 8588 8938 8712
rect 9062 8588 9338 8712
rect 9462 8588 9738 8712
rect 9862 8588 10138 8712
rect 10262 8588 10538 8712
rect 10662 8588 10938 8712
rect 11062 8588 11338 8712
rect 11462 8588 11738 8712
rect 11862 8588 12138 8712
rect 12262 8588 12538 8712
rect 12662 8588 12938 8712
rect 13062 8588 13338 8712
rect 13462 8588 13738 8712
rect 13862 8588 14138 8712
rect 14262 8588 14538 8712
rect 14662 8588 14938 8712
rect 15062 8588 15220 8712
rect 780 8460 15220 8588
rect 15600 8460 15620 8840
rect 0 8440 16000 8460
rect 380 8060 400 8440
rect 780 8312 15220 8440
rect 780 8188 938 8312
rect 1062 8188 1338 8312
rect 1462 8188 1738 8312
rect 1862 8188 2138 8312
rect 2262 8188 2538 8312
rect 2662 8188 2938 8312
rect 3062 8188 3338 8312
rect 3462 8188 3738 8312
rect 3862 8188 4138 8312
rect 4262 8188 4538 8312
rect 4662 8188 4938 8312
rect 5062 8188 5338 8312
rect 5462 8188 5738 8312
rect 5862 8188 6138 8312
rect 6262 8188 6538 8312
rect 6662 8188 6938 8312
rect 7062 8188 7338 8312
rect 7462 8188 7738 8312
rect 7862 8188 8138 8312
rect 8262 8188 8538 8312
rect 8662 8188 8938 8312
rect 9062 8188 9338 8312
rect 9462 8188 9738 8312
rect 9862 8188 10138 8312
rect 10262 8188 10538 8312
rect 10662 8188 10938 8312
rect 11062 8188 11338 8312
rect 11462 8188 11738 8312
rect 11862 8188 12138 8312
rect 12262 8188 12538 8312
rect 12662 8188 12938 8312
rect 13062 8188 13338 8312
rect 13462 8188 13738 8312
rect 13862 8188 14138 8312
rect 14262 8188 14538 8312
rect 14662 8188 14938 8312
rect 15062 8188 15220 8312
rect 780 8060 15220 8188
rect 15600 8060 15620 8440
rect 0 8040 16000 8060
rect 380 7660 400 8040
rect 780 7912 15220 8040
rect 780 7788 938 7912
rect 1062 7788 1338 7912
rect 1462 7788 1738 7912
rect 1862 7788 2138 7912
rect 2262 7788 2538 7912
rect 2662 7788 2938 7912
rect 3062 7788 3338 7912
rect 3462 7788 3738 7912
rect 3862 7788 4138 7912
rect 4262 7788 4538 7912
rect 4662 7788 4938 7912
rect 5062 7788 5338 7912
rect 5462 7788 5738 7912
rect 5862 7788 6138 7912
rect 6262 7788 6538 7912
rect 6662 7788 6938 7912
rect 7062 7788 7338 7912
rect 7462 7788 7738 7912
rect 7862 7788 8138 7912
rect 8262 7788 8538 7912
rect 8662 7788 8938 7912
rect 9062 7788 9338 7912
rect 9462 7788 9738 7912
rect 9862 7788 10138 7912
rect 10262 7788 10538 7912
rect 10662 7788 10938 7912
rect 11062 7788 11338 7912
rect 11462 7788 11738 7912
rect 11862 7788 12138 7912
rect 12262 7788 12538 7912
rect 12662 7788 12938 7912
rect 13062 7788 13338 7912
rect 13462 7788 13738 7912
rect 13862 7788 14138 7912
rect 14262 7788 14538 7912
rect 14662 7788 14938 7912
rect 15062 7788 15220 7912
rect 780 7660 15220 7788
rect 15600 7660 15620 8040
rect 0 7640 16000 7660
rect 380 7260 400 7640
rect 780 7512 15220 7640
rect 780 7388 938 7512
rect 1062 7388 1338 7512
rect 1462 7388 1738 7512
rect 1862 7388 2138 7512
rect 2262 7388 2538 7512
rect 2662 7388 2938 7512
rect 3062 7388 3338 7512
rect 3462 7388 3738 7512
rect 3862 7388 4138 7512
rect 4262 7388 4538 7512
rect 4662 7388 4938 7512
rect 5062 7388 5338 7512
rect 5462 7388 5738 7512
rect 5862 7388 6138 7512
rect 6262 7388 6538 7512
rect 6662 7388 6938 7512
rect 7062 7388 7338 7512
rect 7462 7388 7738 7512
rect 7862 7388 8138 7512
rect 8262 7388 8538 7512
rect 8662 7388 8938 7512
rect 9062 7388 9338 7512
rect 9462 7388 9738 7512
rect 9862 7388 10138 7512
rect 10262 7388 10538 7512
rect 10662 7388 10938 7512
rect 11062 7388 11338 7512
rect 11462 7388 11738 7512
rect 11862 7388 12138 7512
rect 12262 7388 12538 7512
rect 12662 7388 12938 7512
rect 13062 7388 13338 7512
rect 13462 7388 13738 7512
rect 13862 7388 14138 7512
rect 14262 7388 14538 7512
rect 14662 7388 14938 7512
rect 15062 7388 15220 7512
rect 780 7260 15220 7388
rect 15600 7260 15620 7640
rect 0 6900 16000 7260
rect 0 6140 16000 6500
rect 380 5760 400 6140
rect 780 6012 15220 6140
rect 780 5888 938 6012
rect 1062 5888 1338 6012
rect 1462 5888 1738 6012
rect 1862 5888 2138 6012
rect 2262 5888 2538 6012
rect 2662 5888 2938 6012
rect 3062 5888 3338 6012
rect 3462 5888 3738 6012
rect 3862 5888 4138 6012
rect 4262 5888 4538 6012
rect 4662 5888 4938 6012
rect 5062 5888 5338 6012
rect 5462 5888 5738 6012
rect 5862 5888 6138 6012
rect 6262 5888 6538 6012
rect 6662 5888 6938 6012
rect 7062 5888 7338 6012
rect 7462 5888 7738 6012
rect 7862 5888 8138 6012
rect 8262 5888 8538 6012
rect 8662 5888 8938 6012
rect 9062 5888 9338 6012
rect 9462 5888 9738 6012
rect 9862 5888 10138 6012
rect 10262 5888 10538 6012
rect 10662 5888 10938 6012
rect 11062 5888 11338 6012
rect 11462 5888 11738 6012
rect 11862 5888 12138 6012
rect 12262 5888 12538 6012
rect 12662 5888 12938 6012
rect 13062 5888 13338 6012
rect 13462 5888 13738 6012
rect 13862 5888 14138 6012
rect 14262 5888 14538 6012
rect 14662 5888 14938 6012
rect 15062 5888 15220 6012
rect 780 5760 15220 5888
rect 15600 5760 15620 6140
rect 0 5740 16000 5760
rect 380 5360 400 5740
rect 780 5612 15220 5740
rect 780 5488 938 5612
rect 1062 5488 1338 5612
rect 1462 5488 1738 5612
rect 1862 5488 2138 5612
rect 2262 5488 2538 5612
rect 2662 5488 2938 5612
rect 3062 5488 3338 5612
rect 3462 5488 3738 5612
rect 3862 5488 4138 5612
rect 4262 5488 4538 5612
rect 4662 5488 4938 5612
rect 5062 5488 5338 5612
rect 5462 5488 5738 5612
rect 5862 5488 6138 5612
rect 6262 5488 6538 5612
rect 6662 5488 6938 5612
rect 7062 5488 7338 5612
rect 7462 5488 7738 5612
rect 7862 5488 8138 5612
rect 8262 5488 8538 5612
rect 8662 5488 8938 5612
rect 9062 5488 9338 5612
rect 9462 5488 9738 5612
rect 9862 5488 10138 5612
rect 10262 5488 10538 5612
rect 10662 5488 10938 5612
rect 11062 5488 11338 5612
rect 11462 5488 11738 5612
rect 11862 5488 12138 5612
rect 12262 5488 12538 5612
rect 12662 5488 12938 5612
rect 13062 5488 13338 5612
rect 13462 5488 13738 5612
rect 13862 5488 14138 5612
rect 14262 5488 14538 5612
rect 14662 5488 14938 5612
rect 15062 5488 15220 5612
rect 780 5360 15220 5488
rect 15600 5360 15620 5740
rect 0 5340 16000 5360
rect 380 4960 400 5340
rect 780 5212 15220 5340
rect 780 5088 938 5212
rect 1062 5088 1338 5212
rect 1462 5088 1738 5212
rect 1862 5088 2138 5212
rect 2262 5088 2538 5212
rect 2662 5088 2938 5212
rect 3062 5088 3338 5212
rect 3462 5088 3738 5212
rect 3862 5088 4138 5212
rect 4262 5088 4538 5212
rect 4662 5088 4938 5212
rect 5062 5088 5338 5212
rect 5462 5088 5738 5212
rect 5862 5088 6138 5212
rect 6262 5088 6538 5212
rect 6662 5088 6938 5212
rect 7062 5088 7338 5212
rect 7462 5088 7738 5212
rect 7862 5088 8138 5212
rect 8262 5088 8538 5212
rect 8662 5088 8938 5212
rect 9062 5088 9338 5212
rect 9462 5088 9738 5212
rect 9862 5088 10138 5212
rect 10262 5088 10538 5212
rect 10662 5088 10938 5212
rect 11062 5088 11338 5212
rect 11462 5088 11738 5212
rect 11862 5088 12138 5212
rect 12262 5088 12538 5212
rect 12662 5088 12938 5212
rect 13062 5088 13338 5212
rect 13462 5088 13738 5212
rect 13862 5088 14138 5212
rect 14262 5088 14538 5212
rect 14662 5088 14938 5212
rect 15062 5088 15220 5212
rect 780 4960 15220 5088
rect 15600 4960 15620 5340
rect 0 4940 16000 4960
rect 380 4560 400 4940
rect 780 4812 15220 4940
rect 780 4688 938 4812
rect 1062 4688 1338 4812
rect 1462 4688 1738 4812
rect 1862 4688 2138 4812
rect 2262 4688 2538 4812
rect 2662 4688 2938 4812
rect 3062 4688 3338 4812
rect 3462 4688 3738 4812
rect 3862 4688 4138 4812
rect 4262 4688 4538 4812
rect 4662 4688 4938 4812
rect 5062 4688 5338 4812
rect 5462 4688 5738 4812
rect 5862 4688 6138 4812
rect 6262 4688 6538 4812
rect 6662 4688 6938 4812
rect 7062 4688 7338 4812
rect 7462 4688 7738 4812
rect 7862 4688 8138 4812
rect 8262 4688 8538 4812
rect 8662 4688 8938 4812
rect 9062 4688 9338 4812
rect 9462 4688 9738 4812
rect 9862 4688 10138 4812
rect 10262 4688 10538 4812
rect 10662 4688 10938 4812
rect 11062 4688 11338 4812
rect 11462 4688 11738 4812
rect 11862 4688 12138 4812
rect 12262 4688 12538 4812
rect 12662 4688 12938 4812
rect 13062 4688 13338 4812
rect 13462 4688 13738 4812
rect 13862 4688 14138 4812
rect 14262 4688 14538 4812
rect 14662 4688 14938 4812
rect 15062 4688 15220 4812
rect 780 4560 15220 4688
rect 15600 4560 15620 4940
rect 0 4540 16000 4560
rect 380 4160 400 4540
rect 780 4412 15220 4540
rect 780 4288 938 4412
rect 1062 4288 1338 4412
rect 1462 4288 1738 4412
rect 1862 4288 2138 4412
rect 2262 4288 2538 4412
rect 2662 4288 2938 4412
rect 3062 4288 3338 4412
rect 3462 4288 3738 4412
rect 3862 4288 4138 4412
rect 4262 4288 4538 4412
rect 4662 4288 4938 4412
rect 5062 4288 5338 4412
rect 5462 4288 5738 4412
rect 5862 4288 6138 4412
rect 6262 4288 6538 4412
rect 6662 4288 6938 4412
rect 7062 4288 7338 4412
rect 7462 4288 7738 4412
rect 7862 4288 8138 4412
rect 8262 4288 8538 4412
rect 8662 4288 8938 4412
rect 9062 4288 9338 4412
rect 9462 4288 9738 4412
rect 9862 4288 10138 4412
rect 10262 4288 10538 4412
rect 10662 4288 10938 4412
rect 11062 4288 11338 4412
rect 11462 4288 11738 4412
rect 11862 4288 12138 4412
rect 12262 4288 12538 4412
rect 12662 4288 12938 4412
rect 13062 4288 13338 4412
rect 13462 4288 13738 4412
rect 13862 4288 14138 4412
rect 14262 4288 14538 4412
rect 14662 4288 14938 4412
rect 15062 4288 15220 4412
rect 780 4160 15220 4288
rect 15600 4160 15620 4540
rect 0 4140 16000 4160
rect 380 3760 400 4140
rect 780 4012 15220 4140
rect 780 3888 938 4012
rect 1062 3888 1338 4012
rect 1462 3888 1738 4012
rect 1862 3888 2138 4012
rect 2262 3888 2538 4012
rect 2662 3888 2938 4012
rect 3062 3888 3338 4012
rect 3462 3888 3738 4012
rect 3862 3888 4138 4012
rect 4262 3888 4538 4012
rect 4662 3888 4938 4012
rect 5062 3888 5338 4012
rect 5462 3888 5738 4012
rect 5862 3888 6138 4012
rect 6262 3888 6538 4012
rect 6662 3888 6938 4012
rect 7062 3888 7338 4012
rect 7462 3888 7738 4012
rect 7862 3888 8138 4012
rect 8262 3888 8538 4012
rect 8662 3888 8938 4012
rect 9062 3888 9338 4012
rect 9462 3888 9738 4012
rect 9862 3888 10138 4012
rect 10262 3888 10538 4012
rect 10662 3888 10938 4012
rect 11062 3888 11338 4012
rect 11462 3888 11738 4012
rect 11862 3888 12138 4012
rect 12262 3888 12538 4012
rect 12662 3888 12938 4012
rect 13062 3888 13338 4012
rect 13462 3888 13738 4012
rect 13862 3888 14138 4012
rect 14262 3888 14538 4012
rect 14662 3888 14938 4012
rect 15062 3888 15220 4012
rect 780 3760 15220 3888
rect 15600 3760 15620 4140
rect 0 3740 16000 3760
rect 380 3360 400 3740
rect 780 3612 15220 3740
rect 780 3488 938 3612
rect 1062 3488 1338 3612
rect 1462 3488 1738 3612
rect 1862 3488 2138 3612
rect 2262 3488 2538 3612
rect 2662 3488 2938 3612
rect 3062 3488 3338 3612
rect 3462 3488 3738 3612
rect 3862 3488 4138 3612
rect 4262 3488 4538 3612
rect 4662 3488 4938 3612
rect 5062 3488 5338 3612
rect 5462 3488 5738 3612
rect 5862 3488 6138 3612
rect 6262 3488 6538 3612
rect 6662 3488 6938 3612
rect 7062 3488 7338 3612
rect 7462 3488 7738 3612
rect 7862 3488 8138 3612
rect 8262 3488 8538 3612
rect 8662 3488 8938 3612
rect 9062 3488 9338 3612
rect 9462 3488 9738 3612
rect 9862 3488 10138 3612
rect 10262 3488 10538 3612
rect 10662 3488 10938 3612
rect 11062 3488 11338 3612
rect 11462 3488 11738 3612
rect 11862 3488 12138 3612
rect 12262 3488 12538 3612
rect 12662 3488 12938 3612
rect 13062 3488 13338 3612
rect 13462 3488 13738 3612
rect 13862 3488 14138 3612
rect 14262 3488 14538 3612
rect 14662 3488 14938 3612
rect 15062 3488 15220 3612
rect 780 3360 15220 3488
rect 15600 3360 15620 3740
rect 0 3340 16000 3360
rect 380 2960 400 3340
rect 780 3212 15220 3340
rect 780 3088 938 3212
rect 1062 3088 1338 3212
rect 1462 3088 1738 3212
rect 1862 3088 2138 3212
rect 2262 3088 2538 3212
rect 2662 3088 2938 3212
rect 3062 3088 3338 3212
rect 3462 3088 3738 3212
rect 3862 3088 4138 3212
rect 4262 3088 4538 3212
rect 4662 3088 4938 3212
rect 5062 3088 5338 3212
rect 5462 3088 5738 3212
rect 5862 3088 6138 3212
rect 6262 3088 6538 3212
rect 6662 3088 6938 3212
rect 7062 3088 7338 3212
rect 7462 3088 7738 3212
rect 7862 3088 8138 3212
rect 8262 3088 8538 3212
rect 8662 3088 8938 3212
rect 9062 3088 9338 3212
rect 9462 3088 9738 3212
rect 9862 3088 10138 3212
rect 10262 3088 10538 3212
rect 10662 3088 10938 3212
rect 11062 3088 11338 3212
rect 11462 3088 11738 3212
rect 11862 3088 12138 3212
rect 12262 3088 12538 3212
rect 12662 3088 12938 3212
rect 13062 3088 13338 3212
rect 13462 3088 13738 3212
rect 13862 3088 14138 3212
rect 14262 3088 14538 3212
rect 14662 3088 14938 3212
rect 15062 3088 15220 3212
rect 780 2960 15220 3088
rect 15600 2960 15620 3340
rect 0 2940 16000 2960
rect 380 2560 400 2940
rect 780 2812 15220 2940
rect 780 2688 938 2812
rect 1062 2688 1338 2812
rect 1462 2688 1738 2812
rect 1862 2688 2138 2812
rect 2262 2688 2538 2812
rect 2662 2688 2938 2812
rect 3062 2688 3338 2812
rect 3462 2688 3738 2812
rect 3862 2688 4138 2812
rect 4262 2688 4538 2812
rect 4662 2688 4938 2812
rect 5062 2688 5338 2812
rect 5462 2688 5738 2812
rect 5862 2688 6138 2812
rect 6262 2688 6538 2812
rect 6662 2688 6938 2812
rect 7062 2688 7338 2812
rect 7462 2688 7738 2812
rect 7862 2688 8138 2812
rect 8262 2688 8538 2812
rect 8662 2688 8938 2812
rect 9062 2688 9338 2812
rect 9462 2688 9738 2812
rect 9862 2688 10138 2812
rect 10262 2688 10538 2812
rect 10662 2688 10938 2812
rect 11062 2688 11338 2812
rect 11462 2688 11738 2812
rect 11862 2688 12138 2812
rect 12262 2688 12538 2812
rect 12662 2688 12938 2812
rect 13062 2688 13338 2812
rect 13462 2688 13738 2812
rect 13862 2688 14138 2812
rect 14262 2688 14538 2812
rect 14662 2688 14938 2812
rect 15062 2688 15220 2812
rect 780 2560 15220 2688
rect 15600 2560 15620 2940
rect 0 2540 16000 2560
rect 380 2160 400 2540
rect 780 2412 15220 2540
rect 780 2288 938 2412
rect 1062 2288 1338 2412
rect 1462 2288 1738 2412
rect 1862 2288 2138 2412
rect 2262 2288 2538 2412
rect 2662 2288 2938 2412
rect 3062 2288 3338 2412
rect 3462 2288 3738 2412
rect 3862 2288 4138 2412
rect 4262 2288 4538 2412
rect 4662 2288 4938 2412
rect 5062 2288 5338 2412
rect 5462 2288 5738 2412
rect 5862 2288 6138 2412
rect 6262 2288 6538 2412
rect 6662 2288 6938 2412
rect 7062 2288 7338 2412
rect 7462 2288 7738 2412
rect 7862 2288 8138 2412
rect 8262 2288 8538 2412
rect 8662 2288 8938 2412
rect 9062 2288 9338 2412
rect 9462 2288 9738 2412
rect 9862 2288 10138 2412
rect 10262 2288 10538 2412
rect 10662 2288 10938 2412
rect 11062 2288 11338 2412
rect 11462 2288 11738 2412
rect 11862 2288 12138 2412
rect 12262 2288 12538 2412
rect 12662 2288 12938 2412
rect 13062 2288 13338 2412
rect 13462 2288 13738 2412
rect 13862 2288 14138 2412
rect 14262 2288 14538 2412
rect 14662 2288 14938 2412
rect 15062 2288 15220 2412
rect 780 2160 15220 2288
rect 15600 2160 15620 2540
rect 0 2140 16000 2160
rect 380 1760 400 2140
rect 780 2012 15220 2140
rect 780 1888 938 2012
rect 1062 1888 1338 2012
rect 1462 1888 1738 2012
rect 1862 1888 2138 2012
rect 2262 1888 2538 2012
rect 2662 1888 2938 2012
rect 3062 1888 3338 2012
rect 3462 1888 3738 2012
rect 3862 1888 4138 2012
rect 4262 1888 4538 2012
rect 4662 1888 4938 2012
rect 5062 1888 5338 2012
rect 5462 1888 5738 2012
rect 5862 1888 6138 2012
rect 6262 1888 6538 2012
rect 6662 1888 6938 2012
rect 7062 1888 7338 2012
rect 7462 1888 7738 2012
rect 7862 1888 8138 2012
rect 8262 1888 8538 2012
rect 8662 1888 8938 2012
rect 9062 1888 9338 2012
rect 9462 1888 9738 2012
rect 9862 1888 10138 2012
rect 10262 1888 10538 2012
rect 10662 1888 10938 2012
rect 11062 1888 11338 2012
rect 11462 1888 11738 2012
rect 11862 1888 12138 2012
rect 12262 1888 12538 2012
rect 12662 1888 12938 2012
rect 13062 1888 13338 2012
rect 13462 1888 13738 2012
rect 13862 1888 14138 2012
rect 14262 1888 14538 2012
rect 14662 1888 14938 2012
rect 15062 1888 15220 2012
rect 780 1760 15220 1888
rect 15600 1760 15620 2140
rect 0 1400 16000 1760
rect 1000 490 15000 600
rect 1000 110 1010 490
rect 1390 110 1410 490
rect 1790 110 1810 490
rect 2190 110 2210 490
rect 2590 110 2610 490
rect 2990 110 3010 490
rect 3390 110 3410 490
rect 3790 110 3810 490
rect 4190 110 4210 490
rect 4590 110 4610 490
rect 4990 110 5010 490
rect 5390 110 5410 490
rect 5790 110 5810 490
rect 6190 110 6210 490
rect 6590 110 6610 490
rect 6990 110 7010 490
rect 7390 110 7410 490
rect 7790 110 7810 490
rect 8190 110 8210 490
rect 8590 110 8610 490
rect 8990 110 9010 490
rect 9390 110 9410 490
rect 9790 110 9810 490
rect 10190 110 10210 490
rect 10590 110 10610 490
rect 10990 110 11010 490
rect 11390 110 11410 490
rect 11790 110 11810 490
rect 12190 110 12210 490
rect 12590 110 12610 490
rect 12990 110 13010 490
rect 13390 110 13410 490
rect 13790 110 13810 490
rect 14190 110 14210 490
rect 14590 110 14610 490
rect 14990 110 15000 490
rect 1000 0 15000 110
<< via6 >>
rect 410 26138 538 26190
rect 538 26138 662 26190
rect 662 26138 790 26190
rect 410 25862 790 26138
rect 410 25810 538 25862
rect 538 25810 662 25862
rect 662 25810 790 25862
rect 810 26138 938 26190
rect 938 26138 1062 26190
rect 1062 26138 1190 26190
rect 810 25862 1190 26138
rect 810 25810 938 25862
rect 938 25810 1062 25862
rect 1062 25810 1190 25862
rect 1210 26138 1338 26190
rect 1338 26138 1462 26190
rect 1462 26138 1590 26190
rect 1210 25862 1590 26138
rect 1210 25810 1338 25862
rect 1338 25810 1462 25862
rect 1462 25810 1590 25862
rect 1610 26138 1738 26190
rect 1738 26138 1862 26190
rect 1862 26138 1990 26190
rect 1610 25862 1990 26138
rect 1610 25810 1738 25862
rect 1738 25810 1862 25862
rect 1862 25810 1990 25862
rect 2010 26138 2138 26190
rect 2138 26138 2262 26190
rect 2262 26138 2390 26190
rect 2010 25862 2390 26138
rect 2010 25810 2138 25862
rect 2138 25810 2262 25862
rect 2262 25810 2390 25862
rect 2410 26138 2538 26190
rect 2538 26138 2662 26190
rect 2662 26138 2790 26190
rect 2410 25862 2790 26138
rect 2410 25810 2538 25862
rect 2538 25810 2662 25862
rect 2662 25810 2790 25862
rect 2810 26138 2938 26190
rect 2938 26138 3062 26190
rect 3062 26138 3190 26190
rect 2810 25862 3190 26138
rect 2810 25810 2938 25862
rect 2938 25810 3062 25862
rect 3062 25810 3190 25862
rect 3210 26138 3338 26190
rect 3338 26138 3462 26190
rect 3462 26138 3590 26190
rect 3210 25862 3590 26138
rect 3210 25810 3338 25862
rect 3338 25810 3462 25862
rect 3462 25810 3590 25862
rect 3610 26138 3738 26190
rect 3738 26138 3862 26190
rect 3862 26138 3990 26190
rect 3610 25862 3990 26138
rect 3610 25810 3738 25862
rect 3738 25810 3862 25862
rect 3862 25810 3990 25862
rect 4010 26138 4138 26190
rect 4138 26138 4262 26190
rect 4262 26138 4390 26190
rect 4010 25862 4390 26138
rect 4010 25810 4138 25862
rect 4138 25810 4262 25862
rect 4262 25810 4390 25862
rect 4410 26138 4538 26190
rect 4538 26138 4662 26190
rect 4662 26138 4790 26190
rect 4410 25862 4790 26138
rect 4410 25810 4538 25862
rect 4538 25810 4662 25862
rect 4662 25810 4790 25862
rect 4810 26138 4938 26190
rect 4938 26138 5062 26190
rect 5062 26138 5190 26190
rect 4810 25862 5190 26138
rect 4810 25810 4938 25862
rect 4938 25810 5062 25862
rect 5062 25810 5190 25862
rect 5210 26138 5338 26190
rect 5338 26138 5462 26190
rect 5462 26138 5590 26190
rect 5210 25862 5590 26138
rect 5210 25810 5338 25862
rect 5338 25810 5462 25862
rect 5462 25810 5590 25862
rect 5610 26138 5738 26190
rect 5738 26138 5862 26190
rect 5862 26138 5990 26190
rect 5610 25862 5990 26138
rect 5610 25810 5738 25862
rect 5738 25810 5862 25862
rect 5862 25810 5990 25862
rect 6010 26138 6138 26190
rect 6138 26138 6262 26190
rect 6262 26138 6390 26190
rect 6010 25862 6390 26138
rect 6010 25810 6138 25862
rect 6138 25810 6262 25862
rect 6262 25810 6390 25862
rect 6410 26138 6538 26190
rect 6538 26138 6662 26190
rect 6662 26138 6790 26190
rect 6410 25862 6790 26138
rect 6410 25810 6538 25862
rect 6538 25810 6662 25862
rect 6662 25810 6790 25862
rect 6810 26138 6938 26190
rect 6938 26138 7062 26190
rect 7062 26138 7190 26190
rect 6810 25862 7190 26138
rect 6810 25810 6938 25862
rect 6938 25810 7062 25862
rect 7062 25810 7190 25862
rect 7210 26138 7338 26190
rect 7338 26138 7462 26190
rect 7462 26138 7590 26190
rect 7210 25862 7590 26138
rect 7210 25810 7338 25862
rect 7338 25810 7462 25862
rect 7462 25810 7590 25862
rect 7610 26138 7738 26190
rect 7738 26138 7862 26190
rect 7862 26138 7990 26190
rect 7610 25862 7990 26138
rect 7610 25810 7738 25862
rect 7738 25810 7862 25862
rect 7862 25810 7990 25862
rect 8010 26138 8138 26190
rect 8138 26138 8262 26190
rect 8262 26138 8390 26190
rect 8010 25862 8390 26138
rect 8010 25810 8138 25862
rect 8138 25810 8262 25862
rect 8262 25810 8390 25862
rect 8410 26138 8538 26190
rect 8538 26138 8662 26190
rect 8662 26138 8790 26190
rect 8410 25862 8790 26138
rect 8410 25810 8538 25862
rect 8538 25810 8662 25862
rect 8662 25810 8790 25862
rect 8810 26138 8938 26190
rect 8938 26138 9062 26190
rect 9062 26138 9190 26190
rect 8810 25862 9190 26138
rect 8810 25810 8938 25862
rect 8938 25810 9062 25862
rect 9062 25810 9190 25862
rect 9210 26138 9338 26190
rect 9338 26138 9462 26190
rect 9462 26138 9590 26190
rect 9210 25862 9590 26138
rect 9210 25810 9338 25862
rect 9338 25810 9462 25862
rect 9462 25810 9590 25862
rect 9610 26138 9738 26190
rect 9738 26138 9862 26190
rect 9862 26138 9990 26190
rect 9610 25862 9990 26138
rect 9610 25810 9738 25862
rect 9738 25810 9862 25862
rect 9862 25810 9990 25862
rect 10010 26138 10138 26190
rect 10138 26138 10262 26190
rect 10262 26138 10390 26190
rect 10010 25862 10390 26138
rect 10010 25810 10138 25862
rect 10138 25810 10262 25862
rect 10262 25810 10390 25862
rect 10410 26138 10538 26190
rect 10538 26138 10662 26190
rect 10662 26138 10790 26190
rect 10410 25862 10790 26138
rect 10410 25810 10538 25862
rect 10538 25810 10662 25862
rect 10662 25810 10790 25862
rect 10810 26138 10938 26190
rect 10938 26138 11062 26190
rect 11062 26138 11190 26190
rect 10810 25862 11190 26138
rect 10810 25810 10938 25862
rect 10938 25810 11062 25862
rect 11062 25810 11190 25862
rect 11210 26138 11338 26190
rect 11338 26138 11462 26190
rect 11462 26138 11590 26190
rect 11210 25862 11590 26138
rect 11210 25810 11338 25862
rect 11338 25810 11462 25862
rect 11462 25810 11590 25862
rect 11610 26138 11738 26190
rect 11738 26138 11862 26190
rect 11862 26138 11990 26190
rect 11610 25862 11990 26138
rect 11610 25810 11738 25862
rect 11738 25810 11862 25862
rect 11862 25810 11990 25862
rect 12010 26138 12138 26190
rect 12138 26138 12262 26190
rect 12262 26138 12390 26190
rect 12010 25862 12390 26138
rect 12010 25810 12138 25862
rect 12138 25810 12262 25862
rect 12262 25810 12390 25862
rect 12410 26138 12538 26190
rect 12538 26138 12662 26190
rect 12662 26138 12790 26190
rect 12410 25862 12790 26138
rect 12410 25810 12538 25862
rect 12538 25810 12662 25862
rect 12662 25810 12790 25862
rect 12810 26138 12938 26190
rect 12938 26138 13062 26190
rect 13062 26138 13190 26190
rect 12810 25862 13190 26138
rect 12810 25810 12938 25862
rect 12938 25810 13062 25862
rect 13062 25810 13190 25862
rect 13210 26138 13338 26190
rect 13338 26138 13462 26190
rect 13462 26138 13590 26190
rect 13210 25862 13590 26138
rect 13210 25810 13338 25862
rect 13338 25810 13462 25862
rect 13462 25810 13590 25862
rect 13610 26138 13738 26190
rect 13738 26138 13862 26190
rect 13862 26138 13990 26190
rect 13610 25862 13990 26138
rect 13610 25810 13738 25862
rect 13738 25810 13862 25862
rect 13862 25810 13990 25862
rect 14010 26138 14138 26190
rect 14138 26138 14262 26190
rect 14262 26138 14390 26190
rect 14010 25862 14390 26138
rect 14010 25810 14138 25862
rect 14138 25810 14262 25862
rect 14262 25810 14390 25862
rect 14410 26138 14538 26190
rect 14538 26138 14662 26190
rect 14662 26138 14790 26190
rect 14410 25862 14790 26138
rect 14410 25810 14538 25862
rect 14538 25810 14662 25862
rect 14662 25810 14790 25862
rect 14810 26138 14938 26190
rect 14938 26138 15062 26190
rect 15062 26138 15190 26190
rect 14810 25862 15190 26138
rect 14810 25810 14938 25862
rect 14938 25810 15062 25862
rect 15062 25810 15190 25862
rect 15210 26138 15338 26190
rect 15338 26138 15462 26190
rect 15462 26138 15590 26190
rect 15210 25862 15590 26138
rect 15210 25810 15338 25862
rect 15338 25810 15462 25862
rect 15462 25810 15590 25862
rect 410 23188 538 23240
rect 538 23188 662 23240
rect 662 23188 790 23240
rect 410 22912 790 23188
rect 410 22860 538 22912
rect 538 22860 662 22912
rect 662 22860 790 22912
rect 810 23188 938 23240
rect 938 23188 1062 23240
rect 1062 23188 1190 23240
rect 810 22912 1190 23188
rect 810 22860 938 22912
rect 938 22860 1062 22912
rect 1062 22860 1190 22912
rect 1210 23188 1338 23240
rect 1338 23188 1462 23240
rect 1462 23188 1590 23240
rect 1210 22912 1590 23188
rect 1210 22860 1338 22912
rect 1338 22860 1462 22912
rect 1462 22860 1590 22912
rect 1610 23188 1738 23240
rect 1738 23188 1862 23240
rect 1862 23188 1990 23240
rect 1610 22912 1990 23188
rect 1610 22860 1738 22912
rect 1738 22860 1862 22912
rect 1862 22860 1990 22912
rect 2010 23188 2138 23240
rect 2138 23188 2262 23240
rect 2262 23188 2390 23240
rect 2010 22912 2390 23188
rect 2010 22860 2138 22912
rect 2138 22860 2262 22912
rect 2262 22860 2390 22912
rect 2410 23188 2538 23240
rect 2538 23188 2662 23240
rect 2662 23188 2790 23240
rect 2410 22912 2790 23188
rect 2410 22860 2538 22912
rect 2538 22860 2662 22912
rect 2662 22860 2790 22912
rect 2810 23188 2938 23240
rect 2938 23188 3062 23240
rect 3062 23188 3190 23240
rect 2810 22912 3190 23188
rect 2810 22860 2938 22912
rect 2938 22860 3062 22912
rect 3062 22860 3190 22912
rect 3210 23188 3338 23240
rect 3338 23188 3462 23240
rect 3462 23188 3590 23240
rect 3210 22912 3590 23188
rect 3210 22860 3338 22912
rect 3338 22860 3462 22912
rect 3462 22860 3590 22912
rect 3610 23188 3738 23240
rect 3738 23188 3862 23240
rect 3862 23188 3990 23240
rect 3610 22912 3990 23188
rect 3610 22860 3738 22912
rect 3738 22860 3862 22912
rect 3862 22860 3990 22912
rect 4010 23188 4138 23240
rect 4138 23188 4262 23240
rect 4262 23188 4390 23240
rect 4010 22912 4390 23188
rect 4010 22860 4138 22912
rect 4138 22860 4262 22912
rect 4262 22860 4390 22912
rect 4410 23188 4538 23240
rect 4538 23188 4662 23240
rect 4662 23188 4790 23240
rect 4410 22912 4790 23188
rect 4410 22860 4538 22912
rect 4538 22860 4662 22912
rect 4662 22860 4790 22912
rect 4810 23188 4938 23240
rect 4938 23188 5062 23240
rect 5062 23188 5190 23240
rect 4810 22912 5190 23188
rect 4810 22860 4938 22912
rect 4938 22860 5062 22912
rect 5062 22860 5190 22912
rect 5210 23188 5338 23240
rect 5338 23188 5462 23240
rect 5462 23188 5590 23240
rect 5210 22912 5590 23188
rect 5210 22860 5338 22912
rect 5338 22860 5462 22912
rect 5462 22860 5590 22912
rect 5610 23188 5738 23240
rect 5738 23188 5862 23240
rect 5862 23188 5990 23240
rect 5610 22912 5990 23188
rect 5610 22860 5738 22912
rect 5738 22860 5862 22912
rect 5862 22860 5990 22912
rect 6010 23188 6138 23240
rect 6138 23188 6262 23240
rect 6262 23188 6390 23240
rect 6010 22912 6390 23188
rect 6010 22860 6138 22912
rect 6138 22860 6262 22912
rect 6262 22860 6390 22912
rect 6410 23188 6538 23240
rect 6538 23188 6662 23240
rect 6662 23188 6790 23240
rect 6410 22912 6790 23188
rect 6410 22860 6538 22912
rect 6538 22860 6662 22912
rect 6662 22860 6790 22912
rect 6810 23188 6938 23240
rect 6938 23188 7062 23240
rect 7062 23188 7190 23240
rect 6810 22912 7190 23188
rect 6810 22860 6938 22912
rect 6938 22860 7062 22912
rect 7062 22860 7190 22912
rect 7210 23188 7338 23240
rect 7338 23188 7462 23240
rect 7462 23188 7590 23240
rect 7210 22912 7590 23188
rect 7210 22860 7338 22912
rect 7338 22860 7462 22912
rect 7462 22860 7590 22912
rect 7610 23188 7738 23240
rect 7738 23188 7862 23240
rect 7862 23188 7990 23240
rect 7610 22912 7990 23188
rect 7610 22860 7738 22912
rect 7738 22860 7862 22912
rect 7862 22860 7990 22912
rect 8010 23188 8138 23240
rect 8138 23188 8262 23240
rect 8262 23188 8390 23240
rect 8010 22912 8390 23188
rect 8010 22860 8138 22912
rect 8138 22860 8262 22912
rect 8262 22860 8390 22912
rect 8410 23188 8538 23240
rect 8538 23188 8662 23240
rect 8662 23188 8790 23240
rect 8410 22912 8790 23188
rect 8410 22860 8538 22912
rect 8538 22860 8662 22912
rect 8662 22860 8790 22912
rect 8810 23188 8938 23240
rect 8938 23188 9062 23240
rect 9062 23188 9190 23240
rect 8810 22912 9190 23188
rect 8810 22860 8938 22912
rect 8938 22860 9062 22912
rect 9062 22860 9190 22912
rect 9210 23188 9338 23240
rect 9338 23188 9462 23240
rect 9462 23188 9590 23240
rect 9210 22912 9590 23188
rect 9210 22860 9338 22912
rect 9338 22860 9462 22912
rect 9462 22860 9590 22912
rect 9610 23188 9738 23240
rect 9738 23188 9862 23240
rect 9862 23188 9990 23240
rect 9610 22912 9990 23188
rect 9610 22860 9738 22912
rect 9738 22860 9862 22912
rect 9862 22860 9990 22912
rect 10010 23188 10138 23240
rect 10138 23188 10262 23240
rect 10262 23188 10390 23240
rect 10010 22912 10390 23188
rect 10010 22860 10138 22912
rect 10138 22860 10262 22912
rect 10262 22860 10390 22912
rect 10410 23188 10538 23240
rect 10538 23188 10662 23240
rect 10662 23188 10790 23240
rect 10410 22912 10790 23188
rect 10410 22860 10538 22912
rect 10538 22860 10662 22912
rect 10662 22860 10790 22912
rect 10810 23188 10938 23240
rect 10938 23188 11062 23240
rect 11062 23188 11190 23240
rect 10810 22912 11190 23188
rect 10810 22860 10938 22912
rect 10938 22860 11062 22912
rect 11062 22860 11190 22912
rect 11210 23188 11338 23240
rect 11338 23188 11462 23240
rect 11462 23188 11590 23240
rect 11210 22912 11590 23188
rect 11210 22860 11338 22912
rect 11338 22860 11462 22912
rect 11462 22860 11590 22912
rect 11610 23188 11738 23240
rect 11738 23188 11862 23240
rect 11862 23188 11990 23240
rect 11610 22912 11990 23188
rect 11610 22860 11738 22912
rect 11738 22860 11862 22912
rect 11862 22860 11990 22912
rect 12010 23188 12138 23240
rect 12138 23188 12262 23240
rect 12262 23188 12390 23240
rect 12010 22912 12390 23188
rect 12010 22860 12138 22912
rect 12138 22860 12262 22912
rect 12262 22860 12390 22912
rect 12410 23188 12538 23240
rect 12538 23188 12662 23240
rect 12662 23188 12790 23240
rect 12410 22912 12790 23188
rect 12410 22860 12538 22912
rect 12538 22860 12662 22912
rect 12662 22860 12790 22912
rect 12810 23188 12938 23240
rect 12938 23188 13062 23240
rect 13062 23188 13190 23240
rect 12810 22912 13190 23188
rect 12810 22860 12938 22912
rect 12938 22860 13062 22912
rect 13062 22860 13190 22912
rect 13210 23188 13338 23240
rect 13338 23188 13462 23240
rect 13462 23188 13590 23240
rect 13210 22912 13590 23188
rect 13210 22860 13338 22912
rect 13338 22860 13462 22912
rect 13462 22860 13590 22912
rect 13610 23188 13738 23240
rect 13738 23188 13862 23240
rect 13862 23188 13990 23240
rect 13610 22912 13990 23188
rect 13610 22860 13738 22912
rect 13738 22860 13862 22912
rect 13862 22860 13990 22912
rect 14010 23188 14138 23240
rect 14138 23188 14262 23240
rect 14262 23188 14390 23240
rect 14010 22912 14390 23188
rect 14010 22860 14138 22912
rect 14138 22860 14262 22912
rect 14262 22860 14390 22912
rect 14410 23188 14538 23240
rect 14538 23188 14662 23240
rect 14662 23188 14790 23240
rect 14410 22912 14790 23188
rect 14410 22860 14538 22912
rect 14538 22860 14662 22912
rect 14662 22860 14790 22912
rect 14810 23188 14938 23240
rect 14938 23188 15062 23240
rect 15062 23188 15190 23240
rect 14810 22912 15190 23188
rect 14810 22860 14938 22912
rect 14938 22860 15062 22912
rect 15062 22860 15190 22912
rect 15210 23188 15338 23240
rect 15338 23188 15462 23240
rect 15462 23188 15590 23240
rect 15210 22912 15590 23188
rect 15210 22860 15338 22912
rect 15338 22860 15462 22912
rect 15462 22860 15590 22912
rect 410 22788 538 22840
rect 538 22788 662 22840
rect 662 22788 790 22840
rect 410 22512 790 22788
rect 410 22460 538 22512
rect 538 22460 662 22512
rect 662 22460 790 22512
rect 810 22788 938 22840
rect 938 22788 1062 22840
rect 1062 22788 1190 22840
rect 810 22512 1190 22788
rect 810 22460 938 22512
rect 938 22460 1062 22512
rect 1062 22460 1190 22512
rect 1210 22788 1338 22840
rect 1338 22788 1462 22840
rect 1462 22788 1590 22840
rect 1210 22512 1590 22788
rect 1210 22460 1338 22512
rect 1338 22460 1462 22512
rect 1462 22460 1590 22512
rect 1610 22788 1738 22840
rect 1738 22788 1862 22840
rect 1862 22788 1990 22840
rect 1610 22512 1990 22788
rect 1610 22460 1738 22512
rect 1738 22460 1862 22512
rect 1862 22460 1990 22512
rect 2010 22788 2138 22840
rect 2138 22788 2262 22840
rect 2262 22788 2390 22840
rect 2010 22512 2390 22788
rect 2010 22460 2138 22512
rect 2138 22460 2262 22512
rect 2262 22460 2390 22512
rect 2410 22788 2538 22840
rect 2538 22788 2662 22840
rect 2662 22788 2790 22840
rect 2410 22512 2790 22788
rect 2410 22460 2538 22512
rect 2538 22460 2662 22512
rect 2662 22460 2790 22512
rect 2810 22788 2938 22840
rect 2938 22788 3062 22840
rect 3062 22788 3190 22840
rect 2810 22512 3190 22788
rect 2810 22460 2938 22512
rect 2938 22460 3062 22512
rect 3062 22460 3190 22512
rect 3210 22788 3338 22840
rect 3338 22788 3462 22840
rect 3462 22788 3590 22840
rect 3210 22512 3590 22788
rect 3210 22460 3338 22512
rect 3338 22460 3462 22512
rect 3462 22460 3590 22512
rect 3610 22788 3738 22840
rect 3738 22788 3862 22840
rect 3862 22788 3990 22840
rect 3610 22512 3990 22788
rect 3610 22460 3738 22512
rect 3738 22460 3862 22512
rect 3862 22460 3990 22512
rect 4010 22788 4138 22840
rect 4138 22788 4262 22840
rect 4262 22788 4390 22840
rect 4010 22512 4390 22788
rect 4010 22460 4138 22512
rect 4138 22460 4262 22512
rect 4262 22460 4390 22512
rect 4410 22788 4538 22840
rect 4538 22788 4662 22840
rect 4662 22788 4790 22840
rect 4410 22512 4790 22788
rect 4410 22460 4538 22512
rect 4538 22460 4662 22512
rect 4662 22460 4790 22512
rect 4810 22788 4938 22840
rect 4938 22788 5062 22840
rect 5062 22788 5190 22840
rect 4810 22512 5190 22788
rect 4810 22460 4938 22512
rect 4938 22460 5062 22512
rect 5062 22460 5190 22512
rect 5210 22788 5338 22840
rect 5338 22788 5462 22840
rect 5462 22788 5590 22840
rect 5210 22512 5590 22788
rect 5210 22460 5338 22512
rect 5338 22460 5462 22512
rect 5462 22460 5590 22512
rect 5610 22788 5738 22840
rect 5738 22788 5862 22840
rect 5862 22788 5990 22840
rect 5610 22512 5990 22788
rect 5610 22460 5738 22512
rect 5738 22460 5862 22512
rect 5862 22460 5990 22512
rect 6010 22788 6138 22840
rect 6138 22788 6262 22840
rect 6262 22788 6390 22840
rect 6010 22512 6390 22788
rect 6010 22460 6138 22512
rect 6138 22460 6262 22512
rect 6262 22460 6390 22512
rect 6410 22788 6538 22840
rect 6538 22788 6662 22840
rect 6662 22788 6790 22840
rect 6410 22512 6790 22788
rect 6410 22460 6538 22512
rect 6538 22460 6662 22512
rect 6662 22460 6790 22512
rect 6810 22788 6938 22840
rect 6938 22788 7062 22840
rect 7062 22788 7190 22840
rect 6810 22512 7190 22788
rect 6810 22460 6938 22512
rect 6938 22460 7062 22512
rect 7062 22460 7190 22512
rect 7210 22788 7338 22840
rect 7338 22788 7462 22840
rect 7462 22788 7590 22840
rect 7210 22512 7590 22788
rect 7210 22460 7338 22512
rect 7338 22460 7462 22512
rect 7462 22460 7590 22512
rect 7610 22788 7738 22840
rect 7738 22788 7862 22840
rect 7862 22788 7990 22840
rect 7610 22512 7990 22788
rect 7610 22460 7738 22512
rect 7738 22460 7862 22512
rect 7862 22460 7990 22512
rect 8010 22788 8138 22840
rect 8138 22788 8262 22840
rect 8262 22788 8390 22840
rect 8010 22512 8390 22788
rect 8010 22460 8138 22512
rect 8138 22460 8262 22512
rect 8262 22460 8390 22512
rect 8410 22788 8538 22840
rect 8538 22788 8662 22840
rect 8662 22788 8790 22840
rect 8410 22512 8790 22788
rect 8410 22460 8538 22512
rect 8538 22460 8662 22512
rect 8662 22460 8790 22512
rect 8810 22788 8938 22840
rect 8938 22788 9062 22840
rect 9062 22788 9190 22840
rect 8810 22512 9190 22788
rect 8810 22460 8938 22512
rect 8938 22460 9062 22512
rect 9062 22460 9190 22512
rect 9210 22788 9338 22840
rect 9338 22788 9462 22840
rect 9462 22788 9590 22840
rect 9210 22512 9590 22788
rect 9210 22460 9338 22512
rect 9338 22460 9462 22512
rect 9462 22460 9590 22512
rect 9610 22788 9738 22840
rect 9738 22788 9862 22840
rect 9862 22788 9990 22840
rect 9610 22512 9990 22788
rect 9610 22460 9738 22512
rect 9738 22460 9862 22512
rect 9862 22460 9990 22512
rect 10010 22788 10138 22840
rect 10138 22788 10262 22840
rect 10262 22788 10390 22840
rect 10010 22512 10390 22788
rect 10010 22460 10138 22512
rect 10138 22460 10262 22512
rect 10262 22460 10390 22512
rect 10410 22788 10538 22840
rect 10538 22788 10662 22840
rect 10662 22788 10790 22840
rect 10410 22512 10790 22788
rect 10410 22460 10538 22512
rect 10538 22460 10662 22512
rect 10662 22460 10790 22512
rect 10810 22788 10938 22840
rect 10938 22788 11062 22840
rect 11062 22788 11190 22840
rect 10810 22512 11190 22788
rect 10810 22460 10938 22512
rect 10938 22460 11062 22512
rect 11062 22460 11190 22512
rect 11210 22788 11338 22840
rect 11338 22788 11462 22840
rect 11462 22788 11590 22840
rect 11210 22512 11590 22788
rect 11210 22460 11338 22512
rect 11338 22460 11462 22512
rect 11462 22460 11590 22512
rect 11610 22788 11738 22840
rect 11738 22788 11862 22840
rect 11862 22788 11990 22840
rect 11610 22512 11990 22788
rect 11610 22460 11738 22512
rect 11738 22460 11862 22512
rect 11862 22460 11990 22512
rect 12010 22788 12138 22840
rect 12138 22788 12262 22840
rect 12262 22788 12390 22840
rect 12010 22512 12390 22788
rect 12010 22460 12138 22512
rect 12138 22460 12262 22512
rect 12262 22460 12390 22512
rect 12410 22788 12538 22840
rect 12538 22788 12662 22840
rect 12662 22788 12790 22840
rect 12410 22512 12790 22788
rect 12410 22460 12538 22512
rect 12538 22460 12662 22512
rect 12662 22460 12790 22512
rect 12810 22788 12938 22840
rect 12938 22788 13062 22840
rect 13062 22788 13190 22840
rect 12810 22512 13190 22788
rect 12810 22460 12938 22512
rect 12938 22460 13062 22512
rect 13062 22460 13190 22512
rect 13210 22788 13338 22840
rect 13338 22788 13462 22840
rect 13462 22788 13590 22840
rect 13210 22512 13590 22788
rect 13210 22460 13338 22512
rect 13338 22460 13462 22512
rect 13462 22460 13590 22512
rect 13610 22788 13738 22840
rect 13738 22788 13862 22840
rect 13862 22788 13990 22840
rect 13610 22512 13990 22788
rect 13610 22460 13738 22512
rect 13738 22460 13862 22512
rect 13862 22460 13990 22512
rect 14010 22788 14138 22840
rect 14138 22788 14262 22840
rect 14262 22788 14390 22840
rect 14010 22512 14390 22788
rect 14010 22460 14138 22512
rect 14138 22460 14262 22512
rect 14262 22460 14390 22512
rect 14410 22788 14538 22840
rect 14538 22788 14662 22840
rect 14662 22788 14790 22840
rect 14410 22512 14790 22788
rect 14410 22460 14538 22512
rect 14538 22460 14662 22512
rect 14662 22460 14790 22512
rect 14810 22788 14938 22840
rect 14938 22788 15062 22840
rect 15062 22788 15190 22840
rect 14810 22512 15190 22788
rect 14810 22460 14938 22512
rect 14938 22460 15062 22512
rect 15062 22460 15190 22512
rect 15210 22788 15338 22840
rect 15338 22788 15462 22840
rect 15462 22788 15590 22840
rect 15210 22512 15590 22788
rect 15210 22460 15338 22512
rect 15338 22460 15462 22512
rect 15462 22460 15590 22512
rect 410 22388 538 22440
rect 538 22388 662 22440
rect 662 22388 790 22440
rect 410 22112 790 22388
rect 410 22060 538 22112
rect 538 22060 662 22112
rect 662 22060 790 22112
rect 810 22388 938 22440
rect 938 22388 1062 22440
rect 1062 22388 1190 22440
rect 810 22112 1190 22388
rect 810 22060 938 22112
rect 938 22060 1062 22112
rect 1062 22060 1190 22112
rect 1210 22388 1338 22440
rect 1338 22388 1462 22440
rect 1462 22388 1590 22440
rect 1210 22112 1590 22388
rect 1210 22060 1338 22112
rect 1338 22060 1462 22112
rect 1462 22060 1590 22112
rect 1610 22388 1738 22440
rect 1738 22388 1862 22440
rect 1862 22388 1990 22440
rect 1610 22112 1990 22388
rect 1610 22060 1738 22112
rect 1738 22060 1862 22112
rect 1862 22060 1990 22112
rect 2010 22388 2138 22440
rect 2138 22388 2262 22440
rect 2262 22388 2390 22440
rect 2010 22112 2390 22388
rect 2010 22060 2138 22112
rect 2138 22060 2262 22112
rect 2262 22060 2390 22112
rect 2410 22388 2538 22440
rect 2538 22388 2662 22440
rect 2662 22388 2790 22440
rect 2410 22112 2790 22388
rect 2410 22060 2538 22112
rect 2538 22060 2662 22112
rect 2662 22060 2790 22112
rect 2810 22388 2938 22440
rect 2938 22388 3062 22440
rect 3062 22388 3190 22440
rect 2810 22112 3190 22388
rect 2810 22060 2938 22112
rect 2938 22060 3062 22112
rect 3062 22060 3190 22112
rect 3210 22388 3338 22440
rect 3338 22388 3462 22440
rect 3462 22388 3590 22440
rect 3210 22112 3590 22388
rect 3210 22060 3338 22112
rect 3338 22060 3462 22112
rect 3462 22060 3590 22112
rect 3610 22388 3738 22440
rect 3738 22388 3862 22440
rect 3862 22388 3990 22440
rect 3610 22112 3990 22388
rect 3610 22060 3738 22112
rect 3738 22060 3862 22112
rect 3862 22060 3990 22112
rect 4010 22388 4138 22440
rect 4138 22388 4262 22440
rect 4262 22388 4390 22440
rect 4010 22112 4390 22388
rect 4010 22060 4138 22112
rect 4138 22060 4262 22112
rect 4262 22060 4390 22112
rect 4410 22388 4538 22440
rect 4538 22388 4662 22440
rect 4662 22388 4790 22440
rect 4410 22112 4790 22388
rect 4410 22060 4538 22112
rect 4538 22060 4662 22112
rect 4662 22060 4790 22112
rect 4810 22388 4938 22440
rect 4938 22388 5062 22440
rect 5062 22388 5190 22440
rect 4810 22112 5190 22388
rect 4810 22060 4938 22112
rect 4938 22060 5062 22112
rect 5062 22060 5190 22112
rect 5210 22388 5338 22440
rect 5338 22388 5462 22440
rect 5462 22388 5590 22440
rect 5210 22112 5590 22388
rect 5210 22060 5338 22112
rect 5338 22060 5462 22112
rect 5462 22060 5590 22112
rect 5610 22388 5738 22440
rect 5738 22388 5862 22440
rect 5862 22388 5990 22440
rect 5610 22112 5990 22388
rect 5610 22060 5738 22112
rect 5738 22060 5862 22112
rect 5862 22060 5990 22112
rect 6010 22388 6138 22440
rect 6138 22388 6262 22440
rect 6262 22388 6390 22440
rect 6010 22112 6390 22388
rect 6010 22060 6138 22112
rect 6138 22060 6262 22112
rect 6262 22060 6390 22112
rect 6410 22388 6538 22440
rect 6538 22388 6662 22440
rect 6662 22388 6790 22440
rect 6410 22112 6790 22388
rect 6410 22060 6538 22112
rect 6538 22060 6662 22112
rect 6662 22060 6790 22112
rect 6810 22388 6938 22440
rect 6938 22388 7062 22440
rect 7062 22388 7190 22440
rect 6810 22112 7190 22388
rect 6810 22060 6938 22112
rect 6938 22060 7062 22112
rect 7062 22060 7190 22112
rect 7210 22388 7338 22440
rect 7338 22388 7462 22440
rect 7462 22388 7590 22440
rect 7210 22112 7590 22388
rect 7210 22060 7338 22112
rect 7338 22060 7462 22112
rect 7462 22060 7590 22112
rect 7610 22388 7738 22440
rect 7738 22388 7862 22440
rect 7862 22388 7990 22440
rect 7610 22112 7990 22388
rect 7610 22060 7738 22112
rect 7738 22060 7862 22112
rect 7862 22060 7990 22112
rect 8010 22388 8138 22440
rect 8138 22388 8262 22440
rect 8262 22388 8390 22440
rect 8010 22112 8390 22388
rect 8010 22060 8138 22112
rect 8138 22060 8262 22112
rect 8262 22060 8390 22112
rect 8410 22388 8538 22440
rect 8538 22388 8662 22440
rect 8662 22388 8790 22440
rect 8410 22112 8790 22388
rect 8410 22060 8538 22112
rect 8538 22060 8662 22112
rect 8662 22060 8790 22112
rect 8810 22388 8938 22440
rect 8938 22388 9062 22440
rect 9062 22388 9190 22440
rect 8810 22112 9190 22388
rect 8810 22060 8938 22112
rect 8938 22060 9062 22112
rect 9062 22060 9190 22112
rect 9210 22388 9338 22440
rect 9338 22388 9462 22440
rect 9462 22388 9590 22440
rect 9210 22112 9590 22388
rect 9210 22060 9338 22112
rect 9338 22060 9462 22112
rect 9462 22060 9590 22112
rect 9610 22388 9738 22440
rect 9738 22388 9862 22440
rect 9862 22388 9990 22440
rect 9610 22112 9990 22388
rect 9610 22060 9738 22112
rect 9738 22060 9862 22112
rect 9862 22060 9990 22112
rect 10010 22388 10138 22440
rect 10138 22388 10262 22440
rect 10262 22388 10390 22440
rect 10010 22112 10390 22388
rect 10010 22060 10138 22112
rect 10138 22060 10262 22112
rect 10262 22060 10390 22112
rect 10410 22388 10538 22440
rect 10538 22388 10662 22440
rect 10662 22388 10790 22440
rect 10410 22112 10790 22388
rect 10410 22060 10538 22112
rect 10538 22060 10662 22112
rect 10662 22060 10790 22112
rect 10810 22388 10938 22440
rect 10938 22388 11062 22440
rect 11062 22388 11190 22440
rect 10810 22112 11190 22388
rect 10810 22060 10938 22112
rect 10938 22060 11062 22112
rect 11062 22060 11190 22112
rect 11210 22388 11338 22440
rect 11338 22388 11462 22440
rect 11462 22388 11590 22440
rect 11210 22112 11590 22388
rect 11210 22060 11338 22112
rect 11338 22060 11462 22112
rect 11462 22060 11590 22112
rect 11610 22388 11738 22440
rect 11738 22388 11862 22440
rect 11862 22388 11990 22440
rect 11610 22112 11990 22388
rect 11610 22060 11738 22112
rect 11738 22060 11862 22112
rect 11862 22060 11990 22112
rect 12010 22388 12138 22440
rect 12138 22388 12262 22440
rect 12262 22388 12390 22440
rect 12010 22112 12390 22388
rect 12010 22060 12138 22112
rect 12138 22060 12262 22112
rect 12262 22060 12390 22112
rect 12410 22388 12538 22440
rect 12538 22388 12662 22440
rect 12662 22388 12790 22440
rect 12410 22112 12790 22388
rect 12410 22060 12538 22112
rect 12538 22060 12662 22112
rect 12662 22060 12790 22112
rect 12810 22388 12938 22440
rect 12938 22388 13062 22440
rect 13062 22388 13190 22440
rect 12810 22112 13190 22388
rect 12810 22060 12938 22112
rect 12938 22060 13062 22112
rect 13062 22060 13190 22112
rect 13210 22388 13338 22440
rect 13338 22388 13462 22440
rect 13462 22388 13590 22440
rect 13210 22112 13590 22388
rect 13210 22060 13338 22112
rect 13338 22060 13462 22112
rect 13462 22060 13590 22112
rect 13610 22388 13738 22440
rect 13738 22388 13862 22440
rect 13862 22388 13990 22440
rect 13610 22112 13990 22388
rect 13610 22060 13738 22112
rect 13738 22060 13862 22112
rect 13862 22060 13990 22112
rect 14010 22388 14138 22440
rect 14138 22388 14262 22440
rect 14262 22388 14390 22440
rect 14010 22112 14390 22388
rect 14010 22060 14138 22112
rect 14138 22060 14262 22112
rect 14262 22060 14390 22112
rect 14410 22388 14538 22440
rect 14538 22388 14662 22440
rect 14662 22388 14790 22440
rect 14410 22112 14790 22388
rect 14410 22060 14538 22112
rect 14538 22060 14662 22112
rect 14662 22060 14790 22112
rect 14810 22388 14938 22440
rect 14938 22388 15062 22440
rect 15062 22388 15190 22440
rect 14810 22112 15190 22388
rect 14810 22060 14938 22112
rect 14938 22060 15062 22112
rect 15062 22060 15190 22112
rect 15210 22388 15338 22440
rect 15338 22388 15462 22440
rect 15462 22388 15590 22440
rect 15210 22112 15590 22388
rect 15210 22060 15338 22112
rect 15338 22060 15462 22112
rect 15462 22060 15590 22112
rect 410 21988 538 22040
rect 538 21988 662 22040
rect 662 21988 790 22040
rect 410 21712 790 21988
rect 410 21660 538 21712
rect 538 21660 662 21712
rect 662 21660 790 21712
rect 810 21988 938 22040
rect 938 21988 1062 22040
rect 1062 21988 1190 22040
rect 810 21712 1190 21988
rect 810 21660 938 21712
rect 938 21660 1062 21712
rect 1062 21660 1190 21712
rect 1210 21988 1338 22040
rect 1338 21988 1462 22040
rect 1462 21988 1590 22040
rect 1210 21712 1590 21988
rect 1210 21660 1338 21712
rect 1338 21660 1462 21712
rect 1462 21660 1590 21712
rect 1610 21988 1738 22040
rect 1738 21988 1862 22040
rect 1862 21988 1990 22040
rect 1610 21712 1990 21988
rect 1610 21660 1738 21712
rect 1738 21660 1862 21712
rect 1862 21660 1990 21712
rect 2010 21988 2138 22040
rect 2138 21988 2262 22040
rect 2262 21988 2390 22040
rect 2010 21712 2390 21988
rect 2010 21660 2138 21712
rect 2138 21660 2262 21712
rect 2262 21660 2390 21712
rect 2410 21988 2538 22040
rect 2538 21988 2662 22040
rect 2662 21988 2790 22040
rect 2410 21712 2790 21988
rect 2410 21660 2538 21712
rect 2538 21660 2662 21712
rect 2662 21660 2790 21712
rect 2810 21988 2938 22040
rect 2938 21988 3062 22040
rect 3062 21988 3190 22040
rect 2810 21712 3190 21988
rect 2810 21660 2938 21712
rect 2938 21660 3062 21712
rect 3062 21660 3190 21712
rect 3210 21988 3338 22040
rect 3338 21988 3462 22040
rect 3462 21988 3590 22040
rect 3210 21712 3590 21988
rect 3210 21660 3338 21712
rect 3338 21660 3462 21712
rect 3462 21660 3590 21712
rect 3610 21988 3738 22040
rect 3738 21988 3862 22040
rect 3862 21988 3990 22040
rect 3610 21712 3990 21988
rect 3610 21660 3738 21712
rect 3738 21660 3862 21712
rect 3862 21660 3990 21712
rect 4010 21988 4138 22040
rect 4138 21988 4262 22040
rect 4262 21988 4390 22040
rect 4010 21712 4390 21988
rect 4010 21660 4138 21712
rect 4138 21660 4262 21712
rect 4262 21660 4390 21712
rect 4410 21988 4538 22040
rect 4538 21988 4662 22040
rect 4662 21988 4790 22040
rect 4410 21712 4790 21988
rect 4410 21660 4538 21712
rect 4538 21660 4662 21712
rect 4662 21660 4790 21712
rect 4810 21988 4938 22040
rect 4938 21988 5062 22040
rect 5062 21988 5190 22040
rect 4810 21712 5190 21988
rect 4810 21660 4938 21712
rect 4938 21660 5062 21712
rect 5062 21660 5190 21712
rect 5210 21988 5338 22040
rect 5338 21988 5462 22040
rect 5462 21988 5590 22040
rect 5210 21712 5590 21988
rect 5210 21660 5338 21712
rect 5338 21660 5462 21712
rect 5462 21660 5590 21712
rect 5610 21988 5738 22040
rect 5738 21988 5862 22040
rect 5862 21988 5990 22040
rect 5610 21712 5990 21988
rect 5610 21660 5738 21712
rect 5738 21660 5862 21712
rect 5862 21660 5990 21712
rect 6010 21988 6138 22040
rect 6138 21988 6262 22040
rect 6262 21988 6390 22040
rect 6010 21712 6390 21988
rect 6010 21660 6138 21712
rect 6138 21660 6262 21712
rect 6262 21660 6390 21712
rect 6410 21988 6538 22040
rect 6538 21988 6662 22040
rect 6662 21988 6790 22040
rect 6410 21712 6790 21988
rect 6410 21660 6538 21712
rect 6538 21660 6662 21712
rect 6662 21660 6790 21712
rect 6810 21988 6938 22040
rect 6938 21988 7062 22040
rect 7062 21988 7190 22040
rect 6810 21712 7190 21988
rect 6810 21660 6938 21712
rect 6938 21660 7062 21712
rect 7062 21660 7190 21712
rect 7210 21988 7338 22040
rect 7338 21988 7462 22040
rect 7462 21988 7590 22040
rect 7210 21712 7590 21988
rect 7210 21660 7338 21712
rect 7338 21660 7462 21712
rect 7462 21660 7590 21712
rect 7610 21988 7738 22040
rect 7738 21988 7862 22040
rect 7862 21988 7990 22040
rect 7610 21712 7990 21988
rect 7610 21660 7738 21712
rect 7738 21660 7862 21712
rect 7862 21660 7990 21712
rect 8010 21988 8138 22040
rect 8138 21988 8262 22040
rect 8262 21988 8390 22040
rect 8010 21712 8390 21988
rect 8010 21660 8138 21712
rect 8138 21660 8262 21712
rect 8262 21660 8390 21712
rect 8410 21988 8538 22040
rect 8538 21988 8662 22040
rect 8662 21988 8790 22040
rect 8410 21712 8790 21988
rect 8410 21660 8538 21712
rect 8538 21660 8662 21712
rect 8662 21660 8790 21712
rect 8810 21988 8938 22040
rect 8938 21988 9062 22040
rect 9062 21988 9190 22040
rect 8810 21712 9190 21988
rect 8810 21660 8938 21712
rect 8938 21660 9062 21712
rect 9062 21660 9190 21712
rect 9210 21988 9338 22040
rect 9338 21988 9462 22040
rect 9462 21988 9590 22040
rect 9210 21712 9590 21988
rect 9210 21660 9338 21712
rect 9338 21660 9462 21712
rect 9462 21660 9590 21712
rect 9610 21988 9738 22040
rect 9738 21988 9862 22040
rect 9862 21988 9990 22040
rect 9610 21712 9990 21988
rect 9610 21660 9738 21712
rect 9738 21660 9862 21712
rect 9862 21660 9990 21712
rect 10010 21988 10138 22040
rect 10138 21988 10262 22040
rect 10262 21988 10390 22040
rect 10010 21712 10390 21988
rect 10010 21660 10138 21712
rect 10138 21660 10262 21712
rect 10262 21660 10390 21712
rect 10410 21988 10538 22040
rect 10538 21988 10662 22040
rect 10662 21988 10790 22040
rect 10410 21712 10790 21988
rect 10410 21660 10538 21712
rect 10538 21660 10662 21712
rect 10662 21660 10790 21712
rect 10810 21988 10938 22040
rect 10938 21988 11062 22040
rect 11062 21988 11190 22040
rect 10810 21712 11190 21988
rect 10810 21660 10938 21712
rect 10938 21660 11062 21712
rect 11062 21660 11190 21712
rect 11210 21988 11338 22040
rect 11338 21988 11462 22040
rect 11462 21988 11590 22040
rect 11210 21712 11590 21988
rect 11210 21660 11338 21712
rect 11338 21660 11462 21712
rect 11462 21660 11590 21712
rect 11610 21988 11738 22040
rect 11738 21988 11862 22040
rect 11862 21988 11990 22040
rect 11610 21712 11990 21988
rect 11610 21660 11738 21712
rect 11738 21660 11862 21712
rect 11862 21660 11990 21712
rect 12010 21988 12138 22040
rect 12138 21988 12262 22040
rect 12262 21988 12390 22040
rect 12010 21712 12390 21988
rect 12010 21660 12138 21712
rect 12138 21660 12262 21712
rect 12262 21660 12390 21712
rect 12410 21988 12538 22040
rect 12538 21988 12662 22040
rect 12662 21988 12790 22040
rect 12410 21712 12790 21988
rect 12410 21660 12538 21712
rect 12538 21660 12662 21712
rect 12662 21660 12790 21712
rect 12810 21988 12938 22040
rect 12938 21988 13062 22040
rect 13062 21988 13190 22040
rect 12810 21712 13190 21988
rect 12810 21660 12938 21712
rect 12938 21660 13062 21712
rect 13062 21660 13190 21712
rect 13210 21988 13338 22040
rect 13338 21988 13462 22040
rect 13462 21988 13590 22040
rect 13210 21712 13590 21988
rect 13210 21660 13338 21712
rect 13338 21660 13462 21712
rect 13462 21660 13590 21712
rect 13610 21988 13738 22040
rect 13738 21988 13862 22040
rect 13862 21988 13990 22040
rect 13610 21712 13990 21988
rect 13610 21660 13738 21712
rect 13738 21660 13862 21712
rect 13862 21660 13990 21712
rect 14010 21988 14138 22040
rect 14138 21988 14262 22040
rect 14262 21988 14390 22040
rect 14010 21712 14390 21988
rect 14010 21660 14138 21712
rect 14138 21660 14262 21712
rect 14262 21660 14390 21712
rect 14410 21988 14538 22040
rect 14538 21988 14662 22040
rect 14662 21988 14790 22040
rect 14410 21712 14790 21988
rect 14410 21660 14538 21712
rect 14538 21660 14662 21712
rect 14662 21660 14790 21712
rect 14810 21988 14938 22040
rect 14938 21988 15062 22040
rect 15062 21988 15190 22040
rect 14810 21712 15190 21988
rect 14810 21660 14938 21712
rect 14938 21660 15062 21712
rect 15062 21660 15190 21712
rect 15210 21988 15338 22040
rect 15338 21988 15462 22040
rect 15462 21988 15590 22040
rect 15210 21712 15590 21988
rect 15210 21660 15338 21712
rect 15338 21660 15462 21712
rect 15462 21660 15590 21712
rect 410 21588 538 21640
rect 538 21588 662 21640
rect 662 21588 790 21640
rect 410 21312 790 21588
rect 410 21260 538 21312
rect 538 21260 662 21312
rect 662 21260 790 21312
rect 810 21588 938 21640
rect 938 21588 1062 21640
rect 1062 21588 1190 21640
rect 810 21312 1190 21588
rect 810 21260 938 21312
rect 938 21260 1062 21312
rect 1062 21260 1190 21312
rect 1210 21588 1338 21640
rect 1338 21588 1462 21640
rect 1462 21588 1590 21640
rect 1210 21312 1590 21588
rect 1210 21260 1338 21312
rect 1338 21260 1462 21312
rect 1462 21260 1590 21312
rect 1610 21588 1738 21640
rect 1738 21588 1862 21640
rect 1862 21588 1990 21640
rect 1610 21312 1990 21588
rect 1610 21260 1738 21312
rect 1738 21260 1862 21312
rect 1862 21260 1990 21312
rect 2010 21588 2138 21640
rect 2138 21588 2262 21640
rect 2262 21588 2390 21640
rect 2010 21312 2390 21588
rect 2010 21260 2138 21312
rect 2138 21260 2262 21312
rect 2262 21260 2390 21312
rect 2410 21588 2538 21640
rect 2538 21588 2662 21640
rect 2662 21588 2790 21640
rect 2410 21312 2790 21588
rect 2410 21260 2538 21312
rect 2538 21260 2662 21312
rect 2662 21260 2790 21312
rect 2810 21588 2938 21640
rect 2938 21588 3062 21640
rect 3062 21588 3190 21640
rect 2810 21312 3190 21588
rect 2810 21260 2938 21312
rect 2938 21260 3062 21312
rect 3062 21260 3190 21312
rect 3210 21588 3338 21640
rect 3338 21588 3462 21640
rect 3462 21588 3590 21640
rect 3210 21312 3590 21588
rect 3210 21260 3338 21312
rect 3338 21260 3462 21312
rect 3462 21260 3590 21312
rect 3610 21588 3738 21640
rect 3738 21588 3862 21640
rect 3862 21588 3990 21640
rect 3610 21312 3990 21588
rect 3610 21260 3738 21312
rect 3738 21260 3862 21312
rect 3862 21260 3990 21312
rect 4010 21588 4138 21640
rect 4138 21588 4262 21640
rect 4262 21588 4390 21640
rect 4010 21312 4390 21588
rect 4010 21260 4138 21312
rect 4138 21260 4262 21312
rect 4262 21260 4390 21312
rect 4410 21588 4538 21640
rect 4538 21588 4662 21640
rect 4662 21588 4790 21640
rect 4410 21312 4790 21588
rect 4410 21260 4538 21312
rect 4538 21260 4662 21312
rect 4662 21260 4790 21312
rect 4810 21588 4938 21640
rect 4938 21588 5062 21640
rect 5062 21588 5190 21640
rect 4810 21312 5190 21588
rect 4810 21260 4938 21312
rect 4938 21260 5062 21312
rect 5062 21260 5190 21312
rect 5210 21588 5338 21640
rect 5338 21588 5462 21640
rect 5462 21588 5590 21640
rect 5210 21312 5590 21588
rect 5210 21260 5338 21312
rect 5338 21260 5462 21312
rect 5462 21260 5590 21312
rect 5610 21588 5738 21640
rect 5738 21588 5862 21640
rect 5862 21588 5990 21640
rect 5610 21312 5990 21588
rect 5610 21260 5738 21312
rect 5738 21260 5862 21312
rect 5862 21260 5990 21312
rect 6010 21588 6138 21640
rect 6138 21588 6262 21640
rect 6262 21588 6390 21640
rect 6010 21312 6390 21588
rect 6010 21260 6138 21312
rect 6138 21260 6262 21312
rect 6262 21260 6390 21312
rect 6410 21588 6538 21640
rect 6538 21588 6662 21640
rect 6662 21588 6790 21640
rect 6410 21312 6790 21588
rect 6410 21260 6538 21312
rect 6538 21260 6662 21312
rect 6662 21260 6790 21312
rect 6810 21588 6938 21640
rect 6938 21588 7062 21640
rect 7062 21588 7190 21640
rect 6810 21312 7190 21588
rect 6810 21260 6938 21312
rect 6938 21260 7062 21312
rect 7062 21260 7190 21312
rect 7210 21588 7338 21640
rect 7338 21588 7462 21640
rect 7462 21588 7590 21640
rect 7210 21312 7590 21588
rect 7210 21260 7338 21312
rect 7338 21260 7462 21312
rect 7462 21260 7590 21312
rect 7610 21588 7738 21640
rect 7738 21588 7862 21640
rect 7862 21588 7990 21640
rect 7610 21312 7990 21588
rect 7610 21260 7738 21312
rect 7738 21260 7862 21312
rect 7862 21260 7990 21312
rect 8010 21588 8138 21640
rect 8138 21588 8262 21640
rect 8262 21588 8390 21640
rect 8010 21312 8390 21588
rect 8010 21260 8138 21312
rect 8138 21260 8262 21312
rect 8262 21260 8390 21312
rect 8410 21588 8538 21640
rect 8538 21588 8662 21640
rect 8662 21588 8790 21640
rect 8410 21312 8790 21588
rect 8410 21260 8538 21312
rect 8538 21260 8662 21312
rect 8662 21260 8790 21312
rect 8810 21588 8938 21640
rect 8938 21588 9062 21640
rect 9062 21588 9190 21640
rect 8810 21312 9190 21588
rect 8810 21260 8938 21312
rect 8938 21260 9062 21312
rect 9062 21260 9190 21312
rect 9210 21588 9338 21640
rect 9338 21588 9462 21640
rect 9462 21588 9590 21640
rect 9210 21312 9590 21588
rect 9210 21260 9338 21312
rect 9338 21260 9462 21312
rect 9462 21260 9590 21312
rect 9610 21588 9738 21640
rect 9738 21588 9862 21640
rect 9862 21588 9990 21640
rect 9610 21312 9990 21588
rect 9610 21260 9738 21312
rect 9738 21260 9862 21312
rect 9862 21260 9990 21312
rect 10010 21588 10138 21640
rect 10138 21588 10262 21640
rect 10262 21588 10390 21640
rect 10010 21312 10390 21588
rect 10010 21260 10138 21312
rect 10138 21260 10262 21312
rect 10262 21260 10390 21312
rect 10410 21588 10538 21640
rect 10538 21588 10662 21640
rect 10662 21588 10790 21640
rect 10410 21312 10790 21588
rect 10410 21260 10538 21312
rect 10538 21260 10662 21312
rect 10662 21260 10790 21312
rect 10810 21588 10938 21640
rect 10938 21588 11062 21640
rect 11062 21588 11190 21640
rect 10810 21312 11190 21588
rect 10810 21260 10938 21312
rect 10938 21260 11062 21312
rect 11062 21260 11190 21312
rect 11210 21588 11338 21640
rect 11338 21588 11462 21640
rect 11462 21588 11590 21640
rect 11210 21312 11590 21588
rect 11210 21260 11338 21312
rect 11338 21260 11462 21312
rect 11462 21260 11590 21312
rect 11610 21588 11738 21640
rect 11738 21588 11862 21640
rect 11862 21588 11990 21640
rect 11610 21312 11990 21588
rect 11610 21260 11738 21312
rect 11738 21260 11862 21312
rect 11862 21260 11990 21312
rect 12010 21588 12138 21640
rect 12138 21588 12262 21640
rect 12262 21588 12390 21640
rect 12010 21312 12390 21588
rect 12010 21260 12138 21312
rect 12138 21260 12262 21312
rect 12262 21260 12390 21312
rect 12410 21588 12538 21640
rect 12538 21588 12662 21640
rect 12662 21588 12790 21640
rect 12410 21312 12790 21588
rect 12410 21260 12538 21312
rect 12538 21260 12662 21312
rect 12662 21260 12790 21312
rect 12810 21588 12938 21640
rect 12938 21588 13062 21640
rect 13062 21588 13190 21640
rect 12810 21312 13190 21588
rect 12810 21260 12938 21312
rect 12938 21260 13062 21312
rect 13062 21260 13190 21312
rect 13210 21588 13338 21640
rect 13338 21588 13462 21640
rect 13462 21588 13590 21640
rect 13210 21312 13590 21588
rect 13210 21260 13338 21312
rect 13338 21260 13462 21312
rect 13462 21260 13590 21312
rect 13610 21588 13738 21640
rect 13738 21588 13862 21640
rect 13862 21588 13990 21640
rect 13610 21312 13990 21588
rect 13610 21260 13738 21312
rect 13738 21260 13862 21312
rect 13862 21260 13990 21312
rect 14010 21588 14138 21640
rect 14138 21588 14262 21640
rect 14262 21588 14390 21640
rect 14010 21312 14390 21588
rect 14010 21260 14138 21312
rect 14138 21260 14262 21312
rect 14262 21260 14390 21312
rect 14410 21588 14538 21640
rect 14538 21588 14662 21640
rect 14662 21588 14790 21640
rect 14410 21312 14790 21588
rect 14410 21260 14538 21312
rect 14538 21260 14662 21312
rect 14662 21260 14790 21312
rect 14810 21588 14938 21640
rect 14938 21588 15062 21640
rect 15062 21588 15190 21640
rect 14810 21312 15190 21588
rect 14810 21260 14938 21312
rect 14938 21260 15062 21312
rect 15062 21260 15190 21312
rect 15210 21588 15338 21640
rect 15338 21588 15462 21640
rect 15462 21588 15590 21640
rect 15210 21312 15590 21588
rect 15210 21260 15338 21312
rect 15338 21260 15462 21312
rect 15462 21260 15590 21312
rect 410 21188 538 21240
rect 538 21188 662 21240
rect 662 21188 790 21240
rect 410 20912 790 21188
rect 410 20860 538 20912
rect 538 20860 662 20912
rect 662 20860 790 20912
rect 810 21188 938 21240
rect 938 21188 1062 21240
rect 1062 21188 1190 21240
rect 810 20912 1190 21188
rect 810 20860 938 20912
rect 938 20860 1062 20912
rect 1062 20860 1190 20912
rect 1210 21188 1338 21240
rect 1338 21188 1462 21240
rect 1462 21188 1590 21240
rect 1210 20912 1590 21188
rect 1210 20860 1338 20912
rect 1338 20860 1462 20912
rect 1462 20860 1590 20912
rect 1610 21188 1738 21240
rect 1738 21188 1862 21240
rect 1862 21188 1990 21240
rect 1610 20912 1990 21188
rect 1610 20860 1738 20912
rect 1738 20860 1862 20912
rect 1862 20860 1990 20912
rect 2010 21188 2138 21240
rect 2138 21188 2262 21240
rect 2262 21188 2390 21240
rect 2010 20912 2390 21188
rect 2010 20860 2138 20912
rect 2138 20860 2262 20912
rect 2262 20860 2390 20912
rect 2410 21188 2538 21240
rect 2538 21188 2662 21240
rect 2662 21188 2790 21240
rect 2410 20912 2790 21188
rect 2410 20860 2538 20912
rect 2538 20860 2662 20912
rect 2662 20860 2790 20912
rect 2810 21188 2938 21240
rect 2938 21188 3062 21240
rect 3062 21188 3190 21240
rect 2810 20912 3190 21188
rect 2810 20860 2938 20912
rect 2938 20860 3062 20912
rect 3062 20860 3190 20912
rect 3210 21188 3338 21240
rect 3338 21188 3462 21240
rect 3462 21188 3590 21240
rect 3210 20912 3590 21188
rect 3210 20860 3338 20912
rect 3338 20860 3462 20912
rect 3462 20860 3590 20912
rect 3610 21188 3738 21240
rect 3738 21188 3862 21240
rect 3862 21188 3990 21240
rect 3610 20912 3990 21188
rect 3610 20860 3738 20912
rect 3738 20860 3862 20912
rect 3862 20860 3990 20912
rect 4010 21188 4138 21240
rect 4138 21188 4262 21240
rect 4262 21188 4390 21240
rect 4010 20912 4390 21188
rect 4010 20860 4138 20912
rect 4138 20860 4262 20912
rect 4262 20860 4390 20912
rect 4410 21188 4538 21240
rect 4538 21188 4662 21240
rect 4662 21188 4790 21240
rect 4410 20912 4790 21188
rect 4410 20860 4538 20912
rect 4538 20860 4662 20912
rect 4662 20860 4790 20912
rect 4810 21188 4938 21240
rect 4938 21188 5062 21240
rect 5062 21188 5190 21240
rect 4810 20912 5190 21188
rect 4810 20860 4938 20912
rect 4938 20860 5062 20912
rect 5062 20860 5190 20912
rect 5210 21188 5338 21240
rect 5338 21188 5462 21240
rect 5462 21188 5590 21240
rect 5210 20912 5590 21188
rect 5210 20860 5338 20912
rect 5338 20860 5462 20912
rect 5462 20860 5590 20912
rect 5610 21188 5738 21240
rect 5738 21188 5862 21240
rect 5862 21188 5990 21240
rect 5610 20912 5990 21188
rect 5610 20860 5738 20912
rect 5738 20860 5862 20912
rect 5862 20860 5990 20912
rect 6010 21188 6138 21240
rect 6138 21188 6262 21240
rect 6262 21188 6390 21240
rect 6010 20912 6390 21188
rect 6010 20860 6138 20912
rect 6138 20860 6262 20912
rect 6262 20860 6390 20912
rect 6410 21188 6538 21240
rect 6538 21188 6662 21240
rect 6662 21188 6790 21240
rect 6410 20912 6790 21188
rect 6410 20860 6538 20912
rect 6538 20860 6662 20912
rect 6662 20860 6790 20912
rect 6810 21188 6938 21240
rect 6938 21188 7062 21240
rect 7062 21188 7190 21240
rect 6810 20912 7190 21188
rect 6810 20860 6938 20912
rect 6938 20860 7062 20912
rect 7062 20860 7190 20912
rect 7210 21188 7338 21240
rect 7338 21188 7462 21240
rect 7462 21188 7590 21240
rect 7210 20912 7590 21188
rect 7210 20860 7338 20912
rect 7338 20860 7462 20912
rect 7462 20860 7590 20912
rect 7610 21188 7738 21240
rect 7738 21188 7862 21240
rect 7862 21188 7990 21240
rect 7610 20912 7990 21188
rect 7610 20860 7738 20912
rect 7738 20860 7862 20912
rect 7862 20860 7990 20912
rect 8010 21188 8138 21240
rect 8138 21188 8262 21240
rect 8262 21188 8390 21240
rect 8010 20912 8390 21188
rect 8010 20860 8138 20912
rect 8138 20860 8262 20912
rect 8262 20860 8390 20912
rect 8410 21188 8538 21240
rect 8538 21188 8662 21240
rect 8662 21188 8790 21240
rect 8410 20912 8790 21188
rect 8410 20860 8538 20912
rect 8538 20860 8662 20912
rect 8662 20860 8790 20912
rect 8810 21188 8938 21240
rect 8938 21188 9062 21240
rect 9062 21188 9190 21240
rect 8810 20912 9190 21188
rect 8810 20860 8938 20912
rect 8938 20860 9062 20912
rect 9062 20860 9190 20912
rect 9210 21188 9338 21240
rect 9338 21188 9462 21240
rect 9462 21188 9590 21240
rect 9210 20912 9590 21188
rect 9210 20860 9338 20912
rect 9338 20860 9462 20912
rect 9462 20860 9590 20912
rect 9610 21188 9738 21240
rect 9738 21188 9862 21240
rect 9862 21188 9990 21240
rect 9610 20912 9990 21188
rect 9610 20860 9738 20912
rect 9738 20860 9862 20912
rect 9862 20860 9990 20912
rect 10010 21188 10138 21240
rect 10138 21188 10262 21240
rect 10262 21188 10390 21240
rect 10010 20912 10390 21188
rect 10010 20860 10138 20912
rect 10138 20860 10262 20912
rect 10262 20860 10390 20912
rect 10410 21188 10538 21240
rect 10538 21188 10662 21240
rect 10662 21188 10790 21240
rect 10410 20912 10790 21188
rect 10410 20860 10538 20912
rect 10538 20860 10662 20912
rect 10662 20860 10790 20912
rect 10810 21188 10938 21240
rect 10938 21188 11062 21240
rect 11062 21188 11190 21240
rect 10810 20912 11190 21188
rect 10810 20860 10938 20912
rect 10938 20860 11062 20912
rect 11062 20860 11190 20912
rect 11210 21188 11338 21240
rect 11338 21188 11462 21240
rect 11462 21188 11590 21240
rect 11210 20912 11590 21188
rect 11210 20860 11338 20912
rect 11338 20860 11462 20912
rect 11462 20860 11590 20912
rect 11610 21188 11738 21240
rect 11738 21188 11862 21240
rect 11862 21188 11990 21240
rect 11610 20912 11990 21188
rect 11610 20860 11738 20912
rect 11738 20860 11862 20912
rect 11862 20860 11990 20912
rect 12010 21188 12138 21240
rect 12138 21188 12262 21240
rect 12262 21188 12390 21240
rect 12010 20912 12390 21188
rect 12010 20860 12138 20912
rect 12138 20860 12262 20912
rect 12262 20860 12390 20912
rect 12410 21188 12538 21240
rect 12538 21188 12662 21240
rect 12662 21188 12790 21240
rect 12410 20912 12790 21188
rect 12410 20860 12538 20912
rect 12538 20860 12662 20912
rect 12662 20860 12790 20912
rect 12810 21188 12938 21240
rect 12938 21188 13062 21240
rect 13062 21188 13190 21240
rect 12810 20912 13190 21188
rect 12810 20860 12938 20912
rect 12938 20860 13062 20912
rect 13062 20860 13190 20912
rect 13210 21188 13338 21240
rect 13338 21188 13462 21240
rect 13462 21188 13590 21240
rect 13210 20912 13590 21188
rect 13210 20860 13338 20912
rect 13338 20860 13462 20912
rect 13462 20860 13590 20912
rect 13610 21188 13738 21240
rect 13738 21188 13862 21240
rect 13862 21188 13990 21240
rect 13610 20912 13990 21188
rect 13610 20860 13738 20912
rect 13738 20860 13862 20912
rect 13862 20860 13990 20912
rect 14010 21188 14138 21240
rect 14138 21188 14262 21240
rect 14262 21188 14390 21240
rect 14010 20912 14390 21188
rect 14010 20860 14138 20912
rect 14138 20860 14262 20912
rect 14262 20860 14390 20912
rect 14410 21188 14538 21240
rect 14538 21188 14662 21240
rect 14662 21188 14790 21240
rect 14410 20912 14790 21188
rect 14410 20860 14538 20912
rect 14538 20860 14662 20912
rect 14662 20860 14790 20912
rect 14810 21188 14938 21240
rect 14938 21188 15062 21240
rect 15062 21188 15190 21240
rect 14810 20912 15190 21188
rect 14810 20860 14938 20912
rect 14938 20860 15062 20912
rect 15062 20860 15190 20912
rect 15210 21188 15338 21240
rect 15338 21188 15462 21240
rect 15462 21188 15590 21240
rect 15210 20912 15590 21188
rect 15210 20860 15338 20912
rect 15338 20860 15462 20912
rect 15462 20860 15590 20912
rect 410 20788 538 20840
rect 538 20788 662 20840
rect 662 20788 790 20840
rect 410 20512 790 20788
rect 410 20460 538 20512
rect 538 20460 662 20512
rect 662 20460 790 20512
rect 810 20788 938 20840
rect 938 20788 1062 20840
rect 1062 20788 1190 20840
rect 810 20512 1190 20788
rect 810 20460 938 20512
rect 938 20460 1062 20512
rect 1062 20460 1190 20512
rect 1210 20788 1338 20840
rect 1338 20788 1462 20840
rect 1462 20788 1590 20840
rect 1210 20512 1590 20788
rect 1210 20460 1338 20512
rect 1338 20460 1462 20512
rect 1462 20460 1590 20512
rect 1610 20788 1738 20840
rect 1738 20788 1862 20840
rect 1862 20788 1990 20840
rect 1610 20512 1990 20788
rect 1610 20460 1738 20512
rect 1738 20460 1862 20512
rect 1862 20460 1990 20512
rect 2010 20788 2138 20840
rect 2138 20788 2262 20840
rect 2262 20788 2390 20840
rect 2010 20512 2390 20788
rect 2010 20460 2138 20512
rect 2138 20460 2262 20512
rect 2262 20460 2390 20512
rect 2410 20788 2538 20840
rect 2538 20788 2662 20840
rect 2662 20788 2790 20840
rect 2410 20512 2790 20788
rect 2410 20460 2538 20512
rect 2538 20460 2662 20512
rect 2662 20460 2790 20512
rect 2810 20788 2938 20840
rect 2938 20788 3062 20840
rect 3062 20788 3190 20840
rect 2810 20512 3190 20788
rect 2810 20460 2938 20512
rect 2938 20460 3062 20512
rect 3062 20460 3190 20512
rect 3210 20788 3338 20840
rect 3338 20788 3462 20840
rect 3462 20788 3590 20840
rect 3210 20512 3590 20788
rect 3210 20460 3338 20512
rect 3338 20460 3462 20512
rect 3462 20460 3590 20512
rect 3610 20788 3738 20840
rect 3738 20788 3862 20840
rect 3862 20788 3990 20840
rect 3610 20512 3990 20788
rect 3610 20460 3738 20512
rect 3738 20460 3862 20512
rect 3862 20460 3990 20512
rect 4010 20788 4138 20840
rect 4138 20788 4262 20840
rect 4262 20788 4390 20840
rect 4010 20512 4390 20788
rect 4010 20460 4138 20512
rect 4138 20460 4262 20512
rect 4262 20460 4390 20512
rect 4410 20788 4538 20840
rect 4538 20788 4662 20840
rect 4662 20788 4790 20840
rect 4410 20512 4790 20788
rect 4410 20460 4538 20512
rect 4538 20460 4662 20512
rect 4662 20460 4790 20512
rect 4810 20788 4938 20840
rect 4938 20788 5062 20840
rect 5062 20788 5190 20840
rect 4810 20512 5190 20788
rect 4810 20460 4938 20512
rect 4938 20460 5062 20512
rect 5062 20460 5190 20512
rect 5210 20788 5338 20840
rect 5338 20788 5462 20840
rect 5462 20788 5590 20840
rect 5210 20512 5590 20788
rect 5210 20460 5338 20512
rect 5338 20460 5462 20512
rect 5462 20460 5590 20512
rect 5610 20788 5738 20840
rect 5738 20788 5862 20840
rect 5862 20788 5990 20840
rect 5610 20512 5990 20788
rect 5610 20460 5738 20512
rect 5738 20460 5862 20512
rect 5862 20460 5990 20512
rect 6010 20788 6138 20840
rect 6138 20788 6262 20840
rect 6262 20788 6390 20840
rect 6010 20512 6390 20788
rect 6010 20460 6138 20512
rect 6138 20460 6262 20512
rect 6262 20460 6390 20512
rect 6410 20788 6538 20840
rect 6538 20788 6662 20840
rect 6662 20788 6790 20840
rect 6410 20512 6790 20788
rect 6410 20460 6538 20512
rect 6538 20460 6662 20512
rect 6662 20460 6790 20512
rect 6810 20788 6938 20840
rect 6938 20788 7062 20840
rect 7062 20788 7190 20840
rect 6810 20512 7190 20788
rect 6810 20460 6938 20512
rect 6938 20460 7062 20512
rect 7062 20460 7190 20512
rect 7210 20788 7338 20840
rect 7338 20788 7462 20840
rect 7462 20788 7590 20840
rect 7210 20512 7590 20788
rect 7210 20460 7338 20512
rect 7338 20460 7462 20512
rect 7462 20460 7590 20512
rect 7610 20788 7738 20840
rect 7738 20788 7862 20840
rect 7862 20788 7990 20840
rect 7610 20512 7990 20788
rect 7610 20460 7738 20512
rect 7738 20460 7862 20512
rect 7862 20460 7990 20512
rect 8010 20788 8138 20840
rect 8138 20788 8262 20840
rect 8262 20788 8390 20840
rect 8010 20512 8390 20788
rect 8010 20460 8138 20512
rect 8138 20460 8262 20512
rect 8262 20460 8390 20512
rect 8410 20788 8538 20840
rect 8538 20788 8662 20840
rect 8662 20788 8790 20840
rect 8410 20512 8790 20788
rect 8410 20460 8538 20512
rect 8538 20460 8662 20512
rect 8662 20460 8790 20512
rect 8810 20788 8938 20840
rect 8938 20788 9062 20840
rect 9062 20788 9190 20840
rect 8810 20512 9190 20788
rect 8810 20460 8938 20512
rect 8938 20460 9062 20512
rect 9062 20460 9190 20512
rect 9210 20788 9338 20840
rect 9338 20788 9462 20840
rect 9462 20788 9590 20840
rect 9210 20512 9590 20788
rect 9210 20460 9338 20512
rect 9338 20460 9462 20512
rect 9462 20460 9590 20512
rect 9610 20788 9738 20840
rect 9738 20788 9862 20840
rect 9862 20788 9990 20840
rect 9610 20512 9990 20788
rect 9610 20460 9738 20512
rect 9738 20460 9862 20512
rect 9862 20460 9990 20512
rect 10010 20788 10138 20840
rect 10138 20788 10262 20840
rect 10262 20788 10390 20840
rect 10010 20512 10390 20788
rect 10010 20460 10138 20512
rect 10138 20460 10262 20512
rect 10262 20460 10390 20512
rect 10410 20788 10538 20840
rect 10538 20788 10662 20840
rect 10662 20788 10790 20840
rect 10410 20512 10790 20788
rect 10410 20460 10538 20512
rect 10538 20460 10662 20512
rect 10662 20460 10790 20512
rect 10810 20788 10938 20840
rect 10938 20788 11062 20840
rect 11062 20788 11190 20840
rect 10810 20512 11190 20788
rect 10810 20460 10938 20512
rect 10938 20460 11062 20512
rect 11062 20460 11190 20512
rect 11210 20788 11338 20840
rect 11338 20788 11462 20840
rect 11462 20788 11590 20840
rect 11210 20512 11590 20788
rect 11210 20460 11338 20512
rect 11338 20460 11462 20512
rect 11462 20460 11590 20512
rect 11610 20788 11738 20840
rect 11738 20788 11862 20840
rect 11862 20788 11990 20840
rect 11610 20512 11990 20788
rect 11610 20460 11738 20512
rect 11738 20460 11862 20512
rect 11862 20460 11990 20512
rect 12010 20788 12138 20840
rect 12138 20788 12262 20840
rect 12262 20788 12390 20840
rect 12010 20512 12390 20788
rect 12010 20460 12138 20512
rect 12138 20460 12262 20512
rect 12262 20460 12390 20512
rect 12410 20788 12538 20840
rect 12538 20788 12662 20840
rect 12662 20788 12790 20840
rect 12410 20512 12790 20788
rect 12410 20460 12538 20512
rect 12538 20460 12662 20512
rect 12662 20460 12790 20512
rect 12810 20788 12938 20840
rect 12938 20788 13062 20840
rect 13062 20788 13190 20840
rect 12810 20512 13190 20788
rect 12810 20460 12938 20512
rect 12938 20460 13062 20512
rect 13062 20460 13190 20512
rect 13210 20788 13338 20840
rect 13338 20788 13462 20840
rect 13462 20788 13590 20840
rect 13210 20512 13590 20788
rect 13210 20460 13338 20512
rect 13338 20460 13462 20512
rect 13462 20460 13590 20512
rect 13610 20788 13738 20840
rect 13738 20788 13862 20840
rect 13862 20788 13990 20840
rect 13610 20512 13990 20788
rect 13610 20460 13738 20512
rect 13738 20460 13862 20512
rect 13862 20460 13990 20512
rect 14010 20788 14138 20840
rect 14138 20788 14262 20840
rect 14262 20788 14390 20840
rect 14010 20512 14390 20788
rect 14010 20460 14138 20512
rect 14138 20460 14262 20512
rect 14262 20460 14390 20512
rect 14410 20788 14538 20840
rect 14538 20788 14662 20840
rect 14662 20788 14790 20840
rect 14410 20512 14790 20788
rect 14410 20460 14538 20512
rect 14538 20460 14662 20512
rect 14662 20460 14790 20512
rect 14810 20788 14938 20840
rect 14938 20788 15062 20840
rect 15062 20788 15190 20840
rect 14810 20512 15190 20788
rect 14810 20460 14938 20512
rect 14938 20460 15062 20512
rect 15062 20460 15190 20512
rect 15210 20788 15338 20840
rect 15338 20788 15462 20840
rect 15462 20788 15590 20840
rect 15210 20512 15590 20788
rect 15210 20460 15338 20512
rect 15338 20460 15462 20512
rect 15462 20460 15590 20512
rect 410 20388 538 20440
rect 538 20388 662 20440
rect 662 20388 790 20440
rect 410 20112 790 20388
rect 410 20060 538 20112
rect 538 20060 662 20112
rect 662 20060 790 20112
rect 810 20388 938 20440
rect 938 20388 1062 20440
rect 1062 20388 1190 20440
rect 810 20112 1190 20388
rect 810 20060 938 20112
rect 938 20060 1062 20112
rect 1062 20060 1190 20112
rect 1210 20388 1338 20440
rect 1338 20388 1462 20440
rect 1462 20388 1590 20440
rect 1210 20112 1590 20388
rect 1210 20060 1338 20112
rect 1338 20060 1462 20112
rect 1462 20060 1590 20112
rect 1610 20388 1738 20440
rect 1738 20388 1862 20440
rect 1862 20388 1990 20440
rect 1610 20112 1990 20388
rect 1610 20060 1738 20112
rect 1738 20060 1862 20112
rect 1862 20060 1990 20112
rect 2010 20388 2138 20440
rect 2138 20388 2262 20440
rect 2262 20388 2390 20440
rect 2010 20112 2390 20388
rect 2010 20060 2138 20112
rect 2138 20060 2262 20112
rect 2262 20060 2390 20112
rect 2410 20388 2538 20440
rect 2538 20388 2662 20440
rect 2662 20388 2790 20440
rect 2410 20112 2790 20388
rect 2410 20060 2538 20112
rect 2538 20060 2662 20112
rect 2662 20060 2790 20112
rect 2810 20388 2938 20440
rect 2938 20388 3062 20440
rect 3062 20388 3190 20440
rect 2810 20112 3190 20388
rect 2810 20060 2938 20112
rect 2938 20060 3062 20112
rect 3062 20060 3190 20112
rect 3210 20388 3338 20440
rect 3338 20388 3462 20440
rect 3462 20388 3590 20440
rect 3210 20112 3590 20388
rect 3210 20060 3338 20112
rect 3338 20060 3462 20112
rect 3462 20060 3590 20112
rect 3610 20388 3738 20440
rect 3738 20388 3862 20440
rect 3862 20388 3990 20440
rect 3610 20112 3990 20388
rect 3610 20060 3738 20112
rect 3738 20060 3862 20112
rect 3862 20060 3990 20112
rect 4010 20388 4138 20440
rect 4138 20388 4262 20440
rect 4262 20388 4390 20440
rect 4010 20112 4390 20388
rect 4010 20060 4138 20112
rect 4138 20060 4262 20112
rect 4262 20060 4390 20112
rect 4410 20388 4538 20440
rect 4538 20388 4662 20440
rect 4662 20388 4790 20440
rect 4410 20112 4790 20388
rect 4410 20060 4538 20112
rect 4538 20060 4662 20112
rect 4662 20060 4790 20112
rect 4810 20388 4938 20440
rect 4938 20388 5062 20440
rect 5062 20388 5190 20440
rect 4810 20112 5190 20388
rect 4810 20060 4938 20112
rect 4938 20060 5062 20112
rect 5062 20060 5190 20112
rect 5210 20388 5338 20440
rect 5338 20388 5462 20440
rect 5462 20388 5590 20440
rect 5210 20112 5590 20388
rect 5210 20060 5338 20112
rect 5338 20060 5462 20112
rect 5462 20060 5590 20112
rect 5610 20388 5738 20440
rect 5738 20388 5862 20440
rect 5862 20388 5990 20440
rect 5610 20112 5990 20388
rect 5610 20060 5738 20112
rect 5738 20060 5862 20112
rect 5862 20060 5990 20112
rect 6010 20388 6138 20440
rect 6138 20388 6262 20440
rect 6262 20388 6390 20440
rect 6010 20112 6390 20388
rect 6010 20060 6138 20112
rect 6138 20060 6262 20112
rect 6262 20060 6390 20112
rect 6410 20388 6538 20440
rect 6538 20388 6662 20440
rect 6662 20388 6790 20440
rect 6410 20112 6790 20388
rect 6410 20060 6538 20112
rect 6538 20060 6662 20112
rect 6662 20060 6790 20112
rect 6810 20388 6938 20440
rect 6938 20388 7062 20440
rect 7062 20388 7190 20440
rect 6810 20112 7190 20388
rect 6810 20060 6938 20112
rect 6938 20060 7062 20112
rect 7062 20060 7190 20112
rect 7210 20388 7338 20440
rect 7338 20388 7462 20440
rect 7462 20388 7590 20440
rect 7210 20112 7590 20388
rect 7210 20060 7338 20112
rect 7338 20060 7462 20112
rect 7462 20060 7590 20112
rect 7610 20388 7738 20440
rect 7738 20388 7862 20440
rect 7862 20388 7990 20440
rect 7610 20112 7990 20388
rect 7610 20060 7738 20112
rect 7738 20060 7862 20112
rect 7862 20060 7990 20112
rect 8010 20388 8138 20440
rect 8138 20388 8262 20440
rect 8262 20388 8390 20440
rect 8010 20112 8390 20388
rect 8010 20060 8138 20112
rect 8138 20060 8262 20112
rect 8262 20060 8390 20112
rect 8410 20388 8538 20440
rect 8538 20388 8662 20440
rect 8662 20388 8790 20440
rect 8410 20112 8790 20388
rect 8410 20060 8538 20112
rect 8538 20060 8662 20112
rect 8662 20060 8790 20112
rect 8810 20388 8938 20440
rect 8938 20388 9062 20440
rect 9062 20388 9190 20440
rect 8810 20112 9190 20388
rect 8810 20060 8938 20112
rect 8938 20060 9062 20112
rect 9062 20060 9190 20112
rect 9210 20388 9338 20440
rect 9338 20388 9462 20440
rect 9462 20388 9590 20440
rect 9210 20112 9590 20388
rect 9210 20060 9338 20112
rect 9338 20060 9462 20112
rect 9462 20060 9590 20112
rect 9610 20388 9738 20440
rect 9738 20388 9862 20440
rect 9862 20388 9990 20440
rect 9610 20112 9990 20388
rect 9610 20060 9738 20112
rect 9738 20060 9862 20112
rect 9862 20060 9990 20112
rect 10010 20388 10138 20440
rect 10138 20388 10262 20440
rect 10262 20388 10390 20440
rect 10010 20112 10390 20388
rect 10010 20060 10138 20112
rect 10138 20060 10262 20112
rect 10262 20060 10390 20112
rect 10410 20388 10538 20440
rect 10538 20388 10662 20440
rect 10662 20388 10790 20440
rect 10410 20112 10790 20388
rect 10410 20060 10538 20112
rect 10538 20060 10662 20112
rect 10662 20060 10790 20112
rect 10810 20388 10938 20440
rect 10938 20388 11062 20440
rect 11062 20388 11190 20440
rect 10810 20112 11190 20388
rect 10810 20060 10938 20112
rect 10938 20060 11062 20112
rect 11062 20060 11190 20112
rect 11210 20388 11338 20440
rect 11338 20388 11462 20440
rect 11462 20388 11590 20440
rect 11210 20112 11590 20388
rect 11210 20060 11338 20112
rect 11338 20060 11462 20112
rect 11462 20060 11590 20112
rect 11610 20388 11738 20440
rect 11738 20388 11862 20440
rect 11862 20388 11990 20440
rect 11610 20112 11990 20388
rect 11610 20060 11738 20112
rect 11738 20060 11862 20112
rect 11862 20060 11990 20112
rect 12010 20388 12138 20440
rect 12138 20388 12262 20440
rect 12262 20388 12390 20440
rect 12010 20112 12390 20388
rect 12010 20060 12138 20112
rect 12138 20060 12262 20112
rect 12262 20060 12390 20112
rect 12410 20388 12538 20440
rect 12538 20388 12662 20440
rect 12662 20388 12790 20440
rect 12410 20112 12790 20388
rect 12410 20060 12538 20112
rect 12538 20060 12662 20112
rect 12662 20060 12790 20112
rect 12810 20388 12938 20440
rect 12938 20388 13062 20440
rect 13062 20388 13190 20440
rect 12810 20112 13190 20388
rect 12810 20060 12938 20112
rect 12938 20060 13062 20112
rect 13062 20060 13190 20112
rect 13210 20388 13338 20440
rect 13338 20388 13462 20440
rect 13462 20388 13590 20440
rect 13210 20112 13590 20388
rect 13210 20060 13338 20112
rect 13338 20060 13462 20112
rect 13462 20060 13590 20112
rect 13610 20388 13738 20440
rect 13738 20388 13862 20440
rect 13862 20388 13990 20440
rect 13610 20112 13990 20388
rect 13610 20060 13738 20112
rect 13738 20060 13862 20112
rect 13862 20060 13990 20112
rect 14010 20388 14138 20440
rect 14138 20388 14262 20440
rect 14262 20388 14390 20440
rect 14010 20112 14390 20388
rect 14010 20060 14138 20112
rect 14138 20060 14262 20112
rect 14262 20060 14390 20112
rect 14410 20388 14538 20440
rect 14538 20388 14662 20440
rect 14662 20388 14790 20440
rect 14410 20112 14790 20388
rect 14410 20060 14538 20112
rect 14538 20060 14662 20112
rect 14662 20060 14790 20112
rect 14810 20388 14938 20440
rect 14938 20388 15062 20440
rect 15062 20388 15190 20440
rect 14810 20112 15190 20388
rect 14810 20060 14938 20112
rect 14938 20060 15062 20112
rect 15062 20060 15190 20112
rect 15210 20388 15338 20440
rect 15338 20388 15462 20440
rect 15462 20388 15590 20440
rect 15210 20112 15590 20388
rect 15210 20060 15338 20112
rect 15338 20060 15462 20112
rect 15462 20060 15590 20112
rect 410 19988 538 20040
rect 538 19988 662 20040
rect 662 19988 790 20040
rect 410 19712 790 19988
rect 410 19660 538 19712
rect 538 19660 662 19712
rect 662 19660 790 19712
rect 810 19988 938 20040
rect 938 19988 1062 20040
rect 1062 19988 1190 20040
rect 810 19712 1190 19988
rect 810 19660 938 19712
rect 938 19660 1062 19712
rect 1062 19660 1190 19712
rect 1210 19988 1338 20040
rect 1338 19988 1462 20040
rect 1462 19988 1590 20040
rect 1210 19712 1590 19988
rect 1210 19660 1338 19712
rect 1338 19660 1462 19712
rect 1462 19660 1590 19712
rect 1610 19988 1738 20040
rect 1738 19988 1862 20040
rect 1862 19988 1990 20040
rect 1610 19712 1990 19988
rect 1610 19660 1738 19712
rect 1738 19660 1862 19712
rect 1862 19660 1990 19712
rect 2010 19988 2138 20040
rect 2138 19988 2262 20040
rect 2262 19988 2390 20040
rect 2010 19712 2390 19988
rect 2010 19660 2138 19712
rect 2138 19660 2262 19712
rect 2262 19660 2390 19712
rect 2410 19988 2538 20040
rect 2538 19988 2662 20040
rect 2662 19988 2790 20040
rect 2410 19712 2790 19988
rect 2410 19660 2538 19712
rect 2538 19660 2662 19712
rect 2662 19660 2790 19712
rect 2810 19988 2938 20040
rect 2938 19988 3062 20040
rect 3062 19988 3190 20040
rect 2810 19712 3190 19988
rect 2810 19660 2938 19712
rect 2938 19660 3062 19712
rect 3062 19660 3190 19712
rect 3210 19988 3338 20040
rect 3338 19988 3462 20040
rect 3462 19988 3590 20040
rect 3210 19712 3590 19988
rect 3210 19660 3338 19712
rect 3338 19660 3462 19712
rect 3462 19660 3590 19712
rect 3610 19988 3738 20040
rect 3738 19988 3862 20040
rect 3862 19988 3990 20040
rect 3610 19712 3990 19988
rect 3610 19660 3738 19712
rect 3738 19660 3862 19712
rect 3862 19660 3990 19712
rect 4010 19988 4138 20040
rect 4138 19988 4262 20040
rect 4262 19988 4390 20040
rect 4010 19712 4390 19988
rect 4010 19660 4138 19712
rect 4138 19660 4262 19712
rect 4262 19660 4390 19712
rect 4410 19988 4538 20040
rect 4538 19988 4662 20040
rect 4662 19988 4790 20040
rect 4410 19712 4790 19988
rect 4410 19660 4538 19712
rect 4538 19660 4662 19712
rect 4662 19660 4790 19712
rect 4810 19988 4938 20040
rect 4938 19988 5062 20040
rect 5062 19988 5190 20040
rect 4810 19712 5190 19988
rect 4810 19660 4938 19712
rect 4938 19660 5062 19712
rect 5062 19660 5190 19712
rect 5210 19988 5338 20040
rect 5338 19988 5462 20040
rect 5462 19988 5590 20040
rect 5210 19712 5590 19988
rect 5210 19660 5338 19712
rect 5338 19660 5462 19712
rect 5462 19660 5590 19712
rect 5610 19988 5738 20040
rect 5738 19988 5862 20040
rect 5862 19988 5990 20040
rect 5610 19712 5990 19988
rect 5610 19660 5738 19712
rect 5738 19660 5862 19712
rect 5862 19660 5990 19712
rect 6010 19988 6138 20040
rect 6138 19988 6262 20040
rect 6262 19988 6390 20040
rect 6010 19712 6390 19988
rect 6010 19660 6138 19712
rect 6138 19660 6262 19712
rect 6262 19660 6390 19712
rect 6410 19988 6538 20040
rect 6538 19988 6662 20040
rect 6662 19988 6790 20040
rect 6410 19712 6790 19988
rect 6410 19660 6538 19712
rect 6538 19660 6662 19712
rect 6662 19660 6790 19712
rect 6810 19988 6938 20040
rect 6938 19988 7062 20040
rect 7062 19988 7190 20040
rect 6810 19712 7190 19988
rect 6810 19660 6938 19712
rect 6938 19660 7062 19712
rect 7062 19660 7190 19712
rect 7210 19988 7338 20040
rect 7338 19988 7462 20040
rect 7462 19988 7590 20040
rect 7210 19712 7590 19988
rect 7210 19660 7338 19712
rect 7338 19660 7462 19712
rect 7462 19660 7590 19712
rect 7610 19988 7738 20040
rect 7738 19988 7862 20040
rect 7862 19988 7990 20040
rect 7610 19712 7990 19988
rect 7610 19660 7738 19712
rect 7738 19660 7862 19712
rect 7862 19660 7990 19712
rect 8010 19988 8138 20040
rect 8138 19988 8262 20040
rect 8262 19988 8390 20040
rect 8010 19712 8390 19988
rect 8010 19660 8138 19712
rect 8138 19660 8262 19712
rect 8262 19660 8390 19712
rect 8410 19988 8538 20040
rect 8538 19988 8662 20040
rect 8662 19988 8790 20040
rect 8410 19712 8790 19988
rect 8410 19660 8538 19712
rect 8538 19660 8662 19712
rect 8662 19660 8790 19712
rect 8810 19988 8938 20040
rect 8938 19988 9062 20040
rect 9062 19988 9190 20040
rect 8810 19712 9190 19988
rect 8810 19660 8938 19712
rect 8938 19660 9062 19712
rect 9062 19660 9190 19712
rect 9210 19988 9338 20040
rect 9338 19988 9462 20040
rect 9462 19988 9590 20040
rect 9210 19712 9590 19988
rect 9210 19660 9338 19712
rect 9338 19660 9462 19712
rect 9462 19660 9590 19712
rect 9610 19988 9738 20040
rect 9738 19988 9862 20040
rect 9862 19988 9990 20040
rect 9610 19712 9990 19988
rect 9610 19660 9738 19712
rect 9738 19660 9862 19712
rect 9862 19660 9990 19712
rect 10010 19988 10138 20040
rect 10138 19988 10262 20040
rect 10262 19988 10390 20040
rect 10010 19712 10390 19988
rect 10010 19660 10138 19712
rect 10138 19660 10262 19712
rect 10262 19660 10390 19712
rect 10410 19988 10538 20040
rect 10538 19988 10662 20040
rect 10662 19988 10790 20040
rect 10410 19712 10790 19988
rect 10410 19660 10538 19712
rect 10538 19660 10662 19712
rect 10662 19660 10790 19712
rect 10810 19988 10938 20040
rect 10938 19988 11062 20040
rect 11062 19988 11190 20040
rect 10810 19712 11190 19988
rect 10810 19660 10938 19712
rect 10938 19660 11062 19712
rect 11062 19660 11190 19712
rect 11210 19988 11338 20040
rect 11338 19988 11462 20040
rect 11462 19988 11590 20040
rect 11210 19712 11590 19988
rect 11210 19660 11338 19712
rect 11338 19660 11462 19712
rect 11462 19660 11590 19712
rect 11610 19988 11738 20040
rect 11738 19988 11862 20040
rect 11862 19988 11990 20040
rect 11610 19712 11990 19988
rect 11610 19660 11738 19712
rect 11738 19660 11862 19712
rect 11862 19660 11990 19712
rect 12010 19988 12138 20040
rect 12138 19988 12262 20040
rect 12262 19988 12390 20040
rect 12010 19712 12390 19988
rect 12010 19660 12138 19712
rect 12138 19660 12262 19712
rect 12262 19660 12390 19712
rect 12410 19988 12538 20040
rect 12538 19988 12662 20040
rect 12662 19988 12790 20040
rect 12410 19712 12790 19988
rect 12410 19660 12538 19712
rect 12538 19660 12662 19712
rect 12662 19660 12790 19712
rect 12810 19988 12938 20040
rect 12938 19988 13062 20040
rect 13062 19988 13190 20040
rect 12810 19712 13190 19988
rect 12810 19660 12938 19712
rect 12938 19660 13062 19712
rect 13062 19660 13190 19712
rect 13210 19988 13338 20040
rect 13338 19988 13462 20040
rect 13462 19988 13590 20040
rect 13210 19712 13590 19988
rect 13210 19660 13338 19712
rect 13338 19660 13462 19712
rect 13462 19660 13590 19712
rect 13610 19988 13738 20040
rect 13738 19988 13862 20040
rect 13862 19988 13990 20040
rect 13610 19712 13990 19988
rect 13610 19660 13738 19712
rect 13738 19660 13862 19712
rect 13862 19660 13990 19712
rect 14010 19988 14138 20040
rect 14138 19988 14262 20040
rect 14262 19988 14390 20040
rect 14010 19712 14390 19988
rect 14010 19660 14138 19712
rect 14138 19660 14262 19712
rect 14262 19660 14390 19712
rect 14410 19988 14538 20040
rect 14538 19988 14662 20040
rect 14662 19988 14790 20040
rect 14410 19712 14790 19988
rect 14410 19660 14538 19712
rect 14538 19660 14662 19712
rect 14662 19660 14790 19712
rect 14810 19988 14938 20040
rect 14938 19988 15062 20040
rect 15062 19988 15190 20040
rect 14810 19712 15190 19988
rect 14810 19660 14938 19712
rect 14938 19660 15062 19712
rect 15062 19660 15190 19712
rect 15210 19988 15338 20040
rect 15338 19988 15462 20040
rect 15462 19988 15590 20040
rect 15210 19712 15590 19988
rect 15210 19660 15338 19712
rect 15338 19660 15462 19712
rect 15462 19660 15590 19712
rect 410 19588 538 19640
rect 538 19588 662 19640
rect 662 19588 790 19640
rect 410 19312 790 19588
rect 410 19260 538 19312
rect 538 19260 662 19312
rect 662 19260 790 19312
rect 810 19588 938 19640
rect 938 19588 1062 19640
rect 1062 19588 1190 19640
rect 810 19312 1190 19588
rect 810 19260 938 19312
rect 938 19260 1062 19312
rect 1062 19260 1190 19312
rect 1210 19588 1338 19640
rect 1338 19588 1462 19640
rect 1462 19588 1590 19640
rect 1210 19312 1590 19588
rect 1210 19260 1338 19312
rect 1338 19260 1462 19312
rect 1462 19260 1590 19312
rect 1610 19588 1738 19640
rect 1738 19588 1862 19640
rect 1862 19588 1990 19640
rect 1610 19312 1990 19588
rect 1610 19260 1738 19312
rect 1738 19260 1862 19312
rect 1862 19260 1990 19312
rect 2010 19588 2138 19640
rect 2138 19588 2262 19640
rect 2262 19588 2390 19640
rect 2010 19312 2390 19588
rect 2010 19260 2138 19312
rect 2138 19260 2262 19312
rect 2262 19260 2390 19312
rect 2410 19588 2538 19640
rect 2538 19588 2662 19640
rect 2662 19588 2790 19640
rect 2410 19312 2790 19588
rect 2410 19260 2538 19312
rect 2538 19260 2662 19312
rect 2662 19260 2790 19312
rect 2810 19588 2938 19640
rect 2938 19588 3062 19640
rect 3062 19588 3190 19640
rect 2810 19312 3190 19588
rect 2810 19260 2938 19312
rect 2938 19260 3062 19312
rect 3062 19260 3190 19312
rect 3210 19588 3338 19640
rect 3338 19588 3462 19640
rect 3462 19588 3590 19640
rect 3210 19312 3590 19588
rect 3210 19260 3338 19312
rect 3338 19260 3462 19312
rect 3462 19260 3590 19312
rect 3610 19588 3738 19640
rect 3738 19588 3862 19640
rect 3862 19588 3990 19640
rect 3610 19312 3990 19588
rect 3610 19260 3738 19312
rect 3738 19260 3862 19312
rect 3862 19260 3990 19312
rect 4010 19588 4138 19640
rect 4138 19588 4262 19640
rect 4262 19588 4390 19640
rect 4010 19312 4390 19588
rect 4010 19260 4138 19312
rect 4138 19260 4262 19312
rect 4262 19260 4390 19312
rect 4410 19588 4538 19640
rect 4538 19588 4662 19640
rect 4662 19588 4790 19640
rect 4410 19312 4790 19588
rect 4410 19260 4538 19312
rect 4538 19260 4662 19312
rect 4662 19260 4790 19312
rect 4810 19588 4938 19640
rect 4938 19588 5062 19640
rect 5062 19588 5190 19640
rect 4810 19312 5190 19588
rect 4810 19260 4938 19312
rect 4938 19260 5062 19312
rect 5062 19260 5190 19312
rect 5210 19588 5338 19640
rect 5338 19588 5462 19640
rect 5462 19588 5590 19640
rect 5210 19312 5590 19588
rect 5210 19260 5338 19312
rect 5338 19260 5462 19312
rect 5462 19260 5590 19312
rect 5610 19588 5738 19640
rect 5738 19588 5862 19640
rect 5862 19588 5990 19640
rect 5610 19312 5990 19588
rect 5610 19260 5738 19312
rect 5738 19260 5862 19312
rect 5862 19260 5990 19312
rect 6010 19588 6138 19640
rect 6138 19588 6262 19640
rect 6262 19588 6390 19640
rect 6010 19312 6390 19588
rect 6010 19260 6138 19312
rect 6138 19260 6262 19312
rect 6262 19260 6390 19312
rect 6410 19588 6538 19640
rect 6538 19588 6662 19640
rect 6662 19588 6790 19640
rect 6410 19312 6790 19588
rect 6410 19260 6538 19312
rect 6538 19260 6662 19312
rect 6662 19260 6790 19312
rect 6810 19588 6938 19640
rect 6938 19588 7062 19640
rect 7062 19588 7190 19640
rect 6810 19312 7190 19588
rect 6810 19260 6938 19312
rect 6938 19260 7062 19312
rect 7062 19260 7190 19312
rect 7210 19588 7338 19640
rect 7338 19588 7462 19640
rect 7462 19588 7590 19640
rect 7210 19312 7590 19588
rect 7210 19260 7338 19312
rect 7338 19260 7462 19312
rect 7462 19260 7590 19312
rect 7610 19588 7738 19640
rect 7738 19588 7862 19640
rect 7862 19588 7990 19640
rect 7610 19312 7990 19588
rect 7610 19260 7738 19312
rect 7738 19260 7862 19312
rect 7862 19260 7990 19312
rect 8010 19588 8138 19640
rect 8138 19588 8262 19640
rect 8262 19588 8390 19640
rect 8010 19312 8390 19588
rect 8010 19260 8138 19312
rect 8138 19260 8262 19312
rect 8262 19260 8390 19312
rect 8410 19588 8538 19640
rect 8538 19588 8662 19640
rect 8662 19588 8790 19640
rect 8410 19312 8790 19588
rect 8410 19260 8538 19312
rect 8538 19260 8662 19312
rect 8662 19260 8790 19312
rect 8810 19588 8938 19640
rect 8938 19588 9062 19640
rect 9062 19588 9190 19640
rect 8810 19312 9190 19588
rect 8810 19260 8938 19312
rect 8938 19260 9062 19312
rect 9062 19260 9190 19312
rect 9210 19588 9338 19640
rect 9338 19588 9462 19640
rect 9462 19588 9590 19640
rect 9210 19312 9590 19588
rect 9210 19260 9338 19312
rect 9338 19260 9462 19312
rect 9462 19260 9590 19312
rect 9610 19588 9738 19640
rect 9738 19588 9862 19640
rect 9862 19588 9990 19640
rect 9610 19312 9990 19588
rect 9610 19260 9738 19312
rect 9738 19260 9862 19312
rect 9862 19260 9990 19312
rect 10010 19588 10138 19640
rect 10138 19588 10262 19640
rect 10262 19588 10390 19640
rect 10010 19312 10390 19588
rect 10010 19260 10138 19312
rect 10138 19260 10262 19312
rect 10262 19260 10390 19312
rect 10410 19588 10538 19640
rect 10538 19588 10662 19640
rect 10662 19588 10790 19640
rect 10410 19312 10790 19588
rect 10410 19260 10538 19312
rect 10538 19260 10662 19312
rect 10662 19260 10790 19312
rect 10810 19588 10938 19640
rect 10938 19588 11062 19640
rect 11062 19588 11190 19640
rect 10810 19312 11190 19588
rect 10810 19260 10938 19312
rect 10938 19260 11062 19312
rect 11062 19260 11190 19312
rect 11210 19588 11338 19640
rect 11338 19588 11462 19640
rect 11462 19588 11590 19640
rect 11210 19312 11590 19588
rect 11210 19260 11338 19312
rect 11338 19260 11462 19312
rect 11462 19260 11590 19312
rect 11610 19588 11738 19640
rect 11738 19588 11862 19640
rect 11862 19588 11990 19640
rect 11610 19312 11990 19588
rect 11610 19260 11738 19312
rect 11738 19260 11862 19312
rect 11862 19260 11990 19312
rect 12010 19588 12138 19640
rect 12138 19588 12262 19640
rect 12262 19588 12390 19640
rect 12010 19312 12390 19588
rect 12010 19260 12138 19312
rect 12138 19260 12262 19312
rect 12262 19260 12390 19312
rect 12410 19588 12538 19640
rect 12538 19588 12662 19640
rect 12662 19588 12790 19640
rect 12410 19312 12790 19588
rect 12410 19260 12538 19312
rect 12538 19260 12662 19312
rect 12662 19260 12790 19312
rect 12810 19588 12938 19640
rect 12938 19588 13062 19640
rect 13062 19588 13190 19640
rect 12810 19312 13190 19588
rect 12810 19260 12938 19312
rect 12938 19260 13062 19312
rect 13062 19260 13190 19312
rect 13210 19588 13338 19640
rect 13338 19588 13462 19640
rect 13462 19588 13590 19640
rect 13210 19312 13590 19588
rect 13210 19260 13338 19312
rect 13338 19260 13462 19312
rect 13462 19260 13590 19312
rect 13610 19588 13738 19640
rect 13738 19588 13862 19640
rect 13862 19588 13990 19640
rect 13610 19312 13990 19588
rect 13610 19260 13738 19312
rect 13738 19260 13862 19312
rect 13862 19260 13990 19312
rect 14010 19588 14138 19640
rect 14138 19588 14262 19640
rect 14262 19588 14390 19640
rect 14010 19312 14390 19588
rect 14010 19260 14138 19312
rect 14138 19260 14262 19312
rect 14262 19260 14390 19312
rect 14410 19588 14538 19640
rect 14538 19588 14662 19640
rect 14662 19588 14790 19640
rect 14410 19312 14790 19588
rect 14410 19260 14538 19312
rect 14538 19260 14662 19312
rect 14662 19260 14790 19312
rect 14810 19588 14938 19640
rect 14938 19588 15062 19640
rect 15062 19588 15190 19640
rect 14810 19312 15190 19588
rect 14810 19260 14938 19312
rect 14938 19260 15062 19312
rect 15062 19260 15190 19312
rect 15210 19588 15338 19640
rect 15338 19588 15462 19640
rect 15462 19588 15590 19640
rect 15210 19312 15590 19588
rect 15210 19260 15338 19312
rect 15338 19260 15462 19312
rect 15462 19260 15590 19312
rect 410 17688 538 17740
rect 538 17688 662 17740
rect 662 17688 790 17740
rect 410 17412 790 17688
rect 410 17360 538 17412
rect 538 17360 662 17412
rect 662 17360 790 17412
rect 810 17688 938 17740
rect 938 17688 1062 17740
rect 1062 17688 1190 17740
rect 810 17412 1190 17688
rect 810 17360 938 17412
rect 938 17360 1062 17412
rect 1062 17360 1190 17412
rect 1210 17688 1338 17740
rect 1338 17688 1462 17740
rect 1462 17688 1590 17740
rect 1210 17412 1590 17688
rect 1210 17360 1338 17412
rect 1338 17360 1462 17412
rect 1462 17360 1590 17412
rect 1610 17688 1738 17740
rect 1738 17688 1862 17740
rect 1862 17688 1990 17740
rect 1610 17412 1990 17688
rect 1610 17360 1738 17412
rect 1738 17360 1862 17412
rect 1862 17360 1990 17412
rect 2010 17688 2138 17740
rect 2138 17688 2262 17740
rect 2262 17688 2390 17740
rect 2010 17412 2390 17688
rect 2010 17360 2138 17412
rect 2138 17360 2262 17412
rect 2262 17360 2390 17412
rect 2410 17688 2538 17740
rect 2538 17688 2662 17740
rect 2662 17688 2790 17740
rect 2410 17412 2790 17688
rect 2410 17360 2538 17412
rect 2538 17360 2662 17412
rect 2662 17360 2790 17412
rect 2810 17688 2938 17740
rect 2938 17688 3062 17740
rect 3062 17688 3190 17740
rect 2810 17412 3190 17688
rect 2810 17360 2938 17412
rect 2938 17360 3062 17412
rect 3062 17360 3190 17412
rect 3210 17688 3338 17740
rect 3338 17688 3462 17740
rect 3462 17688 3590 17740
rect 3210 17412 3590 17688
rect 3210 17360 3338 17412
rect 3338 17360 3462 17412
rect 3462 17360 3590 17412
rect 3610 17688 3738 17740
rect 3738 17688 3862 17740
rect 3862 17688 3990 17740
rect 3610 17412 3990 17688
rect 3610 17360 3738 17412
rect 3738 17360 3862 17412
rect 3862 17360 3990 17412
rect 4010 17688 4138 17740
rect 4138 17688 4262 17740
rect 4262 17688 4390 17740
rect 4010 17412 4390 17688
rect 4010 17360 4138 17412
rect 4138 17360 4262 17412
rect 4262 17360 4390 17412
rect 4410 17688 4538 17740
rect 4538 17688 4662 17740
rect 4662 17688 4790 17740
rect 4410 17412 4790 17688
rect 4410 17360 4538 17412
rect 4538 17360 4662 17412
rect 4662 17360 4790 17412
rect 4810 17688 4938 17740
rect 4938 17688 5062 17740
rect 5062 17688 5190 17740
rect 4810 17412 5190 17688
rect 4810 17360 4938 17412
rect 4938 17360 5062 17412
rect 5062 17360 5190 17412
rect 5210 17688 5338 17740
rect 5338 17688 5462 17740
rect 5462 17688 5590 17740
rect 5210 17412 5590 17688
rect 5210 17360 5338 17412
rect 5338 17360 5462 17412
rect 5462 17360 5590 17412
rect 5610 17688 5738 17740
rect 5738 17688 5862 17740
rect 5862 17688 5990 17740
rect 5610 17412 5990 17688
rect 5610 17360 5738 17412
rect 5738 17360 5862 17412
rect 5862 17360 5990 17412
rect 6010 17688 6138 17740
rect 6138 17688 6262 17740
rect 6262 17688 6390 17740
rect 6010 17412 6390 17688
rect 6010 17360 6138 17412
rect 6138 17360 6262 17412
rect 6262 17360 6390 17412
rect 6410 17688 6538 17740
rect 6538 17688 6662 17740
rect 6662 17688 6790 17740
rect 6410 17412 6790 17688
rect 6410 17360 6538 17412
rect 6538 17360 6662 17412
rect 6662 17360 6790 17412
rect 6810 17688 6938 17740
rect 6938 17688 7062 17740
rect 7062 17688 7190 17740
rect 6810 17412 7190 17688
rect 6810 17360 6938 17412
rect 6938 17360 7062 17412
rect 7062 17360 7190 17412
rect 7210 17688 7338 17740
rect 7338 17688 7462 17740
rect 7462 17688 7590 17740
rect 7210 17412 7590 17688
rect 7210 17360 7338 17412
rect 7338 17360 7462 17412
rect 7462 17360 7590 17412
rect 7610 17688 7738 17740
rect 7738 17688 7862 17740
rect 7862 17688 7990 17740
rect 7610 17412 7990 17688
rect 7610 17360 7738 17412
rect 7738 17360 7862 17412
rect 7862 17360 7990 17412
rect 8010 17688 8138 17740
rect 8138 17688 8262 17740
rect 8262 17688 8390 17740
rect 8010 17412 8390 17688
rect 8010 17360 8138 17412
rect 8138 17360 8262 17412
rect 8262 17360 8390 17412
rect 8410 17688 8538 17740
rect 8538 17688 8662 17740
rect 8662 17688 8790 17740
rect 8410 17412 8790 17688
rect 8410 17360 8538 17412
rect 8538 17360 8662 17412
rect 8662 17360 8790 17412
rect 8810 17688 8938 17740
rect 8938 17688 9062 17740
rect 9062 17688 9190 17740
rect 8810 17412 9190 17688
rect 8810 17360 8938 17412
rect 8938 17360 9062 17412
rect 9062 17360 9190 17412
rect 9210 17688 9338 17740
rect 9338 17688 9462 17740
rect 9462 17688 9590 17740
rect 9210 17412 9590 17688
rect 9210 17360 9338 17412
rect 9338 17360 9462 17412
rect 9462 17360 9590 17412
rect 9610 17688 9738 17740
rect 9738 17688 9862 17740
rect 9862 17688 9990 17740
rect 9610 17412 9990 17688
rect 9610 17360 9738 17412
rect 9738 17360 9862 17412
rect 9862 17360 9990 17412
rect 10010 17688 10138 17740
rect 10138 17688 10262 17740
rect 10262 17688 10390 17740
rect 10010 17412 10390 17688
rect 10010 17360 10138 17412
rect 10138 17360 10262 17412
rect 10262 17360 10390 17412
rect 10410 17688 10538 17740
rect 10538 17688 10662 17740
rect 10662 17688 10790 17740
rect 10410 17412 10790 17688
rect 10410 17360 10538 17412
rect 10538 17360 10662 17412
rect 10662 17360 10790 17412
rect 10810 17688 10938 17740
rect 10938 17688 11062 17740
rect 11062 17688 11190 17740
rect 10810 17412 11190 17688
rect 10810 17360 10938 17412
rect 10938 17360 11062 17412
rect 11062 17360 11190 17412
rect 11210 17688 11338 17740
rect 11338 17688 11462 17740
rect 11462 17688 11590 17740
rect 11210 17412 11590 17688
rect 11210 17360 11338 17412
rect 11338 17360 11462 17412
rect 11462 17360 11590 17412
rect 11610 17688 11738 17740
rect 11738 17688 11862 17740
rect 11862 17688 11990 17740
rect 11610 17412 11990 17688
rect 11610 17360 11738 17412
rect 11738 17360 11862 17412
rect 11862 17360 11990 17412
rect 12010 17688 12138 17740
rect 12138 17688 12262 17740
rect 12262 17688 12390 17740
rect 12010 17412 12390 17688
rect 12010 17360 12138 17412
rect 12138 17360 12262 17412
rect 12262 17360 12390 17412
rect 12410 17688 12538 17740
rect 12538 17688 12662 17740
rect 12662 17688 12790 17740
rect 12410 17412 12790 17688
rect 12410 17360 12538 17412
rect 12538 17360 12662 17412
rect 12662 17360 12790 17412
rect 12810 17688 12938 17740
rect 12938 17688 13062 17740
rect 13062 17688 13190 17740
rect 12810 17412 13190 17688
rect 12810 17360 12938 17412
rect 12938 17360 13062 17412
rect 13062 17360 13190 17412
rect 13210 17688 13338 17740
rect 13338 17688 13462 17740
rect 13462 17688 13590 17740
rect 13210 17412 13590 17688
rect 13210 17360 13338 17412
rect 13338 17360 13462 17412
rect 13462 17360 13590 17412
rect 13610 17688 13738 17740
rect 13738 17688 13862 17740
rect 13862 17688 13990 17740
rect 13610 17412 13990 17688
rect 13610 17360 13738 17412
rect 13738 17360 13862 17412
rect 13862 17360 13990 17412
rect 14010 17688 14138 17740
rect 14138 17688 14262 17740
rect 14262 17688 14390 17740
rect 14010 17412 14390 17688
rect 14010 17360 14138 17412
rect 14138 17360 14262 17412
rect 14262 17360 14390 17412
rect 14410 17688 14538 17740
rect 14538 17688 14662 17740
rect 14662 17688 14790 17740
rect 14410 17412 14790 17688
rect 14410 17360 14538 17412
rect 14538 17360 14662 17412
rect 14662 17360 14790 17412
rect 14810 17688 14938 17740
rect 14938 17688 15062 17740
rect 15062 17688 15190 17740
rect 14810 17412 15190 17688
rect 14810 17360 14938 17412
rect 14938 17360 15062 17412
rect 15062 17360 15190 17412
rect 15210 17688 15338 17740
rect 15338 17688 15462 17740
rect 15462 17688 15590 17740
rect 15210 17412 15590 17688
rect 15210 17360 15338 17412
rect 15338 17360 15462 17412
rect 15462 17360 15590 17412
rect 410 17288 538 17340
rect 538 17288 662 17340
rect 662 17288 790 17340
rect 410 17012 790 17288
rect 410 16960 538 17012
rect 538 16960 662 17012
rect 662 16960 790 17012
rect 810 17288 938 17340
rect 938 17288 1062 17340
rect 1062 17288 1190 17340
rect 810 17012 1190 17288
rect 810 16960 938 17012
rect 938 16960 1062 17012
rect 1062 16960 1190 17012
rect 1210 17288 1338 17340
rect 1338 17288 1462 17340
rect 1462 17288 1590 17340
rect 1210 17012 1590 17288
rect 1210 16960 1338 17012
rect 1338 16960 1462 17012
rect 1462 16960 1590 17012
rect 1610 17288 1738 17340
rect 1738 17288 1862 17340
rect 1862 17288 1990 17340
rect 1610 17012 1990 17288
rect 1610 16960 1738 17012
rect 1738 16960 1862 17012
rect 1862 16960 1990 17012
rect 2010 17288 2138 17340
rect 2138 17288 2262 17340
rect 2262 17288 2390 17340
rect 2010 17012 2390 17288
rect 2010 16960 2138 17012
rect 2138 16960 2262 17012
rect 2262 16960 2390 17012
rect 2410 17288 2538 17340
rect 2538 17288 2662 17340
rect 2662 17288 2790 17340
rect 2410 17012 2790 17288
rect 2410 16960 2538 17012
rect 2538 16960 2662 17012
rect 2662 16960 2790 17012
rect 2810 17288 2938 17340
rect 2938 17288 3062 17340
rect 3062 17288 3190 17340
rect 2810 17012 3190 17288
rect 2810 16960 2938 17012
rect 2938 16960 3062 17012
rect 3062 16960 3190 17012
rect 3210 17288 3338 17340
rect 3338 17288 3462 17340
rect 3462 17288 3590 17340
rect 3210 17012 3590 17288
rect 3210 16960 3338 17012
rect 3338 16960 3462 17012
rect 3462 16960 3590 17012
rect 3610 17288 3738 17340
rect 3738 17288 3862 17340
rect 3862 17288 3990 17340
rect 3610 17012 3990 17288
rect 3610 16960 3738 17012
rect 3738 16960 3862 17012
rect 3862 16960 3990 17012
rect 4010 17288 4138 17340
rect 4138 17288 4262 17340
rect 4262 17288 4390 17340
rect 4010 17012 4390 17288
rect 4010 16960 4138 17012
rect 4138 16960 4262 17012
rect 4262 16960 4390 17012
rect 4410 17288 4538 17340
rect 4538 17288 4662 17340
rect 4662 17288 4790 17340
rect 4410 17012 4790 17288
rect 4410 16960 4538 17012
rect 4538 16960 4662 17012
rect 4662 16960 4790 17012
rect 4810 17288 4938 17340
rect 4938 17288 5062 17340
rect 5062 17288 5190 17340
rect 4810 17012 5190 17288
rect 4810 16960 4938 17012
rect 4938 16960 5062 17012
rect 5062 16960 5190 17012
rect 5210 17288 5338 17340
rect 5338 17288 5462 17340
rect 5462 17288 5590 17340
rect 5210 17012 5590 17288
rect 5210 16960 5338 17012
rect 5338 16960 5462 17012
rect 5462 16960 5590 17012
rect 5610 17288 5738 17340
rect 5738 17288 5862 17340
rect 5862 17288 5990 17340
rect 5610 17012 5990 17288
rect 5610 16960 5738 17012
rect 5738 16960 5862 17012
rect 5862 16960 5990 17012
rect 6010 17288 6138 17340
rect 6138 17288 6262 17340
rect 6262 17288 6390 17340
rect 6010 17012 6390 17288
rect 6010 16960 6138 17012
rect 6138 16960 6262 17012
rect 6262 16960 6390 17012
rect 6410 17288 6538 17340
rect 6538 17288 6662 17340
rect 6662 17288 6790 17340
rect 6410 17012 6790 17288
rect 6410 16960 6538 17012
rect 6538 16960 6662 17012
rect 6662 16960 6790 17012
rect 6810 17288 6938 17340
rect 6938 17288 7062 17340
rect 7062 17288 7190 17340
rect 6810 17012 7190 17288
rect 6810 16960 6938 17012
rect 6938 16960 7062 17012
rect 7062 16960 7190 17012
rect 7210 17288 7338 17340
rect 7338 17288 7462 17340
rect 7462 17288 7590 17340
rect 7210 17012 7590 17288
rect 7210 16960 7338 17012
rect 7338 16960 7462 17012
rect 7462 16960 7590 17012
rect 7610 17288 7738 17340
rect 7738 17288 7862 17340
rect 7862 17288 7990 17340
rect 7610 17012 7990 17288
rect 7610 16960 7738 17012
rect 7738 16960 7862 17012
rect 7862 16960 7990 17012
rect 8010 17288 8138 17340
rect 8138 17288 8262 17340
rect 8262 17288 8390 17340
rect 8010 17012 8390 17288
rect 8010 16960 8138 17012
rect 8138 16960 8262 17012
rect 8262 16960 8390 17012
rect 8410 17288 8538 17340
rect 8538 17288 8662 17340
rect 8662 17288 8790 17340
rect 8410 17012 8790 17288
rect 8410 16960 8538 17012
rect 8538 16960 8662 17012
rect 8662 16960 8790 17012
rect 8810 17288 8938 17340
rect 8938 17288 9062 17340
rect 9062 17288 9190 17340
rect 8810 17012 9190 17288
rect 8810 16960 8938 17012
rect 8938 16960 9062 17012
rect 9062 16960 9190 17012
rect 9210 17288 9338 17340
rect 9338 17288 9462 17340
rect 9462 17288 9590 17340
rect 9210 17012 9590 17288
rect 9210 16960 9338 17012
rect 9338 16960 9462 17012
rect 9462 16960 9590 17012
rect 9610 17288 9738 17340
rect 9738 17288 9862 17340
rect 9862 17288 9990 17340
rect 9610 17012 9990 17288
rect 9610 16960 9738 17012
rect 9738 16960 9862 17012
rect 9862 16960 9990 17012
rect 10010 17288 10138 17340
rect 10138 17288 10262 17340
rect 10262 17288 10390 17340
rect 10010 17012 10390 17288
rect 10010 16960 10138 17012
rect 10138 16960 10262 17012
rect 10262 16960 10390 17012
rect 10410 17288 10538 17340
rect 10538 17288 10662 17340
rect 10662 17288 10790 17340
rect 10410 17012 10790 17288
rect 10410 16960 10538 17012
rect 10538 16960 10662 17012
rect 10662 16960 10790 17012
rect 10810 17288 10938 17340
rect 10938 17288 11062 17340
rect 11062 17288 11190 17340
rect 10810 17012 11190 17288
rect 10810 16960 10938 17012
rect 10938 16960 11062 17012
rect 11062 16960 11190 17012
rect 11210 17288 11338 17340
rect 11338 17288 11462 17340
rect 11462 17288 11590 17340
rect 11210 17012 11590 17288
rect 11210 16960 11338 17012
rect 11338 16960 11462 17012
rect 11462 16960 11590 17012
rect 11610 17288 11738 17340
rect 11738 17288 11862 17340
rect 11862 17288 11990 17340
rect 11610 17012 11990 17288
rect 11610 16960 11738 17012
rect 11738 16960 11862 17012
rect 11862 16960 11990 17012
rect 12010 17288 12138 17340
rect 12138 17288 12262 17340
rect 12262 17288 12390 17340
rect 12010 17012 12390 17288
rect 12010 16960 12138 17012
rect 12138 16960 12262 17012
rect 12262 16960 12390 17012
rect 12410 17288 12538 17340
rect 12538 17288 12662 17340
rect 12662 17288 12790 17340
rect 12410 17012 12790 17288
rect 12410 16960 12538 17012
rect 12538 16960 12662 17012
rect 12662 16960 12790 17012
rect 12810 17288 12938 17340
rect 12938 17288 13062 17340
rect 13062 17288 13190 17340
rect 12810 17012 13190 17288
rect 12810 16960 12938 17012
rect 12938 16960 13062 17012
rect 13062 16960 13190 17012
rect 13210 17288 13338 17340
rect 13338 17288 13462 17340
rect 13462 17288 13590 17340
rect 13210 17012 13590 17288
rect 13210 16960 13338 17012
rect 13338 16960 13462 17012
rect 13462 16960 13590 17012
rect 13610 17288 13738 17340
rect 13738 17288 13862 17340
rect 13862 17288 13990 17340
rect 13610 17012 13990 17288
rect 13610 16960 13738 17012
rect 13738 16960 13862 17012
rect 13862 16960 13990 17012
rect 14010 17288 14138 17340
rect 14138 17288 14262 17340
rect 14262 17288 14390 17340
rect 14010 17012 14390 17288
rect 14010 16960 14138 17012
rect 14138 16960 14262 17012
rect 14262 16960 14390 17012
rect 14410 17288 14538 17340
rect 14538 17288 14662 17340
rect 14662 17288 14790 17340
rect 14410 17012 14790 17288
rect 14410 16960 14538 17012
rect 14538 16960 14662 17012
rect 14662 16960 14790 17012
rect 14810 17288 14938 17340
rect 14938 17288 15062 17340
rect 15062 17288 15190 17340
rect 14810 17012 15190 17288
rect 14810 16960 14938 17012
rect 14938 16960 15062 17012
rect 15062 16960 15190 17012
rect 15210 17288 15338 17340
rect 15338 17288 15462 17340
rect 15462 17288 15590 17340
rect 15210 17012 15590 17288
rect 15210 16960 15338 17012
rect 15338 16960 15462 17012
rect 15462 16960 15590 17012
rect 410 16888 538 16940
rect 538 16888 662 16940
rect 662 16888 790 16940
rect 410 16612 790 16888
rect 410 16560 538 16612
rect 538 16560 662 16612
rect 662 16560 790 16612
rect 810 16888 938 16940
rect 938 16888 1062 16940
rect 1062 16888 1190 16940
rect 810 16612 1190 16888
rect 810 16560 938 16612
rect 938 16560 1062 16612
rect 1062 16560 1190 16612
rect 1210 16888 1338 16940
rect 1338 16888 1462 16940
rect 1462 16888 1590 16940
rect 1210 16612 1590 16888
rect 1210 16560 1338 16612
rect 1338 16560 1462 16612
rect 1462 16560 1590 16612
rect 1610 16888 1738 16940
rect 1738 16888 1862 16940
rect 1862 16888 1990 16940
rect 1610 16612 1990 16888
rect 1610 16560 1738 16612
rect 1738 16560 1862 16612
rect 1862 16560 1990 16612
rect 2010 16888 2138 16940
rect 2138 16888 2262 16940
rect 2262 16888 2390 16940
rect 2010 16612 2390 16888
rect 2010 16560 2138 16612
rect 2138 16560 2262 16612
rect 2262 16560 2390 16612
rect 2410 16888 2538 16940
rect 2538 16888 2662 16940
rect 2662 16888 2790 16940
rect 2410 16612 2790 16888
rect 2410 16560 2538 16612
rect 2538 16560 2662 16612
rect 2662 16560 2790 16612
rect 2810 16888 2938 16940
rect 2938 16888 3062 16940
rect 3062 16888 3190 16940
rect 2810 16612 3190 16888
rect 2810 16560 2938 16612
rect 2938 16560 3062 16612
rect 3062 16560 3190 16612
rect 3210 16888 3338 16940
rect 3338 16888 3462 16940
rect 3462 16888 3590 16940
rect 3210 16612 3590 16888
rect 3210 16560 3338 16612
rect 3338 16560 3462 16612
rect 3462 16560 3590 16612
rect 3610 16888 3738 16940
rect 3738 16888 3862 16940
rect 3862 16888 3990 16940
rect 3610 16612 3990 16888
rect 3610 16560 3738 16612
rect 3738 16560 3862 16612
rect 3862 16560 3990 16612
rect 4010 16888 4138 16940
rect 4138 16888 4262 16940
rect 4262 16888 4390 16940
rect 4010 16612 4390 16888
rect 4010 16560 4138 16612
rect 4138 16560 4262 16612
rect 4262 16560 4390 16612
rect 4410 16888 4538 16940
rect 4538 16888 4662 16940
rect 4662 16888 4790 16940
rect 4410 16612 4790 16888
rect 4410 16560 4538 16612
rect 4538 16560 4662 16612
rect 4662 16560 4790 16612
rect 4810 16888 4938 16940
rect 4938 16888 5062 16940
rect 5062 16888 5190 16940
rect 4810 16612 5190 16888
rect 4810 16560 4938 16612
rect 4938 16560 5062 16612
rect 5062 16560 5190 16612
rect 5210 16888 5338 16940
rect 5338 16888 5462 16940
rect 5462 16888 5590 16940
rect 5210 16612 5590 16888
rect 5210 16560 5338 16612
rect 5338 16560 5462 16612
rect 5462 16560 5590 16612
rect 5610 16888 5738 16940
rect 5738 16888 5862 16940
rect 5862 16888 5990 16940
rect 5610 16612 5990 16888
rect 5610 16560 5738 16612
rect 5738 16560 5862 16612
rect 5862 16560 5990 16612
rect 6010 16888 6138 16940
rect 6138 16888 6262 16940
rect 6262 16888 6390 16940
rect 6010 16612 6390 16888
rect 6010 16560 6138 16612
rect 6138 16560 6262 16612
rect 6262 16560 6390 16612
rect 6410 16888 6538 16940
rect 6538 16888 6662 16940
rect 6662 16888 6790 16940
rect 6410 16612 6790 16888
rect 6410 16560 6538 16612
rect 6538 16560 6662 16612
rect 6662 16560 6790 16612
rect 6810 16888 6938 16940
rect 6938 16888 7062 16940
rect 7062 16888 7190 16940
rect 6810 16612 7190 16888
rect 6810 16560 6938 16612
rect 6938 16560 7062 16612
rect 7062 16560 7190 16612
rect 7210 16888 7338 16940
rect 7338 16888 7462 16940
rect 7462 16888 7590 16940
rect 7210 16612 7590 16888
rect 7210 16560 7338 16612
rect 7338 16560 7462 16612
rect 7462 16560 7590 16612
rect 7610 16888 7738 16940
rect 7738 16888 7862 16940
rect 7862 16888 7990 16940
rect 7610 16612 7990 16888
rect 7610 16560 7738 16612
rect 7738 16560 7862 16612
rect 7862 16560 7990 16612
rect 8010 16888 8138 16940
rect 8138 16888 8262 16940
rect 8262 16888 8390 16940
rect 8010 16612 8390 16888
rect 8010 16560 8138 16612
rect 8138 16560 8262 16612
rect 8262 16560 8390 16612
rect 8410 16888 8538 16940
rect 8538 16888 8662 16940
rect 8662 16888 8790 16940
rect 8410 16612 8790 16888
rect 8410 16560 8538 16612
rect 8538 16560 8662 16612
rect 8662 16560 8790 16612
rect 8810 16888 8938 16940
rect 8938 16888 9062 16940
rect 9062 16888 9190 16940
rect 8810 16612 9190 16888
rect 8810 16560 8938 16612
rect 8938 16560 9062 16612
rect 9062 16560 9190 16612
rect 9210 16888 9338 16940
rect 9338 16888 9462 16940
rect 9462 16888 9590 16940
rect 9210 16612 9590 16888
rect 9210 16560 9338 16612
rect 9338 16560 9462 16612
rect 9462 16560 9590 16612
rect 9610 16888 9738 16940
rect 9738 16888 9862 16940
rect 9862 16888 9990 16940
rect 9610 16612 9990 16888
rect 9610 16560 9738 16612
rect 9738 16560 9862 16612
rect 9862 16560 9990 16612
rect 10010 16888 10138 16940
rect 10138 16888 10262 16940
rect 10262 16888 10390 16940
rect 10010 16612 10390 16888
rect 10010 16560 10138 16612
rect 10138 16560 10262 16612
rect 10262 16560 10390 16612
rect 10410 16888 10538 16940
rect 10538 16888 10662 16940
rect 10662 16888 10790 16940
rect 10410 16612 10790 16888
rect 10410 16560 10538 16612
rect 10538 16560 10662 16612
rect 10662 16560 10790 16612
rect 10810 16888 10938 16940
rect 10938 16888 11062 16940
rect 11062 16888 11190 16940
rect 10810 16612 11190 16888
rect 10810 16560 10938 16612
rect 10938 16560 11062 16612
rect 11062 16560 11190 16612
rect 11210 16888 11338 16940
rect 11338 16888 11462 16940
rect 11462 16888 11590 16940
rect 11210 16612 11590 16888
rect 11210 16560 11338 16612
rect 11338 16560 11462 16612
rect 11462 16560 11590 16612
rect 11610 16888 11738 16940
rect 11738 16888 11862 16940
rect 11862 16888 11990 16940
rect 11610 16612 11990 16888
rect 11610 16560 11738 16612
rect 11738 16560 11862 16612
rect 11862 16560 11990 16612
rect 12010 16888 12138 16940
rect 12138 16888 12262 16940
rect 12262 16888 12390 16940
rect 12010 16612 12390 16888
rect 12010 16560 12138 16612
rect 12138 16560 12262 16612
rect 12262 16560 12390 16612
rect 12410 16888 12538 16940
rect 12538 16888 12662 16940
rect 12662 16888 12790 16940
rect 12410 16612 12790 16888
rect 12410 16560 12538 16612
rect 12538 16560 12662 16612
rect 12662 16560 12790 16612
rect 12810 16888 12938 16940
rect 12938 16888 13062 16940
rect 13062 16888 13190 16940
rect 12810 16612 13190 16888
rect 12810 16560 12938 16612
rect 12938 16560 13062 16612
rect 13062 16560 13190 16612
rect 13210 16888 13338 16940
rect 13338 16888 13462 16940
rect 13462 16888 13590 16940
rect 13210 16612 13590 16888
rect 13210 16560 13338 16612
rect 13338 16560 13462 16612
rect 13462 16560 13590 16612
rect 13610 16888 13738 16940
rect 13738 16888 13862 16940
rect 13862 16888 13990 16940
rect 13610 16612 13990 16888
rect 13610 16560 13738 16612
rect 13738 16560 13862 16612
rect 13862 16560 13990 16612
rect 14010 16888 14138 16940
rect 14138 16888 14262 16940
rect 14262 16888 14390 16940
rect 14010 16612 14390 16888
rect 14010 16560 14138 16612
rect 14138 16560 14262 16612
rect 14262 16560 14390 16612
rect 14410 16888 14538 16940
rect 14538 16888 14662 16940
rect 14662 16888 14790 16940
rect 14410 16612 14790 16888
rect 14410 16560 14538 16612
rect 14538 16560 14662 16612
rect 14662 16560 14790 16612
rect 14810 16888 14938 16940
rect 14938 16888 15062 16940
rect 15062 16888 15190 16940
rect 14810 16612 15190 16888
rect 14810 16560 14938 16612
rect 14938 16560 15062 16612
rect 15062 16560 15190 16612
rect 15210 16888 15338 16940
rect 15338 16888 15462 16940
rect 15462 16888 15590 16940
rect 15210 16612 15590 16888
rect 15210 16560 15338 16612
rect 15338 16560 15462 16612
rect 15462 16560 15590 16612
rect 410 16488 538 16540
rect 538 16488 662 16540
rect 662 16488 790 16540
rect 410 16212 790 16488
rect 410 16160 538 16212
rect 538 16160 662 16212
rect 662 16160 790 16212
rect 810 16488 938 16540
rect 938 16488 1062 16540
rect 1062 16488 1190 16540
rect 810 16212 1190 16488
rect 810 16160 938 16212
rect 938 16160 1062 16212
rect 1062 16160 1190 16212
rect 1210 16488 1338 16540
rect 1338 16488 1462 16540
rect 1462 16488 1590 16540
rect 1210 16212 1590 16488
rect 1210 16160 1338 16212
rect 1338 16160 1462 16212
rect 1462 16160 1590 16212
rect 1610 16488 1738 16540
rect 1738 16488 1862 16540
rect 1862 16488 1990 16540
rect 1610 16212 1990 16488
rect 1610 16160 1738 16212
rect 1738 16160 1862 16212
rect 1862 16160 1990 16212
rect 2010 16488 2138 16540
rect 2138 16488 2262 16540
rect 2262 16488 2390 16540
rect 2010 16212 2390 16488
rect 2010 16160 2138 16212
rect 2138 16160 2262 16212
rect 2262 16160 2390 16212
rect 2410 16488 2538 16540
rect 2538 16488 2662 16540
rect 2662 16488 2790 16540
rect 2410 16212 2790 16488
rect 2410 16160 2538 16212
rect 2538 16160 2662 16212
rect 2662 16160 2790 16212
rect 2810 16488 2938 16540
rect 2938 16488 3062 16540
rect 3062 16488 3190 16540
rect 2810 16212 3190 16488
rect 2810 16160 2938 16212
rect 2938 16160 3062 16212
rect 3062 16160 3190 16212
rect 3210 16488 3338 16540
rect 3338 16488 3462 16540
rect 3462 16488 3590 16540
rect 3210 16212 3590 16488
rect 3210 16160 3338 16212
rect 3338 16160 3462 16212
rect 3462 16160 3590 16212
rect 3610 16488 3738 16540
rect 3738 16488 3862 16540
rect 3862 16488 3990 16540
rect 3610 16212 3990 16488
rect 3610 16160 3738 16212
rect 3738 16160 3862 16212
rect 3862 16160 3990 16212
rect 4010 16488 4138 16540
rect 4138 16488 4262 16540
rect 4262 16488 4390 16540
rect 4010 16212 4390 16488
rect 4010 16160 4138 16212
rect 4138 16160 4262 16212
rect 4262 16160 4390 16212
rect 4410 16488 4538 16540
rect 4538 16488 4662 16540
rect 4662 16488 4790 16540
rect 4410 16212 4790 16488
rect 4410 16160 4538 16212
rect 4538 16160 4662 16212
rect 4662 16160 4790 16212
rect 4810 16488 4938 16540
rect 4938 16488 5062 16540
rect 5062 16488 5190 16540
rect 4810 16212 5190 16488
rect 4810 16160 4938 16212
rect 4938 16160 5062 16212
rect 5062 16160 5190 16212
rect 5210 16488 5338 16540
rect 5338 16488 5462 16540
rect 5462 16488 5590 16540
rect 5210 16212 5590 16488
rect 5210 16160 5338 16212
rect 5338 16160 5462 16212
rect 5462 16160 5590 16212
rect 5610 16488 5738 16540
rect 5738 16488 5862 16540
rect 5862 16488 5990 16540
rect 5610 16212 5990 16488
rect 5610 16160 5738 16212
rect 5738 16160 5862 16212
rect 5862 16160 5990 16212
rect 6010 16488 6138 16540
rect 6138 16488 6262 16540
rect 6262 16488 6390 16540
rect 6010 16212 6390 16488
rect 6010 16160 6138 16212
rect 6138 16160 6262 16212
rect 6262 16160 6390 16212
rect 6410 16488 6538 16540
rect 6538 16488 6662 16540
rect 6662 16488 6790 16540
rect 6410 16212 6790 16488
rect 6410 16160 6538 16212
rect 6538 16160 6662 16212
rect 6662 16160 6790 16212
rect 6810 16488 6938 16540
rect 6938 16488 7062 16540
rect 7062 16488 7190 16540
rect 6810 16212 7190 16488
rect 6810 16160 6938 16212
rect 6938 16160 7062 16212
rect 7062 16160 7190 16212
rect 7210 16488 7338 16540
rect 7338 16488 7462 16540
rect 7462 16488 7590 16540
rect 7210 16212 7590 16488
rect 7210 16160 7338 16212
rect 7338 16160 7462 16212
rect 7462 16160 7590 16212
rect 7610 16488 7738 16540
rect 7738 16488 7862 16540
rect 7862 16488 7990 16540
rect 7610 16212 7990 16488
rect 7610 16160 7738 16212
rect 7738 16160 7862 16212
rect 7862 16160 7990 16212
rect 8010 16488 8138 16540
rect 8138 16488 8262 16540
rect 8262 16488 8390 16540
rect 8010 16212 8390 16488
rect 8010 16160 8138 16212
rect 8138 16160 8262 16212
rect 8262 16160 8390 16212
rect 8410 16488 8538 16540
rect 8538 16488 8662 16540
rect 8662 16488 8790 16540
rect 8410 16212 8790 16488
rect 8410 16160 8538 16212
rect 8538 16160 8662 16212
rect 8662 16160 8790 16212
rect 8810 16488 8938 16540
rect 8938 16488 9062 16540
rect 9062 16488 9190 16540
rect 8810 16212 9190 16488
rect 8810 16160 8938 16212
rect 8938 16160 9062 16212
rect 9062 16160 9190 16212
rect 9210 16488 9338 16540
rect 9338 16488 9462 16540
rect 9462 16488 9590 16540
rect 9210 16212 9590 16488
rect 9210 16160 9338 16212
rect 9338 16160 9462 16212
rect 9462 16160 9590 16212
rect 9610 16488 9738 16540
rect 9738 16488 9862 16540
rect 9862 16488 9990 16540
rect 9610 16212 9990 16488
rect 9610 16160 9738 16212
rect 9738 16160 9862 16212
rect 9862 16160 9990 16212
rect 10010 16488 10138 16540
rect 10138 16488 10262 16540
rect 10262 16488 10390 16540
rect 10010 16212 10390 16488
rect 10010 16160 10138 16212
rect 10138 16160 10262 16212
rect 10262 16160 10390 16212
rect 10410 16488 10538 16540
rect 10538 16488 10662 16540
rect 10662 16488 10790 16540
rect 10410 16212 10790 16488
rect 10410 16160 10538 16212
rect 10538 16160 10662 16212
rect 10662 16160 10790 16212
rect 10810 16488 10938 16540
rect 10938 16488 11062 16540
rect 11062 16488 11190 16540
rect 10810 16212 11190 16488
rect 10810 16160 10938 16212
rect 10938 16160 11062 16212
rect 11062 16160 11190 16212
rect 11210 16488 11338 16540
rect 11338 16488 11462 16540
rect 11462 16488 11590 16540
rect 11210 16212 11590 16488
rect 11210 16160 11338 16212
rect 11338 16160 11462 16212
rect 11462 16160 11590 16212
rect 11610 16488 11738 16540
rect 11738 16488 11862 16540
rect 11862 16488 11990 16540
rect 11610 16212 11990 16488
rect 11610 16160 11738 16212
rect 11738 16160 11862 16212
rect 11862 16160 11990 16212
rect 12010 16488 12138 16540
rect 12138 16488 12262 16540
rect 12262 16488 12390 16540
rect 12010 16212 12390 16488
rect 12010 16160 12138 16212
rect 12138 16160 12262 16212
rect 12262 16160 12390 16212
rect 12410 16488 12538 16540
rect 12538 16488 12662 16540
rect 12662 16488 12790 16540
rect 12410 16212 12790 16488
rect 12410 16160 12538 16212
rect 12538 16160 12662 16212
rect 12662 16160 12790 16212
rect 12810 16488 12938 16540
rect 12938 16488 13062 16540
rect 13062 16488 13190 16540
rect 12810 16212 13190 16488
rect 12810 16160 12938 16212
rect 12938 16160 13062 16212
rect 13062 16160 13190 16212
rect 13210 16488 13338 16540
rect 13338 16488 13462 16540
rect 13462 16488 13590 16540
rect 13210 16212 13590 16488
rect 13210 16160 13338 16212
rect 13338 16160 13462 16212
rect 13462 16160 13590 16212
rect 13610 16488 13738 16540
rect 13738 16488 13862 16540
rect 13862 16488 13990 16540
rect 13610 16212 13990 16488
rect 13610 16160 13738 16212
rect 13738 16160 13862 16212
rect 13862 16160 13990 16212
rect 14010 16488 14138 16540
rect 14138 16488 14262 16540
rect 14262 16488 14390 16540
rect 14010 16212 14390 16488
rect 14010 16160 14138 16212
rect 14138 16160 14262 16212
rect 14262 16160 14390 16212
rect 14410 16488 14538 16540
rect 14538 16488 14662 16540
rect 14662 16488 14790 16540
rect 14410 16212 14790 16488
rect 14410 16160 14538 16212
rect 14538 16160 14662 16212
rect 14662 16160 14790 16212
rect 14810 16488 14938 16540
rect 14938 16488 15062 16540
rect 15062 16488 15190 16540
rect 14810 16212 15190 16488
rect 14810 16160 14938 16212
rect 14938 16160 15062 16212
rect 15062 16160 15190 16212
rect 15210 16488 15338 16540
rect 15338 16488 15462 16540
rect 15462 16488 15590 16540
rect 15210 16212 15590 16488
rect 15210 16160 15338 16212
rect 15338 16160 15462 16212
rect 15462 16160 15590 16212
rect 410 16088 538 16140
rect 538 16088 662 16140
rect 662 16088 790 16140
rect 410 15812 790 16088
rect 410 15760 538 15812
rect 538 15760 662 15812
rect 662 15760 790 15812
rect 810 16088 938 16140
rect 938 16088 1062 16140
rect 1062 16088 1190 16140
rect 810 15812 1190 16088
rect 810 15760 938 15812
rect 938 15760 1062 15812
rect 1062 15760 1190 15812
rect 1210 16088 1338 16140
rect 1338 16088 1462 16140
rect 1462 16088 1590 16140
rect 1210 15812 1590 16088
rect 1210 15760 1338 15812
rect 1338 15760 1462 15812
rect 1462 15760 1590 15812
rect 1610 16088 1738 16140
rect 1738 16088 1862 16140
rect 1862 16088 1990 16140
rect 1610 15812 1990 16088
rect 1610 15760 1738 15812
rect 1738 15760 1862 15812
rect 1862 15760 1990 15812
rect 2010 16088 2138 16140
rect 2138 16088 2262 16140
rect 2262 16088 2390 16140
rect 2010 15812 2390 16088
rect 2010 15760 2138 15812
rect 2138 15760 2262 15812
rect 2262 15760 2390 15812
rect 2410 16088 2538 16140
rect 2538 16088 2662 16140
rect 2662 16088 2790 16140
rect 2410 15812 2790 16088
rect 2410 15760 2538 15812
rect 2538 15760 2662 15812
rect 2662 15760 2790 15812
rect 2810 16088 2938 16140
rect 2938 16088 3062 16140
rect 3062 16088 3190 16140
rect 2810 15812 3190 16088
rect 2810 15760 2938 15812
rect 2938 15760 3062 15812
rect 3062 15760 3190 15812
rect 3210 16088 3338 16140
rect 3338 16088 3462 16140
rect 3462 16088 3590 16140
rect 3210 15812 3590 16088
rect 3210 15760 3338 15812
rect 3338 15760 3462 15812
rect 3462 15760 3590 15812
rect 3610 16088 3738 16140
rect 3738 16088 3862 16140
rect 3862 16088 3990 16140
rect 3610 15812 3990 16088
rect 3610 15760 3738 15812
rect 3738 15760 3862 15812
rect 3862 15760 3990 15812
rect 4010 16088 4138 16140
rect 4138 16088 4262 16140
rect 4262 16088 4390 16140
rect 4010 15812 4390 16088
rect 4010 15760 4138 15812
rect 4138 15760 4262 15812
rect 4262 15760 4390 15812
rect 4410 16088 4538 16140
rect 4538 16088 4662 16140
rect 4662 16088 4790 16140
rect 4410 15812 4790 16088
rect 4410 15760 4538 15812
rect 4538 15760 4662 15812
rect 4662 15760 4790 15812
rect 4810 16088 4938 16140
rect 4938 16088 5062 16140
rect 5062 16088 5190 16140
rect 4810 15812 5190 16088
rect 4810 15760 4938 15812
rect 4938 15760 5062 15812
rect 5062 15760 5190 15812
rect 5210 16088 5338 16140
rect 5338 16088 5462 16140
rect 5462 16088 5590 16140
rect 5210 15812 5590 16088
rect 5210 15760 5338 15812
rect 5338 15760 5462 15812
rect 5462 15760 5590 15812
rect 5610 16088 5738 16140
rect 5738 16088 5862 16140
rect 5862 16088 5990 16140
rect 5610 15812 5990 16088
rect 5610 15760 5738 15812
rect 5738 15760 5862 15812
rect 5862 15760 5990 15812
rect 6010 16088 6138 16140
rect 6138 16088 6262 16140
rect 6262 16088 6390 16140
rect 6010 15812 6390 16088
rect 6010 15760 6138 15812
rect 6138 15760 6262 15812
rect 6262 15760 6390 15812
rect 6410 16088 6538 16140
rect 6538 16088 6662 16140
rect 6662 16088 6790 16140
rect 6410 15812 6790 16088
rect 6410 15760 6538 15812
rect 6538 15760 6662 15812
rect 6662 15760 6790 15812
rect 6810 16088 6938 16140
rect 6938 16088 7062 16140
rect 7062 16088 7190 16140
rect 6810 15812 7190 16088
rect 6810 15760 6938 15812
rect 6938 15760 7062 15812
rect 7062 15760 7190 15812
rect 7210 16088 7338 16140
rect 7338 16088 7462 16140
rect 7462 16088 7590 16140
rect 7210 15812 7590 16088
rect 7210 15760 7338 15812
rect 7338 15760 7462 15812
rect 7462 15760 7590 15812
rect 7610 16088 7738 16140
rect 7738 16088 7862 16140
rect 7862 16088 7990 16140
rect 7610 15812 7990 16088
rect 7610 15760 7738 15812
rect 7738 15760 7862 15812
rect 7862 15760 7990 15812
rect 8010 16088 8138 16140
rect 8138 16088 8262 16140
rect 8262 16088 8390 16140
rect 8010 15812 8390 16088
rect 8010 15760 8138 15812
rect 8138 15760 8262 15812
rect 8262 15760 8390 15812
rect 8410 16088 8538 16140
rect 8538 16088 8662 16140
rect 8662 16088 8790 16140
rect 8410 15812 8790 16088
rect 8410 15760 8538 15812
rect 8538 15760 8662 15812
rect 8662 15760 8790 15812
rect 8810 16088 8938 16140
rect 8938 16088 9062 16140
rect 9062 16088 9190 16140
rect 8810 15812 9190 16088
rect 8810 15760 8938 15812
rect 8938 15760 9062 15812
rect 9062 15760 9190 15812
rect 9210 16088 9338 16140
rect 9338 16088 9462 16140
rect 9462 16088 9590 16140
rect 9210 15812 9590 16088
rect 9210 15760 9338 15812
rect 9338 15760 9462 15812
rect 9462 15760 9590 15812
rect 9610 16088 9738 16140
rect 9738 16088 9862 16140
rect 9862 16088 9990 16140
rect 9610 15812 9990 16088
rect 9610 15760 9738 15812
rect 9738 15760 9862 15812
rect 9862 15760 9990 15812
rect 10010 16088 10138 16140
rect 10138 16088 10262 16140
rect 10262 16088 10390 16140
rect 10010 15812 10390 16088
rect 10010 15760 10138 15812
rect 10138 15760 10262 15812
rect 10262 15760 10390 15812
rect 10410 16088 10538 16140
rect 10538 16088 10662 16140
rect 10662 16088 10790 16140
rect 10410 15812 10790 16088
rect 10410 15760 10538 15812
rect 10538 15760 10662 15812
rect 10662 15760 10790 15812
rect 10810 16088 10938 16140
rect 10938 16088 11062 16140
rect 11062 16088 11190 16140
rect 10810 15812 11190 16088
rect 10810 15760 10938 15812
rect 10938 15760 11062 15812
rect 11062 15760 11190 15812
rect 11210 16088 11338 16140
rect 11338 16088 11462 16140
rect 11462 16088 11590 16140
rect 11210 15812 11590 16088
rect 11210 15760 11338 15812
rect 11338 15760 11462 15812
rect 11462 15760 11590 15812
rect 11610 16088 11738 16140
rect 11738 16088 11862 16140
rect 11862 16088 11990 16140
rect 11610 15812 11990 16088
rect 11610 15760 11738 15812
rect 11738 15760 11862 15812
rect 11862 15760 11990 15812
rect 12010 16088 12138 16140
rect 12138 16088 12262 16140
rect 12262 16088 12390 16140
rect 12010 15812 12390 16088
rect 12010 15760 12138 15812
rect 12138 15760 12262 15812
rect 12262 15760 12390 15812
rect 12410 16088 12538 16140
rect 12538 16088 12662 16140
rect 12662 16088 12790 16140
rect 12410 15812 12790 16088
rect 12410 15760 12538 15812
rect 12538 15760 12662 15812
rect 12662 15760 12790 15812
rect 12810 16088 12938 16140
rect 12938 16088 13062 16140
rect 13062 16088 13190 16140
rect 12810 15812 13190 16088
rect 12810 15760 12938 15812
rect 12938 15760 13062 15812
rect 13062 15760 13190 15812
rect 13210 16088 13338 16140
rect 13338 16088 13462 16140
rect 13462 16088 13590 16140
rect 13210 15812 13590 16088
rect 13210 15760 13338 15812
rect 13338 15760 13462 15812
rect 13462 15760 13590 15812
rect 13610 16088 13738 16140
rect 13738 16088 13862 16140
rect 13862 16088 13990 16140
rect 13610 15812 13990 16088
rect 13610 15760 13738 15812
rect 13738 15760 13862 15812
rect 13862 15760 13990 15812
rect 14010 16088 14138 16140
rect 14138 16088 14262 16140
rect 14262 16088 14390 16140
rect 14010 15812 14390 16088
rect 14010 15760 14138 15812
rect 14138 15760 14262 15812
rect 14262 15760 14390 15812
rect 14410 16088 14538 16140
rect 14538 16088 14662 16140
rect 14662 16088 14790 16140
rect 14410 15812 14790 16088
rect 14410 15760 14538 15812
rect 14538 15760 14662 15812
rect 14662 15760 14790 15812
rect 14810 16088 14938 16140
rect 14938 16088 15062 16140
rect 15062 16088 15190 16140
rect 14810 15812 15190 16088
rect 14810 15760 14938 15812
rect 14938 15760 15062 15812
rect 15062 15760 15190 15812
rect 15210 16088 15338 16140
rect 15338 16088 15462 16140
rect 15462 16088 15590 16140
rect 15210 15812 15590 16088
rect 15210 15760 15338 15812
rect 15338 15760 15462 15812
rect 15462 15760 15590 15812
rect 410 15688 538 15740
rect 538 15688 662 15740
rect 662 15688 790 15740
rect 410 15412 790 15688
rect 410 15360 538 15412
rect 538 15360 662 15412
rect 662 15360 790 15412
rect 810 15688 938 15740
rect 938 15688 1062 15740
rect 1062 15688 1190 15740
rect 810 15412 1190 15688
rect 810 15360 938 15412
rect 938 15360 1062 15412
rect 1062 15360 1190 15412
rect 1210 15688 1338 15740
rect 1338 15688 1462 15740
rect 1462 15688 1590 15740
rect 1210 15412 1590 15688
rect 1210 15360 1338 15412
rect 1338 15360 1462 15412
rect 1462 15360 1590 15412
rect 1610 15688 1738 15740
rect 1738 15688 1862 15740
rect 1862 15688 1990 15740
rect 1610 15412 1990 15688
rect 1610 15360 1738 15412
rect 1738 15360 1862 15412
rect 1862 15360 1990 15412
rect 2010 15688 2138 15740
rect 2138 15688 2262 15740
rect 2262 15688 2390 15740
rect 2010 15412 2390 15688
rect 2010 15360 2138 15412
rect 2138 15360 2262 15412
rect 2262 15360 2390 15412
rect 2410 15688 2538 15740
rect 2538 15688 2662 15740
rect 2662 15688 2790 15740
rect 2410 15412 2790 15688
rect 2410 15360 2538 15412
rect 2538 15360 2662 15412
rect 2662 15360 2790 15412
rect 2810 15688 2938 15740
rect 2938 15688 3062 15740
rect 3062 15688 3190 15740
rect 2810 15412 3190 15688
rect 2810 15360 2938 15412
rect 2938 15360 3062 15412
rect 3062 15360 3190 15412
rect 3210 15688 3338 15740
rect 3338 15688 3462 15740
rect 3462 15688 3590 15740
rect 3210 15412 3590 15688
rect 3210 15360 3338 15412
rect 3338 15360 3462 15412
rect 3462 15360 3590 15412
rect 3610 15688 3738 15740
rect 3738 15688 3862 15740
rect 3862 15688 3990 15740
rect 3610 15412 3990 15688
rect 3610 15360 3738 15412
rect 3738 15360 3862 15412
rect 3862 15360 3990 15412
rect 4010 15688 4138 15740
rect 4138 15688 4262 15740
rect 4262 15688 4390 15740
rect 4010 15412 4390 15688
rect 4010 15360 4138 15412
rect 4138 15360 4262 15412
rect 4262 15360 4390 15412
rect 4410 15688 4538 15740
rect 4538 15688 4662 15740
rect 4662 15688 4790 15740
rect 4410 15412 4790 15688
rect 4410 15360 4538 15412
rect 4538 15360 4662 15412
rect 4662 15360 4790 15412
rect 4810 15688 4938 15740
rect 4938 15688 5062 15740
rect 5062 15688 5190 15740
rect 4810 15412 5190 15688
rect 4810 15360 4938 15412
rect 4938 15360 5062 15412
rect 5062 15360 5190 15412
rect 5210 15688 5338 15740
rect 5338 15688 5462 15740
rect 5462 15688 5590 15740
rect 5210 15412 5590 15688
rect 5210 15360 5338 15412
rect 5338 15360 5462 15412
rect 5462 15360 5590 15412
rect 5610 15688 5738 15740
rect 5738 15688 5862 15740
rect 5862 15688 5990 15740
rect 5610 15412 5990 15688
rect 5610 15360 5738 15412
rect 5738 15360 5862 15412
rect 5862 15360 5990 15412
rect 6010 15688 6138 15740
rect 6138 15688 6262 15740
rect 6262 15688 6390 15740
rect 6010 15412 6390 15688
rect 6010 15360 6138 15412
rect 6138 15360 6262 15412
rect 6262 15360 6390 15412
rect 6410 15688 6538 15740
rect 6538 15688 6662 15740
rect 6662 15688 6790 15740
rect 6410 15412 6790 15688
rect 6410 15360 6538 15412
rect 6538 15360 6662 15412
rect 6662 15360 6790 15412
rect 6810 15688 6938 15740
rect 6938 15688 7062 15740
rect 7062 15688 7190 15740
rect 6810 15412 7190 15688
rect 6810 15360 6938 15412
rect 6938 15360 7062 15412
rect 7062 15360 7190 15412
rect 7210 15688 7338 15740
rect 7338 15688 7462 15740
rect 7462 15688 7590 15740
rect 7210 15412 7590 15688
rect 7210 15360 7338 15412
rect 7338 15360 7462 15412
rect 7462 15360 7590 15412
rect 7610 15688 7738 15740
rect 7738 15688 7862 15740
rect 7862 15688 7990 15740
rect 7610 15412 7990 15688
rect 7610 15360 7738 15412
rect 7738 15360 7862 15412
rect 7862 15360 7990 15412
rect 8010 15688 8138 15740
rect 8138 15688 8262 15740
rect 8262 15688 8390 15740
rect 8010 15412 8390 15688
rect 8010 15360 8138 15412
rect 8138 15360 8262 15412
rect 8262 15360 8390 15412
rect 8410 15688 8538 15740
rect 8538 15688 8662 15740
rect 8662 15688 8790 15740
rect 8410 15412 8790 15688
rect 8410 15360 8538 15412
rect 8538 15360 8662 15412
rect 8662 15360 8790 15412
rect 8810 15688 8938 15740
rect 8938 15688 9062 15740
rect 9062 15688 9190 15740
rect 8810 15412 9190 15688
rect 8810 15360 8938 15412
rect 8938 15360 9062 15412
rect 9062 15360 9190 15412
rect 9210 15688 9338 15740
rect 9338 15688 9462 15740
rect 9462 15688 9590 15740
rect 9210 15412 9590 15688
rect 9210 15360 9338 15412
rect 9338 15360 9462 15412
rect 9462 15360 9590 15412
rect 9610 15688 9738 15740
rect 9738 15688 9862 15740
rect 9862 15688 9990 15740
rect 9610 15412 9990 15688
rect 9610 15360 9738 15412
rect 9738 15360 9862 15412
rect 9862 15360 9990 15412
rect 10010 15688 10138 15740
rect 10138 15688 10262 15740
rect 10262 15688 10390 15740
rect 10010 15412 10390 15688
rect 10010 15360 10138 15412
rect 10138 15360 10262 15412
rect 10262 15360 10390 15412
rect 10410 15688 10538 15740
rect 10538 15688 10662 15740
rect 10662 15688 10790 15740
rect 10410 15412 10790 15688
rect 10410 15360 10538 15412
rect 10538 15360 10662 15412
rect 10662 15360 10790 15412
rect 10810 15688 10938 15740
rect 10938 15688 11062 15740
rect 11062 15688 11190 15740
rect 10810 15412 11190 15688
rect 10810 15360 10938 15412
rect 10938 15360 11062 15412
rect 11062 15360 11190 15412
rect 11210 15688 11338 15740
rect 11338 15688 11462 15740
rect 11462 15688 11590 15740
rect 11210 15412 11590 15688
rect 11210 15360 11338 15412
rect 11338 15360 11462 15412
rect 11462 15360 11590 15412
rect 11610 15688 11738 15740
rect 11738 15688 11862 15740
rect 11862 15688 11990 15740
rect 11610 15412 11990 15688
rect 11610 15360 11738 15412
rect 11738 15360 11862 15412
rect 11862 15360 11990 15412
rect 12010 15688 12138 15740
rect 12138 15688 12262 15740
rect 12262 15688 12390 15740
rect 12010 15412 12390 15688
rect 12010 15360 12138 15412
rect 12138 15360 12262 15412
rect 12262 15360 12390 15412
rect 12410 15688 12538 15740
rect 12538 15688 12662 15740
rect 12662 15688 12790 15740
rect 12410 15412 12790 15688
rect 12410 15360 12538 15412
rect 12538 15360 12662 15412
rect 12662 15360 12790 15412
rect 12810 15688 12938 15740
rect 12938 15688 13062 15740
rect 13062 15688 13190 15740
rect 12810 15412 13190 15688
rect 12810 15360 12938 15412
rect 12938 15360 13062 15412
rect 13062 15360 13190 15412
rect 13210 15688 13338 15740
rect 13338 15688 13462 15740
rect 13462 15688 13590 15740
rect 13210 15412 13590 15688
rect 13210 15360 13338 15412
rect 13338 15360 13462 15412
rect 13462 15360 13590 15412
rect 13610 15688 13738 15740
rect 13738 15688 13862 15740
rect 13862 15688 13990 15740
rect 13610 15412 13990 15688
rect 13610 15360 13738 15412
rect 13738 15360 13862 15412
rect 13862 15360 13990 15412
rect 14010 15688 14138 15740
rect 14138 15688 14262 15740
rect 14262 15688 14390 15740
rect 14010 15412 14390 15688
rect 14010 15360 14138 15412
rect 14138 15360 14262 15412
rect 14262 15360 14390 15412
rect 14410 15688 14538 15740
rect 14538 15688 14662 15740
rect 14662 15688 14790 15740
rect 14410 15412 14790 15688
rect 14410 15360 14538 15412
rect 14538 15360 14662 15412
rect 14662 15360 14790 15412
rect 14810 15688 14938 15740
rect 14938 15688 15062 15740
rect 15062 15688 15190 15740
rect 14810 15412 15190 15688
rect 14810 15360 14938 15412
rect 14938 15360 15062 15412
rect 15062 15360 15190 15412
rect 15210 15688 15338 15740
rect 15338 15688 15462 15740
rect 15462 15688 15590 15740
rect 15210 15412 15590 15688
rect 15210 15360 15338 15412
rect 15338 15360 15462 15412
rect 15462 15360 15590 15412
rect 410 15288 538 15340
rect 538 15288 662 15340
rect 662 15288 790 15340
rect 410 15012 790 15288
rect 410 14960 538 15012
rect 538 14960 662 15012
rect 662 14960 790 15012
rect 810 15288 938 15340
rect 938 15288 1062 15340
rect 1062 15288 1190 15340
rect 810 15012 1190 15288
rect 810 14960 938 15012
rect 938 14960 1062 15012
rect 1062 14960 1190 15012
rect 1210 15288 1338 15340
rect 1338 15288 1462 15340
rect 1462 15288 1590 15340
rect 1210 15012 1590 15288
rect 1210 14960 1338 15012
rect 1338 14960 1462 15012
rect 1462 14960 1590 15012
rect 1610 15288 1738 15340
rect 1738 15288 1862 15340
rect 1862 15288 1990 15340
rect 1610 15012 1990 15288
rect 1610 14960 1738 15012
rect 1738 14960 1862 15012
rect 1862 14960 1990 15012
rect 2010 15288 2138 15340
rect 2138 15288 2262 15340
rect 2262 15288 2390 15340
rect 2010 15012 2390 15288
rect 2010 14960 2138 15012
rect 2138 14960 2262 15012
rect 2262 14960 2390 15012
rect 2410 15288 2538 15340
rect 2538 15288 2662 15340
rect 2662 15288 2790 15340
rect 2410 15012 2790 15288
rect 2410 14960 2538 15012
rect 2538 14960 2662 15012
rect 2662 14960 2790 15012
rect 2810 15288 2938 15340
rect 2938 15288 3062 15340
rect 3062 15288 3190 15340
rect 2810 15012 3190 15288
rect 2810 14960 2938 15012
rect 2938 14960 3062 15012
rect 3062 14960 3190 15012
rect 3210 15288 3338 15340
rect 3338 15288 3462 15340
rect 3462 15288 3590 15340
rect 3210 15012 3590 15288
rect 3210 14960 3338 15012
rect 3338 14960 3462 15012
rect 3462 14960 3590 15012
rect 3610 15288 3738 15340
rect 3738 15288 3862 15340
rect 3862 15288 3990 15340
rect 3610 15012 3990 15288
rect 3610 14960 3738 15012
rect 3738 14960 3862 15012
rect 3862 14960 3990 15012
rect 4010 15288 4138 15340
rect 4138 15288 4262 15340
rect 4262 15288 4390 15340
rect 4010 15012 4390 15288
rect 4010 14960 4138 15012
rect 4138 14960 4262 15012
rect 4262 14960 4390 15012
rect 4410 15288 4538 15340
rect 4538 15288 4662 15340
rect 4662 15288 4790 15340
rect 4410 15012 4790 15288
rect 4410 14960 4538 15012
rect 4538 14960 4662 15012
rect 4662 14960 4790 15012
rect 4810 15288 4938 15340
rect 4938 15288 5062 15340
rect 5062 15288 5190 15340
rect 4810 15012 5190 15288
rect 4810 14960 4938 15012
rect 4938 14960 5062 15012
rect 5062 14960 5190 15012
rect 5210 15288 5338 15340
rect 5338 15288 5462 15340
rect 5462 15288 5590 15340
rect 5210 15012 5590 15288
rect 5210 14960 5338 15012
rect 5338 14960 5462 15012
rect 5462 14960 5590 15012
rect 5610 15288 5738 15340
rect 5738 15288 5862 15340
rect 5862 15288 5990 15340
rect 5610 15012 5990 15288
rect 5610 14960 5738 15012
rect 5738 14960 5862 15012
rect 5862 14960 5990 15012
rect 6010 15288 6138 15340
rect 6138 15288 6262 15340
rect 6262 15288 6390 15340
rect 6010 15012 6390 15288
rect 6010 14960 6138 15012
rect 6138 14960 6262 15012
rect 6262 14960 6390 15012
rect 6410 15288 6538 15340
rect 6538 15288 6662 15340
rect 6662 15288 6790 15340
rect 6410 15012 6790 15288
rect 6410 14960 6538 15012
rect 6538 14960 6662 15012
rect 6662 14960 6790 15012
rect 6810 15288 6938 15340
rect 6938 15288 7062 15340
rect 7062 15288 7190 15340
rect 6810 15012 7190 15288
rect 6810 14960 6938 15012
rect 6938 14960 7062 15012
rect 7062 14960 7190 15012
rect 7210 15288 7338 15340
rect 7338 15288 7462 15340
rect 7462 15288 7590 15340
rect 7210 15012 7590 15288
rect 7210 14960 7338 15012
rect 7338 14960 7462 15012
rect 7462 14960 7590 15012
rect 7610 15288 7738 15340
rect 7738 15288 7862 15340
rect 7862 15288 7990 15340
rect 7610 15012 7990 15288
rect 7610 14960 7738 15012
rect 7738 14960 7862 15012
rect 7862 14960 7990 15012
rect 8010 15288 8138 15340
rect 8138 15288 8262 15340
rect 8262 15288 8390 15340
rect 8010 15012 8390 15288
rect 8010 14960 8138 15012
rect 8138 14960 8262 15012
rect 8262 14960 8390 15012
rect 8410 15288 8538 15340
rect 8538 15288 8662 15340
rect 8662 15288 8790 15340
rect 8410 15012 8790 15288
rect 8410 14960 8538 15012
rect 8538 14960 8662 15012
rect 8662 14960 8790 15012
rect 8810 15288 8938 15340
rect 8938 15288 9062 15340
rect 9062 15288 9190 15340
rect 8810 15012 9190 15288
rect 8810 14960 8938 15012
rect 8938 14960 9062 15012
rect 9062 14960 9190 15012
rect 9210 15288 9338 15340
rect 9338 15288 9462 15340
rect 9462 15288 9590 15340
rect 9210 15012 9590 15288
rect 9210 14960 9338 15012
rect 9338 14960 9462 15012
rect 9462 14960 9590 15012
rect 9610 15288 9738 15340
rect 9738 15288 9862 15340
rect 9862 15288 9990 15340
rect 9610 15012 9990 15288
rect 9610 14960 9738 15012
rect 9738 14960 9862 15012
rect 9862 14960 9990 15012
rect 10010 15288 10138 15340
rect 10138 15288 10262 15340
rect 10262 15288 10390 15340
rect 10010 15012 10390 15288
rect 10010 14960 10138 15012
rect 10138 14960 10262 15012
rect 10262 14960 10390 15012
rect 10410 15288 10538 15340
rect 10538 15288 10662 15340
rect 10662 15288 10790 15340
rect 10410 15012 10790 15288
rect 10410 14960 10538 15012
rect 10538 14960 10662 15012
rect 10662 14960 10790 15012
rect 10810 15288 10938 15340
rect 10938 15288 11062 15340
rect 11062 15288 11190 15340
rect 10810 15012 11190 15288
rect 10810 14960 10938 15012
rect 10938 14960 11062 15012
rect 11062 14960 11190 15012
rect 11210 15288 11338 15340
rect 11338 15288 11462 15340
rect 11462 15288 11590 15340
rect 11210 15012 11590 15288
rect 11210 14960 11338 15012
rect 11338 14960 11462 15012
rect 11462 14960 11590 15012
rect 11610 15288 11738 15340
rect 11738 15288 11862 15340
rect 11862 15288 11990 15340
rect 11610 15012 11990 15288
rect 11610 14960 11738 15012
rect 11738 14960 11862 15012
rect 11862 14960 11990 15012
rect 12010 15288 12138 15340
rect 12138 15288 12262 15340
rect 12262 15288 12390 15340
rect 12010 15012 12390 15288
rect 12010 14960 12138 15012
rect 12138 14960 12262 15012
rect 12262 14960 12390 15012
rect 12410 15288 12538 15340
rect 12538 15288 12662 15340
rect 12662 15288 12790 15340
rect 12410 15012 12790 15288
rect 12410 14960 12538 15012
rect 12538 14960 12662 15012
rect 12662 14960 12790 15012
rect 12810 15288 12938 15340
rect 12938 15288 13062 15340
rect 13062 15288 13190 15340
rect 12810 15012 13190 15288
rect 12810 14960 12938 15012
rect 12938 14960 13062 15012
rect 13062 14960 13190 15012
rect 13210 15288 13338 15340
rect 13338 15288 13462 15340
rect 13462 15288 13590 15340
rect 13210 15012 13590 15288
rect 13210 14960 13338 15012
rect 13338 14960 13462 15012
rect 13462 14960 13590 15012
rect 13610 15288 13738 15340
rect 13738 15288 13862 15340
rect 13862 15288 13990 15340
rect 13610 15012 13990 15288
rect 13610 14960 13738 15012
rect 13738 14960 13862 15012
rect 13862 14960 13990 15012
rect 14010 15288 14138 15340
rect 14138 15288 14262 15340
rect 14262 15288 14390 15340
rect 14010 15012 14390 15288
rect 14010 14960 14138 15012
rect 14138 14960 14262 15012
rect 14262 14960 14390 15012
rect 14410 15288 14538 15340
rect 14538 15288 14662 15340
rect 14662 15288 14790 15340
rect 14410 15012 14790 15288
rect 14410 14960 14538 15012
rect 14538 14960 14662 15012
rect 14662 14960 14790 15012
rect 14810 15288 14938 15340
rect 14938 15288 15062 15340
rect 15062 15288 15190 15340
rect 14810 15012 15190 15288
rect 14810 14960 14938 15012
rect 14938 14960 15062 15012
rect 15062 14960 15190 15012
rect 15210 15288 15338 15340
rect 15338 15288 15462 15340
rect 15462 15288 15590 15340
rect 15210 15012 15590 15288
rect 15210 14960 15338 15012
rect 15338 14960 15462 15012
rect 15462 14960 15590 15012
rect 410 14888 538 14940
rect 538 14888 662 14940
rect 662 14888 790 14940
rect 410 14612 790 14888
rect 410 14560 538 14612
rect 538 14560 662 14612
rect 662 14560 790 14612
rect 810 14888 938 14940
rect 938 14888 1062 14940
rect 1062 14888 1190 14940
rect 810 14612 1190 14888
rect 810 14560 938 14612
rect 938 14560 1062 14612
rect 1062 14560 1190 14612
rect 1210 14888 1338 14940
rect 1338 14888 1462 14940
rect 1462 14888 1590 14940
rect 1210 14612 1590 14888
rect 1210 14560 1338 14612
rect 1338 14560 1462 14612
rect 1462 14560 1590 14612
rect 1610 14888 1738 14940
rect 1738 14888 1862 14940
rect 1862 14888 1990 14940
rect 1610 14612 1990 14888
rect 1610 14560 1738 14612
rect 1738 14560 1862 14612
rect 1862 14560 1990 14612
rect 2010 14888 2138 14940
rect 2138 14888 2262 14940
rect 2262 14888 2390 14940
rect 2010 14612 2390 14888
rect 2010 14560 2138 14612
rect 2138 14560 2262 14612
rect 2262 14560 2390 14612
rect 2410 14888 2538 14940
rect 2538 14888 2662 14940
rect 2662 14888 2790 14940
rect 2410 14612 2790 14888
rect 2410 14560 2538 14612
rect 2538 14560 2662 14612
rect 2662 14560 2790 14612
rect 2810 14888 2938 14940
rect 2938 14888 3062 14940
rect 3062 14888 3190 14940
rect 2810 14612 3190 14888
rect 2810 14560 2938 14612
rect 2938 14560 3062 14612
rect 3062 14560 3190 14612
rect 3210 14888 3338 14940
rect 3338 14888 3462 14940
rect 3462 14888 3590 14940
rect 3210 14612 3590 14888
rect 3210 14560 3338 14612
rect 3338 14560 3462 14612
rect 3462 14560 3590 14612
rect 3610 14888 3738 14940
rect 3738 14888 3862 14940
rect 3862 14888 3990 14940
rect 3610 14612 3990 14888
rect 3610 14560 3738 14612
rect 3738 14560 3862 14612
rect 3862 14560 3990 14612
rect 4010 14888 4138 14940
rect 4138 14888 4262 14940
rect 4262 14888 4390 14940
rect 4010 14612 4390 14888
rect 4010 14560 4138 14612
rect 4138 14560 4262 14612
rect 4262 14560 4390 14612
rect 4410 14888 4538 14940
rect 4538 14888 4662 14940
rect 4662 14888 4790 14940
rect 4410 14612 4790 14888
rect 4410 14560 4538 14612
rect 4538 14560 4662 14612
rect 4662 14560 4790 14612
rect 4810 14888 4938 14940
rect 4938 14888 5062 14940
rect 5062 14888 5190 14940
rect 4810 14612 5190 14888
rect 4810 14560 4938 14612
rect 4938 14560 5062 14612
rect 5062 14560 5190 14612
rect 5210 14888 5338 14940
rect 5338 14888 5462 14940
rect 5462 14888 5590 14940
rect 5210 14612 5590 14888
rect 5210 14560 5338 14612
rect 5338 14560 5462 14612
rect 5462 14560 5590 14612
rect 5610 14888 5738 14940
rect 5738 14888 5862 14940
rect 5862 14888 5990 14940
rect 5610 14612 5990 14888
rect 5610 14560 5738 14612
rect 5738 14560 5862 14612
rect 5862 14560 5990 14612
rect 6010 14888 6138 14940
rect 6138 14888 6262 14940
rect 6262 14888 6390 14940
rect 6010 14612 6390 14888
rect 6010 14560 6138 14612
rect 6138 14560 6262 14612
rect 6262 14560 6390 14612
rect 6410 14888 6538 14940
rect 6538 14888 6662 14940
rect 6662 14888 6790 14940
rect 6410 14612 6790 14888
rect 6410 14560 6538 14612
rect 6538 14560 6662 14612
rect 6662 14560 6790 14612
rect 6810 14888 6938 14940
rect 6938 14888 7062 14940
rect 7062 14888 7190 14940
rect 6810 14612 7190 14888
rect 6810 14560 6938 14612
rect 6938 14560 7062 14612
rect 7062 14560 7190 14612
rect 7210 14888 7338 14940
rect 7338 14888 7462 14940
rect 7462 14888 7590 14940
rect 7210 14612 7590 14888
rect 7210 14560 7338 14612
rect 7338 14560 7462 14612
rect 7462 14560 7590 14612
rect 7610 14888 7738 14940
rect 7738 14888 7862 14940
rect 7862 14888 7990 14940
rect 7610 14612 7990 14888
rect 7610 14560 7738 14612
rect 7738 14560 7862 14612
rect 7862 14560 7990 14612
rect 8010 14888 8138 14940
rect 8138 14888 8262 14940
rect 8262 14888 8390 14940
rect 8010 14612 8390 14888
rect 8010 14560 8138 14612
rect 8138 14560 8262 14612
rect 8262 14560 8390 14612
rect 8410 14888 8538 14940
rect 8538 14888 8662 14940
rect 8662 14888 8790 14940
rect 8410 14612 8790 14888
rect 8410 14560 8538 14612
rect 8538 14560 8662 14612
rect 8662 14560 8790 14612
rect 8810 14888 8938 14940
rect 8938 14888 9062 14940
rect 9062 14888 9190 14940
rect 8810 14612 9190 14888
rect 8810 14560 8938 14612
rect 8938 14560 9062 14612
rect 9062 14560 9190 14612
rect 9210 14888 9338 14940
rect 9338 14888 9462 14940
rect 9462 14888 9590 14940
rect 9210 14612 9590 14888
rect 9210 14560 9338 14612
rect 9338 14560 9462 14612
rect 9462 14560 9590 14612
rect 9610 14888 9738 14940
rect 9738 14888 9862 14940
rect 9862 14888 9990 14940
rect 9610 14612 9990 14888
rect 9610 14560 9738 14612
rect 9738 14560 9862 14612
rect 9862 14560 9990 14612
rect 10010 14888 10138 14940
rect 10138 14888 10262 14940
rect 10262 14888 10390 14940
rect 10010 14612 10390 14888
rect 10010 14560 10138 14612
rect 10138 14560 10262 14612
rect 10262 14560 10390 14612
rect 10410 14888 10538 14940
rect 10538 14888 10662 14940
rect 10662 14888 10790 14940
rect 10410 14612 10790 14888
rect 10410 14560 10538 14612
rect 10538 14560 10662 14612
rect 10662 14560 10790 14612
rect 10810 14888 10938 14940
rect 10938 14888 11062 14940
rect 11062 14888 11190 14940
rect 10810 14612 11190 14888
rect 10810 14560 10938 14612
rect 10938 14560 11062 14612
rect 11062 14560 11190 14612
rect 11210 14888 11338 14940
rect 11338 14888 11462 14940
rect 11462 14888 11590 14940
rect 11210 14612 11590 14888
rect 11210 14560 11338 14612
rect 11338 14560 11462 14612
rect 11462 14560 11590 14612
rect 11610 14888 11738 14940
rect 11738 14888 11862 14940
rect 11862 14888 11990 14940
rect 11610 14612 11990 14888
rect 11610 14560 11738 14612
rect 11738 14560 11862 14612
rect 11862 14560 11990 14612
rect 12010 14888 12138 14940
rect 12138 14888 12262 14940
rect 12262 14888 12390 14940
rect 12010 14612 12390 14888
rect 12010 14560 12138 14612
rect 12138 14560 12262 14612
rect 12262 14560 12390 14612
rect 12410 14888 12538 14940
rect 12538 14888 12662 14940
rect 12662 14888 12790 14940
rect 12410 14612 12790 14888
rect 12410 14560 12538 14612
rect 12538 14560 12662 14612
rect 12662 14560 12790 14612
rect 12810 14888 12938 14940
rect 12938 14888 13062 14940
rect 13062 14888 13190 14940
rect 12810 14612 13190 14888
rect 12810 14560 12938 14612
rect 12938 14560 13062 14612
rect 13062 14560 13190 14612
rect 13210 14888 13338 14940
rect 13338 14888 13462 14940
rect 13462 14888 13590 14940
rect 13210 14612 13590 14888
rect 13210 14560 13338 14612
rect 13338 14560 13462 14612
rect 13462 14560 13590 14612
rect 13610 14888 13738 14940
rect 13738 14888 13862 14940
rect 13862 14888 13990 14940
rect 13610 14612 13990 14888
rect 13610 14560 13738 14612
rect 13738 14560 13862 14612
rect 13862 14560 13990 14612
rect 14010 14888 14138 14940
rect 14138 14888 14262 14940
rect 14262 14888 14390 14940
rect 14010 14612 14390 14888
rect 14010 14560 14138 14612
rect 14138 14560 14262 14612
rect 14262 14560 14390 14612
rect 14410 14888 14538 14940
rect 14538 14888 14662 14940
rect 14662 14888 14790 14940
rect 14410 14612 14790 14888
rect 14410 14560 14538 14612
rect 14538 14560 14662 14612
rect 14662 14560 14790 14612
rect 14810 14888 14938 14940
rect 14938 14888 15062 14940
rect 15062 14888 15190 14940
rect 14810 14612 15190 14888
rect 14810 14560 14938 14612
rect 14938 14560 15062 14612
rect 15062 14560 15190 14612
rect 15210 14888 15338 14940
rect 15338 14888 15462 14940
rect 15462 14888 15590 14940
rect 15210 14612 15590 14888
rect 15210 14560 15338 14612
rect 15338 14560 15462 14612
rect 15462 14560 15590 14612
rect 410 14488 538 14540
rect 538 14488 662 14540
rect 662 14488 790 14540
rect 410 14212 790 14488
rect 410 14160 538 14212
rect 538 14160 662 14212
rect 662 14160 790 14212
rect 810 14488 938 14540
rect 938 14488 1062 14540
rect 1062 14488 1190 14540
rect 810 14212 1190 14488
rect 810 14160 938 14212
rect 938 14160 1062 14212
rect 1062 14160 1190 14212
rect 1210 14488 1338 14540
rect 1338 14488 1462 14540
rect 1462 14488 1590 14540
rect 1210 14212 1590 14488
rect 1210 14160 1338 14212
rect 1338 14160 1462 14212
rect 1462 14160 1590 14212
rect 1610 14488 1738 14540
rect 1738 14488 1862 14540
rect 1862 14488 1990 14540
rect 1610 14212 1990 14488
rect 1610 14160 1738 14212
rect 1738 14160 1862 14212
rect 1862 14160 1990 14212
rect 2010 14488 2138 14540
rect 2138 14488 2262 14540
rect 2262 14488 2390 14540
rect 2010 14212 2390 14488
rect 2010 14160 2138 14212
rect 2138 14160 2262 14212
rect 2262 14160 2390 14212
rect 2410 14488 2538 14540
rect 2538 14488 2662 14540
rect 2662 14488 2790 14540
rect 2410 14212 2790 14488
rect 2410 14160 2538 14212
rect 2538 14160 2662 14212
rect 2662 14160 2790 14212
rect 2810 14488 2938 14540
rect 2938 14488 3062 14540
rect 3062 14488 3190 14540
rect 2810 14212 3190 14488
rect 2810 14160 2938 14212
rect 2938 14160 3062 14212
rect 3062 14160 3190 14212
rect 3210 14488 3338 14540
rect 3338 14488 3462 14540
rect 3462 14488 3590 14540
rect 3210 14212 3590 14488
rect 3210 14160 3338 14212
rect 3338 14160 3462 14212
rect 3462 14160 3590 14212
rect 3610 14488 3738 14540
rect 3738 14488 3862 14540
rect 3862 14488 3990 14540
rect 3610 14212 3990 14488
rect 3610 14160 3738 14212
rect 3738 14160 3862 14212
rect 3862 14160 3990 14212
rect 4010 14488 4138 14540
rect 4138 14488 4262 14540
rect 4262 14488 4390 14540
rect 4010 14212 4390 14488
rect 4010 14160 4138 14212
rect 4138 14160 4262 14212
rect 4262 14160 4390 14212
rect 4410 14488 4538 14540
rect 4538 14488 4662 14540
rect 4662 14488 4790 14540
rect 4410 14212 4790 14488
rect 4410 14160 4538 14212
rect 4538 14160 4662 14212
rect 4662 14160 4790 14212
rect 4810 14488 4938 14540
rect 4938 14488 5062 14540
rect 5062 14488 5190 14540
rect 4810 14212 5190 14488
rect 4810 14160 4938 14212
rect 4938 14160 5062 14212
rect 5062 14160 5190 14212
rect 5210 14488 5338 14540
rect 5338 14488 5462 14540
rect 5462 14488 5590 14540
rect 5210 14212 5590 14488
rect 5210 14160 5338 14212
rect 5338 14160 5462 14212
rect 5462 14160 5590 14212
rect 5610 14488 5738 14540
rect 5738 14488 5862 14540
rect 5862 14488 5990 14540
rect 5610 14212 5990 14488
rect 5610 14160 5738 14212
rect 5738 14160 5862 14212
rect 5862 14160 5990 14212
rect 6010 14488 6138 14540
rect 6138 14488 6262 14540
rect 6262 14488 6390 14540
rect 6010 14212 6390 14488
rect 6010 14160 6138 14212
rect 6138 14160 6262 14212
rect 6262 14160 6390 14212
rect 6410 14488 6538 14540
rect 6538 14488 6662 14540
rect 6662 14488 6790 14540
rect 6410 14212 6790 14488
rect 6410 14160 6538 14212
rect 6538 14160 6662 14212
rect 6662 14160 6790 14212
rect 6810 14488 6938 14540
rect 6938 14488 7062 14540
rect 7062 14488 7190 14540
rect 6810 14212 7190 14488
rect 6810 14160 6938 14212
rect 6938 14160 7062 14212
rect 7062 14160 7190 14212
rect 7210 14488 7338 14540
rect 7338 14488 7462 14540
rect 7462 14488 7590 14540
rect 7210 14212 7590 14488
rect 7210 14160 7338 14212
rect 7338 14160 7462 14212
rect 7462 14160 7590 14212
rect 7610 14488 7738 14540
rect 7738 14488 7862 14540
rect 7862 14488 7990 14540
rect 7610 14212 7990 14488
rect 7610 14160 7738 14212
rect 7738 14160 7862 14212
rect 7862 14160 7990 14212
rect 8010 14488 8138 14540
rect 8138 14488 8262 14540
rect 8262 14488 8390 14540
rect 8010 14212 8390 14488
rect 8010 14160 8138 14212
rect 8138 14160 8262 14212
rect 8262 14160 8390 14212
rect 8410 14488 8538 14540
rect 8538 14488 8662 14540
rect 8662 14488 8790 14540
rect 8410 14212 8790 14488
rect 8410 14160 8538 14212
rect 8538 14160 8662 14212
rect 8662 14160 8790 14212
rect 8810 14488 8938 14540
rect 8938 14488 9062 14540
rect 9062 14488 9190 14540
rect 8810 14212 9190 14488
rect 8810 14160 8938 14212
rect 8938 14160 9062 14212
rect 9062 14160 9190 14212
rect 9210 14488 9338 14540
rect 9338 14488 9462 14540
rect 9462 14488 9590 14540
rect 9210 14212 9590 14488
rect 9210 14160 9338 14212
rect 9338 14160 9462 14212
rect 9462 14160 9590 14212
rect 9610 14488 9738 14540
rect 9738 14488 9862 14540
rect 9862 14488 9990 14540
rect 9610 14212 9990 14488
rect 9610 14160 9738 14212
rect 9738 14160 9862 14212
rect 9862 14160 9990 14212
rect 10010 14488 10138 14540
rect 10138 14488 10262 14540
rect 10262 14488 10390 14540
rect 10010 14212 10390 14488
rect 10010 14160 10138 14212
rect 10138 14160 10262 14212
rect 10262 14160 10390 14212
rect 10410 14488 10538 14540
rect 10538 14488 10662 14540
rect 10662 14488 10790 14540
rect 10410 14212 10790 14488
rect 10410 14160 10538 14212
rect 10538 14160 10662 14212
rect 10662 14160 10790 14212
rect 10810 14488 10938 14540
rect 10938 14488 11062 14540
rect 11062 14488 11190 14540
rect 10810 14212 11190 14488
rect 10810 14160 10938 14212
rect 10938 14160 11062 14212
rect 11062 14160 11190 14212
rect 11210 14488 11338 14540
rect 11338 14488 11462 14540
rect 11462 14488 11590 14540
rect 11210 14212 11590 14488
rect 11210 14160 11338 14212
rect 11338 14160 11462 14212
rect 11462 14160 11590 14212
rect 11610 14488 11738 14540
rect 11738 14488 11862 14540
rect 11862 14488 11990 14540
rect 11610 14212 11990 14488
rect 11610 14160 11738 14212
rect 11738 14160 11862 14212
rect 11862 14160 11990 14212
rect 12010 14488 12138 14540
rect 12138 14488 12262 14540
rect 12262 14488 12390 14540
rect 12010 14212 12390 14488
rect 12010 14160 12138 14212
rect 12138 14160 12262 14212
rect 12262 14160 12390 14212
rect 12410 14488 12538 14540
rect 12538 14488 12662 14540
rect 12662 14488 12790 14540
rect 12410 14212 12790 14488
rect 12410 14160 12538 14212
rect 12538 14160 12662 14212
rect 12662 14160 12790 14212
rect 12810 14488 12938 14540
rect 12938 14488 13062 14540
rect 13062 14488 13190 14540
rect 12810 14212 13190 14488
rect 12810 14160 12938 14212
rect 12938 14160 13062 14212
rect 13062 14160 13190 14212
rect 13210 14488 13338 14540
rect 13338 14488 13462 14540
rect 13462 14488 13590 14540
rect 13210 14212 13590 14488
rect 13210 14160 13338 14212
rect 13338 14160 13462 14212
rect 13462 14160 13590 14212
rect 13610 14488 13738 14540
rect 13738 14488 13862 14540
rect 13862 14488 13990 14540
rect 13610 14212 13990 14488
rect 13610 14160 13738 14212
rect 13738 14160 13862 14212
rect 13862 14160 13990 14212
rect 14010 14488 14138 14540
rect 14138 14488 14262 14540
rect 14262 14488 14390 14540
rect 14010 14212 14390 14488
rect 14010 14160 14138 14212
rect 14138 14160 14262 14212
rect 14262 14160 14390 14212
rect 14410 14488 14538 14540
rect 14538 14488 14662 14540
rect 14662 14488 14790 14540
rect 14410 14212 14790 14488
rect 14410 14160 14538 14212
rect 14538 14160 14662 14212
rect 14662 14160 14790 14212
rect 14810 14488 14938 14540
rect 14938 14488 15062 14540
rect 15062 14488 15190 14540
rect 14810 14212 15190 14488
rect 14810 14160 14938 14212
rect 14938 14160 15062 14212
rect 15062 14160 15190 14212
rect 15210 14488 15338 14540
rect 15338 14488 15462 14540
rect 15462 14488 15590 14540
rect 15210 14212 15590 14488
rect 15210 14160 15338 14212
rect 15338 14160 15462 14212
rect 15462 14160 15590 14212
rect 410 14088 538 14140
rect 538 14088 662 14140
rect 662 14088 790 14140
rect 410 13812 790 14088
rect 410 13760 538 13812
rect 538 13760 662 13812
rect 662 13760 790 13812
rect 810 14088 938 14140
rect 938 14088 1062 14140
rect 1062 14088 1190 14140
rect 810 13812 1190 14088
rect 810 13760 938 13812
rect 938 13760 1062 13812
rect 1062 13760 1190 13812
rect 1210 14088 1338 14140
rect 1338 14088 1462 14140
rect 1462 14088 1590 14140
rect 1210 13812 1590 14088
rect 1210 13760 1338 13812
rect 1338 13760 1462 13812
rect 1462 13760 1590 13812
rect 1610 14088 1738 14140
rect 1738 14088 1862 14140
rect 1862 14088 1990 14140
rect 1610 13812 1990 14088
rect 1610 13760 1738 13812
rect 1738 13760 1862 13812
rect 1862 13760 1990 13812
rect 2010 14088 2138 14140
rect 2138 14088 2262 14140
rect 2262 14088 2390 14140
rect 2010 13812 2390 14088
rect 2010 13760 2138 13812
rect 2138 13760 2262 13812
rect 2262 13760 2390 13812
rect 2410 14088 2538 14140
rect 2538 14088 2662 14140
rect 2662 14088 2790 14140
rect 2410 13812 2790 14088
rect 2410 13760 2538 13812
rect 2538 13760 2662 13812
rect 2662 13760 2790 13812
rect 2810 14088 2938 14140
rect 2938 14088 3062 14140
rect 3062 14088 3190 14140
rect 2810 13812 3190 14088
rect 2810 13760 2938 13812
rect 2938 13760 3062 13812
rect 3062 13760 3190 13812
rect 3210 14088 3338 14140
rect 3338 14088 3462 14140
rect 3462 14088 3590 14140
rect 3210 13812 3590 14088
rect 3210 13760 3338 13812
rect 3338 13760 3462 13812
rect 3462 13760 3590 13812
rect 3610 14088 3738 14140
rect 3738 14088 3862 14140
rect 3862 14088 3990 14140
rect 3610 13812 3990 14088
rect 3610 13760 3738 13812
rect 3738 13760 3862 13812
rect 3862 13760 3990 13812
rect 4010 14088 4138 14140
rect 4138 14088 4262 14140
rect 4262 14088 4390 14140
rect 4010 13812 4390 14088
rect 4010 13760 4138 13812
rect 4138 13760 4262 13812
rect 4262 13760 4390 13812
rect 4410 14088 4538 14140
rect 4538 14088 4662 14140
rect 4662 14088 4790 14140
rect 4410 13812 4790 14088
rect 4410 13760 4538 13812
rect 4538 13760 4662 13812
rect 4662 13760 4790 13812
rect 4810 14088 4938 14140
rect 4938 14088 5062 14140
rect 5062 14088 5190 14140
rect 4810 13812 5190 14088
rect 4810 13760 4938 13812
rect 4938 13760 5062 13812
rect 5062 13760 5190 13812
rect 5210 14088 5338 14140
rect 5338 14088 5462 14140
rect 5462 14088 5590 14140
rect 5210 13812 5590 14088
rect 5210 13760 5338 13812
rect 5338 13760 5462 13812
rect 5462 13760 5590 13812
rect 5610 14088 5738 14140
rect 5738 14088 5862 14140
rect 5862 14088 5990 14140
rect 5610 13812 5990 14088
rect 5610 13760 5738 13812
rect 5738 13760 5862 13812
rect 5862 13760 5990 13812
rect 6010 14088 6138 14140
rect 6138 14088 6262 14140
rect 6262 14088 6390 14140
rect 6010 13812 6390 14088
rect 6010 13760 6138 13812
rect 6138 13760 6262 13812
rect 6262 13760 6390 13812
rect 6410 14088 6538 14140
rect 6538 14088 6662 14140
rect 6662 14088 6790 14140
rect 6410 13812 6790 14088
rect 6410 13760 6538 13812
rect 6538 13760 6662 13812
rect 6662 13760 6790 13812
rect 6810 14088 6938 14140
rect 6938 14088 7062 14140
rect 7062 14088 7190 14140
rect 6810 13812 7190 14088
rect 6810 13760 6938 13812
rect 6938 13760 7062 13812
rect 7062 13760 7190 13812
rect 7210 14088 7338 14140
rect 7338 14088 7462 14140
rect 7462 14088 7590 14140
rect 7210 13812 7590 14088
rect 7210 13760 7338 13812
rect 7338 13760 7462 13812
rect 7462 13760 7590 13812
rect 7610 14088 7738 14140
rect 7738 14088 7862 14140
rect 7862 14088 7990 14140
rect 7610 13812 7990 14088
rect 7610 13760 7738 13812
rect 7738 13760 7862 13812
rect 7862 13760 7990 13812
rect 8010 14088 8138 14140
rect 8138 14088 8262 14140
rect 8262 14088 8390 14140
rect 8010 13812 8390 14088
rect 8010 13760 8138 13812
rect 8138 13760 8262 13812
rect 8262 13760 8390 13812
rect 8410 14088 8538 14140
rect 8538 14088 8662 14140
rect 8662 14088 8790 14140
rect 8410 13812 8790 14088
rect 8410 13760 8538 13812
rect 8538 13760 8662 13812
rect 8662 13760 8790 13812
rect 8810 14088 8938 14140
rect 8938 14088 9062 14140
rect 9062 14088 9190 14140
rect 8810 13812 9190 14088
rect 8810 13760 8938 13812
rect 8938 13760 9062 13812
rect 9062 13760 9190 13812
rect 9210 14088 9338 14140
rect 9338 14088 9462 14140
rect 9462 14088 9590 14140
rect 9210 13812 9590 14088
rect 9210 13760 9338 13812
rect 9338 13760 9462 13812
rect 9462 13760 9590 13812
rect 9610 14088 9738 14140
rect 9738 14088 9862 14140
rect 9862 14088 9990 14140
rect 9610 13812 9990 14088
rect 9610 13760 9738 13812
rect 9738 13760 9862 13812
rect 9862 13760 9990 13812
rect 10010 14088 10138 14140
rect 10138 14088 10262 14140
rect 10262 14088 10390 14140
rect 10010 13812 10390 14088
rect 10010 13760 10138 13812
rect 10138 13760 10262 13812
rect 10262 13760 10390 13812
rect 10410 14088 10538 14140
rect 10538 14088 10662 14140
rect 10662 14088 10790 14140
rect 10410 13812 10790 14088
rect 10410 13760 10538 13812
rect 10538 13760 10662 13812
rect 10662 13760 10790 13812
rect 10810 14088 10938 14140
rect 10938 14088 11062 14140
rect 11062 14088 11190 14140
rect 10810 13812 11190 14088
rect 10810 13760 10938 13812
rect 10938 13760 11062 13812
rect 11062 13760 11190 13812
rect 11210 14088 11338 14140
rect 11338 14088 11462 14140
rect 11462 14088 11590 14140
rect 11210 13812 11590 14088
rect 11210 13760 11338 13812
rect 11338 13760 11462 13812
rect 11462 13760 11590 13812
rect 11610 14088 11738 14140
rect 11738 14088 11862 14140
rect 11862 14088 11990 14140
rect 11610 13812 11990 14088
rect 11610 13760 11738 13812
rect 11738 13760 11862 13812
rect 11862 13760 11990 13812
rect 12010 14088 12138 14140
rect 12138 14088 12262 14140
rect 12262 14088 12390 14140
rect 12010 13812 12390 14088
rect 12010 13760 12138 13812
rect 12138 13760 12262 13812
rect 12262 13760 12390 13812
rect 12410 14088 12538 14140
rect 12538 14088 12662 14140
rect 12662 14088 12790 14140
rect 12410 13812 12790 14088
rect 12410 13760 12538 13812
rect 12538 13760 12662 13812
rect 12662 13760 12790 13812
rect 12810 14088 12938 14140
rect 12938 14088 13062 14140
rect 13062 14088 13190 14140
rect 12810 13812 13190 14088
rect 12810 13760 12938 13812
rect 12938 13760 13062 13812
rect 13062 13760 13190 13812
rect 13210 14088 13338 14140
rect 13338 14088 13462 14140
rect 13462 14088 13590 14140
rect 13210 13812 13590 14088
rect 13210 13760 13338 13812
rect 13338 13760 13462 13812
rect 13462 13760 13590 13812
rect 13610 14088 13738 14140
rect 13738 14088 13862 14140
rect 13862 14088 13990 14140
rect 13610 13812 13990 14088
rect 13610 13760 13738 13812
rect 13738 13760 13862 13812
rect 13862 13760 13990 13812
rect 14010 14088 14138 14140
rect 14138 14088 14262 14140
rect 14262 14088 14390 14140
rect 14010 13812 14390 14088
rect 14010 13760 14138 13812
rect 14138 13760 14262 13812
rect 14262 13760 14390 13812
rect 14410 14088 14538 14140
rect 14538 14088 14662 14140
rect 14662 14088 14790 14140
rect 14410 13812 14790 14088
rect 14410 13760 14538 13812
rect 14538 13760 14662 13812
rect 14662 13760 14790 13812
rect 14810 14088 14938 14140
rect 14938 14088 15062 14140
rect 15062 14088 15190 14140
rect 14810 13812 15190 14088
rect 14810 13760 14938 13812
rect 14938 13760 15062 13812
rect 15062 13760 15190 13812
rect 15210 14088 15338 14140
rect 15338 14088 15462 14140
rect 15462 14088 15590 14140
rect 15210 13812 15590 14088
rect 15210 13760 15338 13812
rect 15338 13760 15462 13812
rect 15462 13760 15590 13812
rect 0 11260 380 11640
rect 400 11512 780 11640
rect 15220 11512 15600 11640
rect 400 11388 538 11512
rect 538 11388 662 11512
rect 662 11388 780 11512
rect 15220 11388 15338 11512
rect 15338 11388 15462 11512
rect 15462 11388 15600 11512
rect 400 11260 780 11388
rect 15220 11260 15600 11388
rect 15620 11260 16000 11640
rect 0 10860 380 11240
rect 400 11112 780 11240
rect 15220 11112 15600 11240
rect 400 10988 538 11112
rect 538 10988 662 11112
rect 662 10988 780 11112
rect 15220 10988 15338 11112
rect 15338 10988 15462 11112
rect 15462 10988 15600 11112
rect 400 10860 780 10988
rect 15220 10860 15600 10988
rect 15620 10860 16000 11240
rect 0 10460 380 10840
rect 400 10712 780 10840
rect 15220 10712 15600 10840
rect 400 10588 538 10712
rect 538 10588 662 10712
rect 662 10588 780 10712
rect 15220 10588 15338 10712
rect 15338 10588 15462 10712
rect 15462 10588 15600 10712
rect 400 10460 780 10588
rect 15220 10460 15600 10588
rect 15620 10460 16000 10840
rect 0 10060 380 10440
rect 400 10312 780 10440
rect 15220 10312 15600 10440
rect 400 10188 538 10312
rect 538 10188 662 10312
rect 662 10188 780 10312
rect 15220 10188 15338 10312
rect 15338 10188 15462 10312
rect 15462 10188 15600 10312
rect 400 10060 780 10188
rect 15220 10060 15600 10188
rect 15620 10060 16000 10440
rect 0 9660 380 10040
rect 400 9912 780 10040
rect 15220 9912 15600 10040
rect 400 9788 538 9912
rect 538 9788 662 9912
rect 662 9788 780 9912
rect 15220 9788 15338 9912
rect 15338 9788 15462 9912
rect 15462 9788 15600 9912
rect 400 9660 780 9788
rect 15220 9660 15600 9788
rect 15620 9660 16000 10040
rect 0 9260 380 9640
rect 400 9512 780 9640
rect 15220 9512 15600 9640
rect 400 9388 538 9512
rect 538 9388 662 9512
rect 662 9388 780 9512
rect 15220 9388 15338 9512
rect 15338 9388 15462 9512
rect 15462 9388 15600 9512
rect 400 9260 780 9388
rect 15220 9260 15600 9388
rect 15620 9260 16000 9640
rect 0 8860 380 9240
rect 400 9112 780 9240
rect 15220 9112 15600 9240
rect 400 8988 538 9112
rect 538 8988 662 9112
rect 662 8988 780 9112
rect 15220 8988 15338 9112
rect 15338 8988 15462 9112
rect 15462 8988 15600 9112
rect 400 8860 780 8988
rect 15220 8860 15600 8988
rect 15620 8860 16000 9240
rect 0 8460 380 8840
rect 400 8712 780 8840
rect 15220 8712 15600 8840
rect 400 8588 538 8712
rect 538 8588 662 8712
rect 662 8588 780 8712
rect 15220 8588 15338 8712
rect 15338 8588 15462 8712
rect 15462 8588 15600 8712
rect 400 8460 780 8588
rect 15220 8460 15600 8588
rect 15620 8460 16000 8840
rect 0 8060 380 8440
rect 400 8312 780 8440
rect 15220 8312 15600 8440
rect 400 8188 538 8312
rect 538 8188 662 8312
rect 662 8188 780 8312
rect 15220 8188 15338 8312
rect 15338 8188 15462 8312
rect 15462 8188 15600 8312
rect 400 8060 780 8188
rect 15220 8060 15600 8188
rect 15620 8060 16000 8440
rect 0 7660 380 8040
rect 400 7912 780 8040
rect 15220 7912 15600 8040
rect 400 7788 538 7912
rect 538 7788 662 7912
rect 662 7788 780 7912
rect 15220 7788 15338 7912
rect 15338 7788 15462 7912
rect 15462 7788 15600 7912
rect 400 7660 780 7788
rect 15220 7660 15600 7788
rect 15620 7660 16000 8040
rect 0 7260 380 7640
rect 400 7512 780 7640
rect 15220 7512 15600 7640
rect 400 7388 538 7512
rect 538 7388 662 7512
rect 662 7388 780 7512
rect 15220 7388 15338 7512
rect 15338 7388 15462 7512
rect 15462 7388 15600 7512
rect 400 7260 780 7388
rect 15220 7260 15600 7388
rect 15620 7260 16000 7640
rect 0 5760 380 6140
rect 400 6012 780 6140
rect 15220 6012 15600 6140
rect 400 5888 538 6012
rect 538 5888 662 6012
rect 662 5888 780 6012
rect 15220 5888 15338 6012
rect 15338 5888 15462 6012
rect 15462 5888 15600 6012
rect 400 5760 780 5888
rect 15220 5760 15600 5888
rect 15620 5760 16000 6140
rect 0 5360 380 5740
rect 400 5612 780 5740
rect 15220 5612 15600 5740
rect 400 5488 538 5612
rect 538 5488 662 5612
rect 662 5488 780 5612
rect 15220 5488 15338 5612
rect 15338 5488 15462 5612
rect 15462 5488 15600 5612
rect 400 5360 780 5488
rect 15220 5360 15600 5488
rect 15620 5360 16000 5740
rect 0 4960 380 5340
rect 400 5212 780 5340
rect 15220 5212 15600 5340
rect 400 5088 538 5212
rect 538 5088 662 5212
rect 662 5088 780 5212
rect 15220 5088 15338 5212
rect 15338 5088 15462 5212
rect 15462 5088 15600 5212
rect 400 4960 780 5088
rect 15220 4960 15600 5088
rect 15620 4960 16000 5340
rect 0 4560 380 4940
rect 400 4812 780 4940
rect 15220 4812 15600 4940
rect 400 4688 538 4812
rect 538 4688 662 4812
rect 662 4688 780 4812
rect 15220 4688 15338 4812
rect 15338 4688 15462 4812
rect 15462 4688 15600 4812
rect 400 4560 780 4688
rect 15220 4560 15600 4688
rect 15620 4560 16000 4940
rect 0 4160 380 4540
rect 400 4412 780 4540
rect 15220 4412 15600 4540
rect 400 4288 538 4412
rect 538 4288 662 4412
rect 662 4288 780 4412
rect 15220 4288 15338 4412
rect 15338 4288 15462 4412
rect 15462 4288 15600 4412
rect 400 4160 780 4288
rect 15220 4160 15600 4288
rect 15620 4160 16000 4540
rect 0 3760 380 4140
rect 400 4012 780 4140
rect 15220 4012 15600 4140
rect 400 3888 538 4012
rect 538 3888 662 4012
rect 662 3888 780 4012
rect 15220 3888 15338 4012
rect 15338 3888 15462 4012
rect 15462 3888 15600 4012
rect 400 3760 780 3888
rect 15220 3760 15600 3888
rect 15620 3760 16000 4140
rect 0 3360 380 3740
rect 400 3612 780 3740
rect 15220 3612 15600 3740
rect 400 3488 538 3612
rect 538 3488 662 3612
rect 662 3488 780 3612
rect 15220 3488 15338 3612
rect 15338 3488 15462 3612
rect 15462 3488 15600 3612
rect 400 3360 780 3488
rect 15220 3360 15600 3488
rect 15620 3360 16000 3740
rect 0 2960 380 3340
rect 400 3212 780 3340
rect 15220 3212 15600 3340
rect 400 3088 538 3212
rect 538 3088 662 3212
rect 662 3088 780 3212
rect 15220 3088 15338 3212
rect 15338 3088 15462 3212
rect 15462 3088 15600 3212
rect 400 2960 780 3088
rect 15220 2960 15600 3088
rect 15620 2960 16000 3340
rect 0 2560 380 2940
rect 400 2812 780 2940
rect 15220 2812 15600 2940
rect 400 2688 538 2812
rect 538 2688 662 2812
rect 662 2688 780 2812
rect 15220 2688 15338 2812
rect 15338 2688 15462 2812
rect 15462 2688 15600 2812
rect 400 2560 780 2688
rect 15220 2560 15600 2688
rect 15620 2560 16000 2940
rect 0 2160 380 2540
rect 400 2412 780 2540
rect 15220 2412 15600 2540
rect 400 2288 538 2412
rect 538 2288 662 2412
rect 662 2288 780 2412
rect 15220 2288 15338 2412
rect 15338 2288 15462 2412
rect 15462 2288 15600 2412
rect 400 2160 780 2288
rect 15220 2160 15600 2288
rect 15620 2160 16000 2540
rect 0 1760 380 2140
rect 400 2012 780 2140
rect 15220 2012 15600 2140
rect 400 1888 538 2012
rect 538 1888 662 2012
rect 662 1888 780 2012
rect 15220 1888 15338 2012
rect 15338 1888 15462 2012
rect 15462 1888 15600 2012
rect 400 1760 780 1888
rect 15220 1760 15600 1888
rect 15620 1760 16000 2140
rect 1010 362 1390 490
rect 1010 238 1138 362
rect 1138 238 1262 362
rect 1262 238 1390 362
rect 1010 110 1390 238
rect 1410 362 1790 490
rect 1410 238 1538 362
rect 1538 238 1662 362
rect 1662 238 1790 362
rect 1410 110 1790 238
rect 1810 362 2190 490
rect 1810 238 1938 362
rect 1938 238 2062 362
rect 2062 238 2190 362
rect 1810 110 2190 238
rect 2210 362 2590 490
rect 2210 238 2338 362
rect 2338 238 2462 362
rect 2462 238 2590 362
rect 2210 110 2590 238
rect 2610 362 2990 490
rect 2610 238 2738 362
rect 2738 238 2862 362
rect 2862 238 2990 362
rect 2610 110 2990 238
rect 3010 362 3390 490
rect 3010 238 3138 362
rect 3138 238 3262 362
rect 3262 238 3390 362
rect 3010 110 3390 238
rect 3410 362 3790 490
rect 3410 238 3538 362
rect 3538 238 3662 362
rect 3662 238 3790 362
rect 3410 110 3790 238
rect 3810 362 4190 490
rect 3810 238 3938 362
rect 3938 238 4062 362
rect 4062 238 4190 362
rect 3810 110 4190 238
rect 4210 362 4590 490
rect 4210 238 4338 362
rect 4338 238 4462 362
rect 4462 238 4590 362
rect 4210 110 4590 238
rect 4610 362 4990 490
rect 4610 238 4738 362
rect 4738 238 4862 362
rect 4862 238 4990 362
rect 4610 110 4990 238
rect 5010 362 5390 490
rect 5010 238 5138 362
rect 5138 238 5262 362
rect 5262 238 5390 362
rect 5010 110 5390 238
rect 5410 362 5790 490
rect 5410 238 5538 362
rect 5538 238 5662 362
rect 5662 238 5790 362
rect 5410 110 5790 238
rect 5810 362 6190 490
rect 5810 238 5938 362
rect 5938 238 6062 362
rect 6062 238 6190 362
rect 5810 110 6190 238
rect 6210 362 6590 490
rect 6210 238 6338 362
rect 6338 238 6462 362
rect 6462 238 6590 362
rect 6210 110 6590 238
rect 6610 362 6990 490
rect 6610 238 6738 362
rect 6738 238 6862 362
rect 6862 238 6990 362
rect 6610 110 6990 238
rect 7010 362 7390 490
rect 7010 238 7138 362
rect 7138 238 7262 362
rect 7262 238 7390 362
rect 7010 110 7390 238
rect 7410 362 7790 490
rect 7410 238 7538 362
rect 7538 238 7662 362
rect 7662 238 7790 362
rect 7410 110 7790 238
rect 7810 362 8190 490
rect 7810 238 7938 362
rect 7938 238 8062 362
rect 8062 238 8190 362
rect 7810 110 8190 238
rect 8210 362 8590 490
rect 8210 238 8338 362
rect 8338 238 8462 362
rect 8462 238 8590 362
rect 8210 110 8590 238
rect 8610 362 8990 490
rect 8610 238 8738 362
rect 8738 238 8862 362
rect 8862 238 8990 362
rect 8610 110 8990 238
rect 9010 362 9390 490
rect 9010 238 9138 362
rect 9138 238 9262 362
rect 9262 238 9390 362
rect 9010 110 9390 238
rect 9410 362 9790 490
rect 9410 238 9538 362
rect 9538 238 9662 362
rect 9662 238 9790 362
rect 9410 110 9790 238
rect 9810 362 10190 490
rect 9810 238 9938 362
rect 9938 238 10062 362
rect 10062 238 10190 362
rect 9810 110 10190 238
rect 10210 362 10590 490
rect 10210 238 10338 362
rect 10338 238 10462 362
rect 10462 238 10590 362
rect 10210 110 10590 238
rect 10610 362 10990 490
rect 10610 238 10738 362
rect 10738 238 10862 362
rect 10862 238 10990 362
rect 10610 110 10990 238
rect 11010 362 11390 490
rect 11010 238 11138 362
rect 11138 238 11262 362
rect 11262 238 11390 362
rect 11010 110 11390 238
rect 11410 362 11790 490
rect 11410 238 11538 362
rect 11538 238 11662 362
rect 11662 238 11790 362
rect 11410 110 11790 238
rect 11810 362 12190 490
rect 11810 238 11938 362
rect 11938 238 12062 362
rect 12062 238 12190 362
rect 11810 110 12190 238
rect 12210 362 12590 490
rect 12210 238 12338 362
rect 12338 238 12462 362
rect 12462 238 12590 362
rect 12210 110 12590 238
rect 12610 362 12990 490
rect 12610 238 12738 362
rect 12738 238 12862 362
rect 12862 238 12990 362
rect 12610 110 12990 238
rect 13010 362 13390 490
rect 13010 238 13138 362
rect 13138 238 13262 362
rect 13262 238 13390 362
rect 13010 110 13390 238
rect 13410 362 13790 490
rect 13410 238 13538 362
rect 13538 238 13662 362
rect 13662 238 13790 362
rect 13410 110 13790 238
rect 13810 362 14190 490
rect 13810 238 13938 362
rect 13938 238 14062 362
rect 14062 238 14190 362
rect 13810 110 14190 238
rect 14210 362 14590 490
rect 14210 238 14338 362
rect 14338 238 14462 362
rect 14462 238 14590 362
rect 14210 110 14590 238
rect 14610 362 14990 490
rect 14610 238 14738 362
rect 14738 238 14862 362
rect 14862 238 14990 362
rect 14610 110 14990 238
<< metal7 >>
rect 0 26190 16000 26500
rect 0 25810 410 26190
rect 790 25810 810 26190
rect 1190 25810 1210 26190
rect 1590 25810 1610 26190
rect 1990 25810 2010 26190
rect 2390 25810 2410 26190
rect 2790 25810 2810 26190
rect 3190 25810 3210 26190
rect 3590 25810 3610 26190
rect 3990 25810 4010 26190
rect 4390 25810 4410 26190
rect 4790 25810 4810 26190
rect 5190 25810 5210 26190
rect 5590 25810 5610 26190
rect 5990 25810 6010 26190
rect 6390 25810 6410 26190
rect 6790 25810 6810 26190
rect 7190 25810 7210 26190
rect 7590 25810 7610 26190
rect 7990 25810 8010 26190
rect 8390 25810 8410 26190
rect 8790 25810 8810 26190
rect 9190 25810 9210 26190
rect 9590 25810 9610 26190
rect 9990 25810 10010 26190
rect 10390 25810 10410 26190
rect 10790 25810 10810 26190
rect 11190 25810 11210 26190
rect 11590 25810 11610 26190
rect 11990 25810 12010 26190
rect 12390 25810 12410 26190
rect 12790 25810 12810 26190
rect 13190 25810 13210 26190
rect 13590 25810 13610 26190
rect 13990 25810 14010 26190
rect 14390 25810 14410 26190
rect 14790 25810 14810 26190
rect 15190 25810 15210 26190
rect 15590 25810 16000 26190
rect 0 25500 16000 25810
rect 0 23240 16000 23500
rect 0 22860 410 23240
rect 790 22860 810 23240
rect 1190 22860 1210 23240
rect 1590 22860 1610 23240
rect 1990 22860 2010 23240
rect 2390 22860 2410 23240
rect 2790 22860 2810 23240
rect 3190 22860 3210 23240
rect 3590 22860 3610 23240
rect 3990 22860 4010 23240
rect 4390 22860 4410 23240
rect 4790 22860 4810 23240
rect 5190 22860 5210 23240
rect 5590 22860 5610 23240
rect 5990 22860 6010 23240
rect 6390 22860 6410 23240
rect 6790 22860 6810 23240
rect 7190 22860 7210 23240
rect 7590 22860 7610 23240
rect 7990 22860 8010 23240
rect 8390 22860 8410 23240
rect 8790 22860 8810 23240
rect 9190 22860 9210 23240
rect 9590 22860 9610 23240
rect 9990 22860 10010 23240
rect 10390 22860 10410 23240
rect 10790 22860 10810 23240
rect 11190 22860 11210 23240
rect 11590 22860 11610 23240
rect 11990 22860 12010 23240
rect 12390 22860 12410 23240
rect 12790 22860 12810 23240
rect 13190 22860 13210 23240
rect 13590 22860 13610 23240
rect 13990 22860 14010 23240
rect 14390 22860 14410 23240
rect 14790 22860 14810 23240
rect 15190 22860 15210 23240
rect 15590 22860 16000 23240
rect 0 22840 16000 22860
rect 0 22460 410 22840
rect 790 22460 810 22840
rect 1190 22460 1210 22840
rect 1590 22460 1610 22840
rect 1990 22460 2010 22840
rect 2390 22460 2410 22840
rect 2790 22460 2810 22840
rect 3190 22460 3210 22840
rect 3590 22460 3610 22840
rect 3990 22460 4010 22840
rect 4390 22460 4410 22840
rect 4790 22460 4810 22840
rect 5190 22460 5210 22840
rect 5590 22460 5610 22840
rect 5990 22460 6010 22840
rect 6390 22460 6410 22840
rect 6790 22460 6810 22840
rect 7190 22460 7210 22840
rect 7590 22460 7610 22840
rect 7990 22460 8010 22840
rect 8390 22460 8410 22840
rect 8790 22460 8810 22840
rect 9190 22460 9210 22840
rect 9590 22460 9610 22840
rect 9990 22460 10010 22840
rect 10390 22460 10410 22840
rect 10790 22460 10810 22840
rect 11190 22460 11210 22840
rect 11590 22460 11610 22840
rect 11990 22460 12010 22840
rect 12390 22460 12410 22840
rect 12790 22460 12810 22840
rect 13190 22460 13210 22840
rect 13590 22460 13610 22840
rect 13990 22460 14010 22840
rect 14390 22460 14410 22840
rect 14790 22460 14810 22840
rect 15190 22460 15210 22840
rect 15590 22460 16000 22840
rect 0 22440 16000 22460
rect 0 22060 410 22440
rect 790 22060 810 22440
rect 1190 22060 1210 22440
rect 1590 22060 1610 22440
rect 1990 22060 2010 22440
rect 2390 22060 2410 22440
rect 2790 22060 2810 22440
rect 3190 22060 3210 22440
rect 3590 22060 3610 22440
rect 3990 22060 4010 22440
rect 4390 22060 4410 22440
rect 4790 22060 4810 22440
rect 5190 22060 5210 22440
rect 5590 22060 5610 22440
rect 5990 22060 6010 22440
rect 6390 22060 6410 22440
rect 6790 22060 6810 22440
rect 7190 22060 7210 22440
rect 7590 22060 7610 22440
rect 7990 22060 8010 22440
rect 8390 22060 8410 22440
rect 8790 22060 8810 22440
rect 9190 22060 9210 22440
rect 9590 22060 9610 22440
rect 9990 22060 10010 22440
rect 10390 22060 10410 22440
rect 10790 22060 10810 22440
rect 11190 22060 11210 22440
rect 11590 22060 11610 22440
rect 11990 22060 12010 22440
rect 12390 22060 12410 22440
rect 12790 22060 12810 22440
rect 13190 22060 13210 22440
rect 13590 22060 13610 22440
rect 13990 22060 14010 22440
rect 14390 22060 14410 22440
rect 14790 22060 14810 22440
rect 15190 22060 15210 22440
rect 15590 22060 16000 22440
rect 0 22040 16000 22060
rect 0 21660 410 22040
rect 790 21660 810 22040
rect 1190 21660 1210 22040
rect 1590 21660 1610 22040
rect 1990 21660 2010 22040
rect 2390 21660 2410 22040
rect 2790 21660 2810 22040
rect 3190 21660 3210 22040
rect 3590 21660 3610 22040
rect 3990 21660 4010 22040
rect 4390 21660 4410 22040
rect 4790 21660 4810 22040
rect 5190 21660 5210 22040
rect 5590 21660 5610 22040
rect 5990 21660 6010 22040
rect 6390 21660 6410 22040
rect 6790 21660 6810 22040
rect 7190 21660 7210 22040
rect 7590 21660 7610 22040
rect 7990 21660 8010 22040
rect 8390 21660 8410 22040
rect 8790 21660 8810 22040
rect 9190 21660 9210 22040
rect 9590 21660 9610 22040
rect 9990 21660 10010 22040
rect 10390 21660 10410 22040
rect 10790 21660 10810 22040
rect 11190 21660 11210 22040
rect 11590 21660 11610 22040
rect 11990 21660 12010 22040
rect 12390 21660 12410 22040
rect 12790 21660 12810 22040
rect 13190 21660 13210 22040
rect 13590 21660 13610 22040
rect 13990 21660 14010 22040
rect 14390 21660 14410 22040
rect 14790 21660 14810 22040
rect 15190 21660 15210 22040
rect 15590 21660 16000 22040
rect 0 21640 16000 21660
rect 0 21260 410 21640
rect 790 21260 810 21640
rect 1190 21260 1210 21640
rect 1590 21260 1610 21640
rect 1990 21260 2010 21640
rect 2390 21260 2410 21640
rect 2790 21260 2810 21640
rect 3190 21260 3210 21640
rect 3590 21260 3610 21640
rect 3990 21260 4010 21640
rect 4390 21260 4410 21640
rect 4790 21260 4810 21640
rect 5190 21260 5210 21640
rect 5590 21260 5610 21640
rect 5990 21260 6010 21640
rect 6390 21260 6410 21640
rect 6790 21260 6810 21640
rect 7190 21260 7210 21640
rect 7590 21260 7610 21640
rect 7990 21260 8010 21640
rect 8390 21260 8410 21640
rect 8790 21260 8810 21640
rect 9190 21260 9210 21640
rect 9590 21260 9610 21640
rect 9990 21260 10010 21640
rect 10390 21260 10410 21640
rect 10790 21260 10810 21640
rect 11190 21260 11210 21640
rect 11590 21260 11610 21640
rect 11990 21260 12010 21640
rect 12390 21260 12410 21640
rect 12790 21260 12810 21640
rect 13190 21260 13210 21640
rect 13590 21260 13610 21640
rect 13990 21260 14010 21640
rect 14390 21260 14410 21640
rect 14790 21260 14810 21640
rect 15190 21260 15210 21640
rect 15590 21260 16000 21640
rect 0 21240 16000 21260
rect 0 20860 410 21240
rect 790 20860 810 21240
rect 1190 20860 1210 21240
rect 1590 20860 1610 21240
rect 1990 20860 2010 21240
rect 2390 20860 2410 21240
rect 2790 20860 2810 21240
rect 3190 20860 3210 21240
rect 3590 20860 3610 21240
rect 3990 20860 4010 21240
rect 4390 20860 4410 21240
rect 4790 20860 4810 21240
rect 5190 20860 5210 21240
rect 5590 20860 5610 21240
rect 5990 20860 6010 21240
rect 6390 20860 6410 21240
rect 6790 20860 6810 21240
rect 7190 20860 7210 21240
rect 7590 20860 7610 21240
rect 7990 20860 8010 21240
rect 8390 20860 8410 21240
rect 8790 20860 8810 21240
rect 9190 20860 9210 21240
rect 9590 20860 9610 21240
rect 9990 20860 10010 21240
rect 10390 20860 10410 21240
rect 10790 20860 10810 21240
rect 11190 20860 11210 21240
rect 11590 20860 11610 21240
rect 11990 20860 12010 21240
rect 12390 20860 12410 21240
rect 12790 20860 12810 21240
rect 13190 20860 13210 21240
rect 13590 20860 13610 21240
rect 13990 20860 14010 21240
rect 14390 20860 14410 21240
rect 14790 20860 14810 21240
rect 15190 20860 15210 21240
rect 15590 20860 16000 21240
rect 0 20840 16000 20860
rect 0 20460 410 20840
rect 790 20460 810 20840
rect 1190 20460 1210 20840
rect 1590 20460 1610 20840
rect 1990 20460 2010 20840
rect 2390 20460 2410 20840
rect 2790 20460 2810 20840
rect 3190 20460 3210 20840
rect 3590 20460 3610 20840
rect 3990 20460 4010 20840
rect 4390 20460 4410 20840
rect 4790 20460 4810 20840
rect 5190 20460 5210 20840
rect 5590 20460 5610 20840
rect 5990 20460 6010 20840
rect 6390 20460 6410 20840
rect 6790 20460 6810 20840
rect 7190 20460 7210 20840
rect 7590 20460 7610 20840
rect 7990 20460 8010 20840
rect 8390 20460 8410 20840
rect 8790 20460 8810 20840
rect 9190 20460 9210 20840
rect 9590 20460 9610 20840
rect 9990 20460 10010 20840
rect 10390 20460 10410 20840
rect 10790 20460 10810 20840
rect 11190 20460 11210 20840
rect 11590 20460 11610 20840
rect 11990 20460 12010 20840
rect 12390 20460 12410 20840
rect 12790 20460 12810 20840
rect 13190 20460 13210 20840
rect 13590 20460 13610 20840
rect 13990 20460 14010 20840
rect 14390 20460 14410 20840
rect 14790 20460 14810 20840
rect 15190 20460 15210 20840
rect 15590 20460 16000 20840
rect 0 20440 16000 20460
rect 0 20060 410 20440
rect 790 20060 810 20440
rect 1190 20060 1210 20440
rect 1590 20060 1610 20440
rect 1990 20060 2010 20440
rect 2390 20060 2410 20440
rect 2790 20060 2810 20440
rect 3190 20060 3210 20440
rect 3590 20060 3610 20440
rect 3990 20060 4010 20440
rect 4390 20060 4410 20440
rect 4790 20060 4810 20440
rect 5190 20060 5210 20440
rect 5590 20060 5610 20440
rect 5990 20060 6010 20440
rect 6390 20060 6410 20440
rect 6790 20060 6810 20440
rect 7190 20060 7210 20440
rect 7590 20060 7610 20440
rect 7990 20060 8010 20440
rect 8390 20060 8410 20440
rect 8790 20060 8810 20440
rect 9190 20060 9210 20440
rect 9590 20060 9610 20440
rect 9990 20060 10010 20440
rect 10390 20060 10410 20440
rect 10790 20060 10810 20440
rect 11190 20060 11210 20440
rect 11590 20060 11610 20440
rect 11990 20060 12010 20440
rect 12390 20060 12410 20440
rect 12790 20060 12810 20440
rect 13190 20060 13210 20440
rect 13590 20060 13610 20440
rect 13990 20060 14010 20440
rect 14390 20060 14410 20440
rect 14790 20060 14810 20440
rect 15190 20060 15210 20440
rect 15590 20060 16000 20440
rect 0 20040 16000 20060
rect 0 19660 410 20040
rect 790 19660 810 20040
rect 1190 19660 1210 20040
rect 1590 19660 1610 20040
rect 1990 19660 2010 20040
rect 2390 19660 2410 20040
rect 2790 19660 2810 20040
rect 3190 19660 3210 20040
rect 3590 19660 3610 20040
rect 3990 19660 4010 20040
rect 4390 19660 4410 20040
rect 4790 19660 4810 20040
rect 5190 19660 5210 20040
rect 5590 19660 5610 20040
rect 5990 19660 6010 20040
rect 6390 19660 6410 20040
rect 6790 19660 6810 20040
rect 7190 19660 7210 20040
rect 7590 19660 7610 20040
rect 7990 19660 8010 20040
rect 8390 19660 8410 20040
rect 8790 19660 8810 20040
rect 9190 19660 9210 20040
rect 9590 19660 9610 20040
rect 9990 19660 10010 20040
rect 10390 19660 10410 20040
rect 10790 19660 10810 20040
rect 11190 19660 11210 20040
rect 11590 19660 11610 20040
rect 11990 19660 12010 20040
rect 12390 19660 12410 20040
rect 12790 19660 12810 20040
rect 13190 19660 13210 20040
rect 13590 19660 13610 20040
rect 13990 19660 14010 20040
rect 14390 19660 14410 20040
rect 14790 19660 14810 20040
rect 15190 19660 15210 20040
rect 15590 19660 16000 20040
rect 0 19640 16000 19660
rect 0 19260 410 19640
rect 790 19260 810 19640
rect 1190 19260 1210 19640
rect 1590 19260 1610 19640
rect 1990 19260 2010 19640
rect 2390 19260 2410 19640
rect 2790 19260 2810 19640
rect 3190 19260 3210 19640
rect 3590 19260 3610 19640
rect 3990 19260 4010 19640
rect 4390 19260 4410 19640
rect 4790 19260 4810 19640
rect 5190 19260 5210 19640
rect 5590 19260 5610 19640
rect 5990 19260 6010 19640
rect 6390 19260 6410 19640
rect 6790 19260 6810 19640
rect 7190 19260 7210 19640
rect 7590 19260 7610 19640
rect 7990 19260 8010 19640
rect 8390 19260 8410 19640
rect 8790 19260 8810 19640
rect 9190 19260 9210 19640
rect 9590 19260 9610 19640
rect 9990 19260 10010 19640
rect 10390 19260 10410 19640
rect 10790 19260 10810 19640
rect 11190 19260 11210 19640
rect 11590 19260 11610 19640
rect 11990 19260 12010 19640
rect 12390 19260 12410 19640
rect 12790 19260 12810 19640
rect 13190 19260 13210 19640
rect 13590 19260 13610 19640
rect 13990 19260 14010 19640
rect 14390 19260 14410 19640
rect 14790 19260 14810 19640
rect 15190 19260 15210 19640
rect 15590 19260 16000 19640
rect 0 19000 16000 19260
rect 1500 18000 5166 19000
rect 6166 18000 9832 19000
rect 10834 18000 14500 19000
rect 0 17740 16000 18000
rect 0 17360 410 17740
rect 790 17360 810 17740
rect 1190 17360 1210 17740
rect 1590 17360 1610 17740
rect 1990 17360 2010 17740
rect 2390 17360 2410 17740
rect 2790 17360 2810 17740
rect 3190 17360 3210 17740
rect 3590 17360 3610 17740
rect 3990 17360 4010 17740
rect 4390 17360 4410 17740
rect 4790 17360 4810 17740
rect 5190 17360 5210 17740
rect 5590 17360 5610 17740
rect 5990 17360 6010 17740
rect 6390 17360 6410 17740
rect 6790 17360 6810 17740
rect 7190 17360 7210 17740
rect 7590 17360 7610 17740
rect 7990 17360 8010 17740
rect 8390 17360 8410 17740
rect 8790 17360 8810 17740
rect 9190 17360 9210 17740
rect 9590 17360 9610 17740
rect 9990 17360 10010 17740
rect 10390 17360 10410 17740
rect 10790 17360 10810 17740
rect 11190 17360 11210 17740
rect 11590 17360 11610 17740
rect 11990 17360 12010 17740
rect 12390 17360 12410 17740
rect 12790 17360 12810 17740
rect 13190 17360 13210 17740
rect 13590 17360 13610 17740
rect 13990 17360 14010 17740
rect 14390 17360 14410 17740
rect 14790 17360 14810 17740
rect 15190 17360 15210 17740
rect 15590 17360 16000 17740
rect 0 17340 16000 17360
rect 0 16960 410 17340
rect 790 16960 810 17340
rect 1190 16960 1210 17340
rect 1590 16960 1610 17340
rect 1990 16960 2010 17340
rect 2390 16960 2410 17340
rect 2790 16960 2810 17340
rect 3190 16960 3210 17340
rect 3590 16960 3610 17340
rect 3990 16960 4010 17340
rect 4390 16960 4410 17340
rect 4790 16960 4810 17340
rect 5190 16960 5210 17340
rect 5590 16960 5610 17340
rect 5990 16960 6010 17340
rect 6390 16960 6410 17340
rect 6790 16960 6810 17340
rect 7190 16960 7210 17340
rect 7590 16960 7610 17340
rect 7990 16960 8010 17340
rect 8390 16960 8410 17340
rect 8790 16960 8810 17340
rect 9190 16960 9210 17340
rect 9590 16960 9610 17340
rect 9990 16960 10010 17340
rect 10390 16960 10410 17340
rect 10790 16960 10810 17340
rect 11190 16960 11210 17340
rect 11590 16960 11610 17340
rect 11990 16960 12010 17340
rect 12390 16960 12410 17340
rect 12790 16960 12810 17340
rect 13190 16960 13210 17340
rect 13590 16960 13610 17340
rect 13990 16960 14010 17340
rect 14390 16960 14410 17340
rect 14790 16960 14810 17340
rect 15190 16960 15210 17340
rect 15590 16960 16000 17340
rect 0 16940 16000 16960
rect 0 16560 410 16940
rect 790 16560 810 16940
rect 1190 16560 1210 16940
rect 1590 16560 1610 16940
rect 1990 16560 2010 16940
rect 2390 16560 2410 16940
rect 2790 16560 2810 16940
rect 3190 16560 3210 16940
rect 3590 16560 3610 16940
rect 3990 16560 4010 16940
rect 4390 16560 4410 16940
rect 4790 16560 4810 16940
rect 5190 16560 5210 16940
rect 5590 16560 5610 16940
rect 5990 16560 6010 16940
rect 6390 16560 6410 16940
rect 6790 16560 6810 16940
rect 7190 16560 7210 16940
rect 7590 16560 7610 16940
rect 7990 16560 8010 16940
rect 8390 16560 8410 16940
rect 8790 16560 8810 16940
rect 9190 16560 9210 16940
rect 9590 16560 9610 16940
rect 9990 16560 10010 16940
rect 10390 16560 10410 16940
rect 10790 16560 10810 16940
rect 11190 16560 11210 16940
rect 11590 16560 11610 16940
rect 11990 16560 12010 16940
rect 12390 16560 12410 16940
rect 12790 16560 12810 16940
rect 13190 16560 13210 16940
rect 13590 16560 13610 16940
rect 13990 16560 14010 16940
rect 14390 16560 14410 16940
rect 14790 16560 14810 16940
rect 15190 16560 15210 16940
rect 15590 16560 16000 16940
rect 0 16540 16000 16560
rect 0 16160 410 16540
rect 790 16160 810 16540
rect 1190 16160 1210 16540
rect 1590 16160 1610 16540
rect 1990 16160 2010 16540
rect 2390 16160 2410 16540
rect 2790 16160 2810 16540
rect 3190 16160 3210 16540
rect 3590 16160 3610 16540
rect 3990 16160 4010 16540
rect 4390 16160 4410 16540
rect 4790 16160 4810 16540
rect 5190 16160 5210 16540
rect 5590 16160 5610 16540
rect 5990 16160 6010 16540
rect 6390 16160 6410 16540
rect 6790 16160 6810 16540
rect 7190 16160 7210 16540
rect 7590 16160 7610 16540
rect 7990 16160 8010 16540
rect 8390 16160 8410 16540
rect 8790 16160 8810 16540
rect 9190 16160 9210 16540
rect 9590 16160 9610 16540
rect 9990 16160 10010 16540
rect 10390 16160 10410 16540
rect 10790 16160 10810 16540
rect 11190 16160 11210 16540
rect 11590 16160 11610 16540
rect 11990 16160 12010 16540
rect 12390 16160 12410 16540
rect 12790 16160 12810 16540
rect 13190 16160 13210 16540
rect 13590 16160 13610 16540
rect 13990 16160 14010 16540
rect 14390 16160 14410 16540
rect 14790 16160 14810 16540
rect 15190 16160 15210 16540
rect 15590 16160 16000 16540
rect 0 16140 16000 16160
rect 0 15760 410 16140
rect 790 15760 810 16140
rect 1190 15760 1210 16140
rect 1590 15760 1610 16140
rect 1990 15760 2010 16140
rect 2390 15760 2410 16140
rect 2790 15760 2810 16140
rect 3190 15760 3210 16140
rect 3590 15760 3610 16140
rect 3990 15760 4010 16140
rect 4390 15760 4410 16140
rect 4790 15760 4810 16140
rect 5190 15760 5210 16140
rect 5590 15760 5610 16140
rect 5990 15760 6010 16140
rect 6390 15760 6410 16140
rect 6790 15760 6810 16140
rect 7190 15760 7210 16140
rect 7590 15760 7610 16140
rect 7990 15760 8010 16140
rect 8390 15760 8410 16140
rect 8790 15760 8810 16140
rect 9190 15760 9210 16140
rect 9590 15760 9610 16140
rect 9990 15760 10010 16140
rect 10390 15760 10410 16140
rect 10790 15760 10810 16140
rect 11190 15760 11210 16140
rect 11590 15760 11610 16140
rect 11990 15760 12010 16140
rect 12390 15760 12410 16140
rect 12790 15760 12810 16140
rect 13190 15760 13210 16140
rect 13590 15760 13610 16140
rect 13990 15760 14010 16140
rect 14390 15760 14410 16140
rect 14790 15760 14810 16140
rect 15190 15760 15210 16140
rect 15590 15760 16000 16140
rect 0 15740 16000 15760
rect 0 15360 410 15740
rect 790 15360 810 15740
rect 1190 15360 1210 15740
rect 1590 15360 1610 15740
rect 1990 15360 2010 15740
rect 2390 15360 2410 15740
rect 2790 15360 2810 15740
rect 3190 15360 3210 15740
rect 3590 15360 3610 15740
rect 3990 15360 4010 15740
rect 4390 15360 4410 15740
rect 4790 15360 4810 15740
rect 5190 15360 5210 15740
rect 5590 15360 5610 15740
rect 5990 15360 6010 15740
rect 6390 15360 6410 15740
rect 6790 15360 6810 15740
rect 7190 15360 7210 15740
rect 7590 15360 7610 15740
rect 7990 15360 8010 15740
rect 8390 15360 8410 15740
rect 8790 15360 8810 15740
rect 9190 15360 9210 15740
rect 9590 15360 9610 15740
rect 9990 15360 10010 15740
rect 10390 15360 10410 15740
rect 10790 15360 10810 15740
rect 11190 15360 11210 15740
rect 11590 15360 11610 15740
rect 11990 15360 12010 15740
rect 12390 15360 12410 15740
rect 12790 15360 12810 15740
rect 13190 15360 13210 15740
rect 13590 15360 13610 15740
rect 13990 15360 14010 15740
rect 14390 15360 14410 15740
rect 14790 15360 14810 15740
rect 15190 15360 15210 15740
rect 15590 15360 16000 15740
rect 0 15340 16000 15360
rect 0 14960 410 15340
rect 790 14960 810 15340
rect 1190 14960 1210 15340
rect 1590 14960 1610 15340
rect 1990 14960 2010 15340
rect 2390 14960 2410 15340
rect 2790 14960 2810 15340
rect 3190 14960 3210 15340
rect 3590 14960 3610 15340
rect 3990 14960 4010 15340
rect 4390 14960 4410 15340
rect 4790 14960 4810 15340
rect 5190 14960 5210 15340
rect 5590 14960 5610 15340
rect 5990 14960 6010 15340
rect 6390 14960 6410 15340
rect 6790 14960 6810 15340
rect 7190 14960 7210 15340
rect 7590 14960 7610 15340
rect 7990 14960 8010 15340
rect 8390 14960 8410 15340
rect 8790 14960 8810 15340
rect 9190 14960 9210 15340
rect 9590 14960 9610 15340
rect 9990 14960 10010 15340
rect 10390 14960 10410 15340
rect 10790 14960 10810 15340
rect 11190 14960 11210 15340
rect 11590 14960 11610 15340
rect 11990 14960 12010 15340
rect 12390 14960 12410 15340
rect 12790 14960 12810 15340
rect 13190 14960 13210 15340
rect 13590 14960 13610 15340
rect 13990 14960 14010 15340
rect 14390 14960 14410 15340
rect 14790 14960 14810 15340
rect 15190 14960 15210 15340
rect 15590 14960 16000 15340
rect 0 14940 16000 14960
rect 0 14560 410 14940
rect 790 14560 810 14940
rect 1190 14560 1210 14940
rect 1590 14560 1610 14940
rect 1990 14560 2010 14940
rect 2390 14560 2410 14940
rect 2790 14560 2810 14940
rect 3190 14560 3210 14940
rect 3590 14560 3610 14940
rect 3990 14560 4010 14940
rect 4390 14560 4410 14940
rect 4790 14560 4810 14940
rect 5190 14560 5210 14940
rect 5590 14560 5610 14940
rect 5990 14560 6010 14940
rect 6390 14560 6410 14940
rect 6790 14560 6810 14940
rect 7190 14560 7210 14940
rect 7590 14560 7610 14940
rect 7990 14560 8010 14940
rect 8390 14560 8410 14940
rect 8790 14560 8810 14940
rect 9190 14560 9210 14940
rect 9590 14560 9610 14940
rect 9990 14560 10010 14940
rect 10390 14560 10410 14940
rect 10790 14560 10810 14940
rect 11190 14560 11210 14940
rect 11590 14560 11610 14940
rect 11990 14560 12010 14940
rect 12390 14560 12410 14940
rect 12790 14560 12810 14940
rect 13190 14560 13210 14940
rect 13590 14560 13610 14940
rect 13990 14560 14010 14940
rect 14390 14560 14410 14940
rect 14790 14560 14810 14940
rect 15190 14560 15210 14940
rect 15590 14560 16000 14940
rect 0 14540 16000 14560
rect 0 14160 410 14540
rect 790 14160 810 14540
rect 1190 14160 1210 14540
rect 1590 14160 1610 14540
rect 1990 14160 2010 14540
rect 2390 14160 2410 14540
rect 2790 14160 2810 14540
rect 3190 14160 3210 14540
rect 3590 14160 3610 14540
rect 3990 14160 4010 14540
rect 4390 14160 4410 14540
rect 4790 14160 4810 14540
rect 5190 14160 5210 14540
rect 5590 14160 5610 14540
rect 5990 14160 6010 14540
rect 6390 14160 6410 14540
rect 6790 14160 6810 14540
rect 7190 14160 7210 14540
rect 7590 14160 7610 14540
rect 7990 14160 8010 14540
rect 8390 14160 8410 14540
rect 8790 14160 8810 14540
rect 9190 14160 9210 14540
rect 9590 14160 9610 14540
rect 9990 14160 10010 14540
rect 10390 14160 10410 14540
rect 10790 14160 10810 14540
rect 11190 14160 11210 14540
rect 11590 14160 11610 14540
rect 11990 14160 12010 14540
rect 12390 14160 12410 14540
rect 12790 14160 12810 14540
rect 13190 14160 13210 14540
rect 13590 14160 13610 14540
rect 13990 14160 14010 14540
rect 14390 14160 14410 14540
rect 14790 14160 14810 14540
rect 15190 14160 15210 14540
rect 15590 14160 16000 14540
rect 0 14140 16000 14160
rect 0 13760 410 14140
rect 790 13760 810 14140
rect 1190 13760 1210 14140
rect 1590 13760 1610 14140
rect 1990 13760 2010 14140
rect 2390 13760 2410 14140
rect 2790 13760 2810 14140
rect 3190 13760 3210 14140
rect 3590 13760 3610 14140
rect 3990 13760 4010 14140
rect 4390 13760 4410 14140
rect 4790 13760 4810 14140
rect 5190 13760 5210 14140
rect 5590 13760 5610 14140
rect 5990 13760 6010 14140
rect 6390 13760 6410 14140
rect 6790 13760 6810 14140
rect 7190 13760 7210 14140
rect 7590 13760 7610 14140
rect 7990 13760 8010 14140
rect 8390 13760 8410 14140
rect 8790 13760 8810 14140
rect 9190 13760 9210 14140
rect 9590 13760 9610 14140
rect 9990 13760 10010 14140
rect 10390 13760 10410 14140
rect 10790 13760 10810 14140
rect 11190 13760 11210 14140
rect 11590 13760 11610 14140
rect 11990 13760 12010 14140
rect 12390 13760 12410 14140
rect 12790 13760 12810 14140
rect 13190 13760 13210 14140
rect 13590 13760 13610 14140
rect 13990 13760 14010 14140
rect 14390 13760 14410 14140
rect 14790 13760 14810 14140
rect 15190 13760 15210 14140
rect 15590 13760 16000 14140
rect 0 13500 16000 13760
rect 0 11640 780 11700
rect 380 11260 400 11640
rect 0 11240 780 11260
rect 380 10860 400 11240
rect 0 10840 780 10860
rect 380 10460 400 10840
rect 0 10440 780 10460
rect 380 10060 400 10440
rect 0 10040 780 10060
rect 380 9660 400 10040
rect 0 9640 780 9660
rect 380 9260 400 9640
rect 0 9240 780 9260
rect 380 8860 400 9240
rect 0 8840 780 8860
rect 380 8460 400 8840
rect 0 8440 780 8460
rect 380 8060 400 8440
rect 0 8040 780 8060
rect 380 7660 400 8040
rect 0 7640 780 7660
rect 380 7260 400 7640
rect 0 7200 780 7260
rect 0 6140 780 6200
rect 380 5760 400 6140
rect 0 5740 780 5760
rect 380 5360 400 5740
rect 0 5340 780 5360
rect 380 4960 400 5340
rect 0 4940 780 4960
rect 380 4560 400 4940
rect 0 4540 780 4560
rect 380 4160 400 4540
rect 0 4140 780 4160
rect 380 3760 400 4140
rect 0 3740 780 3760
rect 380 3360 400 3740
rect 0 3340 780 3360
rect 380 2960 400 3340
rect 0 2940 780 2960
rect 380 2560 400 2940
rect 0 2540 780 2560
rect 380 2160 400 2540
rect 0 2140 780 2160
rect 380 1760 400 2140
rect 0 1700 780 1760
rect 1500 600 5166 13500
rect 6166 600 9832 13500
rect 10834 600 14500 13500
rect 15220 11640 16000 11700
rect 15600 11260 15620 11640
rect 15220 11240 16000 11260
rect 15600 10860 15620 11240
rect 15220 10840 16000 10860
rect 15600 10460 15620 10840
rect 15220 10440 16000 10460
rect 15600 10060 15620 10440
rect 15220 10040 16000 10060
rect 15600 9660 15620 10040
rect 15220 9640 16000 9660
rect 15600 9260 15620 9640
rect 15220 9240 16000 9260
rect 15600 8860 15620 9240
rect 15220 8840 16000 8860
rect 15600 8460 15620 8840
rect 15220 8440 16000 8460
rect 15600 8060 15620 8440
rect 15220 8040 16000 8060
rect 15600 7660 15620 8040
rect 15220 7640 16000 7660
rect 15600 7260 15620 7640
rect 15220 7200 16000 7260
rect 15220 6140 16000 6200
rect 15600 5760 15620 6140
rect 15220 5740 16000 5760
rect 15600 5360 15620 5740
rect 15220 5340 16000 5360
rect 15600 4960 15620 5340
rect 15220 4940 16000 4960
rect 15600 4560 15620 4940
rect 15220 4540 16000 4560
rect 15600 4160 15620 4540
rect 15220 4140 16000 4160
rect 15600 3760 15620 4140
rect 15220 3740 16000 3760
rect 15600 3360 15620 3740
rect 15220 3340 16000 3360
rect 15600 2960 15620 3340
rect 15220 2940 16000 2960
rect 15600 2560 15620 2940
rect 15220 2540 16000 2560
rect 15600 2160 15620 2540
rect 15220 2140 16000 2160
rect 15600 1760 15620 2140
rect 15220 1700 16000 1760
rect 1000 490 15000 600
rect 1000 110 1010 490
rect 1390 110 1410 490
rect 1790 110 1810 490
rect 2190 110 2210 490
rect 2590 110 2610 490
rect 2990 110 3010 490
rect 3390 110 3410 490
rect 3790 110 3810 490
rect 4190 110 4210 490
rect 4590 110 4610 490
rect 4990 110 5010 490
rect 5390 110 5410 490
rect 5790 110 5810 490
rect 6190 110 6210 490
rect 6590 110 6610 490
rect 6990 110 7010 490
rect 7390 110 7410 490
rect 7790 110 7810 490
rect 8190 110 8210 490
rect 8590 110 8610 490
rect 8990 110 9010 490
rect 9390 110 9410 490
rect 9790 110 9810 490
rect 10190 110 10210 490
rect 10590 110 10610 490
rect 10990 110 11010 490
rect 11390 110 11410 490
rect 11790 110 11810 490
rect 12190 110 12210 490
rect 12590 110 12610 490
rect 12990 110 13010 490
rect 13390 110 13410 490
rect 13790 110 13810 490
rect 14190 110 14210 490
rect 14590 110 14610 490
rect 14990 110 15000 490
rect 1000 0 15000 110
use sg13g2_Clamp_N43N43D4R  sg13g2_Clamp_N43N43D4R_0
timestamp 1755542813
transform 1 0 0 0 1 1200
box -124 -124 16124 5008
use sg13g2_RCClampInverter  sg13g2_RCClampInverter_0
timestamp 1755542813
transform -1 0 16000 0 1 13000
box -26 -26 16026 7214
use sg13g2_RCClampResistor  sg13g2_RCClampResistor_0
timestamp 1755542813
transform 1 0 3775 0 -1 11628
box 0 -2 8450 4174
<< labels >>
rlabel metal2 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal3 s 0 32000 16000 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 16000 31600 4 vss
port 1 nsew
rlabel metal3 s 0 13200 16000 18300 4 iovdd
port 4 nsew
rlabel metal3 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal3 s 0 18700 16000 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 6900 16000 12000 4 iovss
port 3 nsew
rlabel metal3 s 0 25200 16000 26800 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 16000 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 16000 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 16000 35600 4 vss
port 1 nsew
rlabel metal4 s 0 13200 16000 18300 4 iovdd
port 4 nsew
rlabel metal4 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal4 s 0 18700 16000 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 6900 16000 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 25200 16000 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 16000 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 16000 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 16000 35600 4 vss
port 1 nsew
rlabel metal5 s 0 13200 16000 18300 4 iovdd
port 4 nsew
rlabel metal5 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal5 s 0 18700 16000 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 6900 16000 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 25200 16000 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 16000 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 16000 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 16000 35600 4 vss
port 1 nsew
rlabel metal6 s 0 13200 16000 18300 4 iovdd
port 4 nsew
rlabel metal6 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal6 s 0 18700 16000 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 6900 16000 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 25200 16000 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 16000 6500 4 iovss
port 3 nsew
rlabel metal7 s 1000 0 15000 600 4 iovdd
port 4 nsew
rlabel metal7 s 0 19000 16000 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 13500 16000 18000 4 iovdd
port 4 nsew
rlabel metal7 s 15220 1700 16000 6200 4 iovss
port 3 nsew
rlabel metal7 s 0 25500 16000 26500 4 iovss
port 3 nsew
rlabel metal7 s 15220 7200 16000 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 1700 780 6200 4 iovss
port 3 nsew
rlabel metal7 s 0 7200 780 11700 4 iovss
port 3 nsew
flabel comment s 15626 31404 15626 31404 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string FIXED_BBOX 0 0 16000 36000
string GDS_END 4087230
string GDS_FILE sg13g2_io.gds
string GDS_START 2434280
<< end >>
