magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752936403
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 23 56 543 292
rect -26 -56 602 56
<< nmos >>
rect 117 118 143 266
rect 219 118 245 266
rect 321 118 347 266
rect 423 118 449 266
<< pmos >>
rect 117 412 143 636
rect 219 412 245 636
rect 321 412 347 636
rect 423 412 449 636
<< ndiff >>
rect 49 232 117 266
rect 49 200 63 232
rect 95 200 117 232
rect 49 164 117 200
rect 49 132 63 164
rect 95 132 117 164
rect 49 118 117 132
rect 143 232 219 266
rect 143 200 165 232
rect 197 200 219 232
rect 143 164 219 200
rect 143 132 165 164
rect 197 132 219 164
rect 143 118 219 132
rect 245 164 321 266
rect 245 132 267 164
rect 299 132 321 164
rect 245 118 321 132
rect 347 232 423 266
rect 347 200 369 232
rect 401 200 423 232
rect 347 164 423 200
rect 347 132 369 164
rect 401 132 423 164
rect 347 118 423 132
rect 449 164 517 266
rect 449 132 471 164
rect 503 132 517 164
rect 449 118 517 132
<< pdiff >>
rect 49 621 117 636
rect 49 589 63 621
rect 95 589 117 621
rect 49 553 117 589
rect 49 521 63 553
rect 95 521 117 553
rect 49 483 117 521
rect 49 451 63 483
rect 95 451 117 483
rect 49 412 117 451
rect 143 621 219 636
rect 143 589 165 621
rect 197 589 219 621
rect 143 553 219 589
rect 143 521 165 553
rect 197 521 219 553
rect 143 483 219 521
rect 143 451 165 483
rect 197 451 219 483
rect 143 412 219 451
rect 245 621 321 636
rect 245 589 267 621
rect 299 589 321 621
rect 245 551 321 589
rect 245 519 267 551
rect 299 519 321 551
rect 245 412 321 519
rect 347 621 423 636
rect 347 589 369 621
rect 401 589 423 621
rect 347 553 423 589
rect 347 521 369 553
rect 401 521 423 553
rect 347 483 423 521
rect 347 451 369 483
rect 401 451 423 483
rect 347 412 423 451
rect 449 621 517 636
rect 449 589 471 621
rect 503 589 517 621
rect 449 551 517 589
rect 449 519 471 551
rect 503 519 517 551
rect 449 412 517 519
<< ndiffc >>
rect 63 200 95 232
rect 63 132 95 164
rect 165 200 197 232
rect 165 132 197 164
rect 267 132 299 164
rect 369 200 401 232
rect 369 132 401 164
rect 471 132 503 164
<< pdiffc >>
rect 63 589 95 621
rect 63 521 95 553
rect 63 451 95 483
rect 165 589 197 621
rect 165 521 197 553
rect 165 451 197 483
rect 267 589 299 621
rect 267 519 299 551
rect 369 589 401 621
rect 369 521 401 553
rect 369 451 401 483
rect 471 589 503 621
rect 471 519 503 551
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 117 636 143 672
rect 219 636 245 672
rect 321 636 347 672
rect 423 636 449 672
rect 117 380 143 412
rect 219 380 245 412
rect 321 380 347 412
rect 423 380 449 412
rect 117 363 449 380
rect 117 331 147 363
rect 179 331 215 363
rect 247 331 283 363
rect 315 331 351 363
rect 383 331 449 363
rect 117 314 449 331
rect 117 266 143 314
rect 219 266 245 314
rect 321 266 347 314
rect 423 266 449 314
rect 117 82 143 118
rect 219 82 245 118
rect 321 82 347 118
rect 423 82 449 118
<< polycont >>
rect 147 331 179 363
rect 215 331 247 363
rect 283 331 315 363
rect 351 331 383 363
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 53 621 105 712
rect 53 589 63 621
rect 95 589 105 621
rect 53 553 105 589
rect 53 521 63 553
rect 95 521 105 553
rect 53 483 105 521
rect 53 451 63 483
rect 95 451 105 483
rect 53 441 105 451
rect 155 621 207 631
rect 155 589 165 621
rect 197 589 207 621
rect 155 553 207 589
rect 155 521 165 553
rect 197 521 207 553
rect 155 483 207 521
rect 257 621 309 712
rect 257 589 267 621
rect 299 589 309 621
rect 257 551 309 589
rect 257 519 267 551
rect 299 519 309 551
rect 257 509 309 519
rect 359 621 411 631
rect 359 589 369 621
rect 401 589 411 621
rect 359 553 411 589
rect 359 521 369 553
rect 401 521 411 553
rect 155 451 165 483
rect 197 468 207 483
rect 359 483 411 521
rect 461 621 513 712
rect 461 589 471 621
rect 503 589 513 621
rect 461 551 513 589
rect 461 519 471 551
rect 503 519 513 551
rect 461 509 513 519
rect 359 468 369 483
rect 197 451 369 468
rect 401 468 411 483
rect 401 451 508 468
rect 155 434 508 451
rect 96 363 400 380
rect 96 331 147 363
rect 179 331 215 363
rect 247 331 283 363
rect 315 331 351 363
rect 383 331 400 363
rect 96 304 400 331
rect 449 242 508 434
rect 53 232 105 242
rect 53 200 63 232
rect 95 200 105 232
rect 53 164 105 200
rect 53 132 63 164
rect 95 132 105 164
rect 53 44 105 132
rect 155 232 508 242
rect 155 200 165 232
rect 197 210 369 232
rect 197 200 207 210
rect 155 164 207 200
rect 359 200 369 210
rect 401 210 508 232
rect 401 200 411 210
rect 155 132 165 164
rect 197 132 207 164
rect 155 122 207 132
rect 256 164 310 174
rect 256 132 267 164
rect 299 132 310 164
rect 256 44 310 132
rect 359 164 411 200
rect 359 132 369 164
rect 401 132 411 164
rect 359 122 411 132
rect 461 164 513 174
rect 461 132 471 164
rect 503 132 513 164
rect 461 44 513 132
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 96 304 400 380 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 449 210 508 468 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 328610
string GDS_FILE sg13g2_stdcell.gds
string GDS_START 323594
<< end >>
