magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 31 56 560 285
rect -26 -56 602 56
<< nmos >>
rect 132 115 158 259
rect 234 115 260 259
rect 338 115 364 259
rect 440 115 466 259
<< pmos >>
rect 132 412 158 636
rect 234 412 260 636
rect 338 412 364 636
rect 440 412 466 636
<< ndiff >>
rect 57 230 132 259
rect 57 198 75 230
rect 107 198 132 230
rect 57 162 132 198
rect 57 130 76 162
rect 108 130 132 162
rect 57 115 132 130
rect 158 161 234 259
rect 158 129 180 161
rect 212 129 234 161
rect 158 115 234 129
rect 260 233 338 259
rect 260 201 282 233
rect 314 201 338 233
rect 260 164 338 201
rect 260 132 282 164
rect 314 132 338 164
rect 260 115 338 132
rect 364 242 440 259
rect 364 210 386 242
rect 418 210 440 242
rect 364 115 440 210
rect 466 230 534 259
rect 466 198 488 230
rect 520 198 534 230
rect 466 162 534 198
rect 466 130 488 162
rect 520 130 534 162
rect 466 115 534 130
<< pdiff >>
rect 60 622 132 636
rect 60 590 74 622
rect 106 590 132 622
rect 60 540 132 590
rect 60 508 74 540
rect 106 508 132 540
rect 60 458 132 508
rect 60 426 74 458
rect 106 426 132 458
rect 60 412 132 426
rect 158 622 234 636
rect 158 590 180 622
rect 212 590 234 622
rect 158 542 234 590
rect 158 510 180 542
rect 212 510 234 542
rect 158 412 234 510
rect 260 622 338 636
rect 260 590 282 622
rect 314 590 338 622
rect 260 412 338 590
rect 364 622 440 636
rect 364 590 386 622
rect 418 590 440 622
rect 364 542 440 590
rect 364 510 386 542
rect 418 510 440 542
rect 364 412 440 510
rect 466 622 536 636
rect 466 590 488 622
rect 520 590 536 622
rect 466 542 536 590
rect 466 510 488 542
rect 520 510 536 542
rect 466 474 536 510
rect 466 442 488 474
rect 520 442 536 474
rect 466 412 536 442
<< ndiffc >>
rect 75 198 107 230
rect 76 130 108 162
rect 180 129 212 161
rect 282 201 314 233
rect 282 132 314 164
rect 386 210 418 242
rect 488 198 520 230
rect 488 130 520 162
<< pdiffc >>
rect 74 590 106 622
rect 74 508 106 540
rect 74 426 106 458
rect 180 590 212 622
rect 180 510 212 542
rect 282 590 314 622
rect 386 590 418 622
rect 386 510 418 542
rect 488 590 520 622
rect 488 510 520 542
rect 488 442 520 474
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 132 636 158 672
rect 234 636 260 672
rect 338 636 364 672
rect 440 636 466 672
rect 132 375 158 412
rect 234 375 260 412
rect 132 360 260 375
rect 132 328 180 360
rect 212 328 260 360
rect 132 313 260 328
rect 132 259 158 313
rect 234 259 260 313
rect 338 398 364 412
rect 440 398 466 412
rect 338 384 466 398
rect 338 352 386 384
rect 418 352 466 384
rect 338 338 466 352
rect 338 259 364 338
rect 440 259 466 338
rect 132 79 158 115
rect 234 79 260 115
rect 338 79 364 115
rect 440 79 466 115
<< polycont >>
rect 180 328 212 360
rect 386 352 418 384
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 64 622 116 712
rect 64 590 74 622
rect 106 590 116 622
rect 64 540 116 590
rect 64 508 74 540
rect 106 508 116 540
rect 64 458 116 508
rect 170 622 222 632
rect 170 590 180 622
rect 212 590 222 622
rect 170 544 222 590
rect 272 622 324 712
rect 272 590 282 622
rect 314 590 324 622
rect 272 580 324 590
rect 376 622 428 632
rect 376 590 386 622
rect 418 590 428 622
rect 376 544 428 590
rect 170 542 428 544
rect 170 510 180 542
rect 212 510 386 542
rect 418 510 428 542
rect 170 500 428 510
rect 478 622 530 712
rect 478 590 488 622
rect 520 590 530 622
rect 478 542 530 590
rect 478 510 488 542
rect 520 510 530 542
rect 64 426 74 458
rect 106 426 116 458
rect 64 416 116 426
rect 164 360 220 380
rect 164 328 180 360
rect 212 328 220 360
rect 164 287 220 328
rect 264 310 312 500
rect 478 474 530 510
rect 358 396 410 464
rect 478 442 488 474
rect 520 442 530 474
rect 478 432 530 442
rect 358 384 434 396
rect 358 352 386 384
rect 418 352 434 384
rect 358 346 434 352
rect 264 278 428 310
rect 376 242 428 278
rect 65 233 324 240
rect 65 230 282 233
rect 65 198 75 230
rect 107 207 282 230
rect 107 198 117 207
rect 65 162 117 198
rect 270 201 282 207
rect 314 201 324 233
rect 65 130 76 162
rect 108 130 117 162
rect 65 100 117 130
rect 170 161 222 171
rect 170 129 180 161
rect 212 129 222 161
rect 170 44 222 129
rect 270 164 324 201
rect 376 210 386 242
rect 418 210 428 242
rect 376 200 428 210
rect 474 230 530 240
rect 270 132 282 164
rect 314 152 324 164
rect 474 198 488 230
rect 520 198 530 230
rect 474 162 530 198
rect 474 152 488 162
rect 314 132 488 152
rect 270 130 488 132
rect 520 130 530 162
rect 270 106 530 130
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 264 278 312 472 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 358 346 410 464 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 164 287 220 380 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 197062
string GDS_FILE 6_final.gds
string GDS_START 192320
<< end >>
