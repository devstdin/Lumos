magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< nwell >>
rect 13769 149 13958 209
rect 17333 149 17525 202
<< metal1 >>
rect 13405 13357 17939 14105
rect 13405 13179 14083 13357
rect 14161 13211 17133 13263
rect 13405 11207 14135 13179
rect 13405 10995 14083 11207
rect 15547 11175 15747 13211
rect 17159 11207 17291 13179
rect 14161 11027 17133 11175
rect 13405 9023 14135 10995
rect 13405 8811 14083 9023
rect 15547 8991 15747 11027
rect 17211 10995 17291 11207
rect 17159 9023 17291 10995
rect 14161 8843 17133 8991
rect 13405 6839 14135 8811
rect 13405 6627 14083 6839
rect 15547 6807 15747 8843
rect 17211 8811 17291 9023
rect 17159 6839 17291 8811
rect 14161 6659 17133 6807
rect 13405 4655 14135 6627
rect 13405 4443 14083 4655
rect 15547 4623 15747 6659
rect 17211 6627 17291 6839
rect 17159 4655 17291 6627
rect 14161 4475 17133 4623
rect 13405 2471 14135 4443
rect 13405 2259 14083 2471
rect 15547 2439 15747 4475
rect 17211 4443 17291 4655
rect 17159 2471 17291 4443
rect 14161 2291 17133 2439
rect 13405 327 14135 2259
rect 13897 287 14135 327
rect 15547 255 15747 2291
rect 17211 2259 17291 2471
rect 17159 287 17291 2259
rect 17366 327 17939 13357
rect 14161 203 17133 255
rect 15547 138 15747 203
rect 15547 -16 15557 138
rect 15737 -16 15747 138
rect 15547 -26 15747 -16
rect 17211 149 17291 287
rect 17211 -120 17398 149
rect 17049 -637 17939 -120
<< via1 >>
rect 15557 -16 15737 138
<< metal2 >>
rect 13299 138 17938 148
rect 13299 -16 15557 138
rect 15737 -16 17938 138
rect 13299 -26 17938 -16
use hvpmos_NE86AY  hvpmos_NE86AY_4
timestamp 1757240632
transform 1 0 15647 0 1 1273
box -1878 -1124 1878 12229
<< labels >>
flabel metal2 17545 -26 17938 148 0 FreeSans 800 0 0 0 VSOURCE
port 4 nsew
flabel metal1 17422 -637 17939 -120 0 FreeSans 800 0 0 0 ISOURCE
port 5 nsew
flabel metal1 17563 13544 17939 14105 0 FreeSans 800 0 0 0 VDD
port 6 nsew
<< end >>
