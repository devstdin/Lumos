magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757364080
<< nwell >>
rect -3926 2579 -3442 2618
rect 2714 1139 3709 1248
rect 3715 1143 3877 1248
rect 3776 1139 3877 1143
rect 2714 829 3877 1139
rect 2714 764 4273 829
rect 3600 -336 4272 -284
rect -3926 -1132 -3442 -1085
<< metal1 >>
rect -4492 2644 -3740 2905
rect -4492 -1153 -4232 2644
rect -3564 2640 -1337 2905
rect -3564 2555 -3400 2640
rect -1599 2618 -1337 2640
rect -3343 2395 -2722 2564
rect -3343 -1153 -3189 2395
rect -2805 2341 -2722 2395
rect -1599 2392 4631 2618
rect -2805 1999 -2569 2341
rect -1599 2310 -1304 2392
rect 4396 2310 4631 2392
rect -2414 2241 -2342 2251
rect -2414 2197 -2404 2241
rect -2352 2197 -2342 2241
rect -2414 2187 -2342 2197
rect -2502 1999 -2456 2174
rect -2394 2101 -2362 2187
rect -2300 2177 -2227 2187
rect -2300 2111 -2290 2177
rect -2237 2111 -2227 2177
rect -2300 2101 -2227 2111
rect -2414 2049 -2342 2101
rect -2805 1845 -2135 1999
rect -2805 1505 -2569 1845
rect -2420 1743 -2348 1795
rect -2528 1701 -2456 1725
rect -2528 1649 -2518 1701
rect -2466 1649 -2456 1701
rect -2528 1625 -2456 1649
rect -2400 1607 -2368 1743
rect -2420 1597 -2348 1607
rect -2420 1554 -2410 1597
rect -2358 1554 -2348 1597
rect -2420 1544 -2348 1554
rect -2312 1505 -2266 1725
rect -2199 1505 -2135 1845
rect -2805 1351 -1725 1505
rect -2805 911 -2569 1351
rect -2420 1249 -2348 1301
rect -1998 1249 -1926 1301
rect -2525 1207 -2456 1231
rect -2525 1055 -2515 1207
rect -2466 1055 -2456 1207
rect -2525 1031 -2456 1055
rect -2400 1013 -2368 1249
rect -2420 1003 -2348 1013
rect -2420 960 -2410 1003
rect -2358 960 -2348 1003
rect -2420 950 -2348 960
rect -2312 911 -2266 1231
rect -2103 1207 -2034 1231
rect -2103 1055 -2093 1207
rect -2044 1055 -2034 1207
rect -2103 1031 -2034 1055
rect -1978 1013 -1946 1249
rect -1998 1003 -1926 1013
rect -1998 960 -1988 1003
rect -1936 960 -1926 1003
rect -1998 950 -1926 960
rect -1890 911 -1844 1227
rect -2805 757 -1725 911
rect -2805 317 -2569 757
rect -2420 655 -2348 707
rect -2142 655 -2070 707
rect -2508 613 -2456 637
rect -2508 461 -2498 613
rect -2458 461 -2456 613
rect -2508 437 -2456 461
rect -2400 419 -2368 655
rect -2420 409 -2348 419
rect -2420 364 -2410 409
rect -2358 364 -2348 409
rect -2420 354 -2348 364
rect -2312 317 -2266 637
rect -2230 613 -2178 637
rect -2230 461 -2220 613
rect -2180 461 -2178 613
rect -2230 437 -2178 461
rect -2122 419 -2090 655
rect -2142 409 -2070 419
rect -2142 364 -2132 409
rect -2080 364 -2070 409
rect -2142 354 -2070 364
rect -2034 317 -1988 637
rect -1921 317 -1725 757
rect -1599 821 -1402 2310
rect 1354 1896 1646 1953
rect 1354 1807 1508 1896
rect 3814 1796 3891 1946
rect 4434 1907 4631 2310
rect 4386 1554 4631 1642
rect -399 1321 -338 1331
rect -1292 1274 -1207 1284
rect -1292 1218 -1282 1274
rect -1217 1218 -1207 1274
rect -863 1218 -559 1294
rect -399 1229 -389 1321
rect -348 1229 -338 1321
rect 3701 1359 3785 1369
rect -399 1219 -338 1229
rect 2576 1289 2647 1323
rect -1292 1208 -1207 1218
rect -592 1130 -559 1218
rect 2576 1247 2789 1289
rect 2576 1227 2647 1247
rect -399 1162 -315 1172
rect -614 1120 -540 1130
rect -614 952 -604 1120
rect -550 952 -540 1120
rect -399 1032 -389 1162
rect -325 1032 -315 1162
rect 2747 1081 2789 1247
rect 3701 1143 3715 1359
rect 3775 1143 3785 1359
rect 4125 1284 4355 1294
rect 4125 1228 4301 1284
rect 4345 1228 4355 1284
rect 4125 1218 4355 1228
rect 3701 1130 3785 1143
rect 2747 1071 3679 1081
rect 2747 1039 3627 1071
rect -399 1022 -315 1032
rect 3617 988 3627 1039
rect 3669 988 3679 1071
rect 3617 978 3679 988
rect -614 942 -540 952
rect 2681 821 4225 886
rect -1599 798 4225 821
rect -1599 502 3485 798
rect 4391 631 4631 1554
rect -517 395 -145 502
rect 147 395 519 502
rect 811 395 1183 502
rect 1475 395 1847 502
rect 2139 395 2511 502
rect 2803 395 3175 502
rect -601 360 -549 369
rect -601 320 -591 360
rect -551 349 -549 360
rect -113 360 -61 369
rect -113 349 -111 360
rect -551 320 -111 349
rect -71 320 -61 360
rect -601 317 -61 320
rect -2805 163 -1167 317
rect -601 297 -549 317
rect -113 297 -61 317
rect 63 360 115 369
rect 63 320 73 360
rect 113 349 115 360
rect 551 360 603 369
rect 551 349 553 360
rect 113 320 553 349
rect 593 320 603 360
rect 63 317 603 320
rect 63 297 115 317
rect 551 297 603 317
rect 727 360 779 369
rect 727 320 737 360
rect 777 349 779 360
rect 1215 360 1267 369
rect 1215 349 1217 360
rect 777 320 1217 349
rect 1257 320 1267 360
rect 727 317 1267 320
rect 727 297 779 317
rect 1215 297 1267 317
rect 1391 360 1443 369
rect 1391 320 1401 360
rect 1441 349 1443 360
rect 1879 360 1931 369
rect 1879 349 1881 360
rect 1441 320 1881 349
rect 1921 320 1931 360
rect 1391 317 1931 320
rect 1391 297 1443 317
rect 1879 297 1931 317
rect 2055 360 2107 369
rect 2055 320 2065 360
rect 2105 349 2107 360
rect 2543 360 2595 369
rect 2543 349 2545 360
rect 2105 320 2545 349
rect 2585 320 2595 360
rect 2055 317 2595 320
rect 2055 297 2107 317
rect 2543 297 2595 317
rect 2719 360 2771 369
rect 2719 320 2729 360
rect 2769 349 2771 360
rect 3207 360 3259 369
rect 3207 349 3209 360
rect 2769 320 3209 349
rect 3249 320 3259 360
rect 2719 317 3259 320
rect 2719 297 2771 317
rect 3207 297 3259 317
rect -517 261 -145 271
rect -517 218 -507 261
rect -155 218 -145 261
rect -517 215 -145 218
rect 147 261 519 271
rect 147 218 157 261
rect 509 218 519 261
rect 147 215 519 218
rect 811 261 1183 271
rect 811 218 821 261
rect 1173 218 1183 261
rect 811 215 1183 218
rect 1475 261 1847 271
rect 1475 218 1485 261
rect 1837 218 1847 261
rect 1475 215 1847 218
rect 2139 261 2511 271
rect 2139 218 2149 261
rect 2501 218 2511 261
rect 2139 215 2511 218
rect 2803 261 3175 271
rect 2803 218 2813 261
rect 3165 218 3175 261
rect 2803 215 3175 218
rect -2805 -1153 -2569 163
rect -2420 61 -2348 113
rect -2142 61 -2070 113
rect -1864 61 -1792 113
rect -1586 61 -1514 113
rect -2508 19 -2456 43
rect -2508 -133 -2498 19
rect -2458 -133 -2456 19
rect -2508 -157 -2456 -133
rect -2400 -175 -2368 61
rect -2420 -185 -2348 -175
rect -2420 -228 -2410 -185
rect -2358 -228 -2348 -185
rect -2420 -238 -2348 -228
rect -2312 -284 -2266 43
rect -2230 19 -2178 43
rect -2230 -133 -2220 19
rect -2180 -133 -2178 19
rect -2230 -157 -2178 -133
rect -2122 -175 -2090 61
rect -2142 -185 -2070 -175
rect -2142 -228 -2132 -185
rect -2080 -228 -2070 -185
rect -2142 -238 -2070 -228
rect -2034 -284 -1988 43
rect -1952 19 -1900 43
rect -1952 -133 -1942 19
rect -1902 -133 -1900 19
rect -1952 -157 -1900 -133
rect -1844 -175 -1812 61
rect -1864 -185 -1792 -175
rect -1864 -228 -1854 -185
rect -1802 -228 -1792 -185
rect -1864 -238 -1792 -228
rect -1756 -284 -1710 43
rect -1674 19 -1622 43
rect -1674 -133 -1664 19
rect -1624 -133 -1622 19
rect -1674 -157 -1622 -133
rect -1566 -175 -1534 61
rect -1586 -185 -1514 -175
rect -1586 -228 -1576 -185
rect -1524 -228 -1514 -185
rect -1586 -238 -1514 -228
rect -1478 -284 -1432 43
rect -2420 -431 -2348 -379
rect -2508 -473 -2456 -449
rect -2508 -625 -2498 -473
rect -2458 -625 -2456 -473
rect -2508 -649 -2456 -625
rect -2400 -667 -2368 -431
rect -2312 -649 -2266 -325
rect -2142 -431 -2070 -379
rect -2230 -473 -2178 -449
rect -2230 -625 -2220 -473
rect -2180 -625 -2178 -473
rect -2230 -649 -2178 -625
rect -2122 -667 -2090 -431
rect -2034 -649 -1988 -325
rect -1864 -431 -1792 -379
rect -1952 -473 -1900 -449
rect -1952 -625 -1942 -473
rect -1902 -625 -1900 -473
rect -1952 -649 -1900 -625
rect -1844 -667 -1812 -431
rect -1756 -649 -1710 -325
rect -1586 -431 -1514 -379
rect -1674 -473 -1622 -449
rect -1674 -625 -1664 -473
rect -1624 -625 -1622 -473
rect -1674 -649 -1622 -625
rect -1566 -667 -1534 -431
rect -1478 -649 -1432 -325
rect -2420 -719 -2348 -667
rect -2420 -763 -2410 -719
rect -2358 -763 -2348 -719
rect -2420 -815 -2348 -763
rect -2142 -719 -2070 -667
rect -2142 -763 -2132 -719
rect -2080 -763 -2070 -719
rect -2142 -815 -2070 -763
rect -1864 -719 -1792 -667
rect -1864 -763 -1854 -719
rect -1802 -763 -1792 -719
rect -1864 -815 -1792 -763
rect -1586 -719 -1514 -667
rect -1586 -763 -1576 -719
rect -1524 -763 -1514 -719
rect -1586 -815 -1514 -763
rect -2508 -857 -2456 -833
rect -2508 -1009 -2498 -857
rect -2458 -1009 -2456 -857
rect -2508 -1033 -2456 -1009
rect -2400 -1051 -2368 -815
rect -2420 -1103 -2348 -1051
rect -2312 -1153 -2266 -833
rect -2230 -857 -2178 -833
rect -2230 -1009 -2220 -857
rect -2180 -1009 -2178 -857
rect -2230 -1033 -2178 -1009
rect -2122 -1051 -2090 -815
rect -2142 -1103 -2070 -1051
rect -2034 -1153 -1988 -833
rect -1952 -857 -1900 -833
rect -1952 -1009 -1942 -857
rect -1902 -1009 -1900 -857
rect -1952 -1033 -1900 -1009
rect -1844 -1051 -1812 -815
rect -1864 -1103 -1792 -1051
rect -1756 -1153 -1710 -833
rect -1674 -857 -1622 -833
rect -1674 -1009 -1664 -857
rect -1624 -1009 -1622 -857
rect -1674 -1033 -1622 -1009
rect -1566 -1051 -1534 -815
rect -1586 -1103 -1514 -1051
rect -1478 -1153 -1432 -833
rect -1365 -1153 -1167 163
rect 147 70 519 71
rect 147 25 157 70
rect 509 25 519 70
rect 147 15 519 25
rect 811 70 1183 71
rect 811 25 821 70
rect 1173 25 1183 70
rect 811 15 1183 25
rect 1475 70 1847 71
rect 1475 25 1485 70
rect 1837 25 1847 70
rect 1475 15 1847 25
rect 2139 70 2511 71
rect 2139 25 2149 70
rect 2501 25 2511 70
rect 2139 15 2511 25
rect 2803 70 3175 71
rect 2803 25 2813 70
rect 3165 25 3175 70
rect 2803 15 3175 25
rect 63 -21 115 -11
rect 63 -73 64 -21
rect 105 -31 115 -21
rect 551 -31 603 -11
rect 105 -63 603 -31
rect 105 -73 115 -63
rect 63 -83 115 -73
rect 551 -83 603 -63
rect 727 -21 779 -11
rect 727 -73 728 -21
rect 769 -31 779 -21
rect 1215 -31 1267 -11
rect 769 -63 1267 -31
rect 769 -73 779 -63
rect 727 -83 779 -73
rect 1215 -83 1267 -63
rect 1391 -21 1443 -11
rect 1391 -73 1392 -21
rect 1433 -31 1443 -21
rect 1879 -31 1931 -11
rect 1433 -63 1931 -31
rect 1433 -73 1443 -63
rect 1391 -83 1443 -73
rect 1879 -83 1931 -63
rect 2055 -21 2107 -11
rect 2055 -73 2056 -21
rect 2097 -31 2107 -21
rect 2543 -31 2595 -11
rect 2097 -63 2595 -31
rect 2097 -73 2107 -63
rect 2055 -83 2107 -73
rect 2543 -83 2595 -63
rect 2719 -21 2771 -11
rect 2719 -73 2720 -21
rect 2761 -31 2771 -21
rect 3207 -31 3259 -11
rect 2761 -63 3259 -31
rect 2761 -73 2771 -63
rect 2719 -83 2771 -73
rect 3207 -83 3259 -63
rect 147 -119 519 -109
rect 147 -163 157 -119
rect 509 -163 519 -119
rect 147 -165 519 -163
rect 811 -119 1183 -109
rect 811 -163 821 -119
rect 1173 -163 1183 -119
rect 811 -165 1183 -163
rect 1475 -119 1847 -109
rect 1475 -163 1485 -119
rect 1837 -163 1847 -119
rect 1475 -165 1847 -163
rect 2139 -119 2511 -109
rect 2139 -163 2149 -119
rect 2501 -163 2511 -119
rect 2139 -165 2511 -163
rect 2803 -119 3175 -109
rect 2803 -163 2813 -119
rect 3165 -163 3175 -119
rect 3304 -138 3485 502
rect 3648 498 4631 631
rect 3632 301 3775 311
rect 3632 82 3642 301
rect 3765 82 3775 301
rect 4124 169 4325 216
rect 3632 72 3775 82
rect 2803 -165 3175 -163
rect 3305 -172 3485 -138
rect 3305 -263 4224 -172
rect -528 -309 -436 -300
rect 1847 -305 3452 -302
rect -528 -310 -156 -309
rect -528 -355 -518 -310
rect -446 -355 -156 -310
rect 1847 -346 1863 -305
rect 2023 -346 3452 -305
rect 1847 -349 3452 -346
rect -528 -365 -156 -355
rect -612 -401 -560 -391
rect -612 -453 -611 -401
rect -570 -411 -560 -401
rect -124 -411 -72 -391
rect -570 -443 -72 -411
rect -570 -453 -560 -443
rect -612 -463 -560 -453
rect -124 -463 -72 -443
rect 147 -489 519 -486
rect -528 -499 -156 -489
rect -528 -541 -229 -499
rect -171 -541 -156 -499
rect -528 -545 -156 -541
rect 147 -532 157 -489
rect 509 -532 519 -489
rect 147 -542 519 -532
rect 811 -489 1183 -486
rect 811 -532 821 -489
rect 1173 -532 1183 -489
rect 811 -542 1183 -532
rect 1475 -489 1847 -486
rect 1475 -532 1485 -489
rect 1837 -532 1847 -489
rect 1475 -542 1847 -532
rect 2139 -489 2511 -486
rect 2139 -532 2149 -489
rect 2501 -532 2511 -489
rect 2139 -542 2511 -532
rect 2803 -489 3175 -486
rect 2803 -532 2813 -489
rect 3165 -532 3175 -489
rect 2803 -542 3175 -532
rect -239 -551 -161 -545
rect -612 -576 -560 -567
rect -612 -630 -611 -576
rect -570 -587 -560 -576
rect -124 -587 -72 -567
rect -570 -619 -72 -587
rect -570 -630 -560 -619
rect -612 -639 -560 -630
rect -124 -639 -72 -619
rect 63 -578 115 -568
rect 63 -630 64 -578
rect 105 -588 115 -578
rect 551 -588 603 -568
rect 105 -620 603 -588
rect 105 -630 115 -620
rect 63 -640 115 -630
rect 551 -640 603 -620
rect 727 -578 779 -568
rect 727 -630 728 -578
rect 769 -588 779 -578
rect 1215 -588 1267 -568
rect 769 -620 1267 -588
rect 769 -630 779 -620
rect 727 -640 779 -630
rect 1215 -640 1267 -620
rect 1391 -578 1443 -568
rect 1391 -630 1392 -578
rect 1433 -588 1443 -578
rect 1879 -588 1931 -568
rect 1433 -620 1931 -588
rect 1433 -630 1443 -620
rect 1391 -640 1443 -630
rect 1879 -640 1931 -620
rect 2055 -578 2107 -568
rect 2055 -630 2056 -578
rect 2097 -588 2107 -578
rect 2543 -588 2595 -568
rect 2097 -620 2595 -588
rect 2097 -630 2107 -620
rect 2055 -640 2107 -630
rect 2543 -640 2595 -620
rect 2719 -578 2771 -568
rect 2719 -630 2720 -578
rect 2761 -588 2771 -578
rect 3207 -588 3259 -568
rect 2761 -620 3259 -588
rect 2761 -630 2771 -620
rect 2719 -640 2771 -630
rect 3207 -640 3259 -620
rect -528 -777 -156 -665
rect 147 -675 519 -666
rect 147 -718 157 -675
rect 509 -718 519 -675
rect 147 -722 519 -718
rect 811 -675 1183 -666
rect 811 -718 821 -675
rect 1173 -718 1183 -675
rect 811 -722 1183 -718
rect 1475 -675 1847 -666
rect 1475 -718 1485 -675
rect 1837 -718 1847 -675
rect 1475 -722 1847 -718
rect 2139 -675 2511 -666
rect 2139 -718 2149 -675
rect 2501 -718 2511 -675
rect 2139 -722 2511 -718
rect 2803 -675 3175 -666
rect 2803 -718 2813 -675
rect 3165 -718 3175 -675
rect 2803 -722 3175 -718
rect 3405 -786 3452 -349
rect 3505 -446 4224 -263
rect 4278 -786 4325 169
rect 3405 -833 3748 -786
rect 4114 -833 4325 -786
rect -517 -869 -145 -866
rect -517 -912 -507 -869
rect -155 -912 -145 -869
rect -517 -922 -145 -912
rect 147 -869 519 -866
rect 147 -912 157 -869
rect 509 -912 519 -869
rect 147 -922 519 -912
rect 811 -869 1183 -866
rect 811 -912 821 -869
rect 1173 -912 1183 -869
rect 811 -922 1183 -912
rect 1475 -869 1847 -866
rect 1475 -912 1485 -869
rect 1837 -912 1847 -869
rect 1475 -922 1847 -912
rect 2139 -869 2511 -866
rect 2139 -912 2149 -869
rect 2501 -912 2511 -869
rect 2139 -922 2511 -912
rect 2803 -869 3175 -866
rect 2803 -912 2813 -869
rect 3165 -912 3175 -869
rect 2803 -922 3175 -912
rect -601 -968 -549 -948
rect -113 -968 -61 -948
rect -601 -971 -61 -968
rect -601 -1011 -591 -971
rect -551 -1000 -111 -971
rect -551 -1011 -549 -1000
rect -601 -1020 -549 -1011
rect -113 -1011 -111 -1000
rect -71 -1011 -61 -971
rect -113 -1020 -61 -1011
rect 63 -968 115 -948
rect 551 -968 603 -948
rect 63 -971 603 -968
rect 63 -1011 73 -971
rect 113 -1000 553 -971
rect 113 -1011 115 -1000
rect 63 -1020 115 -1011
rect 551 -1011 553 -1000
rect 593 -1011 603 -971
rect 551 -1020 603 -1011
rect 727 -968 779 -948
rect 1215 -968 1267 -948
rect 727 -971 1267 -968
rect 727 -1011 737 -971
rect 777 -1000 1217 -971
rect 777 -1011 779 -1000
rect 727 -1020 779 -1011
rect 1215 -1011 1217 -1000
rect 1257 -1011 1267 -971
rect 1215 -1020 1267 -1011
rect 1391 -968 1443 -948
rect 1879 -968 1931 -948
rect 1391 -971 1931 -968
rect 1391 -1011 1401 -971
rect 1441 -1000 1881 -971
rect 1441 -1011 1443 -1000
rect 1391 -1020 1443 -1011
rect 1879 -1011 1881 -1000
rect 1921 -1011 1931 -971
rect 1879 -1020 1931 -1011
rect 2055 -968 2107 -948
rect 2543 -968 2595 -948
rect 2055 -971 2595 -968
rect 2055 -1011 2065 -971
rect 2105 -1000 2545 -971
rect 2105 -1011 2107 -1000
rect 2055 -1020 2107 -1011
rect 2543 -1011 2545 -1000
rect 2585 -1011 2595 -971
rect 2543 -1020 2595 -1011
rect 2719 -968 2771 -948
rect 3207 -968 3259 -948
rect 2719 -971 3259 -968
rect 2719 -1011 2729 -971
rect 2769 -1000 3209 -971
rect 2769 -1011 2771 -1000
rect 2719 -1020 2771 -1011
rect 3207 -1011 3209 -1000
rect 3249 -1011 3259 -971
rect 4247 -971 4257 -833
rect 4315 -971 4325 -833
rect 4247 -981 4325 -971
rect 3207 -1020 3259 -1011
rect -517 -1153 -145 -1046
rect 147 -1153 519 -1046
rect 811 -1153 1183 -1046
rect 1475 -1153 1847 -1046
rect 2139 -1153 2511 -1046
rect 2803 -1153 3175 -1046
rect 4391 -1153 4631 498
rect -4492 -1414 4631 -1153
<< via1 >>
rect -2404 2197 -2352 2241
rect -2290 2111 -2237 2177
rect -2518 1649 -2466 1701
rect -2410 1554 -2358 1597
rect -2515 1055 -2466 1207
rect -2410 960 -2358 1003
rect -2093 1055 -2044 1207
rect -1988 960 -1936 1003
rect -2498 461 -2458 613
rect -2410 364 -2358 409
rect -2220 461 -2180 613
rect -2132 364 -2080 409
rect -1273 1883 -1222 1959
rect -884 1910 -794 1981
rect -51 1875 54 1975
rect 1996 1926 2086 1981
rect 2829 1866 2934 1975
rect 4250 1817 4330 1886
rect -1282 1218 -1217 1274
rect -389 1229 -348 1321
rect -134 1310 0 1379
rect 1310 1221 1415 1321
rect 2158 1215 2248 1286
rect -604 952 -550 1120
rect -389 1032 -325 1162
rect 3715 1143 3775 1359
rect 4301 1228 4345 1284
rect 3627 988 3669 1071
rect -591 320 -551 360
rect -111 320 -71 360
rect 73 320 113 360
rect 553 320 593 360
rect 737 320 777 360
rect 1217 320 1257 360
rect 1401 320 1441 360
rect 1881 320 1921 360
rect 2065 320 2105 360
rect 2545 320 2585 360
rect 2729 320 2769 360
rect 3209 320 3249 360
rect -507 218 -155 261
rect 157 218 509 261
rect 821 218 1173 261
rect 1485 218 1837 261
rect 2149 218 2501 261
rect 2813 218 3165 261
rect -2498 -133 -2458 19
rect -2410 -228 -2358 -185
rect -2220 -133 -2180 19
rect -2132 -228 -2080 -185
rect -1942 -133 -1902 19
rect -1854 -228 -1802 -185
rect -1664 -133 -1624 19
rect -1576 -228 -1524 -185
rect -2498 -625 -2458 -473
rect -2220 -625 -2180 -473
rect -1942 -625 -1902 -473
rect -1664 -625 -1624 -473
rect -2410 -763 -2358 -719
rect -2132 -763 -2080 -719
rect -1854 -763 -1802 -719
rect -1576 -763 -1524 -719
rect -2498 -1009 -2458 -857
rect -2220 -1009 -2180 -857
rect -1942 -1009 -1902 -857
rect -1664 -1009 -1624 -857
rect 157 25 509 70
rect 821 25 1173 70
rect 1485 25 1837 70
rect 2149 25 2501 70
rect 2813 25 3165 70
rect 64 -73 105 -21
rect 728 -73 769 -21
rect 1392 -73 1433 -21
rect 2056 -73 2097 -21
rect 2720 -73 2761 -21
rect 157 -163 509 -119
rect 821 -163 1173 -119
rect 1485 -163 1837 -119
rect 2149 -163 2501 -119
rect 2813 -163 3165 -119
rect 3642 82 3765 301
rect -518 -355 -446 -310
rect 1863 -346 2023 -305
rect -611 -453 -570 -401
rect -229 -541 -171 -499
rect 157 -532 509 -489
rect 821 -532 1173 -489
rect 1485 -532 1837 -489
rect 2149 -532 2501 -489
rect 2813 -532 3165 -489
rect -611 -630 -570 -576
rect 64 -630 105 -578
rect 728 -630 769 -578
rect 1392 -630 1433 -578
rect 2056 -630 2097 -578
rect 2720 -630 2761 -578
rect 157 -718 509 -675
rect 821 -718 1173 -675
rect 1485 -718 1837 -675
rect 2149 -718 2501 -675
rect 2813 -718 3165 -675
rect -507 -912 -155 -869
rect 157 -912 509 -869
rect 821 -912 1173 -869
rect 1485 -912 1837 -869
rect 2149 -912 2501 -869
rect 2813 -912 3165 -869
rect -591 -1011 -551 -971
rect -111 -1011 -71 -971
rect 73 -1011 113 -971
rect 553 -1011 593 -971
rect 737 -1011 777 -971
rect 1217 -1011 1257 -971
rect 1401 -1011 1441 -971
rect 1881 -1011 1921 -971
rect 2065 -1011 2105 -971
rect 2545 -1011 2585 -971
rect 2729 -1011 2769 -971
rect 3209 -1011 3249 -971
rect 4257 -971 4315 -833
<< metal2 >>
rect -2228 2432 -2028 2593
rect -2104 2376 -2028 2432
rect -2829 2323 -2028 2376
rect -2751 2241 -2342 2251
rect -2751 2197 -2404 2241
rect -2352 2197 -2342 2241
rect -2751 2162 -2697 2197
rect -2414 2187 -2342 2197
rect -2826 2081 -2697 2162
rect -2300 2177 -2227 2187
rect -2300 2111 -2290 2177
rect -2237 2164 -2227 2177
rect -2104 2164 -2028 2323
rect -2237 2124 -2028 2164
rect -2237 2111 -2227 2124
rect -2300 2101 -2227 2111
rect -4492 1956 -4357 2037
rect -2885 1695 -2708 1776
rect -2528 1701 -2456 1711
rect -2528 1695 -2518 1701
rect -2749 1655 -2518 1695
rect -2528 1649 -2518 1655
rect -2466 1695 -2456 1701
rect -2104 1695 -2028 2124
rect -1839 1969 -1626 2593
rect -865 2126 3701 2173
rect -865 1991 -818 2126
rect 2023 1991 2070 2126
rect -894 1981 -784 1991
rect -1839 1959 -1212 1969
rect -1839 1883 -1273 1959
rect -1222 1883 -1212 1959
rect -894 1910 -884 1981
rect -794 1910 -784 1981
rect -894 1900 -784 1910
rect -61 1975 64 1985
rect -1839 1873 -1212 1883
rect -2466 1655 -2028 1695
rect -2466 1649 -2456 1655
rect -2528 1639 -2456 1649
rect -2104 1611 -2028 1655
rect -2420 1597 -2348 1607
rect -2420 1590 -2410 1597
rect -2749 1562 -2410 1590
rect -2892 1554 -2410 1562
rect -2358 1554 -2348 1597
rect -2892 1544 -2348 1554
rect -2892 1481 -2702 1544
rect -2104 1535 -1624 1611
rect -4492 1356 -4357 1437
rect -2525 1207 -2456 1217
rect -2885 1157 -2749 1176
rect -2525 1157 -2515 1207
rect -2885 1105 -2515 1157
rect -2885 1095 -2749 1105
rect -2525 1055 -2515 1105
rect -2466 1157 -2456 1207
rect -2103 1207 -2034 1217
rect -2103 1157 -2093 1207
rect -2466 1105 -2093 1157
rect -2466 1055 -2456 1105
rect -2525 1045 -2456 1055
rect -2103 1055 -2093 1105
rect -2044 1157 -2034 1207
rect -1700 1157 -1624 1535
rect -1283 1537 -1212 1873
rect -61 1875 -51 1975
rect 54 1920 64 1975
rect 1986 1981 2096 1991
rect 1986 1926 1996 1981
rect 2086 1926 2096 1981
rect 54 1875 251 1920
rect 1986 1916 2096 1926
rect 2819 1975 2944 1985
rect -61 1871 251 1875
rect -61 1865 64 1871
rect 202 1864 251 1871
rect 202 1815 1356 1864
rect -1283 1496 -348 1537
rect -399 1331 -348 1496
rect -144 1379 10 1389
rect -399 1321 -338 1331
rect -1292 1274 -1207 1284
rect -1292 1218 -1282 1274
rect -1217 1218 -1207 1274
rect -399 1229 -389 1321
rect -348 1229 -338 1321
rect -399 1219 -338 1229
rect -144 1310 -134 1379
rect 0 1310 10 1379
rect 1307 1331 1356 1815
rect -144 1300 10 1310
rect 1300 1321 1425 1331
rect -1292 1208 -1207 1218
rect -2044 1105 -1624 1157
rect -2044 1055 -2034 1105
rect -2103 1045 -2034 1055
rect -2420 1003 -2348 1013
rect -2420 993 -2410 1003
rect -2749 962 -2410 993
rect -2885 960 -2410 962
rect -2358 960 -2348 1003
rect -2885 950 -2348 960
rect -2103 993 -2058 1045
rect -1998 1003 -1926 1013
rect -1998 993 -1988 1003
rect -2103 960 -1988 993
rect -1936 960 -1926 1003
rect -2103 950 -1926 960
rect -2885 881 -2706 950
rect -4492 756 -4357 837
rect -2508 613 -2449 623
rect -2885 563 -2749 576
rect -2508 563 -2498 613
rect -2885 511 -2498 563
rect -2885 495 -2749 511
rect -2508 461 -2498 511
rect -2458 563 -2449 613
rect -2230 613 -2171 623
rect -2230 563 -2220 613
rect -2458 511 -2220 563
rect -2458 461 -2449 511
rect -2508 451 -2449 461
rect -2230 461 -2220 511
rect -2180 563 -2171 613
rect -1700 563 -1624 1105
rect -1269 759 -1229 1208
rect -144 1172 -93 1300
rect 1300 1221 1310 1321
rect 1415 1221 1425 1321
rect 2023 1277 2070 1916
rect 2819 1866 2829 1975
rect 2934 1866 2944 1975
rect 2819 1864 2944 1866
rect 2819 1815 3569 1864
rect 2148 1286 2258 1296
rect 2148 1277 2158 1286
rect 2023 1230 2158 1277
rect 1300 1211 1425 1221
rect 2148 1215 2158 1230
rect 2248 1215 2258 1286
rect -399 1162 -93 1172
rect -614 1120 -540 1130
rect -614 952 -604 1120
rect -550 952 -540 1120
rect -399 1032 -389 1162
rect -325 1118 -93 1162
rect -325 1032 -315 1118
rect -399 1022 -315 1032
rect -614 942 -540 952
rect 1328 960 1388 1211
rect 2148 1205 2258 1215
rect 3509 960 3569 1815
rect 3654 1369 3701 2126
rect 4240 1886 4340 1896
rect 4240 1817 4250 1886
rect 4330 1817 4340 1886
rect 4240 1807 4340 1817
rect 4240 1491 4280 1807
rect 4191 1451 4280 1491
rect 3654 1359 3785 1369
rect 3654 1143 3715 1359
rect 3775 1143 3785 1359
rect 3654 1130 3785 1143
rect -1269 719 -838 759
rect -614 758 -574 942
rect 1328 900 3569 960
rect 3617 1071 3679 1081
rect 3617 988 3627 1071
rect 3669 988 3679 1071
rect 3617 941 3679 988
rect 4191 941 4231 1451
rect 4391 1294 4631 1347
rect 4291 1284 4631 1294
rect 4291 1228 4301 1284
rect 4345 1228 4631 1284
rect 4291 1218 4631 1228
rect 4391 1208 4631 1218
rect 3617 901 4231 941
rect -2180 511 -1624 563
rect -2180 461 -2171 511
rect -2230 451 -2171 461
rect -1700 423 -1624 511
rect -2420 409 -2348 419
rect -2420 398 -2410 409
rect -2749 364 -2410 398
rect -2358 398 -2348 409
rect -2142 409 -2070 419
rect -2142 398 -2132 409
rect -2358 364 -2132 398
rect -2080 364 -2070 409
rect -2749 362 -2070 364
rect -2885 354 -2070 362
rect -2885 281 -2705 354
rect -1700 347 -1066 423
rect -4492 156 -4357 237
rect -2508 19 -2449 29
rect -2885 -31 -2749 -24
rect -2508 -31 -2498 19
rect -2885 -83 -2498 -31
rect -2885 -105 -2749 -83
rect -2508 -133 -2498 -83
rect -2458 -31 -2449 19
rect -2230 19 -2171 29
rect -2230 -31 -2220 19
rect -2458 -83 -2220 -31
rect -2458 -133 -2449 -83
rect -2508 -143 -2449 -133
rect -2230 -133 -2220 -83
rect -2180 -31 -2171 19
rect -1952 19 -1893 29
rect -1952 -31 -1942 19
rect -2180 -83 -1942 -31
rect -2180 -133 -2171 -83
rect -2230 -143 -2171 -133
rect -1952 -133 -1942 -83
rect -1902 -31 -1893 19
rect -1674 19 -1615 29
rect -1674 -31 -1664 19
rect -1902 -83 -1664 -31
rect -1902 -133 -1893 -83
rect -1952 -143 -1893 -133
rect -1674 -133 -1664 -83
rect -1624 -31 -1615 19
rect -1142 -31 -1066 347
rect -1624 -83 -1066 -31
rect -1624 -133 -1615 -83
rect -1674 -143 -1615 -133
rect -2420 -185 -2348 -175
rect -2420 -196 -2410 -185
rect -2749 -228 -2410 -196
rect -2358 -196 -2348 -185
rect -2142 -185 -2070 -175
rect -2142 -196 -2132 -185
rect -2358 -228 -2132 -196
rect -2080 -196 -2070 -185
rect -1864 -185 -1792 -175
rect -1864 -196 -1854 -185
rect -2080 -228 -1854 -196
rect -1802 -196 -1792 -185
rect -1586 -185 -1514 -175
rect -1586 -196 -1576 -185
rect -1802 -228 -1576 -196
rect -1524 -228 -1514 -185
rect -2749 -238 -1514 -228
rect -2885 -319 -2707 -238
rect -4492 -444 -4357 -363
rect -2508 -473 -2449 -463
rect -2508 -523 -2498 -473
rect -2749 -575 -2498 -523
rect -2749 -624 -2697 -575
rect -2885 -705 -2697 -624
rect -2508 -625 -2498 -575
rect -2458 -523 -2449 -473
rect -2230 -473 -2171 -463
rect -2230 -523 -2220 -473
rect -2458 -575 -2220 -523
rect -2458 -625 -2449 -575
rect -2508 -635 -2449 -625
rect -2230 -625 -2220 -575
rect -2180 -523 -2171 -473
rect -1952 -473 -1893 -463
rect -1952 -523 -1942 -473
rect -2180 -575 -1942 -523
rect -2180 -625 -2171 -575
rect -2230 -635 -2171 -625
rect -1952 -625 -1942 -575
rect -1902 -523 -1893 -473
rect -1674 -473 -1615 -463
rect -1674 -523 -1664 -473
rect -1902 -575 -1664 -523
rect -1902 -625 -1893 -575
rect -1952 -635 -1893 -625
rect -1674 -625 -1664 -575
rect -1624 -523 -1615 -473
rect -1142 -523 -1066 -83
rect -878 -65 -838 719
rect -794 718 -574 758
rect -794 24 -754 718
rect -702 572 3395 619
rect -702 116 -655 572
rect -601 320 -591 360
rect -551 320 -111 360
rect -71 320 73 360
rect 113 320 553 360
rect 593 320 737 360
rect 777 320 1217 360
rect 1257 320 1401 360
rect 1441 320 1881 360
rect 1921 320 2065 360
rect 2105 320 2545 360
rect 2585 320 2729 360
rect 2769 320 3209 360
rect 3249 320 3259 360
rect -601 271 -549 320
rect -601 261 -145 271
rect -601 218 -507 261
rect -155 218 -145 261
rect -601 215 -145 218
rect -517 169 -145 215
rect 147 261 519 271
rect 147 218 157 261
rect 509 218 519 261
rect -702 69 -466 116
rect -794 -16 -576 24
rect -878 -105 -659 -65
rect -1624 -575 -1066 -523
rect -1624 -625 -1615 -575
rect -1674 -635 -1615 -625
rect -2420 -716 -2348 -709
rect -2142 -716 -2070 -709
rect -1864 -716 -1792 -709
rect -1586 -716 -1514 -709
rect -2633 -719 -1514 -716
rect -2633 -763 -2410 -719
rect -2358 -763 -2132 -719
rect -2080 -763 -1854 -719
rect -1802 -763 -1576 -719
rect -1524 -763 -1514 -719
rect -2633 -766 -1514 -763
rect -2633 -838 -2583 -766
rect -2420 -773 -2348 -766
rect -2142 -773 -2070 -766
rect -1864 -773 -1792 -766
rect -1586 -773 -1514 -766
rect -2885 -919 -2583 -838
rect -2508 -857 -2449 -847
rect -4492 -1044 -4357 -963
rect -2508 -1009 -2498 -857
rect -2458 -907 -2449 -857
rect -2230 -857 -2171 -847
rect -2230 -907 -2220 -857
rect -2458 -959 -2220 -907
rect -2458 -1009 -2449 -959
rect -2508 -1019 -2449 -1009
rect -2230 -1009 -2220 -959
rect -2180 -907 -2171 -857
rect -1952 -857 -1893 -847
rect -1952 -907 -1942 -857
rect -2180 -959 -1942 -907
rect -2180 -1009 -2171 -959
rect -2230 -1019 -2171 -1009
rect -1952 -1009 -1942 -959
rect -1902 -907 -1893 -857
rect -1674 -857 -1615 -847
rect -1674 -907 -1664 -857
rect -1902 -959 -1664 -907
rect -1902 -1009 -1893 -959
rect -1952 -1019 -1893 -1009
rect -1674 -1009 -1664 -959
rect -1624 -907 -1615 -857
rect -1142 -907 -1066 -575
rect -699 -582 -659 -105
rect -616 -377 -576 -16
rect -513 -300 -466 69
rect -528 -310 -436 -300
rect -528 -355 -518 -310
rect -446 -355 -436 -310
rect -528 -365 -436 -355
rect -616 -401 -570 -377
rect -616 -453 -611 -401
rect -616 -463 -570 -453
rect -616 -576 -570 -553
rect -616 -582 -611 -576
rect -699 -622 -611 -582
rect -616 -630 -611 -622
rect -616 -639 -570 -630
rect -390 -820 -294 169
rect 147 70 519 218
rect 147 25 157 70
rect 509 25 519 70
rect 147 15 519 25
rect 811 261 1183 271
rect 811 218 821 261
rect 1173 218 1183 261
rect 811 70 1183 218
rect 811 25 821 70
rect 1173 25 1183 70
rect 811 15 1183 25
rect 1475 261 1847 271
rect 1475 218 1485 261
rect 1837 218 1847 261
rect 1475 70 1847 218
rect 1475 25 1485 70
rect 1837 25 1847 70
rect 1475 15 1847 25
rect 2139 261 2511 271
rect 2139 218 2149 261
rect 2501 218 2511 261
rect 2139 70 2511 218
rect 2139 25 2149 70
rect 2501 25 2511 70
rect 2139 15 2511 25
rect 2803 261 3175 271
rect 2803 218 2813 261
rect 3165 218 3175 261
rect 2803 70 3175 218
rect 2803 25 2813 70
rect 3165 25 3175 70
rect 2803 15 3175 25
rect 59 -21 105 3
rect 59 -73 64 -21
rect 59 -97 105 -73
rect 723 -21 769 3
rect 723 -73 728 -21
rect 723 -97 769 -73
rect 1387 -21 1433 3
rect 1387 -73 1392 -21
rect 1387 -97 1433 -73
rect 2051 -21 2097 3
rect 2051 -73 2056 -21
rect 2051 -97 2097 -73
rect 2715 -21 2761 3
rect 2715 -73 2720 -21
rect 2715 -97 2761 -73
rect 59 -489 99 -97
rect -239 -499 99 -489
rect -239 -541 -229 -499
rect -171 -531 99 -499
rect -171 -541 -161 -531
rect -239 -551 -161 -541
rect 59 -554 99 -531
rect 147 -119 519 -109
rect 147 -163 157 -119
rect 509 -163 519 -119
rect 147 -302 519 -163
rect 723 -302 763 -97
rect 147 -349 763 -302
rect 147 -489 519 -349
rect 147 -532 157 -489
rect 509 -532 519 -489
rect 147 -542 519 -532
rect 723 -554 763 -349
rect 811 -119 1183 -109
rect 811 -163 821 -119
rect 1173 -163 1183 -119
rect 811 -302 1183 -163
rect 1387 -302 1427 -97
rect 811 -349 1427 -302
rect 811 -489 1183 -349
rect 811 -532 821 -489
rect 1173 -532 1183 -489
rect 811 -542 1183 -532
rect 1387 -554 1427 -349
rect 1475 -119 1847 -109
rect 1475 -163 1485 -119
rect 1837 -163 1847 -119
rect 1475 -302 1847 -163
rect 2051 -302 2091 -97
rect 1475 -305 2091 -302
rect 1475 -346 1863 -305
rect 2023 -346 2091 -305
rect 1475 -349 2091 -346
rect 1475 -489 1847 -349
rect 1475 -532 1485 -489
rect 1837 -532 1847 -489
rect 1475 -542 1847 -532
rect 2051 -554 2091 -349
rect 2139 -119 2511 -109
rect 2139 -163 2149 -119
rect 2501 -163 2511 -119
rect 2139 -302 2511 -163
rect 2715 -302 2755 -97
rect 2139 -349 2755 -302
rect 2139 -489 2511 -349
rect 2139 -532 2149 -489
rect 2501 -532 2511 -489
rect 2139 -542 2511 -532
rect 2715 -554 2755 -349
rect 2803 -119 3175 -109
rect 2803 -163 2813 -119
rect 3165 -163 3175 -119
rect 2803 -302 3175 -163
rect 3345 -302 3395 572
rect 3509 311 3569 900
rect 3509 301 3775 311
rect 3509 82 3642 301
rect 3765 82 3775 301
rect 3509 72 3775 82
rect 2803 -349 3395 -302
rect 2803 -489 3175 -349
rect 2803 -532 2813 -489
rect 3165 -532 3175 -489
rect 2803 -542 3175 -532
rect 59 -578 105 -554
rect 59 -630 64 -578
rect 59 -654 105 -630
rect 723 -578 769 -554
rect 723 -630 728 -578
rect 723 -654 769 -630
rect 1387 -578 1433 -554
rect 1387 -630 1392 -578
rect 1387 -654 1433 -630
rect 2051 -578 2097 -554
rect 2051 -630 2056 -578
rect 2051 -654 2097 -630
rect 2715 -578 2761 -554
rect 2715 -630 2720 -578
rect 2715 -654 2761 -630
rect 147 -675 519 -666
rect 147 -718 157 -675
rect 509 -718 519 -675
rect -1624 -959 -1066 -907
rect -517 -869 -145 -820
rect -517 -912 -507 -869
rect -155 -912 -145 -869
rect -517 -922 -145 -912
rect 147 -869 519 -718
rect 147 -912 157 -869
rect 509 -912 519 -869
rect 147 -922 519 -912
rect 811 -675 1183 -666
rect 811 -718 821 -675
rect 1173 -718 1183 -675
rect 811 -869 1183 -718
rect 811 -912 821 -869
rect 1173 -912 1183 -869
rect 811 -922 1183 -912
rect 1475 -675 1847 -666
rect 1475 -718 1485 -675
rect 1837 -718 1847 -675
rect 1475 -869 1847 -718
rect 1475 -912 1485 -869
rect 1837 -912 1847 -869
rect 1475 -922 1847 -912
rect 2139 -675 2511 -666
rect 2139 -718 2149 -675
rect 2501 -718 2511 -675
rect 2139 -869 2511 -718
rect 2139 -912 2149 -869
rect 2501 -912 2511 -869
rect 2139 -922 2511 -912
rect 2803 -675 3175 -666
rect 2803 -718 2813 -675
rect 3165 -718 3175 -675
rect 2803 -869 3175 -718
rect 2803 -912 2813 -869
rect 3165 -912 3175 -869
rect 2803 -922 3175 -912
rect 4247 -833 4631 -823
rect -1624 -1009 -1615 -959
rect -1674 -1019 -1615 -1009
rect -1142 -971 -1066 -959
rect 4247 -971 4257 -833
rect 4315 -971 4631 -833
rect -1142 -1011 -591 -971
rect -551 -1011 -111 -971
rect -71 -1011 73 -971
rect 113 -1011 553 -971
rect 593 -1011 737 -971
rect 777 -1011 1217 -971
rect 1257 -1011 1401 -971
rect 1441 -1011 1881 -971
rect 1921 -1011 2065 -971
rect 2105 -1011 2545 -971
rect 2585 -1011 2729 -971
rect 2769 -1011 3209 -971
rect 3249 -1011 3259 -971
rect 4247 -981 4631 -971
use lvnmos_4S7S6F  lvnmos_4S7S6F_0
timestamp 1752866318
transform -1 0 -1550 0 -1 -549
box -241 -276 1075 660
use lvnmos_5S7A3R  lvnmos_5S7A3R_0
timestamp 1752864670
transform -1 0 -2106 0 -1 537
box -241 -276 519 276
use lvnmos_5S7JXQ  lvnmos_5S7JXQ_0
timestamp 1752864670
transform -1 0 -2384 0 -1 1131
box -241 -276 241 276
use lvnmos_5S7JXQ  lvnmos_5S7JXQ_1
timestamp 1752864670
transform -1 0 -1962 0 -1 1131
box -241 -276 241 276
use lvnmos_5S7S6P  lvnmos_5S7S6P_0
timestamp 1752864670
transform 1 0 -2384 0 1 -57
box -241 -276 1075 276
use lvnmos_5SCLEP  lvnmos_5SCLEP_0
timestamp 1752865035
transform -1 0 -2384 0 -1 1675
box -241 -226 241 226
use lvnmos_5SUVYP  lvnmos_5SUVYP_0
timestamp 1752865035
transform -1 0 -2378 0 -1 2144
box -247 -201 247 201
use lvnmos_BBXWCS  lvnmos_BBXWCS_0
timestamp 1749294910
transform 0 1 -342 -1 0 -427
box -118 -274 118 274
use lvnmos_BBXWCS  lvnmos_BBXWCS_1
timestamp 1749294910
transform 0 1 -342 -1 0 -603
box -118 -274 118 274
use lvnmos_S23XCS  lvnmos_S23XCS_0
timestamp 1749147318
transform 0 1 333 -1 0 -984
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_1
timestamp 1749147318
transform 0 1 997 -1 0 -604
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_2
timestamp 1749147318
transform 0 1 333 -1 0 -604
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_3
timestamp 1749147318
transform 0 1 1661 -1 0 -604
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_4
timestamp 1749147318
transform 0 1 2325 -1 0 -604
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_5
timestamp 1749147318
transform 0 1 2989 -1 0 -604
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_6
timestamp 1749147318
transform 0 1 2989 -1 0 -984
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_7
timestamp 1749147318
transform 0 1 997 -1 0 -984
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_8
timestamp 1749147318
transform 0 1 1661 -1 0 -984
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_9
timestamp 1749147318
transform 0 1 2325 -1 0 -984
box -220 -362 220 362
use lvnmos_S23XCS  lvnmos_S23XCS_12
timestamp 1749147318
transform 0 1 -331 -1 0 -984
box -220 -362 220 362
use lvpmos_S23XCS  lvpmos_S23XCS_0
timestamp 1749294910
transform 0 1 1661 -1 0 -47
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_1
timestamp 1749294910
transform 0 1 2989 -1 0 333
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_2
timestamp 1749294910
transform 0 1 333 -1 0 333
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_3
timestamp 1749294910
transform 0 1 997 -1 0 333
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_4
timestamp 1749294910
transform 0 1 1661 -1 0 333
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_5
timestamp 1749294910
transform 0 1 2325 -1 0 333
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_6
timestamp 1749294910
transform 0 1 333 -1 0 -47
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_7
timestamp 1749294910
transform 0 1 997 -1 0 -47
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_8
timestamp 1749294910
transform 0 1 2325 -1 0 -47
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_9
timestamp 1749294910
transform 0 1 2989 -1 0 -47
box -268 -410 268 410
use lvpmos_S23XCS  lvpmos_S23XCS_10
timestamp 1749294910
transform 0 1 -331 -1 0 333
box -268 -410 268 410
use sg13g2_dfrbp_2  sg13g2_dfrbp_2_0
timestamp 1752936403
transform 1 0 1546 0 1 1598
box -48 -56 2928 834
use sg13g2_dfrbp_2  sg13g2_dfrbp_2_1
timestamp 1752936403
transform -1 0 2698 0 -1 1598
box -48 -56 2928 834
use sg13g2_dfrbp_2  sg13g2_dfrbp_2_2
timestamp 1752936403
transform 1 0 -1334 0 1 1598
box -48 -56 2928 834
use sg13g2_inv_4  sg13g2_inv_4_0
timestamp 1752936403
transform -1 0 4224 0 -1 540
box -48 -56 624 834
use sg13g2_inv_4  sg13g2_inv_4_1
timestamp 1752936403
transform -1 0 -758 0 -1 1598
box -48 -56 624 834
use sg13g2_inv_4  sg13g2_inv_4_2
timestamp 1752936403
transform 1 0 3648 0 1 -1158
box -48 -56 624 834
use sg13g2_inv_4  sg13g2_inv_4_3
timestamp 1752936403
transform -1 0 4234 0 -1 1598
box -48 -56 624 834
use sg13g2_or2_2  sg13g2_or2_2_0
timestamp 1752937939
transform -1 0 -182 0 -1 1598
box -48 -56 624 834
use trimsw  trimsw_0
timestamp 1757363851
transform 1 0 5032 0 1 -426
box -9524 -779 -7781 38
use trimsw  trimsw_1
timestamp 1757363851
transform 1 0 5032 0 1 174
box -9524 -779 -7781 38
use trimsw  trimsw_2
timestamp 1757363851
transform 1 0 5032 0 1 774
box -9524 -779 -7781 38
use trimsw  trimsw_3
timestamp 1757363851
transform 1 0 5032 0 1 1374
box -9524 -779 -7781 38
use trimsw  trimsw_4
timestamp 1757363851
transform 1 0 5032 0 1 1974
box -9524 -779 -7781 38
use trimsw  trimsw_5
timestamp 1757363851
transform 1 0 5032 0 1 2574
box -9524 -779 -7781 38
<< labels >>
flabel metal2 4387 -981 4631 -823 0 FreeSans 800 0 0 0 OSC
port 2 nsew
flabel metal2 4391 1208 4631 1347 0 FreeSans 400 0 0 0 RESET
port 4 nsew
flabel metal1 4391 -1414 4631 -1084 0 FreeSans 400 0 0 0 VSS
port 9 nsew
flabel metal2 3670 1439 3670 1439 0 FreeSans 320 0 0 0 RESETB
flabel metal1 -726 1259 -726 1259 0 FreeSans 160 0 0 0 ENA2
flabel metal2 -860 436 -860 436 0 FreeSans 160 0 0 0 ENA1
flabel metal2 -1839 2453 -1632 2593 0 FreeSans 800 0 0 0 EN
port 0 nsew
flabel metal1 4434 1993 4631 2391 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal2 -2227 2432 -2030 2593 0 FreeSans 800 0 0 0 IB
port 7 nsew
flabel metal1 3847 1893 3847 1893 0 FreeSans 160 0 0 0 ENA_D1
flabel metal2 -4492 1956 -4357 2037 0 FreeSans 320 0 0 0 T0
port 10 nsew
flabel metal2 -4492 1356 -4357 1437 0 FreeSans 320 0 0 0 T1
port 11 nsew
flabel metal2 -4492 756 -4357 837 0 FreeSans 320 0 0 0 T2
port 12 nsew
flabel metal2 -4492 156 -4357 237 0 FreeSans 320 0 0 0 T3
port 13 nsew
flabel metal2 -4492 -444 -4357 -363 0 FreeSans 320 0 0 0 T4
port 14 nsew
flabel metal2 -4492 -1044 -4357 -963 0 FreeSans 320 0 0 0 T5
port 15 nsew
<< end >>
