magic
tech ihp-sg13g2
timestamp 1748598742
<< dnwell >>
rect -174 -174 174 174
<< nbase >>
rect -193 -193 193 193
<< pdiff >>
rect -100 93 100 100
rect -100 -93 -93 93
rect 93 -93 100 93
rect -100 -100 100 -93
<< pdiffc >>
rect -93 -93 93 93
<< psubdiff >>
rect -254 247 254 254
rect -254 231 -217 247
rect 217 231 254 247
rect -254 224 254 231
rect -254 217 -224 224
rect -254 -217 -247 217
rect -231 -217 -224 217
rect 224 217 254 224
rect -254 -224 -224 -217
rect 224 -217 231 217
rect 247 -217 254 217
rect 224 -224 254 -217
rect -254 -231 254 -224
rect -254 -247 -217 -231
rect 217 -247 254 -231
rect -254 -254 254 -247
<< nsubdiff >>
rect -169 162 169 169
rect -169 146 -132 162
rect 132 146 169 162
rect -169 139 169 146
rect -169 132 -139 139
rect -169 -132 -162 132
rect -146 -132 -139 132
rect 139 132 169 139
rect -169 -139 -139 -132
rect 139 -132 146 132
rect 162 -132 169 132
rect 139 -139 169 -132
rect -169 -146 169 -139
rect -169 -162 -132 -146
rect 132 -162 169 -146
rect -169 -169 169 -162
<< psubdiffcont >>
rect -217 231 217 247
rect -247 -217 -231 217
rect 231 -217 247 217
rect -217 -247 217 -231
<< nsubdiffcont >>
rect -132 146 132 162
rect -162 -132 -146 132
rect 146 -132 162 132
rect -132 -162 132 -146
<< metal1 >>
rect -252 247 252 252
rect -252 231 -217 247
rect 217 231 252 247
rect -252 226 252 231
rect -252 217 -226 226
rect -252 -217 -247 217
rect -231 -217 -226 217
rect 226 217 252 226
rect -167 162 167 167
rect -167 146 -132 162
rect 132 146 167 162
rect -167 141 167 146
rect -167 132 -141 141
rect -167 -132 -162 132
rect -146 -132 -141 132
rect 141 132 167 141
rect -98 93 98 98
rect -98 -93 -93 93
rect 93 -93 98 93
rect -98 -98 98 -93
rect -167 -141 -141 -132
rect 141 -132 146 132
rect 162 -132 167 132
rect 141 -141 167 -132
rect -167 -146 167 -141
rect -167 -162 -132 -146
rect 132 -162 167 -146
rect -167 -167 167 -162
rect -252 -226 -226 -217
rect 226 -217 231 217
rect 247 -217 252 217
rect 226 -226 252 -217
rect -252 -231 252 -226
rect -252 -247 -217 -231
rect 217 -247 252 -231
rect -252 -252 252 -247
<< properties >>
string gencell pnpmpa
string library sg13g2_devstdin
string parameters w 2 l 2 nx 1 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class bjt glc 0 grc 0 gtc 0 gbc 0
<< end >>
