magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 17 56 741 292
rect -26 -56 794 56
<< nmos >>
rect 111 118 137 266
rect 213 118 239 266
rect 315 118 341 266
rect 417 118 443 266
rect 621 118 647 266
<< pmos >>
rect 111 412 137 636
rect 213 412 239 636
rect 315 412 341 636
rect 417 412 443 636
rect 519 412 545 580
rect 621 412 647 580
<< ndiff >>
rect 43 232 111 266
rect 43 200 57 232
rect 89 200 111 232
rect 43 164 111 200
rect 43 132 57 164
rect 89 132 111 164
rect 43 118 111 132
rect 137 232 213 266
rect 137 200 159 232
rect 191 200 213 232
rect 137 164 213 200
rect 137 132 159 164
rect 191 132 213 164
rect 137 118 213 132
rect 239 164 315 266
rect 239 132 261 164
rect 293 132 315 164
rect 239 118 315 132
rect 341 232 417 266
rect 341 200 363 232
rect 395 200 417 232
rect 341 164 417 200
rect 341 132 363 164
rect 395 132 417 164
rect 341 118 417 132
rect 443 164 621 266
rect 443 132 485 164
rect 517 132 553 164
rect 585 132 621 164
rect 443 118 621 132
rect 647 232 715 266
rect 647 200 669 232
rect 701 200 715 232
rect 647 164 715 200
rect 647 132 669 164
rect 701 132 715 164
rect 647 118 715 132
<< pdiff >>
rect 43 622 111 636
rect 43 590 57 622
rect 89 590 111 622
rect 43 540 111 590
rect 43 508 57 540
rect 89 508 111 540
rect 43 458 111 508
rect 43 426 57 458
rect 89 426 111 458
rect 43 412 111 426
rect 137 622 213 636
rect 137 590 159 622
rect 191 590 213 622
rect 137 540 213 590
rect 137 508 159 540
rect 191 508 213 540
rect 137 458 213 508
rect 137 426 159 458
rect 191 426 213 458
rect 137 412 213 426
rect 239 622 315 636
rect 239 590 261 622
rect 293 590 315 622
rect 239 540 315 590
rect 239 508 261 540
rect 293 508 315 540
rect 239 412 315 508
rect 341 622 417 636
rect 341 590 363 622
rect 395 590 417 622
rect 341 540 417 590
rect 341 508 363 540
rect 395 508 417 540
rect 341 458 417 508
rect 341 426 363 458
rect 395 426 417 458
rect 341 412 417 426
rect 443 580 505 636
rect 443 540 519 580
rect 443 508 465 540
rect 497 508 519 540
rect 443 458 519 508
rect 443 426 465 458
rect 497 426 519 458
rect 443 412 519 426
rect 545 540 621 580
rect 545 508 567 540
rect 599 508 621 540
rect 545 472 621 508
rect 545 440 567 472
rect 599 440 621 472
rect 545 412 621 440
rect 647 566 715 580
rect 647 534 669 566
rect 701 534 715 566
rect 647 412 715 534
<< ndiffc >>
rect 57 200 89 232
rect 57 132 89 164
rect 159 200 191 232
rect 159 132 191 164
rect 261 132 293 164
rect 363 200 395 232
rect 363 132 395 164
rect 485 132 517 164
rect 553 132 585 164
rect 669 200 701 232
rect 669 132 701 164
<< pdiffc >>
rect 57 590 89 622
rect 57 508 89 540
rect 57 426 89 458
rect 159 590 191 622
rect 159 508 191 540
rect 159 426 191 458
rect 261 590 293 622
rect 261 508 293 540
rect 363 590 395 622
rect 363 508 395 540
rect 363 426 395 458
rect 465 508 497 540
rect 465 426 497 458
rect 567 508 599 540
rect 567 440 599 472
rect 669 534 701 566
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 111 636 137 672
rect 213 636 239 672
rect 315 636 341 672
rect 417 636 443 672
rect 519 580 545 616
rect 621 580 647 616
rect 111 334 137 412
rect 213 334 239 412
rect 315 364 341 412
rect 417 364 443 412
rect 519 380 545 412
rect 621 380 647 412
rect 315 350 460 364
rect 519 363 647 380
rect 519 350 581 363
rect 315 334 346 350
rect 111 318 346 334
rect 378 318 414 350
rect 446 318 460 350
rect 111 304 460 318
rect 564 331 581 350
rect 613 331 647 363
rect 564 314 647 331
rect 111 266 137 304
rect 213 266 239 304
rect 315 266 341 304
rect 417 266 443 304
rect 621 266 647 314
rect 111 82 137 118
rect 213 82 239 118
rect 315 82 341 118
rect 417 82 443 118
rect 621 82 647 118
<< polycont >>
rect 346 318 378 350
rect 414 318 446 350
rect 581 331 613 363
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 47 622 99 712
rect 47 590 57 622
rect 89 590 99 622
rect 47 540 99 590
rect 47 508 57 540
rect 89 508 99 540
rect 47 458 99 508
rect 47 426 57 458
rect 89 426 99 458
rect 47 423 99 426
rect 149 622 201 626
rect 149 590 159 622
rect 191 590 201 622
rect 149 540 201 590
rect 149 508 159 540
rect 191 508 201 540
rect 149 458 201 508
rect 251 622 303 712
rect 251 590 261 622
rect 293 590 303 622
rect 251 540 303 590
rect 251 508 261 540
rect 293 508 303 540
rect 251 498 303 508
rect 353 622 405 626
rect 353 590 363 622
rect 395 590 405 622
rect 353 540 405 590
rect 353 508 363 540
rect 395 508 405 540
rect 149 426 159 458
rect 191 433 201 458
rect 353 458 405 508
rect 353 433 363 458
rect 191 426 363 433
rect 395 426 405 458
rect 149 399 405 426
rect 455 540 507 712
rect 659 566 711 712
rect 455 508 465 540
rect 497 508 507 540
rect 455 458 507 508
rect 455 426 465 458
rect 497 426 507 458
rect 557 540 609 554
rect 557 508 567 540
rect 599 508 609 540
rect 659 534 669 566
rect 701 534 711 566
rect 659 528 711 534
rect 557 484 609 508
rect 557 472 718 484
rect 557 440 567 472
rect 599 440 718 472
rect 557 430 718 440
rect 455 416 507 426
rect 149 368 201 399
rect 64 305 201 368
rect 540 363 630 377
rect 336 350 486 360
rect 336 318 346 350
rect 378 318 414 350
rect 446 318 486 350
rect 336 308 486 318
rect 149 245 201 305
rect 47 232 99 242
rect 47 200 57 232
rect 89 200 99 232
rect 47 164 99 200
rect 47 132 57 164
rect 89 132 99 164
rect 47 44 99 132
rect 149 232 405 245
rect 149 200 159 232
rect 191 213 363 232
rect 191 200 201 213
rect 149 164 201 200
rect 353 200 363 213
rect 395 200 405 232
rect 453 242 486 308
rect 540 331 581 363
rect 613 331 630 363
rect 540 295 630 331
rect 680 242 718 430
rect 453 232 718 242
rect 453 210 669 232
rect 149 132 159 164
rect 191 132 201 164
rect 149 121 201 132
rect 251 164 303 174
rect 251 132 261 164
rect 293 132 303 164
rect 251 44 303 132
rect 353 164 405 200
rect 649 200 669 210
rect 701 200 718 232
rect 353 132 363 164
rect 395 132 405 164
rect 353 129 405 132
rect 475 164 595 174
rect 475 132 485 164
rect 517 132 553 164
rect 585 132 595 164
rect 475 122 595 132
rect 649 164 718 200
rect 649 132 669 164
rect 701 132 718 164
rect 649 128 718 132
rect 509 44 561 122
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 64 305 201 368 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 540 295 630 377 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 128046
string GDS_FILE 6_final.gds
string GDS_START 121798
<< end >>
