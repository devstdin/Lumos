magic
tech ihp-sg13g2
timestamp 1752520737
<< error_p >>
rect -18 2036 -13 2041
rect 13 2036 18 2041
rect 82 2036 87 2041
rect 113 2036 118 2041
rect -23 2031 23 2036
rect 77 2031 123 2036
rect -18 2025 18 2031
rect 82 2025 118 2031
rect -23 2020 23 2025
rect 77 2020 123 2025
rect -18 2015 -13 2020
rect 13 2015 18 2020
rect 82 2015 87 2020
rect 113 2015 118 2020
rect -18 -2020 -13 -2015
rect 13 -2020 18 -2015
rect 82 -2020 87 -2015
rect 113 -2020 118 -2015
rect -23 -2025 23 -2020
rect 77 -2025 123 -2020
rect -18 -2031 18 -2025
rect 82 -2031 118 -2025
rect -23 -2036 23 -2031
rect 77 -2036 123 -2031
rect -18 -2041 -13 -2036
rect 13 -2041 18 -2036
rect 82 -2041 87 -2036
rect 113 -2041 118 -2036
<< psubdiff >>
rect -115 2126 215 2133
rect -115 2110 -78 2126
rect 178 2110 215 2126
rect -115 2103 215 2110
rect -115 2096 -85 2103
rect -115 -2096 -108 2096
rect -92 -2096 -85 2096
rect 185 2096 215 2103
rect -115 -2103 -85 -2096
rect 185 -2096 192 2096
rect 208 -2096 215 2096
rect 185 -2103 215 -2096
rect -115 -2110 215 -2103
rect -115 -2126 -78 -2110
rect 178 -2126 215 -2110
rect -115 -2133 215 -2126
<< psubdiffcont >>
rect -78 2110 178 2126
rect -108 -2096 -92 2096
rect 192 -2096 208 2096
rect -78 -2126 178 -2110
<< poly >>
rect -25 2036 25 2043
rect -25 2020 -18 2036
rect 18 2020 25 2036
rect -25 2000 25 2020
rect -25 -2020 25 -2000
rect -25 -2036 -18 -2020
rect 18 -2036 25 -2020
rect -25 -2043 25 -2036
rect 75 2036 125 2043
rect 75 2020 82 2036
rect 118 2020 125 2036
rect 75 2000 125 2020
rect 75 -2020 125 -2000
rect 75 -2036 82 -2020
rect 118 -2036 125 -2020
rect 75 -2043 125 -2036
<< polycont >>
rect -18 2020 18 2036
rect -18 -2036 18 -2020
rect 82 2020 118 2036
rect 82 -2036 118 -2020
<< xpolyres >>
rect -25 -2000 25 2000
rect 75 -2000 125 2000
<< metal1 >>
rect -113 2126 213 2131
rect -113 2110 -78 2126
rect 178 2110 213 2126
rect -113 2105 213 2110
rect -113 2096 -87 2105
rect -113 -2096 -108 2096
rect -92 -2096 -87 2096
rect 187 2096 213 2105
rect -113 -2105 -87 -2096
rect 187 -2096 192 2096
rect 208 -2096 213 2096
rect 187 -2105 213 -2096
rect -113 -2110 213 -2105
rect -113 -2126 -78 -2110
rect 178 -2126 213 -2110
rect -113 -2131 213 -2126
<< properties >>
string gencell rhigh
string library sg13g2_devstdin
string parameters w 0.5 l 40 nx 2 dx 0.5 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class resistor endcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
