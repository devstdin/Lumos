magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< metal1 >>
rect 1460 21880 23980 21968
rect 60 21124 25380 21212
rect 1460 20368 23980 20456
rect 60 19612 25380 19700
rect 1460 18856 23980 18944
rect 60 18100 25380 18188
rect 1460 17344 23980 17432
rect 60 16588 25380 16676
rect 1460 15832 23980 15920
rect 60 15076 25380 15164
rect 1460 14320 23980 14408
rect 60 13564 25380 13652
rect 1460 12808 23980 12896
rect 60 12052 25380 12140
rect 1460 11296 23980 11384
rect 60 10540 25380 10628
rect 1460 9784 23980 9872
rect 60 9028 25380 9116
rect 1460 8272 23980 8360
rect 60 7516 25380 7604
rect 1460 6760 23980 6848
rect 60 6004 25380 6092
rect 1460 5248 23980 5336
rect 60 4492 25380 4580
rect 1460 3736 23980 3824
<< metal2 >>
rect 5146 17356 5186 17684
rect 5272 17300 5312 24212
rect 5104 17260 5312 17300
rect 4852 17068 4892 17204
rect 4768 15572 4808 17059
rect 4768 15532 4892 15572
rect 4516 15342 4556 15456
rect 4684 14668 4724 14900
rect 4852 14380 4892 14708
rect 5104 14516 5144 17260
rect 5242 17020 5312 17060
rect 5272 16052 5312 17020
rect 5356 16244 5396 21716
rect 5524 17740 5564 18356
rect 5440 17145 5480 17684
rect 5776 17108 5816 18740
rect 6112 18700 6236 18740
rect 6196 18657 6236 18700
rect 6280 18556 6320 18740
rect 6028 18414 6068 18528
rect 6364 17876 6404 24404
rect 6448 18452 6488 24884
rect 6586 20716 6656 20756
rect 6448 18412 6572 18452
rect 6364 17836 6488 17876
rect 5524 17068 5816 17108
rect 5944 16876 5984 17300
rect 6280 16878 6320 16992
rect 5356 16204 5564 16244
rect 5272 16012 5396 16052
rect 5272 14574 5312 14688
rect 5104 14476 5312 14516
rect 4404 13652 4444 14043
rect 4404 13612 4472 13652
rect 4432 13036 4472 13612
rect 4516 11980 4556 13844
rect 4600 13230 4640 13344
rect 4684 13132 4724 13953
rect 5104 13902 5168 14036
rect 4768 13132 4808 13268
rect 5104 12596 5144 13902
rect 5188 13204 5228 13364
rect 5032 12556 5144 12596
rect 5032 12212 5072 12556
rect 5032 12172 5090 12212
rect 5050 12116 5090 12172
rect 5050 12076 5144 12116
rect 4852 11406 4892 11520
rect 4768 10156 4808 10868
rect 4390 9966 4430 10080
rect 5104 9044 5144 12076
rect 5272 11692 5312 14476
rect 5356 13996 5396 16012
rect 5776 15342 5816 16244
rect 5896 16204 5936 16340
rect 6196 16204 6236 16340
rect 6364 16204 6404 17684
rect 6448 17108 6488 17836
rect 6532 17164 6572 18412
rect 6616 18356 6656 20716
rect 6784 20180 6824 20660
rect 6868 20524 6908 20756
rect 6700 20140 6824 20180
rect 6700 18796 6740 20140
rect 6868 19852 6908 20084
rect 6952 19564 6992 24596
rect 7288 20524 7328 20660
rect 7036 19604 7076 19988
rect 7162 19950 7202 20064
rect 7288 20044 7328 20180
rect 7036 19564 7160 19604
rect 7120 19412 7160 19564
rect 6994 19372 7160 19412
rect 7372 19316 7412 25268
rect 7456 20526 7496 20640
rect 7540 20044 7790 20084
rect 7540 19948 7580 20044
rect 7876 19988 7916 20756
rect 7624 19948 7916 19988
rect 8044 19988 8084 21524
rect 8447 21140 8487 21521
rect 8447 21100 8504 21140
rect 8464 20524 8504 21100
rect 8128 20044 8168 20276
rect 8212 19988 8252 20180
rect 8044 19948 8252 19988
rect 7624 19468 7664 19948
rect 6784 18700 6824 19316
rect 7204 19276 7412 19316
rect 7288 19180 8084 19220
rect 6700 18508 6908 18548
rect 6700 18412 6740 18508
rect 6616 18316 6740 18356
rect 6448 17068 6572 17108
rect 6280 16052 6320 16119
rect 6280 16012 6404 16052
rect 6364 15724 6404 16012
rect 6448 15572 6488 16916
rect 6532 16244 6572 17068
rect 6700 16876 6740 18316
rect 6784 16686 6824 16800
rect 6616 16300 6824 16340
rect 6532 16204 6656 16244
rect 6784 16204 6824 16300
rect 6112 15532 6404 15572
rect 6448 15532 6512 15572
rect 5944 15244 6152 15284
rect 6112 14668 6152 15244
rect 5776 14228 5816 14420
rect 6364 14228 6404 15532
rect 6616 15476 6656 16204
rect 6700 15633 6740 15764
rect 5524 14092 5564 14227
rect 5776 14188 5900 14228
rect 6196 14188 6404 14228
rect 6448 15436 6656 15476
rect 5440 12556 5480 14036
rect 5776 12652 5816 13268
rect 6028 13038 6068 13152
rect 6196 12980 6236 14188
rect 6280 13420 6320 14036
rect 6196 12940 6404 12980
rect 5356 12460 5480 12500
rect 5440 10772 5480 12460
rect 5734 11790 5774 11904
rect 5524 10828 5564 11732
rect 5860 11540 5900 12692
rect 5944 12417 5984 12596
rect 6364 12460 6404 12940
rect 6448 12404 6488 15436
rect 6784 14956 6824 15572
rect 7120 14996 7160 18836
rect 7288 18548 7328 19180
rect 7372 19084 7580 19124
rect 7204 18508 7328 18548
rect 7204 16974 7244 18508
rect 7540 18452 7580 19084
rect 8128 18556 8168 19948
rect 8548 19700 8588 25172
rect 9052 21620 9092 23444
rect 9556 21676 9596 25446
rect 9976 23060 10016 25446
rect 10396 23060 10436 25446
rect 10816 24172 10856 25446
rect 11236 23060 11276 25446
rect 9976 23020 10100 23060
rect 10396 23020 10520 23060
rect 11236 23020 11444 23060
rect 9010 21580 9092 21620
rect 8632 21294 8672 21408
rect 8716 20140 8756 20756
rect 8447 19660 8588 19700
rect 8447 19299 8487 19660
rect 8632 19278 8672 19392
rect 7540 18412 8168 18452
rect 7624 17644 7664 17779
rect 8044 17356 8084 17724
rect 8128 17723 8168 18412
rect 8548 17876 8588 18740
rect 8528 17836 8588 17876
rect 8528 17741 8568 17836
rect 8632 17740 8672 18932
rect 8716 17204 8756 19892
rect 8800 19180 8840 21524
rect 9010 21484 9050 21580
rect 9304 21390 9344 21504
rect 8968 20044 9008 20180
rect 8884 18508 8924 19796
rect 9178 19243 9218 19378
rect 9094 19124 9134 19143
rect 8968 19084 9134 19124
rect 8968 17644 9008 19084
rect 9220 17780 9260 19028
rect 9304 17836 9344 18356
rect 9094 17740 9260 17780
rect 9136 17644 9260 17684
rect 8632 17164 8756 17204
rect 7456 17068 7832 17108
rect 7204 15916 7244 16820
rect 7456 15532 7496 15668
rect 7204 15244 7580 15284
rect 7120 14956 7328 14996
rect 6574 13997 6614 14132
rect 7120 14092 7160 14956
rect 7540 14668 7580 15244
rect 6112 12364 6488 12404
rect 6532 12384 6572 12498
rect 6616 12308 6656 13460
rect 6532 12268 6656 12308
rect 6112 11884 6152 12116
rect 6532 12020 6572 12268
rect 6532 11980 6656 12020
rect 5944 11743 5984 11878
rect 6280 11596 6572 11636
rect 5776 11500 5900 11540
rect 5776 11252 5816 11500
rect 5776 11212 6152 11252
rect 6112 11020 6152 11212
rect 5836 10868 5876 11012
rect 6028 10868 6068 10992
rect 5836 10828 6068 10868
rect 5440 10732 5564 10772
rect 5075 9004 5144 9044
rect 5188 9484 5264 9524
rect 5440 9486 5480 9600
rect 5524 9484 5564 10732
rect 5608 10156 5732 10196
rect 4936 8852 4976 8976
rect 4684 8812 4976 8852
rect 4684 8756 4724 8812
rect 4403 8716 4724 8756
rect 4403 8647 4443 8716
rect 4516 8620 4640 8660
rect 4768 8640 4808 8754
rect 3928 7084 3968 8468
rect 4516 8428 4556 8620
rect 4600 8524 4724 8564
rect 4600 8428 4640 8524
rect 4978 8276 5018 8754
rect 5075 8637 5115 9004
rect 5188 8524 5228 9484
rect 4978 8236 5144 8276
rect 4012 6988 4052 7988
rect 4474 7854 4514 7968
rect 4222 7124 4262 7153
rect 4096 6604 4136 7124
rect 4222 7084 4514 7124
rect 4852 7086 4892 7988
rect 4474 6892 4514 7084
rect 5104 6836 5144 8236
rect 5083 6796 5144 6836
rect 4012 6340 4052 6475
rect 4959 6412 4999 6547
rect 5083 6460 5123 6796
rect 5272 6452 5312 8852
rect 5356 8640 5396 8754
rect 5554 8668 5594 8948
rect 5440 8524 5480 8660
rect 5692 7084 5732 10156
rect 5776 9676 5816 10100
rect 6028 9964 6068 10828
rect 6196 10004 6236 11137
rect 6532 11116 6572 11596
rect 6616 10924 6656 11980
rect 6700 11828 6740 14036
rect 7036 13996 7286 14036
rect 7624 13844 7664 15764
rect 7708 15673 7748 17012
rect 7792 16052 7832 17068
rect 7876 16108 7916 17036
rect 8044 16110 8084 16224
rect 7792 16012 8168 16052
rect 7708 15633 7790 15673
rect 7750 15555 7790 15633
rect 7876 14708 7916 15956
rect 8128 15340 8168 16012
rect 8338 15532 8378 15860
rect 8422 15532 8462 15668
rect 7876 14668 8000 14708
rect 7204 13804 7664 13844
rect 7204 12980 7244 13804
rect 6784 11924 6824 12980
rect 7120 12940 7244 12980
rect 7120 12748 7160 12940
rect 6952 12268 6992 12596
rect 7078 12461 7118 12596
rect 7456 12364 7496 13172
rect 6784 11884 6992 11924
rect 6700 11788 6908 11828
rect 6700 11598 6740 11712
rect 6196 9964 6404 10004
rect 5944 9582 5984 9696
rect 6364 9620 6404 9964
rect 6112 9580 6404 9620
rect 6784 9580 6824 10004
rect 6112 9481 6152 9580
rect 6248 9389 6288 9524
rect 6448 9294 6488 9408
rect 6700 9292 6740 9476
rect 6868 9004 6908 11788
rect 6952 10868 6992 11884
rect 7066 10924 7106 11059
rect 7372 10988 7412 12308
rect 7540 11502 7580 11616
rect 6952 10828 7076 10868
rect 6952 10060 6992 10196
rect 7036 9580 7076 10828
rect 7204 10252 7328 10292
rect 5776 8814 5816 8928
rect 6952 8908 6992 9476
rect 7204 9390 7244 10252
rect 7372 9964 7412 10196
rect 7456 10060 7496 11108
rect 7372 9388 7412 9523
rect 7540 9484 7580 9620
rect 5776 8468 5816 8592
rect 6028 8526 6068 8640
rect 6700 8620 6740 8852
rect 5776 8428 5900 8468
rect 6224 8430 6264 8544
rect 5776 7028 5816 8428
rect 6868 7508 6908 8660
rect 7036 8620 7076 8756
rect 7204 8526 7244 8640
rect 6952 7948 7076 7988
rect 6868 7468 6992 7508
rect 5608 6988 5816 7028
rect 5188 6412 5312 6452
rect 5524 6356 5564 6487
rect 5608 6412 5648 6988
rect 5692 6556 5732 6932
rect 5776 6473 5816 6644
rect 6952 6604 6992 7468
rect 7036 6548 7076 7948
rect 7204 7854 7244 7968
rect 7372 7220 7412 8852
rect 7540 8660 7580 9332
rect 7456 8620 7580 8660
rect 7456 7316 7496 8620
rect 7624 7988 7664 12500
rect 7708 11884 7748 14036
rect 7876 13204 7916 14668
rect 8128 12366 8168 12480
rect 7960 11596 8000 12308
rect 8044 10995 8084 12020
rect 8243 10995 8283 11130
rect 8380 10868 8420 14612
rect 8464 13132 8504 14036
rect 8548 12980 8588 13364
rect 8506 12940 8588 12980
rect 8632 12980 8672 17164
rect 8716 14708 8756 17060
rect 9136 15572 9176 17644
rect 9220 16206 9260 17300
rect 9388 16724 9428 19412
rect 9472 18932 9512 21620
rect 9685 21580 9725 21716
rect 9934 21140 9974 21572
rect 9556 21100 9974 21140
rect 9556 19468 9596 21100
rect 9724 20524 9932 20564
rect 9724 18988 9764 20524
rect 9892 19283 9932 20084
rect 10060 19283 10100 23020
rect 10312 20140 10352 21620
rect 10144 19852 10268 19892
rect 9868 19243 9932 19283
rect 9976 19243 10100 19283
rect 9868 19228 9908 19243
rect 9472 18892 9722 18932
rect 9682 18700 9722 18892
rect 9976 18644 10016 19243
rect 10144 19180 10184 19700
rect 10060 18700 10100 19143
rect 10228 18892 10268 19852
rect 9808 18604 10016 18644
rect 9472 17260 9512 18497
rect 9808 17876 9848 18604
rect 9946 18508 10016 18548
rect 9724 17836 9848 17876
rect 9976 17836 10016 18508
rect 10144 17932 10184 18692
rect 10228 17972 10268 18557
rect 10228 17932 10352 17972
rect 10396 17876 10436 22964
rect 10144 17836 10436 17876
rect 9622 17548 9662 17749
rect 9388 16684 9596 16724
rect 9556 16628 9596 16684
rect 9556 16588 9616 16628
rect 9100 15532 9176 15572
rect 9388 15532 9428 16532
rect 9472 15764 9512 16244
rect 9576 16219 9616 16588
rect 9472 15724 9680 15764
rect 9472 15534 9512 15648
rect 8800 15340 9008 15380
rect 8716 14668 8840 14708
rect 8716 13172 8756 13212
rect 8716 13132 8840 13172
rect 8632 12940 8756 12980
rect 8506 12516 8546 12940
rect 8616 12172 8656 12509
rect 8716 12116 8756 12940
rect 8632 12076 8756 12116
rect 8212 10828 8420 10868
rect 7792 10196 7832 10772
rect 7750 10156 7832 10196
rect 7750 10108 7790 10156
rect 8128 10062 8168 10176
rect 8128 9580 8168 9908
rect 7792 9292 7832 9476
rect 8086 9428 8126 9476
rect 7876 9388 8126 9428
rect 7876 8544 7916 9388
rect 8296 9140 8336 9524
rect 8128 9100 8336 9140
rect 8128 8756 8168 9100
rect 8086 8716 8168 8756
rect 8086 8668 8126 8716
rect 8212 8668 8252 8948
rect 7624 7948 7685 7988
rect 7456 7276 7664 7316
rect 7540 7228 7580 7276
rect 7372 7180 7497 7220
rect 7457 6796 7497 7180
rect 5751 6412 5816 6473
rect 6983 6508 7076 6548
rect 6983 6412 7023 6508
rect 7204 6460 7244 6644
rect 7456 6412 7496 6644
rect 5356 6316 5564 6356
rect 7204 6222 7244 6336
rect 7624 6260 7664 7276
rect 7792 7084 7958 7124
rect 8212 6460 8252 8564
rect 8380 8084 8420 8756
rect 8464 8620 8504 11732
rect 8632 11692 8672 12076
rect 8716 10964 8756 11732
rect 8800 11596 8840 13132
rect 8884 11540 8924 14708
rect 8968 13228 9008 15340
rect 9136 13132 9176 15532
rect 9640 14036 9680 15724
rect 9724 15572 9764 17836
rect 9808 17740 10058 17780
rect 10018 17705 10058 17740
rect 9808 16204 9848 17300
rect 9892 16436 9932 17012
rect 9892 16396 10100 16436
rect 9976 16204 10016 16340
rect 10060 16252 10100 16396
rect 9808 15628 9974 15668
rect 9724 15532 9848 15572
rect 9640 13996 9764 14036
rect 9808 12980 9848 15532
rect 9976 14862 10016 14976
rect 9724 12940 9848 12980
rect 9010 12461 9050 12596
rect 9579 12500 9619 12692
rect 9136 12460 9260 12500
rect 9220 11732 9260 12460
rect 9556 12460 9619 12500
rect 8548 10924 8756 10964
rect 8800 11500 8924 11540
rect 8548 10772 8588 10924
rect 8800 10868 8840 11500
rect 8632 10828 8840 10868
rect 8548 10732 8672 10772
rect 8632 9484 8672 10732
rect 8884 9868 8924 11060
rect 8968 10156 9008 11636
rect 9082 11598 9122 11712
rect 9220 11692 9428 11732
rect 9388 11596 9428 11692
rect 9472 11540 9512 11636
rect 9304 11500 9512 11540
rect 9178 11020 9218 11156
rect 9304 11020 9344 11500
rect 9556 11116 9596 12460
rect 9724 11444 9764 12940
rect 9892 12556 9932 13076
rect 9934 11540 9974 11636
rect 9808 11500 9974 11540
rect 9724 11404 10016 11444
rect 9556 10972 9806 11012
rect 9556 10828 9596 10972
rect 9136 9524 9176 10196
rect 9556 9676 9596 10676
rect 8380 8044 8457 8084
rect 8296 7796 8336 7988
rect 8417 7852 8457 8044
rect 8296 7756 8420 7796
rect 8296 7085 8336 7220
rect 8380 6556 8420 7756
rect 8548 7180 8588 9476
rect 8464 6473 8504 6836
rect 7708 6318 7748 6432
rect 8439 6412 8504 6473
rect 8632 6356 8672 9044
rect 8800 8814 8840 8928
rect 8744 8660 8784 8671
rect 8968 8660 9008 9524
rect 9094 9484 9176 9524
rect 9094 9340 9134 9484
rect 9808 9390 9848 9504
rect 8744 8620 9008 8660
rect 9304 8620 9344 8852
rect 9556 8756 9596 8852
rect 9892 8812 9932 10292
rect 9556 8716 9932 8756
rect 9556 8620 9615 8660
rect 8884 7892 8924 7988
rect 8716 7852 8924 7892
rect 8968 7796 9008 8620
rect 8884 7756 9008 7796
rect 8884 6460 8924 7756
rect 9052 6556 9092 7220
rect 9136 7084 9176 7988
rect 9304 7084 9344 7988
rect 9556 6836 9596 8620
rect 9808 8564 9848 8612
rect 9724 8524 9848 8564
rect 9892 8428 9932 8716
rect 9976 8660 10016 11404
rect 10060 10636 10100 16052
rect 10144 14708 10184 17836
rect 10354 17646 10394 17760
rect 10228 16588 10268 16820
rect 10396 16396 10436 17588
rect 10480 17068 10520 23020
rect 11236 21484 11276 21620
rect 10564 20814 10604 20928
rect 11110 20764 11150 21044
rect 10816 20622 10856 20736
rect 10648 20044 10772 20084
rect 10564 19758 10604 19872
rect 10648 19508 10688 20044
rect 10564 19468 10688 19508
rect 10900 18452 10940 19412
rect 10984 18604 11024 20756
rect 11152 20044 11192 20180
rect 11135 19028 11175 19339
rect 11135 18988 11192 19028
rect 10900 18412 11108 18452
rect 10648 18316 11024 18356
rect 10480 16340 10520 16820
rect 10564 16396 10604 17745
rect 10816 17646 10856 17760
rect 10900 17684 10940 18260
rect 10984 17740 11024 18316
rect 10900 17644 11024 17684
rect 10648 17068 10688 17300
rect 10732 16492 10772 17588
rect 10312 16300 10520 16340
rect 10312 15532 10352 16300
rect 10816 16244 10856 17300
rect 10551 16204 10856 16244
rect 10564 14956 10604 16204
rect 10144 14668 10394 14708
rect 10144 14478 10184 14592
rect 10354 14188 10394 14668
rect 10564 14574 10604 14688
rect 10144 13420 10184 13961
rect 10648 13420 10688 16148
rect 10900 14284 10940 17204
rect 10984 14132 11024 17644
rect 11068 16780 11108 18412
rect 11152 17260 11192 18988
rect 11236 18452 11276 19892
rect 11320 19278 11360 19392
rect 11404 18452 11444 23020
rect 11656 21044 11696 25446
rect 11572 21004 11696 21044
rect 11488 20812 11528 20948
rect 11488 18528 11528 18642
rect 11236 18412 11360 18452
rect 11404 18412 11528 18452
rect 11236 18222 11276 18336
rect 11320 17780 11360 18412
rect 11320 17740 11444 17780
rect 11068 16012 11108 16244
rect 10900 14092 11024 14132
rect 10816 13900 10856 14036
rect 10900 13804 10940 14092
rect 11152 14036 11192 17108
rect 11278 17068 11318 17300
rect 11404 17068 11444 17204
rect 11488 17012 11528 18412
rect 11320 16972 11528 17012
rect 11236 16302 11276 16416
rect 11236 15438 11276 15552
rect 11320 15380 11360 16972
rect 11404 15820 11444 16820
rect 11488 16204 11528 16340
rect 11053 13996 11192 14036
rect 11236 15340 11360 15380
rect 10438 13324 11024 13364
rect 10144 12788 10184 13193
rect 10451 13161 10604 13201
rect 10312 12788 10352 12980
rect 10144 12748 10268 12788
rect 10312 12748 10436 12788
rect 10228 12692 10268 12748
rect 10228 12652 10352 12692
rect 10396 11732 10436 12748
rect 10144 11692 10436 11732
rect 10144 10997 10184 11692
rect 10144 8852 10184 10128
rect 10354 10062 10394 10176
rect 10438 9966 10478 10080
rect 10228 8908 10268 9524
rect 10564 8852 10604 13161
rect 10732 10348 10772 13172
rect 10900 13036 10940 13171
rect 10984 13132 11024 13324
rect 11152 12366 11192 13748
rect 11236 12980 11276 15340
rect 11404 14188 11444 14708
rect 11404 13708 11444 13844
rect 11236 12940 11360 12980
rect 10900 12268 11024 12308
rect 10984 10924 11024 12268
rect 11236 10924 11276 11684
rect 11320 10868 11360 12940
rect 11404 12556 11444 13364
rect 11236 10828 11360 10868
rect 11152 10156 11192 10292
rect 10648 9044 10688 9524
rect 11236 9292 11276 10828
rect 11488 10156 11528 13844
rect 11572 12980 11612 21004
rect 11656 20716 11696 20852
rect 11740 19316 11780 25076
rect 12076 24364 12116 25446
rect 11656 19276 11780 19316
rect 11824 18740 11864 22964
rect 12496 21580 12536 25446
rect 12916 23060 12956 25446
rect 12832 23020 12956 23060
rect 13000 25324 13292 25364
rect 11992 20044 12032 21524
rect 12076 21484 12200 21524
rect 12664 21484 12788 21524
rect 12076 20140 12116 21484
rect 12664 21332 12704 21484
rect 12370 21292 12704 21332
rect 11908 19276 12304 19316
rect 12160 18796 12200 19220
rect 12264 19215 12304 19276
rect 12664 19182 12704 21292
rect 12832 21044 12872 23020
rect 12916 21812 12956 21852
rect 13000 21812 13040 25324
rect 13252 25268 13292 25324
rect 13336 25268 13376 25446
rect 13252 25228 13376 25268
rect 13420 23060 13460 24980
rect 12916 21772 13040 21812
rect 13336 23020 13460 23060
rect 13210 21236 13250 21620
rect 12748 21004 12872 21044
rect 13168 21196 13250 21236
rect 12748 19948 12788 21004
rect 12748 19276 12788 19700
rect 11656 17260 11696 18740
rect 11824 18700 11948 18740
rect 11782 18509 11822 18644
rect 11740 16782 11780 16896
rect 11656 16014 11696 16128
rect 11824 13902 11864 14016
rect 11824 13652 11864 13844
rect 11807 13612 11864 13652
rect 11807 13251 11847 13612
rect 11908 12980 11948 18700
rect 12328 18452 12368 18644
rect 12832 18548 12872 20948
rect 13168 20756 13208 21196
rect 12916 20716 13208 20756
rect 13168 19468 13208 19892
rect 13252 19412 13292 21044
rect 13239 19372 13292 19412
rect 13239 19243 13279 19372
rect 12748 18508 12872 18548
rect 12160 18412 12368 18452
rect 11992 16244 12032 18356
rect 12244 17645 12284 17780
rect 13168 17644 13208 18644
rect 12076 16972 12116 17108
rect 12664 17070 12704 17184
rect 12244 16686 12284 16800
rect 11992 16204 12116 16244
rect 12370 15534 12410 15648
rect 12496 14996 12536 15668
rect 12652 15532 12692 15764
rect 12748 15476 12788 17012
rect 12916 16110 12956 16224
rect 12832 15648 12872 15762
rect 12664 15436 12788 15476
rect 12916 15438 12956 15552
rect 12496 14956 12620 14996
rect 11992 13326 12032 13440
rect 12076 13132 12116 14036
rect 11572 12940 11780 12980
rect 11908 12940 12116 12980
rect 11320 9484 11528 9524
rect 10648 9004 11192 9044
rect 10144 8812 10520 8852
rect 10564 8812 10688 8852
rect 11068 8814 11108 8928
rect 10060 8716 10352 8756
rect 9976 8620 10100 8660
rect 9976 8430 10016 8544
rect 9087 6356 9127 6473
rect 9388 6460 9428 6836
rect 9556 6796 9602 6836
rect 9562 6451 9602 6796
rect 9724 6356 9764 8276
rect 10060 7084 10100 8620
rect 10186 8236 10226 8623
rect 10144 7854 10184 7968
rect 8632 6316 9127 6356
rect 9556 6316 9764 6356
rect 10312 6316 10352 8716
rect 10480 8660 10520 8812
rect 10480 8620 10856 8660
rect 11152 7756 11192 9004
rect 11320 7892 11360 9484
rect 11572 9140 11612 10964
rect 11740 10292 11780 12940
rect 11824 12364 11864 12500
rect 12076 11828 12116 12940
rect 12160 11884 12200 14036
rect 12328 13998 12368 14324
rect 12454 14044 12494 14324
rect 12244 13132 12284 13652
rect 12328 13132 12368 13556
rect 12580 13220 12620 14132
rect 12538 13180 12620 13220
rect 12538 13164 12578 13180
rect 12538 12980 12578 13095
rect 12664 13076 12704 15436
rect 12748 14668 12956 14708
rect 12916 13940 12956 14668
rect 13000 14420 13040 17204
rect 13126 16876 13166 17060
rect 13252 14804 13292 18836
rect 13336 16532 13376 23020
rect 13756 21772 13796 25446
rect 13504 21332 13544 21620
rect 13924 21484 13964 21620
rect 13504 21292 14048 21332
rect 13420 19950 13460 20064
rect 13588 20045 13628 20180
rect 13672 19948 13712 20084
rect 14008 19988 14048 21292
rect 14092 20910 14132 21024
rect 14008 19948 14132 19988
rect 14092 19276 14132 19508
rect 13756 18604 13796 19265
rect 13924 18990 13964 19104
rect 14176 18796 14216 25446
rect 14596 23020 14636 25446
rect 15016 23060 15056 25446
rect 14932 23020 15056 23060
rect 14470 20428 14510 20753
rect 14596 20276 14636 21812
rect 14764 21486 14804 21600
rect 14764 20736 14804 20850
rect 14512 20236 14636 20276
rect 14764 20620 14888 20660
rect 14260 19374 14300 19488
rect 14344 18644 14384 20084
rect 14428 19604 14468 20084
rect 14512 19988 14552 20236
rect 14638 20064 14678 20178
rect 14512 19948 14720 19988
rect 14428 19564 14498 19604
rect 14458 19299 14498 19564
rect 14596 19220 14636 19892
rect 14680 19468 14720 19948
rect 14008 18604 14384 18644
rect 14428 19180 14636 19220
rect 13588 18414 13628 18528
rect 13420 17838 13460 17952
rect 13798 17740 13964 17780
rect 13504 16780 13544 17044
rect 13336 16492 13544 16532
rect 13336 15724 13376 16148
rect 13504 15436 13544 16492
rect 13714 15264 13754 15378
rect 13252 14764 13376 14804
rect 13168 14668 13292 14708
rect 13000 14380 13063 14420
rect 13023 14019 13063 14380
rect 13126 14094 13166 14208
rect 12832 13900 12956 13940
rect 12916 13324 13166 13364
rect 13126 13180 13166 13324
rect 13252 13132 13292 14668
rect 13336 13420 13376 14764
rect 13924 14036 13964 17740
rect 14008 16340 14048 18604
rect 14092 17740 14132 17972
rect 14092 17644 14216 17684
rect 14092 16396 14132 17644
rect 14344 17108 14384 18548
rect 14428 17492 14468 19180
rect 14680 17836 14720 19316
rect 14764 18508 14804 20620
rect 14848 19852 14888 20468
rect 14848 19084 14888 19241
rect 14764 17740 14888 17780
rect 14764 17644 14804 17740
rect 14932 17684 14972 23020
rect 15184 20620 15350 20660
rect 15100 20044 15266 20084
rect 15131 19225 15171 19360
rect 15058 19084 15224 19124
rect 15184 18260 15224 19084
rect 15436 18644 15476 25446
rect 15856 24844 15896 25446
rect 16276 23404 16316 25446
rect 16696 23060 16736 25446
rect 16696 23020 16820 23060
rect 15352 18604 15476 18644
rect 15268 18318 15308 18432
rect 15142 18220 15224 18260
rect 15142 17740 15182 18220
rect 14848 17644 14972 17684
rect 14512 17548 14804 17588
rect 14428 17452 14720 17492
rect 14176 17068 14384 17108
rect 14008 16300 14132 16340
rect 14008 14574 14048 15476
rect 13840 13996 13964 14036
rect 14092 14036 14132 16300
rect 14176 15724 14216 17068
rect 14470 16409 14510 16820
rect 14389 15092 14429 15648
rect 14680 15572 14720 17452
rect 14764 16204 14804 17548
rect 14680 15532 14804 15572
rect 14389 15052 14636 15092
rect 14092 13996 14216 14036
rect 14344 13997 14384 14132
rect 13588 13806 13628 13920
rect 13840 13902 13880 13996
rect 14470 13804 14510 14036
rect 13504 13196 13544 13331
rect 12664 13036 12788 13076
rect 12538 12940 12620 12980
rect 12580 12788 12620 12940
rect 12748 12912 12788 13036
rect 12580 12748 12884 12788
rect 12844 12692 12884 12748
rect 12832 12652 12884 12692
rect 13840 12652 13880 13076
rect 12076 11788 12620 11828
rect 12370 11500 12410 11636
rect 12160 11022 12200 11136
rect 12328 10924 12368 11156
rect 12580 11116 12620 11788
rect 12160 10350 12200 10464
rect 11656 10196 11696 10292
rect 11740 10252 12116 10292
rect 11656 10156 11822 10196
rect 11824 9332 11864 10071
rect 11824 9292 12032 9332
rect 11572 9100 11810 9140
rect 11404 8620 11444 8755
rect 11488 8621 11528 8756
rect 11770 8719 11810 9100
rect 11614 8334 11654 8448
rect 11908 8180 11948 9236
rect 11992 8524 12032 9292
rect 11656 8140 11948 8180
rect 11236 7796 11276 7892
rect 11320 7852 11444 7892
rect 11236 7756 11360 7796
rect 11404 7180 11444 7852
rect 11698 7796 11738 7988
rect 11488 7756 11738 7796
rect 10396 6796 10436 7146
rect 10732 6990 10772 7104
rect 11488 7028 11528 7756
rect 11908 7180 11948 7796
rect 12076 7372 12116 10252
rect 12244 10252 12464 10292
rect 12244 8620 12284 10252
rect 12328 7988 12368 10196
rect 12424 10156 12464 10252
rect 12664 10060 12704 12525
rect 12748 11692 12788 12500
rect 12832 11404 12872 12652
rect 12748 10444 12788 11060
rect 12832 10196 12872 11156
rect 12748 10156 12872 10196
rect 12916 10156 12956 11540
rect 13126 10964 13166 11012
rect 13000 10924 13166 10964
rect 12832 9966 12872 10080
rect 13000 9620 13040 10924
rect 13168 10350 13208 10464
rect 12832 9580 13040 9620
rect 12664 9102 12704 9216
rect 12538 8668 12578 8803
rect 12664 8524 12704 8660
rect 12244 7948 12368 7988
rect 12244 7132 12284 7948
rect 12832 7756 12872 9580
rect 13252 9524 13292 10292
rect 13336 10196 13376 11828
rect 13840 10868 13880 11732
rect 13924 10964 13964 11636
rect 14008 11020 14048 13076
rect 14092 12366 14132 12480
rect 14260 11656 14300 13172
rect 14344 13036 14384 13172
rect 14512 12366 14552 12480
rect 14596 12364 14636 15052
rect 14680 11732 14720 15532
rect 14848 14188 14888 17644
rect 15016 17550 15056 17664
rect 15184 16204 15224 16916
rect 14932 14092 14972 15860
rect 15352 15572 15392 18604
rect 15436 17972 15476 18548
rect 15520 18068 15560 21716
rect 15688 20756 15728 21524
rect 15604 20716 15728 20756
rect 15604 20044 15644 20716
rect 15940 19948 15980 21524
rect 16192 21486 16232 21600
rect 16528 20756 16568 21620
rect 16612 21580 16652 21716
rect 16444 20716 16652 20756
rect 15604 19200 15644 19314
rect 16108 19276 16148 20084
rect 16444 20044 16484 20716
rect 16192 19339 16232 19988
rect 16696 19604 16736 20756
rect 16695 19564 16736 19604
rect 16192 19299 16274 19339
rect 16234 19276 16274 19299
rect 16695 19243 16735 19564
rect 16780 19468 16820 23020
rect 17116 21772 17156 25446
rect 17536 23060 17576 25446
rect 17368 23020 17576 23060
rect 16864 21004 16904 21524
rect 17074 21484 17114 21620
rect 17200 19412 17240 22964
rect 17284 21390 17324 21504
rect 17116 19372 17240 19412
rect 15720 19086 15760 19200
rect 15856 18412 15896 18548
rect 15520 18028 15644 18068
rect 15436 17932 15560 17972
rect 15604 17876 15644 18028
rect 15520 17836 15644 17876
rect 15436 15628 15476 15764
rect 15016 15436 15056 15572
rect 15352 15532 15476 15572
rect 15520 15532 15560 17836
rect 15814 17740 15854 17876
rect 15711 17396 15751 17732
rect 16024 17705 16064 17876
rect 15688 17356 15751 17396
rect 15688 17164 15728 17356
rect 15604 15820 15644 17060
rect 16024 16782 16064 16896
rect 16108 16244 16148 17588
rect 16360 17548 16400 17780
rect 16276 16780 16400 16820
rect 16024 16204 16148 16244
rect 15604 15534 15644 15648
rect 15016 14284 15056 14516
rect 15100 14324 15140 14708
rect 15184 14496 15224 14610
rect 15310 14420 15350 14612
rect 15226 14380 15350 14420
rect 15226 14324 15266 14380
rect 15436 14324 15476 15532
rect 15100 14284 15170 14324
rect 15226 14284 15308 14324
rect 15130 13948 15170 14284
rect 15268 13844 15308 14284
rect 14848 13804 15308 13844
rect 15352 12980 15392 14324
rect 15436 14284 15560 14324
rect 15184 12940 15392 12980
rect 14638 11692 14720 11732
rect 14092 11212 14132 11540
rect 13924 10924 14048 10964
rect 13840 10828 13964 10868
rect 13924 10196 13964 10828
rect 13336 10156 13460 10196
rect 12916 8908 12956 9524
rect 13252 9484 13376 9524
rect 13420 9236 13460 10156
rect 13588 10031 13628 10166
rect 13672 10156 13964 10196
rect 13336 9196 13460 9236
rect 13336 8660 13376 9196
rect 13336 8620 13460 8660
rect 13672 8620 13712 8948
rect 13588 8430 13628 8544
rect 14008 7900 14048 10924
rect 14260 10388 14300 11540
rect 14638 11348 14678 11692
rect 14764 11500 14804 12500
rect 14932 11683 14972 12788
rect 14848 11404 14888 11583
rect 14092 10348 14300 10388
rect 14596 11308 14678 11348
rect 14176 9484 14216 10196
rect 14260 8948 14300 10100
rect 14092 8908 14300 8948
rect 14596 8756 14636 11308
rect 14680 10156 14720 11252
rect 14596 8716 14678 8756
rect 14638 8668 14678 8716
rect 14176 8046 14216 8160
rect 14764 7900 14804 8756
rect 14932 8620 14972 9236
rect 14848 8430 14888 8544
rect 15016 8180 15056 12020
rect 15184 11212 15224 12940
rect 15436 11980 15476 14228
rect 15520 11884 15560 14284
rect 15604 14132 15644 15284
rect 15688 14284 15728 15572
rect 16024 15438 16064 15552
rect 15856 14284 15896 14516
rect 15604 14092 15728 14132
rect 15688 14084 15728 14092
rect 15688 14044 15760 14084
rect 15604 13364 15644 14036
rect 16108 13902 16148 14228
rect 16234 13996 16274 14324
rect 16360 13940 16400 16780
rect 16528 13996 16568 18644
rect 16696 18556 16736 18740
rect 16654 17645 16694 17780
rect 16696 16974 16736 17088
rect 16780 16396 16820 17684
rect 17032 17068 17072 17876
rect 16612 14574 16652 14688
rect 16696 14420 16736 15476
rect 16864 14668 16904 15572
rect 16695 14380 16736 14420
rect 16695 14009 16735 14380
rect 16276 13900 16400 13940
rect 15604 13324 15728 13364
rect 15184 8524 15224 10772
rect 14932 8140 15056 8180
rect 15268 8140 15308 11828
rect 15352 11788 15560 11828
rect 15520 11692 15560 11788
rect 15604 11404 15644 13194
rect 15688 13172 15728 13324
rect 15688 13132 15938 13172
rect 16008 13132 16148 13172
rect 15436 10444 15476 11060
rect 15520 10062 15560 10176
rect 15688 10004 15728 13132
rect 16024 12508 16064 12980
rect 16108 12652 16148 13132
rect 16276 12460 16316 13900
rect 16402 12980 16442 13172
rect 16360 12940 16442 12980
rect 15940 11252 15980 11732
rect 15856 11212 15980 11252
rect 15856 10997 15896 11212
rect 15688 9964 15770 10004
rect 15730 9492 15770 9964
rect 15352 8716 15392 9428
rect 15814 9140 15854 9493
rect 15688 9100 15854 9140
rect 15520 8468 15560 8564
rect 15688 8524 15728 9100
rect 15940 8620 15980 11212
rect 16360 11116 16400 12940
rect 16528 11692 16568 13268
rect 16959 12980 16999 13207
rect 16948 12940 16999 12980
rect 16948 12748 16988 12940
rect 16738 11636 16778 11684
rect 16696 11596 16778 11636
rect 16696 10196 16736 11596
rect 17116 10964 17156 19372
rect 17200 18604 17240 19261
rect 17368 19220 17408 23020
rect 17452 21678 17492 21792
rect 17818 21236 17858 21521
rect 17746 21196 17858 21236
rect 17746 20620 17786 21196
rect 17620 19872 17660 19986
rect 17823 19700 17863 20083
rect 17956 19988 17996 25446
rect 18376 23020 18416 25446
rect 18628 23060 18668 23252
rect 18796 23116 18836 25446
rect 18460 23020 18668 23060
rect 18040 21390 18080 21504
rect 17956 19948 18080 19988
rect 17620 19660 17863 19700
rect 17284 19180 17408 19220
rect 17284 19028 17324 19180
rect 17536 19124 17576 19241
rect 17368 19084 17576 19124
rect 17284 18988 17576 19028
rect 17284 16972 17324 17780
rect 17452 17045 17492 18836
rect 17536 16492 17576 18988
rect 17620 17742 17660 19660
rect 17830 19488 17870 19602
rect 17819 19181 17859 19316
rect 17704 17684 17744 18932
rect 17956 18700 17996 19892
rect 18040 18892 18080 19948
rect 18208 18796 18248 19412
rect 18292 18836 18332 19508
rect 18376 19182 18416 19296
rect 18292 18796 18416 18836
rect 18124 18548 18164 18567
rect 18040 18508 18164 18548
rect 17872 17740 17912 18356
rect 17620 17644 17744 17684
rect 17200 16302 17240 16416
rect 17368 14284 17408 16292
rect 17536 14188 17576 14516
rect 17368 14092 17576 14132
rect 17200 13902 17240 14016
rect 17368 13036 17408 13940
rect 17326 12404 17366 12452
rect 17284 12364 17366 12404
rect 17284 12308 17324 12364
rect 17200 12268 17324 12308
rect 17200 11692 17240 12268
rect 17074 10924 17156 10964
rect 17074 10444 17114 10924
rect 16864 10196 16904 10244
rect 16612 10156 16736 10196
rect 16780 10156 16904 10196
rect 17320 10156 17360 10388
rect 16318 9484 16358 9620
rect 16192 9294 16232 9408
rect 16612 8660 16652 10156
rect 16780 10004 16820 10156
rect 17452 10100 17492 14036
rect 17536 13996 17576 14092
rect 17620 12692 17660 17644
rect 18040 16436 18080 18508
rect 18292 18452 18332 18596
rect 18376 18556 18416 18796
rect 18124 16532 18164 18452
rect 18208 18412 18332 18452
rect 18208 17260 18248 18412
rect 18292 17043 18332 18356
rect 18460 18068 18500 23020
rect 18544 18412 18584 20180
rect 19216 19372 19256 25446
rect 19636 23444 19676 25446
rect 19552 23404 19676 23444
rect 19552 21388 19592 23404
rect 18628 19086 18668 19200
rect 19384 18508 19424 18643
rect 18376 18028 18500 18068
rect 18544 18316 18836 18356
rect 18880 18316 19214 18356
rect 18124 16492 18248 16532
rect 18040 16396 18164 16436
rect 17746 14496 17786 14610
rect 17872 14420 17912 15572
rect 18040 15342 18080 16292
rect 18124 15572 18164 16396
rect 18376 15668 18416 18028
rect 18544 17972 18584 18316
rect 18502 17932 18584 17972
rect 18502 17740 18542 17932
rect 18880 17740 18920 18316
rect 19468 18222 19508 18336
rect 19468 17068 19508 17204
rect 18712 16396 19340 16436
rect 19300 16204 19340 16396
rect 18880 16108 19172 16148
rect 18376 15628 18584 15668
rect 18124 15532 18416 15572
rect 18292 14708 18332 15532
rect 18544 15476 18584 15628
rect 18670 15552 18710 15666
rect 18544 15436 18668 15476
rect 17746 14380 17912 14420
rect 18208 14668 18332 14708
rect 18376 14668 18416 15284
rect 18502 14669 18542 14804
rect 17746 14188 17786 14380
rect 17819 13708 17859 14039
rect 18208 13996 18248 14668
rect 18544 14121 18584 14256
rect 17704 13228 17855 13268
rect 17815 13169 17855 13228
rect 18123 13132 18164 13194
rect 17872 12788 17912 13076
rect 17536 12652 17660 12692
rect 17836 12748 17912 12788
rect 17836 12508 17876 12748
rect 18040 12500 18080 13076
rect 18123 13061 18163 13132
rect 18208 12556 18248 13844
rect 18502 13804 18542 14021
rect 18292 12980 18332 13172
rect 18292 12940 18584 12980
rect 18040 12460 18164 12500
rect 17956 11406 17996 11520
rect 17872 11022 17912 11136
rect 16696 9964 16820 10004
rect 17284 10060 17492 10100
rect 16696 8908 16736 9964
rect 16780 9196 16820 9524
rect 17284 9475 17324 10060
rect 17536 9964 17576 10099
rect 17620 10060 17660 10196
rect 17704 9676 17744 10964
rect 18040 10868 18080 12404
rect 18292 11884 18332 12884
rect 18376 11500 18416 12788
rect 18544 12652 18584 12940
rect 18628 11732 18668 15436
rect 18796 14764 18836 15860
rect 19132 15724 19172 16108
rect 19468 15532 19508 16820
rect 18880 14132 18920 14900
rect 19216 14574 19256 14688
rect 18880 14092 19088 14132
rect 19468 13900 19508 14036
rect 18712 13036 18752 13195
rect 18880 12980 18920 13748
rect 19552 13036 19592 13197
rect 18460 11692 18668 11732
rect 18712 12940 18920 12980
rect 18124 10944 18164 11058
rect 18040 10828 18164 10868
rect 17452 9484 17492 9620
rect 17788 9580 17828 10772
rect 18040 10156 18080 10292
rect 18124 9484 18164 10828
rect 18208 10062 18248 10176
rect 18376 9390 18416 9504
rect 17956 8908 17996 9236
rect 16612 8620 16820 8660
rect 18208 8620 18248 9332
rect 18460 8756 18500 11692
rect 18712 11636 18752 12940
rect 19552 12366 19592 12480
rect 19384 12174 19424 12288
rect 18586 11596 18752 11636
rect 18880 10348 18920 11060
rect 18964 10828 19004 11732
rect 19048 11020 19088 11636
rect 19174 10964 19214 10997
rect 19132 10924 19214 10964
rect 18628 10062 18668 10176
rect 18712 9716 18752 10100
rect 18628 9676 18752 9716
rect 18712 9484 18752 9620
rect 19048 9524 19088 10196
rect 19132 9964 19172 10924
rect 19300 9908 19340 10196
rect 19284 9868 19340 9908
rect 19048 9484 19130 9524
rect 19090 9340 19130 9484
rect 19284 9475 19324 9868
rect 19468 9716 19508 10196
rect 19384 9676 19508 9716
rect 19552 9580 19592 10772
rect 19636 9332 19676 22964
rect 20056 21580 20096 25446
rect 19839 18508 19879 18643
rect 19804 18316 20012 18356
rect 19804 17780 19844 18316
rect 19762 17740 19844 17780
rect 19762 17715 19802 17740
rect 20140 17396 20180 23156
rect 20476 21484 20516 25446
rect 20896 20140 20936 25446
rect 21316 23060 21356 25446
rect 21316 23020 21608 23060
rect 21736 23020 21776 25446
rect 22156 24556 22196 25446
rect 22576 25132 22616 25446
rect 22996 25228 23036 25446
rect 23416 25036 23456 25446
rect 19888 17356 20180 17396
rect 19720 16972 19760 17108
rect 19888 17012 19928 17356
rect 20014 17068 20054 17300
rect 20896 17260 20936 17588
rect 19888 16972 20012 17012
rect 20140 16974 20180 17088
rect 19888 15438 19928 15552
rect 19972 12413 20012 16972
rect 20628 16916 20668 17067
rect 20628 16876 20852 16916
rect 20392 16686 20432 16800
rect 20560 16780 20768 16820
rect 20560 16532 20600 16780
rect 20140 16492 20600 16532
rect 20140 16204 20180 16492
rect 20812 16148 20852 16876
rect 21568 16244 21608 23020
rect 23836 22388 23876 25446
rect 24256 24940 24296 25446
rect 24676 23116 24716 25446
rect 25096 23212 25136 25446
rect 23836 22348 24044 22388
rect 24004 19276 24044 22348
rect 21484 16148 21524 16244
rect 21568 16204 21692 16244
rect 20644 16108 21524 16148
rect 20224 14668 20432 14708
rect 20140 12558 20180 12672
rect 20224 12308 20264 14668
rect 20644 14612 20684 16108
rect 20728 15532 20768 16052
rect 20896 16012 21356 16052
rect 20896 15820 20936 16012
rect 21568 15918 21608 16032
rect 21652 15860 21692 16204
rect 21568 15820 21692 15860
rect 20644 14572 20768 14612
rect 20308 13902 20348 14016
rect 20392 12980 20432 13076
rect 20392 12940 20474 12980
rect 20434 12652 20474 12940
rect 20350 12525 20390 12535
rect 20644 12525 20684 14572
rect 20896 13844 20936 15572
rect 21484 14094 21524 14208
rect 20728 13420 20768 13844
rect 20896 13804 21146 13844
rect 21106 13385 21146 13804
rect 21568 13460 21608 15820
rect 21904 15150 21944 15264
rect 21778 14708 21818 14852
rect 21778 14668 21944 14708
rect 21652 13996 21692 14132
rect 21778 13902 21818 14016
rect 21904 13900 21944 14668
rect 21484 13420 21608 13460
rect 21316 12980 21356 13268
rect 21316 12940 21524 12980
rect 21484 12748 21524 12940
rect 20350 12485 20684 12525
rect 20224 12268 20348 12308
rect 19804 11597 19844 11732
rect 20308 11020 20348 12268
rect 19972 10734 20012 10848
rect 20812 10156 20852 11540
rect 20980 11500 21020 11636
rect 21183 11500 21223 11684
rect 21316 11598 21356 11712
rect 21087 10176 21127 10290
rect 20644 9870 20684 9984
rect 20812 9964 21230 10004
rect 19972 9390 20012 9504
rect 20812 9484 20852 9964
rect 21652 9484 21692 10868
rect 19174 9292 19676 9332
rect 18460 8716 18668 8756
rect 18964 8716 19004 9236
rect 19174 8908 19214 9292
rect 18418 8526 18458 8640
rect 21988 8620 22028 9236
rect 15352 8428 15560 8468
rect 18796 8430 18836 8544
rect 12370 7086 12410 7200
rect 11404 6988 11528 7028
rect 11404 6894 11444 6988
rect 7456 6220 7664 6260
<< metal3 >>
rect 7372 25228 23036 25268
rect 8548 25132 22616 25172
rect 11740 25036 23456 25076
rect 13420 24940 24296 24980
rect 6448 24844 15896 24884
rect 6952 24556 22196 24596
rect 6364 24364 12116 24404
rect 5272 24172 10856 24212
rect 9052 23404 16316 23444
rect 18628 23212 25136 23252
rect 10900 23116 18836 23156
rect 20140 23116 24716 23156
rect 10900 22964 10940 23116
rect 14596 22964 14636 23060
rect 18376 22964 18416 23060
rect 21736 22964 21776 23060
rect 10396 22924 10940 22964
rect 11824 22924 14636 22964
rect 17200 22924 18416 22964
rect 19636 22924 21776 22964
rect 13756 21772 14636 21812
rect 17116 21772 17492 21812
rect 5356 21676 9596 21716
rect 9685 21676 16652 21716
rect 9472 21580 12536 21620
rect 13210 21580 16568 21620
rect 17074 21580 20096 21620
rect 8044 21484 12032 21524
rect 12160 21484 15728 21524
rect 15940 21484 17324 21524
rect 18040 21484 20516 21524
rect 8632 21388 19592 21428
rect 11110 21004 16904 21044
rect 10564 20908 12872 20948
rect 11488 20812 11696 20852
rect 6616 20716 12980 20756
rect 14764 20716 17786 20756
rect 12940 20660 12980 20716
rect 7288 20620 7496 20660
rect 12940 20620 14510 20660
rect 6868 20524 9764 20564
rect 14470 20428 14888 20468
rect 7876 20236 10352 20276
rect 10312 20180 10352 20236
rect 6784 20140 7328 20180
rect 8212 20140 9008 20180
rect 10312 20140 12116 20180
rect 13588 20140 14804 20180
rect 18544 20140 20936 20180
rect 7162 20044 8840 20084
rect 9892 20044 13460 20084
rect 14428 20044 16148 20084
rect 7036 19948 12788 19988
rect 13672 19948 16232 19988
rect 6868 19852 9932 19892
rect 10564 19852 11276 19892
rect 12940 19852 14384 19892
rect 14596 19852 14888 19892
rect 16108 19852 17660 19892
rect 12940 19796 12980 19852
rect 8884 19756 12980 19796
rect 10144 19660 13208 19700
rect 6858 19564 6972 19604
rect 13168 19468 14132 19508
rect 14260 19468 16820 19508
rect 17830 19468 18332 19508
rect 8632 19372 9428 19412
rect 11320 19372 19256 19412
rect 9178 19276 12704 19316
rect 14680 19276 17859 19316
rect 18376 19276 24044 19316
rect 8800 18932 8840 19220
rect 12160 19180 15644 19220
rect 15720 19180 18668 19220
rect 13924 19084 14888 19124
rect 9220 18988 9764 19028
rect 8632 18892 10268 18932
rect 17704 18892 18080 18932
rect 6112 18796 7160 18836
rect 10648 18796 12200 18836
rect 13252 18796 14216 18836
rect 17452 18796 18248 18836
rect 6112 18740 6152 18796
rect 5776 18700 6152 18740
rect 6280 18700 8588 18740
rect 8968 18700 10100 18740
rect 11656 18700 14804 18740
rect 16696 18700 17996 18740
rect 10060 18644 10100 18700
rect 10060 18604 11822 18644
rect 13168 18604 17240 18644
rect 5776 18508 8924 18548
rect 11488 18452 11528 18548
rect 13588 18508 14384 18548
rect 17620 18508 19879 18548
rect 10900 18412 11528 18452
rect 15268 18412 15896 18452
rect 18124 18412 18584 18452
rect 10900 18220 10940 18412
rect 11236 18316 12032 18356
rect 18292 18316 19508 18356
rect 10144 17932 14132 17972
rect 8528 17836 9344 17876
rect 9976 17684 10016 17876
rect 10816 17836 14720 17876
rect 16024 17836 17660 17876
rect 10816 17780 10856 17836
rect 10354 17740 10856 17780
rect 12244 17740 15854 17780
rect 16528 17740 17912 17780
rect 16528 17684 16568 17740
rect 5440 17644 9008 17684
rect 9220 17644 10016 17684
rect 12940 17644 13208 17684
rect 12940 17588 12980 17644
rect 9622 17548 12980 17588
rect 14764 17588 14804 17684
rect 15016 17644 16568 17684
rect 14764 17548 18080 17588
rect 5146 17356 5816 17396
rect 8044 17356 9848 17396
rect 5776 17300 5816 17356
rect 9808 17300 9848 17356
rect 5776 17260 5984 17300
rect 9220 17260 9512 17300
rect 9808 17260 10688 17300
rect 10816 17260 11192 17300
rect 11278 17260 11696 17300
rect 18208 17260 20936 17300
rect 10900 17164 11444 17204
rect 12664 17164 15728 17204
rect 4852 17068 7244 17108
rect 10480 17068 16736 17108
rect 19468 17068 20180 17108
rect 6280 16972 9932 17012
rect 12076 16972 17324 17012
rect 18040 16972 19760 17012
rect 6448 16876 6740 16916
rect 11740 16876 13166 16916
rect 15184 16876 16064 16916
rect 6784 16780 7244 16820
rect 10480 16780 11108 16820
rect 11404 16780 12284 16820
rect 13504 16780 14510 16820
rect 19468 16780 20432 16820
rect 4768 16684 11024 16724
rect 10228 16588 10688 16628
rect 9388 16492 10772 16532
rect 5776 16300 5936 16340
rect 6196 16300 10016 16340
rect 5776 16204 8756 16244
rect 9472 16204 9848 16244
rect 7876 15956 7916 16148
rect 10396 16052 10436 16436
rect 10564 16396 11276 16436
rect 16780 16396 17240 16436
rect 11488 16204 12956 16244
rect 10554 16108 10668 16148
rect 11656 16108 13376 16148
rect 10060 16012 11108 16052
rect 20728 16012 21608 16052
rect 7204 15916 7916 15956
rect 8338 15820 11444 15860
rect 14932 15820 15644 15860
rect 18796 15820 20936 15860
rect 6364 15724 7664 15764
rect 12652 15724 13964 15764
rect 7456 15628 8672 15668
rect 9472 15628 12410 15668
rect 12496 15628 12872 15668
rect 15436 15628 15644 15668
rect 12328 15572 12368 15628
rect 8422 15532 11276 15572
rect 12328 15532 12956 15572
rect 14389 15532 15560 15572
rect 15688 15532 16064 15572
rect 17872 15532 18710 15572
rect 19888 15532 20936 15572
rect 4516 15436 5816 15476
rect 15016 15436 18080 15476
rect 13714 15244 15644 15284
rect 18376 15244 21944 15284
rect 6784 14956 10604 14996
rect 18502 14764 18836 14804
rect 4684 14668 5312 14708
rect 8884 14668 10604 14708
rect 14008 14668 16904 14708
rect 19216 14668 20264 14708
rect 8380 14572 10184 14612
rect 15016 14476 15896 14516
rect 17536 14476 17786 14516
rect 4852 14380 5816 14420
rect 10900 14284 12368 14324
rect 12454 14284 15056 14324
rect 15352 14284 15728 14324
rect 15856 14284 17408 14324
rect 11404 14188 13166 14228
rect 14848 14188 15476 14228
rect 16108 14188 17576 14228
rect 18544 14188 21524 14228
rect 5524 14092 7160 14132
rect 12328 14092 14972 14132
rect 20644 14092 21692 14132
rect 5128 13996 5396 14036
rect 10816 13996 11864 14036
rect 12076 13996 13880 14036
rect 14470 13996 16148 14036
rect 16528 13996 17492 14036
rect 18208 13940 18248 14036
rect 20308 13996 21818 14036
rect 13588 13900 18248 13940
rect 19468 13900 21944 13940
rect 10900 13804 11528 13844
rect 11824 13804 14510 13844
rect 18208 13804 20768 13844
rect 11152 13708 14636 13748
rect 17788 13708 17923 13748
rect 11488 13612 12284 13652
rect 7876 13516 12368 13556
rect 6280 13420 6656 13460
rect 10164 13420 10278 13460
rect 10648 13420 10716 13460
rect 11992 13420 13376 13460
rect 10648 13364 10688 13420
rect 4600 13324 5228 13364
rect 6700 13324 15728 13364
rect 4768 13228 5816 13268
rect 8968 13228 13544 13268
rect 4684 13132 8840 13172
rect 9136 13132 12116 13172
rect 12328 13132 14300 13172
rect 17788 13132 18164 13172
rect 4432 13036 12980 13076
rect 12940 12980 12980 13036
rect 13084 13036 13880 13076
rect 14008 13036 16064 13076
rect 17368 13036 17912 13076
rect 18040 13036 18752 13076
rect 19552 13036 20432 13076
rect 13084 12980 13124 13036
rect 16024 12980 16064 13036
rect 5776 12940 6824 12980
rect 10218 12940 10332 12980
rect 10470 12940 10584 12980
rect 8716 12844 12200 12884
rect 5440 12748 7160 12788
rect 5860 12692 5900 12748
rect 5860 12652 5928 12692
rect 9579 12652 10184 12692
rect 5944 12556 9932 12596
rect 12748 12500 12788 12980
rect 12940 12940 13124 12980
rect 15996 12940 16064 12980
rect 18040 12884 18080 13036
rect 18040 12844 18332 12884
rect 14932 12748 21524 12788
rect 16108 12652 20180 12692
rect 6364 12460 11192 12500
rect 12748 12460 14132 12500
rect 14512 12460 19592 12500
rect 6532 12364 11864 12404
rect 14596 12364 18080 12404
rect 5440 12268 7412 12308
rect 19384 12268 20348 12308
rect 6112 12172 8656 12212
rect 6112 12076 6152 12172
rect 4516 11980 8084 12020
rect 15016 11980 15476 12020
rect 5734 11884 7748 11924
rect 12160 11884 12980 11924
rect 12940 11828 12980 11884
rect 15268 11884 15560 11924
rect 5944 11788 6992 11828
rect 12940 11788 13376 11828
rect 15268 11788 15308 11884
rect 5524 11692 6740 11732
rect 8464 11692 9122 11732
rect 13840 11692 17240 11732
rect 19804 11692 21356 11732
rect 7540 11596 9008 11636
rect 9388 11596 13964 11636
rect 19048 11596 21020 11636
rect 4852 11500 5480 11540
rect 7372 11500 9344 11540
rect 11236 11500 14048 11540
rect 14260 11500 14804 11540
rect 17956 11500 18416 11540
rect 20812 11500 21223 11540
rect 12822 11404 15644 11444
rect 14092 11212 15896 11252
rect 9178 11116 12200 11156
rect 12328 11116 17912 11156
rect 8243 11020 10772 11060
rect 6028 10924 7106 10964
rect 10984 10924 11612 10964
rect 17704 10924 18164 10964
rect 18964 10828 20012 10868
rect 10564 10732 17828 10772
rect 9556 10636 10100 10676
rect 12160 10444 12788 10484
rect 13168 10444 15476 10484
rect 11152 10348 18920 10388
rect 11152 10292 11192 10348
rect 9892 10252 11192 10292
rect 11656 10252 12956 10292
rect 13252 10252 14720 10292
rect 8128 10156 9176 10196
rect 10354 10156 12956 10196
rect 14176 10156 17744 10196
rect 18040 10156 18248 10196
rect 18628 10156 19088 10196
rect 19300 10156 21127 10196
rect 4390 10060 5816 10100
rect 6952 10060 10184 10100
rect 10438 10060 12704 10100
rect 12792 10060 13628 10100
rect 17620 10060 18752 10100
rect 5776 9964 6068 10004
rect 6784 9964 7412 10004
rect 17536 9964 20684 10004
rect 8128 9868 14636 9908
rect 6364 9772 8672 9812
rect 5776 9676 5984 9716
rect 5440 9580 6824 9620
rect 7036 9580 12284 9620
rect 16318 9580 16736 9620
rect 17788 9580 18752 9620
rect 6248 9484 6908 9524
rect 7204 9484 8336 9524
rect 8632 9484 9848 9524
rect 17452 9484 18416 9524
rect 19972 9484 21692 9524
rect 6448 9388 7412 9428
rect 15352 9388 16232 9428
rect 6700 9292 7832 9332
rect 11236 9292 18248 9332
rect 11908 9196 12704 9236
rect 14932 9196 19004 9236
rect 6868 9004 8672 9044
rect 4936 8908 5594 8948
rect 5682 8908 5796 8948
rect 8212 8908 8840 8948
rect 10228 8908 11108 8948
rect 13672 8908 16736 8948
rect 4768 8812 9344 8852
rect 4768 8620 4808 8812
rect 5188 8716 8420 8756
rect 5188 8660 5228 8716
rect 4978 8620 5228 8660
rect 5356 8620 6908 8660
rect 7204 8620 7916 8660
rect 9892 8564 9932 8852
rect 10312 8716 11528 8756
rect 12538 8716 15392 8756
rect 11404 8620 11948 8660
rect 18418 8620 22028 8660
rect 4684 8524 5228 8564
rect 5440 8524 5816 8564
rect 5944 8524 9764 8564
rect 9892 8524 10016 8564
rect 11992 8524 15224 8564
rect 15688 8524 18836 8564
rect 5944 8468 5984 8524
rect 3928 8428 5984 8468
rect 9892 8428 11654 8468
rect 9724 8236 10226 8276
rect 14176 8140 15308 8180
rect 4012 7948 4514 7988
rect 5692 7948 10184 7988
rect 8417 7852 11276 7892
rect 11152 7756 11528 7796
rect 4852 7180 8336 7220
rect 8548 7180 9092 7220
rect 11404 7180 12410 7220
rect 8296 7124 8336 7180
rect 8296 7084 9344 7124
rect 10060 7084 10772 7124
rect 9304 7028 9344 7084
rect 9304 6988 11444 7028
rect 4474 6892 5732 6932
rect 7457 6796 10436 6836
rect 5776 6604 7496 6644
rect 4012 6412 7748 6452
rect 7204 6316 10352 6356
<< metal4 >>
rect 5776 12940 5816 18548
rect 6952 11788 6992 19604
rect 10144 12652 10184 13460
rect 10312 12940 10352 13556
rect 10564 12940 10604 17780
rect 10648 17260 10688 18836
rect 10648 16108 10688 16628
rect 12916 10060 12956 11444
rect 17788 10732 17828 13748
rect 5776 8908 5816 10004
<< metal5 >>
rect 1480 21862 2440 21986
rect 5887 21862 6273 21986
rect 21007 21862 21393 21986
rect 23000 21862 23960 21986
rect 80 21106 1040 21230
rect 13447 21106 13833 21230
rect 24400 21106 25360 21230
rect 1480 20350 2440 20474
rect 5887 20350 6273 20474
rect 21007 20350 21393 20474
rect 23000 20350 23960 20474
rect 80 19594 1040 19718
rect 13447 19594 13833 19718
rect 24400 19594 25360 19718
rect 1480 18838 2440 18962
rect 5887 18838 6273 18962
rect 21007 18838 21393 18962
rect 23000 18838 23960 18962
rect 80 18082 1040 18206
rect 13447 18082 13833 18206
rect 24400 18082 25360 18206
rect 1480 17326 2440 17450
rect 5887 17326 6273 17450
rect 21007 17326 21393 17450
rect 23000 17326 23960 17450
rect 80 16570 1040 16694
rect 13447 16570 13833 16694
rect 24400 16570 25360 16694
rect 1480 15814 2440 15938
rect 5887 15814 6273 15938
rect 21007 15814 21393 15938
rect 23000 15814 23960 15938
rect 80 15058 1040 15182
rect 13447 15058 13833 15182
rect 24400 15058 25360 15182
rect 1480 14302 2440 14426
rect 5887 14302 6273 14426
rect 21007 14302 21393 14426
rect 23000 14302 23960 14426
rect 80 13546 1040 13670
rect 13447 13546 13833 13670
rect 24400 13546 25360 13670
rect 1480 12790 2440 12914
rect 5887 12790 6273 12914
rect 21007 12790 21393 12914
rect 23000 12790 23960 12914
rect 80 12034 1040 12158
rect 13447 12034 13833 12158
rect 24400 12034 25360 12158
rect 1480 11278 2440 11402
rect 5887 11278 6273 11402
rect 21007 11278 21393 11402
rect 23000 11278 23960 11402
rect 80 10522 1040 10646
rect 13447 10522 13833 10646
rect 24400 10522 25360 10646
rect 1480 9766 2440 9890
rect 5887 9766 6273 9890
rect 21007 9766 21393 9890
rect 23000 9766 23960 9890
rect 80 9010 1040 9134
rect 13447 9010 13833 9134
rect 24400 9010 25360 9134
rect 1480 8254 2440 8378
rect 5887 8254 6273 8378
rect 21007 8254 21393 8378
rect 23000 8254 23960 8378
rect 80 7498 1040 7622
rect 13447 7498 13833 7622
rect 24400 7498 25360 7622
rect 1480 6742 2440 6866
rect 5887 6742 6273 6866
rect 21007 6742 21393 6866
rect 23000 6742 23960 6866
rect 80 5986 1040 6110
rect 13447 5986 13833 6110
rect 24400 5986 25360 6110
rect 1480 5230 2440 5354
rect 5887 5230 6273 5354
rect 21007 5230 21393 5354
rect 23000 5230 23960 5354
rect 80 4474 1040 4598
rect 13447 4474 13833 4598
rect 24400 4474 25360 4598
rect 1480 3718 2440 3842
rect 5887 3718 6273 3842
rect 21007 3718 21393 3842
rect 23000 3718 23960 3842
<< metal6 >>
rect 60 480 1060 25224
rect 1460 1880 2460 23824
rect 5860 480 6300 25224
rect 13420 480 13860 25224
rect 20980 480 21420 25224
rect 22980 1880 23980 23824
rect 24380 480 25380 25224
<< metal7 >>
rect 60 24224 25380 25224
rect 1460 22824 23980 23824
rect 60 21394 25380 21834
rect 60 13834 25380 14274
rect 60 6274 25380 6714
rect 1460 1880 23980 2880
rect 60 480 25380 1480
use sg13g2_a21o_1  sg13g2_a21o_1_0
timestamp 1754861848
transform 1 0 11040 0 1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  sg13g2_a21oi_1_0
timestamp 1754861848
transform 1 0 3840 0 1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  sg13g2_a22oi_1_0
timestamp 1754861848
transform 1 0 9696 0 1 8316
box -48 -56 624 834
use sg13g2_and2_1  sg13g2_and2_1_0
timestamp 1754861848
transform 1 0 11520 0 -1 8316
box -48 -56 528 834
use sg13g2_and2_2  sg13g2_and2_2_0
timestamp 1754861848
transform 1 0 5856 0 1 8316
box -48 -56 624 834
use sg13g2_buf_1  sg13g2_buf_1_0
timestamp 1754861848
transform 1 0 16800 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_1
timestamp 1754861848
transform 1 0 18048 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_2
timestamp 1754861848
transform 1 0 13920 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_3
timestamp 1754861848
transform 1 0 14688 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_4
timestamp 1754861848
transform 1 0 18528 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_5
timestamp 1754861848
transform 1 0 18912 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_6
timestamp 1754861848
transform 1 0 11808 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_7
timestamp 1754861848
transform 1 0 5856 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_8
timestamp 1754861848
transform 1 0 12288 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_9
timestamp 1754861848
transform 1 0 11712 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_10
timestamp 1754861848
transform 1 0 10080 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_11
timestamp 1754861848
transform 1 0 4608 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_12
timestamp 1754861848
transform 1 0 4416 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_13
timestamp 1754861848
transform 1 0 7104 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_14
timestamp 1754861848
transform 1 0 6720 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_15
timestamp 1754861848
transform 1 0 11040 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_16
timestamp 1754861848
transform 1 0 8352 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_17
timestamp 1754861848
transform 1 0 8352 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_18
timestamp 1754861848
transform 1 0 9408 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_19
timestamp 1754861848
transform 1 0 8736 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_20
timestamp 1754861848
transform 1 0 11616 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_21
timestamp 1754861848
transform 1 0 6240 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_22
timestamp 1754861848
transform 1 0 7968 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_23
timestamp 1754861848
transform 1 0 17952 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_24
timestamp 1754861848
transform 1 0 13440 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_25
timestamp 1754861848
transform 1 0 15072 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_26
timestamp 1754861848
transform 1 0 16800 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_27
timestamp 1754861848
transform 1 0 14400 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_28
timestamp 1754861848
transform 1 0 14016 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_29
timestamp 1754861848
transform 1 0 17760 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_30
timestamp 1754861848
transform 1 0 18336 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_31
timestamp 1754861848
transform 1 0 17184 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_32
timestamp 1754861848
transform 1 0 17280 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_33
timestamp 1754861848
transform 1 0 17280 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_34
timestamp 1754861848
transform 1 0 5856 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_35
timestamp 1754861848
transform 1 0 12672 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_36
timestamp 1754861848
transform 1 0 19872 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_37
timestamp 1754861848
transform 1 0 11712 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  sg13g2_buf_1_38
timestamp 1754861848
transform 1 0 21216 0 1 12852
box -48 -56 432 834
use sg13g2_buf_2  sg13g2_buf_2_0
timestamp 1754861848
transform 1 0 18048 0 1 8316
box -48 -56 528 834
use sg13g2_buf_4  sg13g2_buf_4_0
timestamp 1754861848
transform 1 0 13728 0 1 11340
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_1
timestamp 1754861848
transform 1 0 17568 0 -1 9828
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_2
timestamp 1754861848
transform 1 0 4704 0 1 11340
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_3
timestamp 1754861848
transform 1 0 10560 0 1 9828
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_4
timestamp 1754861848
transform 1 0 9216 0 -1 9828
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_5
timestamp 1754861848
transform 1 0 7104 0 -1 8316
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_6
timestamp 1754861848
transform 1 0 10272 0 1 8316
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_7
timestamp 1754861848
transform 1 0 11232 0 -1 14364
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_8
timestamp 1754861848
transform 1 0 10464 0 -1 14364
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_9
timestamp 1754861848
transform 1 0 4800 0 -1 15876
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_10
timestamp 1754861848
transform 1 0 4992 0 1 15876
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_11
timestamp 1754861848
transform 1 0 5568 0 -1 15876
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_12
timestamp 1754861848
transform 1 0 9120 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_13
timestamp 1754861848
transform 1 0 10080 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_14
timestamp 1754861848
transform 1 0 6624 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_15
timestamp 1754861848
transform 1 0 7488 0 1 18900
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_16
timestamp 1754861848
transform 1 0 13824 0 -1 15876
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_17
timestamp 1754861848
transform 1 0 13248 0 -1 14364
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_18
timestamp 1754861848
transform 1 0 16032 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_19
timestamp 1754861848
transform 1 0 16128 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_20
timestamp 1754861848
transform 1 0 13920 0 -1 12852
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_21
timestamp 1754861848
transform 1 0 19008 0 -1 12852
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_22
timestamp 1754861848
transform 1 0 7584 0 -1 12852
box -48 -56 816 834
use sg13g2_buf_4  sg13g2_buf_4_23
timestamp 1754861848
transform 1 0 10560 0 -1 12852
box -48 -56 816 834
use sg13g2_buf_8  sg13g2_buf_8_0
timestamp 1754861848
transform 1 0 20160 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_1
timestamp 1754861848
transform 1 0 10560 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_2
timestamp 1754861848
transform 1 0 19008 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_3
timestamp 1754861848
transform 1 0 20256 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_4
timestamp 1754861848
transform 1 0 17184 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_5
timestamp 1754861848
transform 1 0 11808 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  sg13g2_buf_8_6
timestamp 1754861848
transform 1 0 12480 0 1 11340
box -48 -56 1296 834
use sg13g2_decap_4  sg13g2_decap_4_0
timestamp 1754861848
transform 1 0 21504 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_1
timestamp 1754861848
transform 1 0 21504 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_2
timestamp 1754861848
transform 1 0 21504 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_3
timestamp 1754861848
transform 1 0 14304 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_4
timestamp 1754861848
transform 1 0 6528 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_5
timestamp 1754861848
transform 1 0 4224 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_6
timestamp 1754861848
transform 1 0 3360 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_7
timestamp 1754861848
transform 1 0 3360 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_8
timestamp 1754861848
transform 1 0 4704 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_9
timestamp 1754861848
transform 1 0 4896 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_10
timestamp 1754861848
transform 1 0 4032 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_11
timestamp 1754861848
transform 1 0 4032 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_12
timestamp 1754861848
transform 1 0 4032 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_13
timestamp 1754861848
transform 1 0 4032 0 1 14364
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_14
timestamp 1754861848
transform 1 0 4704 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_15
timestamp 1754861848
transform 1 0 7392 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_16
timestamp 1754861848
transform 1 0 6048 0 1 20412
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_17
timestamp 1754861848
transform 1 0 4704 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_18
timestamp 1754861848
transform 1 0 21696 0 1 15876
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_19
timestamp 1754861848
transform 1 0 21504 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_20
timestamp 1754861848
transform 1 0 21504 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_21
timestamp 1754861848
transform 1 0 21696 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_22
timestamp 1754861848
transform 1 0 18624 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_4  sg13g2_decap_4_23
timestamp 1754861848
transform 1 0 21600 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  sg13g2_decap_8_0
timestamp 1754861848
transform 1 0 18144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_1
timestamp 1754861848
transform 1 0 18816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_2
timestamp 1754861848
transform 1 0 19488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_3
timestamp 1754861848
transform 1 0 21216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_4
timestamp 1754861848
transform 1 0 20832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_5
timestamp 1754861848
transform 1 0 20160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_6
timestamp 1754861848
transform 1 0 20544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_7
timestamp 1754861848
transform 1 0 19488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_8
timestamp 1754861848
transform 1 0 19872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_9
timestamp 1754861848
transform 1 0 18432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_10
timestamp 1754861848
transform 1 0 19104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_11
timestamp 1754861848
transform 1 0 19776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_12
timestamp 1754861848
transform 1 0 19488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_13
timestamp 1754861848
transform 1 0 20448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_14
timestamp 1754861848
transform 1 0 20160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_15
timestamp 1754861848
transform 1 0 18816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_16
timestamp 1754861848
transform 1 0 20832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_17
timestamp 1754861848
transform 1 0 18144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_18
timestamp 1754861848
transform 1 0 18816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_19
timestamp 1754861848
transform 1 0 19200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_20
timestamp 1754861848
transform 1 0 17856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_21
timestamp 1754861848
transform 1 0 18528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_22
timestamp 1754861848
transform 1 0 21120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_23
timestamp 1754861848
transform 1 0 17472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_24
timestamp 1754861848
transform 1 0 18144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_25
timestamp 1754861848
transform 1 0 20832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_26
timestamp 1754861848
transform 1 0 17472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_27
timestamp 1754861848
transform 1 0 20160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_28
timestamp 1754861848
transform 1 0 17472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_29
timestamp 1754861848
transform 1 0 17760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_30
timestamp 1754861848
transform 1 0 13824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_31
timestamp 1754861848
transform 1 0 13152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_32
timestamp 1754861848
transform 1 0 12768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_33
timestamp 1754861848
transform 1 0 16128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_34
timestamp 1754861848
transform 1 0 16512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_35
timestamp 1754861848
transform 1 0 12768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_36
timestamp 1754861848
transform 1 0 13440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_37
timestamp 1754861848
transform 1 0 16128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_38
timestamp 1754861848
transform 1 0 15456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_39
timestamp 1754861848
transform 1 0 15456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_40
timestamp 1754861848
transform 1 0 14784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_41
timestamp 1754861848
transform 1 0 13056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_42
timestamp 1754861848
transform 1 0 13440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_43
timestamp 1754861848
transform 1 0 16416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_44
timestamp 1754861848
transform 1 0 14112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_45
timestamp 1754861848
transform 1 0 14784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_46
timestamp 1754861848
transform 1 0 14112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_47
timestamp 1754861848
transform 1 0 15840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_48
timestamp 1754861848
transform 1 0 14784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_49
timestamp 1754861848
transform 1 0 15744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_50
timestamp 1754861848
transform 1 0 14112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_51
timestamp 1754861848
transform 1 0 13728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_52
timestamp 1754861848
transform 1 0 16128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_53
timestamp 1754861848
transform 1 0 13440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_54
timestamp 1754861848
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_55
timestamp 1754861848
transform 1 0 15168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_56
timestamp 1754861848
transform 1 0 15456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_57
timestamp 1754861848
transform 1 0 12768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_58
timestamp 1754861848
transform 1 0 14496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_59
timestamp 1754861848
transform 1 0 15072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_60
timestamp 1754861848
transform 1 0 21312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_61
timestamp 1754861848
transform 1 0 21408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_62
timestamp 1754861848
transform 1 0 17088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_63
timestamp 1754861848
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_64
timestamp 1754861848
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_65
timestamp 1754861848
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_66
timestamp 1754861848
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_67
timestamp 1754861848
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_68
timestamp 1754861848
transform 1 0 18432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_69
timestamp 1754861848
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_70
timestamp 1754861848
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_71
timestamp 1754861848
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_72
timestamp 1754861848
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_73
timestamp 1754861848
transform 1 0 16800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_74
timestamp 1754861848
transform 1 0 12960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_75
timestamp 1754861848
transform 1 0 17184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_76
timestamp 1754861848
transform 1 0 16800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_77
timestamp 1754861848
transform 1 0 21312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_78
timestamp 1754861848
transform 1 0 20640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_79
timestamp 1754861848
transform 1 0 19968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_80
timestamp 1754861848
transform 1 0 19296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_81
timestamp 1754861848
transform 1 0 16800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_82
timestamp 1754861848
transform 1 0 11040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_83
timestamp 1754861848
transform 1 0 9408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_84
timestamp 1754861848
transform 1 0 10752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_85
timestamp 1754861848
transform 1 0 9696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_86
timestamp 1754861848
transform 1 0 11424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_87
timestamp 1754861848
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_88
timestamp 1754861848
transform 1 0 10752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_89
timestamp 1754861848
transform 1 0 10752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_90
timestamp 1754861848
transform 1 0 8064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_91
timestamp 1754861848
transform 1 0 11424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_92
timestamp 1754861848
transform 1 0 8736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_93
timestamp 1754861848
transform 1 0 9408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_94
timestamp 1754861848
transform 1 0 10080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_95
timestamp 1754861848
transform 1 0 8064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_96
timestamp 1754861848
transform 1 0 11712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_97
timestamp 1754861848
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_98
timestamp 1754861848
transform 1 0 10080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_99
timestamp 1754861848
transform 1 0 9408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_100
timestamp 1754861848
transform 1 0 8736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_101
timestamp 1754861848
transform 1 0 8064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_102
timestamp 1754861848
transform 1 0 10368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_103
timestamp 1754861848
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_104
timestamp 1754861848
transform 1 0 3360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_105
timestamp 1754861848
transform 1 0 6720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_106
timestamp 1754861848
transform 1 0 6048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_107
timestamp 1754861848
transform 1 0 4032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_108
timestamp 1754861848
transform 1 0 4032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_109
timestamp 1754861848
transform 1 0 3360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_110
timestamp 1754861848
transform 1 0 6720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_111
timestamp 1754861848
transform 1 0 3360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_112
timestamp 1754861848
transform 1 0 5376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_113
timestamp 1754861848
transform 1 0 4704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_114
timestamp 1754861848
transform 1 0 5856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_115
timestamp 1754861848
transform 1 0 4704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_116
timestamp 1754861848
transform 1 0 4032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_117
timestamp 1754861848
transform 1 0 6048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_118
timestamp 1754861848
transform 1 0 5376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_119
timestamp 1754861848
transform 1 0 4704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_120
timestamp 1754861848
transform 1 0 6720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_121
timestamp 1754861848
transform 1 0 5376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_122
timestamp 1754861848
transform 1 0 6048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_123
timestamp 1754861848
transform 1 0 4032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_124
timestamp 1754861848
transform 1 0 3360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_125
timestamp 1754861848
transform 1 0 3360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_126
timestamp 1754861848
transform 1 0 3360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_127
timestamp 1754861848
transform 1 0 3360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_128
timestamp 1754861848
transform 1 0 4032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_129
timestamp 1754861848
transform 1 0 7392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_130
timestamp 1754861848
transform 1 0 7392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_131
timestamp 1754861848
transform 1 0 3360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_132
timestamp 1754861848
transform 1 0 7392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_133
timestamp 1754861848
transform 1 0 3360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_134
timestamp 1754861848
transform 1 0 3360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_135
timestamp 1754861848
transform 1 0 3360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_136
timestamp 1754861848
transform 1 0 3360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_137
timestamp 1754861848
transform 1 0 3360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_138
timestamp 1754861848
transform 1 0 4032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_139
timestamp 1754861848
transform 1 0 6720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_140
timestamp 1754861848
transform 1 0 4032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_141
timestamp 1754861848
transform 1 0 5376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_142
timestamp 1754861848
transform 1 0 4032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_143
timestamp 1754861848
transform 1 0 5376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_144
timestamp 1754861848
transform 1 0 4032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_145
timestamp 1754861848
transform 1 0 4704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_146
timestamp 1754861848
transform 1 0 6048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_147
timestamp 1754861848
transform 1 0 3360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_148
timestamp 1754861848
transform 1 0 3360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_149
timestamp 1754861848
transform 1 0 5376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_150
timestamp 1754861848
transform 1 0 4704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_151
timestamp 1754861848
transform 1 0 3360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_152
timestamp 1754861848
transform 1 0 4704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_153
timestamp 1754861848
transform 1 0 6048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_154
timestamp 1754861848
transform 1 0 3360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_155
timestamp 1754861848
transform 1 0 4032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_156
timestamp 1754861848
transform 1 0 6048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_157
timestamp 1754861848
transform 1 0 4032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_158
timestamp 1754861848
transform 1 0 5376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_159
timestamp 1754861848
transform 1 0 4704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_160
timestamp 1754861848
transform 1 0 3360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_161
timestamp 1754861848
transform 1 0 4032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_162
timestamp 1754861848
transform 1 0 3360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_163
timestamp 1754861848
transform 1 0 4032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_164
timestamp 1754861848
transform 1 0 3360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_165
timestamp 1754861848
transform 1 0 18816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_166
timestamp 1754861848
transform 1 0 18528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_167
timestamp 1754861848
transform 1 0 19488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_168
timestamp 1754861848
transform 1 0 17856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_169
timestamp 1754861848
transform 1 0 21408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_170
timestamp 1754861848
transform 1 0 20064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_171
timestamp 1754861848
transform 1 0 20736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_172
timestamp 1754861848
transform 1 0 20064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_173
timestamp 1754861848
transform 1 0 19392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_174
timestamp 1754861848
transform 1 0 20160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_175
timestamp 1754861848
transform 1 0 18720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_176
timestamp 1754861848
transform 1 0 20064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_177
timestamp 1754861848
transform 1 0 20832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_178
timestamp 1754861848
transform 1 0 19392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_179
timestamp 1754861848
transform 1 0 20736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_180
timestamp 1754861848
transform 1 0 18720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_181
timestamp 1754861848
transform 1 0 20544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_182
timestamp 1754861848
transform 1 0 19200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_183
timestamp 1754861848
transform 1 0 21408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_184
timestamp 1754861848
transform 1 0 21216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_185
timestamp 1754861848
transform 1 0 21408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_186
timestamp 1754861848
transform 1 0 18048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_187
timestamp 1754861848
transform 1 0 19872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_188
timestamp 1754861848
transform 1 0 20736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_189
timestamp 1754861848
transform 1 0 18144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_190
timestamp 1754861848
transform 1 0 21024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_191
timestamp 1754861848
transform 1 0 20832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_192
timestamp 1754861848
transform 1 0 12096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_193
timestamp 1754861848
transform 1 0 12384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_194
timestamp 1754861848
transform 1 0 4032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_195
timestamp 1754861848
transform 1 0 21216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_196
timestamp 1754861848
transform 1 0 20544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_197
timestamp 1754861848
transform 1 0 3360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_198
timestamp 1754861848
transform 1 0 12096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_199
timestamp 1754861848
transform 1 0 3360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_200
timestamp 1754861848
transform 1 0 12096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  sg13g2_decap_8_201
timestamp 1754861848
transform 1 0 12480 0 1 6804
box -48 -56 720 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_0
timestamp 1754861848
transform 1 0 14208 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_1
timestamp 1754861848
transform 1 0 12864 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_2
timestamp 1754861848
transform 1 0 19488 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_3
timestamp 1754861848
transform 1 0 18144 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_4
timestamp 1754861848
transform 1 0 18528 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_5
timestamp 1754861848
transform 1 0 15456 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_6
timestamp 1754861848
transform 1 0 15456 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_7
timestamp 1754861848
transform 1 0 4320 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_8
timestamp 1754861848
transform 1 0 9696 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_9
timestamp 1754861848
transform 1 0 9888 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_10
timestamp 1754861848
transform 1 0 7680 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_11
timestamp 1754861848
transform 1 0 9888 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_12
timestamp 1754861848
transform 1 0 10080 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_13
timestamp 1754861848
transform 1 0 9888 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_14
timestamp 1754861848
transform 1 0 7680 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_15
timestamp 1754861848
transform 1 0 6816 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_16
timestamp 1754861848
transform 1 0 7392 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_17
timestamp 1754861848
transform 1 0 7392 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_18
timestamp 1754861848
transform 1 0 6720 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_19
timestamp 1754861848
transform 1 0 7488 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_20
timestamp 1754861848
transform 1 0 18816 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_21
timestamp 1754861848
transform 1 0 19392 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_22
timestamp 1754861848
transform 1 0 19008 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_23
timestamp 1754861848
transform 1 0 14688 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_24
timestamp 1754861848
transform 1 0 13440 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_25
timestamp 1754861848
transform 1 0 16992 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_26
timestamp 1754861848
transform 1 0 15360 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_27
timestamp 1754861848
transform 1 0 15552 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_28
timestamp 1754861848
transform 1 0 15168 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_29
timestamp 1754861848
transform 1 0 15264 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_30
timestamp 1754861848
transform 1 0 15264 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_31
timestamp 1754861848
transform 1 0 18432 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_32
timestamp 1754861848
transform 1 0 10176 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_33
timestamp 1754861848
transform 1 0 11328 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_34
timestamp 1754861848
transform 1 0 10656 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_35
timestamp 1754861848
transform 1 0 14688 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_36
timestamp 1754861848
transform 1 0 12672 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_37
timestamp 1754861848
transform 1 0 11616 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_38
timestamp 1754861848
transform 1 0 7392 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_39
timestamp 1754861848
transform 1 0 10944 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_40
timestamp 1754861848
transform 1 0 18240 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  sg13g2_dfrbpq_1_41
timestamp 1754861848
transform 1 0 11616 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_0
timestamp 1754861848
transform 1 0 15360 0 -1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_1
timestamp 1754861848
transform 1 0 4416 0 1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_2
timestamp 1754861848
transform 1 0 4416 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_3
timestamp 1754861848
transform 1 0 8832 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_4
timestamp 1754861848
transform 1 0 7872 0 1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_5
timestamp 1754861848
transform 1 0 6240 0 1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_6
timestamp 1754861848
transform 1 0 4800 0 1 14364
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_7
timestamp 1754861848
transform 1 0 7200 0 -1 14364
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_8
timestamp 1754861848
transform 1 0 5088 0 1 17388
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_9
timestamp 1754861848
transform 1 0 13056 0 -1 17388
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_10
timestamp 1754861848
transform 1 0 12288 0 -1 18900
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_11
timestamp 1754861848
transform 1 0 12672 0 -1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_12
timestamp 1754861848
transform 1 0 13056 0 1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_2  sg13g2_dfrbpq_2_13
timestamp 1754861848
transform 1 0 4704 0 1 12852
box -48 -56 2736 834
use sg13g2_fill_1  sg13g2_fill_1_0
timestamp 1754861848
transform 1 0 21984 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_1
timestamp 1754861848
transform 1 0 12768 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_2
timestamp 1754861848
transform 1 0 15456 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_3
timestamp 1754861848
transform 1 0 21984 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_4
timestamp 1754861848
transform 1 0 18432 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_5
timestamp 1754861848
transform 1 0 18624 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_6
timestamp 1754861848
transform 1 0 20064 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_7
timestamp 1754861848
transform 1 0 21984 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_8
timestamp 1754861848
transform 1 0 21984 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_9
timestamp 1754861848
transform 1 0 13824 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_10
timestamp 1754861848
transform 1 0 14400 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_11
timestamp 1754861848
transform 1 0 21984 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_12
timestamp 1754861848
transform 1 0 8736 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_13
timestamp 1754861848
transform 1 0 9216 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_14
timestamp 1754861848
transform 1 0 8064 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_15
timestamp 1754861848
transform 1 0 4320 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_16
timestamp 1754861848
transform 1 0 3744 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_17
timestamp 1754861848
transform 1 0 6816 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_18
timestamp 1754861848
transform 1 0 7872 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_19
timestamp 1754861848
transform 1 0 4224 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_20
timestamp 1754861848
transform 1 0 4416 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_21
timestamp 1754861848
transform 1 0 4224 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_22
timestamp 1754861848
transform 1 0 4224 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_23
timestamp 1754861848
transform 1 0 7104 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_24
timestamp 1754861848
transform 1 0 4896 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_25
timestamp 1754861848
transform 1 0 10176 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_26
timestamp 1754861848
transform 1 0 8256 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_27
timestamp 1754861848
transform 1 0 9984 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_28
timestamp 1754861848
transform 1 0 7776 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_29
timestamp 1754861848
transform 1 0 9888 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_30
timestamp 1754861848
transform 1 0 17856 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_31
timestamp 1754861848
transform 1 0 21984 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_32
timestamp 1754861848
transform 1 0 18336 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_33
timestamp 1754861848
transform 1 0 17952 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_34
timestamp 1754861848
transform 1 0 18144 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_35
timestamp 1754861848
transform 1 0 14592 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_36
timestamp 1754861848
transform 1 0 14976 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_37
timestamp 1754861848
transform 1 0 13056 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_38
timestamp 1754861848
transform 1 0 14208 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_39
timestamp 1754861848
transform 1 0 13536 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_40
timestamp 1754861848
transform 1 0 14592 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_41
timestamp 1754861848
transform 1 0 16896 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_42
timestamp 1754861848
transform 1 0 19776 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_43
timestamp 1754861848
transform 1 0 4224 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_44
timestamp 1754861848
transform 1 0 21984 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  sg13g2_fill_1_45
timestamp 1754861848
transform 1 0 9984 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  sg13g2_fill_2_0
timestamp 1754861848
transform 1 0 21888 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_1
timestamp 1754861848
transform 1 0 21888 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_2
timestamp 1754861848
transform 1 0 21792 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_3
timestamp 1754861848
transform 1 0 21888 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_4
timestamp 1754861848
transform 1 0 21888 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_5
timestamp 1754861848
transform 1 0 18432 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_6
timestamp 1754861848
transform 1 0 21792 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_7
timestamp 1754861848
transform 1 0 13632 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_8
timestamp 1754861848
transform 1 0 21792 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_9
timestamp 1754861848
transform 1 0 13056 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_10
timestamp 1754861848
transform 1 0 14208 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_11
timestamp 1754861848
transform 1 0 8544 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_12
timestamp 1754861848
transform 1 0 3744 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_13
timestamp 1754861848
transform 1 0 4608 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_14
timestamp 1754861848
transform 1 0 6624 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_15
timestamp 1754861848
transform 1 0 4032 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_16
timestamp 1754861848
transform 1 0 9984 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_17
timestamp 1754861848
transform 1 0 7872 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_18
timestamp 1754861848
transform 1 0 7872 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_19
timestamp 1754861848
transform 1 0 12000 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_20
timestamp 1754861848
transform 1 0 9024 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_21
timestamp 1754861848
transform 1 0 6432 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_22
timestamp 1754861848
transform 1 0 4032 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_23
timestamp 1754861848
transform 1 0 9888 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_24
timestamp 1754861848
transform 1 0 5952 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_25
timestamp 1754861848
transform 1 0 4704 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_26
timestamp 1754861848
transform 1 0 4032 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_27
timestamp 1754861848
transform 1 0 7776 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_28
timestamp 1754861848
transform 1 0 5088 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_29
timestamp 1754861848
transform 1 0 5664 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_30
timestamp 1754861848
transform 1 0 12480 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_31
timestamp 1754861848
transform 1 0 9984 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_32
timestamp 1754861848
transform 1 0 10752 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_33
timestamp 1754861848
transform 1 0 11424 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_34
timestamp 1754861848
transform 1 0 6048 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_35
timestamp 1754861848
transform 1 0 19200 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_36
timestamp 1754861848
transform 1 0 21888 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_37
timestamp 1754861848
transform 1 0 17664 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_38
timestamp 1754861848
transform 1 0 21888 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_39
timestamp 1754861848
transform 1 0 17856 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_40
timestamp 1754861848
transform 1 0 15264 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_41
timestamp 1754861848
transform 1 0 17568 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_42
timestamp 1754861848
transform 1 0 21888 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_43
timestamp 1754861848
transform 1 0 19584 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_44
timestamp 1754861848
transform 1 0 21888 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_45
timestamp 1754861848
transform 1 0 21888 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_46
timestamp 1754861848
transform 1 0 21888 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_47
timestamp 1754861848
transform 1 0 4704 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_48
timestamp 1754861848
transform 1 0 10368 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_49
timestamp 1754861848
transform 1 0 11520 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  sg13g2_fill_2_50
timestamp 1754861848
transform 1 0 4032 0 1 12852
box -48 -56 240 834
use sg13g2_inv_1  sg13g2_inv_1_0
timestamp 1754861848
transform 1 0 19200 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_1
timestamp 1754861848
transform 1 0 21024 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_2
timestamp 1754861848
transform 1 0 21120 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_3
timestamp 1754861848
transform 1 0 20736 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_4
timestamp 1754861848
transform 1 0 12192 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_5
timestamp 1754861848
transform 1 0 3936 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_6
timestamp 1754861848
transform 1 0 10272 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_7
timestamp 1754861848
transform 1 0 8256 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_8
timestamp 1754861848
transform 1 0 11328 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_9
timestamp 1754861848
transform 1 0 4320 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_10
timestamp 1754861848
transform 1 0 21408 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_11
timestamp 1754861848
transform 1 0 21600 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_12
timestamp 1754861848
transform 1 0 12960 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_13
timestamp 1754861848
transform 1 0 13152 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_14
timestamp 1754861848
transform 1 0 17760 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_15
timestamp 1754861848
transform 1 0 19776 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_16
timestamp 1754861848
transform 1 0 19296 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_17
timestamp 1754861848
transform 1 0 20544 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_18
timestamp 1754861848
transform 1 0 15648 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_19
timestamp 1754861848
transform 1 0 15936 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  sg13g2_inv_1_20
timestamp 1754861848
transform 1 0 20256 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_2  sg13g2_inv_2_0
timestamp 1754861848
transform 1 0 12192 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_2  sg13g2_inv_2_1
timestamp 1754861848
transform 1 0 4704 0 -1 17388
box -48 -56 432 834
use sg13g2_mux2_1  sg13g2_mux2_1_0
timestamp 1754861848
transform 1 0 14496 0 1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_1
timestamp 1754861848
transform 1 0 13248 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_2
timestamp 1754861848
transform 1 0 18720 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_3
timestamp 1754861848
transform 1 0 13248 0 1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_4
timestamp 1754861848
transform 1 0 14496 0 1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_5
timestamp 1754861848
transform 1 0 17184 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_6
timestamp 1754861848
transform 1 0 5088 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_7
timestamp 1754861848
transform 1 0 5664 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_8
timestamp 1754861848
transform 1 0 6912 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_9
timestamp 1754861848
transform 1 0 8928 0 1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_10
timestamp 1754861848
transform 1 0 11328 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_11
timestamp 1754861848
transform 1 0 8736 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_12
timestamp 1754861848
transform 1 0 8928 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_13
timestamp 1754861848
transform 1 0 6336 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_14
timestamp 1754861848
transform 1 0 6144 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_15
timestamp 1754861848
transform 1 0 4992 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_16
timestamp 1754861848
transform 1 0 5760 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_17
timestamp 1754861848
transform 1 0 5856 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_18
timestamp 1754861848
transform 1 0 6432 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_19
timestamp 1754861848
transform 1 0 6720 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_20
timestamp 1754861848
transform 1 0 10656 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_21
timestamp 1754861848
transform 1 0 11328 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_22
timestamp 1754861848
transform 1 0 9696 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_23
timestamp 1754861848
transform 1 0 9792 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_24
timestamp 1754861848
transform 1 0 8736 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_25
timestamp 1754861848
transform 1 0 7296 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_26
timestamp 1754861848
transform 1 0 5088 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_27
timestamp 1754861848
transform 1 0 10848 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_28
timestamp 1754861848
transform 1 0 18240 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_29
timestamp 1754861848
transform 1 0 18048 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_30
timestamp 1754861848
transform 1 0 18048 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_31
timestamp 1754861848
transform 1 0 14016 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_32
timestamp 1754861848
transform 1 0 14592 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_33
timestamp 1754861848
transform 1 0 13248 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_34
timestamp 1754861848
transform 1 0 14304 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_35
timestamp 1754861848
transform 1 0 14208 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_36
timestamp 1754861848
transform 1 0 17952 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_37
timestamp 1754861848
transform 1 0 19584 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_38
timestamp 1754861848
transform 1 0 13632 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_39
timestamp 1754861848
transform 1 0 16224 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_40
timestamp 1754861848
transform 1 0 14688 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_41
timestamp 1754861848
transform 1 0 6624 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_42
timestamp 1754861848
transform 1 0 12000 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_43
timestamp 1754861848
transform 1 0 17664 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_44
timestamp 1754861848
transform 1 0 12480 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_45
timestamp 1754861848
transform 1 0 4896 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_46
timestamp 1754861848
transform 1 0 12288 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_47
timestamp 1754861848
transform 1 0 12096 0 1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_48
timestamp 1754861848
transform 1 0 12096 0 1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  sg13g2_mux2_1_49
timestamp 1754861848
transform 1 0 10560 0 1 12852
box -48 -56 1008 834
use sg13g2_mux4_1  sg13g2_mux4_1_0
timestamp 1754861848
transform 1 0 15552 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_1
timestamp 1754861848
transform 1 0 9312 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_2
timestamp 1754861848
transform 1 0 7872 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_3
timestamp 1754861848
transform 1 0 15456 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_4
timestamp 1754861848
transform 1 0 15456 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_5
timestamp 1754861848
transform 1 0 8352 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_6
timestamp 1754861848
transform 1 0 15744 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  sg13g2_mux4_1_7
timestamp 1754861848
transform 1 0 12000 0 1 18900
box -48 -56 2064 834
use sg13g2_nand2_1  sg13g2_nand2_1_0
timestamp 1754861848
transform 1 0 8160 0 -1 6804
box -48 -56 432 834
use sg13g2_nand2_1  sg13g2_nand2_1_1
timestamp 1754861848
transform 1 0 8832 0 -1 6804
box -48 -56 432 834
use sg13g2_nand2_1  sg13g2_nand2_1_2
timestamp 1754861848
transform 1 0 5472 0 -1 6804
box -48 -56 432 834
use sg13g2_nand2_1  sg13g2_nand2_1_3
timestamp 1754861848
transform 1 0 4320 0 1 8316
box -48 -56 432 834
use sg13g2_nand2_2  sg13g2_nand2_2_0
timestamp 1754861848
transform 1 0 7296 0 -1 6804
box -48 -56 624 834
use sg13g2_nand2b_1  sg13g2_nand2b_1_0
timestamp 1754861848
transform 1 0 6048 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  sg13g2_nand2b_1_1
timestamp 1754861848
transform 1 0 8544 0 1 8316
box -48 -56 528 834
use sg13g2_nand2b_2  sg13g2_nand2b_2_0
timestamp 1754861848
transform 1 0 6912 0 1 9828
box -48 -56 816 834
use sg13g2_nand2b_2  sg13g2_nand2b_2_1
timestamp 1754861848
transform 1 0 6624 0 1 8316
box -48 -56 816 834
use sg13g2_nand3b_1  sg13g2_nand3b_1_0
timestamp 1754861848
transform 1 0 4800 0 -1 6804
box -48 -56 720 834
use sg13g2_nand3b_1  sg13g2_nand3b_1_1
timestamp 1754861848
transform 1 0 5184 0 1 8316
box -48 -56 720 834
use sg13g2_nor2_1  sg13g2_nor2_1_0
timestamp 1754861848
transform 1 0 9312 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  sg13g2_nor2_1_1
timestamp 1754861848
transform 1 0 6912 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  sg13g2_nor2_1_2
timestamp 1754861848
transform 1 0 7968 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_0
timestamp 1754861848
transform 1 0 18336 0 -1 9828
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_1
timestamp 1754861848
transform 1 0 9216 0 1 8316
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_2
timestamp 1754861848
transform 1 0 9984 0 1 17388
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_3
timestamp 1754861848
transform 1 0 10464 0 1 17388
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_4
timestamp 1754861848
transform 1 0 14784 0 1 18900
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_5
timestamp 1754861848
transform 1 0 17472 0 -1 14364
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_6
timestamp 1754861848
transform 1 0 17472 0 1 18900
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_7
timestamp 1754861848
transform 1 0 17760 0 1 12852
box -54 -56 528 834
use sg13g2_nor2b_1  sg13g2_nor2b_1_8
timestamp 1754861848
transform 1 0 10080 0 1 12852
box -54 -56 528 834
use sg13g2_nor3_1  sg13g2_nor3_1_0
timestamp 1754861848
transform 1 0 4704 0 1 8316
box -48 -56 528 834
use sg13g2_nor4_2  sg13g2_nor4_2_0
timestamp 1754861848
transform 1 0 6528 0 -1 9828
box -48 -56 1200 834
use sg13g2_nor4_2  sg13g2_nor4_2_1
timestamp 1754861848
transform 1 0 7680 0 -1 9828
box -48 -56 1200 834
use sg13g2_nor4_2  sg13g2_nor4_2_2
timestamp 1754861848
transform 1 0 7392 0 1 8316
box -48 -56 1200 834
use sg13g2_tiehi  sg13g2_tiehi_0
timestamp 1754861848
transform 1 0 18816 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_1
timestamp 1754861848
transform 1 0 19680 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_2
timestamp 1754861848
transform 1 0 21408 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_3
timestamp 1754861848
transform 1 0 18048 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_4
timestamp 1754861848
transform 1 0 4512 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_5
timestamp 1754861848
transform 1 0 5280 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_6
timestamp 1754861848
transform 1 0 5472 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_7
timestamp 1754861848
transform 1 0 8352 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_8
timestamp 1754861848
transform 1 0 8832 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_9
timestamp 1754861848
transform 1 0 8544 0 -1 15876
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_10
timestamp 1754861848
transform 1 0 4416 0 1 14364
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_11
timestamp 1754861848
transform 1 0 5280 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_12
timestamp 1754861848
transform 1 0 10272 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_13
timestamp 1754861848
transform 1 0 10944 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_14
timestamp 1754861848
transform 1 0 10656 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_15
timestamp 1754861848
transform 1 0 10272 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_16
timestamp 1754861848
transform 1 0 18432 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_17
timestamp 1754861848
transform 1 0 21504 0 1 14364
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_18
timestamp 1754861848
transform 1 0 14208 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_19
timestamp 1754861848
transform 1 0 14976 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_20
timestamp 1754861848
transform 1 0 18912 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_21
timestamp 1754861848
transform 1 0 17952 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_22
timestamp 1754861848
transform 1 0 15744 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_23
timestamp 1754861848
transform 1 0 12576 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_24
timestamp 1754861848
transform 1 0 6240 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_25
timestamp 1754861848
transform 1 0 4320 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  sg13g2_tiehi_26
timestamp 1754861848
transform 1 0 20832 0 1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  sg13g2_xnor2_1_0
timestamp 1754861848
transform 1 0 7104 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  sg13g2_xnor2_1_1
timestamp 1754861848
transform 1 0 8064 0 -1 8316
box -48 -56 816 834
use spi_DEF_FILL  spi_DEF_FILL_0
timestamp 1754861848
transform 1 0 0 0 1 0
box 3360 3780 21984 21836
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_0
timestamp 1754861848
transform 1 0 21200 0 1 5292
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_1
timestamp 1754861848
transform 1 0 21200 0 1 3780
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_2
timestamp 1754861848
transform 1 0 13640 0 1 4536
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_3
timestamp 1754861848
transform 1 0 13640 0 1 6048
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_4
timestamp 1754861848
transform 1 0 13640 0 1 7560
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_5
timestamp 1754861848
transform 1 0 13640 0 1 9072
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_6
timestamp 1754861848
transform 1 0 13640 0 1 10584
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_7
timestamp 1754861848
transform 1 0 13640 0 1 12096
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_8
timestamp 1754861848
transform 1 0 21200 0 1 6804
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_9
timestamp 1754861848
transform 1 0 21200 0 1 8316
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_10
timestamp 1754861848
transform 1 0 21200 0 1 11340
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_11
timestamp 1754861848
transform 1 0 21200 0 1 9828
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_12
timestamp 1754861848
transform 1 0 6080 0 1 3780
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_13
timestamp 1754861848
transform 1 0 6080 0 1 5292
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_14
timestamp 1754861848
transform 1 0 6080 0 1 6804
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_15
timestamp 1754861848
transform 1 0 6080 0 1 8316
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_16
timestamp 1754861848
transform 1 0 6080 0 1 9828
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_17
timestamp 1754861848
transform 1 0 6080 0 1 11340
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_18
timestamp 1754861848
transform 1 0 6080 0 1 15876
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_19
timestamp 1754861848
transform 1 0 6080 0 1 14364
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_20
timestamp 1754861848
transform 1 0 6080 0 1 18900
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_21
timestamp 1754861848
transform 1 0 6080 0 1 17388
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_22
timestamp 1754861848
transform 1 0 6080 0 1 21924
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_23
timestamp 1754861848
transform 1 0 6080 0 1 20412
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_24
timestamp 1754861848
transform 1 0 21200 0 1 15876
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_25
timestamp 1754861848
transform 1 0 21200 0 1 14364
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_26
timestamp 1754861848
transform 1 0 21200 0 1 17388
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_27
timestamp 1754861848
transform 1 0 21200 0 1 18900
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_28
timestamp 1754861848
transform 1 0 13640 0 1 15120
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_29
timestamp 1754861848
transform 1 0 13640 0 1 13608
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_30
timestamp 1754861848
transform 1 0 13640 0 1 18144
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_31
timestamp 1754861848
transform 1 0 13640 0 1 16632
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_32
timestamp 1754861848
transform 1 0 13640 0 1 21168
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_33
timestamp 1754861848
transform 1 0 13640 0 1 19656
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_34
timestamp 1754861848
transform 1 0 21200 0 1 21924
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_35
timestamp 1754861848
transform 1 0 21200 0 1 20412
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_36
timestamp 1754861848
transform 1 0 6080 0 1 12852
box -193 -44 193 44
use VIA_via1_2_2200_440_1_5_410_410  VIA_via1_2_2200_440_1_5_410_410_37
timestamp 1754861848
transform 1 0 21200 0 1 12852
box -193 -44 193 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_0
timestamp 1754861848
transform 1 0 24880 0 1 4536
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_1
timestamp 1754861848
transform 1 0 23480 0 1 5292
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_2
timestamp 1754861848
transform 1 0 23480 0 1 3780
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_3
timestamp 1754861848
transform 1 0 24880 0 1 6048
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_4
timestamp 1754861848
transform 1 0 24880 0 1 9072
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_5
timestamp 1754861848
transform 1 0 23480 0 1 6804
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_6
timestamp 1754861848
transform 1 0 24880 0 1 7560
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_7
timestamp 1754861848
transform 1 0 23480 0 1 8316
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_8
timestamp 1754861848
transform 1 0 23480 0 1 11340
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_9
timestamp 1754861848
transform 1 0 23480 0 1 9828
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_10
timestamp 1754861848
transform 1 0 24880 0 1 10584
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_11
timestamp 1754861848
transform 1 0 24880 0 1 12096
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_12
timestamp 1754861848
transform 1 0 560 0 1 6048
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_13
timestamp 1754861848
transform 1 0 1960 0 1 5292
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_14
timestamp 1754861848
transform 1 0 1960 0 1 3780
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_15
timestamp 1754861848
transform 1 0 560 0 1 4536
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_16
timestamp 1754861848
transform 1 0 1960 0 1 8316
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_17
timestamp 1754861848
transform 1 0 1960 0 1 6804
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_18
timestamp 1754861848
transform 1 0 560 0 1 7560
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_19
timestamp 1754861848
transform 1 0 560 0 1 9072
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_20
timestamp 1754861848
transform 1 0 560 0 1 12096
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_21
timestamp 1754861848
transform 1 0 1960 0 1 11340
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_22
timestamp 1754861848
transform 1 0 1960 0 1 9828
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_23
timestamp 1754861848
transform 1 0 560 0 1 10584
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_24
timestamp 1754861848
transform 1 0 1960 0 1 14364
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_25
timestamp 1754861848
transform 1 0 560 0 1 15120
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_26
timestamp 1754861848
transform 1 0 1960 0 1 15876
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_27
timestamp 1754861848
transform 1 0 560 0 1 13608
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_28
timestamp 1754861848
transform 1 0 1960 0 1 17388
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_29
timestamp 1754861848
transform 1 0 560 0 1 16632
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_30
timestamp 1754861848
transform 1 0 560 0 1 18144
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_31
timestamp 1754861848
transform 1 0 1960 0 1 18900
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_32
timestamp 1754861848
transform 1 0 1960 0 1 21924
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_33
timestamp 1754861848
transform 1 0 1960 0 1 20412
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_34
timestamp 1754861848
transform 1 0 560 0 1 19656
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_35
timestamp 1754861848
transform 1 0 560 0 1 21168
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_36
timestamp 1754861848
transform 1 0 24880 0 1 13608
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_37
timestamp 1754861848
transform 1 0 24880 0 1 15120
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_38
timestamp 1754861848
transform 1 0 23480 0 1 15876
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_39
timestamp 1754861848
transform 1 0 23480 0 1 14364
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_40
timestamp 1754861848
transform 1 0 24880 0 1 18144
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_41
timestamp 1754861848
transform 1 0 23480 0 1 17388
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_42
timestamp 1754861848
transform 1 0 24880 0 1 16632
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_43
timestamp 1754861848
transform 1 0 23480 0 1 18900
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_44
timestamp 1754861848
transform 1 0 24880 0 1 21168
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_45
timestamp 1754861848
transform 1 0 23480 0 1 21924
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_46
timestamp 1754861848
transform 1 0 23480 0 1 20412
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_47
timestamp 1754861848
transform 1 0 24880 0 1 19656
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_48
timestamp 1754861848
transform 1 0 1960 0 1 12852
box -480 -44 480 44
use VIA_via1_2_5000_440_1_12_410_410  VIA_via1_2_5000_440_1_12_410_410_49
timestamp 1754861848
transform 1 0 23480 0 1 12852
box -480 -44 480 44
use VIA_Via1_XY  VIA_Via1_XY_0
timestamp 1754861848
transform 1 0 18732 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_1
timestamp 1754861848
transform 1 0 15960 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_2
timestamp 1754861848
transform 1 0 16800 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_3
timestamp 1754861848
transform 1 0 18228 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_4
timestamp 1754861848
transform 1 0 16338 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_5
timestamp 1754861848
transform 1 0 18144 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_6
timestamp 1754861848
transform 1 0 18648 0 1 9696
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_7
timestamp 1754861848
transform 1 0 16800 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_8
timestamp 1754861848
transform 1 0 18438 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_9
timestamp 1754861848
transform 1 0 17304 0 1 9495
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_10
timestamp 1754861848
transform 1 0 18396 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_11
timestamp 1754861848
transform 1 0 13356 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_12
timestamp 1754861848
transform 1 0 13608 0 1 8544
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_13
timestamp 1754861848
transform 1 0 14028 0 1 7920
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_14
timestamp 1754861848
transform 1 0 14112 0 1 8928
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_15
timestamp 1754861848
transform 1 0 14868 0 1 8544
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_16
timestamp 1754861848
transform 1 0 15372 0 1 9216
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_17
timestamp 1754861848
transform 1 0 14196 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_18
timestamp 1754861848
transform 1 0 14784 0 1 7920
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_19
timestamp 1754861848
transform 1 0 15540 0 1 8544
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_20
timestamp 1754861848
transform 1 0 13440 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_21
timestamp 1754861848
transform 1 0 14658 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_22
timestamp 1754861848
transform 1 0 14952 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_23
timestamp 1754861848
transform 1 0 14112 0 1 10368
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_24
timestamp 1754861848
transform 1 0 15204 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_25
timestamp 1754861848
transform 1 0 13146 0 1 10992
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_26
timestamp 1754861848
transform 1 0 13440 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_27
timestamp 1754861848
transform 1 0 14952 0 1 11703
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_28
timestamp 1754861848
transform 1 0 14868 0 1 11563
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_29
timestamp 1754861848
transform 1 0 14532 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_30
timestamp 1754861848
transform 1 0 13608 0 1 10051
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_31
timestamp 1754861848
transform 1 0 14700 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_32
timestamp 1754861848
transform 1 0 15540 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_33
timestamp 1754861848
transform 1 0 14028 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_34
timestamp 1754861848
transform 1 0 14658 0 1 11661
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_35
timestamp 1754861848
transform 1 0 15540 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_36
timestamp 1754861848
transform 1 0 12768 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_37
timestamp 1754861848
transform 1 0 15372 0 1 11808
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_38
timestamp 1754861848
transform 1 0 17856 0 1 12528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_39
timestamp 1754861848
transform 1 0 16716 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_40
timestamp 1754861848
transform 1 0 17556 0 1 10051
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_41
timestamp 1754861848
transform 1 0 18900 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_42
timestamp 1754861848
transform 1 0 18984 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_43
timestamp 1754861848
transform 1 0 17340 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_44
timestamp 1754861848
transform 1 0 15960 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_45
timestamp 1754861848
transform 1 0 18648 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_46
timestamp 1754861848
transform 1 0 18060 0 1 10272
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_47
timestamp 1754861848
transform 1 0 18144 0 1 10944
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_48
timestamp 1754861848
transform 1 0 17640 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_49
timestamp 1754861848
transform 1 0 16716 0 1 9984
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_50
timestamp 1754861848
transform 1 0 18228 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_51
timestamp 1754861848
transform 1 0 16044 0 1 12528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_52
timestamp 1754861848
transform 1 0 15876 0 1 11017
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_53
timestamp 1754861848
transform 1 0 19992 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_54
timestamp 1754861848
transform 1 0 20832 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_55
timestamp 1754861848
transform 1 0 19572 0 1 9600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_56
timestamp 1754861848
transform 1 0 19572 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_57
timestamp 1754861848
transform 1 0 19488 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_58
timestamp 1754861848
transform 1 0 19194 0 1 10977
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_59
timestamp 1754861848
transform 1 0 20328 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_60
timestamp 1754861848
transform 1 0 20832 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_61
timestamp 1754861848
transform 1 0 7476 0 1 6432
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_62
timestamp 1754861848
transform 1 0 8400 0 1 6576
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_63
timestamp 1754861848
transform 1 0 9072 0 1 6576
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_64
timestamp 1754861848
transform 1 0 7728 0 1 6432
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_65
timestamp 1754861848
transform 1 0 9576 0 1 6336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_66
timestamp 1754861848
transform 1 0 4032 0 1 6455
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_67
timestamp 1754861848
transform 1 0 5208 0 1 6432
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_68
timestamp 1754861848
transform 1 0 5376 0 1 6336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_69
timestamp 1754861848
transform 1 0 5712 0 1 6576
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_70
timestamp 1754861848
transform 1 0 5244 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_71
timestamp 1754861848
transform 1 0 5460 0 1 9600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_72
timestamp 1754861848
transform 1 0 5574 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_73
timestamp 1754861848
transform 1 0 6048 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_74
timestamp 1754861848
transform 1 0 5544 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_75
timestamp 1754861848
transform 1 0 6132 0 1 9501
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_76
timestamp 1754861848
transform 1 0 4956 0 1 8832
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_77
timestamp 1754861848
transform 1 0 6244 0 1 8544
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_78
timestamp 1754861848
transform 1 0 4788 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_79
timestamp 1754861848
transform 1 0 5052 0 1 12528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_80
timestamp 1754861848
transform 1 0 6132 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_81
timestamp 1754861848
transform 1 0 6216 0 1 11117
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_82
timestamp 1754861848
transform 1 0 5754 0 1 11904
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_83
timestamp 1754861848
transform 1 0 4410 0 1 10080
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_84
timestamp 1754861848
transform 1 0 5856 0 1 10992
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_85
timestamp 1754861848
transform 1 0 5292 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_86
timestamp 1754861848
transform 1 0 12264 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_87
timestamp 1754861848
transform 1 0 11424 0 1 7008
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_88
timestamp 1754861848
transform 1 0 11508 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_89
timestamp 1754861848
transform 1 0 9595 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_90
timestamp 1754861848
transform 1 0 9828 0 1 8592
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_91
timestamp 1754861848
transform 1 0 10206 0 1 8603
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_92
timestamp 1754861848
transform 1 0 9912 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_93
timestamp 1754861848
transform 1 0 10752 0 1 7104
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_94
timestamp 1754861848
transform 1 0 12558 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_95
timestamp 1754861848
transform 1 0 10164 0 1 7968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_96
timestamp 1754861848
transform 1 0 12684 0 1 9216
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_97
timestamp 1754861848
transform 1 0 11928 0 1 7776
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_98
timestamp 1754861848
transform 1 0 11718 0 1 7968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_99
timestamp 1754861848
transform 1 0 10668 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_100
timestamp 1754861848
transform 1 0 10416 0 1 7126
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_101
timestamp 1754861848
transform 1 0 6972 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_102
timestamp 1754861848
transform 1 0 8106 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_103
timestamp 1754861848
transform 1 0 7392 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_104
timestamp 1754861848
transform 1 0 6972 0 1 7152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_105
timestamp 1754861848
transform 1 0 7560 0 1 7248
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_106
timestamp 1754861848
transform 1 0 8232 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_107
timestamp 1754861848
transform 1 0 7812 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_108
timestamp 1754861848
transform 1 0 6720 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_109
timestamp 1754861848
transform 1 0 7896 0 1 8688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_110
timestamp 1754861848
transform 1 0 7224 0 1 7968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_111
timestamp 1754861848
transform 1 0 7560 0 1 8649
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_112
timestamp 1754861848
transform 1 0 7224 0 1 9495
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_113
timestamp 1754861848
transform 1 0 8568 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_114
timestamp 1754861848
transform 1 0 9324 0 1 7968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_115
timestamp 1754861848
transform 1 0 8484 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_116
timestamp 1754861848
transform 1 0 8736 0 1 7872
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_117
timestamp 1754861848
transform 1 0 6972 0 1 7968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_118
timestamp 1754861848
transform 1 0 7560 0 1 9504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_119
timestamp 1754861848
transform 1 0 9324 0 1 8640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_120
timestamp 1754861848
transform 1 0 8106 0 1 9456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_121
timestamp 1754861848
transform 1 0 8232 0 1 10848
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_122
timestamp 1754861848
transform 1 0 9030 0 1 12528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_123
timestamp 1754861848
transform 1 0 6720 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_124
timestamp 1754861848
transform 1 0 7086 0 1 10992
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_125
timestamp 1754861848
transform 1 0 7560 0 1 11616
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_126
timestamp 1754861848
transform 1 0 7770 0 1 10128
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_127
timestamp 1754861848
transform 1 0 7392 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_128
timestamp 1754861848
transform 1 0 6804 0 1 9984
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_129
timestamp 1754861848
transform 1 0 6972 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_130
timestamp 1754861848
transform 1 0 8148 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_131
timestamp 1754861848
transform 1 0 6804 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_132
timestamp 1754861848
transform 1 0 8636 0 1 12489
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_133
timestamp 1754861848
transform 1 0 9198 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_134
timestamp 1754861848
transform 1 0 8148 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_135
timestamp 1754861848
transform 1 0 9102 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_136
timestamp 1754861848
transform 1 0 8904 0 1 11040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_137
timestamp 1754861848
transform 1 0 7308 0 1 10272
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_138
timestamp 1754861848
transform 1 0 7098 0 1 12551
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_139
timestamp 1754861848
transform 1 0 11172 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_140
timestamp 1754861848
transform 1 0 11802 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_141
timestamp 1754861848
transform 1 0 12684 0 1 12505
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_142
timestamp 1754861848
transform 1 0 10374 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_143
timestamp 1754861848
transform 1 0 12390 0 1 11520
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_144
timestamp 1754861848
transform 1 0 10164 0 1 9984
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_145
timestamp 1754861848
transform 1 0 11508 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_146
timestamp 1754861848
transform 1 0 12180 0 1 10464
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_147
timestamp 1754861848
transform 1 0 11256 0 1 11664
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_148
timestamp 1754861848
transform 1 0 11844 0 1 10051
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_149
timestamp 1754861848
transform 1 0 11844 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_150
timestamp 1754861848
transform 1 0 9786 0 1 10992
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_151
timestamp 1754861848
transform 1 0 10332 0 1 11712
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_152
timestamp 1754861848
transform 1 0 12180 0 1 11136
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_153
timestamp 1754861848
transform 1 0 9599 0 1 12480
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_154
timestamp 1754861848
transform 1 0 12444 0 1 10176
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_155
timestamp 1754861848
transform 1 0 10164 0 1 11017
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_156
timestamp 1754861848
transform 1 0 11256 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_157
timestamp 1754861848
transform 1 0 12474 0 1 14064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_158
timestamp 1754861848
transform 1 0 10836 0 1 13920
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_159
timestamp 1754861848
transform 1 0 11004 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_160
timestamp 1754861848
transform 1 0 12180 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_161
timestamp 1754861848
transform 1 0 10458 0 1 13344
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_162
timestamp 1754861848
transform 1 0 12558 0 1 13184
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_163
timestamp 1754861848
transform 1 0 10920 0 1 13075
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_164
timestamp 1754861848
transform 1 0 12264 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_165
timestamp 1754861848
transform 1 0 10164 0 1 13173
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_166
timestamp 1754861848
transform 1 0 10752 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_167
timestamp 1754861848
transform 1 0 11424 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_168
timestamp 1754861848
transform 1 0 11424 0 1 13344
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_169
timestamp 1754861848
transform 1 0 10584 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_170
timestamp 1754861848
transform 1 0 10164 0 1 14592
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_171
timestamp 1754861848
transform 1 0 12672 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_172
timestamp 1754861848
transform 1 0 9954 0 1 15648
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_173
timestamp 1754861848
transform 1 0 9744 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_174
timestamp 1754861848
transform 1 0 10332 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_175
timestamp 1754861848
transform 1 0 12558 0 1 13075
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_176
timestamp 1754861848
transform 1 0 9996 0 1 14976
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_177
timestamp 1754861848
transform 1 0 6804 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_178
timestamp 1754861848
transform 1 0 6720 0 1 15653
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_179
timestamp 1754861848
transform 1 0 7476 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_180
timestamp 1754861848
transform 1 0 9120 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_181
timestamp 1754861848
transform 1 0 8820 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_182
timestamp 1754861848
transform 1 0 8358 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_183
timestamp 1754861848
transform 1 0 7896 0 1 13224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_184
timestamp 1754861848
transform 1 0 8736 0 1 13177
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_185
timestamp 1754861848
transform 1 0 7308 0 1 14976
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_186
timestamp 1754861848
transform 1 0 7980 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_187
timestamp 1754861848
transform 1 0 6594 0 1 14064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_188
timestamp 1754861848
transform 1 0 6492 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_189
timestamp 1754861848
transform 1 0 7770 0 1 15575
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_190
timestamp 1754861848
transform 1 0 7224 0 1 15264
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_191
timestamp 1754861848
transform 1 0 9492 0 1 15648
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_192
timestamp 1754861848
transform 1 0 7476 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_193
timestamp 1754861848
transform 1 0 9324 0 1 18336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_194
timestamp 1754861848
transform 1 0 8652 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_195
timestamp 1754861848
transform 1 0 9114 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_196
timestamp 1754861848
transform 1 0 8148 0 1 18576
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_197
timestamp 1754861848
transform 1 0 7476 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_198
timestamp 1754861848
transform 1 0 8736 0 1 17040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_199
timestamp 1754861848
transform 1 0 7644 0 1 17710
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_200
timestamp 1754861848
transform 1 0 9492 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_201
timestamp 1754861848
transform 1 0 6804 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_202
timestamp 1754861848
transform 1 0 7224 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_203
timestamp 1754861848
transform 1 0 7224 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_204
timestamp 1754861848
transform 1 0 8064 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_205
timestamp 1754861848
transform 1 0 6720 0 1 18432
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_206
timestamp 1754861848
transform 1 0 7308 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_207
timestamp 1754861848
transform 1 0 7896 0 1 17016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_208
timestamp 1754861848
transform 1 0 6636 0 1 16320
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_209
timestamp 1754861848
transform 1 0 8548 0 1 17808
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_210
timestamp 1754861848
transform 1 0 10164 0 1 18672
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_211
timestamp 1754861848
transform 1 0 9966 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_212
timestamp 1754861848
transform 1 0 11802 0 1 18599
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_213
timestamp 1754861848
transform 1 0 10836 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_214
timestamp 1754861848
transform 1 0 11298 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_215
timestamp 1754861848
transform 1 0 10668 0 1 18336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_216
timestamp 1754861848
transform 1 0 11508 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_217
timestamp 1754861848
transform 1 0 11424 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_218
timestamp 1754861848
transform 1 0 12264 0 1 17735
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_219
timestamp 1754861848
transform 1 0 11424 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_220
timestamp 1754861848
transform 1 0 11004 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_221
timestamp 1754861848
transform 1 0 9596 0 1 16239
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_222
timestamp 1754861848
transform 1 0 12096 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_223
timestamp 1754861848
transform 1 0 10248 0 1 18537
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_224
timestamp 1754861848
transform 1 0 10668 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_225
timestamp 1754861848
transform 1 0 12096 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_226
timestamp 1754861848
transform 1 0 4788 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_227
timestamp 1754861848
transform 1 0 6132 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_228
timestamp 1754861848
transform 1 0 5544 0 1 14141
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_229
timestamp 1754861848
transform 1 0 5208 0 1 13224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_230
timestamp 1754861848
transform 1 0 5460 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_231
timestamp 1754861848
transform 1 0 4704 0 1 13933
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_232
timestamp 1754861848
transform 1 0 5148 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_233
timestamp 1754861848
transform 1 0 6048 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_234
timestamp 1754861848
transform 1 0 5796 0 1 15456
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_235
timestamp 1754861848
transform 1 0 5292 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_236
timestamp 1754861848
transform 1 0 5376 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_237
timestamp 1754861848
transform 1 0 6300 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_238
timestamp 1754861848
transform 1 0 5916 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_239
timestamp 1754861848
transform 1 0 5262 0 1 17040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_240
timestamp 1754861848
transform 1 0 6216 0 1 18677
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_241
timestamp 1754861848
transform 1 0 4788 0 1 17039
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_242
timestamp 1754861848
transform 1 0 5544 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_243
timestamp 1754861848
transform 1 0 5460 0 1 17165
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_244
timestamp 1754861848
transform 1 0 6048 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_245
timestamp 1754861848
transform 1 0 5964 0 1 16896
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_246
timestamp 1754861848
transform 1 0 6300 0 1 16099
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_247
timestamp 1754861848
transform 1 0 5544 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_248
timestamp 1754861848
transform 1 0 6216 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_249
timestamp 1754861848
transform 1 0 12284 0 1 19235
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_250
timestamp 1754861848
transform 1 0 12012 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_251
timestamp 1754861848
transform 1 0 11256 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_252
timestamp 1754861848
transform 1 0 10836 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_253
timestamp 1754861848
transform 1 0 10584 0 1 19488
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_254
timestamp 1754861848
transform 1 0 9705 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_255
timestamp 1754861848
transform 1 0 9888 0 1 19248
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_256
timestamp 1754861848
transform 1 0 11130 0 1 20784
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_257
timestamp 1754861848
transform 1 0 12096 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_258
timestamp 1754861848
transform 1 0 10080 0 1 19123
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_259
timestamp 1754861848
transform 1 0 12390 0 1 21312
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_260
timestamp 1754861848
transform 1 0 10164 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_261
timestamp 1754861848
transform 1 0 11172 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_262
timestamp 1754861848
transform 1 0 12180 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_263
timestamp 1754861848
transform 1 0 10332 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_264
timestamp 1754861848
transform 1 0 8064 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_265
timestamp 1754861848
transform 1 0 6804 0 1 20640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_266
timestamp 1754861848
transform 1 0 7770 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_267
timestamp 1754861848
transform 1 0 7896 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_268
timestamp 1754861848
transform 1 0 8148 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_269
timestamp 1754861848
transform 1 0 6888 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_270
timestamp 1754861848
transform 1 0 6606 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_271
timestamp 1754861848
transform 1 0 9114 0 1 19123
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_272
timestamp 1754861848
transform 1 0 9198 0 1 19263
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_273
timestamp 1754861848
transform 1 0 6888 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_274
timestamp 1754861848
transform 1 0 7476 0 1 20640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_275
timestamp 1754861848
transform 1 0 8736 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_276
timestamp 1754861848
transform 1 0 8064 0 1 21504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_277
timestamp 1754861848
transform 1 0 8904 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_278
timestamp 1754861848
transform 1 0 7182 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_279
timestamp 1754861848
transform 1 0 6384 0 1 17664
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_280
timestamp 1754861848
transform 1 0 19488 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_281
timestamp 1754861848
transform 1 0 19908 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_282
timestamp 1754861848
transform 1 0 21504 0 1 14208
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_283
timestamp 1754861848
transform 1 0 19572 0 1 13177
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_284
timestamp 1754861848
transform 1 0 19236 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_285
timestamp 1754861848
transform 1 0 20412 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_286
timestamp 1754861848
transform 1 0 20328 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_287
timestamp 1754861848
transform 1 0 20748 0 1 13440
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_288
timestamp 1754861848
transform 1 0 20748 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_289
timestamp 1754861848
transform 1 0 19320 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_290
timestamp 1754861848
transform 1 0 20034 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_291
timestamp 1754861848
transform 1 0 20160 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_292
timestamp 1754861848
transform 1 0 19782 0 1 17735
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_293
timestamp 1754861848
transform 1 0 19740 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_294
timestamp 1754861848
transform 1 0 20916 0 1 17568
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_295
timestamp 1754861848
transform 1 0 19194 0 1 18336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_296
timestamp 1754861848
transform 1 0 19488 0 1 17184
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_297
timestamp 1754861848
transform 1 0 21504 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_298
timestamp 1754861848
transform 1 0 16028 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_299
timestamp 1754861848
transform 1 0 16632 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_300
timestamp 1754861848
transform 1 0 18732 0 1 13175
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_301
timestamp 1754861848
transform 1 0 17556 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_302
timestamp 1754861848
transform 1 0 16884 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_303
timestamp 1754861848
transform 1 0 18900 0 1 13728
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_304
timestamp 1754861848
transform 1 0 16422 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_305
timestamp 1754861848
transform 1 0 18522 0 1 14001
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_306
timestamp 1754861848
transform 1 0 18143 0 1 13173
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_307
timestamp 1754861848
transform 1 0 18228 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_308
timestamp 1754861848
transform 1 0 18564 0 1 14141
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_309
timestamp 1754861848
transform 1 0 18522 0 1 14736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_310
timestamp 1754861848
transform 1 0 17766 0 1 14496
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_311
timestamp 1754861848
transform 1 0 18396 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_312
timestamp 1754861848
transform 1 0 18228 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_313
timestamp 1754861848
transform 1 0 15918 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_314
timestamp 1754861848
transform 1 0 16044 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_315
timestamp 1754861848
transform 1 0 14952 0 1 15648
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_316
timestamp 1754861848
transform 1 0 14409 0 1 15504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_317
timestamp 1754861848
transform 1 0 15624 0 1 15648
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_318
timestamp 1754861848
transform 1 0 14490 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_319
timestamp 1754861848
transform 1 0 12852 0 1 15648
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_320
timestamp 1754861848
transform 1 0 15708 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_321
timestamp 1754861848
transform 1 0 15330 0 1 14592
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_322
timestamp 1754861848
transform 1 0 13608 0 1 13920
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_323
timestamp 1754861848
transform 1 0 15740 0 1 14064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_324
timestamp 1754861848
transform 1 0 13188 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_325
timestamp 1754861848
transform 1 0 14364 0 1 13152
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_326
timestamp 1754861848
transform 1 0 14196 0 1 15744
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_327
timestamp 1754861848
transform 1 0 14028 0 1 14688
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_328
timestamp 1754861848
transform 1 0 12936 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_329
timestamp 1754861848
transform 1 0 14196 0 1 14016
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_330
timestamp 1754861848
transform 1 0 15624 0 1 13174
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_331
timestamp 1754861848
transform 1 0 13146 0 1 13200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_332
timestamp 1754861848
transform 1 0 14784 0 1 15552
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_333
timestamp 1754861848
transform 1 0 13440 0 1 17952
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_334
timestamp 1754861848
transform 1 0 13818 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_335
timestamp 1754861848
transform 1 0 13608 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_336
timestamp 1754861848
transform 1 0 15162 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_337
timestamp 1754861848
transform 1 0 12936 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_338
timestamp 1754861848
transform 1 0 14112 0 1 16416
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_339
timestamp 1754861848
transform 1 0 15624 0 1 17040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_340
timestamp 1754861848
transform 1 0 15204 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_341
timestamp 1754861848
transform 1 0 14868 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_342
timestamp 1754861848
transform 1 0 12768 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_343
timestamp 1754861848
transform 1 0 13146 0 1 17040
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_344
timestamp 1754861848
transform 1 0 14364 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_345
timestamp 1754861848
transform 1 0 16380 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_346
timestamp 1754861848
transform 1 0 16716 0 1 18576
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_347
timestamp 1754861848
transform 1 0 18900 0 1 16128
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_348
timestamp 1754861848
transform 1 0 18522 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_349
timestamp 1754861848
transform 1 0 18060 0 1 16272
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_350
timestamp 1754861848
transform 1 0 18816 0 1 18336
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_351
timestamp 1754861848
transform 1 0 18312 0 1 17063
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_352
timestamp 1754861848
transform 1 0 17388 0 1 16272
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_353
timestamp 1754861848
transform 1 0 16716 0 1 17088
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_354
timestamp 1754861848
transform 1 0 17556 0 1 16512
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_355
timestamp 1754861848
transform 1 0 17304 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_356
timestamp 1754861848
transform 1 0 18228 0 1 16512
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_357
timestamp 1754861848
transform 1 0 16044 0 1 16224
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_358
timestamp 1754861848
transform 1 0 18900 0 1 17760
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_359
timestamp 1754861848
transform 1 0 17472 0 1 17065
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_360
timestamp 1754861848
transform 1 0 18144 0 1 18547
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_361
timestamp 1754861848
transform 1 0 15876 0 1 18528
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_362
timestamp 1754861848
transform 1 0 16632 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_363
timestamp 1754861848
transform 1 0 16632 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_364
timestamp 1754861848
transform 1 0 17850 0 1 19488
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_365
timestamp 1754861848
transform 1 0 17556 0 1 19221
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_366
timestamp 1754861848
transform 1 0 12936 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_367
timestamp 1754861848
transform 1 0 14868 0 1 20640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_368
timestamp 1754861848
transform 1 0 14364 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_369
timestamp 1754861848
transform 1 0 14112 0 1 19968
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_370
timestamp 1754861848
transform 1 0 13524 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_371
timestamp 1754861848
transform 1 0 15330 0 1 20640
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_372
timestamp 1754861848
transform 1 0 15740 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_373
timestamp 1754861848
transform 1 0 14112 0 1 21024
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_374
timestamp 1754861848
transform 1 0 14490 0 1 20733
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_375
timestamp 1754861848
transform 1 0 13440 0 1 20064
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_376
timestamp 1754861848
transform 1 0 15624 0 1 19200
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_377
timestamp 1754861848
transform 1 0 12768 0 1 21504
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_378
timestamp 1754861848
transform 1 0 15708 0 1 20736
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_379
timestamp 1754861848
transform 1 0 14868 0 1 19221
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_380
timestamp 1754861848
transform 1 0 13944 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_381
timestamp 1754861848
transform 1 0 14784 0 1 21600
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_382
timestamp 1754861848
transform 1 0 14112 0 1 19296
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_383
timestamp 1754861848
transform 1 0 13944 0 1 19104
box -29 -29 29 29
use VIA_Via1_XY  VIA_Via1_XY_384
timestamp 1754861848
transform 1 0 17388 0 1 19104
box -29 -29 29 29
use VIA_Via1_YY  VIA_Via1_YY_0
timestamp 1754861848
transform 1 0 17976 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_1
timestamp 1754861848
transform 1 0 17724 0 1 9696
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_2
timestamp 1754861848
transform 1 0 17472 0 1 9600
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_3
timestamp 1754861848
transform 1 0 18816 0 1 8544
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_4
timestamp 1754861848
transform 1 0 16212 0 1 9408
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_5
timestamp 1754861848
transform 1 0 18648 0 1 8736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_6
timestamp 1754861848
transform 1 0 18984 0 1 8736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_7
timestamp 1754861848
transform 1 0 12936 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_8
timestamp 1754861848
transform 1 0 13692 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_9
timestamp 1754861848
transform 1 0 15372 0 1 8448
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_10
timestamp 1754861848
transform 1 0 14952 0 1 8160
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_11
timestamp 1754861848
transform 1 0 12936 0 1 9504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_12
timestamp 1754861848
transform 1 0 14196 0 1 8160
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_13
timestamp 1754861848
transform 1 0 12852 0 1 7776
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_14
timestamp 1754861848
transform 1 0 15750 0 1 9512
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_15
timestamp 1754861848
transform 1 0 15834 0 1 9473
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_16
timestamp 1754861848
transform 1 0 14280 0 1 11676
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_17
timestamp 1754861848
transform 1 0 14280 0 1 10080
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_18
timestamp 1754861848
transform 1 0 12936 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_19
timestamp 1754861848
transform 1 0 14784 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_20
timestamp 1754861848
transform 1 0 14112 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_21
timestamp 1754861848
transform 1 0 13692 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_22
timestamp 1754861848
transform 1 0 12852 0 1 10080
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_23
timestamp 1754861848
transform 1 0 15456 0 1 11040
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_24
timestamp 1754861848
transform 1 0 12768 0 1 11040
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_25
timestamp 1754861848
transform 1 0 13860 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_26
timestamp 1754861848
transform 1 0 12768 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_27
timestamp 1754861848
transform 1 0 13188 0 1 10464
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_28
timestamp 1754861848
transform 1 0 14112 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_29
timestamp 1754861848
transform 1 0 15204 0 1 10752
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_30
timestamp 1754861848
transform 1 0 16758 0 1 11664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_31
timestamp 1754861848
transform 1 0 17556 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_32
timestamp 1754861848
transform 1 0 18606 0 1 11616
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_33
timestamp 1754861848
transform 1 0 17094 0 1 10464
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_34
timestamp 1754861848
transform 1 0 17346 0 1 12432
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_35
timestamp 1754861848
transform 1 0 17220 0 1 12288
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_36
timestamp 1754861848
transform 1 0 16884 0 1 10224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_37
timestamp 1754861848
transform 1 0 18564 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_38
timestamp 1754861848
transform 1 0 18312 0 1 11904
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_39
timestamp 1754861848
transform 1 0 17892 0 1 11136
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_40
timestamp 1754861848
transform 1 0 18228 0 1 12576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_41
timestamp 1754861848
transform 1 0 18144 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_42
timestamp 1754861848
transform 1 0 17976 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_43
timestamp 1754861848
transform 1 0 22008 0 1 9216
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_44
timestamp 1754861848
transform 1 0 19404 0 1 9696
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_45
timestamp 1754861848
transform 1 0 19194 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_46
timestamp 1754861848
transform 1 0 19304 0 1 9495
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_47
timestamp 1754861848
transform 1 0 19110 0 1 9360
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_48
timestamp 1754861848
transform 1 0 21336 0 1 11712
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_49
timestamp 1754861848
transform 1 0 19992 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_50
timestamp 1754861848
transform 1 0 19572 0 1 10752
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_51
timestamp 1754861848
transform 1 0 19824 0 1 11676
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_52
timestamp 1754861848
transform 1 0 20832 0 1 10752
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_53
timestamp 1754861848
transform 1 0 21107 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_54
timestamp 1754861848
transform 1 0 20370 0 1 12515
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_55
timestamp 1754861848
transform 1 0 20664 0 1 9984
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_56
timestamp 1754861848
transform 1 0 21203 0 1 11664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_57
timestamp 1754861848
transform 1 0 19992 0 1 12433
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_58
timestamp 1754861848
transform 1 0 21672 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_59
timestamp 1754861848
transform 1 0 19404 0 1 12288
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_60
timestamp 1754861848
transform 1 0 20160 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_61
timestamp 1754861848
transform 1 0 20454 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_62
timestamp 1754861848
transform 1 0 21000 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_63
timestamp 1754861848
transform 1 0 21210 0 1 9984
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_64
timestamp 1754861848
transform 1 0 19068 0 1 11040
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_65
timestamp 1754861848
transform 1 0 7003 0 1 6455
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_66
timestamp 1754861848
transform 1 0 7224 0 1 6336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_67
timestamp 1754861848
transform 1 0 7476 0 1 6240
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_68
timestamp 1754861848
transform 1 0 7224 0 1 6480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_69
timestamp 1754861848
transform 1 0 9107 0 1 6453
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_70
timestamp 1754861848
transform 1 0 8232 0 1 6480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_71
timestamp 1754861848
transform 1 0 9582 0 1 6471
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_72
timestamp 1754861848
transform 1 0 9408 0 1 6480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_73
timestamp 1754861848
transform 1 0 8904 0 1 6480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_74
timestamp 1754861848
transform 1 0 8459 0 1 6453
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_75
timestamp 1754861848
transform 1 0 4116 0 1 6624
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_76
timestamp 1754861848
transform 1 0 5103 0 1 6480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_77
timestamp 1754861848
transform 1 0 5544 0 1 6467
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_78
timestamp 1754861848
transform 1 0 4979 0 1 6453
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_79
timestamp 1754861848
transform 1 0 5771 0 1 6453
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_80
timestamp 1754861848
transform 1 0 5796 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_81
timestamp 1754861848
transform 1 0 4620 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_82
timestamp 1754861848
transform 1 0 4788 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_83
timestamp 1754861848
transform 1 0 4116 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_84
timestamp 1754861848
transform 1 0 4423 0 1 8667
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_85
timestamp 1754861848
transform 1 0 5460 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_86
timestamp 1754861848
transform 1 0 5712 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_87
timestamp 1754861848
transform 1 0 4998 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_88
timestamp 1754861848
transform 1 0 4494 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_89
timestamp 1754861848
transform 1 0 5964 0 1 9696
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_90
timestamp 1754861848
transform 1 0 5376 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_91
timestamp 1754861848
transform 1 0 5880 0 1 8448
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_92
timestamp 1754861848
transform 1 0 4242 0 1 7133
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_93
timestamp 1754861848
transform 1 0 4620 0 1 8448
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_94
timestamp 1754861848
transform 1 0 3948 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_95
timestamp 1754861848
transform 1 0 4032 0 1 7008
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_96
timestamp 1754861848
transform 1 0 4494 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_97
timestamp 1754861848
transform 1 0 4872 0 1 7152
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_98
timestamp 1754861848
transform 1 0 4872 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_99
timestamp 1754861848
transform 1 0 5712 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_100
timestamp 1754861848
transform 1 0 5095 0 1 8657
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_101
timestamp 1754861848
transform 1 0 6268 0 1 9493
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_102
timestamp 1754861848
transform 1 0 6132 0 1 11904
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_103
timestamp 1754861848
transform 1 0 5964 0 1 12437
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_104
timestamp 1754861848
transform 1 0 6132 0 1 12384
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_105
timestamp 1754861848
transform 1 0 6300 0 1 11616
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_106
timestamp 1754861848
transform 1 0 5796 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_107
timestamp 1754861848
transform 1 0 4788 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_108
timestamp 1754861848
transform 1 0 5964 0 1 11763
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_109
timestamp 1754861848
transform 1 0 5376 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_110
timestamp 1754861848
transform 1 0 5628 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_111
timestamp 1754861848
transform 1 0 5460 0 1 12576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_112
timestamp 1754861848
transform 1 0 4872 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_113
timestamp 1754861848
transform 1 0 5544 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_114
timestamp 1754861848
transform 1 0 11424 0 1 8668
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_115
timestamp 1754861848
transform 1 0 11340 0 1 7776
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_116
timestamp 1754861848
transform 1 0 10668 0 1 8832
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_117
timestamp 1754861848
transform 1 0 11508 0 1 8688
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_118
timestamp 1754861848
transform 1 0 11634 0 1 8448
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_119
timestamp 1754861848
transform 1 0 12390 0 1 7200
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_120
timestamp 1754861848
transform 1 0 10248 0 1 9504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_121
timestamp 1754861848
transform 1 0 9576 0 1 8832
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_122
timestamp 1754861848
transform 1 0 11790 0 1 8739
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_123
timestamp 1754861848
transform 1 0 10080 0 1 8736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_124
timestamp 1754861848
transform 1 0 9576 0 1 9696
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_125
timestamp 1754861848
transform 1 0 11928 0 1 7200
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_126
timestamp 1754861848
transform 1 0 11088 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_127
timestamp 1754861848
transform 1 0 9996 0 1 8544
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_128
timestamp 1754861848
transform 1 0 10836 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_129
timestamp 1754861848
transform 1 0 12684 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_130
timestamp 1754861848
transform 1 0 11676 0 1 8160
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_131
timestamp 1754861848
transform 1 0 9828 0 1 9504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_132
timestamp 1754861848
transform 1 0 12096 0 1 7392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_133
timestamp 1754861848
transform 1 0 12264 0 1 7152
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_134
timestamp 1754861848
transform 1 0 12264 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_135
timestamp 1754861848
transform 1 0 8764 0 1 8651
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_136
timestamp 1754861848
transform 1 0 7056 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_137
timestamp 1754861848
transform 1 0 8316 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_138
timestamp 1754861848
transform 1 0 8437 0 1 7982
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_139
timestamp 1754861848
transform 1 0 9114 0 1 9360
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_140
timestamp 1754861848
transform 1 0 8316 0 1 7152
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_141
timestamp 1754861848
transform 1 0 9156 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_142
timestamp 1754861848
transform 1 0 6468 0 1 9408
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_143
timestamp 1754861848
transform 1 0 8316 0 1 9484
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_144
timestamp 1754861848
transform 1 0 8148 0 1 9600
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_145
timestamp 1754861848
transform 1 0 7938 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_146
timestamp 1754861848
transform 1 0 7812 0 1 7104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_147
timestamp 1754861848
transform 1 0 7665 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_148
timestamp 1754861848
transform 1 0 8820 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_149
timestamp 1754861848
transform 1 0 8904 0 1 7968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_150
timestamp 1754861848
transform 1 0 7224 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_151
timestamp 1754861848
transform 1 0 6972 0 1 8928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_152
timestamp 1754861848
transform 1 0 8652 0 1 8652
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_153
timestamp 1754861848
transform 1 0 7477 0 1 7155
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_154
timestamp 1754861848
transform 1 0 6720 0 1 8640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_155
timestamp 1754861848
transform 1 0 9408 0 1 11712
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_156
timestamp 1754861848
transform 1 0 9324 0 1 11040
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_157
timestamp 1754861848
transform 1 0 8988 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_158
timestamp 1754861848
transform 1 0 9156 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_159
timestamp 1754861848
transform 1 0 7980 0 1 12288
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_160
timestamp 1754861848
transform 1 0 8263 0 1 11015
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_161
timestamp 1754861848
transform 1 0 8064 0 1 11015
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_162
timestamp 1754861848
transform 1 0 6972 0 1 12576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_163
timestamp 1754861848
transform 1 0 8652 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_164
timestamp 1754861848
transform 1 0 7476 0 1 12384
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_165
timestamp 1754861848
transform 1 0 7476 0 1 11088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_166
timestamp 1754861848
transform 1 0 9492 0 1 11616
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_167
timestamp 1754861848
transform 1 0 8526 0 1 12536
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_168
timestamp 1754861848
transform 1 0 6552 0 1 12384
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_169
timestamp 1754861848
transform 1 0 7392 0 1 11008
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_170
timestamp 1754861848
transform 1 0 8736 0 1 11712
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_171
timestamp 1754861848
transform 1 0 6552 0 1 11136
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_172
timestamp 1754861848
transform 1 0 7812 0 1 10752
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_173
timestamp 1754861848
transform 1 0 12348 0 1 10944
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_174
timestamp 1754861848
transform 1 0 12600 0 1 11136
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_175
timestamp 1754861848
transform 1 0 9576 0 1 10848
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_176
timestamp 1754861848
transform 1 0 11004 0 1 10992
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_177
timestamp 1754861848
transform 1 0 10920 0 1 12288
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_178
timestamp 1754861848
transform 1 0 10080 0 1 12480
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_179
timestamp 1754861848
transform 1 0 9828 0 1 11520
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_180
timestamp 1754861848
transform 1 0 9954 0 1 11616
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_181
timestamp 1754861848
transform 1 0 10752 0 1 10368
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_182
timestamp 1754861848
transform 1 0 11424 0 1 12576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_183
timestamp 1754861848
transform 1 0 10458 0 1 10080
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_184
timestamp 1754861848
transform 1 0 11172 0 1 10176
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_185
timestamp 1754861848
transform 1 0 10332 0 1 12672
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_186
timestamp 1754861848
transform 1 0 12012 0 1 13440
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_187
timestamp 1754861848
transform 1 0 11073 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_188
timestamp 1754861848
transform 1 0 12348 0 1 14088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_189
timestamp 1754861848
transform 1 0 11424 0 1 13824
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_190
timestamp 1754861848
transform 1 0 12390 0 1 15648
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_191
timestamp 1754861848
transform 1 0 11844 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_192
timestamp 1754861848
transform 1 0 9912 0 1 13056
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_193
timestamp 1754861848
transform 1 0 10164 0 1 13941
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_194
timestamp 1754861848
transform 1 0 12600 0 1 14976
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_195
timestamp 1754861848
transform 1 0 10471 0 1 13181
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_196
timestamp 1754861848
transform 1 0 11827 0 1 13271
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_197
timestamp 1754861848
transform 1 0 10374 0 1 14208
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_198
timestamp 1754861848
transform 1 0 9828 0 1 15648
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_199
timestamp 1754861848
transform 1 0 7266 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_200
timestamp 1754861848
transform 1 0 9408 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_201
timestamp 1754861848
transform 1 0 7056 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_202
timestamp 1754861848
transform 1 0 8148 0 1 15360
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_203
timestamp 1754861848
transform 1 0 7560 0 1 14688
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_204
timestamp 1754861848
transform 1 0 8442 0 1 15648
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_205
timestamp 1754861848
transform 1 0 8484 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_206
timestamp 1754861848
transform 1 0 8820 0 1 15360
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_207
timestamp 1754861848
transform 1 0 7728 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_208
timestamp 1754861848
transform 1 0 7644 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_209
timestamp 1754861848
transform 1 0 7224 0 1 13440
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_210
timestamp 1754861848
transform 1 0 6720 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_211
timestamp 1754861848
transform 1 0 6552 0 1 17184
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_212
timestamp 1754861848
transform 1 0 8064 0 1 17704
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_213
timestamp 1754861848
transform 1 0 9492 0 1 18477
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_214
timestamp 1754861848
transform 1 0 6804 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_215
timestamp 1754861848
transform 1 0 9240 0 1 16320
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_216
timestamp 1754861848
transform 1 0 8148 0 1 17743
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_217
timestamp 1754861848
transform 1 0 6888 0 1 18528
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_218
timestamp 1754861848
transform 1 0 12684 0 1 17184
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_219
timestamp 1754861848
transform 1 0 12264 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_220
timestamp 1754861848
transform 1 0 10080 0 1 16272
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_221
timestamp 1754861848
transform 1 0 9912 0 1 16992
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_222
timestamp 1754861848
transform 1 0 9642 0 1 17729
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_223
timestamp 1754861848
transform 1 0 10038 0 1 17725
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_224
timestamp 1754861848
transform 1 0 9828 0 1 17760
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_225
timestamp 1754861848
transform 1 0 10332 0 1 17952
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_226
timestamp 1754861848
transform 1 0 11256 0 1 16416
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_227
timestamp 1754861848
transform 1 0 10584 0 1 17725
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_228
timestamp 1754861848
transform 1 0 10752 0 1 17568
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_229
timestamp 1754861848
transform 1 0 10571 0 1 16224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_230
timestamp 1754861848
transform 1 0 9996 0 1 16224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_231
timestamp 1754861848
transform 1 0 11088 0 1 16224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_232
timestamp 1754861848
transform 1 0 12180 0 1 18432
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_233
timestamp 1754861848
transform 1 0 11256 0 1 18336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_234
timestamp 1754861848
transform 1 0 10248 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_235
timestamp 1754861848
transform 1 0 10374 0 1 17760
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_236
timestamp 1754861848
transform 1 0 11676 0 1 18624
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_237
timestamp 1754861848
transform 1 0 11424 0 1 17088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_238
timestamp 1754861848
transform 1 0 11676 0 1 16128
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_239
timestamp 1754861848
transform 1 0 9702 0 1 18720
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_240
timestamp 1754861848
transform 1 0 11760 0 1 16896
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_241
timestamp 1754861848
transform 1 0 12348 0 1 18624
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_242
timestamp 1754861848
transform 1 0 11508 0 1 16320
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_243
timestamp 1754861848
transform 1 0 11004 0 1 17760
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_244
timestamp 1754861848
transform 1 0 5964 0 1 15264
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_245
timestamp 1754861848
transform 1 0 4536 0 1 15456
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_246
timestamp 1754861848
transform 1 0 5880 0 1 14208
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_247
timestamp 1754861848
transform 1 0 4424 0 1 14023
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_248
timestamp 1754861848
transform 1 0 4704 0 1 14880
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_249
timestamp 1754861848
transform 1 0 4620 0 1 13344
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_250
timestamp 1754861848
transform 1 0 6132 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_251
timestamp 1754861848
transform 1 0 4872 0 1 14688
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_252
timestamp 1754861848
transform 1 0 4536 0 1 13824
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_253
timestamp 1754861848
transform 1 0 4872 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_254
timestamp 1754861848
transform 1 0 6300 0 1 16992
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_255
timestamp 1754861848
transform 1 0 6300 0 1 18576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_256
timestamp 1754861848
transform 1 0 5166 0 1 17664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_257
timestamp 1754861848
transform 1 0 5544 0 1 16224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_258
timestamp 1754861848
transform 1 0 5544 0 1 18336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_259
timestamp 1754861848
transform 1 0 4872 0 1 17184
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_260
timestamp 1754861848
transform 1 0 5376 0 1 16032
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_261
timestamp 1754861848
transform 1 0 10164 0 1 19872
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_262
timestamp 1754861848
transform 1 0 11004 0 1 20736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_263
timestamp 1754861848
transform 1 0 9576 0 1 19488
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_264
timestamp 1754861848
transform 1 0 12684 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_265
timestamp 1754861848
transform 1 0 9954 0 1 21552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_266
timestamp 1754861848
transform 1 0 11340 0 1 19392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_267
timestamp 1754861848
transform 1 0 10752 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_268
timestamp 1754861848
transform 1 0 10920 0 1 19392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_269
timestamp 1754861848
transform 1 0 11676 0 1 20736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_270
timestamp 1754861848
transform 1 0 11508 0 1 20928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_271
timestamp 1754861848
transform 1 0 10584 0 1 19872
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_272
timestamp 1754861848
transform 1 0 10584 0 1 20928
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_273
timestamp 1754861848
transform 1 0 11928 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_274
timestamp 1754861848
transform 1 0 9912 0 1 20544
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_275
timestamp 1754861848
transform 1 0 11676 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_276
timestamp 1754861848
transform 1 0 11155 0 1 19319
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_277
timestamp 1754861848
transform 1 0 8988 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_278
timestamp 1754861848
transform 1 0 9324 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_279
timestamp 1754861848
transform 1 0 8820 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_280
timestamp 1754861848
transform 1 0 8652 0 1 19392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_281
timestamp 1754861848
transform 1 0 6804 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_282
timestamp 1754861848
transform 1 0 7014 0 1 19392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_283
timestamp 1754861848
transform 1 0 7308 0 1 20544
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_284
timestamp 1754861848
transform 1 0 9030 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_285
timestamp 1754861848
transform 1 0 7644 0 1 19488
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_286
timestamp 1754861848
transform 1 0 7308 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_287
timestamp 1754861848
transform 1 0 7224 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_288
timestamp 1754861848
transform 1 0 7560 0 1 19968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_289
timestamp 1754861848
transform 1 0 8467 0 1 19319
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_290
timestamp 1754861848
transform 1 0 8467 0 1 21501
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_291
timestamp 1754861848
transform 1 0 8652 0 1 21408
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_292
timestamp 1754861848
transform 1 0 7392 0 1 19104
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_293
timestamp 1754861848
transform 1 0 21924 0 1 15264
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_294
timestamp 1754861848
transform 1 0 21336 0 1 13248
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_295
timestamp 1754861848
transform 1 0 21504 0 1 13440
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_296
timestamp 1754861848
transform 1 0 21798 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_297
timestamp 1754861848
transform 1 0 19152 0 1 15744
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_298
timestamp 1754861848
transform 1 0 19488 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_299
timestamp 1754861848
transform 1 0 20748 0 1 14592
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_300
timestamp 1754861848
transform 1 0 21672 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_301
timestamp 1754861848
transform 1 0 21126 0 1 13405
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_302
timestamp 1754861848
transform 1 0 21798 0 1 14832
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_303
timestamp 1754861848
transform 1 0 21336 0 1 16032
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_304
timestamp 1754861848
transform 1 0 20160 0 1 17088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_305
timestamp 1754861848
transform 1 0 20748 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_306
timestamp 1754861848
transform 1 0 19992 0 1 18336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_307
timestamp 1754861848
transform 1 0 19488 0 1 18336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_308
timestamp 1754861848
transform 1 0 21588 0 1 16032
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_309
timestamp 1754861848
transform 1 0 20412 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_310
timestamp 1754861848
transform 1 0 19859 0 1 18551
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_311
timestamp 1754861848
transform 1 0 19404 0 1 18563
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_312
timestamp 1754861848
transform 1 0 20648 0 1 17047
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_313
timestamp 1754861848
transform 1 0 18816 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_314
timestamp 1754861848
transform 1 0 16128 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_315
timestamp 1754861848
transform 1 0 17766 0 1 14208
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_316
timestamp 1754861848
transform 1 0 18060 0 1 13056
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_317
timestamp 1754861848
transform 1 0 18690 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_318
timestamp 1754861848
transform 1 0 18312 0 1 13152
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_319
timestamp 1754861848
transform 1 0 16715 0 1 14029
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_320
timestamp 1754861848
transform 1 0 17388 0 1 14112
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_321
timestamp 1754861848
transform 1 0 18396 0 1 14688
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_322
timestamp 1754861848
transform 1 0 17220 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_323
timestamp 1754861848
transform 1 0 18060 0 1 15456
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_324
timestamp 1754861848
transform 1 0 16979 0 1 13187
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_325
timestamp 1754861848
transform 1 0 17835 0 1 13189
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_326
timestamp 1754861848
transform 1 0 16254 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_327
timestamp 1754861848
transform 1 0 16548 0 1 13248
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_328
timestamp 1754861848
transform 1 0 17472 0 1 13202
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_329
timestamp 1754861848
transform 1 0 17839 0 1 14019
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_330
timestamp 1754861848
transform 1 0 18900 0 1 14880
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_331
timestamp 1754861848
transform 1 0 17724 0 1 13248
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_332
timestamp 1754861848
transform 1 0 15204 0 1 14496
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_333
timestamp 1754861848
transform 1 0 15150 0 1 13968
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_334
timestamp 1754861848
transform 1 0 14868 0 1 13824
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_335
timestamp 1754861848
transform 1 0 15624 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_336
timestamp 1754861848
transform 1 0 12768 0 1 14688
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_337
timestamp 1754861848
transform 1 0 13356 0 1 15744
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_338
timestamp 1754861848
transform 1 0 13043 0 1 14039
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_339
timestamp 1754861848
transform 1 0 15036 0 1 15552
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_340
timestamp 1754861848
transform 1 0 15456 0 1 15744
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_341
timestamp 1754861848
transform 1 0 14364 0 1 14088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_342
timestamp 1754861848
transform 1 0 12936 0 1 13344
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_343
timestamp 1754861848
transform 1 0 14028 0 1 15456
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_344
timestamp 1754861848
transform 1 0 13146 0 1 14208
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_345
timestamp 1754861848
transform 1 0 13524 0 1 15456
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_346
timestamp 1754861848
transform 1 0 13734 0 1 15264
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_347
timestamp 1754861848
transform 1 0 12852 0 1 13920
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_348
timestamp 1754861848
transform 1 0 13860 0 1 14016
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_349
timestamp 1754861848
transform 1 0 13524 0 1 13216
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_350
timestamp 1754861848
transform 1 0 15540 0 1 17952
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_351
timestamp 1754861848
transform 1 0 13524 0 1 17024
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_352
timestamp 1754861848
transform 1 0 14490 0 1 16429
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_353
timestamp 1754861848
transform 1 0 14532 0 1 17568
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_354
timestamp 1754861848
transform 1 0 14784 0 1 16224
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_355
timestamp 1754861848
transform 1 0 15036 0 1 17664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_356
timestamp 1754861848
transform 1 0 15288 0 1 18432
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_357
timestamp 1754861848
transform 1 0 14112 0 1 17760
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_358
timestamp 1754861848
transform 1 0 14784 0 1 18528
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_359
timestamp 1754861848
transform 1 0 14196 0 1 17664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_360
timestamp 1754861848
transform 1 0 15731 0 1 17712
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_361
timestamp 1754861848
transform 1 0 15456 0 1 18528
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_362
timestamp 1754861848
transform 1 0 15834 0 1 17856
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_363
timestamp 1754861848
transform 1 0 18396 0 1 18576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_364
timestamp 1754861848
transform 1 0 18312 0 1 18576
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_365
timestamp 1754861848
transform 1 0 16674 0 1 17743
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_366
timestamp 1754861848
transform 1 0 17892 0 1 18336
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_367
timestamp 1754861848
transform 1 0 16800 0 1 17664
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_368
timestamp 1754861848
transform 1 0 17220 0 1 16416
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_369
timestamp 1754861848
transform 1 0 17052 0 1 17856
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_370
timestamp 1754861848
transform 1 0 16128 0 1 17568
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_371
timestamp 1754861848
transform 1 0 16044 0 1 16896
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_372
timestamp 1754861848
transform 1 0 18732 0 1 16416
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_373
timestamp 1754861848
transform 1 0 17052 0 1 17088
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_374
timestamp 1754861848
transform 1 0 16296 0 1 16800
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_375
timestamp 1754861848
transform 1 0 16044 0 1 17725
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_376
timestamp 1754861848
transform 1 0 17640 0 1 17856
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_377
timestamp 1754861848
transform 1 0 17640 0 1 19872
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_378
timestamp 1754861848
transform 1 0 16128 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_379
timestamp 1754861848
transform 1 0 17839 0 1 19245
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_380
timestamp 1754861848
transform 1 0 16254 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_381
timestamp 1754861848
transform 1 0 17766 0 1 20640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_382
timestamp 1754861848
transform 1 0 17220 0 1 19241
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_383
timestamp 1754861848
transform 1 0 17304 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_384
timestamp 1754861848
transform 1 0 16884 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_385
timestamp 1754861848
transform 1 0 16715 0 1 19263
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_386
timestamp 1754861848
transform 1 0 17838 0 1 21501
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_387
timestamp 1754861848
transform 1 0 15960 0 1 21312
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_388
timestamp 1754861848
transform 1 0 17976 0 1 19872
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_389
timestamp 1754861848
transform 1 0 18648 0 1 19200
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_390
timestamp 1754861848
transform 1 0 18228 0 1 19392
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_391
timestamp 1754861848
transform 1 0 17472 0 1 21792
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_392
timestamp 1754861848
transform 1 0 18396 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_393
timestamp 1754861848
transform 1 0 17094 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_394
timestamp 1754861848
transform 1 0 18060 0 1 21504
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_395
timestamp 1754861848
transform 1 0 17843 0 1 20063
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_396
timestamp 1754861848
transform 1 0 16464 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_397
timestamp 1754861848
transform 1 0 16212 0 1 21600
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_398
timestamp 1754861848
transform 1 0 15151 0 1 19245
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_399
timestamp 1754861848
transform 1 0 13776 0 1 19245
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_400
timestamp 1754861848
transform 1 0 14784 0 1 20736
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_401
timestamp 1754861848
transform 1 0 13259 0 1 19263
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_402
timestamp 1754861848
transform 1 0 14280 0 1 19488
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_403
timestamp 1754861848
transform 1 0 12936 0 1 21792
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_404
timestamp 1754861848
transform 1 0 14700 0 1 19488
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_405
timestamp 1754861848
transform 1 0 13230 0 1 21600
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_406
timestamp 1754861848
transform 1 0 12768 0 1 19296
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_407
timestamp 1754861848
transform 1 0 13188 0 1 19872
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_408
timestamp 1754861848
transform 1 0 13692 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_409
timestamp 1754861848
transform 1 0 14478 0 1 19319
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_410
timestamp 1754861848
transform 1 0 14658 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_411
timestamp 1754861848
transform 1 0 15624 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_412
timestamp 1754861848
transform 1 0 15204 0 1 20640
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_413
timestamp 1754861848
transform 1 0 14784 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_414
timestamp 1754861848
transform 1 0 13608 0 1 20092
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_415
timestamp 1754861848
transform 1 0 15246 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_416
timestamp 1754861848
transform 1 0 15120 0 1 20064
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_417
timestamp 1754861848
transform 1 0 19068 0 1 14112
box -21 -29 21 29
use VIA_Via1_YY  VIA_Via1_YY_418
timestamp 1754861848
transform 1 0 15078 0 1 19104
box -21 -29 21 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_0
timestamp 1754861848
transform 1 0 21200 0 1 5292
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_1
timestamp 1754861848
transform 1 0 21200 0 1 3780
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_2
timestamp 1754861848
transform 1 0 13640 0 1 4536
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_3
timestamp 1754861848
transform 1 0 13640 0 1 6048
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_4
timestamp 1754861848
transform 1 0 13640 0 1 9072
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_5
timestamp 1754861848
transform 1 0 13640 0 1 7560
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_6
timestamp 1754861848
transform 1 0 13640 0 1 12096
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_7
timestamp 1754861848
transform 1 0 13640 0 1 10584
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_8
timestamp 1754861848
transform 1 0 21200 0 1 6804
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_9
timestamp 1754861848
transform 1 0 21200 0 1 8316
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_10
timestamp 1754861848
transform 1 0 21200 0 1 9828
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_11
timestamp 1754861848
transform 1 0 21200 0 1 11340
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_12
timestamp 1754861848
transform 1 0 6080 0 1 3780
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_13
timestamp 1754861848
transform 1 0 6080 0 1 5292
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_14
timestamp 1754861848
transform 1 0 6080 0 1 8316
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_15
timestamp 1754861848
transform 1 0 6080 0 1 6804
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_16
timestamp 1754861848
transform 1 0 6080 0 1 11340
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_17
timestamp 1754861848
transform 1 0 6080 0 1 9828
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_18
timestamp 1754861848
transform 1 0 6080 0 1 15876
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_19
timestamp 1754861848
transform 1 0 6080 0 1 14364
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_20
timestamp 1754861848
transform 1 0 6080 0 1 18900
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_21
timestamp 1754861848
transform 1 0 6080 0 1 17388
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_22
timestamp 1754861848
transform 1 0 6080 0 1 20412
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_23
timestamp 1754861848
transform 1 0 6080 0 1 21924
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_24
timestamp 1754861848
transform 1 0 21200 0 1 15876
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_25
timestamp 1754861848
transform 1 0 21200 0 1 14364
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_26
timestamp 1754861848
transform 1 0 21200 0 1 17388
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_27
timestamp 1754861848
transform 1 0 21200 0 1 18900
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_28
timestamp 1754861848
transform 1 0 13640 0 1 13608
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_29
timestamp 1754861848
transform 1 0 13640 0 1 15120
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_30
timestamp 1754861848
transform 1 0 13640 0 1 16632
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_31
timestamp 1754861848
transform 1 0 13640 0 1 18144
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_32
timestamp 1754861848
transform 1 0 13640 0 1 19656
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_33
timestamp 1754861848
transform 1 0 13640 0 1 21168
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_34
timestamp 1754861848
transform 1 0 21200 0 1 21924
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_35
timestamp 1754861848
transform 1 0 21200 0 1 20412
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_36
timestamp 1754861848
transform 1 0 21200 0 1 12852
box -193 -29 193 29
use VIA_via2_3_2200_440_1_5_410_410  VIA_via2_3_2200_440_1_5_410_410_37
timestamp 1754861848
transform 1 0 6080 0 1 12852
box -193 -29 193 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_0
timestamp 1754861848
transform 1 0 23480 0 1 5292
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_1
timestamp 1754861848
transform 1 0 23480 0 1 3780
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_2
timestamp 1754861848
transform 1 0 24880 0 1 6048
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_3
timestamp 1754861848
transform 1 0 24880 0 1 4536
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_4
timestamp 1754861848
transform 1 0 23480 0 1 6804
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_5
timestamp 1754861848
transform 1 0 24880 0 1 9072
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_6
timestamp 1754861848
transform 1 0 23480 0 1 8316
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_7
timestamp 1754861848
transform 1 0 24880 0 1 7560
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_8
timestamp 1754861848
transform 1 0 24880 0 1 12096
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_9
timestamp 1754861848
transform 1 0 24880 0 1 10584
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_10
timestamp 1754861848
transform 1 0 23480 0 1 11340
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_11
timestamp 1754861848
transform 1 0 23480 0 1 9828
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_12
timestamp 1754861848
transform 1 0 1960 0 1 5292
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_13
timestamp 1754861848
transform 1 0 560 0 1 4536
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_14
timestamp 1754861848
transform 1 0 560 0 1 6048
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_15
timestamp 1754861848
transform 1 0 1960 0 1 3780
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_16
timestamp 1754861848
transform 1 0 1960 0 1 6804
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_17
timestamp 1754861848
transform 1 0 560 0 1 7560
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_18
timestamp 1754861848
transform 1 0 560 0 1 9072
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_19
timestamp 1754861848
transform 1 0 1960 0 1 8316
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_20
timestamp 1754861848
transform 1 0 1960 0 1 9828
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_21
timestamp 1754861848
transform 1 0 560 0 1 10584
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_22
timestamp 1754861848
transform 1 0 560 0 1 12096
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_23
timestamp 1754861848
transform 1 0 1960 0 1 11340
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_24
timestamp 1754861848
transform 1 0 560 0 1 15120
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_25
timestamp 1754861848
transform 1 0 1960 0 1 15876
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_26
timestamp 1754861848
transform 1 0 1960 0 1 14364
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_27
timestamp 1754861848
transform 1 0 560 0 1 13608
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_28
timestamp 1754861848
transform 1 0 1960 0 1 18900
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_29
timestamp 1754861848
transform 1 0 1960 0 1 17388
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_30
timestamp 1754861848
transform 1 0 560 0 1 16632
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_31
timestamp 1754861848
transform 1 0 560 0 1 18144
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_32
timestamp 1754861848
transform 1 0 1960 0 1 20412
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_33
timestamp 1754861848
transform 1 0 560 0 1 21168
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_34
timestamp 1754861848
transform 1 0 560 0 1 19656
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_35
timestamp 1754861848
transform 1 0 1960 0 1 21924
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_36
timestamp 1754861848
transform 1 0 23480 0 1 15876
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_37
timestamp 1754861848
transform 1 0 24880 0 1 15120
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_38
timestamp 1754861848
transform 1 0 23480 0 1 14364
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_39
timestamp 1754861848
transform 1 0 24880 0 1 13608
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_40
timestamp 1754861848
transform 1 0 23480 0 1 17388
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_41
timestamp 1754861848
transform 1 0 24880 0 1 16632
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_42
timestamp 1754861848
transform 1 0 24880 0 1 18144
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_43
timestamp 1754861848
transform 1 0 23480 0 1 18900
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_44
timestamp 1754861848
transform 1 0 23480 0 1 21924
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_45
timestamp 1754861848
transform 1 0 24880 0 1 19656
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_46
timestamp 1754861848
transform 1 0 24880 0 1 21168
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_47
timestamp 1754861848
transform 1 0 23480 0 1 20412
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_48
timestamp 1754861848
transform 1 0 23480 0 1 12852
box -480 -29 480 29
use VIA_via2_3_5000_440_1_12_410_410  VIA_via2_3_5000_440_1_12_410_410_49
timestamp 1754861848
transform 1 0 1960 0 1 12852
box -480 -29 480 29
use VIA_Via2_YX  VIA_Via2_YX_0
timestamp 1754861848
transform 1 0 17472 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_1
timestamp 1754861848
transform 1 0 18984 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_2
timestamp 1754861848
transform 1 0 16212 0 1 9408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_3
timestamp 1754861848
transform 1 0 16800 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_4
timestamp 1754861848
transform 1 0 16716 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_5
timestamp 1754861848
transform 1 0 17976 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_6
timestamp 1754861848
transform 1 0 18228 0 1 9312
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_7
timestamp 1754861848
transform 1 0 16338 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_8
timestamp 1754861848
transform 1 0 18816 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_9
timestamp 1754861848
transform 1 0 17808 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_10
timestamp 1754861848
transform 1 0 18732 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_11
timestamp 1754861848
transform 1 0 18396 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_12
timestamp 1754861848
transform 1 0 16716 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_13
timestamp 1754861848
transform 1 0 18438 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_14
timestamp 1754861848
transform 1 0 14784 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_15
timestamp 1754861848
transform 1 0 15372 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_16
timestamp 1754861848
transform 1 0 15372 0 1 9408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_17
timestamp 1754861848
transform 1 0 14196 0 1 8160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_18
timestamp 1754861848
transform 1 0 15288 0 1 8160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_19
timestamp 1754861848
transform 1 0 14868 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_20
timestamp 1754861848
transform 1 0 15204 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_21
timestamp 1754861848
transform 1 0 13608 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_22
timestamp 1754861848
transform 1 0 15708 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_23
timestamp 1754861848
transform 1 0 13692 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_24
timestamp 1754861848
transform 1 0 14952 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_25
timestamp 1754861848
transform 1 0 12768 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_26
timestamp 1754861848
transform 1 0 14616 0 1 9888
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_27
timestamp 1754861848
transform 1 0 14700 0 1 10272
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_28
timestamp 1754861848
transform 1 0 15288 0 1 11808
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_29
timestamp 1754861848
transform 1 0 15540 0 1 11904
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_30
timestamp 1754861848
transform 1 0 13188 0 1 10464
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_31
timestamp 1754861848
transform 1 0 14532 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_32
timestamp 1754861848
transform 1 0 12852 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_33
timestamp 1754861848
transform 1 0 14784 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_34
timestamp 1754861848
transform 1 0 14280 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_35
timestamp 1754861848
transform 1 0 14112 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_36
timestamp 1754861848
transform 1 0 13272 0 1 10272
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_37
timestamp 1754861848
transform 1 0 14112 0 1 11232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_38
timestamp 1754861848
transform 1 0 14700 0 1 11232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_39
timestamp 1754861848
transform 1 0 12768 0 1 10464
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_40
timestamp 1754861848
transform 1 0 15540 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_41
timestamp 1754861848
transform 1 0 14196 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_42
timestamp 1754861848
transform 1 0 13860 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_43
timestamp 1754861848
transform 1 0 14028 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_44
timestamp 1754861848
transform 1 0 14616 0 1 12384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_45
timestamp 1754861848
transform 1 0 15456 0 1 10464
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_46
timestamp 1754861848
transform 1 0 15204 0 1 11232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_47
timestamp 1754861848
transform 1 0 13356 0 1 11808
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_48
timestamp 1754861848
transform 1 0 15036 0 1 12000
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_49
timestamp 1754861848
transform 1 0 12936 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_50
timestamp 1754861848
transform 1 0 13608 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_51
timestamp 1754861848
transform 1 0 14868 0 1 11424
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_52
timestamp 1754861848
transform 1 0 15624 0 1 11424
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_53
timestamp 1754861848
transform 1 0 12852 0 1 11424
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_54
timestamp 1754861848
transform 1 0 12852 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_55
timestamp 1754861848
transform 1 0 13944 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_56
timestamp 1754861848
transform 1 0 15456 0 1 12000
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_57
timestamp 1754861848
transform 1 0 14952 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_58
timestamp 1754861848
transform 1 0 18732 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_59
timestamp 1754861848
transform 1 0 17640 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_60
timestamp 1754861848
transform 1 0 16380 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_61
timestamp 1754861848
transform 1 0 17892 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_62
timestamp 1754861848
transform 1 0 16296 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_63
timestamp 1754861848
transform 1 0 17808 0 1 10752
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_64
timestamp 1754861848
transform 1 0 16716 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_65
timestamp 1754861848
transform 1 0 17724 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_66
timestamp 1754861848
transform 1 0 18144 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_67
timestamp 1754861848
transform 1 0 17724 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_68
timestamp 1754861848
transform 1 0 18060 0 1 12384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_69
timestamp 1754861848
transform 1 0 18228 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_70
timestamp 1754861848
transform 1 0 18060 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_71
timestamp 1754861848
transform 1 0 18900 0 1 10368
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_72
timestamp 1754861848
transform 1 0 17340 0 1 10368
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_73
timestamp 1754861848
transform 1 0 16968 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_74
timestamp 1754861848
transform 1 0 17976 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_75
timestamp 1754861848
transform 1 0 18396 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_76
timestamp 1754861848
transform 1 0 18396 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_77
timestamp 1754861848
transform 1 0 17556 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_78
timestamp 1754861848
transform 1 0 18648 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_79
timestamp 1754861848
transform 1 0 16128 0 1 12672
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_80
timestamp 1754861848
transform 1 0 18984 0 1 10848
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_81
timestamp 1754861848
transform 1 0 17220 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_82
timestamp 1754861848
transform 1 0 16548 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_83
timestamp 1754861848
transform 1 0 15876 0 1 11232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_84
timestamp 1754861848
transform 1 0 22008 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_85
timestamp 1754861848
transform 1 0 21672 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_86
timestamp 1754861848
transform 1 0 19992 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_87
timestamp 1754861848
transform 1 0 19404 0 1 12288
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_88
timestamp 1754861848
transform 1 0 20328 0 1 12288
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_89
timestamp 1754861848
transform 1 0 20832 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_90
timestamp 1754861848
transform 1 0 19320 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_91
timestamp 1754861848
transform 1 0 21336 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_92
timestamp 1754861848
transform 1 0 19824 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_93
timestamp 1754861848
transform 1 0 19572 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_94
timestamp 1754861848
transform 1 0 21203 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_95
timestamp 1754861848
transform 1 0 21000 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_96
timestamp 1754861848
transform 1 0 20664 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_97
timestamp 1754861848
transform 1 0 19152 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_98
timestamp 1754861848
transform 1 0 21504 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_99
timestamp 1754861848
transform 1 0 20160 0 1 12672
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_100
timestamp 1754861848
transform 1 0 19992 0 1 10848
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_101
timestamp 1754861848
transform 1 0 20832 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_102
timestamp 1754861848
transform 1 0 21107 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_103
timestamp 1754861848
transform 1 0 19068 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_104
timestamp 1754861848
transform 1 0 19068 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_105
timestamp 1754861848
transform 1 0 7003 0 1 6432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_106
timestamp 1754861848
transform 1 0 7728 0 1 6432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_107
timestamp 1754861848
transform 1 0 6972 0 1 6624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_108
timestamp 1754861848
transform 1 0 7476 0 1 6624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_109
timestamp 1754861848
transform 1 0 7224 0 1 6624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_110
timestamp 1754861848
transform 1 0 10332 0 1 6336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_111
timestamp 1754861848
transform 1 0 7224 0 1 6336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_112
timestamp 1754861848
transform 1 0 5796 0 1 6624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_113
timestamp 1754861848
transform 1 0 4979 0 1 6432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_114
timestamp 1754861848
transform 1 0 4032 0 1 6432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_115
timestamp 1754861848
transform 1 0 5628 0 1 6432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_116
timestamp 1754861848
transform 1 0 5964 0 1 9696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_117
timestamp 1754861848
transform 1 0 4872 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_118
timestamp 1754861848
transform 1 0 4494 0 1 6912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_119
timestamp 1754861848
transform 1 0 5712 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_120
timestamp 1754861848
transform 1 0 4956 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_121
timestamp 1754861848
transform 1 0 4494 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_122
timestamp 1754861848
transform 1 0 4788 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_123
timestamp 1754861848
transform 1 0 4032 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_124
timestamp 1754861848
transform 1 0 5712 0 1 6912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_125
timestamp 1754861848
transform 1 0 5292 0 1 8832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_126
timestamp 1754861848
transform 1 0 5796 0 1 9696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_127
timestamp 1754861848
transform 1 0 6048 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_128
timestamp 1754861848
transform 1 0 5376 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_129
timestamp 1754861848
transform 1 0 5460 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_130
timestamp 1754861848
transform 1 0 3948 0 1 8448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_131
timestamp 1754861848
transform 1 0 6268 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_132
timestamp 1754861848
transform 1 0 6244 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_133
timestamp 1754861848
transform 1 0 5796 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_134
timestamp 1754861848
transform 1 0 4704 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_135
timestamp 1754861848
transform 1 0 4536 0 1 8448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_136
timestamp 1754861848
transform 1 0 5208 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_137
timestamp 1754861848
transform 1 0 4998 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_138
timestamp 1754861848
transform 1 0 5574 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_139
timestamp 1754861848
transform 1 0 5796 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_140
timestamp 1754861848
transform 1 0 5460 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_141
timestamp 1754861848
transform 1 0 5964 0 1 12576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_142
timestamp 1754861848
transform 1 0 4872 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_143
timestamp 1754861848
transform 1 0 5460 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_144
timestamp 1754861848
transform 1 0 5460 0 1 12288
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_145
timestamp 1754861848
transform 1 0 5460 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_146
timestamp 1754861848
transform 1 0 5880 0 1 12672
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_147
timestamp 1754861848
transform 1 0 5796 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_148
timestamp 1754861848
transform 1 0 6132 0 1 12096
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_149
timestamp 1754861848
transform 1 0 5964 0 1 11808
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_150
timestamp 1754861848
transform 1 0 6048 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_151
timestamp 1754861848
transform 1 0 6048 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_152
timestamp 1754861848
transform 1 0 4536 0 1 12000
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_153
timestamp 1754861848
transform 1 0 5754 0 1 11904
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_154
timestamp 1754861848
transform 1 0 5544 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_155
timestamp 1754861848
transform 1 0 4410 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_156
timestamp 1754861848
transform 1 0 10248 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_157
timestamp 1754861848
transform 1 0 11424 0 1 7008
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_158
timestamp 1754861848
transform 1 0 11172 0 1 7776
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_159
timestamp 1754861848
transform 1 0 10164 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_160
timestamp 1754861848
transform 1 0 10080 0 1 7104
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_161
timestamp 1754861848
transform 1 0 10752 0 1 7104
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_162
timestamp 1754861848
transform 1 0 11424 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_163
timestamp 1754861848
transform 1 0 12684 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_164
timestamp 1754861848
transform 1 0 9744 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_165
timestamp 1754861848
transform 1 0 12012 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_166
timestamp 1754861848
transform 1 0 11928 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_167
timestamp 1754861848
transform 1 0 12390 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_168
timestamp 1754861848
transform 1 0 11424 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_169
timestamp 1754861848
transform 1 0 9744 0 1 8256
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_170
timestamp 1754861848
transform 1 0 10206 0 1 8256
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_171
timestamp 1754861848
transform 1 0 11256 0 1 7872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_172
timestamp 1754861848
transform 1 0 9912 0 1 8448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_173
timestamp 1754861848
transform 1 0 9828 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_174
timestamp 1754861848
transform 1 0 11256 0 1 9312
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_175
timestamp 1754861848
transform 1 0 11928 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_176
timestamp 1754861848
transform 1 0 12684 0 1 9216
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_177
timestamp 1754861848
transform 1 0 11634 0 1 8448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_178
timestamp 1754861848
transform 1 0 9912 0 1 8832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_179
timestamp 1754861848
transform 1 0 9996 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_180
timestamp 1754861848
transform 1 0 11508 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_181
timestamp 1754861848
transform 1 0 10332 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_182
timestamp 1754861848
transform 1 0 11508 0 1 7776
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_183
timestamp 1754861848
transform 1 0 12558 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_184
timestamp 1754861848
transform 1 0 10416 0 1 6816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_185
timestamp 1754861848
transform 1 0 11088 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_186
timestamp 1754861848
transform 1 0 12264 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_187
timestamp 1754861848
transform 1 0 8652 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_188
timestamp 1754861848
transform 1 0 7224 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_189
timestamp 1754861848
transform 1 0 7896 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_190
timestamp 1754861848
transform 1 0 7224 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_191
timestamp 1754861848
transform 1 0 7392 0 1 9408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_192
timestamp 1754861848
transform 1 0 6468 0 1 9408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_193
timestamp 1754861848
transform 1 0 7560 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_194
timestamp 1754861848
transform 1 0 7056 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_195
timestamp 1754861848
transform 1 0 8316 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_196
timestamp 1754861848
transform 1 0 8820 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_197
timestamp 1754861848
transform 1 0 8232 0 1 8544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_198
timestamp 1754861848
transform 1 0 6888 0 1 9024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_199
timestamp 1754861848
transform 1 0 6888 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_200
timestamp 1754861848
transform 1 0 8652 0 1 9024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_201
timestamp 1754861848
transform 1 0 7224 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_202
timestamp 1754861848
transform 1 0 6720 0 1 8832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_203
timestamp 1754861848
transform 1 0 7392 0 1 8832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_204
timestamp 1754861848
transform 1 0 8484 0 1 6816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_205
timestamp 1754861848
transform 1 0 7477 0 1 6816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_206
timestamp 1754861848
transform 1 0 9324 0 1 8832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_207
timestamp 1754861848
transform 1 0 9408 0 1 6816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_208
timestamp 1754861848
transform 1 0 7056 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_209
timestamp 1754861848
transform 1 0 9156 0 1 7968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_210
timestamp 1754861848
transform 1 0 9072 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_211
timestamp 1754861848
transform 1 0 8316 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_212
timestamp 1754861848
transform 1 0 9324 0 1 7104
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_213
timestamp 1754861848
transform 1 0 6888 0 1 8640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_214
timestamp 1754861848
transform 1 0 8568 0 1 7200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_215
timestamp 1754861848
transform 1 0 6804 0 1 9600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_216
timestamp 1754861848
transform 1 0 8232 0 1 8928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_217
timestamp 1754861848
transform 1 0 7812 0 1 9312
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_218
timestamp 1754861848
transform 1 0 7560 0 1 9312
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_219
timestamp 1754861848
transform 1 0 8400 0 1 8736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_220
timestamp 1754861848
transform 1 0 8437 0 1 7872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_221
timestamp 1754861848
transform 1 0 6720 0 1 9312
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_222
timestamp 1754861848
transform 1 0 8988 0 1 9504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_223
timestamp 1754861848
transform 1 0 9030 0 1 12576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_224
timestamp 1754861848
transform 1 0 8636 0 1 12192
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_225
timestamp 1754861848
transform 1 0 8820 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_226
timestamp 1754861848
transform 1 0 7098 0 1 12576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_227
timestamp 1754861848
transform 1 0 6972 0 1 12288
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_228
timestamp 1754861848
transform 1 0 9324 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_229
timestamp 1754861848
transform 1 0 7392 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_230
timestamp 1754861848
transform 1 0 7392 0 1 12288
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_231
timestamp 1754861848
transform 1 0 8148 0 1 9888
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_232
timestamp 1754861848
transform 1 0 8263 0 1 11040
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_233
timestamp 1754861848
transform 1 0 7644 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_234
timestamp 1754861848
transform 1 0 9198 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_235
timestamp 1754861848
transform 1 0 8904 0 1 9888
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_236
timestamp 1754861848
transform 1 0 9408 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_237
timestamp 1754861848
transform 1 0 7086 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_238
timestamp 1754861848
transform 1 0 6636 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_239
timestamp 1754861848
transform 1 0 6552 0 1 12384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_240
timestamp 1754861848
transform 1 0 7728 0 1 11904
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_241
timestamp 1754861848
transform 1 0 6720 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_242
timestamp 1754861848
transform 1 0 9102 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_243
timestamp 1754861848
transform 1 0 9156 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_244
timestamp 1754861848
transform 1 0 8148 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_245
timestamp 1754861848
transform 1 0 8148 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_246
timestamp 1754861848
transform 1 0 7476 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_247
timestamp 1754861848
transform 1 0 7392 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_248
timestamp 1754861848
transform 1 0 6804 0 1 9984
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_249
timestamp 1754861848
transform 1 0 8064 0 1 12000
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_250
timestamp 1754861848
transform 1 0 8484 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_251
timestamp 1754861848
transform 1 0 8652 0 1 11712
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_252
timestamp 1754861848
transform 1 0 6972 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_253
timestamp 1754861848
transform 1 0 7140 0 1 12768
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_254
timestamp 1754861848
transform 1 0 7560 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_255
timestamp 1754861848
transform 1 0 8988 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_256
timestamp 1754861848
transform 1 0 7980 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_257
timestamp 1754861848
transform 1 0 9912 0 1 12576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_258
timestamp 1754861848
transform 1 0 10458 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_259
timestamp 1754861848
transform 1 0 12684 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_260
timestamp 1754861848
transform 1 0 10374 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_261
timestamp 1754861848
transform 1 0 12348 0 1 10176
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_262
timestamp 1754861848
transform 1 0 10584 0 1 10752
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_263
timestamp 1754861848
transform 1 0 10752 0 1 11040
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_264
timestamp 1754861848
transform 1 0 11844 0 1 12384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_265
timestamp 1754861848
transform 1 0 9599 0 1 12672
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_266
timestamp 1754861848
transform 1 0 12390 0 1 11616
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_267
timestamp 1754861848
transform 1 0 12180 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_268
timestamp 1754861848
transform 1 0 12180 0 1 10464
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_269
timestamp 1754861848
transform 1 0 11676 0 1 10272
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_270
timestamp 1754861848
transform 1 0 10164 0 1 10080
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_271
timestamp 1754861848
transform 1 0 12348 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_272
timestamp 1754861848
transform 1 0 10080 0 1 10656
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_273
timestamp 1754861848
transform 1 0 11172 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_274
timestamp 1754861848
transform 1 0 11592 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_275
timestamp 1754861848
transform 1 0 11256 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_276
timestamp 1754861848
transform 1 0 11256 0 1 11520
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_277
timestamp 1754861848
transform 1 0 11004 0 1 10944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_278
timestamp 1754861848
transform 1 0 11172 0 1 10272
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_279
timestamp 1754861848
transform 1 0 9912 0 1 10272
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_280
timestamp 1754861848
transform 1 0 12180 0 1 11904
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_281
timestamp 1754861848
transform 1 0 9576 0 1 11136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_282
timestamp 1754861848
transform 1 0 9576 0 1 7872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_283
timestamp 1754861848
transform 1 0 8652 0 1 9792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_284
timestamp 1754861848
transform 1 0 9576 0 1 10656
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_285
timestamp 1754861848
transform 1 0 6384 0 1 9792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_286
timestamp 1754861848
transform 1 0 6384 0 1 12480
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_287
timestamp 1754861848
transform 1 0 11508 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_288
timestamp 1754861848
transform 1 0 10920 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_289
timestamp 1754861848
transform 1 0 12264 0 1 13632
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_290
timestamp 1754861848
transform 1 0 12096 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_291
timestamp 1754861848
transform 1 0 11508 0 1 13632
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_292
timestamp 1754861848
transform 1 0 11424 0 1 13728
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_293
timestamp 1754861848
transform 1 0 11256 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_294
timestamp 1754861848
transform 1 0 11172 0 1 13728
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_295
timestamp 1754861848
transform 1 0 10920 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_296
timestamp 1754861848
transform 1 0 10164 0 1 14592
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_297
timestamp 1754861848
transform 1 0 12348 0 1 13536
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_298
timestamp 1754861848
transform 1 0 12348 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_299
timestamp 1754861848
transform 1 0 9996 0 1 14976
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_300
timestamp 1754861848
transform 1 0 10584 0 1 14976
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_301
timestamp 1754861848
transform 1 0 10668 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_302
timestamp 1754861848
transform 1 0 11844 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_303
timestamp 1754861848
transform 1 0 12474 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_304
timestamp 1754861848
transform 1 0 11424 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_305
timestamp 1754861848
transform 1 0 10332 0 1 12960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_306
timestamp 1754861848
transform 1 0 11844 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_307
timestamp 1754861848
transform 1 0 10584 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_308
timestamp 1754861848
transform 1 0 10836 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_309
timestamp 1754861848
transform 1 0 10584 0 1 12960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_310
timestamp 1754861848
transform 1 0 12516 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_311
timestamp 1754861848
transform 1 0 12012 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_312
timestamp 1754861848
transform 1 0 12348 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_313
timestamp 1754861848
transform 1 0 10164 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_314
timestamp 1754861848
transform 1 0 10920 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_315
timestamp 1754861848
transform 1 0 12348 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_316
timestamp 1754861848
transform 1 0 12600 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_317
timestamp 1754861848
transform 1 0 10752 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_318
timestamp 1754861848
transform 1 0 11424 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_319
timestamp 1754861848
transform 1 0 12096 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_320
timestamp 1754861848
transform 1 0 12672 0 1 15744
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_321
timestamp 1754861848
transform 1 0 12390 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_322
timestamp 1754861848
transform 1 0 9492 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_323
timestamp 1754861848
transform 1 0 8820 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_324
timestamp 1754861848
transform 1 0 8442 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_325
timestamp 1754861848
transform 1 0 8400 0 1 14592
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_326
timestamp 1754861848
transform 1 0 8358 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_327
timestamp 1754861848
transform 1 0 6636 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_328
timestamp 1754861848
transform 1 0 8904 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_329
timestamp 1754861848
transform 1 0 8484 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_330
timestamp 1754861848
transform 1 0 6804 0 1 14976
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_331
timestamp 1754861848
transform 1 0 6804 0 1 12960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_332
timestamp 1754861848
transform 1 0 8568 0 1 13344
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_333
timestamp 1754861848
transform 1 0 6594 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_334
timestamp 1754861848
transform 1 0 7140 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_335
timestamp 1754861848
transform 1 0 6720 0 1 15744
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_336
timestamp 1754861848
transform 1 0 7476 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_337
timestamp 1754861848
transform 1 0 8652 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_338
timestamp 1754861848
transform 1 0 7896 0 1 13536
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_339
timestamp 1754861848
transform 1 0 7224 0 1 15936
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_340
timestamp 1754861848
transform 1 0 7896 0 1 15936
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_341
timestamp 1754861848
transform 1 0 7644 0 1 15744
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_342
timestamp 1754861848
transform 1 0 8988 0 1 13248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_343
timestamp 1754861848
transform 1 0 6720 0 1 13344
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_344
timestamp 1754861848
transform 1 0 9156 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_345
timestamp 1754861848
transform 1 0 7728 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_346
timestamp 1754861848
transform 1 0 9408 0 1 16512
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_347
timestamp 1754861848
transform 1 0 8904 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_348
timestamp 1754861848
transform 1 0 8548 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_349
timestamp 1754861848
transform 1 0 8736 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_350
timestamp 1754861848
transform 1 0 6720 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_351
timestamp 1754861848
transform 1 0 6468 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_352
timestamp 1754861848
transform 1 0 9324 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_353
timestamp 1754861848
transform 1 0 6804 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_354
timestamp 1754861848
transform 1 0 8568 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_355
timestamp 1754861848
transform 1 0 9240 0 1 16320
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_356
timestamp 1754861848
transform 1 0 7644 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_357
timestamp 1754861848
transform 1 0 8988 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_358
timestamp 1754861848
transform 1 0 8988 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_359
timestamp 1754861848
transform 1 0 8652 0 1 18912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_360
timestamp 1754861848
transform 1 0 8064 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_361
timestamp 1754861848
transform 1 0 9492 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_362
timestamp 1754861848
transform 1 0 9492 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_363
timestamp 1754861848
transform 1 0 9240 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_364
timestamp 1754861848
transform 1 0 7896 0 1 16128
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_365
timestamp 1754861848
transform 1 0 6804 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_366
timestamp 1754861848
transform 1 0 8064 0 1 17376
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_367
timestamp 1754861848
transform 1 0 9240 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_368
timestamp 1754861848
transform 1 0 6720 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_369
timestamp 1754861848
transform 1 0 7140 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_370
timestamp 1754861848
transform 1 0 7224 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_371
timestamp 1754861848
transform 1 0 7224 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_372
timestamp 1754861848
transform 1 0 9240 0 1 19008
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_373
timestamp 1754861848
transform 1 0 11760 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_374
timestamp 1754861848
transform 1 0 12264 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_375
timestamp 1754861848
transform 1 0 12012 0 1 18336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_376
timestamp 1754861848
transform 1 0 11256 0 1 18336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_377
timestamp 1754861848
transform 1 0 11508 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_378
timestamp 1754861848
transform 1 0 10374 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_379
timestamp 1754861848
transform 1 0 10836 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_380
timestamp 1754861848
transform 1 0 9996 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_381
timestamp 1754861848
transform 1 0 11676 0 1 16128
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_382
timestamp 1754861848
transform 1 0 9744 0 1 19008
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_383
timestamp 1754861848
transform 1 0 10836 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_384
timestamp 1754861848
transform 1 0 11172 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_385
timestamp 1754861848
transform 1 0 9912 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_386
timestamp 1754861848
transform 1 0 10500 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_387
timestamp 1754861848
transform 1 0 11088 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_388
timestamp 1754861848
transform 1 0 10416 0 1 17568
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_389
timestamp 1754861848
transform 1 0 10668 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_390
timestamp 1754861848
transform 1 0 9828 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_391
timestamp 1754861848
transform 1 0 9828 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_392
timestamp 1754861848
transform 1 0 12180 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_393
timestamp 1754861848
transform 1 0 10500 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_394
timestamp 1754861848
transform 1 0 11172 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_395
timestamp 1754861848
transform 1 0 10920 0 1 17184
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_396
timestamp 1754861848
transform 1 0 11424 0 1 17184
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_397
timestamp 1754861848
transform 1 0 9996 0 1 16320
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_398
timestamp 1754861848
transform 1 0 11298 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_399
timestamp 1754861848
transform 1 0 11676 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_400
timestamp 1754861848
transform 1 0 10080 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_401
timestamp 1754861848
transform 1 0 11802 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_402
timestamp 1754861848
transform 1 0 11004 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_403
timestamp 1754861848
transform 1 0 11676 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_404
timestamp 1754861848
transform 1 0 10248 0 1 18912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_405
timestamp 1754861848
transform 1 0 11088 0 1 16032
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_406
timestamp 1754861848
transform 1 0 10080 0 1 16032
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_407
timestamp 1754861848
transform 1 0 9642 0 1 17568
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_408
timestamp 1754861848
transform 1 0 10416 0 1 16416
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_409
timestamp 1754861848
transform 1 0 10248 0 1 16608
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_410
timestamp 1754861848
transform 1 0 10668 0 1 16128
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_411
timestamp 1754861848
transform 1 0 10164 0 1 17952
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_412
timestamp 1754861848
transform 1 0 11508 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_413
timestamp 1754861848
transform 1 0 10920 0 1 18240
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_414
timestamp 1754861848
transform 1 0 11004 0 1 16704
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_415
timestamp 1754861848
transform 1 0 12096 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_416
timestamp 1754861848
transform 1 0 11256 0 1 16416
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_417
timestamp 1754861848
transform 1 0 10752 0 1 16512
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_418
timestamp 1754861848
transform 1 0 10584 0 1 16416
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_419
timestamp 1754861848
transform 1 0 12264 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_420
timestamp 1754861848
transform 1 0 12684 0 1 17184
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_421
timestamp 1754861848
transform 1 0 11424 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_422
timestamp 1754861848
transform 1 0 6300 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_423
timestamp 1754861848
transform 1 0 4452 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_424
timestamp 1754861848
transform 1 0 6048 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_425
timestamp 1754861848
transform 1 0 5292 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_426
timestamp 1754861848
transform 1 0 4704 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_427
timestamp 1754861848
transform 1 0 5208 0 1 13344
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_428
timestamp 1754861848
transform 1 0 4704 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_429
timestamp 1754861848
transform 1 0 5544 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_430
timestamp 1754861848
transform 1 0 4536 0 1 15456
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_431
timestamp 1754861848
transform 1 0 5796 0 1 14400
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_432
timestamp 1754861848
transform 1 0 5796 0 1 15456
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_433
timestamp 1754861848
transform 1 0 4872 0 1 14400
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_434
timestamp 1754861848
transform 1 0 5796 0 1 13248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_435
timestamp 1754861848
transform 1 0 5376 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_436
timestamp 1754861848
transform 1 0 5148 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_437
timestamp 1754861848
transform 1 0 4788 0 1 13248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_438
timestamp 1754861848
transform 1 0 4620 0 1 13344
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_439
timestamp 1754861848
transform 1 0 6300 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_440
timestamp 1754861848
transform 1 0 6216 0 1 16320
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_441
timestamp 1754861848
transform 1 0 6300 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_442
timestamp 1754861848
transform 1 0 5964 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_443
timestamp 1754861848
transform 1 0 5166 0 1 17376
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_444
timestamp 1754861848
transform 1 0 6132 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_445
timestamp 1754861848
transform 1 0 5796 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_446
timestamp 1754861848
transform 1 0 5460 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_447
timestamp 1754861848
transform 1 0 4788 0 1 16704
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_448
timestamp 1754861848
transform 1 0 4872 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_449
timestamp 1754861848
transform 1 0 5796 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_450
timestamp 1754861848
transform 1 0 6048 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_451
timestamp 1754861848
transform 1 0 5916 0 1 16320
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_452
timestamp 1754861848
transform 1 0 5376 0 1 21696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_453
timestamp 1754861848
transform 1 0 5292 0 1 24192
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_454
timestamp 1754861848
transform 1 0 10836 0 1 20736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_455
timestamp 1754861848
transform 1 0 9912 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_456
timestamp 1754861848
transform 1 0 9912 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_457
timestamp 1754861848
transform 1 0 11130 0 1 21024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_458
timestamp 1754861848
transform 1 0 9744 0 1 20544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_459
timestamp 1754861848
transform 1 0 11256 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_460
timestamp 1754861848
transform 1 0 10584 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_461
timestamp 1754861848
transform 1 0 10584 0 1 20928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_462
timestamp 1754861848
transform 1 0 11340 0 1 19392
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_463
timestamp 1754861848
transform 1 0 12180 0 1 19200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_464
timestamp 1754861848
transform 1 0 12684 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_465
timestamp 1754861848
transform 1 0 11508 0 1 20832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_466
timestamp 1754861848
transform 1 0 11676 0 1 20832
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_467
timestamp 1754861848
transform 1 0 12180 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_468
timestamp 1754861848
transform 1 0 11172 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_469
timestamp 1754861848
transform 1 0 12096 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_470
timestamp 1754861848
transform 1 0 10332 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_471
timestamp 1754861848
transform 1 0 12516 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_472
timestamp 1754861848
transform 1 0 9705 0 1 21696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_473
timestamp 1754861848
transform 1 0 10164 0 1 19680
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_474
timestamp 1754861848
transform 1 0 11256 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_475
timestamp 1754861848
transform 1 0 12012 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_476
timestamp 1754861848
transform 1 0 6888 0 1 20544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_477
timestamp 1754861848
transform 1 0 8484 0 1 20544
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_478
timestamp 1754861848
transform 1 0 6804 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_479
timestamp 1754861848
transform 1 0 7308 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_480
timestamp 1754861848
transform 1 0 8820 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_481
timestamp 1754861848
transform 1 0 8148 0 1 20256
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_482
timestamp 1754861848
transform 1 0 7896 0 1 20256
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_483
timestamp 1754861848
transform 1 0 8232 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_484
timestamp 1754861848
transform 1 0 8736 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_485
timestamp 1754861848
transform 1 0 9324 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_486
timestamp 1754861848
transform 1 0 8064 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_487
timestamp 1754861848
transform 1 0 8988 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_488
timestamp 1754861848
transform 1 0 8904 0 1 19776
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_489
timestamp 1754861848
transform 1 0 6636 0 1 20736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_490
timestamp 1754861848
transform 1 0 6888 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_491
timestamp 1754861848
transform 1 0 8736 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_492
timestamp 1754861848
transform 1 0 9198 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_493
timestamp 1754861848
transform 1 0 9408 0 1 19392
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_494
timestamp 1754861848
transform 1 0 8652 0 1 19392
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_495
timestamp 1754861848
transform 1 0 8820 0 1 19200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_496
timestamp 1754861848
transform 1 0 7182 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_497
timestamp 1754861848
transform 1 0 7056 0 1 19968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_498
timestamp 1754861848
transform 1 0 8652 0 1 21408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_499
timestamp 1754861848
transform 1 0 9492 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_500
timestamp 1754861848
transform 1 0 6972 0 1 19584
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_501
timestamp 1754861848
transform 1 0 7308 0 1 20640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_502
timestamp 1754861848
transform 1 0 7476 0 1 20640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_503
timestamp 1754861848
transform 1 0 9072 0 1 23424
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_504
timestamp 1754861848
transform 1 0 6468 0 1 24864
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_505
timestamp 1754861848
transform 1 0 6972 0 1 24576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_506
timestamp 1754861848
transform 1 0 7392 0 1 25248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_507
timestamp 1754861848
transform 1 0 8568 0 1 25152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_508
timestamp 1754861848
transform 1 0 11760 0 1 25056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_509
timestamp 1754861848
transform 1 0 11844 0 1 22944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_510
timestamp 1754861848
transform 1 0 10416 0 1 22944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_511
timestamp 1754861848
transform 1 0 10836 0 1 24192
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_512
timestamp 1754861848
transform 1 0 12096 0 1 24384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_513
timestamp 1754861848
transform 1 0 9576 0 1 21696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_514
timestamp 1754861848
transform 1 0 6384 0 1 15744
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_515
timestamp 1754861848
transform 1 0 6384 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_516
timestamp 1754861848
transform 1 0 6384 0 1 24384
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_517
timestamp 1754861848
transform 1 0 21672 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_518
timestamp 1754861848
transform 1 0 20328 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_519
timestamp 1754861848
transform 1 0 20664 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_520
timestamp 1754861848
transform 1 0 20412 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_521
timestamp 1754861848
transform 1 0 21798 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_522
timestamp 1754861848
transform 1 0 20916 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_523
timestamp 1754861848
transform 1 0 19908 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_524
timestamp 1754861848
transform 1 0 19488 0 1 13920
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_525
timestamp 1754861848
transform 1 0 21924 0 1 13920
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_526
timestamp 1754861848
transform 1 0 20916 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_527
timestamp 1754861848
transform 1 0 19572 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_528
timestamp 1754861848
transform 1 0 21924 0 1 15264
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_529
timestamp 1754861848
transform 1 0 20748 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_530
timestamp 1754861848
transform 1 0 21504 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_531
timestamp 1754861848
transform 1 0 19236 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_532
timestamp 1754861848
transform 1 0 20244 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_533
timestamp 1754861848
transform 1 0 20916 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_534
timestamp 1754861848
transform 1 0 19488 0 1 18336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_535
timestamp 1754861848
transform 1 0 20748 0 1 16032
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_536
timestamp 1754861848
transform 1 0 21588 0 1 16032
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_537
timestamp 1754861848
transform 1 0 19740 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_538
timestamp 1754861848
transform 1 0 20034 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_539
timestamp 1754861848
transform 1 0 19404 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_540
timestamp 1754861848
transform 1 0 19859 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_541
timestamp 1754861848
transform 1 0 19488 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_542
timestamp 1754861848
transform 1 0 20160 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_543
timestamp 1754861848
transform 1 0 19488 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_544
timestamp 1754861848
transform 1 0 20412 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_545
timestamp 1754861848
transform 1 0 17220 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_546
timestamp 1754861848
transform 1 0 16548 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_547
timestamp 1754861848
transform 1 0 17472 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_548
timestamp 1754861848
transform 1 0 18816 0 1 14784
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_549
timestamp 1754861848
transform 1 0 18522 0 1 14784
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_550
timestamp 1754861848
transform 1 0 18816 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_551
timestamp 1754861848
transform 1 0 17892 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_552
timestamp 1754861848
transform 1 0 17839 0 1 13728
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_553
timestamp 1754861848
transform 1 0 18144 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_554
timestamp 1754861848
transform 1 0 18690 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_555
timestamp 1754861848
transform 1 0 17388 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_556
timestamp 1754861848
transform 1 0 16254 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_557
timestamp 1754861848
transform 1 0 18228 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_558
timestamp 1754861848
transform 1 0 17892 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_559
timestamp 1754861848
transform 1 0 17388 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_560
timestamp 1754861848
transform 1 0 17388 0 1 13920
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_561
timestamp 1754861848
transform 1 0 18396 0 1 15264
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_562
timestamp 1754861848
transform 1 0 18564 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_563
timestamp 1754861848
transform 1 0 16044 0 1 12960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_564
timestamp 1754861848
transform 1 0 16716 0 1 15456
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_565
timestamp 1754861848
transform 1 0 18060 0 1 15456
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_566
timestamp 1754861848
transform 1 0 18732 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_567
timestamp 1754861848
transform 1 0 16884 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_568
timestamp 1754861848
transform 1 0 17556 0 1 14496
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_569
timestamp 1754861848
transform 1 0 17766 0 1 14496
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_570
timestamp 1754861848
transform 1 0 16128 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_571
timestamp 1754861848
transform 1 0 18228 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_572
timestamp 1754861848
transform 1 0 16632 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_573
timestamp 1754861848
transform 1 0 18522 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_574
timestamp 1754861848
transform 1 0 17556 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_575
timestamp 1754861848
transform 1 0 16128 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_576
timestamp 1754861848
transform 1 0 16044 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_577
timestamp 1754861848
transform 1 0 15204 0 1 14496
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_578
timestamp 1754861848
transform 1 0 13734 0 1 15264
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_579
timestamp 1754861848
transform 1 0 15036 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_580
timestamp 1754861848
transform 1 0 15036 0 1 14496
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_581
timestamp 1754861848
transform 1 0 13146 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_582
timestamp 1754861848
transform 1 0 13860 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_583
timestamp 1754861848
transform 1 0 14868 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_584
timestamp 1754861848
transform 1 0 15456 0 1 14208
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_585
timestamp 1754861848
transform 1 0 13944 0 1 15744
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_586
timestamp 1754861848
transform 1 0 13860 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_587
timestamp 1754861848
transform 1 0 15624 0 1 15264
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_588
timestamp 1754861848
transform 1 0 13356 0 1 13440
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_589
timestamp 1754861848
transform 1 0 13608 0 1 13920
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_590
timestamp 1754861848
transform 1 0 12936 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_591
timestamp 1754861848
transform 1 0 15036 0 1 15456
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_592
timestamp 1754861848
transform 1 0 15456 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_593
timestamp 1754861848
transform 1 0 13524 0 1 13248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_594
timestamp 1754861848
transform 1 0 15624 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_595
timestamp 1754861848
transform 1 0 14952 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_596
timestamp 1754861848
transform 1 0 15624 0 1 15840
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_597
timestamp 1754861848
transform 1 0 14364 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_598
timestamp 1754861848
transform 1 0 14952 0 1 14112
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_599
timestamp 1754861848
transform 1 0 12852 0 1 15648
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_600
timestamp 1754861848
transform 1 0 13272 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_601
timestamp 1754861848
transform 1 0 14280 0 1 13152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_602
timestamp 1754861848
transform 1 0 15708 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_603
timestamp 1754861848
transform 1 0 15372 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_604
timestamp 1754861848
transform 1 0 15708 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_605
timestamp 1754861848
transform 1 0 15708 0 1 13344
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_606
timestamp 1754861848
transform 1 0 14616 0 1 13728
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_607
timestamp 1754861848
transform 1 0 15540 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_608
timestamp 1754861848
transform 1 0 12768 0 1 12960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_609
timestamp 1754861848
transform 1 0 14409 0 1 15552
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_610
timestamp 1754861848
transform 1 0 15120 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_611
timestamp 1754861848
transform 1 0 14028 0 1 14688
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_612
timestamp 1754861848
transform 1 0 14028 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_613
timestamp 1754861848
transform 1 0 14364 0 1 13056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_614
timestamp 1754861848
transform 1 0 14490 0 1 14016
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_615
timestamp 1754861848
transform 1 0 14490 0 1 13824
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_616
timestamp 1754861848
transform 1 0 15834 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_617
timestamp 1754861848
transform 1 0 15204 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_618
timestamp 1754861848
transform 1 0 12936 0 1 16224
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_619
timestamp 1754861848
transform 1 0 14784 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_620
timestamp 1754861848
transform 1 0 14700 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_621
timestamp 1754861848
transform 1 0 13188 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_622
timestamp 1754861848
transform 1 0 13188 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_623
timestamp 1754861848
transform 1 0 13776 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_624
timestamp 1754861848
transform 1 0 15288 0 1 18432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_625
timestamp 1754861848
transform 1 0 13524 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_626
timestamp 1754861848
transform 1 0 14490 0 1 16800
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_627
timestamp 1754861848
transform 1 0 14112 0 1 17952
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_628
timestamp 1754861848
transform 1 0 14784 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_629
timestamp 1754861848
transform 1 0 15036 0 1 17664
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_630
timestamp 1754861848
transform 1 0 12768 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_631
timestamp 1754861848
transform 1 0 13440 0 1 17952
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_632
timestamp 1754861848
transform 1 0 14364 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_633
timestamp 1754861848
transform 1 0 13608 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_634
timestamp 1754861848
transform 1 0 13146 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_635
timestamp 1754861848
transform 1 0 13356 0 1 16128
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_636
timestamp 1754861848
transform 1 0 13272 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_637
timestamp 1754861848
transform 1 0 14196 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_638
timestamp 1754861848
transform 1 0 15708 0 1 17184
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_639
timestamp 1754861848
transform 1 0 13020 0 1 17184
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_640
timestamp 1754861848
transform 1 0 16716 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_641
timestamp 1754861848
transform 1 0 17976 0 1 18720
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_642
timestamp 1754861848
transform 1 0 17472 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_643
timestamp 1754861848
transform 1 0 18228 0 1 18816
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_644
timestamp 1754861848
transform 1 0 16044 0 1 16896
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_645
timestamp 1754861848
transform 1 0 18312 0 1 18336
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_646
timestamp 1754861848
transform 1 0 18060 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_647
timestamp 1754861848
transform 1 0 18060 0 1 17568
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_648
timestamp 1754861848
transform 1 0 16380 0 1 17568
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_649
timestamp 1754861848
transform 1 0 17220 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_650
timestamp 1754861848
transform 1 0 16716 0 1 17088
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_651
timestamp 1754861848
transform 1 0 16548 0 1 18624
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_652
timestamp 1754861848
transform 1 0 17304 0 1 16992
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_653
timestamp 1754861848
transform 1 0 17640 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_654
timestamp 1754861848
transform 1 0 16044 0 1 17856
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_655
timestamp 1754861848
transform 1 0 17640 0 1 18528
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_656
timestamp 1754861848
transform 1 0 18144 0 1 18432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_657
timestamp 1754861848
transform 1 0 18564 0 1 18432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_658
timestamp 1754861848
transform 1 0 17724 0 1 18912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_659
timestamp 1754861848
transform 1 0 18060 0 1 18912
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_660
timestamp 1754861848
transform 1 0 17892 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_661
timestamp 1754861848
transform 1 0 16674 0 1 17760
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_662
timestamp 1754861848
transform 1 0 18228 0 1 17280
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_663
timestamp 1754861848
transform 1 0 16800 0 1 16416
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_664
timestamp 1754861848
transform 1 0 17220 0 1 16416
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_665
timestamp 1754861848
transform 1 0 15876 0 1 18432
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_666
timestamp 1754861848
transform 1 0 15876 0 1 14496
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_667
timestamp 1754861848
transform 1 0 15876 0 1 14304
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_668
timestamp 1754861848
transform 1 0 18648 0 1 19200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_669
timestamp 1754861848
transform 1 0 17766 0 1 20736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_670
timestamp 1754861848
transform 1 0 16716 0 1 20736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_671
timestamp 1754861848
transform 1 0 16884 0 1 21024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_672
timestamp 1754861848
transform 1 0 16212 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_673
timestamp 1754861848
transform 1 0 16548 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_674
timestamp 1754861848
transform 1 0 18564 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_675
timestamp 1754861848
transform 1 0 18060 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_676
timestamp 1754861848
transform 1 0 17094 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_677
timestamp 1754861848
transform 1 0 18312 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_678
timestamp 1754861848
transform 1 0 17850 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_679
timestamp 1754861848
transform 1 0 16632 0 1 21696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_680
timestamp 1754861848
transform 1 0 17472 0 1 21792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_681
timestamp 1754861848
transform 1 0 17136 0 1 21792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_682
timestamp 1754861848
transform 1 0 16128 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_683
timestamp 1754861848
transform 1 0 17640 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_684
timestamp 1754861848
transform 1 0 16800 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_685
timestamp 1754861848
transform 1 0 16128 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_686
timestamp 1754861848
transform 1 0 17304 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_687
timestamp 1754861848
transform 1 0 15960 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_688
timestamp 1754861848
transform 1 0 15960 0 1 19968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_689
timestamp 1754861848
transform 1 0 16212 0 1 19968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_690
timestamp 1754861848
transform 1 0 17839 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_691
timestamp 1754861848
transform 1 0 18396 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_692
timestamp 1754861848
transform 1 0 15740 0 1 19200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_693
timestamp 1754861848
transform 1 0 15151 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_694
timestamp 1754861848
transform 1 0 14700 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_695
timestamp 1754861848
transform 1 0 14784 0 1 20736
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_696
timestamp 1754861848
transform 1 0 14112 0 1 21024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_697
timestamp 1754861848
transform 1 0 13272 0 1 21024
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_698
timestamp 1754861848
transform 1 0 12852 0 1 20928
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_699
timestamp 1754861848
transform 1 0 15624 0 1 19200
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_700
timestamp 1754861848
transform 1 0 13608 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_701
timestamp 1754861848
transform 1 0 14784 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_702
timestamp 1754861848
transform 1 0 13944 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_703
timestamp 1754861848
transform 1 0 15708 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_704
timestamp 1754861848
transform 1 0 15540 0 1 21696
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_705
timestamp 1754861848
transform 1 0 14364 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_706
timestamp 1754861848
transform 1 0 14616 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_707
timestamp 1754861848
transform 1 0 14490 0 1 20640
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_708
timestamp 1754861848
transform 1 0 13440 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_709
timestamp 1754861848
transform 1 0 14868 0 1 19872
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_710
timestamp 1754861848
transform 1 0 14490 0 1 20448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_711
timestamp 1754861848
transform 1 0 14868 0 1 20448
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_712
timestamp 1754861848
transform 1 0 14658 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_713
timestamp 1754861848
transform 1 0 14448 0 1 20064
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_714
timestamp 1754861848
transform 1 0 13188 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_715
timestamp 1754861848
transform 1 0 14112 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_716
timestamp 1754861848
transform 1 0 13188 0 1 19680
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_717
timestamp 1754861848
transform 1 0 12768 0 1 19680
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_718
timestamp 1754861848
transform 1 0 13692 0 1 19968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_719
timestamp 1754861848
transform 1 0 14616 0 1 21792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_720
timestamp 1754861848
transform 1 0 13776 0 1 21792
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_721
timestamp 1754861848
transform 1 0 12768 0 1 19968
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_722
timestamp 1754861848
transform 1 0 14784 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_723
timestamp 1754861848
transform 1 0 13230 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_724
timestamp 1754861848
transform 1 0 14280 0 1 19488
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_725
timestamp 1754861848
transform 1 0 13440 0 1 24960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_726
timestamp 1754861848
transform 1 0 14616 0 1 23040
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_727
timestamp 1754861848
transform 1 0 18648 0 1 23232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_728
timestamp 1754861848
transform 1 0 18816 0 1 23136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_729
timestamp 1754861848
transform 1 0 17220 0 1 22944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_730
timestamp 1754861848
transform 1 0 18396 0 1 23040
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_731
timestamp 1754861848
transform 1 0 16296 0 1 23424
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_732
timestamp 1754861848
transform 1 0 15876 0 1 24864
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_733
timestamp 1754861848
transform 1 0 25116 0 1 23232
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_734
timestamp 1754861848
transform 1 0 24696 0 1 23136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_735
timestamp 1754861848
transform 1 0 20916 0 1 20160
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_736
timestamp 1754861848
transform 1 0 20496 0 1 21504
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_737
timestamp 1754861848
transform 1 0 20076 0 1 21600
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_738
timestamp 1754861848
transform 1 0 19572 0 1 21408
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_739
timestamp 1754861848
transform 1 0 19236 0 1 19392
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_740
timestamp 1754861848
transform 1 0 21756 0 1 23040
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_741
timestamp 1754861848
transform 1 0 19656 0 1 22944
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_742
timestamp 1754861848
transform 1 0 22176 0 1 24576
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_743
timestamp 1754861848
transform 1 0 24024 0 1 19296
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_744
timestamp 1754861848
transform 1 0 23436 0 1 25056
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_745
timestamp 1754861848
transform 1 0 20160 0 1 23136
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_746
timestamp 1754861848
transform 1 0 22596 0 1 25152
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_747
timestamp 1754861848
transform 1 0 23016 0 1 25248
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_748
timestamp 1754861848
transform 1 0 24276 0 1 24960
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_749
timestamp 1754861848
transform 1 0 14868 0 1 19104
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_750
timestamp 1754861848
transform 1 0 13944 0 1 19104
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_751
timestamp 1754861848
transform 1 0 18312 0 1 12864
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_752
timestamp 1754861848
transform 1 0 12180 0 1 12864
box -29 -29 29 29
use VIA_Via2_YX  VIA_Via2_YX_753
timestamp 1754861848
transform 1 0 8736 0 1 12864
box -29 -29 29 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_0
timestamp 1754861848
transform 1 0 21200 0 1 5292
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_1
timestamp 1754861848
transform 1 0 21200 0 1 3780
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_2
timestamp 1754861848
transform 1 0 13640 0 1 6048
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_3
timestamp 1754861848
transform 1 0 13640 0 1 4536
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_4
timestamp 1754861848
transform 1 0 13640 0 1 7560
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_5
timestamp 1754861848
transform 1 0 13640 0 1 9072
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_6
timestamp 1754861848
transform 1 0 13640 0 1 10584
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_7
timestamp 1754861848
transform 1 0 13640 0 1 12096
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_8
timestamp 1754861848
transform 1 0 21200 0 1 6804
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_9
timestamp 1754861848
transform 1 0 21200 0 1 8316
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_10
timestamp 1754861848
transform 1 0 21200 0 1 11340
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_11
timestamp 1754861848
transform 1 0 21200 0 1 9828
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_12
timestamp 1754861848
transform 1 0 6080 0 1 3780
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_13
timestamp 1754861848
transform 1 0 6080 0 1 5292
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_14
timestamp 1754861848
transform 1 0 6080 0 1 8316
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_15
timestamp 1754861848
transform 1 0 6080 0 1 6804
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_16
timestamp 1754861848
transform 1 0 6080 0 1 9828
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_17
timestamp 1754861848
transform 1 0 6080 0 1 11340
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_18
timestamp 1754861848
transform 1 0 6080 0 1 14364
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_19
timestamp 1754861848
transform 1 0 6080 0 1 15876
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_20
timestamp 1754861848
transform 1 0 6080 0 1 17388
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_21
timestamp 1754861848
transform 1 0 6080 0 1 18900
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_22
timestamp 1754861848
transform 1 0 6080 0 1 20412
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_23
timestamp 1754861848
transform 1 0 6080 0 1 21924
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_24
timestamp 1754861848
transform 1 0 21200 0 1 15876
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_25
timestamp 1754861848
transform 1 0 21200 0 1 14364
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_26
timestamp 1754861848
transform 1 0 21200 0 1 17388
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_27
timestamp 1754861848
transform 1 0 21200 0 1 18900
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_28
timestamp 1754861848
transform 1 0 13640 0 1 13608
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_29
timestamp 1754861848
transform 1 0 13640 0 1 15120
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_30
timestamp 1754861848
transform 1 0 13640 0 1 16632
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_31
timestamp 1754861848
transform 1 0 13640 0 1 18144
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_32
timestamp 1754861848
transform 1 0 13640 0 1 21168
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_33
timestamp 1754861848
transform 1 0 13640 0 1 19656
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_34
timestamp 1754861848
transform 1 0 21200 0 1 21924
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_35
timestamp 1754861848
transform 1 0 21200 0 1 20412
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_36
timestamp 1754861848
transform 1 0 21200 0 1 12852
box -193 -29 193 29
use VIA_via3_4_2200_440_1_5_410_410  VIA_via3_4_2200_440_1_5_410_410_37
timestamp 1754861848
transform 1 0 6080 0 1 12852
box -193 -29 193 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_0
timestamp 1754861848
transform 1 0 24880 0 1 6048
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_1
timestamp 1754861848
transform 1 0 23480 0 1 5292
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_2
timestamp 1754861848
transform 1 0 24880 0 1 4536
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_3
timestamp 1754861848
transform 1 0 23480 0 1 3780
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_4
timestamp 1754861848
transform 1 0 23480 0 1 8316
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_5
timestamp 1754861848
transform 1 0 24880 0 1 9072
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_6
timestamp 1754861848
transform 1 0 24880 0 1 7560
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_7
timestamp 1754861848
transform 1 0 23480 0 1 6804
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_8
timestamp 1754861848
transform 1 0 23480 0 1 11340
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_9
timestamp 1754861848
transform 1 0 24880 0 1 10584
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_10
timestamp 1754861848
transform 1 0 24880 0 1 12096
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_11
timestamp 1754861848
transform 1 0 23480 0 1 9828
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_12
timestamp 1754861848
transform 1 0 1960 0 1 3780
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_13
timestamp 1754861848
transform 1 0 560 0 1 6048
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_14
timestamp 1754861848
transform 1 0 560 0 1 4536
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_15
timestamp 1754861848
transform 1 0 1960 0 1 5292
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_16
timestamp 1754861848
transform 1 0 560 0 1 7560
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_17
timestamp 1754861848
transform 1 0 1960 0 1 6804
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_18
timestamp 1754861848
transform 1 0 1960 0 1 8316
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_19
timestamp 1754861848
transform 1 0 560 0 1 9072
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_20
timestamp 1754861848
transform 1 0 1960 0 1 9828
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_21
timestamp 1754861848
transform 1 0 560 0 1 10584
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_22
timestamp 1754861848
transform 1 0 1960 0 1 11340
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_23
timestamp 1754861848
transform 1 0 560 0 1 12096
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_24
timestamp 1754861848
transform 1 0 560 0 1 15120
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_25
timestamp 1754861848
transform 1 0 1960 0 1 14364
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_26
timestamp 1754861848
transform 1 0 560 0 1 13608
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_27
timestamp 1754861848
transform 1 0 1960 0 1 15876
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_28
timestamp 1754861848
transform 1 0 560 0 1 18144
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_29
timestamp 1754861848
transform 1 0 1960 0 1 18900
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_30
timestamp 1754861848
transform 1 0 1960 0 1 17388
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_31
timestamp 1754861848
transform 1 0 560 0 1 16632
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_32
timestamp 1754861848
transform 1 0 1960 0 1 20412
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_33
timestamp 1754861848
transform 1 0 560 0 1 21168
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_34
timestamp 1754861848
transform 1 0 560 0 1 19656
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_35
timestamp 1754861848
transform 1 0 1960 0 1 21924
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_36
timestamp 1754861848
transform 1 0 24880 0 1 15120
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_37
timestamp 1754861848
transform 1 0 24880 0 1 13608
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_38
timestamp 1754861848
transform 1 0 23480 0 1 15876
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_39
timestamp 1754861848
transform 1 0 23480 0 1 14364
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_40
timestamp 1754861848
transform 1 0 24880 0 1 18144
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_41
timestamp 1754861848
transform 1 0 23480 0 1 17388
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_42
timestamp 1754861848
transform 1 0 24880 0 1 16632
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_43
timestamp 1754861848
transform 1 0 23480 0 1 18900
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_44
timestamp 1754861848
transform 1 0 23480 0 1 20412
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_45
timestamp 1754861848
transform 1 0 24880 0 1 19656
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_46
timestamp 1754861848
transform 1 0 24880 0 1 21168
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_47
timestamp 1754861848
transform 1 0 23480 0 1 21924
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_48
timestamp 1754861848
transform 1 0 23480 0 1 12852
box -480 -29 480 29
use VIA_via3_4_5000_440_1_12_410_410  VIA_via3_4_5000_440_1_12_410_410_49
timestamp 1754861848
transform 1 0 1960 0 1 12852
box -480 -29 480 29
use VIA_Via3_XY  VIA_Via3_XY_0
timestamp 1754861848
transform 1 0 12936 0 1 10272
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_1
timestamp 1754861848
transform 1 0 12936 0 1 11424
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_2
timestamp 1754861848
transform 1 0 12936 0 1 10080
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_3
timestamp 1754861848
transform 1 0 17808 0 1 10752
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_4
timestamp 1754861848
transform 1 0 5796 0 1 8928
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_5
timestamp 1754861848
transform 1 0 5796 0 1 9984
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_6
timestamp 1754861848
transform 1 0 6972 0 1 11808
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_7
timestamp 1754861848
transform 1 0 10164 0 1 12672
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_8
timestamp 1754861848
transform 1 0 10332 0 1 13536
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_9
timestamp 1754861848
transform 1 0 10584 0 1 12960
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_10
timestamp 1754861848
transform 1 0 10164 0 1 13440
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_11
timestamp 1754861848
transform 1 0 10332 0 1 12960
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_12
timestamp 1754861848
transform 1 0 10668 0 1 18816
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_13
timestamp 1754861848
transform 1 0 10668 0 1 17280
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_14
timestamp 1754861848
transform 1 0 10584 0 1 17760
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_15
timestamp 1754861848
transform 1 0 10668 0 1 16128
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_16
timestamp 1754861848
transform 1 0 10668 0 1 16608
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_17
timestamp 1754861848
transform 1 0 5796 0 1 12960
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_18
timestamp 1754861848
transform 1 0 5796 0 1 16320
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_19
timestamp 1754861848
transform 1 0 5796 0 1 18528
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_20
timestamp 1754861848
transform 1 0 6972 0 1 19584
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_21
timestamp 1754861848
transform 1 0 17808 0 1 13728
box -29 -29 29 29
use VIA_Via3_XY  VIA_Via3_XY_22
timestamp 1754861848
transform 1 0 17808 0 1 13152
box -29 -29 29 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_0
timestamp 1754861848
transform 1 0 21200 0 1 5292
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_1
timestamp 1754861848
transform 1 0 21200 0 1 3780
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_2
timestamp 1754861848
transform 1 0 13640 0 1 6048
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_3
timestamp 1754861848
transform 1 0 13640 0 1 4536
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_4
timestamp 1754861848
transform 1 0 13640 0 1 7560
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_5
timestamp 1754861848
transform 1 0 13640 0 1 9072
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_6
timestamp 1754861848
transform 1 0 13640 0 1 12096
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_7
timestamp 1754861848
transform 1 0 13640 0 1 10584
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_8
timestamp 1754861848
transform 1 0 21200 0 1 6804
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_9
timestamp 1754861848
transform 1 0 21200 0 1 8316
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_10
timestamp 1754861848
transform 1 0 21200 0 1 9828
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_11
timestamp 1754861848
transform 1 0 21200 0 1 11340
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_12
timestamp 1754861848
transform 1 0 6080 0 1 3780
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_13
timestamp 1754861848
transform 1 0 6080 0 1 5292
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_14
timestamp 1754861848
transform 1 0 6080 0 1 6804
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_15
timestamp 1754861848
transform 1 0 6080 0 1 8316
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_16
timestamp 1754861848
transform 1 0 6080 0 1 11340
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_17
timestamp 1754861848
transform 1 0 6080 0 1 9828
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_18
timestamp 1754861848
transform 1 0 6080 0 1 14364
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_19
timestamp 1754861848
transform 1 0 6080 0 1 15876
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_20
timestamp 1754861848
transform 1 0 6080 0 1 17388
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_21
timestamp 1754861848
transform 1 0 6080 0 1 18900
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_22
timestamp 1754861848
transform 1 0 6080 0 1 21924
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_23
timestamp 1754861848
transform 1 0 6080 0 1 20412
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_24
timestamp 1754861848
transform 1 0 21200 0 1 14364
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_25
timestamp 1754861848
transform 1 0 21200 0 1 15876
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_26
timestamp 1754861848
transform 1 0 21200 0 1 18900
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_27
timestamp 1754861848
transform 1 0 21200 0 1 17388
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_28
timestamp 1754861848
transform 1 0 13640 0 1 15120
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_29
timestamp 1754861848
transform 1 0 13640 0 1 13608
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_30
timestamp 1754861848
transform 1 0 13640 0 1 16632
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_31
timestamp 1754861848
transform 1 0 13640 0 1 18144
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_32
timestamp 1754861848
transform 1 0 13640 0 1 19656
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_33
timestamp 1754861848
transform 1 0 13640 0 1 21168
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_34
timestamp 1754861848
transform 1 0 21200 0 1 21924
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_35
timestamp 1754861848
transform 1 0 21200 0 1 20412
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_36
timestamp 1754861848
transform 1 0 21200 0 1 12852
box -193 -29 193 29
use VIA_via4_5_2200_440_1_5_410_410  VIA_via4_5_2200_440_1_5_410_410_37
timestamp 1754861848
transform 1 0 6080 0 1 12852
box -193 -29 193 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_0
timestamp 1754861848
transform 1 0 23480 0 1 3780
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_1
timestamp 1754861848
transform 1 0 23480 0 1 5292
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_2
timestamp 1754861848
transform 1 0 24880 0 1 6048
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_3
timestamp 1754861848
transform 1 0 24880 0 1 4536
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_4
timestamp 1754861848
transform 1 0 24880 0 1 9072
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_5
timestamp 1754861848
transform 1 0 23480 0 1 6804
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_6
timestamp 1754861848
transform 1 0 24880 0 1 7560
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_7
timestamp 1754861848
transform 1 0 23480 0 1 8316
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_8
timestamp 1754861848
transform 1 0 24880 0 1 12096
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_9
timestamp 1754861848
transform 1 0 23480 0 1 11340
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_10
timestamp 1754861848
transform 1 0 24880 0 1 10584
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_11
timestamp 1754861848
transform 1 0 23480 0 1 9828
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_12
timestamp 1754861848
transform 1 0 560 0 1 4536
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_13
timestamp 1754861848
transform 1 0 1960 0 1 5292
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_14
timestamp 1754861848
transform 1 0 1960 0 1 3780
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_15
timestamp 1754861848
transform 1 0 560 0 1 6048
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_16
timestamp 1754861848
transform 1 0 1960 0 1 6804
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_17
timestamp 1754861848
transform 1 0 560 0 1 7560
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_18
timestamp 1754861848
transform 1 0 1960 0 1 8316
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_19
timestamp 1754861848
transform 1 0 560 0 1 9072
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_20
timestamp 1754861848
transform 1 0 1960 0 1 11340
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_21
timestamp 1754861848
transform 1 0 560 0 1 10584
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_22
timestamp 1754861848
transform 1 0 1960 0 1 9828
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_23
timestamp 1754861848
transform 1 0 560 0 1 12096
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_24
timestamp 1754861848
transform 1 0 1960 0 1 14364
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_25
timestamp 1754861848
transform 1 0 560 0 1 13608
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_26
timestamp 1754861848
transform 1 0 560 0 1 15120
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_27
timestamp 1754861848
transform 1 0 1960 0 1 15876
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_28
timestamp 1754861848
transform 1 0 1960 0 1 17388
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_29
timestamp 1754861848
transform 1 0 1960 0 1 18900
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_30
timestamp 1754861848
transform 1 0 560 0 1 18144
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_31
timestamp 1754861848
transform 1 0 560 0 1 16632
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_32
timestamp 1754861848
transform 1 0 1960 0 1 21924
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_33
timestamp 1754861848
transform 1 0 560 0 1 21168
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_34
timestamp 1754861848
transform 1 0 1960 0 1 20412
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_35
timestamp 1754861848
transform 1 0 560 0 1 19656
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_36
timestamp 1754861848
transform 1 0 23480 0 1 15876
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_37
timestamp 1754861848
transform 1 0 23480 0 1 14364
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_38
timestamp 1754861848
transform 1 0 24880 0 1 13608
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_39
timestamp 1754861848
transform 1 0 24880 0 1 15120
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_40
timestamp 1754861848
transform 1 0 24880 0 1 18144
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_41
timestamp 1754861848
transform 1 0 23480 0 1 17388
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_42
timestamp 1754861848
transform 1 0 24880 0 1 16632
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_43
timestamp 1754861848
transform 1 0 23480 0 1 18900
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_44
timestamp 1754861848
transform 1 0 23480 0 1 20412
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_45
timestamp 1754861848
transform 1 0 24880 0 1 19656
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_46
timestamp 1754861848
transform 1 0 24880 0 1 21168
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_47
timestamp 1754861848
transform 1 0 23480 0 1 21924
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_48
timestamp 1754861848
transform 1 0 1960 0 1 12852
box -480 -29 480 29
use VIA_via4_5_5000_440_1_12_410_410  VIA_via4_5_5000_440_1_12_410_410_49
timestamp 1754861848
transform 1 0 23480 0 1 12852
box -480 -29 480 29
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_0
timestamp 1754861848
transform 1 0 21200 0 1 3780
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_1
timestamp 1754861848
transform 1 0 21200 0 1 5292
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_2
timestamp 1754861848
transform 1 0 13640 0 1 6048
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_3
timestamp 1754861848
transform 1 0 13640 0 1 4536
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_4
timestamp 1754861848
transform 1 0 13640 0 1 7560
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_5
timestamp 1754861848
transform 1 0 13640 0 1 9072
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_6
timestamp 1754861848
transform 1 0 13640 0 1 12096
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_7
timestamp 1754861848
transform 1 0 13640 0 1 10584
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_8
timestamp 1754861848
transform 1 0 21200 0 1 8316
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_9
timestamp 1754861848
transform 1 0 21200 0 1 11340
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_10
timestamp 1754861848
transform 1 0 21200 0 1 9828
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_11
timestamp 1754861848
transform 1 0 21200 0 1 6804
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_12
timestamp 1754861848
transform 1 0 6080 0 1 5292
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_13
timestamp 1754861848
transform 1 0 6080 0 1 3780
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_14
timestamp 1754861848
transform 1 0 6080 0 1 8316
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_15
timestamp 1754861848
transform 1 0 6080 0 1 11340
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_16
timestamp 1754861848
transform 1 0 6080 0 1 9828
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_17
timestamp 1754861848
transform 1 0 6080 0 1 6804
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_18
timestamp 1754861848
transform 1 0 6080 0 1 14364
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_19
timestamp 1754861848
transform 1 0 6080 0 1 17388
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_20
timestamp 1754861848
transform 1 0 6080 0 1 18900
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_21
timestamp 1754861848
transform 1 0 6080 0 1 15876
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_22
timestamp 1754861848
transform 1 0 6080 0 1 20412
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_23
timestamp 1754861848
transform 1 0 6080 0 1 21924
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_24
timestamp 1754861848
transform 1 0 21200 0 1 14364
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_25
timestamp 1754861848
transform 1 0 21200 0 1 17388
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_26
timestamp 1754861848
transform 1 0 21200 0 1 18900
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_27
timestamp 1754861848
transform 1 0 21200 0 1 15876
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_28
timestamp 1754861848
transform 1 0 13640 0 1 13608
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_29
timestamp 1754861848
transform 1 0 13640 0 1 15120
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_30
timestamp 1754861848
transform 1 0 13640 0 1 16632
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_31
timestamp 1754861848
transform 1 0 13640 0 1 18144
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_32
timestamp 1754861848
transform 1 0 13640 0 1 21168
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_33
timestamp 1754861848
transform 1 0 13640 0 1 19656
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_34
timestamp 1754861848
transform 1 0 21200 0 1 20412
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_35
timestamp 1754861848
transform 1 0 21200 0 1 21924
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_36
timestamp 1754861848
transform 1 0 21200 0 1 12852
box -220 -126 220 202
use VIA_via5_6_2200_440_1_2_840_840  VIA_via5_6_2200_440_1_2_840_840_37
timestamp 1754861848
transform 1 0 6080 0 1 12852
box -220 -126 220 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_0
timestamp 1754861848
transform 1 0 24880 0 1 6048
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_1
timestamp 1754861848
transform 1 0 23480 0 1 3780
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_2
timestamp 1754861848
transform 1 0 24880 0 1 4536
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_3
timestamp 1754861848
transform 1 0 23480 0 1 5292
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_4
timestamp 1754861848
transform 1 0 24880 0 1 9072
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_5
timestamp 1754861848
transform 1 0 24880 0 1 7560
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_6
timestamp 1754861848
transform 1 0 23480 0 1 8316
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_7
timestamp 1754861848
transform 1 0 24880 0 1 12096
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_8
timestamp 1754861848
transform 1 0 23480 0 1 11340
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_9
timestamp 1754861848
transform 1 0 24880 0 1 10584
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_10
timestamp 1754861848
transform 1 0 23480 0 1 9828
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_11
timestamp 1754861848
transform 1 0 23480 0 1 6804
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_12
timestamp 1754861848
transform 1 0 560 0 1 6048
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_13
timestamp 1754861848
transform 1 0 1960 0 1 3780
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_14
timestamp 1754861848
transform 1 0 560 0 1 4536
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_15
timestamp 1754861848
transform 1 0 1960 0 1 5292
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_16
timestamp 1754861848
transform 1 0 560 0 1 9072
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_17
timestamp 1754861848
transform 1 0 560 0 1 7560
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_18
timestamp 1754861848
transform 1 0 1960 0 1 8316
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_19
timestamp 1754861848
transform 1 0 1960 0 1 11340
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_20
timestamp 1754861848
transform 1 0 560 0 1 12096
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_21
timestamp 1754861848
transform 1 0 560 0 1 10584
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_22
timestamp 1754861848
transform 1 0 1960 0 1 9828
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_23
timestamp 1754861848
transform 1 0 1960 0 1 6804
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_24
timestamp 1754861848
transform 1 0 560 0 1 13608
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_25
timestamp 1754861848
transform 1 0 560 0 1 15120
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_26
timestamp 1754861848
transform 1 0 1960 0 1 14364
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_27
timestamp 1754861848
transform 1 0 1960 0 1 17388
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_28
timestamp 1754861848
transform 1 0 1960 0 1 18900
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_29
timestamp 1754861848
transform 1 0 560 0 1 16632
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_30
timestamp 1754861848
transform 1 0 560 0 1 18144
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_31
timestamp 1754861848
transform 1 0 1960 0 1 15876
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_32
timestamp 1754861848
transform 1 0 1960 0 1 20412
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_33
timestamp 1754861848
transform 1 0 560 0 1 19656
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_34
timestamp 1754861848
transform 1 0 1960 0 1 21924
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_35
timestamp 1754861848
transform 1 0 560 0 1 21168
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_36
timestamp 1754861848
transform 1 0 24880 0 1 13608
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_37
timestamp 1754861848
transform 1 0 23480 0 1 14364
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_38
timestamp 1754861848
transform 1 0 24880 0 1 15120
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_39
timestamp 1754861848
transform 1 0 23480 0 1 18900
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_40
timestamp 1754861848
transform 1 0 24880 0 1 16632
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_41
timestamp 1754861848
transform 1 0 23480 0 1 17388
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_42
timestamp 1754861848
transform 1 0 24880 0 1 18144
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_43
timestamp 1754861848
transform 1 0 23480 0 1 15876
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_44
timestamp 1754861848
transform 1 0 23480 0 1 21924
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_45
timestamp 1754861848
transform 1 0 23480 0 1 20412
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_46
timestamp 1754861848
transform 1 0 24880 0 1 21168
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_47
timestamp 1754861848
transform 1 0 24880 0 1 19656
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_48
timestamp 1754861848
transform 1 0 23480 0 1 12852
box -500 -126 500 202
use VIA_via5_6_5000_440_1_5_840_840  VIA_via5_6_5000_440_1_5_840_840_49
timestamp 1754861848
transform 1 0 1960 0 1 12852
box -500 -126 500 202
use VIA_via6_7_2200_2200_1_1_1960_1960  VIA_via6_7_2200_2200_1_1_1960_1960_0
timestamp 1754861848
transform 1 0 21200 0 1 6494
box -220 -220 220 220
use VIA_via6_7_2200_2200_1_1_1960_1960  VIA_via6_7_2200_2200_1_1_1960_1960_1
timestamp 1754861848
transform 1 0 6080 0 1 6494
box -220 -220 220 220
use VIA_via6_7_2200_2200_1_1_1960_1960  VIA_via6_7_2200_2200_1_1_1960_1960_2
timestamp 1754861848
transform 1 0 6080 0 1 21614
box -220 -220 220 220
use VIA_via6_7_2200_2200_1_1_1960_1960  VIA_via6_7_2200_2200_1_1_1960_1960_3
timestamp 1754861848
transform 1 0 13640 0 1 14054
box -220 -220 220 220
use VIA_via6_7_2200_2200_1_1_1960_1960  VIA_via6_7_2200_2200_1_1_1960_1960_4
timestamp 1754861848
transform 1 0 21200 0 1 21614
box -220 -220 220 220
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_0
timestamp 1754861848
transform 1 0 21200 0 1 2380
box -220 -500 220 500
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_1
timestamp 1754861848
transform 1 0 13640 0 1 980
box -220 -500 220 500
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_2
timestamp 1754861848
transform 1 0 6080 0 1 2380
box -220 -500 220 500
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_3
timestamp 1754861848
transform 1 0 6080 0 1 23324
box -220 -500 220 500
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_4
timestamp 1754861848
transform 1 0 13640 0 1 24724
box -220 -500 220 500
use VIA_via6_7_2200_5000_2_1_1960_1960  VIA_via6_7_2200_5000_2_1_1960_1960_5
timestamp 1754861848
transform 1 0 21200 0 1 23324
box -220 -500 220 500
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_0
timestamp 1754861848
transform 1 0 23480 0 1 6494
box -500 -220 500 220
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_1
timestamp 1754861848
transform 1 0 1960 0 1 6494
box -500 -220 500 220
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_2
timestamp 1754861848
transform 1 0 560 0 1 14054
box -500 -220 500 220
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_3
timestamp 1754861848
transform 1 0 1960 0 1 21614
box -500 -220 500 220
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_4
timestamp 1754861848
transform 1 0 24880 0 1 14054
box -500 -220 500 220
use VIA_via6_7_5000_2200_1_2_1960_1960  VIA_via6_7_5000_2200_1_2_1960_1960_5
timestamp 1754861848
transform 1 0 23480 0 1 21614
box -500 -220 500 220
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_0
timestamp 1754861848
transform 1 0 24880 0 1 980
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_1
timestamp 1754861848
transform 1 0 23480 0 1 2380
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_2
timestamp 1754861848
transform 1 0 1960 0 1 2380
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_3
timestamp 1754861848
transform 1 0 560 0 1 980
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_4
timestamp 1754861848
transform 1 0 560 0 1 24724
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_5
timestamp 1754861848
transform 1 0 1960 0 1 23324
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_6
timestamp 1754861848
transform 1 0 23480 0 1 23324
box -500 -500 500 500
use VIA_via6_7_5000_5000_2_2_1960_1960  VIA_via6_7_5000_5000_2_2_1960_1960_7
timestamp 1754861848
transform 1 0 24880 0 1 24724
box -500 -500 500 500
<< labels >>
rlabel metal2 s 9976 25302 10016 25446 4 cs
port 2 nsew
rlabel metal2 s 15016 25302 15056 25446 4 ctrl0[0]
port 3 nsew
rlabel metal2 s 14596 25302 14636 25446 4 ctrl0[1]
port 4 nsew
rlabel metal2 s 14176 25302 14216 25446 4 ctrl0[2]
port 5 nsew
rlabel metal2 s 13756 25302 13796 25446 4 ctrl0[3]
port 6 nsew
rlabel metal2 s 13336 25302 13376 25446 4 ctrl0[4]
port 7 nsew
rlabel metal2 s 12916 25302 12956 25446 4 ctrl0[5]
port 8 nsew
rlabel metal2 s 12496 25302 12536 25446 4 ctrl0[6]
port 9 nsew
rlabel metal2 s 12076 25302 12116 25446 4 ctrl0[7]
port 10 nsew
rlabel metal2 s 18376 25302 18416 25446 4 ctrl1[0]
port 11 nsew
rlabel metal2 s 17956 25302 17996 25446 4 ctrl1[1]
port 12 nsew
rlabel metal2 s 17536 25302 17576 25446 4 ctrl1[2]
port 13 nsew
rlabel metal2 s 17116 25302 17156 25446 4 ctrl1[3]
port 14 nsew
rlabel metal2 s 16696 25302 16736 25446 4 ctrl1[4]
port 15 nsew
rlabel metal2 s 16276 25302 16316 25446 4 ctrl1[5]
port 16 nsew
rlabel metal2 s 15856 25302 15896 25446 4 ctrl1[6]
port 17 nsew
rlabel metal2 s 15436 25302 15476 25446 4 ctrl1[7]
port 18 nsew
rlabel metal2 s 21736 25302 21776 25446 4 ctrl2[0]
port 19 nsew
rlabel metal2 s 21316 25302 21356 25446 4 ctrl2[1]
port 20 nsew
rlabel metal2 s 20896 25302 20936 25446 4 ctrl2[2]
port 21 nsew
rlabel metal2 s 20476 25302 20516 25446 4 ctrl2[3]
port 22 nsew
rlabel metal2 s 20056 25302 20096 25446 4 ctrl2[4]
port 23 nsew
rlabel metal2 s 19636 25302 19676 25446 4 ctrl2[5]
port 24 nsew
rlabel metal2 s 19216 25302 19256 25446 4 ctrl2[6]
port 25 nsew
rlabel metal2 s 18796 25302 18836 25446 4 ctrl2[7]
port 26 nsew
rlabel metal2 s 10816 25302 10856 25446 4 din
port 27 nsew
rlabel metal2 s 11236 25302 11276 25446 4 dout
port 28 nsew
rlabel metal2 s 11656 25302 11696 25446 4 dout_en
port 29 nsew
rlabel metal2 s 9556 25302 9596 25446 4 reset
port 30 nsew
rlabel metal2 s 10396 25302 10436 25446 4 sclk
port 31 nsew
rlabel metal2 s 25096 25302 25136 25446 4 stat0[0]
port 32 nsew
rlabel metal2 s 24676 25302 24716 25446 4 stat0[1]
port 33 nsew
rlabel metal2 s 24256 25302 24296 25446 4 stat0[2]
port 34 nsew
rlabel metal2 s 23836 25302 23876 25446 4 stat0[3]
port 35 nsew
rlabel metal2 s 23416 25302 23456 25446 4 stat0[4]
port 36 nsew
rlabel metal2 s 22996 25302 23036 25446 4 stat0[5]
port 37 nsew
rlabel metal2 s 22576 25302 22616 25446 4 stat0[6]
port 38 nsew
rlabel metal2 s 22156 25302 22196 25446 4 stat0[7]
port 39 nsew
rlabel metal6 s 60 480 1060 25224 4 VDD
port 41 nsew
rlabel metal6 s 1460 1880 2460 23824 4 VSS
port 42 nsew
rlabel metal7 s 60 480 25380 1480 4 VDD
port 41 nsew
rlabel metal7 s 1460 1880 23980 2880 4 VSS
port 42 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 25446 25446
string GDS_END 529382
string GDS_FILE 6_final.gds
string GDS_START 237050
string path 36.500 59.500 599.500 59.500 
<< end >>
