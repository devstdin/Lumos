magic
tech ihp-sg13g2
timestamp 1754824472
<< metal1 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via1 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal2 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via2 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal3 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via3 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal4 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via4 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal5 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via5 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal6 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< via6 >>
rect 100 6700 6900 6900
rect 100 300 300 6700
rect 6700 300 6900 6700
rect 100 100 6900 300
<< metal7 >>
rect 0 6900 7000 7150
rect 0 100 100 6900
rect 300 6600 6700 6700
rect 300 400 400 6600
rect 6600 400 6700 6600
rect 300 300 6700 400
rect 6900 100 7000 6900
rect 0 0 7000 100
<< pad >>
rect 400 400 6600 6600
<< labels >>
flabel space 0 0 7000 7000 0 FreeSans 800 0 0 0 PAD
port 1 nsew
<< end >>
