magic
tech ihp-sg13g2
timestamp 1748514843
<< error_p >>
rect -93 280 -88 285
rect 88 280 93 285
rect 215 280 220 285
rect 396 280 401 285
rect 523 280 528 285
rect 704 280 709 285
rect 831 280 836 285
rect 1012 280 1017 285
rect 1139 280 1144 285
rect 1320 280 1325 285
rect 1447 280 1452 285
rect 1628 280 1633 285
rect 1755 280 1760 285
rect 1936 280 1941 285
rect 2063 280 2068 285
rect 2244 280 2249 285
rect 2371 280 2376 285
rect 2552 280 2557 285
rect 2679 280 2684 285
rect 2860 280 2865 285
rect 2987 280 2992 285
rect 3168 280 3173 285
rect 3295 280 3300 285
rect 3476 280 3481 285
rect -98 275 -93 280
rect 93 275 98 280
rect 210 275 215 280
rect 401 275 406 280
rect 518 275 523 280
rect 709 275 714 280
rect 826 275 831 280
rect 1017 275 1022 280
rect 1134 275 1139 280
rect 1325 275 1330 280
rect 1442 275 1447 280
rect 1633 275 1638 280
rect 1750 275 1755 280
rect 1941 275 1946 280
rect 2058 275 2063 280
rect 2249 275 2254 280
rect 2366 275 2371 280
rect 2557 275 2562 280
rect 2674 275 2679 280
rect 2865 275 2870 280
rect 2982 275 2987 280
rect 3173 275 3178 280
rect 3290 275 3295 280
rect 3481 275 3486 280
rect -98 264 -93 269
rect 93 264 98 269
rect 210 264 215 269
rect 401 264 406 269
rect 518 264 523 269
rect 709 264 714 269
rect 826 264 831 269
rect 1017 264 1022 269
rect 1134 264 1139 269
rect 1325 264 1330 269
rect 1442 264 1447 269
rect 1633 264 1638 269
rect 1750 264 1755 269
rect 1941 264 1946 269
rect 2058 264 2063 269
rect 2249 264 2254 269
rect 2366 264 2371 269
rect 2557 264 2562 269
rect 2674 264 2679 269
rect 2865 264 2870 269
rect 2982 264 2987 269
rect 3173 264 3178 269
rect 3290 264 3295 269
rect 3481 264 3486 269
rect -93 259 -88 264
rect 88 259 93 264
rect 215 259 220 264
rect 396 259 401 264
rect 523 259 528 264
rect 704 259 709 264
rect 831 259 836 264
rect 1012 259 1017 264
rect 1139 259 1144 264
rect 1320 259 1325 264
rect 1447 259 1452 264
rect 1628 259 1633 264
rect 1755 259 1760 264
rect 1936 259 1941 264
rect 2063 259 2068 264
rect 2244 259 2249 264
rect 2371 259 2376 264
rect 2552 259 2557 264
rect 2679 259 2684 264
rect 2860 259 2865 264
rect 2987 259 2992 264
rect 3168 259 3173 264
rect 3295 259 3300 264
rect 3476 259 3481 264
rect -127 243 -122 248
rect -116 243 -111 248
rect 111 243 116 248
rect 122 243 127 248
rect 181 243 186 248
rect 192 243 197 248
rect 419 243 424 248
rect 430 243 435 248
rect 489 243 494 248
rect 500 243 505 248
rect 727 243 732 248
rect 738 243 743 248
rect 797 243 802 248
rect 808 243 813 248
rect 1035 243 1040 248
rect 1046 243 1051 248
rect 1105 243 1110 248
rect 1116 243 1121 248
rect 1343 243 1348 248
rect 1354 243 1359 248
rect 1413 243 1418 248
rect 1424 243 1429 248
rect 1651 243 1656 248
rect 1662 243 1667 248
rect 1721 243 1726 248
rect 1732 243 1737 248
rect 1959 243 1964 248
rect 1970 243 1975 248
rect 2029 243 2034 248
rect 2040 243 2045 248
rect 2267 243 2272 248
rect 2278 243 2283 248
rect 2337 243 2342 248
rect 2348 243 2353 248
rect 2575 243 2580 248
rect 2586 243 2591 248
rect 2645 243 2650 248
rect 2656 243 2661 248
rect 2883 243 2888 248
rect 2894 243 2899 248
rect 2953 243 2958 248
rect 2964 243 2969 248
rect 3191 243 3196 248
rect 3202 243 3207 248
rect 3261 243 3266 248
rect 3272 243 3277 248
rect 3499 243 3504 248
rect 3510 243 3515 248
rect -132 238 -127 243
rect -111 238 -106 243
rect 106 238 111 243
rect 127 238 132 243
rect 176 238 181 243
rect 197 238 202 243
rect 414 238 419 243
rect 435 238 440 243
rect 484 238 489 243
rect 505 238 510 243
rect 722 238 727 243
rect 743 238 748 243
rect 792 238 797 243
rect 813 238 818 243
rect 1030 238 1035 243
rect 1051 238 1056 243
rect 1100 238 1105 243
rect 1121 238 1126 243
rect 1338 238 1343 243
rect 1359 238 1364 243
rect 1408 238 1413 243
rect 1429 238 1434 243
rect 1646 238 1651 243
rect 1667 238 1672 243
rect 1716 238 1721 243
rect 1737 238 1742 243
rect 1954 238 1959 243
rect 1975 238 1980 243
rect 2024 238 2029 243
rect 2045 238 2050 243
rect 2262 238 2267 243
rect 2283 238 2288 243
rect 2332 238 2337 243
rect 2353 238 2358 243
rect 2570 238 2575 243
rect 2591 238 2596 243
rect 2640 238 2645 243
rect 2661 238 2666 243
rect 2878 238 2883 243
rect 2899 238 2904 243
rect 2948 238 2953 243
rect 2969 238 2974 243
rect 3186 238 3191 243
rect 3207 238 3212 243
rect 3256 238 3261 243
rect 3277 238 3282 243
rect 3494 238 3499 243
rect 3515 238 3520 243
rect -132 -243 -127 -238
rect -111 -243 -106 -238
rect 106 -243 111 -238
rect 127 -243 132 -238
rect 176 -243 181 -238
rect 197 -243 202 -238
rect 414 -243 419 -238
rect 435 -243 440 -238
rect 484 -243 489 -238
rect 505 -243 510 -238
rect 722 -243 727 -238
rect 743 -243 748 -238
rect 792 -243 797 -238
rect 813 -243 818 -238
rect 1030 -243 1035 -238
rect 1051 -243 1056 -238
rect 1100 -243 1105 -238
rect 1121 -243 1126 -238
rect 1338 -243 1343 -238
rect 1359 -243 1364 -238
rect 1408 -243 1413 -238
rect 1429 -243 1434 -238
rect 1646 -243 1651 -238
rect 1667 -243 1672 -238
rect 1716 -243 1721 -238
rect 1737 -243 1742 -238
rect 1954 -243 1959 -238
rect 1975 -243 1980 -238
rect 2024 -243 2029 -238
rect 2045 -243 2050 -238
rect 2262 -243 2267 -238
rect 2283 -243 2288 -238
rect 2332 -243 2337 -238
rect 2353 -243 2358 -238
rect 2570 -243 2575 -238
rect 2591 -243 2596 -238
rect 2640 -243 2645 -238
rect 2661 -243 2666 -238
rect 2878 -243 2883 -238
rect 2899 -243 2904 -238
rect 2948 -243 2953 -238
rect 2969 -243 2974 -238
rect 3186 -243 3191 -238
rect 3207 -243 3212 -238
rect 3256 -243 3261 -238
rect 3277 -243 3282 -238
rect 3494 -243 3499 -238
rect 3515 -243 3520 -238
rect -127 -248 -122 -243
rect -116 -248 -111 -243
rect 111 -248 116 -243
rect 122 -248 127 -243
rect 181 -248 186 -243
rect 192 -248 197 -243
rect 419 -248 424 -243
rect 430 -248 435 -243
rect 489 -248 494 -243
rect 500 -248 505 -243
rect 727 -248 732 -243
rect 738 -248 743 -243
rect 797 -248 802 -243
rect 808 -248 813 -243
rect 1035 -248 1040 -243
rect 1046 -248 1051 -243
rect 1105 -248 1110 -243
rect 1116 -248 1121 -243
rect 1343 -248 1348 -243
rect 1354 -248 1359 -243
rect 1413 -248 1418 -243
rect 1424 -248 1429 -243
rect 1651 -248 1656 -243
rect 1662 -248 1667 -243
rect 1721 -248 1726 -243
rect 1732 -248 1737 -243
rect 1959 -248 1964 -243
rect 1970 -248 1975 -243
rect 2029 -248 2034 -243
rect 2040 -248 2045 -243
rect 2267 -248 2272 -243
rect 2278 -248 2283 -243
rect 2337 -248 2342 -243
rect 2348 -248 2353 -243
rect 2575 -248 2580 -243
rect 2586 -248 2591 -243
rect 2645 -248 2650 -243
rect 2656 -248 2661 -243
rect 2883 -248 2888 -243
rect 2894 -248 2899 -243
rect 2953 -248 2958 -243
rect 2964 -248 2969 -243
rect 3191 -248 3196 -243
rect 3202 -248 3207 -243
rect 3261 -248 3266 -243
rect 3272 -248 3277 -243
rect 3499 -248 3504 -243
rect 3510 -248 3515 -243
rect -93 -264 -88 -259
rect 88 -264 93 -259
rect 215 -264 220 -259
rect 396 -264 401 -259
rect 523 -264 528 -259
rect 704 -264 709 -259
rect 831 -264 836 -259
rect 1012 -264 1017 -259
rect 1139 -264 1144 -259
rect 1320 -264 1325 -259
rect 1447 -264 1452 -259
rect 1628 -264 1633 -259
rect 1755 -264 1760 -259
rect 1936 -264 1941 -259
rect 2063 -264 2068 -259
rect 2244 -264 2249 -259
rect 2371 -264 2376 -259
rect 2552 -264 2557 -259
rect 2679 -264 2684 -259
rect 2860 -264 2865 -259
rect 2987 -264 2992 -259
rect 3168 -264 3173 -259
rect 3295 -264 3300 -259
rect 3476 -264 3481 -259
rect -98 -269 -93 -264
rect 93 -269 98 -264
rect 210 -269 215 -264
rect 401 -269 406 -264
rect 518 -269 523 -264
rect 709 -269 714 -264
rect 826 -269 831 -264
rect 1017 -269 1022 -264
rect 1134 -269 1139 -264
rect 1325 -269 1330 -264
rect 1442 -269 1447 -264
rect 1633 -269 1638 -264
rect 1750 -269 1755 -264
rect 1941 -269 1946 -264
rect 2058 -269 2063 -264
rect 2249 -269 2254 -264
rect 2366 -269 2371 -264
rect 2557 -269 2562 -264
rect 2674 -269 2679 -264
rect 2865 -269 2870 -264
rect 2982 -269 2987 -264
rect 3173 -269 3178 -264
rect 3290 -269 3295 -264
rect 3481 -269 3486 -264
rect -98 -280 -93 -275
rect 93 -280 98 -275
rect 210 -280 215 -275
rect 401 -280 406 -275
rect 518 -280 523 -275
rect 709 -280 714 -275
rect 826 -280 831 -275
rect 1017 -280 1022 -275
rect 1134 -280 1139 -275
rect 1325 -280 1330 -275
rect 1442 -280 1447 -275
rect 1633 -280 1638 -275
rect 1750 -280 1755 -275
rect 1941 -280 1946 -275
rect 2058 -280 2063 -275
rect 2249 -280 2254 -275
rect 2366 -280 2371 -275
rect 2557 -280 2562 -275
rect 2674 -280 2679 -275
rect 2865 -280 2870 -275
rect 2982 -280 2987 -275
rect 3173 -280 3178 -275
rect 3290 -280 3295 -275
rect 3481 -280 3486 -275
rect -93 -285 -88 -280
rect 88 -285 93 -280
rect 215 -285 220 -280
rect 396 -285 401 -280
rect 523 -285 528 -280
rect 704 -285 709 -280
rect 831 -285 836 -280
rect 1012 -285 1017 -280
rect 1139 -285 1144 -280
rect 1320 -285 1325 -280
rect 1447 -285 1452 -280
rect 1628 -285 1633 -280
rect 1755 -285 1760 -280
rect 1936 -285 1941 -280
rect 2063 -285 2068 -280
rect 2244 -285 2249 -280
rect 2371 -285 2376 -280
rect 2552 -285 2557 -280
rect 2679 -285 2684 -280
rect 2860 -285 2865 -280
rect 2987 -285 2992 -280
rect 3168 -285 3173 -280
rect 3295 -285 3300 -280
rect 3476 -285 3481 -280
<< hvnmos >>
rect -100 -250 100 250
rect 208 -250 408 250
rect 516 -250 716 250
rect 824 -250 1024 250
rect 1132 -250 1332 250
rect 1440 -250 1640 250
rect 1748 -250 1948 250
rect 2056 -250 2256 250
rect 2364 -250 2564 250
rect 2672 -250 2872 250
rect 2980 -250 3180 250
rect 3288 -250 3488 250
<< hvndiff >>
rect -134 243 -100 250
rect -134 -243 -127 243
rect -111 -243 -100 243
rect -134 -250 -100 -243
rect 100 243 134 250
rect 100 -243 111 243
rect 127 -243 134 243
rect 100 -250 134 -243
rect 174 243 208 250
rect 174 -243 181 243
rect 197 -243 208 243
rect 174 -250 208 -243
rect 408 243 442 250
rect 408 -243 419 243
rect 435 -243 442 243
rect 408 -250 442 -243
rect 482 243 516 250
rect 482 -243 489 243
rect 505 -243 516 243
rect 482 -250 516 -243
rect 716 243 750 250
rect 716 -243 727 243
rect 743 -243 750 243
rect 716 -250 750 -243
rect 790 243 824 250
rect 790 -243 797 243
rect 813 -243 824 243
rect 790 -250 824 -243
rect 1024 243 1058 250
rect 1024 -243 1035 243
rect 1051 -243 1058 243
rect 1024 -250 1058 -243
rect 1098 243 1132 250
rect 1098 -243 1105 243
rect 1121 -243 1132 243
rect 1098 -250 1132 -243
rect 1332 243 1366 250
rect 1332 -243 1343 243
rect 1359 -243 1366 243
rect 1332 -250 1366 -243
rect 1406 243 1440 250
rect 1406 -243 1413 243
rect 1429 -243 1440 243
rect 1406 -250 1440 -243
rect 1640 243 1674 250
rect 1640 -243 1651 243
rect 1667 -243 1674 243
rect 1640 -250 1674 -243
rect 1714 243 1748 250
rect 1714 -243 1721 243
rect 1737 -243 1748 243
rect 1714 -250 1748 -243
rect 1948 243 1982 250
rect 1948 -243 1959 243
rect 1975 -243 1982 243
rect 1948 -250 1982 -243
rect 2022 243 2056 250
rect 2022 -243 2029 243
rect 2045 -243 2056 243
rect 2022 -250 2056 -243
rect 2256 243 2290 250
rect 2256 -243 2267 243
rect 2283 -243 2290 243
rect 2256 -250 2290 -243
rect 2330 243 2364 250
rect 2330 -243 2337 243
rect 2353 -243 2364 243
rect 2330 -250 2364 -243
rect 2564 243 2598 250
rect 2564 -243 2575 243
rect 2591 -243 2598 243
rect 2564 -250 2598 -243
rect 2638 243 2672 250
rect 2638 -243 2645 243
rect 2661 -243 2672 243
rect 2638 -250 2672 -243
rect 2872 243 2906 250
rect 2872 -243 2883 243
rect 2899 -243 2906 243
rect 2872 -250 2906 -243
rect 2946 243 2980 250
rect 2946 -243 2953 243
rect 2969 -243 2980 243
rect 2946 -250 2980 -243
rect 3180 243 3214 250
rect 3180 -243 3191 243
rect 3207 -243 3214 243
rect 3180 -250 3214 -243
rect 3254 243 3288 250
rect 3254 -243 3261 243
rect 3277 -243 3288 243
rect 3254 -250 3288 -243
rect 3488 243 3522 250
rect 3488 -243 3499 243
rect 3515 -243 3522 243
rect 3488 -250 3522 -243
<< hvndiffc >>
rect -127 -243 -111 243
rect 111 -243 127 243
rect 181 -243 197 243
rect 419 -243 435 243
rect 489 -243 505 243
rect 727 -243 743 243
rect 797 -243 813 243
rect 1035 -243 1051 243
rect 1105 -243 1121 243
rect 1343 -243 1359 243
rect 1413 -243 1429 243
rect 1651 -243 1667 243
rect 1721 -243 1737 243
rect 1959 -243 1975 243
rect 2029 -243 2045 243
rect 2267 -243 2283 243
rect 2337 -243 2353 243
rect 2575 -243 2591 243
rect 2645 -243 2661 243
rect 2883 -243 2899 243
rect 2953 -243 2969 243
rect 3191 -243 3207 243
rect 3261 -243 3277 243
rect 3499 -243 3515 243
<< psubdiff >>
rect -218 332 3606 339
rect -218 316 -181 332
rect 3569 316 3606 332
rect -218 309 3606 316
rect -218 302 -188 309
rect -218 -302 -211 302
rect -195 -302 -188 302
rect 3576 302 3606 309
rect -218 -309 -188 -302
rect 3576 -302 3583 302
rect 3599 -302 3606 302
rect 3576 -309 3606 -302
rect -218 -316 3606 -309
rect -218 -332 -181 -316
rect 3569 -332 3606 -316
rect -218 -339 3606 -332
<< psubdiffcont >>
rect -181 316 3569 332
rect -211 -302 -195 302
rect 3583 -302 3599 302
rect -181 -332 3569 -316
<< poly >>
rect -100 280 100 287
rect -100 264 -93 280
rect 93 264 100 280
rect -100 250 100 264
rect 208 280 408 287
rect 208 264 215 280
rect 401 264 408 280
rect 208 250 408 264
rect 516 280 716 287
rect 516 264 523 280
rect 709 264 716 280
rect 516 250 716 264
rect 824 280 1024 287
rect 824 264 831 280
rect 1017 264 1024 280
rect 824 250 1024 264
rect 1132 280 1332 287
rect 1132 264 1139 280
rect 1325 264 1332 280
rect 1132 250 1332 264
rect 1440 280 1640 287
rect 1440 264 1447 280
rect 1633 264 1640 280
rect 1440 250 1640 264
rect 1748 280 1948 287
rect 1748 264 1755 280
rect 1941 264 1948 280
rect 1748 250 1948 264
rect 2056 280 2256 287
rect 2056 264 2063 280
rect 2249 264 2256 280
rect 2056 250 2256 264
rect 2364 280 2564 287
rect 2364 264 2371 280
rect 2557 264 2564 280
rect 2364 250 2564 264
rect 2672 280 2872 287
rect 2672 264 2679 280
rect 2865 264 2872 280
rect 2672 250 2872 264
rect 2980 280 3180 287
rect 2980 264 2987 280
rect 3173 264 3180 280
rect 2980 250 3180 264
rect 3288 280 3488 287
rect 3288 264 3295 280
rect 3481 264 3488 280
rect 3288 250 3488 264
rect -100 -264 100 -250
rect -100 -280 -93 -264
rect 93 -280 100 -264
rect -100 -287 100 -280
rect 208 -264 408 -250
rect 208 -280 215 -264
rect 401 -280 408 -264
rect 208 -287 408 -280
rect 516 -264 716 -250
rect 516 -280 523 -264
rect 709 -280 716 -264
rect 516 -287 716 -280
rect 824 -264 1024 -250
rect 824 -280 831 -264
rect 1017 -280 1024 -264
rect 824 -287 1024 -280
rect 1132 -264 1332 -250
rect 1132 -280 1139 -264
rect 1325 -280 1332 -264
rect 1132 -287 1332 -280
rect 1440 -264 1640 -250
rect 1440 -280 1447 -264
rect 1633 -280 1640 -264
rect 1440 -287 1640 -280
rect 1748 -264 1948 -250
rect 1748 -280 1755 -264
rect 1941 -280 1948 -264
rect 1748 -287 1948 -280
rect 2056 -264 2256 -250
rect 2056 -280 2063 -264
rect 2249 -280 2256 -264
rect 2056 -287 2256 -280
rect 2364 -264 2564 -250
rect 2364 -280 2371 -264
rect 2557 -280 2564 -264
rect 2364 -287 2564 -280
rect 2672 -264 2872 -250
rect 2672 -280 2679 -264
rect 2865 -280 2872 -264
rect 2672 -287 2872 -280
rect 2980 -264 3180 -250
rect 2980 -280 2987 -264
rect 3173 -280 3180 -264
rect 2980 -287 3180 -280
rect 3288 -264 3488 -250
rect 3288 -280 3295 -264
rect 3481 -280 3488 -264
rect 3288 -287 3488 -280
<< polycont >>
rect -93 264 93 280
rect 215 264 401 280
rect 523 264 709 280
rect 831 264 1017 280
rect 1139 264 1325 280
rect 1447 264 1633 280
rect 1755 264 1941 280
rect 2063 264 2249 280
rect 2371 264 2557 280
rect 2679 264 2865 280
rect 2987 264 3173 280
rect 3295 264 3481 280
rect -93 -280 93 -264
rect 215 -280 401 -264
rect 523 -280 709 -264
rect 831 -280 1017 -264
rect 1139 -280 1325 -264
rect 1447 -280 1633 -264
rect 1755 -280 1941 -264
rect 2063 -280 2249 -264
rect 2371 -280 2557 -264
rect 2679 -280 2865 -264
rect 2987 -280 3173 -264
rect 3295 -280 3481 -264
<< metal1 >>
rect -216 332 3604 337
rect -216 316 -181 332
rect 3569 316 3604 332
rect -216 311 3604 316
rect -216 302 -190 311
rect -216 -302 -211 302
rect -195 -302 -190 302
rect 3578 302 3604 311
rect -216 -311 -190 -302
rect 3578 -302 3583 302
rect 3599 -302 3604 302
rect 3578 -311 3604 -302
rect -216 -316 3604 -311
rect -216 -332 -181 -316
rect 3569 -332 3604 -316
rect -216 -337 3604 -332
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 5 l 2 nf 1 nx 12 dx 0.4 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
