magic
tech ihp-sg13g2
magscale 1 2
timestamp 1748514987
<< metal1 >>
rect 3003 3027 7599 3284
rect 3003 1783 3284 3027
rect 3480 2919 3852 2971
rect 3369 2461 3454 2887
rect 3369 2341 3379 2461
rect 3444 2341 3454 2461
rect 3369 1915 3454 2341
rect 3616 2461 3716 2919
rect 3920 2887 3963 3027
rect 4136 2919 4508 2971
rect 3616 2341 3626 2461
rect 3706 2341 3716 2461
rect 3616 1883 3716 2341
rect 3878 1915 3963 2887
rect 4025 2183 4110 2887
rect 4025 2063 4035 2183
rect 4100 2063 4110 2183
rect 4025 1915 4110 2063
rect 4272 2461 4372 2919
rect 4576 2887 4619 3027
rect 4792 2919 5164 2971
rect 4272 2341 4282 2461
rect 4362 2341 4372 2461
rect 4272 1883 4372 2341
rect 4534 2739 4619 2887
rect 4534 2619 4544 2739
rect 4609 2619 4619 2739
rect 4534 1915 4619 2619
rect 4681 2183 4766 2887
rect 4681 2063 4691 2183
rect 4756 2063 4766 2183
rect 4681 1915 4766 2063
rect 4928 2461 5028 2919
rect 5232 2887 5275 3027
rect 5448 2919 5820 2971
rect 4928 2341 4938 2461
rect 5018 2341 5028 2461
rect 4928 1883 5028 2341
rect 5190 2739 5275 2887
rect 5190 2619 5200 2739
rect 5265 2619 5275 2739
rect 5190 1915 5275 2619
rect 5337 2183 5422 2887
rect 5337 2063 5347 2183
rect 5412 2063 5422 2183
rect 5337 1915 5422 2063
rect 5584 2461 5684 2919
rect 5888 2887 5931 3027
rect 6104 2919 6476 2971
rect 5584 2341 5594 2461
rect 5674 2341 5684 2461
rect 5584 1883 5684 2341
rect 5846 2739 5931 2887
rect 5846 2619 5856 2739
rect 5921 2619 5931 2739
rect 5846 1915 5931 2619
rect 5993 2183 6078 2887
rect 5993 2063 6003 2183
rect 6068 2063 6078 2183
rect 5993 1915 6078 2063
rect 6240 2461 6340 2919
rect 6544 2887 6587 3027
rect 6760 2919 7132 2971
rect 6240 2341 6250 2461
rect 6330 2341 6340 2461
rect 6240 1883 6340 2341
rect 6502 2739 6587 2887
rect 6502 2619 6512 2739
rect 6577 2619 6587 2739
rect 6502 1915 6587 2619
rect 6649 2183 6734 2887
rect 6649 2063 6659 2183
rect 6724 2063 6734 2183
rect 6649 1915 6734 2063
rect 6896 2461 6996 2919
rect 7200 2887 7243 3027
rect 6896 2341 6906 2461
rect 6986 2341 6996 2461
rect 6896 1883 6996 2341
rect 7158 2739 7243 2887
rect 7158 2619 7168 2739
rect 7233 2619 7243 2739
rect 7158 1915 7243 2619
rect 3480 1831 3852 1883
rect 4136 1831 4508 1883
rect 4792 1831 5164 1883
rect 5448 1831 5820 1883
rect 6104 1831 6476 1883
rect 6760 1831 7132 1883
rect -422 1776 3284 1783
rect 7335 1776 7599 3027
rect -422 1428 7599 1776
rect -422 -3096 -54 1428
rect -24 1424 7599 1428
rect 144 1317 316 1369
rect 600 1317 772 1369
rect 1056 1317 1228 1369
rect 1512 1317 1684 1369
rect 1968 1317 2140 1369
rect 2424 1317 2596 1369
rect 2880 1317 3052 1369
rect 3336 1317 3508 1369
rect 3792 1317 3964 1369
rect 4248 1317 4420 1369
rect 4704 1317 4876 1369
rect 5160 1317 5332 1369
rect 5616 1317 5788 1369
rect 6072 1317 6244 1369
rect 6528 1317 6700 1369
rect 6984 1317 7156 1369
rect 31 335 118 1285
rect 31 195 41 335
rect 108 195 118 335
rect 31 -687 118 195
rect 31 -983 76 -687
rect 190 -719 270 1317
rect 342 -687 429 1285
rect 144 -765 316 -719
rect 144 -905 154 -765
rect 306 -905 316 -765
rect 144 -951 316 -905
rect 31 -2955 118 -983
rect 190 -2987 270 -951
rect 384 -983 429 -687
rect 342 -1865 429 -983
rect 342 -2005 352 -1865
rect 419 -2005 429 -1865
rect 342 -2955 429 -2005
rect 487 335 574 1285
rect 487 195 497 335
rect 564 195 574 335
rect 487 -687 574 195
rect 487 -983 532 -687
rect 646 -719 726 1317
rect 798 -687 885 1285
rect 600 -765 772 -719
rect 600 -905 610 -765
rect 762 -905 772 -765
rect 600 -951 772 -905
rect 487 -2955 574 -983
rect 646 -2987 726 -951
rect 840 -983 885 -687
rect 798 -1865 885 -983
rect 798 -2005 808 -1865
rect 875 -2005 885 -1865
rect 798 -2955 885 -2005
rect 943 335 1030 1285
rect 943 195 953 335
rect 1020 195 1030 335
rect 943 -687 1030 195
rect 943 -983 988 -687
rect 1102 -719 1182 1317
rect 1254 -687 1341 1285
rect 1056 -765 1228 -719
rect 1056 -905 1066 -765
rect 1218 -905 1228 -765
rect 1056 -951 1228 -905
rect 943 -2955 1030 -983
rect 1102 -2987 1182 -951
rect 1296 -983 1341 -687
rect 1254 -1865 1341 -983
rect 1254 -2005 1264 -1865
rect 1331 -2005 1341 -1865
rect 1254 -2955 1341 -2005
rect 1399 335 1486 1285
rect 1399 195 1409 335
rect 1476 195 1486 335
rect 1399 -687 1486 195
rect 1399 -983 1444 -687
rect 1558 -719 1638 1317
rect 1710 -687 1797 1285
rect 1512 -765 1684 -719
rect 1512 -905 1522 -765
rect 1674 -905 1684 -765
rect 1512 -951 1684 -905
rect 1399 -2955 1486 -983
rect 1558 -2987 1638 -951
rect 1752 -983 1797 -687
rect 1710 -1865 1797 -983
rect 1710 -2005 1720 -1865
rect 1787 -2005 1797 -1865
rect 1710 -2955 1797 -2005
rect 1855 335 1942 1285
rect 1855 195 1865 335
rect 1932 195 1942 335
rect 1855 -687 1942 195
rect 1855 -983 1900 -687
rect 2014 -719 2094 1317
rect 2166 -687 2253 1285
rect 1968 -765 2140 -719
rect 1968 -905 1978 -765
rect 2130 -905 2140 -765
rect 1968 -951 2140 -905
rect 1855 -2955 1942 -983
rect 2014 -2987 2094 -951
rect 2208 -983 2253 -687
rect 2166 -1865 2253 -983
rect 2166 -2005 2176 -1865
rect 2243 -2005 2253 -1865
rect 2166 -2955 2253 -2005
rect 2311 335 2398 1285
rect 2311 195 2321 335
rect 2388 195 2398 335
rect 2311 -687 2398 195
rect 2311 -983 2356 -687
rect 2470 -719 2550 1317
rect 2622 -687 2709 1285
rect 2424 -765 2596 -719
rect 2424 -905 2434 -765
rect 2586 -905 2596 -765
rect 2424 -951 2596 -905
rect 2311 -2955 2398 -983
rect 2470 -2987 2550 -951
rect 2664 -983 2709 -687
rect 2622 -1865 2709 -983
rect 2622 -2005 2632 -1865
rect 2699 -2005 2709 -1865
rect 2622 -2955 2709 -2005
rect 2767 335 2854 1285
rect 2767 195 2777 335
rect 2844 195 2854 335
rect 2767 -687 2854 195
rect 2767 -983 2812 -687
rect 2926 -719 3006 1317
rect 3078 -687 3165 1285
rect 2880 -765 3052 -719
rect 2880 -905 2890 -765
rect 3042 -905 3052 -765
rect 2880 -951 3052 -905
rect 2767 -2955 2854 -983
rect 2926 -2987 3006 -951
rect 3120 -983 3165 -687
rect 3078 -1865 3165 -983
rect 3078 -2005 3088 -1865
rect 3155 -2005 3165 -1865
rect 3078 -2955 3165 -2005
rect 3223 335 3310 1285
rect 3223 195 3233 335
rect 3300 195 3310 335
rect 3223 -687 3310 195
rect 3223 -983 3268 -687
rect 3382 -719 3462 1317
rect 3534 -687 3621 1285
rect 3336 -765 3508 -719
rect 3336 -905 3346 -765
rect 3498 -905 3508 -765
rect 3336 -951 3508 -905
rect 3223 -2955 3310 -983
rect 3382 -2987 3462 -951
rect 3576 -983 3621 -687
rect 3534 -1865 3621 -983
rect 3534 -2005 3544 -1865
rect 3611 -2005 3621 -1865
rect 3534 -2955 3621 -2005
rect 3679 -687 3766 1285
rect 3679 -983 3724 -687
rect 3838 -719 3918 1317
rect 3990 335 4077 1285
rect 3990 195 4000 335
rect 4067 195 4077 335
rect 3990 -687 4077 195
rect 3792 -765 3964 -719
rect 3792 -905 3802 -765
rect 3954 -905 3964 -765
rect 3792 -951 3964 -905
rect 3679 -1865 3766 -983
rect 3679 -2005 3689 -1865
rect 3756 -2005 3766 -1865
rect 3679 -2955 3766 -2005
rect 3838 -2987 3918 -951
rect 4032 -983 4077 -687
rect 3990 -2955 4077 -983
rect 4135 -687 4222 1285
rect 4135 -983 4180 -687
rect 4294 -719 4374 1317
rect 4446 335 4533 1285
rect 4446 195 4456 335
rect 4523 195 4533 335
rect 4446 -687 4533 195
rect 4248 -765 4420 -719
rect 4248 -905 4258 -765
rect 4410 -905 4420 -765
rect 4248 -951 4420 -905
rect 4135 -1865 4222 -983
rect 4135 -2005 4145 -1865
rect 4212 -2005 4222 -1865
rect 4135 -2955 4222 -2005
rect 4294 -2987 4374 -951
rect 4488 -983 4533 -687
rect 4446 -2955 4533 -983
rect 4591 -687 4678 1285
rect 4591 -983 4636 -687
rect 4750 -719 4830 1317
rect 4902 335 4989 1285
rect 4902 195 4912 335
rect 4979 195 4989 335
rect 4902 -687 4989 195
rect 4704 -765 4876 -719
rect 4704 -905 4714 -765
rect 4866 -905 4876 -765
rect 4704 -951 4876 -905
rect 4591 -1865 4678 -983
rect 4591 -2005 4601 -1865
rect 4668 -2005 4678 -1865
rect 4591 -2955 4678 -2005
rect 4750 -2987 4830 -951
rect 4944 -983 4989 -687
rect 4902 -2955 4989 -983
rect 5047 -687 5134 1285
rect 5047 -983 5092 -687
rect 5206 -719 5286 1317
rect 5358 335 5445 1285
rect 5358 195 5368 335
rect 5435 195 5445 335
rect 5358 -687 5445 195
rect 5160 -765 5332 -719
rect 5160 -905 5170 -765
rect 5322 -905 5332 -765
rect 5160 -951 5332 -905
rect 5047 -1865 5134 -983
rect 5047 -2005 5057 -1865
rect 5124 -2005 5134 -1865
rect 5047 -2955 5134 -2005
rect 5206 -2987 5286 -951
rect 5400 -983 5445 -687
rect 5358 -2955 5445 -983
rect 5503 -687 5590 1285
rect 5503 -983 5548 -687
rect 5662 -719 5742 1317
rect 5814 335 5901 1285
rect 5814 195 5824 335
rect 5891 195 5901 335
rect 5814 -687 5901 195
rect 5616 -765 5788 -719
rect 5616 -905 5626 -765
rect 5778 -905 5788 -765
rect 5616 -951 5788 -905
rect 5503 -1865 5590 -983
rect 5503 -2005 5513 -1865
rect 5580 -2005 5590 -1865
rect 5503 -2955 5590 -2005
rect 5662 -2987 5742 -951
rect 5856 -983 5901 -687
rect 5814 -2955 5901 -983
rect 5959 -687 6046 1285
rect 5959 -983 6004 -687
rect 6118 -719 6198 1317
rect 6270 335 6357 1285
rect 6270 195 6280 335
rect 6347 195 6357 335
rect 6270 -687 6357 195
rect 6072 -765 6244 -719
rect 6072 -905 6082 -765
rect 6234 -905 6244 -765
rect 6072 -951 6244 -905
rect 5959 -1865 6046 -983
rect 5959 -2005 5969 -1865
rect 6036 -2005 6046 -1865
rect 5959 -2955 6046 -2005
rect 6118 -2987 6198 -951
rect 6312 -983 6357 -687
rect 6270 -2955 6357 -983
rect 6415 -687 6502 1285
rect 6415 -983 6460 -687
rect 6574 -719 6654 1317
rect 6726 335 6813 1285
rect 6726 195 6736 335
rect 6803 195 6813 335
rect 6726 -687 6813 195
rect 6528 -765 6700 -719
rect 6528 -905 6538 -765
rect 6690 -905 6700 -765
rect 6528 -951 6700 -905
rect 6415 -1865 6502 -983
rect 6415 -2005 6425 -1865
rect 6492 -2005 6502 -1865
rect 6415 -2955 6502 -2005
rect 6574 -2987 6654 -951
rect 6768 -983 6813 -687
rect 6726 -2955 6813 -983
rect 6871 -687 6958 1285
rect 6871 -983 6916 -687
rect 7030 -719 7110 1317
rect 7182 335 7269 1285
rect 7182 195 7192 335
rect 7259 195 7269 335
rect 7182 -687 7269 195
rect 6984 -765 7156 -719
rect 6984 -905 6994 -765
rect 7146 -905 7156 -765
rect 6984 -951 7156 -905
rect 6871 -1865 6958 -983
rect 6871 -2005 6881 -1865
rect 6948 -2005 6958 -1865
rect 6871 -2955 6958 -2005
rect 7030 -2987 7110 -951
rect 7224 -983 7269 -687
rect 7182 -2955 7269 -983
rect 144 -3039 316 -2987
rect 600 -3039 772 -2987
rect 1056 -3039 1228 -2987
rect 1512 -3039 1684 -2987
rect 1968 -3039 2140 -2987
rect 2424 -3039 2596 -2987
rect 2880 -3039 3052 -2987
rect 3336 -3039 3508 -2987
rect 3792 -3039 3964 -2987
rect 4248 -3039 4420 -2987
rect 4704 -3039 4876 -2987
rect 5160 -3039 5332 -2987
rect 5616 -3039 5788 -2987
rect 6072 -3039 6244 -2987
rect 6528 -3039 6700 -2987
rect 6984 -3039 7156 -2987
rect 7354 -3096 7599 1424
rect -422 -3283 7599 -3096
rect -422 -3610 7599 -3396
rect -422 -4863 -54 -3610
rect 144 -3718 516 -3666
rect 760 -3718 1132 -3666
rect 1376 -3718 1748 -3666
rect 1992 -3718 2364 -3666
rect 2608 -3718 2980 -3666
rect 3224 -3718 3596 -3666
rect 3840 -3718 4212 -3666
rect 4456 -3718 4828 -3666
rect 5072 -3718 5444 -3666
rect 5688 -3718 6060 -3666
rect 6304 -3718 6676 -3666
rect 6920 -3718 7292 -3666
rect 45 -4722 118 -3750
rect 280 -3978 380 -3718
rect 280 -4118 290 -3978
rect 370 -4118 380 -3978
rect 280 -4355 380 -4118
rect 280 -4495 290 -4355
rect 370 -4495 380 -4355
rect 45 -4863 91 -4722
rect 280 -4754 380 -4495
rect 542 -3978 615 -3750
rect 542 -4118 552 -3978
rect 605 -4118 615 -3978
rect 542 -4722 615 -4118
rect 661 -4722 734 -3750
rect 896 -4355 996 -3718
rect 896 -4495 906 -4355
rect 986 -4495 996 -4355
rect 144 -4806 516 -4754
rect 661 -4863 707 -4722
rect 896 -4754 996 -4495
rect 1158 -3978 1231 -3750
rect 1158 -4118 1168 -3978
rect 1221 -4118 1231 -3978
rect 1158 -4722 1231 -4118
rect 1277 -4722 1350 -3750
rect 1512 -4355 1612 -3718
rect 1512 -4495 1522 -4355
rect 1602 -4495 1612 -4355
rect 760 -4806 1132 -4754
rect 1277 -4863 1323 -4722
rect 1512 -4754 1612 -4495
rect 1774 -3978 1847 -3750
rect 1774 -4118 1784 -3978
rect 1837 -4118 1847 -3978
rect 1774 -4722 1847 -4118
rect 1893 -4722 1966 -3750
rect 2128 -4355 2228 -3718
rect 2128 -4495 2138 -4355
rect 2218 -4495 2228 -4355
rect 1376 -4806 1748 -4754
rect 1893 -4863 1939 -4722
rect 2128 -4754 2228 -4495
rect 2390 -3978 2463 -3750
rect 2390 -4118 2400 -3978
rect 2453 -4118 2463 -3978
rect 2390 -4722 2463 -4118
rect 2509 -4722 2582 -3750
rect 2744 -4355 2844 -3718
rect 2744 -4495 2754 -4355
rect 2834 -4495 2844 -4355
rect 1992 -4806 2364 -4754
rect 2509 -4863 2555 -4722
rect 2744 -4754 2844 -4495
rect 3006 -3978 3079 -3750
rect 3006 -4118 3016 -3978
rect 3069 -4118 3079 -3978
rect 3006 -4722 3079 -4118
rect 3125 -4722 3198 -3750
rect 3360 -4355 3460 -3718
rect 3360 -4495 3370 -4355
rect 3450 -4495 3460 -4355
rect 2608 -4806 2980 -4754
rect 3125 -4863 3171 -4722
rect 3360 -4754 3460 -4495
rect 3622 -3978 3695 -3750
rect 3622 -4118 3632 -3978
rect 3685 -4118 3695 -3978
rect 3622 -4722 3695 -4118
rect 3741 -4722 3814 -3750
rect 3976 -4355 4076 -3718
rect 3976 -4495 3986 -4355
rect 4066 -4495 4076 -4355
rect 3224 -4806 3596 -4754
rect 3741 -4863 3787 -4722
rect 3976 -4754 4076 -4495
rect 4238 -3978 4311 -3750
rect 4238 -4118 4248 -3978
rect 4301 -4118 4311 -3978
rect 4238 -4722 4311 -4118
rect 4357 -4722 4430 -3750
rect 4592 -4355 4692 -3718
rect 4592 -4495 4602 -4355
rect 4682 -4495 4692 -4355
rect 3840 -4806 4212 -4754
rect 4357 -4863 4403 -4722
rect 4592 -4754 4692 -4495
rect 4854 -3978 4927 -3750
rect 4854 -4118 4864 -3978
rect 4917 -4118 4927 -3978
rect 4854 -4722 4927 -4118
rect 4973 -4722 5046 -3750
rect 5208 -4355 5308 -3718
rect 5208 -4495 5218 -4355
rect 5298 -4495 5308 -4355
rect 4456 -4806 4828 -4754
rect 4973 -4863 5019 -4722
rect 5208 -4754 5308 -4495
rect 5470 -3978 5543 -3750
rect 5470 -4118 5480 -3978
rect 5533 -4118 5543 -3978
rect 5470 -4722 5543 -4118
rect 5589 -4722 5662 -3750
rect 5824 -4355 5924 -3718
rect 5824 -4495 5834 -4355
rect 5914 -4495 5924 -4355
rect 5072 -4806 5444 -4754
rect 5589 -4863 5635 -4722
rect 5824 -4754 5924 -4495
rect 6086 -3978 6159 -3750
rect 6086 -4118 6096 -3978
rect 6149 -4118 6159 -3978
rect 6086 -4722 6159 -4118
rect 6205 -4722 6278 -3750
rect 6440 -4355 6540 -3718
rect 6440 -4495 6450 -4355
rect 6530 -4495 6540 -4355
rect 5688 -4806 6060 -4754
rect 6205 -4863 6251 -4722
rect 6440 -4754 6540 -4495
rect 6702 -3978 6775 -3750
rect 6702 -4118 6712 -3978
rect 6765 -4118 6775 -3978
rect 6702 -4722 6775 -4118
rect 6821 -4722 6894 -3750
rect 7056 -4355 7156 -3718
rect 7056 -4495 7066 -4355
rect 7146 -4495 7156 -4355
rect 6304 -4806 6676 -4754
rect 6821 -4863 6867 -4722
rect 7056 -4754 7156 -4495
rect 7318 -3978 7391 -3750
rect 7318 -4118 7328 -3978
rect 7381 -4118 7391 -3978
rect 7318 -4722 7391 -4118
rect 6920 -4806 7292 -4754
rect 7490 -4863 7599 -3610
rect -422 -5151 7599 -4863
rect 6203 -5290 6307 -5280
rect 6203 -5362 6213 -5290
rect 6297 -5362 6307 -5290
rect 6203 -5372 6307 -5362
rect 7067 -5290 7171 -5280
rect 7067 -5362 7077 -5290
rect 7161 -5362 7171 -5290
rect 7067 -5372 7171 -5362
<< via1 >>
rect 3379 2341 3444 2461
rect 3626 2341 3706 2461
rect 4035 2063 4100 2183
rect 4282 2341 4362 2461
rect 4544 2619 4609 2739
rect 4691 2063 4756 2183
rect 4938 2341 5018 2461
rect 5200 2619 5265 2739
rect 5347 2063 5412 2183
rect 5594 2341 5674 2461
rect 5856 2619 5921 2739
rect 6003 2063 6068 2183
rect 6250 2341 6330 2461
rect 6512 2619 6577 2739
rect 6659 2063 6724 2183
rect 6906 2341 6986 2461
rect 7168 2619 7233 2739
rect 41 195 108 335
rect 154 -905 306 -765
rect 352 -2005 419 -1865
rect 497 195 564 335
rect 610 -905 762 -765
rect 808 -2005 875 -1865
rect 953 195 1020 335
rect 1066 -905 1218 -765
rect 1264 -2005 1331 -1865
rect 1409 195 1476 335
rect 1522 -905 1674 -765
rect 1720 -2005 1787 -1865
rect 1865 195 1932 335
rect 1978 -905 2130 -765
rect 2176 -2005 2243 -1865
rect 2321 195 2388 335
rect 2434 -905 2586 -765
rect 2632 -2005 2699 -1865
rect 2777 195 2844 335
rect 2890 -905 3042 -765
rect 3088 -2005 3155 -1865
rect 3233 195 3300 335
rect 3346 -905 3498 -765
rect 3544 -2005 3611 -1865
rect 4000 195 4067 335
rect 3802 -905 3954 -765
rect 3689 -2005 3756 -1865
rect 4456 195 4523 335
rect 4258 -905 4410 -765
rect 4145 -2005 4212 -1865
rect 4912 195 4979 335
rect 4714 -905 4866 -765
rect 4601 -2005 4668 -1865
rect 5368 195 5435 335
rect 5170 -905 5322 -765
rect 5057 -2005 5124 -1865
rect 5824 195 5891 335
rect 5626 -905 5778 -765
rect 5513 -2005 5580 -1865
rect 6280 195 6347 335
rect 6082 -905 6234 -765
rect 5969 -2005 6036 -1865
rect 6736 195 6803 335
rect 6538 -905 6690 -765
rect 6425 -2005 6492 -1865
rect 7192 195 7259 335
rect 6994 -905 7146 -765
rect 6881 -2005 6948 -1865
rect 290 -4118 370 -3978
rect 290 -4495 370 -4355
rect 552 -4118 605 -3978
rect 906 -4495 986 -4355
rect 1168 -4118 1221 -3978
rect 1522 -4495 1602 -4355
rect 1784 -4118 1837 -3978
rect 2138 -4495 2218 -4355
rect 2400 -4118 2453 -3978
rect 2754 -4495 2834 -4355
rect 3016 -4118 3069 -3978
rect 3370 -4495 3450 -4355
rect 3632 -4118 3685 -3978
rect 3986 -4495 4066 -4355
rect 4248 -4118 4301 -3978
rect 4602 -4495 4682 -4355
rect 4864 -4118 4917 -3978
rect 5218 -4495 5298 -4355
rect 5480 -4118 5533 -3978
rect 5834 -4495 5914 -4355
rect 6096 -4118 6149 -3978
rect 6450 -4495 6530 -4355
rect 6712 -4118 6765 -3978
rect 7066 -4495 7146 -4355
rect 7328 -4118 7381 -3978
rect 6213 -5362 6297 -5290
rect 7077 -5362 7161 -5290
<< metal2 >>
rect 4025 2739 5275 2749
rect 2541 2471 2897 2663
rect 4025 2619 4544 2739
rect 4609 2619 5200 2739
rect 5265 2619 5275 2739
rect 4025 2609 5275 2619
rect 5337 2739 7243 2749
rect 5337 2619 5856 2739
rect 5921 2619 6512 2739
rect 6577 2619 7168 2739
rect 7233 2619 7243 2739
rect 5337 2609 7243 2619
rect 2541 2461 7243 2471
rect 2541 2341 3379 2461
rect 3444 2341 3626 2461
rect 3706 2341 4282 2461
rect 4362 2341 4938 2461
rect 5018 2341 5594 2461
rect 5674 2341 6250 2461
rect 6330 2341 6906 2461
rect 6986 2341 7243 2461
rect 2541 2331 7243 2341
rect 4025 2183 5275 2193
rect 4025 2063 4035 2183
rect 4100 2063 4691 2183
rect 4756 2063 5275 2183
rect 4025 2053 5275 2063
rect 5337 2183 7674 2193
rect 5337 2063 5347 2183
rect 5412 2063 6003 2183
rect 6068 2063 6659 2183
rect 6724 2063 7674 2183
rect 5337 2053 7674 2063
rect 4590 1657 4710 2053
rect 3576 1534 4710 1657
rect 3576 345 3724 1534
rect 31 335 7269 345
rect 31 195 41 335
rect 108 195 497 335
rect 564 195 953 335
rect 1020 195 1409 335
rect 1476 195 1865 335
rect 1932 195 2321 335
rect 2388 195 2777 335
rect 2844 195 3233 335
rect 3300 195 4000 335
rect 4067 195 4456 335
rect 4523 195 4912 335
rect 4979 195 5368 335
rect 5435 195 5824 335
rect 5891 195 6280 335
rect 6347 195 6736 335
rect 6803 195 7192 335
rect 7259 195 7269 335
rect 31 185 7269 195
rect -422 -627 -191 -527
rect -422 -687 3756 -627
rect 3679 -755 3756 -687
rect -422 -765 3621 -755
rect -422 -905 154 -765
rect 306 -905 610 -765
rect 762 -905 1066 -765
rect 1218 -905 1522 -765
rect 1674 -905 1978 -765
rect 2130 -905 2434 -765
rect 2586 -905 2890 -765
rect 3042 -905 3346 -765
rect 3498 -905 3621 -765
rect -422 -915 3621 -905
rect 3679 -765 7224 -755
rect 3679 -905 3802 -765
rect 3954 -905 4258 -765
rect 4410 -905 4714 -765
rect 4866 -905 5170 -765
rect 5322 -905 5626 -765
rect 5778 -905 6082 -765
rect 6234 -905 6538 -765
rect 6690 -905 6994 -765
rect 7146 -905 7224 -765
rect 3679 -915 7224 -905
rect 3544 -983 3621 -915
rect 3544 -1043 7224 -983
rect 31 -1865 3621 -1855
rect 31 -2005 352 -1865
rect 419 -2005 808 -1865
rect 875 -2005 1264 -1865
rect 1331 -2005 1720 -1865
rect 1787 -2005 2176 -1865
rect 2243 -2005 2632 -1865
rect 2699 -2005 3088 -1865
rect 3155 -2005 3544 -1865
rect 3611 -2005 3621 -1865
rect 31 -2015 3621 -2005
rect 3679 -1865 7269 -1855
rect 3679 -2005 3689 -1865
rect 3756 -2005 4145 -1865
rect 4212 -2005 4601 -1865
rect 4668 -2005 5057 -1865
rect 5124 -2005 5513 -1865
rect 5580 -2005 5969 -1865
rect 6036 -2005 6425 -1865
rect 6492 -2005 6881 -1865
rect 6948 -2005 7269 -1865
rect 3679 -2015 7269 -2005
rect 3120 -3166 3223 -2015
rect 584 -3269 3223 -3166
rect 584 -3968 661 -3269
rect 4032 -3396 4135 -2015
rect 3048 -3499 4135 -3396
rect 3048 -3968 3125 -3499
rect 7478 -3968 7674 2053
rect 76 -3978 2463 -3968
rect 76 -4118 290 -3978
rect 370 -4118 552 -3978
rect 605 -4118 1168 -3978
rect 1221 -4118 1784 -3978
rect 1837 -4118 2400 -3978
rect 2453 -4118 2463 -3978
rect 76 -4128 2463 -4118
rect 2509 -3978 4927 -3968
rect 2509 -4118 3016 -3978
rect 3069 -4118 3632 -3978
rect 3685 -4118 4248 -3978
rect 4301 -4118 4864 -3978
rect 4917 -4118 4927 -3978
rect 2509 -4128 4927 -4118
rect 4973 -3978 7674 -3968
rect 4973 -4118 5480 -3978
rect 5533 -4118 6096 -3978
rect 6149 -4118 6712 -3978
rect 6765 -4118 7328 -3978
rect 7381 -4118 7674 -3978
rect 4973 -4128 7674 -4118
rect 4854 -4205 4927 -4128
rect 4854 -4268 5046 -4205
rect 4973 -4345 5046 -4268
rect 76 -4355 4927 -4345
rect 76 -4495 290 -4355
rect 370 -4495 906 -4355
rect 986 -4495 1522 -4355
rect 1602 -4495 2138 -4355
rect 2218 -4495 2754 -4355
rect 2834 -4495 3370 -4355
rect 3450 -4495 3986 -4355
rect 4066 -4495 4602 -4355
rect 4682 -4495 4927 -4355
rect 76 -4505 4927 -4495
rect 4973 -4355 7360 -4345
rect 4973 -4495 5218 -4355
rect 5298 -4495 5834 -4355
rect 5914 -4495 6450 -4355
rect 6530 -4495 7066 -4355
rect 7146 -4495 7360 -4355
rect 4973 -4505 7360 -4495
rect 5901 -5290 6307 -5280
rect 5901 -5546 5911 -5290
rect 6057 -5362 6213 -5290
rect 6297 -5362 6307 -5290
rect 6057 -5372 6307 -5362
rect 7067 -5290 7171 -4505
rect 7067 -5362 7077 -5290
rect 7161 -5362 7171 -5290
rect 7067 -5372 7171 -5362
rect 6057 -5546 6067 -5372
rect 5901 -5556 6067 -5546
rect 7478 -5789 7674 -4128
rect 6065 -5809 7674 -5789
rect 6065 -6596 6085 -5809
rect 7145 -6596 7674 -5809
rect 6065 -6616 7674 -6596
<< via2 >>
rect 5911 -5546 6057 -5290
rect 6085 -6596 7145 -5809
<< metal3 >>
rect 5901 -5290 6067 -5280
rect 5901 -5546 5911 -5290
rect 6057 -5546 6067 -5290
rect 5901 -5556 6067 -5546
rect 6065 -5809 7165 -5789
rect 6065 -6596 6085 -5809
rect 7145 -6596 7165 -5809
rect 6065 -6616 7165 -6596
<< via3 >>
rect 5911 -5546 6057 -5290
rect 6085 -6596 7145 -5809
<< metal4 >>
rect -422 -5280 5818 -5022
rect -422 -5290 6067 -5280
rect -422 -5546 5911 -5290
rect 6057 -5546 6067 -5290
rect -422 -5556 6067 -5546
rect -422 -9462 5818 -5556
rect 6065 -5809 7165 -5789
rect 6065 -6596 6085 -5809
rect 7145 -6596 7165 -5809
rect 6065 -6616 7165 -6596
<< via4 >>
rect 6085 -6596 7145 -5809
<< metal5 >>
rect 6065 -5809 7165 -5789
rect 6065 -6596 6085 -5809
rect 7145 -6596 7165 -5809
rect 6065 -6616 7165 -6596
<< via5 >>
rect 6185 -6496 7045 -5909
<< metal6 >>
rect -230 -5789 5626 -5214
rect -230 -5909 7165 -5789
rect -230 -6496 6185 -5909
rect 7045 -6496 7165 -5909
rect -230 -6616 7165 -6496
rect -230 -9270 5626 -6616
use cmim_625XFL  cmim_625XFL_0
timestamp 1748298163
transform 1 0 2698 0 1 -7242
box -3120 -2220 3120 2220
use hvnmos_8GWNTL  hvnmos_8GWNTL_0
timestamp 1748514843
transform 1 0 330 0 1 -4236
box -436 -678 7212 678
use hvpmos_QGER4M  hvpmos_QGER4M_0
timestamp 1748514137
transform 1 0 3666 0 1 2401
box -560 -802 3840 802
use hvpmos_Y3H3EP  hvpmos_Y3H3EP_0
timestamp 1748514843
transform 1 0 230 0 1 -1969
box -460 -1302 7300 3570
use rhigh_7UPXCN  rhigh_7UPXCN_0
timestamp 1748298163
transform 0 1 6687 -1 0 -5326
box -230 -616 230 616
<< labels >>
flabel metal2 7478 -6616 7674 -5789 0 FreeSans 800 0 0 0 VOUT
port 0 nsew
flabel metal1 -422 -4926 -125 -3396 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal1 -422 -3283 -125 -1753 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal2 -422 -687 -191 -527 0 FreeSans 800 0 0 0 INP
port 4 nsew
flabel metal2 -422 -915 -191 -755 0 FreeSans 800 0 0 0 INN
port 5 nsew
flabel metal2 2541 2331 2897 2663 0 FreeSans 800 0 0 0 IB
port 1 nsew
<< end >>
