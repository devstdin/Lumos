magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2005 2364 4524
<< nwell >>
rect -124 1152 364 2524
<< pwell >>
rect -5 107 209 1054
rect -114 -5 354 107
<< nmos >>
rect 89 242 115 1028
<< pmos >>
rect 89 1276 115 2158
<< ndiff >>
rect 21 288 89 1028
rect 21 256 35 288
rect 67 256 89 288
rect 21 242 89 256
rect 115 999 183 1028
rect 115 967 137 999
rect 169 967 183 999
rect 115 931 183 967
rect 115 899 137 931
rect 169 899 183 931
rect 115 863 183 899
rect 115 831 137 863
rect 169 831 183 863
rect 115 795 183 831
rect 115 763 137 795
rect 169 763 183 795
rect 115 727 183 763
rect 115 695 137 727
rect 169 695 183 727
rect 115 659 183 695
rect 115 627 137 659
rect 169 627 183 659
rect 115 591 183 627
rect 115 559 137 591
rect 169 559 183 591
rect 115 523 183 559
rect 115 491 137 523
rect 169 491 183 523
rect 115 455 183 491
rect 115 423 137 455
rect 169 423 183 455
rect 115 387 183 423
rect 115 355 137 387
rect 169 355 183 387
rect 115 242 183 355
<< pdiff >>
rect 21 2144 89 2158
rect 21 2112 35 2144
rect 67 2112 89 2144
rect 21 1276 89 2112
rect 115 2031 183 2158
rect 115 1999 137 2031
rect 169 1999 183 2031
rect 115 1963 183 1999
rect 115 1931 137 1963
rect 169 1931 183 1963
rect 115 1895 183 1931
rect 115 1863 137 1895
rect 169 1863 183 1895
rect 115 1827 183 1863
rect 115 1795 137 1827
rect 169 1795 183 1827
rect 115 1759 183 1795
rect 115 1727 137 1759
rect 169 1727 183 1759
rect 115 1691 183 1727
rect 115 1659 137 1691
rect 169 1659 183 1691
rect 115 1623 183 1659
rect 115 1591 137 1623
rect 169 1591 183 1623
rect 115 1555 183 1591
rect 115 1523 137 1555
rect 169 1523 183 1555
rect 115 1487 183 1523
rect 115 1455 137 1487
rect 169 1455 183 1487
rect 115 1419 183 1455
rect 115 1387 137 1419
rect 169 1387 183 1419
rect 115 1351 183 1387
rect 115 1319 137 1351
rect 169 1319 183 1351
rect 115 1276 183 1319
<< ndiffc >>
rect 35 256 67 288
rect 137 967 169 999
rect 137 899 169 931
rect 137 831 169 863
rect 137 763 169 795
rect 137 695 169 727
rect 137 627 169 659
rect 137 559 169 591
rect 137 491 169 523
rect 137 423 169 455
rect 137 355 169 387
<< pdiffc >>
rect 35 2112 67 2144
rect 137 1999 169 2031
rect 137 1931 169 1963
rect 137 1863 169 1895
rect 137 1795 169 1827
rect 137 1727 169 1759
rect 137 1659 169 1691
rect 137 1591 169 1623
rect 137 1523 169 1555
rect 137 1455 169 1487
rect 137 1387 169 1419
rect 137 1319 169 1351
<< psubdiff >>
rect -88 67 328 81
rect -88 35 36 67
rect 68 35 104 67
rect 136 35 172 67
rect 204 35 328 67
rect -88 21 328 35
<< nsubdiff >>
rect 21 2365 219 2379
rect 21 2333 36 2365
rect 68 2333 104 2365
rect 136 2333 172 2365
rect 204 2333 219 2365
rect 21 2319 219 2333
<< psubdiffcont >>
rect 36 35 68 67
rect 104 35 136 67
rect 172 35 204 67
<< nsubdiffcont >>
rect 36 2333 68 2365
rect 104 2333 136 2365
rect 172 2333 204 2365
<< poly >>
rect 89 2158 115 2194
rect 89 1182 115 1276
rect 21 1168 115 1182
rect 21 1136 35 1168
rect 67 1136 115 1168
rect 21 1122 115 1136
rect 89 1028 115 1122
rect 89 206 115 242
<< polycont >>
rect 35 1136 67 1168
<< metal1 >>
rect 0 2365 240 2400
rect 0 2333 36 2365
rect 68 2333 104 2365
rect 136 2333 172 2365
rect 204 2333 240 2365
rect 0 2144 240 2333
rect 0 2112 35 2144
rect 67 2112 240 2144
rect 30 1168 72 2076
rect 30 1136 35 1168
rect 67 1136 72 1168
rect 30 324 72 1136
rect 132 2031 174 2076
rect 132 1999 137 2031
rect 169 1999 174 2031
rect 132 1963 174 1999
rect 132 1931 137 1963
rect 169 1931 174 1963
rect 132 1895 174 1931
rect 132 1863 137 1895
rect 169 1863 174 1895
rect 132 1827 174 1863
rect 132 1795 137 1827
rect 169 1795 174 1827
rect 132 1759 174 1795
rect 132 1727 137 1759
rect 169 1727 174 1759
rect 132 1691 174 1727
rect 132 1659 137 1691
rect 169 1659 174 1691
rect 132 1623 174 1659
rect 132 1591 137 1623
rect 169 1591 174 1623
rect 132 1555 174 1591
rect 132 1523 137 1555
rect 169 1523 174 1555
rect 132 1487 174 1523
rect 132 1455 137 1487
rect 169 1455 174 1487
rect 132 1419 174 1455
rect 132 1387 137 1419
rect 169 1387 174 1419
rect 132 1351 174 1387
rect 132 1319 137 1351
rect 169 1319 174 1351
rect 132 999 174 1319
rect 132 967 137 999
rect 169 967 174 999
rect 132 931 174 967
rect 132 899 137 931
rect 169 899 174 931
rect 132 863 174 899
rect 132 831 137 863
rect 169 831 174 863
rect 132 795 174 831
rect 132 763 137 795
rect 169 763 174 795
rect 132 727 174 763
rect 132 695 137 727
rect 169 695 174 727
rect 132 659 174 695
rect 132 627 137 659
rect 169 627 174 659
rect 132 591 174 627
rect 132 559 137 591
rect 169 559 174 591
rect 132 523 174 559
rect 132 491 137 523
rect 169 491 174 523
rect 132 455 174 491
rect 132 423 137 455
rect 169 423 174 455
rect 132 387 174 423
rect 132 355 137 387
rect 169 355 174 387
rect 132 324 174 355
rect -124 256 35 288
rect 67 256 364 288
rect -124 67 364 256
rect -124 35 36 67
rect 68 35 104 67
rect 136 35 172 67
rect 204 35 364 67
rect -124 0 364 35
<< labels >>
flabel metal1 s 132 324 174 2076 0 FreeSans 800 0 0 0 nq
port 4 nsew
rlabel metal1 s 30 324 72 2076 4 i
port 3 nsew
rlabel metal1 s 0 2112 240 2400 4 vdd
port 1 nsew
rlabel metal1 s 0 0 240 288 4 vss
port 2 nsew
flabel comment s 142 44 142 44 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 22679664
string GDS_FILE sg13g2_io.gds
string GDS_START 22676394
<< end >>
