magic
tech ihp-sg13g2
timestamp 1748517704
<< error_p >>
rect -793 7384 -788 7389
rect 788 7384 793 7389
rect -798 7379 -793 7384
rect 793 7379 798 7384
rect -798 7368 -793 7373
rect 793 7368 798 7373
rect -793 7363 -788 7368
rect 788 7363 793 7368
rect -827 7347 -822 7352
rect -816 7347 -811 7352
rect 811 7347 816 7352
rect 822 7347 827 7352
rect -832 7342 -827 7347
rect -811 7342 -806 7347
rect 806 7342 811 7347
rect 827 7342 832 7347
rect -832 6861 -827 6866
rect -811 6861 -806 6866
rect 806 6861 811 6866
rect 827 6861 832 6866
rect -827 6856 -822 6861
rect -816 6856 -811 6861
rect 811 6856 816 6861
rect 822 6856 827 6861
rect -793 6840 -788 6845
rect 788 6840 793 6845
rect -798 6835 -793 6840
rect 793 6835 798 6840
rect -798 6824 -793 6829
rect 793 6824 798 6829
rect -793 6819 -788 6824
rect 788 6819 793 6824
rect -793 6792 -788 6797
rect 788 6792 793 6797
rect -798 6787 -793 6792
rect 793 6787 798 6792
rect -798 6776 -793 6781
rect 793 6776 798 6781
rect -793 6771 -788 6776
rect 788 6771 793 6776
rect -827 6755 -822 6760
rect -816 6755 -811 6760
rect 811 6755 816 6760
rect 822 6755 827 6760
rect -832 6750 -827 6755
rect -811 6750 -806 6755
rect 806 6750 811 6755
rect 827 6750 832 6755
rect -832 6269 -827 6274
rect -811 6269 -806 6274
rect 806 6269 811 6274
rect 827 6269 832 6274
rect -827 6264 -822 6269
rect -816 6264 -811 6269
rect 811 6264 816 6269
rect 822 6264 827 6269
rect -793 6248 -788 6253
rect 788 6248 793 6253
rect -798 6243 -793 6248
rect 793 6243 798 6248
rect -798 6232 -793 6237
rect 793 6232 798 6237
rect -793 6227 -788 6232
rect 788 6227 793 6232
rect -793 6200 -788 6205
rect 788 6200 793 6205
rect -798 6195 -793 6200
rect 793 6195 798 6200
rect -798 6184 -793 6189
rect 793 6184 798 6189
rect -793 6179 -788 6184
rect 788 6179 793 6184
rect -827 6163 -822 6168
rect -816 6163 -811 6168
rect 811 6163 816 6168
rect 822 6163 827 6168
rect -832 6158 -827 6163
rect -811 6158 -806 6163
rect 806 6158 811 6163
rect 827 6158 832 6163
rect -832 5677 -827 5682
rect -811 5677 -806 5682
rect 806 5677 811 5682
rect 827 5677 832 5682
rect -827 5672 -822 5677
rect -816 5672 -811 5677
rect 811 5672 816 5677
rect 822 5672 827 5677
rect -793 5656 -788 5661
rect 788 5656 793 5661
rect -798 5651 -793 5656
rect 793 5651 798 5656
rect -798 5640 -793 5645
rect 793 5640 798 5645
rect -793 5635 -788 5640
rect 788 5635 793 5640
rect -793 5608 -788 5613
rect 788 5608 793 5613
rect -798 5603 -793 5608
rect 793 5603 798 5608
rect -798 5592 -793 5597
rect 793 5592 798 5597
rect -793 5587 -788 5592
rect 788 5587 793 5592
rect -827 5571 -822 5576
rect -816 5571 -811 5576
rect 811 5571 816 5576
rect 822 5571 827 5576
rect -832 5566 -827 5571
rect -811 5566 -806 5571
rect 806 5566 811 5571
rect 827 5566 832 5571
rect -832 5085 -827 5090
rect -811 5085 -806 5090
rect 806 5085 811 5090
rect 827 5085 832 5090
rect -827 5080 -822 5085
rect -816 5080 -811 5085
rect 811 5080 816 5085
rect 822 5080 827 5085
rect -793 5064 -788 5069
rect 788 5064 793 5069
rect -798 5059 -793 5064
rect 793 5059 798 5064
rect -798 5048 -793 5053
rect 793 5048 798 5053
rect -793 5043 -788 5048
rect 788 5043 793 5048
rect -793 5016 -788 5021
rect 788 5016 793 5021
rect -798 5011 -793 5016
rect 793 5011 798 5016
rect -798 5000 -793 5005
rect 793 5000 798 5005
rect -793 4995 -788 5000
rect 788 4995 793 5000
rect -827 4979 -822 4984
rect -816 4979 -811 4984
rect 811 4979 816 4984
rect 822 4979 827 4984
rect -832 4974 -827 4979
rect -811 4974 -806 4979
rect 806 4974 811 4979
rect 827 4974 832 4979
rect -832 4493 -827 4498
rect -811 4493 -806 4498
rect 806 4493 811 4498
rect 827 4493 832 4498
rect -827 4488 -822 4493
rect -816 4488 -811 4493
rect 811 4488 816 4493
rect 822 4488 827 4493
rect -793 4472 -788 4477
rect 788 4472 793 4477
rect -798 4467 -793 4472
rect 793 4467 798 4472
rect -798 4456 -793 4461
rect 793 4456 798 4461
rect -793 4451 -788 4456
rect 788 4451 793 4456
rect -793 4424 -788 4429
rect 788 4424 793 4429
rect -798 4419 -793 4424
rect 793 4419 798 4424
rect -798 4408 -793 4413
rect 793 4408 798 4413
rect -793 4403 -788 4408
rect 788 4403 793 4408
rect -827 4387 -822 4392
rect -816 4387 -811 4392
rect 811 4387 816 4392
rect 822 4387 827 4392
rect -832 4382 -827 4387
rect -811 4382 -806 4387
rect 806 4382 811 4387
rect 827 4382 832 4387
rect -832 3901 -827 3906
rect -811 3901 -806 3906
rect 806 3901 811 3906
rect 827 3901 832 3906
rect -827 3896 -822 3901
rect -816 3896 -811 3901
rect 811 3896 816 3901
rect 822 3896 827 3901
rect -793 3880 -788 3885
rect 788 3880 793 3885
rect -798 3875 -793 3880
rect 793 3875 798 3880
rect -798 3864 -793 3869
rect 793 3864 798 3869
rect -793 3859 -788 3864
rect 788 3859 793 3864
rect -793 3832 -788 3837
rect 788 3832 793 3837
rect -798 3827 -793 3832
rect 793 3827 798 3832
rect -798 3816 -793 3821
rect 793 3816 798 3821
rect -793 3811 -788 3816
rect 788 3811 793 3816
rect -827 3795 -822 3800
rect -816 3795 -811 3800
rect 811 3795 816 3800
rect 822 3795 827 3800
rect -832 3790 -827 3795
rect -811 3790 -806 3795
rect 806 3790 811 3795
rect 827 3790 832 3795
rect -832 3309 -827 3314
rect -811 3309 -806 3314
rect 806 3309 811 3314
rect 827 3309 832 3314
rect -827 3304 -822 3309
rect -816 3304 -811 3309
rect 811 3304 816 3309
rect 822 3304 827 3309
rect -793 3288 -788 3293
rect 788 3288 793 3293
rect -798 3283 -793 3288
rect 793 3283 798 3288
rect -798 3272 -793 3277
rect 793 3272 798 3277
rect -793 3267 -788 3272
rect 788 3267 793 3272
rect -793 3240 -788 3245
rect 788 3240 793 3245
rect -798 3235 -793 3240
rect 793 3235 798 3240
rect -798 3224 -793 3229
rect 793 3224 798 3229
rect -793 3219 -788 3224
rect 788 3219 793 3224
rect -827 3203 -822 3208
rect -816 3203 -811 3208
rect 811 3203 816 3208
rect 822 3203 827 3208
rect -832 3198 -827 3203
rect -811 3198 -806 3203
rect 806 3198 811 3203
rect 827 3198 832 3203
rect -832 2717 -827 2722
rect -811 2717 -806 2722
rect 806 2717 811 2722
rect 827 2717 832 2722
rect -827 2712 -822 2717
rect -816 2712 -811 2717
rect 811 2712 816 2717
rect 822 2712 827 2717
rect -793 2696 -788 2701
rect 788 2696 793 2701
rect -798 2691 -793 2696
rect 793 2691 798 2696
rect -798 2680 -793 2685
rect 793 2680 798 2685
rect -793 2675 -788 2680
rect 788 2675 793 2680
rect -793 2648 -788 2653
rect 788 2648 793 2653
rect -798 2643 -793 2648
rect 793 2643 798 2648
rect -798 2632 -793 2637
rect 793 2632 798 2637
rect -793 2627 -788 2632
rect 788 2627 793 2632
rect -827 2611 -822 2616
rect -816 2611 -811 2616
rect 811 2611 816 2616
rect 822 2611 827 2616
rect -832 2606 -827 2611
rect -811 2606 -806 2611
rect 806 2606 811 2611
rect 827 2606 832 2611
rect -832 2125 -827 2130
rect -811 2125 -806 2130
rect 806 2125 811 2130
rect 827 2125 832 2130
rect -827 2120 -822 2125
rect -816 2120 -811 2125
rect 811 2120 816 2125
rect 822 2120 827 2125
rect -793 2104 -788 2109
rect 788 2104 793 2109
rect -798 2099 -793 2104
rect 793 2099 798 2104
rect -798 2088 -793 2093
rect 793 2088 798 2093
rect -793 2083 -788 2088
rect 788 2083 793 2088
rect -793 2056 -788 2061
rect 788 2056 793 2061
rect -798 2051 -793 2056
rect 793 2051 798 2056
rect -798 2040 -793 2045
rect 793 2040 798 2045
rect -793 2035 -788 2040
rect 788 2035 793 2040
rect -827 2019 -822 2024
rect -816 2019 -811 2024
rect 811 2019 816 2024
rect 822 2019 827 2024
rect -832 2014 -827 2019
rect -811 2014 -806 2019
rect 806 2014 811 2019
rect 827 2014 832 2019
rect -832 1533 -827 1538
rect -811 1533 -806 1538
rect 806 1533 811 1538
rect 827 1533 832 1538
rect -827 1528 -822 1533
rect -816 1528 -811 1533
rect 811 1528 816 1533
rect 822 1528 827 1533
rect -793 1512 -788 1517
rect 788 1512 793 1517
rect -798 1507 -793 1512
rect 793 1507 798 1512
rect -798 1496 -793 1501
rect 793 1496 798 1501
rect -793 1491 -788 1496
rect 788 1491 793 1496
rect -793 1464 -788 1469
rect 788 1464 793 1469
rect -798 1459 -793 1464
rect 793 1459 798 1464
rect -798 1448 -793 1453
rect 793 1448 798 1453
rect -793 1443 -788 1448
rect 788 1443 793 1448
rect -827 1427 -822 1432
rect -816 1427 -811 1432
rect 811 1427 816 1432
rect 822 1427 827 1432
rect -832 1422 -827 1427
rect -811 1422 -806 1427
rect 806 1422 811 1427
rect 827 1422 832 1427
rect -832 941 -827 946
rect -811 941 -806 946
rect 806 941 811 946
rect 827 941 832 946
rect -827 936 -822 941
rect -816 936 -811 941
rect 811 936 816 941
rect 822 936 827 941
rect -793 920 -788 925
rect 788 920 793 925
rect -798 915 -793 920
rect 793 915 798 920
rect -798 904 -793 909
rect 793 904 798 909
rect -793 899 -788 904
rect 788 899 793 904
rect -793 872 -788 877
rect 788 872 793 877
rect -798 867 -793 872
rect 793 867 798 872
rect -798 856 -793 861
rect 793 856 798 861
rect -793 851 -788 856
rect 788 851 793 856
rect -827 835 -822 840
rect -816 835 -811 840
rect 811 835 816 840
rect 822 835 827 840
rect -832 830 -827 835
rect -811 830 -806 835
rect 806 830 811 835
rect 827 830 832 835
rect -832 349 -827 354
rect -811 349 -806 354
rect 806 349 811 354
rect 827 349 832 354
rect -827 344 -822 349
rect -816 344 -811 349
rect 811 344 816 349
rect 822 344 827 349
rect -793 328 -788 333
rect 788 328 793 333
rect -798 323 -793 328
rect 793 323 798 328
rect -798 312 -793 317
rect 793 312 798 317
rect -793 307 -788 312
rect 788 307 793 312
rect -793 280 -788 285
rect 788 280 793 285
rect -798 275 -793 280
rect 793 275 798 280
rect -798 264 -793 269
rect 793 264 798 269
rect -793 259 -788 264
rect 788 259 793 264
rect -827 243 -822 248
rect -816 243 -811 248
rect 811 243 816 248
rect 822 243 827 248
rect -832 238 -827 243
rect -811 238 -806 243
rect 806 238 811 243
rect 827 238 832 243
rect -832 -243 -827 -238
rect -811 -243 -806 -238
rect 806 -243 811 -238
rect 827 -243 832 -238
rect -827 -248 -822 -243
rect -816 -248 -811 -243
rect 811 -248 816 -243
rect 822 -248 827 -243
rect -793 -264 -788 -259
rect 788 -264 793 -259
rect -798 -269 -793 -264
rect 793 -269 798 -264
rect -798 -280 -793 -275
rect 793 -280 798 -275
rect -793 -285 -788 -280
rect 788 -285 793 -280
<< hvnmos >>
rect -800 6854 800 7354
rect -800 6262 800 6762
rect -800 5670 800 6170
rect -800 5078 800 5578
rect -800 4486 800 4986
rect -800 3894 800 4394
rect -800 3302 800 3802
rect -800 2710 800 3210
rect -800 2118 800 2618
rect -800 1526 800 2026
rect -800 934 800 1434
rect -800 342 800 842
rect -800 -250 800 250
<< hvndiff >>
rect -834 7347 -800 7354
rect -834 6861 -827 7347
rect -811 6861 -800 7347
rect -834 6854 -800 6861
rect 800 7347 834 7354
rect 800 6861 811 7347
rect 827 6861 834 7347
rect 800 6854 834 6861
rect -834 6755 -800 6762
rect -834 6269 -827 6755
rect -811 6269 -800 6755
rect -834 6262 -800 6269
rect 800 6755 834 6762
rect 800 6269 811 6755
rect 827 6269 834 6755
rect 800 6262 834 6269
rect -834 6163 -800 6170
rect -834 5677 -827 6163
rect -811 5677 -800 6163
rect -834 5670 -800 5677
rect 800 6163 834 6170
rect 800 5677 811 6163
rect 827 5677 834 6163
rect 800 5670 834 5677
rect -834 5571 -800 5578
rect -834 5085 -827 5571
rect -811 5085 -800 5571
rect -834 5078 -800 5085
rect 800 5571 834 5578
rect 800 5085 811 5571
rect 827 5085 834 5571
rect 800 5078 834 5085
rect -834 4979 -800 4986
rect -834 4493 -827 4979
rect -811 4493 -800 4979
rect -834 4486 -800 4493
rect 800 4979 834 4986
rect 800 4493 811 4979
rect 827 4493 834 4979
rect 800 4486 834 4493
rect -834 4387 -800 4394
rect -834 3901 -827 4387
rect -811 3901 -800 4387
rect -834 3894 -800 3901
rect 800 4387 834 4394
rect 800 3901 811 4387
rect 827 3901 834 4387
rect 800 3894 834 3901
rect -834 3795 -800 3802
rect -834 3309 -827 3795
rect -811 3309 -800 3795
rect -834 3302 -800 3309
rect 800 3795 834 3802
rect 800 3309 811 3795
rect 827 3309 834 3795
rect 800 3302 834 3309
rect -834 3203 -800 3210
rect -834 2717 -827 3203
rect -811 2717 -800 3203
rect -834 2710 -800 2717
rect 800 3203 834 3210
rect 800 2717 811 3203
rect 827 2717 834 3203
rect 800 2710 834 2717
rect -834 2611 -800 2618
rect -834 2125 -827 2611
rect -811 2125 -800 2611
rect -834 2118 -800 2125
rect 800 2611 834 2618
rect 800 2125 811 2611
rect 827 2125 834 2611
rect 800 2118 834 2125
rect -834 2019 -800 2026
rect -834 1533 -827 2019
rect -811 1533 -800 2019
rect -834 1526 -800 1533
rect 800 2019 834 2026
rect 800 1533 811 2019
rect 827 1533 834 2019
rect 800 1526 834 1533
rect -834 1427 -800 1434
rect -834 941 -827 1427
rect -811 941 -800 1427
rect -834 934 -800 941
rect 800 1427 834 1434
rect 800 941 811 1427
rect 827 941 834 1427
rect 800 934 834 941
rect -834 835 -800 842
rect -834 349 -827 835
rect -811 349 -800 835
rect -834 342 -800 349
rect 800 835 834 842
rect 800 349 811 835
rect 827 349 834 835
rect 800 342 834 349
rect -834 243 -800 250
rect -834 -243 -827 243
rect -811 -243 -800 243
rect -834 -250 -800 -243
rect 800 243 834 250
rect 800 -243 811 243
rect 827 -243 834 243
rect 800 -250 834 -243
<< hvndiffc >>
rect -827 6861 -811 7347
rect 811 6861 827 7347
rect -827 6269 -811 6755
rect 811 6269 827 6755
rect -827 5677 -811 6163
rect 811 5677 827 6163
rect -827 5085 -811 5571
rect 811 5085 827 5571
rect -827 4493 -811 4979
rect 811 4493 827 4979
rect -827 3901 -811 4387
rect 811 3901 827 4387
rect -827 3309 -811 3795
rect 811 3309 827 3795
rect -827 2717 -811 3203
rect 811 2717 827 3203
rect -827 2125 -811 2611
rect 811 2125 827 2611
rect -827 1533 -811 2019
rect 811 1533 827 2019
rect -827 941 -811 1427
rect 811 941 827 1427
rect -827 349 -811 835
rect 811 349 827 835
rect -827 -243 -811 243
rect 811 -243 827 243
<< psubdiff >>
rect -918 7436 918 7443
rect -918 7420 -881 7436
rect 881 7420 918 7436
rect -918 7413 918 7420
rect -918 7406 -888 7413
rect -918 -302 -911 7406
rect -895 -302 -888 7406
rect 888 7406 918 7413
rect -918 -309 -888 -302
rect 888 -302 895 7406
rect 911 -302 918 7406
rect 888 -309 918 -302
rect -918 -316 918 -309
rect -918 -332 -881 -316
rect 881 -332 918 -316
rect -918 -339 918 -332
<< psubdiffcont >>
rect -881 7420 881 7436
rect -911 -302 -895 7406
rect 895 -302 911 7406
rect -881 -332 881 -316
<< poly >>
rect -800 7384 800 7391
rect -800 7368 -793 7384
rect 793 7368 800 7384
rect -800 7354 800 7368
rect -800 6840 800 6854
rect -800 6824 -793 6840
rect 793 6824 800 6840
rect -800 6817 800 6824
rect -800 6792 800 6799
rect -800 6776 -793 6792
rect 793 6776 800 6792
rect -800 6762 800 6776
rect -800 6248 800 6262
rect -800 6232 -793 6248
rect 793 6232 800 6248
rect -800 6225 800 6232
rect -800 6200 800 6207
rect -800 6184 -793 6200
rect 793 6184 800 6200
rect -800 6170 800 6184
rect -800 5656 800 5670
rect -800 5640 -793 5656
rect 793 5640 800 5656
rect -800 5633 800 5640
rect -800 5608 800 5615
rect -800 5592 -793 5608
rect 793 5592 800 5608
rect -800 5578 800 5592
rect -800 5064 800 5078
rect -800 5048 -793 5064
rect 793 5048 800 5064
rect -800 5041 800 5048
rect -800 5016 800 5023
rect -800 5000 -793 5016
rect 793 5000 800 5016
rect -800 4986 800 5000
rect -800 4472 800 4486
rect -800 4456 -793 4472
rect 793 4456 800 4472
rect -800 4449 800 4456
rect -800 4424 800 4431
rect -800 4408 -793 4424
rect 793 4408 800 4424
rect -800 4394 800 4408
rect -800 3880 800 3894
rect -800 3864 -793 3880
rect 793 3864 800 3880
rect -800 3857 800 3864
rect -800 3832 800 3839
rect -800 3816 -793 3832
rect 793 3816 800 3832
rect -800 3802 800 3816
rect -800 3288 800 3302
rect -800 3272 -793 3288
rect 793 3272 800 3288
rect -800 3265 800 3272
rect -800 3240 800 3247
rect -800 3224 -793 3240
rect 793 3224 800 3240
rect -800 3210 800 3224
rect -800 2696 800 2710
rect -800 2680 -793 2696
rect 793 2680 800 2696
rect -800 2673 800 2680
rect -800 2648 800 2655
rect -800 2632 -793 2648
rect 793 2632 800 2648
rect -800 2618 800 2632
rect -800 2104 800 2118
rect -800 2088 -793 2104
rect 793 2088 800 2104
rect -800 2081 800 2088
rect -800 2056 800 2063
rect -800 2040 -793 2056
rect 793 2040 800 2056
rect -800 2026 800 2040
rect -800 1512 800 1526
rect -800 1496 -793 1512
rect 793 1496 800 1512
rect -800 1489 800 1496
rect -800 1464 800 1471
rect -800 1448 -793 1464
rect 793 1448 800 1464
rect -800 1434 800 1448
rect -800 920 800 934
rect -800 904 -793 920
rect 793 904 800 920
rect -800 897 800 904
rect -800 872 800 879
rect -800 856 -793 872
rect 793 856 800 872
rect -800 842 800 856
rect -800 328 800 342
rect -800 312 -793 328
rect 793 312 800 328
rect -800 305 800 312
rect -800 280 800 287
rect -800 264 -793 280
rect 793 264 800 280
rect -800 250 800 264
rect -800 -264 800 -250
rect -800 -280 -793 -264
rect 793 -280 800 -264
rect -800 -287 800 -280
<< polycont >>
rect -793 7368 793 7384
rect -793 6824 793 6840
rect -793 6776 793 6792
rect -793 6232 793 6248
rect -793 6184 793 6200
rect -793 5640 793 5656
rect -793 5592 793 5608
rect -793 5048 793 5064
rect -793 5000 793 5016
rect -793 4456 793 4472
rect -793 4408 793 4424
rect -793 3864 793 3880
rect -793 3816 793 3832
rect -793 3272 793 3288
rect -793 3224 793 3240
rect -793 2680 793 2696
rect -793 2632 793 2648
rect -793 2088 793 2104
rect -793 2040 793 2056
rect -793 1496 793 1512
rect -793 1448 793 1464
rect -793 904 793 920
rect -793 856 793 872
rect -793 312 793 328
rect -793 264 793 280
rect -793 -280 793 -264
<< metal1 >>
rect -916 7436 916 7441
rect -916 7420 -881 7436
rect 881 7420 916 7436
rect -916 7415 916 7420
rect -916 7406 -890 7415
rect -916 -302 -911 7406
rect -895 -302 -890 7406
rect 890 7406 916 7415
rect -916 -311 -890 -302
rect 890 -302 895 7406
rect 911 -302 916 7406
rect 890 -311 916 -302
rect -916 -316 916 -311
rect -916 -332 -881 -316
rect 881 -332 916 -316
rect -916 -337 916 -332
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 5 l 16 nf 1 nx 1 dx 0.22 ny 13 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
