magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752937939
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 225 232 563 270
rect 14 56 563 232
rect -26 -56 602 56
<< nmos >>
rect 108 96 134 206
rect 210 96 236 206
rect 319 96 345 244
rect 435 96 461 244
<< pmos >>
rect 108 492 134 660
rect 210 492 236 660
rect 319 436 345 660
rect 435 436 461 660
<< ndiff >>
rect 251 206 319 244
rect 40 142 108 206
rect 40 110 54 142
rect 86 110 108 142
rect 40 96 108 110
rect 134 142 210 206
rect 134 110 156 142
rect 188 110 210 142
rect 134 96 210 110
rect 236 142 319 206
rect 236 110 265 142
rect 297 110 319 142
rect 236 96 319 110
rect 345 210 435 244
rect 345 178 367 210
rect 399 178 435 210
rect 345 142 435 178
rect 345 110 367 142
rect 399 110 435 142
rect 345 96 435 110
rect 461 210 537 244
rect 461 178 491 210
rect 523 178 537 210
rect 461 142 537 178
rect 461 110 491 142
rect 523 110 537 142
rect 461 96 537 110
<< pdiff >>
rect 40 646 108 660
rect 40 614 54 646
rect 86 614 108 646
rect 40 578 108 614
rect 40 546 54 578
rect 86 546 108 578
rect 40 492 108 546
rect 134 492 210 660
rect 236 646 319 660
rect 236 614 264 646
rect 296 614 319 646
rect 236 578 319 614
rect 236 546 264 578
rect 296 546 319 578
rect 236 510 319 546
rect 236 492 264 510
rect 250 478 264 492
rect 296 478 319 510
rect 250 436 319 478
rect 345 646 435 660
rect 345 614 368 646
rect 400 614 435 646
rect 345 578 435 614
rect 345 546 368 578
rect 400 546 435 578
rect 345 510 435 546
rect 345 478 368 510
rect 400 478 435 510
rect 345 436 435 478
rect 461 646 537 660
rect 461 614 491 646
rect 523 614 537 646
rect 461 578 537 614
rect 461 546 491 578
rect 523 546 537 578
rect 461 510 537 546
rect 461 478 491 510
rect 523 478 537 510
rect 461 436 537 478
<< ndiffc >>
rect 54 110 86 142
rect 156 110 188 142
rect 265 110 297 142
rect 367 178 399 210
rect 367 110 399 142
rect 491 178 523 210
rect 491 110 523 142
<< pdiffc >>
rect 54 614 86 646
rect 54 546 86 578
rect 264 614 296 646
rect 264 546 296 578
rect 264 478 296 510
rect 368 614 400 646
rect 368 546 400 578
rect 368 478 400 510
rect 491 614 523 646
rect 491 546 523 578
rect 491 478 523 510
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 108 660 134 704
rect 210 660 236 705
rect 319 660 345 706
rect 435 660 461 706
rect 108 478 134 492
rect 108 464 174 478
rect 108 432 127 464
rect 159 432 174 464
rect 108 418 174 432
rect 108 206 134 418
rect 210 383 236 492
rect 187 369 247 383
rect 187 337 201 369
rect 233 337 247 369
rect 187 323 247 337
rect 210 206 236 323
rect 319 320 345 436
rect 435 320 461 436
rect 289 306 461 320
rect 289 274 303 306
rect 335 274 461 306
rect 289 260 461 274
rect 319 258 461 260
rect 319 244 345 258
rect 435 244 461 258
rect 108 44 134 96
rect 210 44 236 96
rect 319 44 345 96
rect 435 44 461 96
<< polycont >>
rect 127 432 159 464
rect 201 337 233 369
rect 303 274 335 306
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 44 646 96 656
rect 44 614 54 646
rect 86 614 96 646
rect 44 578 96 614
rect 44 546 54 578
rect 86 546 96 578
rect 254 646 306 712
rect 254 614 264 646
rect 296 614 306 646
rect 254 578 306 614
rect 44 506 96 546
rect 44 225 81 506
rect 168 470 217 576
rect 117 464 217 470
rect 254 546 264 578
rect 296 546 306 578
rect 254 510 306 546
rect 254 478 264 510
rect 296 478 306 510
rect 254 468 306 478
rect 358 646 410 656
rect 358 614 368 646
rect 400 614 410 646
rect 358 578 410 614
rect 358 546 368 578
rect 400 546 410 578
rect 358 510 410 546
rect 358 478 368 510
rect 400 478 410 510
rect 358 468 410 478
rect 481 646 533 712
rect 481 614 491 646
rect 523 614 533 646
rect 481 578 533 614
rect 481 546 491 578
rect 523 546 533 578
rect 481 510 533 546
rect 481 478 491 510
rect 523 478 533 510
rect 481 468 533 478
rect 117 432 127 464
rect 159 432 217 464
rect 117 426 217 432
rect 168 369 243 379
rect 168 337 201 369
rect 233 337 243 369
rect 168 327 243 337
rect 168 267 217 327
rect 285 306 341 316
rect 285 274 303 306
rect 335 274 341 306
rect 285 263 341 274
rect 285 225 319 263
rect 44 189 319 225
rect 377 220 410 468
rect 357 210 410 220
rect 44 142 96 152
rect 44 110 54 142
rect 86 110 96 142
rect 44 44 96 110
rect 146 142 198 189
rect 357 178 367 210
rect 399 178 410 210
rect 146 110 156 142
rect 188 110 198 142
rect 146 100 198 110
rect 255 142 307 152
rect 255 110 265 142
rect 297 110 307 142
rect 255 44 307 110
rect 357 142 410 178
rect 357 110 367 142
rect 399 110 410 142
rect 357 100 410 110
rect 481 210 533 220
rect 481 178 491 210
rect 523 178 533 210
rect 481 142 533 178
rect 481 110 491 142
rect 523 110 533 142
rect 481 44 533 110
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 168 426 217 576 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 168 267 217 379 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 358 468 410 656 0 FreeSans 400 0 0 0 X
port 5 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 464398
string GDS_FILE sg13g2_stdcell.gds
string GDS_START 459992
<< end >>
