magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752864670
<< error_p >>
rect -36 160 -26 170
rect 26 160 36 170
rect 242 160 252 170
rect 304 160 314 170
rect 520 160 530 170
rect 582 160 592 170
rect 798 160 808 170
rect 860 160 870 170
rect -46 150 46 160
rect 232 150 324 160
rect 510 150 602 160
rect 788 150 880 160
rect -36 138 36 150
rect 242 138 314 150
rect 520 138 592 150
rect 798 138 870 150
rect -46 128 46 138
rect 232 128 324 138
rect 510 128 602 138
rect 788 128 880 138
rect -36 118 -26 128
rect 26 118 36 128
rect 242 118 252 128
rect 304 118 314 128
rect 520 118 530 128
rect 582 118 592 128
rect 798 118 808 128
rect 860 118 870 128
rect -104 86 -94 96
rect -82 86 -72 96
rect 72 86 82 96
rect 94 86 104 96
rect 174 86 184 96
rect 196 86 206 96
rect 350 86 360 96
rect 372 86 382 96
rect 452 86 462 96
rect 474 86 484 96
rect 628 86 638 96
rect 650 86 660 96
rect 730 86 740 96
rect 752 86 762 96
rect 906 86 916 96
rect 928 86 938 96
rect -114 76 -104 86
rect -72 76 -62 86
rect 62 76 72 86
rect 104 76 114 86
rect 164 76 174 86
rect 206 76 216 86
rect 340 76 350 86
rect 382 76 392 86
rect 442 76 452 86
rect 484 76 494 86
rect 618 76 628 86
rect 660 76 670 86
rect 720 76 730 86
rect 762 76 772 86
rect 896 76 906 86
rect 938 76 948 86
rect -114 -86 -104 -76
rect -72 -86 -62 -76
rect 62 -86 72 -76
rect 104 -86 114 -76
rect 164 -86 174 -76
rect 206 -86 216 -76
rect 340 -86 350 -76
rect 382 -86 392 -76
rect 442 -86 452 -76
rect 484 -86 494 -76
rect 618 -86 628 -76
rect 660 -86 670 -76
rect 720 -86 730 -76
rect 762 -86 772 -76
rect 896 -86 906 -76
rect 938 -86 948 -76
rect -104 -96 -94 -86
rect -82 -96 -72 -86
rect 72 -96 82 -86
rect 94 -96 104 -86
rect 174 -96 184 -86
rect 196 -96 206 -86
rect 350 -96 360 -86
rect 372 -96 382 -86
rect 452 -96 462 -86
rect 474 -96 484 -86
rect 628 -96 638 -86
rect 650 -96 660 -86
rect 730 -96 740 -86
rect 752 -96 762 -86
rect 906 -96 916 -86
rect 928 -96 938 -86
rect -36 -128 -26 -118
rect 26 -128 36 -118
rect 242 -128 252 -118
rect 304 -128 314 -118
rect 520 -128 530 -118
rect 582 -128 592 -118
rect 798 -128 808 -118
rect 860 -128 870 -118
rect -46 -138 46 -128
rect 232 -138 324 -128
rect 510 -138 602 -128
rect 788 -138 880 -128
rect -36 -150 36 -138
rect 242 -150 314 -138
rect 520 -150 592 -138
rect 798 -150 870 -138
rect -46 -160 46 -150
rect 232 -160 324 -150
rect 510 -160 602 -150
rect 788 -160 880 -150
rect -36 -170 -26 -160
rect 26 -170 36 -160
rect 242 -170 252 -160
rect 304 -170 314 -160
rect 520 -170 530 -160
rect 582 -170 592 -160
rect 798 -170 808 -160
rect 860 -170 870 -160
<< nmos >>
rect -50 -100 50 100
rect 228 -100 328 100
rect 506 -100 606 100
rect 784 -100 884 100
<< ndiff >>
rect -118 86 -50 100
rect -118 -86 -104 86
rect -72 -86 -50 86
rect -118 -100 -50 -86
rect 50 86 118 100
rect 50 -86 72 86
rect 104 -86 118 86
rect 50 -100 118 -86
rect 160 86 228 100
rect 160 -86 174 86
rect 206 -86 228 86
rect 160 -100 228 -86
rect 328 86 396 100
rect 328 -86 350 86
rect 382 -86 396 86
rect 328 -100 396 -86
rect 438 86 506 100
rect 438 -86 452 86
rect 484 -86 506 86
rect 438 -100 506 -86
rect 606 86 674 100
rect 606 -86 628 86
rect 660 -86 674 86
rect 606 -100 674 -86
rect 716 86 784 100
rect 716 -86 730 86
rect 762 -86 784 86
rect 716 -100 784 -86
rect 884 86 952 100
rect 884 -86 906 86
rect 938 -86 952 86
rect 884 -100 952 -86
<< ndiffc >>
rect -104 -86 -72 86
rect 72 -86 104 86
rect 174 -86 206 86
rect 350 -86 382 86
rect 452 -86 484 86
rect 628 -86 660 86
rect 730 -86 762 86
rect 906 -86 938 86
<< psubdiff >>
rect -241 262 1075 276
rect -241 230 -167 262
rect 1001 230 1075 262
rect -241 216 1075 230
rect -241 202 -181 216
rect -241 -202 -227 202
rect -195 -202 -181 202
rect 1015 202 1075 216
rect -241 -216 -181 -202
rect 1015 -202 1029 202
rect 1061 -202 1075 202
rect 1015 -216 1075 -202
rect -241 -230 1075 -216
rect -241 -262 -167 -230
rect 1001 -262 1075 -230
rect -241 -276 1075 -262
<< psubdiffcont >>
rect -167 230 1001 262
rect -227 -202 -195 202
rect 1029 -202 1061 202
rect -167 -262 1001 -230
<< poly >>
rect -50 160 50 174
rect -50 128 -36 160
rect 36 128 50 160
rect -50 100 50 128
rect 228 160 328 174
rect 228 128 242 160
rect 314 128 328 160
rect 228 100 328 128
rect 506 160 606 174
rect 506 128 520 160
rect 592 128 606 160
rect 506 100 606 128
rect 784 160 884 174
rect 784 128 798 160
rect 870 128 884 160
rect 784 100 884 128
rect -50 -128 50 -100
rect -50 -160 -36 -128
rect 36 -160 50 -128
rect -50 -174 50 -160
rect 228 -128 328 -100
rect 228 -160 242 -128
rect 314 -160 328 -128
rect 228 -174 328 -160
rect 506 -128 606 -100
rect 506 -160 520 -128
rect 592 -160 606 -128
rect 506 -174 606 -160
rect 784 -128 884 -100
rect 784 -160 798 -128
rect 870 -160 884 -128
rect 784 -174 884 -160
<< polycont >>
rect -36 128 36 160
rect 242 128 314 160
rect 520 128 592 160
rect 798 128 870 160
rect -36 -160 36 -128
rect 242 -160 314 -128
rect 520 -160 592 -128
rect 798 -160 870 -128
<< metal1 >>
rect -237 262 1071 272
rect -237 230 -167 262
rect 1001 230 1071 262
rect -237 220 1071 230
rect -237 202 -185 220
rect -237 -202 -227 202
rect -195 -202 -185 202
rect 1019 202 1071 220
rect -237 -220 -185 -202
rect 1019 -202 1029 202
rect 1061 -202 1071 202
rect 1019 -220 1071 -202
rect -237 -230 1071 -220
rect -237 -262 -167 -230
rect 1001 -262 1071 -230
rect -237 -272 1071 -262
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 1 l 0.5 nf 1 nx 4 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 1
<< end >>
