magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 50 56 366 292
rect -26 -56 410 56
<< nmos >>
rect 144 118 170 266
rect 246 118 272 266
<< pmos >>
rect 144 412 170 636
rect 212 412 238 636
<< ndiff >>
rect 76 232 144 266
rect 76 200 90 232
rect 122 200 144 232
rect 76 164 144 200
rect 76 132 90 164
rect 122 132 144 164
rect 76 118 144 132
rect 170 232 246 266
rect 170 200 192 232
rect 224 200 246 232
rect 170 164 246 200
rect 170 132 192 164
rect 224 132 246 164
rect 170 118 246 132
rect 272 232 340 266
rect 272 200 294 232
rect 326 200 340 232
rect 272 164 340 200
rect 272 132 294 164
rect 326 132 340 164
rect 272 118 340 132
<< pdiff >>
rect 72 622 144 636
rect 72 590 90 622
rect 122 590 144 622
rect 72 554 144 590
rect 72 522 90 554
rect 122 522 144 554
rect 72 486 144 522
rect 72 454 90 486
rect 122 454 144 486
rect 72 412 144 454
rect 170 412 212 636
rect 238 622 306 636
rect 238 590 260 622
rect 292 590 306 622
rect 238 554 306 590
rect 238 522 260 554
rect 292 522 306 554
rect 238 486 306 522
rect 238 454 260 486
rect 292 454 306 486
rect 238 412 306 454
<< ndiffc >>
rect 90 200 122 232
rect 90 132 122 164
rect 192 200 224 232
rect 192 132 224 164
rect 294 200 326 232
rect 294 132 326 164
<< pdiffc >>
rect 90 590 122 622
rect 90 522 122 554
rect 90 454 122 486
rect 260 590 292 622
rect 260 522 292 554
rect 260 454 292 486
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 144 636 170 672
rect 212 636 238 672
rect 144 370 170 412
rect 70 353 170 370
rect 70 321 87 353
rect 119 321 170 353
rect 70 304 170 321
rect 212 370 238 412
rect 212 353 308 370
rect 212 321 259 353
rect 291 321 308 353
rect 212 304 308 321
rect 144 266 170 304
rect 246 266 272 304
rect 144 82 170 118
rect 246 82 272 118
<< polycont >>
rect 87 321 119 353
rect 259 321 291 353
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 80 622 132 712
rect 80 590 90 622
rect 122 590 132 622
rect 80 554 132 590
rect 80 522 90 554
rect 122 522 132 554
rect 80 486 132 522
rect 250 622 314 632
rect 250 590 260 622
rect 292 590 314 622
rect 250 554 314 590
rect 250 522 260 554
rect 292 522 314 554
rect 250 487 314 522
rect 80 454 90 486
rect 122 454 132 486
rect 80 444 132 454
rect 174 486 314 487
rect 174 454 260 486
rect 292 454 314 486
rect 174 447 314 454
rect 70 353 136 370
rect 70 321 87 353
rect 119 321 136 353
rect 70 304 136 321
rect 174 242 208 447
rect 249 353 316 370
rect 249 321 259 353
rect 291 321 316 353
rect 249 304 316 321
rect 80 232 132 242
rect 80 200 90 232
rect 122 200 132 232
rect 80 164 132 200
rect 80 132 90 164
rect 122 132 132 164
rect 80 44 132 132
rect 174 232 234 242
rect 174 200 192 232
rect 224 200 234 232
rect 174 164 234 200
rect 174 132 192 164
rect 224 132 234 164
rect 174 121 234 132
rect 284 232 336 242
rect 284 200 294 232
rect 326 200 336 232
rect 284 164 336 200
rect 284 132 294 164
rect 326 132 336 164
rect 284 44 336 132
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 70 304 136 370 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 250 447 314 632 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 249 304 316 370 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 219830
string GDS_FILE 6_final.gds
string GDS_START 216064
<< end >>
