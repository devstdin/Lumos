magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2154 2826 5854
<< nwell >>
rect -124 2500 826 3854
rect -124 -154 826 1050
<< pwell >>
rect -5 1756 311 2402
rect -26 1644 728 1756
rect -5 1148 707 1644
<< nmos >>
rect 89 1826 115 2376
<< pmos >>
rect 89 2624 115 3574
<< hvnmos >>
rect 89 1174 179 1554
rect 255 1174 345 1554
rect 523 1174 613 1554
<< hvpmos >>
rect 89 506 179 566
rect 255 506 345 566
rect 523 146 613 926
<< ndiff >>
rect 21 2355 89 2376
rect 21 2323 35 2355
rect 67 2323 89 2355
rect 21 2287 89 2323
rect 21 2255 35 2287
rect 67 2255 89 2287
rect 21 2219 89 2255
rect 21 2187 35 2219
rect 67 2187 89 2219
rect 21 2151 89 2187
rect 21 2119 35 2151
rect 67 2119 89 2151
rect 21 2083 89 2119
rect 21 2051 35 2083
rect 67 2051 89 2083
rect 21 2015 89 2051
rect 21 1983 35 2015
rect 67 1983 89 2015
rect 21 1947 89 1983
rect 21 1915 35 1947
rect 67 1915 89 1947
rect 21 1879 89 1915
rect 21 1847 35 1879
rect 67 1847 89 1879
rect 21 1826 89 1847
rect 115 2321 183 2376
rect 115 2289 137 2321
rect 169 2289 183 2321
rect 115 2253 183 2289
rect 115 2221 137 2253
rect 169 2221 183 2253
rect 115 2185 183 2221
rect 115 2153 137 2185
rect 169 2153 183 2185
rect 115 2117 183 2153
rect 115 2085 137 2117
rect 169 2085 183 2117
rect 115 2049 183 2085
rect 115 2017 137 2049
rect 169 2017 183 2049
rect 115 1981 183 2017
rect 115 1949 137 1981
rect 169 1949 183 1981
rect 115 1913 183 1949
rect 115 1881 137 1913
rect 169 1881 183 1913
rect 115 1826 183 1881
rect 225 2355 285 2376
rect 225 2323 239 2355
rect 271 2323 285 2355
rect 225 2287 285 2323
rect 225 2255 239 2287
rect 271 2255 285 2287
rect 225 2219 285 2255
rect 225 2187 239 2219
rect 271 2187 285 2219
rect 225 2151 285 2187
rect 225 2119 239 2151
rect 271 2119 285 2151
rect 225 2083 285 2119
rect 225 2051 239 2083
rect 271 2051 285 2083
rect 225 2015 285 2051
rect 225 1983 239 2015
rect 271 1983 285 2015
rect 225 1947 285 1983
rect 225 1915 239 1947
rect 271 1915 285 1947
rect 225 1879 285 1915
rect 225 1847 239 1879
rect 271 1847 285 1879
rect 225 1826 285 1847
<< pdiff >>
rect 21 3557 89 3574
rect 21 3525 35 3557
rect 67 3525 89 3557
rect 21 3489 89 3525
rect 21 3457 35 3489
rect 67 3457 89 3489
rect 21 3421 89 3457
rect 21 3389 35 3421
rect 67 3389 89 3421
rect 21 3353 89 3389
rect 21 3321 35 3353
rect 67 3321 89 3353
rect 21 3285 89 3321
rect 21 3253 35 3285
rect 67 3253 89 3285
rect 21 3217 89 3253
rect 21 3185 35 3217
rect 67 3185 89 3217
rect 21 3149 89 3185
rect 21 3117 35 3149
rect 67 3117 89 3149
rect 21 3081 89 3117
rect 21 3049 35 3081
rect 67 3049 89 3081
rect 21 3013 89 3049
rect 21 2981 35 3013
rect 67 2981 89 3013
rect 21 2945 89 2981
rect 21 2913 35 2945
rect 67 2913 89 2945
rect 21 2877 89 2913
rect 21 2845 35 2877
rect 67 2845 89 2877
rect 21 2809 89 2845
rect 21 2777 35 2809
rect 67 2777 89 2809
rect 21 2741 89 2777
rect 21 2709 35 2741
rect 67 2709 89 2741
rect 21 2673 89 2709
rect 21 2641 35 2673
rect 67 2641 89 2673
rect 21 2624 89 2641
rect 115 3523 183 3574
rect 115 3491 137 3523
rect 169 3491 183 3523
rect 115 3455 183 3491
rect 115 3423 137 3455
rect 169 3423 183 3455
rect 115 3387 183 3423
rect 115 3355 137 3387
rect 169 3355 183 3387
rect 115 3319 183 3355
rect 115 3287 137 3319
rect 169 3287 183 3319
rect 115 3251 183 3287
rect 115 3219 137 3251
rect 169 3219 183 3251
rect 115 3183 183 3219
rect 115 3151 137 3183
rect 169 3151 183 3183
rect 115 3115 183 3151
rect 115 3083 137 3115
rect 169 3083 183 3115
rect 115 3047 183 3083
rect 115 3015 137 3047
rect 169 3015 183 3047
rect 115 2979 183 3015
rect 115 2947 137 2979
rect 169 2947 183 2979
rect 115 2911 183 2947
rect 115 2879 137 2911
rect 169 2879 183 2911
rect 115 2843 183 2879
rect 115 2811 137 2843
rect 169 2811 183 2843
rect 115 2775 183 2811
rect 115 2743 137 2775
rect 169 2743 183 2775
rect 115 2707 183 2743
rect 115 2675 137 2707
rect 169 2675 183 2707
rect 115 2624 183 2675
rect 225 3557 285 3574
rect 225 3525 239 3557
rect 271 3525 285 3557
rect 225 3489 285 3525
rect 225 3457 239 3489
rect 271 3457 285 3489
rect 225 3421 285 3457
rect 225 3389 239 3421
rect 271 3389 285 3421
rect 225 3353 285 3389
rect 225 3321 239 3353
rect 271 3321 285 3353
rect 225 3285 285 3321
rect 225 3253 239 3285
rect 271 3253 285 3285
rect 225 3217 285 3253
rect 225 3185 239 3217
rect 271 3185 285 3217
rect 225 3149 285 3185
rect 225 3117 239 3149
rect 271 3117 285 3149
rect 225 3081 285 3117
rect 225 3049 239 3081
rect 271 3049 285 3081
rect 225 3013 285 3049
rect 225 2981 239 3013
rect 271 2981 285 3013
rect 225 2945 285 2981
rect 225 2913 239 2945
rect 271 2913 285 2945
rect 225 2877 285 2913
rect 225 2845 239 2877
rect 271 2845 285 2877
rect 225 2809 285 2845
rect 225 2777 239 2809
rect 271 2777 285 2809
rect 225 2741 285 2777
rect 225 2709 239 2741
rect 271 2709 285 2741
rect 225 2673 285 2709
rect 225 2641 239 2673
rect 271 2641 285 2673
rect 225 2624 285 2641
<< hvndiff >>
rect 21 1516 89 1554
rect 21 1484 35 1516
rect 67 1484 89 1516
rect 21 1448 89 1484
rect 21 1416 35 1448
rect 67 1416 89 1448
rect 21 1380 89 1416
rect 21 1348 35 1380
rect 67 1348 89 1380
rect 21 1312 89 1348
rect 21 1280 35 1312
rect 67 1280 89 1312
rect 21 1244 89 1280
rect 21 1212 35 1244
rect 67 1212 89 1244
rect 21 1174 89 1212
rect 179 1516 255 1554
rect 179 1484 201 1516
rect 233 1484 255 1516
rect 179 1448 255 1484
rect 179 1416 201 1448
rect 233 1416 255 1448
rect 179 1380 255 1416
rect 179 1348 201 1380
rect 233 1348 255 1380
rect 179 1312 255 1348
rect 179 1280 201 1312
rect 233 1280 255 1312
rect 179 1244 255 1280
rect 179 1212 201 1244
rect 233 1212 255 1244
rect 179 1174 255 1212
rect 345 1516 413 1554
rect 345 1484 367 1516
rect 399 1484 413 1516
rect 345 1448 413 1484
rect 345 1416 367 1448
rect 399 1416 413 1448
rect 345 1380 413 1416
rect 345 1348 367 1380
rect 399 1348 413 1380
rect 345 1312 413 1348
rect 345 1280 367 1312
rect 399 1280 413 1312
rect 345 1244 413 1280
rect 345 1212 367 1244
rect 399 1212 413 1244
rect 345 1174 413 1212
rect 455 1516 523 1554
rect 455 1484 469 1516
rect 501 1484 523 1516
rect 455 1448 523 1484
rect 455 1416 469 1448
rect 501 1416 523 1448
rect 455 1380 523 1416
rect 455 1348 469 1380
rect 501 1348 523 1380
rect 455 1312 523 1348
rect 455 1280 469 1312
rect 501 1280 523 1312
rect 455 1244 523 1280
rect 455 1212 469 1244
rect 501 1212 523 1244
rect 455 1174 523 1212
rect 613 1516 681 1554
rect 613 1484 635 1516
rect 667 1484 681 1516
rect 613 1448 681 1484
rect 613 1416 635 1448
rect 667 1416 681 1448
rect 613 1380 681 1416
rect 613 1348 635 1380
rect 667 1348 681 1380
rect 613 1312 681 1348
rect 613 1280 635 1312
rect 667 1280 681 1312
rect 613 1244 681 1280
rect 613 1212 635 1244
rect 667 1212 681 1244
rect 613 1174 681 1212
<< hvpdiff >>
rect 455 892 523 926
rect 455 860 469 892
rect 501 860 523 892
rect 455 824 523 860
rect 455 792 469 824
rect 501 792 523 824
rect 455 756 523 792
rect 455 724 469 756
rect 501 724 523 756
rect 455 688 523 724
rect 455 656 469 688
rect 501 656 523 688
rect 455 620 523 656
rect 455 588 469 620
rect 501 588 523 620
rect 21 552 89 566
rect 21 520 35 552
rect 67 520 89 552
rect 21 506 89 520
rect 179 552 255 566
rect 179 520 201 552
rect 233 520 255 552
rect 179 506 255 520
rect 345 552 413 566
rect 345 520 367 552
rect 399 520 413 552
rect 345 506 413 520
rect 455 552 523 588
rect 455 520 469 552
rect 501 520 523 552
rect 455 484 523 520
rect 455 452 469 484
rect 501 452 523 484
rect 455 416 523 452
rect 455 384 469 416
rect 501 384 523 416
rect 455 348 523 384
rect 455 316 469 348
rect 501 316 523 348
rect 455 280 523 316
rect 455 248 469 280
rect 501 248 523 280
rect 455 212 523 248
rect 455 180 469 212
rect 501 180 523 212
rect 455 146 523 180
rect 613 892 681 926
rect 613 860 635 892
rect 667 860 681 892
rect 613 824 681 860
rect 613 792 635 824
rect 667 792 681 824
rect 613 756 681 792
rect 613 724 635 756
rect 667 724 681 756
rect 613 688 681 724
rect 613 656 635 688
rect 667 656 681 688
rect 613 620 681 656
rect 613 588 635 620
rect 667 588 681 620
rect 613 552 681 588
rect 613 520 635 552
rect 667 520 681 552
rect 613 484 681 520
rect 613 452 635 484
rect 667 452 681 484
rect 613 416 681 452
rect 613 384 635 416
rect 667 384 681 416
rect 613 348 681 384
rect 613 316 635 348
rect 667 316 681 348
rect 613 280 681 316
rect 613 248 635 280
rect 667 248 681 280
rect 613 212 681 248
rect 613 180 635 212
rect 667 180 681 212
rect 613 146 681 180
<< ndiffc >>
rect 35 2323 67 2355
rect 35 2255 67 2287
rect 35 2187 67 2219
rect 35 2119 67 2151
rect 35 2051 67 2083
rect 35 1983 67 2015
rect 35 1915 67 1947
rect 35 1847 67 1879
rect 137 2289 169 2321
rect 137 2221 169 2253
rect 137 2153 169 2185
rect 137 2085 169 2117
rect 137 2017 169 2049
rect 137 1949 169 1981
rect 137 1881 169 1913
rect 239 2323 271 2355
rect 239 2255 271 2287
rect 239 2187 271 2219
rect 239 2119 271 2151
rect 239 2051 271 2083
rect 239 1983 271 2015
rect 239 1915 271 1947
rect 239 1847 271 1879
<< pdiffc >>
rect 35 3525 67 3557
rect 35 3457 67 3489
rect 35 3389 67 3421
rect 35 3321 67 3353
rect 35 3253 67 3285
rect 35 3185 67 3217
rect 35 3117 67 3149
rect 35 3049 67 3081
rect 35 2981 67 3013
rect 35 2913 67 2945
rect 35 2845 67 2877
rect 35 2777 67 2809
rect 35 2709 67 2741
rect 35 2641 67 2673
rect 137 3491 169 3523
rect 137 3423 169 3455
rect 137 3355 169 3387
rect 137 3287 169 3319
rect 137 3219 169 3251
rect 137 3151 169 3183
rect 137 3083 169 3115
rect 137 3015 169 3047
rect 137 2947 169 2979
rect 137 2879 169 2911
rect 137 2811 169 2843
rect 137 2743 169 2775
rect 137 2675 169 2707
rect 239 3525 271 3557
rect 239 3457 271 3489
rect 239 3389 271 3421
rect 239 3321 271 3353
rect 239 3253 271 3285
rect 239 3185 271 3217
rect 239 3117 271 3149
rect 239 3049 271 3081
rect 239 2981 271 3013
rect 239 2913 271 2945
rect 239 2845 271 2877
rect 239 2777 271 2809
rect 239 2709 271 2741
rect 239 2641 271 2673
<< hvndiffc >>
rect 35 1484 67 1516
rect 35 1416 67 1448
rect 35 1348 67 1380
rect 35 1280 67 1312
rect 35 1212 67 1244
rect 201 1484 233 1516
rect 201 1416 233 1448
rect 201 1348 233 1380
rect 201 1280 233 1312
rect 201 1212 233 1244
rect 367 1484 399 1516
rect 367 1416 399 1448
rect 367 1348 399 1380
rect 367 1280 399 1312
rect 367 1212 399 1244
rect 469 1484 501 1516
rect 469 1416 501 1448
rect 469 1348 501 1380
rect 469 1280 501 1312
rect 469 1212 501 1244
rect 635 1484 667 1516
rect 635 1416 667 1448
rect 635 1348 667 1380
rect 635 1280 667 1312
rect 635 1212 667 1244
<< hvpdiffc >>
rect 469 860 501 892
rect 469 792 501 824
rect 469 724 501 756
rect 469 656 501 688
rect 469 588 501 620
rect 35 520 67 552
rect 201 520 233 552
rect 367 520 399 552
rect 469 520 501 552
rect 469 452 501 484
rect 469 384 501 416
rect 469 316 501 348
rect 469 248 501 280
rect 469 180 501 212
rect 635 860 667 892
rect 635 792 667 824
rect 635 724 667 756
rect 635 656 667 688
rect 635 588 667 620
rect 635 520 667 552
rect 635 452 667 484
rect 635 384 667 416
rect 635 316 667 348
rect 635 248 667 280
rect 635 180 667 212
<< psubdiff >>
rect 0 1716 702 1730
rect 0 1684 63 1716
rect 95 1684 131 1716
rect 163 1684 199 1716
rect 231 1684 267 1716
rect 299 1684 335 1716
rect 367 1684 403 1716
rect 435 1684 471 1716
rect 503 1684 539 1716
rect 571 1684 607 1716
rect 639 1684 702 1716
rect 0 1670 702 1684
<< nsubdiff >>
rect 0 3716 702 3730
rect 0 3684 63 3716
rect 95 3684 131 3716
rect 163 3684 199 3716
rect 231 3684 267 3716
rect 299 3684 335 3716
rect 367 3684 403 3716
rect 435 3684 471 3716
rect 503 3684 539 3716
rect 571 3684 607 3716
rect 639 3684 702 3716
rect 0 3670 702 3684
rect 0 16 702 30
rect 0 -16 63 16
rect 95 -16 131 16
rect 163 -16 199 16
rect 231 -16 267 16
rect 299 -16 335 16
rect 367 -16 403 16
rect 435 -16 471 16
rect 503 -16 539 16
rect 571 -16 607 16
rect 639 -16 702 16
rect 0 -30 702 -16
<< psubdiffcont >>
rect 63 1684 95 1716
rect 131 1684 163 1716
rect 199 1684 231 1716
rect 267 1684 299 1716
rect 335 1684 367 1716
rect 403 1684 435 1716
rect 471 1684 503 1716
rect 539 1684 571 1716
rect 607 1684 639 1716
<< nsubdiffcont >>
rect 63 3684 95 3716
rect 131 3684 163 3716
rect 199 3684 231 3716
rect 267 3684 299 3716
rect 335 3684 367 3716
rect 403 3684 435 3716
rect 471 3684 503 3716
rect 539 3684 571 3716
rect 607 3684 639 3716
rect 63 -16 95 16
rect 131 -16 163 16
rect 199 -16 231 16
rect 267 -16 299 16
rect 335 -16 367 16
rect 403 -16 435 16
rect 471 -16 503 16
rect 539 -16 571 16
rect 607 -16 639 16
<< poly >>
rect 89 3574 115 3610
rect 89 2530 115 2624
rect 89 2516 165 2530
rect 89 2484 119 2516
rect 151 2484 165 2516
rect 89 2470 165 2484
rect 89 2376 115 2470
rect 89 1790 115 1826
rect 89 1554 179 1590
rect 255 1554 345 1590
rect 523 1554 613 1590
rect 89 1144 179 1174
rect 89 1112 133 1144
rect 165 1112 179 1144
rect 89 1098 179 1112
rect 255 1144 345 1174
rect 255 1112 269 1144
rect 301 1112 345 1144
rect 255 1098 345 1112
rect 523 1066 613 1174
rect 523 1034 537 1066
rect 569 1034 613 1066
rect 523 926 613 1034
rect 255 736 345 750
rect 255 704 269 736
rect 301 704 345 736
rect 89 636 179 650
rect 89 604 133 636
rect 165 604 179 636
rect 89 566 179 604
rect 255 566 345 704
rect 89 470 179 506
rect 255 470 345 506
rect 523 110 613 146
<< polycont >>
rect 119 2484 151 2516
rect 133 1112 165 1144
rect 269 1112 301 1144
rect 537 1034 569 1066
rect 269 704 301 736
rect 133 604 165 636
<< metal1 >>
rect 0 3716 702 3721
rect 0 3684 63 3716
rect 95 3684 131 3716
rect 163 3684 199 3716
rect 231 3684 267 3716
rect 299 3684 335 3716
rect 367 3684 403 3716
rect 435 3684 471 3716
rect 503 3684 539 3716
rect 571 3684 607 3716
rect 639 3684 702 3716
rect 0 3679 702 3684
rect 25 3557 67 3573
rect 25 3542 35 3557
rect 25 1862 26 3542
rect 66 3489 67 3525
rect 66 3421 67 3457
rect 66 3353 67 3389
rect 66 3285 67 3321
rect 66 3217 67 3253
rect 66 3149 67 3185
rect 66 3081 67 3117
rect 66 3013 67 3049
rect 66 2945 67 2981
rect 66 2877 67 2913
rect 66 2809 67 2845
rect 66 2741 67 2777
rect 66 2673 67 2709
rect 137 3523 169 3679
rect 137 3455 169 3491
rect 137 3387 169 3423
rect 137 3319 169 3355
rect 137 3251 169 3287
rect 137 3183 169 3219
rect 137 3115 169 3151
rect 137 3047 169 3083
rect 137 2979 169 3015
rect 137 2911 169 2947
rect 137 2843 169 2879
rect 137 2775 169 2811
rect 137 2707 169 2743
rect 137 2642 169 2675
rect 234 3557 276 3573
rect 234 3542 239 3557
rect 271 3542 276 3557
rect 66 2355 67 2641
rect 234 2606 235 3542
rect 119 2516 235 2606
rect 151 2484 235 2516
rect 119 2394 235 2484
rect 66 2287 67 2323
rect 66 2219 67 2255
rect 66 2151 67 2187
rect 66 2083 67 2119
rect 66 2015 67 2051
rect 66 1947 67 1983
rect 66 1879 67 1915
rect 25 1847 35 1862
rect 25 1831 67 1847
rect 137 2321 169 2358
rect 137 2253 169 2289
rect 137 2185 169 2221
rect 137 2117 169 2153
rect 137 2049 169 2085
rect 137 1981 169 2017
rect 137 1913 169 1949
rect 137 1721 169 1881
rect 234 1862 235 2394
rect 275 1862 276 3542
rect 234 1847 239 1862
rect 271 1847 276 1862
rect 234 1831 276 1847
rect 0 1716 702 1721
rect 0 1684 63 1716
rect 95 1684 131 1716
rect 163 1684 199 1716
rect 231 1684 267 1716
rect 299 1684 335 1716
rect 367 1684 403 1716
rect 435 1684 471 1716
rect 503 1684 539 1716
rect 571 1684 607 1716
rect 639 1684 702 1716
rect 0 1679 702 1684
rect 35 1516 67 1532
rect 35 1448 67 1484
rect 35 1380 67 1416
rect 35 1312 67 1348
rect 35 1244 67 1280
rect 35 752 67 1212
rect 201 1516 233 1679
rect 201 1448 233 1484
rect 201 1380 233 1416
rect 201 1312 233 1348
rect 201 1244 233 1280
rect 201 1196 233 1212
rect 367 1516 399 1532
rect 367 1448 399 1484
rect 367 1380 399 1416
rect 367 1312 399 1348
rect 367 1244 399 1280
rect 133 1151 175 1160
rect 133 1144 134 1151
rect 133 1029 134 1112
rect 174 1029 175 1151
rect 133 1020 175 1029
rect 259 1151 301 1160
rect 259 1029 260 1151
rect 300 1144 301 1151
rect 300 1029 301 1112
rect 259 1020 301 1029
rect 367 1082 399 1212
rect 469 1516 501 1679
rect 469 1448 501 1484
rect 469 1380 501 1416
rect 469 1312 501 1348
rect 469 1244 501 1280
rect 469 1196 501 1212
rect 635 1516 677 1532
rect 667 1484 677 1516
rect 635 1483 677 1484
rect 635 1448 636 1483
rect 635 1380 636 1416
rect 635 1312 636 1348
rect 635 1244 636 1280
rect 367 1066 569 1082
rect 367 1034 537 1066
rect 367 1018 569 1034
rect 35 736 301 752
rect 35 704 269 736
rect 35 688 301 704
rect 35 552 67 688
rect 367 652 399 1018
rect 133 636 399 652
rect 165 604 399 636
rect 133 588 399 604
rect 367 552 399 588
rect 35 504 67 520
rect 185 520 201 552
rect 233 520 249 552
rect 185 21 249 520
rect 367 504 399 520
rect 469 892 501 908
rect 469 824 501 860
rect 469 756 501 792
rect 469 688 501 724
rect 469 620 501 656
rect 469 552 501 588
rect 469 484 501 520
rect 469 416 501 452
rect 469 348 501 384
rect 469 280 501 316
rect 469 212 501 248
rect 469 21 501 180
rect 635 892 636 1212
rect 635 824 636 860
rect 635 756 636 792
rect 635 688 636 724
rect 635 620 636 656
rect 635 552 636 588
rect 635 484 636 520
rect 635 416 636 452
rect 635 348 636 384
rect 635 280 636 316
rect 635 213 636 248
rect 676 213 677 1483
rect 635 212 677 213
rect 667 180 677 212
rect 635 164 677 180
rect 0 16 702 21
rect 0 -16 63 16
rect 95 -16 131 16
rect 163 -16 199 16
rect 231 -16 267 16
rect 299 -16 335 16
rect 367 -16 403 16
rect 435 -16 471 16
rect 503 -16 539 16
rect 571 -16 607 16
rect 639 -16 702 16
rect 0 -21 702 -16
<< via1 >>
rect 26 3525 35 3542
rect 35 3525 66 3542
rect 26 3489 66 3525
rect 26 3457 35 3489
rect 35 3457 66 3489
rect 26 3421 66 3457
rect 26 3389 35 3421
rect 35 3389 66 3421
rect 26 3353 66 3389
rect 26 3321 35 3353
rect 35 3321 66 3353
rect 26 3285 66 3321
rect 26 3253 35 3285
rect 35 3253 66 3285
rect 26 3217 66 3253
rect 26 3185 35 3217
rect 35 3185 66 3217
rect 26 3149 66 3185
rect 26 3117 35 3149
rect 35 3117 66 3149
rect 26 3081 66 3117
rect 26 3049 35 3081
rect 35 3049 66 3081
rect 26 3013 66 3049
rect 26 2981 35 3013
rect 35 2981 66 3013
rect 26 2945 66 2981
rect 26 2913 35 2945
rect 35 2913 66 2945
rect 26 2877 66 2913
rect 26 2845 35 2877
rect 35 2845 66 2877
rect 26 2809 66 2845
rect 26 2777 35 2809
rect 35 2777 66 2809
rect 26 2741 66 2777
rect 26 2709 35 2741
rect 35 2709 66 2741
rect 26 2673 66 2709
rect 26 2641 35 2673
rect 35 2641 66 2673
rect 26 2355 66 2641
rect 235 3525 239 3542
rect 239 3525 271 3542
rect 271 3525 275 3542
rect 235 3489 275 3525
rect 235 3457 239 3489
rect 239 3457 271 3489
rect 271 3457 275 3489
rect 235 3421 275 3457
rect 235 3389 239 3421
rect 239 3389 271 3421
rect 271 3389 275 3421
rect 235 3353 275 3389
rect 235 3321 239 3353
rect 239 3321 271 3353
rect 271 3321 275 3353
rect 235 3285 275 3321
rect 235 3253 239 3285
rect 239 3253 271 3285
rect 271 3253 275 3285
rect 235 3217 275 3253
rect 235 3185 239 3217
rect 239 3185 271 3217
rect 271 3185 275 3217
rect 235 3149 275 3185
rect 235 3117 239 3149
rect 239 3117 271 3149
rect 271 3117 275 3149
rect 235 3081 275 3117
rect 235 3049 239 3081
rect 239 3049 271 3081
rect 271 3049 275 3081
rect 235 3013 275 3049
rect 235 2981 239 3013
rect 239 2981 271 3013
rect 271 2981 275 3013
rect 235 2945 275 2981
rect 235 2913 239 2945
rect 239 2913 271 2945
rect 271 2913 275 2945
rect 235 2877 275 2913
rect 235 2845 239 2877
rect 239 2845 271 2877
rect 271 2845 275 2877
rect 235 2809 275 2845
rect 235 2777 239 2809
rect 239 2777 271 2809
rect 271 2777 275 2809
rect 235 2741 275 2777
rect 235 2709 239 2741
rect 239 2709 271 2741
rect 271 2709 275 2741
rect 235 2673 275 2709
rect 235 2641 239 2673
rect 239 2641 271 2673
rect 271 2641 275 2673
rect 26 2323 35 2355
rect 35 2323 66 2355
rect 26 2287 66 2323
rect 26 2255 35 2287
rect 35 2255 66 2287
rect 26 2219 66 2255
rect 26 2187 35 2219
rect 35 2187 66 2219
rect 26 2151 66 2187
rect 26 2119 35 2151
rect 35 2119 66 2151
rect 26 2083 66 2119
rect 26 2051 35 2083
rect 35 2051 66 2083
rect 26 2015 66 2051
rect 26 1983 35 2015
rect 35 1983 66 2015
rect 26 1947 66 1983
rect 26 1915 35 1947
rect 35 1915 66 1947
rect 26 1879 66 1915
rect 26 1862 35 1879
rect 35 1862 66 1879
rect 235 2355 275 2641
rect 235 2323 239 2355
rect 239 2323 271 2355
rect 271 2323 275 2355
rect 235 2287 275 2323
rect 235 2255 239 2287
rect 239 2255 271 2287
rect 271 2255 275 2287
rect 235 2219 275 2255
rect 235 2187 239 2219
rect 239 2187 271 2219
rect 271 2187 275 2219
rect 235 2151 275 2187
rect 235 2119 239 2151
rect 239 2119 271 2151
rect 271 2119 275 2151
rect 235 2083 275 2119
rect 235 2051 239 2083
rect 239 2051 271 2083
rect 271 2051 275 2083
rect 235 2015 275 2051
rect 235 1983 239 2015
rect 239 1983 271 2015
rect 271 1983 275 2015
rect 235 1947 275 1983
rect 235 1915 239 1947
rect 239 1915 271 1947
rect 271 1915 275 1947
rect 235 1879 275 1915
rect 235 1862 239 1879
rect 239 1862 271 1879
rect 271 1862 275 1879
rect 134 1144 174 1151
rect 134 1112 165 1144
rect 165 1112 174 1144
rect 134 1029 174 1112
rect 260 1144 300 1151
rect 260 1112 269 1144
rect 269 1112 300 1144
rect 260 1029 300 1112
rect 636 1448 676 1483
rect 636 1416 667 1448
rect 667 1416 676 1448
rect 636 1380 676 1416
rect 636 1348 667 1380
rect 667 1348 676 1380
rect 636 1312 676 1348
rect 636 1280 667 1312
rect 667 1280 676 1312
rect 636 1244 676 1280
rect 636 1212 667 1244
rect 667 1212 676 1244
rect 636 892 676 1212
rect 636 860 667 892
rect 667 860 676 892
rect 636 824 676 860
rect 636 792 667 824
rect 667 792 676 824
rect 636 756 676 792
rect 636 724 667 756
rect 667 724 676 756
rect 636 688 676 724
rect 636 656 667 688
rect 667 656 676 688
rect 636 620 676 656
rect 636 588 667 620
rect 667 588 676 620
rect 636 552 676 588
rect 636 520 667 552
rect 667 520 676 552
rect 636 484 676 520
rect 636 452 667 484
rect 667 452 676 484
rect 636 416 676 452
rect 636 384 667 416
rect 667 384 676 416
rect 636 348 676 384
rect 636 316 667 348
rect 667 316 676 348
rect 636 280 676 316
rect 636 248 667 280
rect 667 248 676 280
rect 636 213 676 248
<< metal2 >>
rect 26 3542 66 3551
rect 235 3542 275 3551
rect 26 900 66 1862
rect 134 1862 235 1873
rect 134 1833 275 1862
rect 134 1151 174 1833
rect 636 1483 676 1492
rect 134 1020 174 1029
rect 260 1151 300 1160
rect 260 900 300 1029
rect 26 860 300 900
rect 636 204 676 213
<< labels >>
rlabel metal2 s 636 204 676 1492 4 o
port 5 nsew
rlabel metal2 s 235 1853 275 3551 4 i
port 4 nsew
rlabel metal1 s 0 -21 702 21 4 iovdd
port 2 nsew
rlabel metal1 s 0 1679 702 1721 4 vss
port 3 nsew
rlabel metal1 s 0 3679 702 3721 4 vdd
port 1 nsew
flabel comment s 650 1702 650 1702 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 29659868
string GDS_FILE sg13g2_io.gds
string GDS_START 29642100
<< end >>
