magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 19 56 437 314
rect -26 -56 506 56
<< nmos >>
rect 113 160 139 288
rect 215 160 241 288
rect 317 140 343 288
<< pmos >>
rect 113 468 139 636
rect 215 468 241 636
rect 317 412 343 636
<< ndiff >>
rect 45 268 113 288
rect 45 236 59 268
rect 91 236 113 268
rect 45 160 113 236
rect 139 160 215 288
rect 241 214 317 288
rect 241 182 263 214
rect 295 182 317 214
rect 241 160 317 182
rect 271 140 317 160
rect 343 254 411 288
rect 343 222 365 254
rect 397 222 411 254
rect 343 186 411 222
rect 343 154 365 186
rect 397 154 411 186
rect 343 140 411 154
<< pdiff >>
rect 45 622 113 636
rect 45 590 59 622
rect 91 590 113 622
rect 45 554 113 590
rect 45 522 59 554
rect 91 522 113 554
rect 45 468 113 522
rect 139 622 215 636
rect 139 590 161 622
rect 193 590 215 622
rect 139 554 215 590
rect 139 522 161 554
rect 193 522 215 554
rect 139 468 215 522
rect 241 622 317 636
rect 241 590 263 622
rect 295 590 317 622
rect 241 554 317 590
rect 241 522 263 554
rect 295 522 317 554
rect 241 468 317 522
rect 271 412 317 468
rect 343 622 411 636
rect 343 590 365 622
rect 397 590 411 622
rect 343 554 411 590
rect 343 522 365 554
rect 397 522 411 554
rect 343 486 411 522
rect 343 454 365 486
rect 397 454 411 486
rect 343 412 411 454
<< ndiffc >>
rect 59 236 91 268
rect 263 182 295 214
rect 365 222 397 254
rect 365 154 397 186
<< pdiffc >>
rect 59 590 91 622
rect 59 522 91 554
rect 161 590 193 622
rect 161 522 193 554
rect 263 590 295 622
rect 263 522 295 554
rect 365 590 397 622
rect 365 522 397 554
rect 365 454 397 486
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 113 636 139 672
rect 215 636 241 672
rect 317 636 343 672
rect 113 288 139 468
rect 215 377 241 468
rect 317 377 343 412
rect 178 363 241 377
rect 178 331 192 363
rect 224 331 241 363
rect 178 317 241 331
rect 291 363 352 377
rect 291 331 306 363
rect 338 331 352 363
rect 291 317 352 331
rect 215 288 241 317
rect 317 288 343 317
rect 113 146 139 160
rect 21 128 155 146
rect 21 96 38 128
rect 70 96 106 128
rect 138 96 155 128
rect 215 124 241 160
rect 317 104 343 140
rect 21 82 155 96
<< polycont >>
rect 192 331 224 363
rect 306 331 338 363
rect 38 96 70 128
rect 106 96 138 128
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 49 622 101 712
rect 49 590 59 622
rect 91 590 101 622
rect 49 554 101 590
rect 49 522 59 554
rect 91 522 101 554
rect 49 512 101 522
rect 151 622 203 632
rect 151 590 161 622
rect 193 590 203 622
rect 151 554 203 590
rect 151 522 161 554
rect 193 522 203 554
rect 151 448 203 522
rect 253 622 305 712
rect 253 590 263 622
rect 295 590 305 622
rect 253 554 305 590
rect 253 522 263 554
rect 295 522 305 554
rect 253 512 305 522
rect 355 622 455 632
rect 355 590 365 622
rect 397 590 455 622
rect 355 554 455 590
rect 355 522 365 554
rect 397 522 455 554
rect 355 486 455 522
rect 355 454 365 486
rect 397 454 455 486
rect 49 410 312 448
rect 355 428 455 454
rect 49 268 101 410
rect 156 363 234 374
rect 156 331 192 363
rect 224 331 234 363
rect 156 287 234 331
rect 280 373 312 410
rect 280 363 348 373
rect 280 331 306 363
rect 338 331 348 363
rect 280 321 348 331
rect 49 236 59 268
rect 91 236 101 268
rect 408 264 455 428
rect 49 228 101 236
rect 355 254 455 264
rect 253 214 305 231
rect 21 128 156 192
rect 21 96 38 128
rect 70 96 106 128
rect 138 96 156 128
rect 21 81 156 96
rect 253 182 263 214
rect 295 182 305 214
rect 253 44 305 182
rect 355 222 365 254
rect 397 222 455 254
rect 355 186 455 222
rect 355 154 365 186
rect 397 154 455 186
rect 355 144 455 154
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 355 428 455 632 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 156 287 234 374 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 s 21 81 156 192 0 FreeSans 400 0 0 0 A
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 132386
string GDS_FILE 6_final.gds
string GDS_START 128092
<< end >>
