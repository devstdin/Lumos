magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757363851
<< error_s >>
rect -8630 10 -8474 38
rect -8582 -38 -8522 -10
rect -8582 -641 -8522 -614
rect -8630 -689 -8474 -662
<< psubdiff >>
rect -9338 -41 -9278 -10
rect -9338 -641 -9278 -613
<< nsubdiff >>
rect -8582 -39 -8522 -10
rect -8582 -641 -8522 -613
<< metal1 >>
rect -9524 -641 -9264 -10
rect -8893 -71 -8673 -61
rect -8893 -145 -8883 -71
rect -8683 -145 -8673 -71
rect -8893 -155 -8673 -145
rect -9004 -409 -8938 -201
rect -8893 -347 -8673 -337
rect -8893 -433 -8883 -347
rect -8683 -433 -8673 -347
rect -8893 -443 -8673 -433
rect -9004 -499 -8938 -489
rect -9004 -608 -8994 -499
rect -8948 -608 -8938 -499
rect -9004 -618 -8938 -608
rect -8596 -641 -8432 -10
rect -8375 -127 -8221 -10
rect -8375 -179 -7785 -127
rect -8375 -727 -8221 -179
rect -8075 -232 -7983 -222
rect -8075 -292 -8065 -232
rect -7993 -292 -7983 -232
rect -8184 -303 -8119 -293
rect -8075 -302 -7983 -292
rect -8184 -364 -8174 -303
rect -8129 -364 -8119 -303
rect -8184 -374 -8119 -364
rect -7943 -369 -7883 -309
rect -8075 -422 -7983 -376
rect -8075 -483 -8065 -422
rect -7993 -483 -7983 -422
rect -8075 -530 -7983 -483
rect -8184 -545 -8119 -535
rect -8184 -620 -8174 -545
rect -8129 -620 -8119 -545
rect -7943 -597 -7883 -537
rect -8184 -630 -8119 -620
rect -8075 -727 -7983 -604
rect -7837 -727 -7785 -179
rect -8375 -779 -7785 -727
<< via1 >>
rect -8883 -145 -8683 -71
rect -8883 -433 -8683 -347
rect -8994 -608 -8948 -499
rect -8065 -292 -7993 -232
rect -8174 -364 -8129 -303
rect -8065 -483 -7993 -422
rect -8174 -620 -8129 -545
<< metal2 >>
rect -8893 -71 -8376 -61
rect -8893 -145 -8883 -71
rect -8683 -111 -8376 -71
rect -8683 -145 -8673 -111
rect -8893 -155 -8673 -145
rect -8426 -247 -8376 -111
rect -8075 -232 -7836 -198
rect -8426 -293 -8119 -247
rect -8184 -303 -8119 -293
rect -8075 -292 -8065 -232
rect -7993 -279 -7836 -232
rect -7993 -292 -7983 -279
rect -8075 -302 -7983 -292
rect -8893 -347 -8375 -337
rect -8893 -433 -8883 -347
rect -8683 -391 -8375 -347
rect -8184 -364 -8174 -303
rect -8129 -364 -8119 -303
rect -8184 -374 -8119 -364
rect -8683 -433 -8673 -391
rect -8893 -443 -8673 -433
rect -9004 -499 -8938 -489
rect -9004 -537 -8994 -499
rect -9524 -608 -8994 -537
rect -8948 -608 -8938 -499
rect -9524 -618 -8938 -608
rect -8429 -556 -8375 -391
rect -8075 -422 -7836 -412
rect -8075 -483 -8065 -422
rect -7993 -483 -7836 -422
rect -8075 -493 -7836 -483
rect -8184 -545 -8119 -535
rect -8184 -556 -8174 -545
rect -8429 -610 -8174 -556
rect -8184 -620 -8174 -610
rect -8129 -620 -8119 -545
rect -8184 -630 -8119 -620
use lvnmos_HKFTVP  lvnmos_HKFTVP_0
timestamp 1752931916
transform 0 1 -8029 -1 0 -339
box -93 -248 93 248
use lvnmos_HKFTVP  lvnmos_HKFTVP_1
timestamp 1752931916
transform 0 1 -8029 -1 0 -567
box -93 -248 93 248
use sg13g2_not_1  sg13g2_inv_1_0
timestamp 1752936403
transform 0 1 -9308 1 0 -326
box -48 -56 336 834
use sg13g2_not_1  sg13g2_inv_1_1
timestamp 1752936403
transform 0 1 -9308 1 0 -614
box -48 -56 336 834
<< labels >>
flabel metal2 -7917 -493 -7836 -412 0 FreeSans 320 0 0 0 G
port 10 nsew
flabel metal2 -7917 -279 -7836 -198 0 FreeSans 320 0 0 0 T
port 11 nsew
flabel metal1 -8375 -106 -8221 -10 0 FreeSans 320 0 0 0 VSS
port 12 nsew
flabel metal1 -8499 -106 -8432 -10 0 FreeSans 320 0 0 0 VDD
port 13 nsew
flabel metal2 -9524 -618 -9389 -537 0 FreeSans 320 0 0 0 EN
port 17 nsew
<< end >>
