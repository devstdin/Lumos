magic
tech ihp-sg13g2
timestamp 1757240632
<< error_p >>
rect -743 5990 -738 5995
rect 738 5990 743 5995
rect -748 5985 -743 5990
rect 743 5985 748 5990
rect -748 5974 -743 5979
rect 743 5974 748 5979
rect -743 5969 -738 5974
rect 738 5969 743 5974
rect -777 5953 -772 5958
rect -766 5953 -761 5958
rect 761 5953 766 5958
rect 772 5953 777 5958
rect -782 5948 -777 5953
rect -761 5948 -756 5953
rect 756 5948 761 5953
rect 777 5948 782 5953
rect -782 4967 -777 4972
rect -761 4967 -756 4972
rect 756 4967 761 4972
rect 777 4967 782 4972
rect -777 4962 -772 4967
rect -766 4962 -761 4967
rect 761 4962 766 4967
rect 772 4962 777 4967
rect -743 4946 -738 4951
rect 738 4946 743 4951
rect -748 4941 -743 4946
rect 743 4941 748 4946
rect -748 4930 -743 4935
rect 743 4930 748 4935
rect -743 4925 -738 4930
rect 738 4925 743 4930
rect -743 4898 -738 4903
rect 738 4898 743 4903
rect -748 4893 -743 4898
rect 743 4893 748 4898
rect -748 4882 -743 4887
rect 743 4882 748 4887
rect -743 4877 -738 4882
rect 738 4877 743 4882
rect -777 4861 -772 4866
rect -766 4861 -761 4866
rect 761 4861 766 4866
rect 772 4861 777 4866
rect -782 4856 -777 4861
rect -761 4856 -756 4861
rect 756 4856 761 4861
rect 777 4856 782 4861
rect -782 3875 -777 3880
rect -761 3875 -756 3880
rect 756 3875 761 3880
rect 777 3875 782 3880
rect -777 3870 -772 3875
rect -766 3870 -761 3875
rect 761 3870 766 3875
rect 772 3870 777 3875
rect -743 3854 -738 3859
rect 738 3854 743 3859
rect -748 3849 -743 3854
rect 743 3849 748 3854
rect -748 3838 -743 3843
rect 743 3838 748 3843
rect -743 3833 -738 3838
rect 738 3833 743 3838
rect -743 3806 -738 3811
rect 738 3806 743 3811
rect -748 3801 -743 3806
rect 743 3801 748 3806
rect -748 3790 -743 3795
rect 743 3790 748 3795
rect -743 3785 -738 3790
rect 738 3785 743 3790
rect -777 3769 -772 3774
rect -766 3769 -761 3774
rect 761 3769 766 3774
rect 772 3769 777 3774
rect -782 3764 -777 3769
rect -761 3764 -756 3769
rect 756 3764 761 3769
rect 777 3764 782 3769
rect -782 2783 -777 2788
rect -761 2783 -756 2788
rect 756 2783 761 2788
rect 777 2783 782 2788
rect -777 2778 -772 2783
rect -766 2778 -761 2783
rect 761 2778 766 2783
rect 772 2778 777 2783
rect -743 2762 -738 2767
rect 738 2762 743 2767
rect -748 2757 -743 2762
rect 743 2757 748 2762
rect -748 2746 -743 2751
rect 743 2746 748 2751
rect -743 2741 -738 2746
rect 738 2741 743 2746
rect -743 2714 -738 2719
rect 738 2714 743 2719
rect -748 2709 -743 2714
rect 743 2709 748 2714
rect -748 2698 -743 2703
rect 743 2698 748 2703
rect -743 2693 -738 2698
rect 738 2693 743 2698
rect -777 2677 -772 2682
rect -766 2677 -761 2682
rect 761 2677 766 2682
rect 772 2677 777 2682
rect -782 2672 -777 2677
rect -761 2672 -756 2677
rect 756 2672 761 2677
rect 777 2672 782 2677
rect -782 1691 -777 1696
rect -761 1691 -756 1696
rect 756 1691 761 1696
rect 777 1691 782 1696
rect -777 1686 -772 1691
rect -766 1686 -761 1691
rect 761 1686 766 1691
rect 772 1686 777 1691
rect -743 1670 -738 1675
rect 738 1670 743 1675
rect -748 1665 -743 1670
rect 743 1665 748 1670
rect -748 1654 -743 1659
rect 743 1654 748 1659
rect -743 1649 -738 1654
rect 738 1649 743 1654
rect -743 1622 -738 1627
rect 738 1622 743 1627
rect -748 1617 -743 1622
rect 743 1617 748 1622
rect -748 1606 -743 1611
rect 743 1606 748 1611
rect -743 1601 -738 1606
rect 738 1601 743 1606
rect -777 1585 -772 1590
rect -766 1585 -761 1590
rect 761 1585 766 1590
rect 772 1585 777 1590
rect -782 1580 -777 1585
rect -761 1580 -756 1585
rect 756 1580 761 1585
rect 777 1580 782 1585
rect -782 599 -777 604
rect -761 599 -756 604
rect 756 599 761 604
rect 777 599 782 604
rect -777 594 -772 599
rect -766 594 -761 599
rect 761 594 766 599
rect 772 594 777 599
rect -743 578 -738 583
rect 738 578 743 583
rect -748 573 -743 578
rect 743 573 748 578
rect -748 562 -743 567
rect 743 562 748 567
rect -743 557 -738 562
rect 738 557 743 562
rect -743 530 -738 535
rect 738 530 743 535
rect -748 525 -743 530
rect 743 525 748 530
rect -748 514 -743 519
rect 743 514 748 519
rect -743 509 -738 514
rect 738 509 743 514
rect -777 493 -772 498
rect -766 493 -761 498
rect 761 493 766 498
rect 772 493 777 498
rect -782 488 -777 493
rect -761 488 -756 493
rect 756 488 761 493
rect 777 488 782 493
rect -782 -493 -777 -488
rect -761 -493 -756 -488
rect 756 -493 761 -488
rect 777 -493 782 -488
rect -777 -498 -772 -493
rect -766 -498 -761 -493
rect 761 -498 766 -493
rect 772 -498 777 -493
rect -743 -514 -738 -509
rect 738 -514 743 -509
rect -748 -519 -743 -514
rect 743 -519 748 -514
rect -748 -530 -743 -525
rect 743 -530 748 -525
rect -743 -535 -738 -530
rect 738 -535 743 -530
<< nmos >>
rect -750 4960 750 5960
rect -750 3868 750 4868
rect -750 2776 750 3776
rect -750 1684 750 2684
rect -750 592 750 1592
rect -750 -500 750 500
<< ndiff >>
rect -784 5953 -750 5960
rect -784 4967 -777 5953
rect -761 4967 -750 5953
rect -784 4960 -750 4967
rect 750 5953 784 5960
rect 750 4967 761 5953
rect 777 4967 784 5953
rect 750 4960 784 4967
rect -784 4861 -750 4868
rect -784 3875 -777 4861
rect -761 3875 -750 4861
rect -784 3868 -750 3875
rect 750 4861 784 4868
rect 750 3875 761 4861
rect 777 3875 784 4861
rect 750 3868 784 3875
rect -784 3769 -750 3776
rect -784 2783 -777 3769
rect -761 2783 -750 3769
rect -784 2776 -750 2783
rect 750 3769 784 3776
rect 750 2783 761 3769
rect 777 2783 784 3769
rect 750 2776 784 2783
rect -784 2677 -750 2684
rect -784 1691 -777 2677
rect -761 1691 -750 2677
rect -784 1684 -750 1691
rect 750 2677 784 2684
rect 750 1691 761 2677
rect 777 1691 784 2677
rect 750 1684 784 1691
rect -784 1585 -750 1592
rect -784 599 -777 1585
rect -761 599 -750 1585
rect -784 592 -750 599
rect 750 1585 784 1592
rect 750 599 761 1585
rect 777 599 784 1585
rect 750 592 784 599
rect -784 493 -750 500
rect -784 -493 -777 493
rect -761 -493 -750 493
rect -784 -500 -750 -493
rect 750 493 784 500
rect 750 -493 761 493
rect 777 -493 784 493
rect 750 -500 784 -493
<< ndiffc >>
rect -777 4967 -761 5953
rect 761 4967 777 5953
rect -777 3875 -761 4861
rect 761 3875 777 4861
rect -777 2783 -761 3769
rect 761 2783 777 3769
rect -777 1691 -761 2677
rect 761 1691 777 2677
rect -777 599 -761 1585
rect 761 599 777 1585
rect -777 -493 -761 493
rect 761 -493 777 493
<< psubdiff >>
rect -877 5990 -847 5997
rect -877 -572 -870 5990
rect -854 -572 -847 5990
rect 847 5990 877 5997
rect -877 -579 -847 -572
rect 847 -572 854 5990
rect 870 -572 877 5990
rect 847 -579 877 -572
rect -877 -586 877 -579
rect -877 -602 -840 -586
rect 840 -602 877 -586
rect -877 -609 877 -602
<< psubdiffcont >>
rect -870 -572 -854 5990
rect 854 -572 870 5990
rect -840 -602 840 -586
<< poly >>
rect -750 5990 750 5997
rect -750 5974 -743 5990
rect 743 5974 750 5990
rect -750 5960 750 5974
rect -750 4946 750 4960
rect -750 4930 -743 4946
rect 743 4930 750 4946
rect -750 4923 750 4930
rect -750 4898 750 4905
rect -750 4882 -743 4898
rect 743 4882 750 4898
rect -750 4868 750 4882
rect -750 3854 750 3868
rect -750 3838 -743 3854
rect 743 3838 750 3854
rect -750 3831 750 3838
rect -750 3806 750 3813
rect -750 3790 -743 3806
rect 743 3790 750 3806
rect -750 3776 750 3790
rect -750 2762 750 2776
rect -750 2746 -743 2762
rect 743 2746 750 2762
rect -750 2739 750 2746
rect -750 2714 750 2721
rect -750 2698 -743 2714
rect 743 2698 750 2714
rect -750 2684 750 2698
rect -750 1670 750 1684
rect -750 1654 -743 1670
rect 743 1654 750 1670
rect -750 1647 750 1654
rect -750 1622 750 1629
rect -750 1606 -743 1622
rect 743 1606 750 1622
rect -750 1592 750 1606
rect -750 578 750 592
rect -750 562 -743 578
rect 743 562 750 578
rect -750 555 750 562
rect -750 530 750 537
rect -750 514 -743 530
rect 743 514 750 530
rect -750 500 750 514
rect -750 -514 750 -500
rect -750 -530 -743 -514
rect 743 -530 750 -514
rect -750 -537 750 -530
<< polycont >>
rect -743 5974 743 5990
rect -743 4930 743 4946
rect -743 4882 743 4898
rect -743 3838 743 3854
rect -743 3790 743 3806
rect -743 2746 743 2762
rect -743 2698 743 2714
rect -743 1654 743 1670
rect -743 1606 743 1622
rect -743 562 743 578
rect -743 514 743 530
rect -743 -530 743 -514
<< metal1 >>
rect -875 5990 -849 5995
rect 849 5990 875 5995
rect -875 -572 -870 5990
rect -854 -572 -849 5990
rect -875 -581 -849 -572
rect 849 -572 854 5990
rect 870 -572 875 5990
rect 849 -581 875 -572
rect -875 -586 875 -581
rect -875 -602 -840 -586
rect 840 -602 875 -586
rect -875 -607 875 -602
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 10 l 15 nf 1 nx 1 dx 0.21 ny 6 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 3 glc 1 grc 1 gtc 0 gbc 1
<< end >>
