magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< metal3 >>
rect -480 -20 -471 20
rect 471 -20 480 20
<< via3 >>
rect -471 -20 471 20
<< metal4 >>
rect -471 20 471 29
rect -471 -29 471 -20
<< properties >>
string GDS_END 6302
string GDS_FILE 6_final.gds
string GDS_START 5402
<< end >>
