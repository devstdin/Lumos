magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2124 18124 4104
<< nwell >>
rect -124 1788 16124 2104
rect -124 192 192 1788
rect 15808 192 16124 1788
rect -124 -124 16124 192
<< pwell >>
rect 334 1526 15666 1646
rect 334 454 454 1526
rect 3944 1244 4152 1526
rect 7642 454 8358 1526
rect 15546 454 15666 1526
rect 334 334 15666 454
<< hvnmos >>
rect 7762 550 7882 1430
rect 8118 550 8238 1430
<< hvndiff >>
rect 7668 1414 7762 1430
rect 7668 1382 7682 1414
rect 7714 1382 7762 1414
rect 7668 1346 7762 1382
rect 7668 1314 7682 1346
rect 7714 1314 7762 1346
rect 7668 1278 7762 1314
rect 7668 1246 7682 1278
rect 7714 1246 7762 1278
rect 7668 1210 7762 1246
rect 7668 1178 7682 1210
rect 7714 1178 7762 1210
rect 7668 1142 7762 1178
rect 7668 1110 7682 1142
rect 7714 1110 7762 1142
rect 7668 1074 7762 1110
rect 7668 1042 7682 1074
rect 7714 1042 7762 1074
rect 7668 1006 7762 1042
rect 7668 974 7682 1006
rect 7714 974 7762 1006
rect 7668 938 7762 974
rect 7668 906 7682 938
rect 7714 906 7762 938
rect 7668 870 7762 906
rect 7668 838 7682 870
rect 7714 838 7762 870
rect 7668 802 7762 838
rect 7668 770 7682 802
rect 7714 770 7762 802
rect 7668 734 7762 770
rect 7668 702 7682 734
rect 7714 702 7762 734
rect 7668 666 7762 702
rect 7668 634 7682 666
rect 7714 634 7762 666
rect 7668 598 7762 634
rect 7668 566 7682 598
rect 7714 566 7762 598
rect 7668 550 7762 566
rect 7882 1414 8118 1430
rect 7882 1382 7984 1414
rect 8016 1382 8118 1414
rect 7882 1346 8118 1382
rect 7882 1314 7984 1346
rect 8016 1314 8118 1346
rect 7882 1278 8118 1314
rect 7882 1246 7984 1278
rect 8016 1246 8118 1278
rect 7882 1210 8118 1246
rect 7882 1178 7984 1210
rect 8016 1178 8118 1210
rect 7882 1142 8118 1178
rect 7882 1110 7984 1142
rect 8016 1110 8118 1142
rect 7882 1074 8118 1110
rect 7882 1042 7984 1074
rect 8016 1042 8118 1074
rect 7882 1006 8118 1042
rect 7882 974 7984 1006
rect 8016 974 8118 1006
rect 7882 938 8118 974
rect 7882 906 7984 938
rect 8016 906 8118 938
rect 7882 870 8118 906
rect 7882 838 7984 870
rect 8016 838 8118 870
rect 7882 802 8118 838
rect 7882 770 7984 802
rect 8016 770 8118 802
rect 7882 734 8118 770
rect 7882 702 7984 734
rect 8016 702 8118 734
rect 7882 666 8118 702
rect 7882 634 7984 666
rect 8016 634 8118 666
rect 7882 598 8118 634
rect 7882 566 7984 598
rect 8016 566 8118 598
rect 7882 550 8118 566
rect 8238 1414 8332 1430
rect 8238 1382 8286 1414
rect 8318 1382 8332 1414
rect 8238 1346 8332 1382
rect 8238 1314 8286 1346
rect 8318 1314 8332 1346
rect 8238 1278 8332 1314
rect 8238 1246 8286 1278
rect 8318 1246 8332 1278
rect 8238 1210 8332 1246
rect 8238 1178 8286 1210
rect 8318 1178 8332 1210
rect 8238 1142 8332 1178
rect 8238 1110 8286 1142
rect 8318 1110 8332 1142
rect 8238 1074 8332 1110
rect 8238 1042 8286 1074
rect 8318 1042 8332 1074
rect 8238 1006 8332 1042
rect 8238 974 8286 1006
rect 8318 974 8332 1006
rect 8238 938 8332 974
rect 8238 906 8286 938
rect 8318 906 8332 938
rect 8238 870 8332 906
rect 8238 838 8286 870
rect 8318 838 8332 870
rect 8238 802 8332 838
rect 8238 770 8286 802
rect 8318 770 8332 802
rect 8238 734 8332 770
rect 8238 702 8286 734
rect 8318 702 8332 734
rect 8238 666 8332 702
rect 8238 634 8286 666
rect 8318 634 8332 666
rect 8238 598 8332 634
rect 8238 566 8286 598
rect 8318 566 8332 598
rect 8238 550 8332 566
<< hvndiffc >>
rect 7682 1382 7714 1414
rect 7682 1314 7714 1346
rect 7682 1246 7714 1278
rect 7682 1178 7714 1210
rect 7682 1110 7714 1142
rect 7682 1042 7714 1074
rect 7682 974 7714 1006
rect 7682 906 7714 938
rect 7682 838 7714 870
rect 7682 770 7714 802
rect 7682 702 7714 734
rect 7682 634 7714 666
rect 7682 566 7714 598
rect 7984 1382 8016 1414
rect 7984 1314 8016 1346
rect 7984 1246 8016 1278
rect 7984 1178 8016 1210
rect 7984 1110 8016 1142
rect 7984 1042 8016 1074
rect 7984 974 8016 1006
rect 7984 906 8016 938
rect 7984 838 8016 870
rect 7984 770 8016 802
rect 7984 702 8016 734
rect 7984 634 8016 666
rect 7984 566 8016 598
rect 8286 1382 8318 1414
rect 8286 1314 8318 1346
rect 8286 1246 8318 1278
rect 8286 1178 8318 1210
rect 8286 1110 8318 1142
rect 8286 1042 8318 1074
rect 8286 974 8318 1006
rect 8286 906 8318 938
rect 8286 838 8318 870
rect 8286 770 8318 802
rect 8286 702 8318 734
rect 8286 634 8318 666
rect 8286 566 8318 598
<< psubdiff >>
rect 360 1602 15640 1620
rect 360 1570 402 1602
rect 434 1570 470 1602
rect 502 1570 538 1602
rect 570 1570 606 1602
rect 638 1570 674 1602
rect 706 1570 742 1602
rect 774 1570 810 1602
rect 842 1570 878 1602
rect 910 1570 946 1602
rect 978 1570 1014 1602
rect 1046 1570 1082 1602
rect 1114 1570 1150 1602
rect 1182 1570 1218 1602
rect 1250 1570 1286 1602
rect 1318 1570 1354 1602
rect 1386 1570 1422 1602
rect 1454 1570 1490 1602
rect 1522 1570 1558 1602
rect 1590 1570 1626 1602
rect 1658 1570 1694 1602
rect 1726 1570 1762 1602
rect 1794 1570 1830 1602
rect 1862 1570 1898 1602
rect 1930 1570 1966 1602
rect 1998 1570 2034 1602
rect 2066 1570 2102 1602
rect 2134 1570 2170 1602
rect 2202 1570 2238 1602
rect 2270 1570 2306 1602
rect 2338 1570 2374 1602
rect 2406 1570 2442 1602
rect 2474 1570 2510 1602
rect 2542 1570 2578 1602
rect 2610 1570 2646 1602
rect 2678 1570 2714 1602
rect 2746 1570 2782 1602
rect 2814 1570 2850 1602
rect 2882 1570 2918 1602
rect 2950 1570 2986 1602
rect 3018 1570 3054 1602
rect 3086 1570 3122 1602
rect 3154 1570 3190 1602
rect 3222 1570 3258 1602
rect 3290 1570 3326 1602
rect 3358 1570 3394 1602
rect 3426 1570 3462 1602
rect 3494 1570 3530 1602
rect 3562 1570 3598 1602
rect 3630 1570 3666 1602
rect 3698 1570 3734 1602
rect 3766 1570 3802 1602
rect 3834 1570 3870 1602
rect 3902 1570 3938 1602
rect 3970 1570 4006 1602
rect 4038 1570 4074 1602
rect 4106 1570 4142 1602
rect 4174 1570 4210 1602
rect 4242 1570 4278 1602
rect 4310 1570 4346 1602
rect 4378 1570 4414 1602
rect 4446 1570 4482 1602
rect 4514 1570 4550 1602
rect 4582 1570 4618 1602
rect 4650 1570 4686 1602
rect 4718 1570 4754 1602
rect 4786 1570 4822 1602
rect 4854 1570 4890 1602
rect 4922 1570 4958 1602
rect 4990 1570 5026 1602
rect 5058 1570 5094 1602
rect 5126 1570 5162 1602
rect 5194 1570 5230 1602
rect 5262 1570 5298 1602
rect 5330 1570 5366 1602
rect 5398 1570 5434 1602
rect 5466 1570 5502 1602
rect 5534 1570 5570 1602
rect 5602 1570 5638 1602
rect 5670 1570 5706 1602
rect 5738 1570 5774 1602
rect 5806 1570 5842 1602
rect 5874 1570 5910 1602
rect 5942 1570 5978 1602
rect 6010 1570 6046 1602
rect 6078 1570 6114 1602
rect 6146 1570 6182 1602
rect 6214 1570 6250 1602
rect 6282 1570 6318 1602
rect 6350 1570 6386 1602
rect 6418 1570 6454 1602
rect 6486 1570 6522 1602
rect 6554 1570 6590 1602
rect 6622 1570 6658 1602
rect 6690 1570 6726 1602
rect 6758 1570 6794 1602
rect 6826 1570 6862 1602
rect 6894 1570 6930 1602
rect 6962 1570 6998 1602
rect 7030 1570 7066 1602
rect 7098 1570 7134 1602
rect 7166 1570 7202 1602
rect 7234 1570 7270 1602
rect 7302 1570 7338 1602
rect 7370 1570 7406 1602
rect 7438 1570 7474 1602
rect 7506 1570 7542 1602
rect 7574 1570 7610 1602
rect 7642 1570 7678 1602
rect 7710 1570 7746 1602
rect 7778 1570 7814 1602
rect 7846 1570 7882 1602
rect 7914 1570 7950 1602
rect 7982 1570 8018 1602
rect 8050 1570 8086 1602
rect 8118 1570 8154 1602
rect 8186 1570 8222 1602
rect 8254 1570 8290 1602
rect 8322 1570 8358 1602
rect 8390 1570 8426 1602
rect 8458 1570 8494 1602
rect 8526 1570 8562 1602
rect 8594 1570 8630 1602
rect 8662 1570 8698 1602
rect 8730 1570 8766 1602
rect 8798 1570 8834 1602
rect 8866 1570 8902 1602
rect 8934 1570 8970 1602
rect 9002 1570 9038 1602
rect 9070 1570 9106 1602
rect 9138 1570 9174 1602
rect 9206 1570 9242 1602
rect 9274 1570 9310 1602
rect 9342 1570 9378 1602
rect 9410 1570 9446 1602
rect 9478 1570 9514 1602
rect 9546 1570 9582 1602
rect 9614 1570 9650 1602
rect 9682 1570 9718 1602
rect 9750 1570 9786 1602
rect 9818 1570 9854 1602
rect 9886 1570 9922 1602
rect 9954 1570 9990 1602
rect 10022 1570 10058 1602
rect 10090 1570 10126 1602
rect 10158 1570 10194 1602
rect 10226 1570 10262 1602
rect 10294 1570 10330 1602
rect 10362 1570 10398 1602
rect 10430 1570 10466 1602
rect 10498 1570 10534 1602
rect 10566 1570 10602 1602
rect 10634 1570 10670 1602
rect 10702 1570 10738 1602
rect 10770 1570 10806 1602
rect 10838 1570 10874 1602
rect 10906 1570 10942 1602
rect 10974 1570 11010 1602
rect 11042 1570 11078 1602
rect 11110 1570 11146 1602
rect 11178 1570 11214 1602
rect 11246 1570 11282 1602
rect 11314 1570 11350 1602
rect 11382 1570 11418 1602
rect 11450 1570 11486 1602
rect 11518 1570 11554 1602
rect 11586 1570 11622 1602
rect 11654 1570 11690 1602
rect 11722 1570 11758 1602
rect 11790 1570 11826 1602
rect 11858 1570 11894 1602
rect 11926 1570 11962 1602
rect 11994 1570 12030 1602
rect 12062 1570 12098 1602
rect 12130 1570 12166 1602
rect 12198 1570 12234 1602
rect 12266 1570 12302 1602
rect 12334 1570 12370 1602
rect 12402 1570 12438 1602
rect 12470 1570 12506 1602
rect 12538 1570 12574 1602
rect 12606 1570 12642 1602
rect 12674 1570 12710 1602
rect 12742 1570 12778 1602
rect 12810 1570 12846 1602
rect 12878 1570 12914 1602
rect 12946 1570 12982 1602
rect 13014 1570 13050 1602
rect 13082 1570 13118 1602
rect 13150 1570 13186 1602
rect 13218 1570 13254 1602
rect 13286 1570 13322 1602
rect 13354 1570 13390 1602
rect 13422 1570 13458 1602
rect 13490 1570 13526 1602
rect 13558 1570 13594 1602
rect 13626 1570 13662 1602
rect 13694 1570 13730 1602
rect 13762 1570 13798 1602
rect 13830 1570 13866 1602
rect 13898 1570 13934 1602
rect 13966 1570 14002 1602
rect 14034 1570 14070 1602
rect 14102 1570 14138 1602
rect 14170 1570 14206 1602
rect 14238 1570 14274 1602
rect 14306 1570 14342 1602
rect 14374 1570 14410 1602
rect 14442 1570 14478 1602
rect 14510 1570 14546 1602
rect 14578 1570 14614 1602
rect 14646 1570 14682 1602
rect 14714 1570 14750 1602
rect 14782 1570 14818 1602
rect 14850 1570 14886 1602
rect 14918 1570 14954 1602
rect 14986 1570 15022 1602
rect 15054 1570 15090 1602
rect 15122 1570 15158 1602
rect 15190 1570 15226 1602
rect 15258 1570 15294 1602
rect 15326 1570 15362 1602
rect 15394 1570 15430 1602
rect 15462 1570 15498 1602
rect 15530 1570 15566 1602
rect 15598 1570 15640 1602
rect 360 1552 15640 1570
rect 360 1516 428 1552
rect 360 1484 378 1516
rect 410 1484 428 1516
rect 15572 1516 15640 1552
rect 360 1448 428 1484
rect 360 1416 378 1448
rect 410 1416 428 1448
rect 15572 1484 15590 1516
rect 15622 1484 15640 1516
rect 15572 1448 15640 1484
rect 360 1380 428 1416
rect 360 1348 378 1380
rect 410 1348 428 1380
rect 360 1312 428 1348
rect 360 1280 378 1312
rect 410 1280 428 1312
rect 360 1244 428 1280
rect 360 1212 378 1244
rect 410 1212 428 1244
rect 360 1176 428 1212
rect 360 1144 378 1176
rect 410 1144 428 1176
rect 360 1108 428 1144
rect 360 1076 378 1108
rect 410 1076 428 1108
rect 360 1040 428 1076
rect 360 1008 378 1040
rect 410 1008 428 1040
rect 360 972 428 1008
rect 360 940 378 972
rect 410 940 428 972
rect 360 904 428 940
rect 360 872 378 904
rect 410 872 428 904
rect 360 836 428 872
rect 360 804 378 836
rect 410 804 428 836
rect 360 768 428 804
rect 360 736 378 768
rect 410 736 428 768
rect 360 700 428 736
rect 360 668 378 700
rect 410 668 428 700
rect 360 632 428 668
rect 360 600 378 632
rect 410 600 428 632
rect 360 564 428 600
rect 360 532 378 564
rect 410 532 428 564
rect 15572 1416 15590 1448
rect 15622 1416 15640 1448
rect 15572 1380 15640 1416
rect 15572 1348 15590 1380
rect 15622 1348 15640 1380
rect 15572 1312 15640 1348
rect 15572 1280 15590 1312
rect 15622 1280 15640 1312
rect 15572 1244 15640 1280
rect 15572 1212 15590 1244
rect 15622 1212 15640 1244
rect 15572 1176 15640 1212
rect 15572 1144 15590 1176
rect 15622 1144 15640 1176
rect 15572 1108 15640 1144
rect 15572 1076 15590 1108
rect 15622 1076 15640 1108
rect 15572 1040 15640 1076
rect 15572 1008 15590 1040
rect 15622 1008 15640 1040
rect 15572 972 15640 1008
rect 15572 940 15590 972
rect 15622 940 15640 972
rect 15572 904 15640 940
rect 15572 872 15590 904
rect 15622 872 15640 904
rect 15572 836 15640 872
rect 15572 804 15590 836
rect 15622 804 15640 836
rect 15572 768 15640 804
rect 15572 736 15590 768
rect 15622 736 15640 768
rect 15572 700 15640 736
rect 15572 668 15590 700
rect 15622 668 15640 700
rect 15572 632 15640 668
rect 15572 600 15590 632
rect 15622 600 15640 632
rect 15572 564 15640 600
rect 360 496 428 532
rect 360 464 378 496
rect 410 464 428 496
rect 15572 532 15590 564
rect 15622 532 15640 564
rect 15572 496 15640 532
rect 360 428 428 464
rect 15572 464 15590 496
rect 15622 464 15640 496
rect 15572 428 15640 464
rect 360 410 15640 428
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 360 15640 378
<< nsubdiff >>
rect 0 1962 16000 1980
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 15932 360 16000 396
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< psubdiffcont >>
rect 402 1570 434 1602
rect 470 1570 502 1602
rect 538 1570 570 1602
rect 606 1570 638 1602
rect 674 1570 706 1602
rect 742 1570 774 1602
rect 810 1570 842 1602
rect 878 1570 910 1602
rect 946 1570 978 1602
rect 1014 1570 1046 1602
rect 1082 1570 1114 1602
rect 1150 1570 1182 1602
rect 1218 1570 1250 1602
rect 1286 1570 1318 1602
rect 1354 1570 1386 1602
rect 1422 1570 1454 1602
rect 1490 1570 1522 1602
rect 1558 1570 1590 1602
rect 1626 1570 1658 1602
rect 1694 1570 1726 1602
rect 1762 1570 1794 1602
rect 1830 1570 1862 1602
rect 1898 1570 1930 1602
rect 1966 1570 1998 1602
rect 2034 1570 2066 1602
rect 2102 1570 2134 1602
rect 2170 1570 2202 1602
rect 2238 1570 2270 1602
rect 2306 1570 2338 1602
rect 2374 1570 2406 1602
rect 2442 1570 2474 1602
rect 2510 1570 2542 1602
rect 2578 1570 2610 1602
rect 2646 1570 2678 1602
rect 2714 1570 2746 1602
rect 2782 1570 2814 1602
rect 2850 1570 2882 1602
rect 2918 1570 2950 1602
rect 2986 1570 3018 1602
rect 3054 1570 3086 1602
rect 3122 1570 3154 1602
rect 3190 1570 3222 1602
rect 3258 1570 3290 1602
rect 3326 1570 3358 1602
rect 3394 1570 3426 1602
rect 3462 1570 3494 1602
rect 3530 1570 3562 1602
rect 3598 1570 3630 1602
rect 3666 1570 3698 1602
rect 3734 1570 3766 1602
rect 3802 1570 3834 1602
rect 3870 1570 3902 1602
rect 3938 1570 3970 1602
rect 4006 1570 4038 1602
rect 4074 1570 4106 1602
rect 4142 1570 4174 1602
rect 4210 1570 4242 1602
rect 4278 1570 4310 1602
rect 4346 1570 4378 1602
rect 4414 1570 4446 1602
rect 4482 1570 4514 1602
rect 4550 1570 4582 1602
rect 4618 1570 4650 1602
rect 4686 1570 4718 1602
rect 4754 1570 4786 1602
rect 4822 1570 4854 1602
rect 4890 1570 4922 1602
rect 4958 1570 4990 1602
rect 5026 1570 5058 1602
rect 5094 1570 5126 1602
rect 5162 1570 5194 1602
rect 5230 1570 5262 1602
rect 5298 1570 5330 1602
rect 5366 1570 5398 1602
rect 5434 1570 5466 1602
rect 5502 1570 5534 1602
rect 5570 1570 5602 1602
rect 5638 1570 5670 1602
rect 5706 1570 5738 1602
rect 5774 1570 5806 1602
rect 5842 1570 5874 1602
rect 5910 1570 5942 1602
rect 5978 1570 6010 1602
rect 6046 1570 6078 1602
rect 6114 1570 6146 1602
rect 6182 1570 6214 1602
rect 6250 1570 6282 1602
rect 6318 1570 6350 1602
rect 6386 1570 6418 1602
rect 6454 1570 6486 1602
rect 6522 1570 6554 1602
rect 6590 1570 6622 1602
rect 6658 1570 6690 1602
rect 6726 1570 6758 1602
rect 6794 1570 6826 1602
rect 6862 1570 6894 1602
rect 6930 1570 6962 1602
rect 6998 1570 7030 1602
rect 7066 1570 7098 1602
rect 7134 1570 7166 1602
rect 7202 1570 7234 1602
rect 7270 1570 7302 1602
rect 7338 1570 7370 1602
rect 7406 1570 7438 1602
rect 7474 1570 7506 1602
rect 7542 1570 7574 1602
rect 7610 1570 7642 1602
rect 7678 1570 7710 1602
rect 7746 1570 7778 1602
rect 7814 1570 7846 1602
rect 7882 1570 7914 1602
rect 7950 1570 7982 1602
rect 8018 1570 8050 1602
rect 8086 1570 8118 1602
rect 8154 1570 8186 1602
rect 8222 1570 8254 1602
rect 8290 1570 8322 1602
rect 8358 1570 8390 1602
rect 8426 1570 8458 1602
rect 8494 1570 8526 1602
rect 8562 1570 8594 1602
rect 8630 1570 8662 1602
rect 8698 1570 8730 1602
rect 8766 1570 8798 1602
rect 8834 1570 8866 1602
rect 8902 1570 8934 1602
rect 8970 1570 9002 1602
rect 9038 1570 9070 1602
rect 9106 1570 9138 1602
rect 9174 1570 9206 1602
rect 9242 1570 9274 1602
rect 9310 1570 9342 1602
rect 9378 1570 9410 1602
rect 9446 1570 9478 1602
rect 9514 1570 9546 1602
rect 9582 1570 9614 1602
rect 9650 1570 9682 1602
rect 9718 1570 9750 1602
rect 9786 1570 9818 1602
rect 9854 1570 9886 1602
rect 9922 1570 9954 1602
rect 9990 1570 10022 1602
rect 10058 1570 10090 1602
rect 10126 1570 10158 1602
rect 10194 1570 10226 1602
rect 10262 1570 10294 1602
rect 10330 1570 10362 1602
rect 10398 1570 10430 1602
rect 10466 1570 10498 1602
rect 10534 1570 10566 1602
rect 10602 1570 10634 1602
rect 10670 1570 10702 1602
rect 10738 1570 10770 1602
rect 10806 1570 10838 1602
rect 10874 1570 10906 1602
rect 10942 1570 10974 1602
rect 11010 1570 11042 1602
rect 11078 1570 11110 1602
rect 11146 1570 11178 1602
rect 11214 1570 11246 1602
rect 11282 1570 11314 1602
rect 11350 1570 11382 1602
rect 11418 1570 11450 1602
rect 11486 1570 11518 1602
rect 11554 1570 11586 1602
rect 11622 1570 11654 1602
rect 11690 1570 11722 1602
rect 11758 1570 11790 1602
rect 11826 1570 11858 1602
rect 11894 1570 11926 1602
rect 11962 1570 11994 1602
rect 12030 1570 12062 1602
rect 12098 1570 12130 1602
rect 12166 1570 12198 1602
rect 12234 1570 12266 1602
rect 12302 1570 12334 1602
rect 12370 1570 12402 1602
rect 12438 1570 12470 1602
rect 12506 1570 12538 1602
rect 12574 1570 12606 1602
rect 12642 1570 12674 1602
rect 12710 1570 12742 1602
rect 12778 1570 12810 1602
rect 12846 1570 12878 1602
rect 12914 1570 12946 1602
rect 12982 1570 13014 1602
rect 13050 1570 13082 1602
rect 13118 1570 13150 1602
rect 13186 1570 13218 1602
rect 13254 1570 13286 1602
rect 13322 1570 13354 1602
rect 13390 1570 13422 1602
rect 13458 1570 13490 1602
rect 13526 1570 13558 1602
rect 13594 1570 13626 1602
rect 13662 1570 13694 1602
rect 13730 1570 13762 1602
rect 13798 1570 13830 1602
rect 13866 1570 13898 1602
rect 13934 1570 13966 1602
rect 14002 1570 14034 1602
rect 14070 1570 14102 1602
rect 14138 1570 14170 1602
rect 14206 1570 14238 1602
rect 14274 1570 14306 1602
rect 14342 1570 14374 1602
rect 14410 1570 14442 1602
rect 14478 1570 14510 1602
rect 14546 1570 14578 1602
rect 14614 1570 14646 1602
rect 14682 1570 14714 1602
rect 14750 1570 14782 1602
rect 14818 1570 14850 1602
rect 14886 1570 14918 1602
rect 14954 1570 14986 1602
rect 15022 1570 15054 1602
rect 15090 1570 15122 1602
rect 15158 1570 15190 1602
rect 15226 1570 15258 1602
rect 15294 1570 15326 1602
rect 15362 1570 15394 1602
rect 15430 1570 15462 1602
rect 15498 1570 15530 1602
rect 15566 1570 15598 1602
rect 378 1484 410 1516
rect 378 1416 410 1448
rect 15590 1484 15622 1516
rect 378 1348 410 1380
rect 378 1280 410 1312
rect 378 1212 410 1244
rect 378 1144 410 1176
rect 378 1076 410 1108
rect 378 1008 410 1040
rect 378 940 410 972
rect 378 872 410 904
rect 378 804 410 836
rect 378 736 410 768
rect 378 668 410 700
rect 378 600 410 632
rect 378 532 410 564
rect 15590 1416 15622 1448
rect 15590 1348 15622 1380
rect 15590 1280 15622 1312
rect 15590 1212 15622 1244
rect 15590 1144 15622 1176
rect 15590 1076 15622 1108
rect 15590 1008 15622 1040
rect 15590 940 15622 972
rect 15590 872 15622 904
rect 15590 804 15622 836
rect 15590 736 15622 768
rect 15590 668 15622 700
rect 15590 600 15622 632
rect 378 464 410 496
rect 15590 532 15622 564
rect 15590 464 15622 496
rect 402 378 434 410
rect 470 378 502 410
rect 538 378 570 410
rect 606 378 638 410
rect 674 378 706 410
rect 742 378 774 410
rect 810 378 842 410
rect 878 378 910 410
rect 946 378 978 410
rect 1014 378 1046 410
rect 1082 378 1114 410
rect 1150 378 1182 410
rect 1218 378 1250 410
rect 1286 378 1318 410
rect 1354 378 1386 410
rect 1422 378 1454 410
rect 1490 378 1522 410
rect 1558 378 1590 410
rect 1626 378 1658 410
rect 1694 378 1726 410
rect 1762 378 1794 410
rect 1830 378 1862 410
rect 1898 378 1930 410
rect 1966 378 1998 410
rect 2034 378 2066 410
rect 2102 378 2134 410
rect 2170 378 2202 410
rect 2238 378 2270 410
rect 2306 378 2338 410
rect 2374 378 2406 410
rect 2442 378 2474 410
rect 2510 378 2542 410
rect 2578 378 2610 410
rect 2646 378 2678 410
rect 2714 378 2746 410
rect 2782 378 2814 410
rect 2850 378 2882 410
rect 2918 378 2950 410
rect 2986 378 3018 410
rect 3054 378 3086 410
rect 3122 378 3154 410
rect 3190 378 3222 410
rect 3258 378 3290 410
rect 3326 378 3358 410
rect 3394 378 3426 410
rect 3462 378 3494 410
rect 3530 378 3562 410
rect 3598 378 3630 410
rect 3666 378 3698 410
rect 3734 378 3766 410
rect 3802 378 3834 410
rect 3870 378 3902 410
rect 3938 378 3970 410
rect 4006 378 4038 410
rect 4074 378 4106 410
rect 4142 378 4174 410
rect 4210 378 4242 410
rect 4278 378 4310 410
rect 4346 378 4378 410
rect 4414 378 4446 410
rect 4482 378 4514 410
rect 4550 378 4582 410
rect 4618 378 4650 410
rect 4686 378 4718 410
rect 4754 378 4786 410
rect 4822 378 4854 410
rect 4890 378 4922 410
rect 4958 378 4990 410
rect 5026 378 5058 410
rect 5094 378 5126 410
rect 5162 378 5194 410
rect 5230 378 5262 410
rect 5298 378 5330 410
rect 5366 378 5398 410
rect 5434 378 5466 410
rect 5502 378 5534 410
rect 5570 378 5602 410
rect 5638 378 5670 410
rect 5706 378 5738 410
rect 5774 378 5806 410
rect 5842 378 5874 410
rect 5910 378 5942 410
rect 5978 378 6010 410
rect 6046 378 6078 410
rect 6114 378 6146 410
rect 6182 378 6214 410
rect 6250 378 6282 410
rect 6318 378 6350 410
rect 6386 378 6418 410
rect 6454 378 6486 410
rect 6522 378 6554 410
rect 6590 378 6622 410
rect 6658 378 6690 410
rect 6726 378 6758 410
rect 6794 378 6826 410
rect 6862 378 6894 410
rect 6930 378 6962 410
rect 6998 378 7030 410
rect 7066 378 7098 410
rect 7134 378 7166 410
rect 7202 378 7234 410
rect 7270 378 7302 410
rect 7338 378 7370 410
rect 7406 378 7438 410
rect 7474 378 7506 410
rect 7542 378 7574 410
rect 7610 378 7642 410
rect 7678 378 7710 410
rect 7746 378 7778 410
rect 7814 378 7846 410
rect 7882 378 7914 410
rect 7950 378 7982 410
rect 8018 378 8050 410
rect 8086 378 8118 410
rect 8154 378 8186 410
rect 8222 378 8254 410
rect 8290 378 8322 410
rect 8358 378 8390 410
rect 8426 378 8458 410
rect 8494 378 8526 410
rect 8562 378 8594 410
rect 8630 378 8662 410
rect 8698 378 8730 410
rect 8766 378 8798 410
rect 8834 378 8866 410
rect 8902 378 8934 410
rect 8970 378 9002 410
rect 9038 378 9070 410
rect 9106 378 9138 410
rect 9174 378 9206 410
rect 9242 378 9274 410
rect 9310 378 9342 410
rect 9378 378 9410 410
rect 9446 378 9478 410
rect 9514 378 9546 410
rect 9582 378 9614 410
rect 9650 378 9682 410
rect 9718 378 9750 410
rect 9786 378 9818 410
rect 9854 378 9886 410
rect 9922 378 9954 410
rect 9990 378 10022 410
rect 10058 378 10090 410
rect 10126 378 10158 410
rect 10194 378 10226 410
rect 10262 378 10294 410
rect 10330 378 10362 410
rect 10398 378 10430 410
rect 10466 378 10498 410
rect 10534 378 10566 410
rect 10602 378 10634 410
rect 10670 378 10702 410
rect 10738 378 10770 410
rect 10806 378 10838 410
rect 10874 378 10906 410
rect 10942 378 10974 410
rect 11010 378 11042 410
rect 11078 378 11110 410
rect 11146 378 11178 410
rect 11214 378 11246 410
rect 11282 378 11314 410
rect 11350 378 11382 410
rect 11418 378 11450 410
rect 11486 378 11518 410
rect 11554 378 11586 410
rect 11622 378 11654 410
rect 11690 378 11722 410
rect 11758 378 11790 410
rect 11826 378 11858 410
rect 11894 378 11926 410
rect 11962 378 11994 410
rect 12030 378 12062 410
rect 12098 378 12130 410
rect 12166 378 12198 410
rect 12234 378 12266 410
rect 12302 378 12334 410
rect 12370 378 12402 410
rect 12438 378 12470 410
rect 12506 378 12538 410
rect 12574 378 12606 410
rect 12642 378 12674 410
rect 12710 378 12742 410
rect 12778 378 12810 410
rect 12846 378 12878 410
rect 12914 378 12946 410
rect 12982 378 13014 410
rect 13050 378 13082 410
rect 13118 378 13150 410
rect 13186 378 13218 410
rect 13254 378 13286 410
rect 13322 378 13354 410
rect 13390 378 13422 410
rect 13458 378 13490 410
rect 13526 378 13558 410
rect 13594 378 13626 410
rect 13662 378 13694 410
rect 13730 378 13762 410
rect 13798 378 13830 410
rect 13866 378 13898 410
rect 13934 378 13966 410
rect 14002 378 14034 410
rect 14070 378 14102 410
rect 14138 378 14170 410
rect 14206 378 14238 410
rect 14274 378 14306 410
rect 14342 378 14374 410
rect 14410 378 14442 410
rect 14478 378 14510 410
rect 14546 378 14578 410
rect 14614 378 14646 410
rect 14682 378 14714 410
rect 14750 378 14782 410
rect 14818 378 14850 410
rect 14886 378 14918 410
rect 14954 378 14986 410
rect 15022 378 15054 410
rect 15090 378 15122 410
rect 15158 378 15190 410
rect 15226 378 15258 410
rect 15294 378 15326 410
rect 15362 378 15394 410
rect 15430 378 15462 410
rect 15498 378 15530 410
rect 15566 378 15598 410
<< nsubdiffcont >>
rect 28 1930 60 1962
rect 96 1930 128 1962
rect 164 1930 196 1962
rect 232 1930 264 1962
rect 300 1930 332 1962
rect 368 1930 400 1962
rect 436 1930 468 1962
rect 504 1930 536 1962
rect 572 1930 604 1962
rect 640 1930 672 1962
rect 708 1930 740 1962
rect 776 1930 808 1962
rect 844 1930 876 1962
rect 912 1930 944 1962
rect 980 1930 1012 1962
rect 1048 1930 1080 1962
rect 1116 1930 1148 1962
rect 1184 1930 1216 1962
rect 1252 1930 1284 1962
rect 1320 1930 1352 1962
rect 1388 1930 1420 1962
rect 1456 1930 1488 1962
rect 1524 1930 1556 1962
rect 1592 1930 1624 1962
rect 1660 1930 1692 1962
rect 1728 1930 1760 1962
rect 1796 1930 1828 1962
rect 1864 1930 1896 1962
rect 1932 1930 1964 1962
rect 2000 1930 2032 1962
rect 2068 1930 2100 1962
rect 2136 1930 2168 1962
rect 2204 1930 2236 1962
rect 2272 1930 2304 1962
rect 2340 1930 2372 1962
rect 2408 1930 2440 1962
rect 2476 1930 2508 1962
rect 2544 1930 2576 1962
rect 2612 1930 2644 1962
rect 2680 1930 2712 1962
rect 2748 1930 2780 1962
rect 2816 1930 2848 1962
rect 2884 1930 2916 1962
rect 2952 1930 2984 1962
rect 3020 1930 3052 1962
rect 3088 1930 3120 1962
rect 3156 1930 3188 1962
rect 3224 1930 3256 1962
rect 3292 1930 3324 1962
rect 3360 1930 3392 1962
rect 3428 1930 3460 1962
rect 3496 1930 3528 1962
rect 3564 1930 3596 1962
rect 3632 1930 3664 1962
rect 3700 1930 3732 1962
rect 3768 1930 3800 1962
rect 3836 1930 3868 1962
rect 3904 1930 3936 1962
rect 3972 1930 4004 1962
rect 4040 1930 4072 1962
rect 4108 1930 4140 1962
rect 4176 1930 4208 1962
rect 4244 1930 4276 1962
rect 4312 1930 4344 1962
rect 4380 1930 4412 1962
rect 4448 1930 4480 1962
rect 4516 1930 4548 1962
rect 4584 1930 4616 1962
rect 4652 1930 4684 1962
rect 4720 1930 4752 1962
rect 4788 1930 4820 1962
rect 4856 1930 4888 1962
rect 4924 1930 4956 1962
rect 4992 1930 5024 1962
rect 5060 1930 5092 1962
rect 5128 1930 5160 1962
rect 5196 1930 5228 1962
rect 5264 1930 5296 1962
rect 5332 1930 5364 1962
rect 5400 1930 5432 1962
rect 5468 1930 5500 1962
rect 5536 1930 5568 1962
rect 5604 1930 5636 1962
rect 5672 1930 5704 1962
rect 5740 1930 5772 1962
rect 5808 1930 5840 1962
rect 5876 1930 5908 1962
rect 5944 1930 5976 1962
rect 6012 1930 6044 1962
rect 6080 1930 6112 1962
rect 6148 1930 6180 1962
rect 6216 1930 6248 1962
rect 6284 1930 6316 1962
rect 6352 1930 6384 1962
rect 6420 1930 6452 1962
rect 6488 1930 6520 1962
rect 6556 1930 6588 1962
rect 6624 1930 6656 1962
rect 6692 1930 6724 1962
rect 6760 1930 6792 1962
rect 6828 1930 6860 1962
rect 6896 1930 6928 1962
rect 6964 1930 6996 1962
rect 7032 1930 7064 1962
rect 7100 1930 7132 1962
rect 7168 1930 7200 1962
rect 7236 1930 7268 1962
rect 7304 1930 7336 1962
rect 7372 1930 7404 1962
rect 7440 1930 7472 1962
rect 7508 1930 7540 1962
rect 7576 1930 7608 1962
rect 7644 1930 7676 1962
rect 7712 1930 7744 1962
rect 7780 1930 7812 1962
rect 7848 1930 7880 1962
rect 7916 1930 7948 1962
rect 7984 1930 8016 1962
rect 8052 1930 8084 1962
rect 8120 1930 8152 1962
rect 8188 1930 8220 1962
rect 8256 1930 8288 1962
rect 8324 1930 8356 1962
rect 8392 1930 8424 1962
rect 8460 1930 8492 1962
rect 8528 1930 8560 1962
rect 8596 1930 8628 1962
rect 8664 1930 8696 1962
rect 8732 1930 8764 1962
rect 8800 1930 8832 1962
rect 8868 1930 8900 1962
rect 8936 1930 8968 1962
rect 9004 1930 9036 1962
rect 9072 1930 9104 1962
rect 9140 1930 9172 1962
rect 9208 1930 9240 1962
rect 9276 1930 9308 1962
rect 9344 1930 9376 1962
rect 9412 1930 9444 1962
rect 9480 1930 9512 1962
rect 9548 1930 9580 1962
rect 9616 1930 9648 1962
rect 9684 1930 9716 1962
rect 9752 1930 9784 1962
rect 9820 1930 9852 1962
rect 9888 1930 9920 1962
rect 9956 1930 9988 1962
rect 10024 1930 10056 1962
rect 10092 1930 10124 1962
rect 10160 1930 10192 1962
rect 10228 1930 10260 1962
rect 10296 1930 10328 1962
rect 10364 1930 10396 1962
rect 10432 1930 10464 1962
rect 10500 1930 10532 1962
rect 10568 1930 10600 1962
rect 10636 1930 10668 1962
rect 10704 1930 10736 1962
rect 10772 1930 10804 1962
rect 10840 1930 10872 1962
rect 10908 1930 10940 1962
rect 10976 1930 11008 1962
rect 11044 1930 11076 1962
rect 11112 1930 11144 1962
rect 11180 1930 11212 1962
rect 11248 1930 11280 1962
rect 11316 1930 11348 1962
rect 11384 1930 11416 1962
rect 11452 1930 11484 1962
rect 11520 1930 11552 1962
rect 11588 1930 11620 1962
rect 11656 1930 11688 1962
rect 11724 1930 11756 1962
rect 11792 1930 11824 1962
rect 11860 1930 11892 1962
rect 11928 1930 11960 1962
rect 11996 1930 12028 1962
rect 12064 1930 12096 1962
rect 12132 1930 12164 1962
rect 12200 1930 12232 1962
rect 12268 1930 12300 1962
rect 12336 1930 12368 1962
rect 12404 1930 12436 1962
rect 12472 1930 12504 1962
rect 12540 1930 12572 1962
rect 12608 1930 12640 1962
rect 12676 1930 12708 1962
rect 12744 1930 12776 1962
rect 12812 1930 12844 1962
rect 12880 1930 12912 1962
rect 12948 1930 12980 1962
rect 13016 1930 13048 1962
rect 13084 1930 13116 1962
rect 13152 1930 13184 1962
rect 13220 1930 13252 1962
rect 13288 1930 13320 1962
rect 13356 1930 13388 1962
rect 13424 1930 13456 1962
rect 13492 1930 13524 1962
rect 13560 1930 13592 1962
rect 13628 1930 13660 1962
rect 13696 1930 13728 1962
rect 13764 1930 13796 1962
rect 13832 1930 13864 1962
rect 13900 1930 13932 1962
rect 13968 1930 14000 1962
rect 14036 1930 14068 1962
rect 14104 1930 14136 1962
rect 14172 1930 14204 1962
rect 14240 1930 14272 1962
rect 14308 1930 14340 1962
rect 14376 1930 14408 1962
rect 14444 1930 14476 1962
rect 14512 1930 14544 1962
rect 14580 1930 14612 1962
rect 14648 1930 14680 1962
rect 14716 1930 14748 1962
rect 14784 1930 14816 1962
rect 14852 1930 14884 1962
rect 14920 1930 14952 1962
rect 14988 1930 15020 1962
rect 15056 1930 15088 1962
rect 15124 1930 15156 1962
rect 15192 1930 15224 1962
rect 15260 1930 15292 1962
rect 15328 1930 15360 1962
rect 15396 1930 15428 1962
rect 15464 1930 15496 1962
rect 15532 1930 15564 1962
rect 15600 1930 15632 1962
rect 15668 1930 15700 1962
rect 15736 1930 15768 1962
rect 15804 1930 15836 1962
rect 15872 1930 15904 1962
rect 15940 1930 15972 1962
rect 18 1824 50 1856
rect 18 1756 50 1788
rect 18 1688 50 1720
rect 18 1620 50 1652
rect 15950 1824 15982 1856
rect 15950 1756 15982 1788
rect 15950 1688 15982 1720
rect 15950 1620 15982 1652
rect 18 1552 50 1584
rect 18 1484 50 1516
rect 18 1416 50 1448
rect 18 1348 50 1380
rect 18 1280 50 1312
rect 18 1212 50 1244
rect 18 1144 50 1176
rect 18 1076 50 1108
rect 18 1008 50 1040
rect 18 940 50 972
rect 18 872 50 904
rect 18 804 50 836
rect 18 736 50 768
rect 18 668 50 700
rect 18 600 50 632
rect 18 532 50 564
rect 18 464 50 496
rect 18 396 50 428
rect 15950 1552 15982 1584
rect 15950 1484 15982 1516
rect 15950 1416 15982 1448
rect 15950 1348 15982 1380
rect 15950 1280 15982 1312
rect 15950 1212 15982 1244
rect 15950 1144 15982 1176
rect 15950 1076 15982 1108
rect 15950 1008 15982 1040
rect 15950 940 15982 972
rect 15950 872 15982 904
rect 15950 804 15982 836
rect 15950 736 15982 768
rect 15950 668 15982 700
rect 15950 600 15982 632
rect 15950 532 15982 564
rect 15950 464 15982 496
rect 15950 396 15982 428
rect 18 328 50 360
rect 18 260 50 292
rect 18 192 50 224
rect 18 124 50 156
rect 15950 328 15982 360
rect 15950 260 15982 292
rect 15950 192 15982 224
rect 15950 124 15982 156
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< poly >>
rect 7762 1490 7882 1504
rect 7762 1458 7806 1490
rect 7838 1458 7882 1490
rect 7762 1430 7882 1458
rect 8118 1490 8238 1504
rect 8118 1458 8162 1490
rect 8194 1458 8238 1490
rect 8118 1430 8238 1458
rect 7762 522 7882 550
rect 7762 490 7806 522
rect 7838 490 7882 522
rect 7762 476 7882 490
rect 8118 522 8238 550
rect 8118 490 8162 522
rect 8194 490 8238 522
rect 8118 476 8238 490
<< polycont >>
rect 7806 1458 7838 1490
rect 8162 1458 8194 1490
rect 7806 490 7838 522
rect 8162 490 8194 522
<< ndiode >>
rect 3970 1398 4126 1426
rect 3970 1366 3998 1398
rect 4030 1366 4066 1398
rect 4098 1366 4126 1398
rect 3970 1330 4126 1366
rect 3970 1298 3998 1330
rect 4030 1298 4066 1330
rect 4098 1298 4126 1330
rect 3970 1270 4126 1298
<< ndiodecont >>
rect 3998 1366 4030 1398
rect 4066 1366 4098 1398
rect 3998 1298 4030 1330
rect 4066 1298 4098 1330
<< metal1 >>
rect 0 1962 16000 1980
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 360 1606 15640 1620
rect 360 1602 7678 1606
rect 7718 1602 8282 1606
rect 8322 1602 15640 1606
rect 360 1570 402 1602
rect 434 1570 470 1602
rect 502 1570 538 1602
rect 570 1570 606 1602
rect 638 1570 674 1602
rect 706 1570 742 1602
rect 774 1570 810 1602
rect 842 1570 878 1602
rect 910 1570 946 1602
rect 978 1570 1014 1602
rect 1046 1570 1082 1602
rect 1114 1570 1150 1602
rect 1182 1570 1218 1602
rect 1250 1570 1286 1602
rect 1318 1570 1354 1602
rect 1386 1570 1422 1602
rect 1454 1570 1490 1602
rect 1522 1570 1558 1602
rect 1590 1570 1626 1602
rect 1658 1570 1694 1602
rect 1726 1570 1762 1602
rect 1794 1570 1830 1602
rect 1862 1570 1898 1602
rect 1930 1570 1966 1602
rect 1998 1570 2034 1602
rect 2066 1570 2102 1602
rect 2134 1570 2170 1602
rect 2202 1570 2238 1602
rect 2270 1570 2306 1602
rect 2338 1570 2374 1602
rect 2406 1570 2442 1602
rect 2474 1570 2510 1602
rect 2542 1570 2578 1602
rect 2610 1570 2646 1602
rect 2678 1570 2714 1602
rect 2746 1570 2782 1602
rect 2814 1570 2850 1602
rect 2882 1570 2918 1602
rect 2950 1570 2986 1602
rect 3018 1570 3054 1602
rect 3086 1570 3122 1602
rect 3154 1570 3190 1602
rect 3222 1570 3258 1602
rect 3290 1570 3326 1602
rect 3358 1570 3394 1602
rect 3426 1570 3462 1602
rect 3494 1570 3530 1602
rect 3562 1570 3598 1602
rect 3630 1570 3666 1602
rect 3698 1570 3734 1602
rect 3766 1570 3802 1602
rect 3834 1570 3870 1602
rect 3902 1570 3938 1602
rect 3970 1570 4006 1602
rect 4038 1570 4074 1602
rect 4106 1570 4142 1602
rect 4174 1570 4210 1602
rect 4242 1570 4278 1602
rect 4310 1570 4346 1602
rect 4378 1570 4414 1602
rect 4446 1570 4482 1602
rect 4514 1570 4550 1602
rect 4582 1570 4618 1602
rect 4650 1570 4686 1602
rect 4718 1570 4754 1602
rect 4786 1570 4822 1602
rect 4854 1570 4890 1602
rect 4922 1570 4958 1602
rect 4990 1570 5026 1602
rect 5058 1570 5094 1602
rect 5126 1570 5162 1602
rect 5194 1570 5230 1602
rect 5262 1570 5298 1602
rect 5330 1570 5366 1602
rect 5398 1570 5434 1602
rect 5466 1570 5502 1602
rect 5534 1570 5570 1602
rect 5602 1570 5638 1602
rect 5670 1570 5706 1602
rect 5738 1570 5774 1602
rect 5806 1570 5842 1602
rect 5874 1570 5910 1602
rect 5942 1570 5978 1602
rect 6010 1570 6046 1602
rect 6078 1570 6114 1602
rect 6146 1570 6182 1602
rect 6214 1570 6250 1602
rect 6282 1570 6318 1602
rect 6350 1570 6386 1602
rect 6418 1570 6454 1602
rect 6486 1570 6522 1602
rect 6554 1570 6590 1602
rect 6622 1570 6658 1602
rect 6690 1570 6726 1602
rect 6758 1570 6794 1602
rect 6826 1570 6862 1602
rect 6894 1570 6930 1602
rect 6962 1570 6998 1602
rect 7030 1570 7066 1602
rect 7098 1570 7134 1602
rect 7166 1570 7202 1602
rect 7234 1570 7270 1602
rect 7302 1570 7338 1602
rect 7370 1570 7406 1602
rect 7438 1570 7474 1602
rect 7506 1570 7542 1602
rect 7574 1570 7610 1602
rect 7642 1570 7678 1602
rect 7718 1570 7746 1602
rect 7778 1570 7814 1602
rect 7846 1570 7882 1602
rect 7914 1570 7950 1602
rect 7982 1570 8018 1602
rect 8050 1570 8086 1602
rect 8118 1570 8154 1602
rect 8186 1570 8222 1602
rect 8254 1570 8282 1602
rect 8322 1570 8358 1602
rect 8390 1570 8426 1602
rect 8458 1570 8494 1602
rect 8526 1570 8562 1602
rect 8594 1570 8630 1602
rect 8662 1570 8698 1602
rect 8730 1570 8766 1602
rect 8798 1570 8834 1602
rect 8866 1570 8902 1602
rect 8934 1570 8970 1602
rect 9002 1570 9038 1602
rect 9070 1570 9106 1602
rect 9138 1570 9174 1602
rect 9206 1570 9242 1602
rect 9274 1570 9310 1602
rect 9342 1570 9378 1602
rect 9410 1570 9446 1602
rect 9478 1570 9514 1602
rect 9546 1570 9582 1602
rect 9614 1570 9650 1602
rect 9682 1570 9718 1602
rect 9750 1570 9786 1602
rect 9818 1570 9854 1602
rect 9886 1570 9922 1602
rect 9954 1570 9990 1602
rect 10022 1570 10058 1602
rect 10090 1570 10126 1602
rect 10158 1570 10194 1602
rect 10226 1570 10262 1602
rect 10294 1570 10330 1602
rect 10362 1570 10398 1602
rect 10430 1570 10466 1602
rect 10498 1570 10534 1602
rect 10566 1570 10602 1602
rect 10634 1570 10670 1602
rect 10702 1570 10738 1602
rect 10770 1570 10806 1602
rect 10838 1570 10874 1602
rect 10906 1570 10942 1602
rect 10974 1570 11010 1602
rect 11042 1570 11078 1602
rect 11110 1570 11146 1602
rect 11178 1570 11214 1602
rect 11246 1570 11282 1602
rect 11314 1570 11350 1602
rect 11382 1570 11418 1602
rect 11450 1570 11486 1602
rect 11518 1570 11554 1602
rect 11586 1570 11622 1602
rect 11654 1570 11690 1602
rect 11722 1570 11758 1602
rect 11790 1570 11826 1602
rect 11858 1570 11894 1602
rect 11926 1570 11962 1602
rect 11994 1570 12030 1602
rect 12062 1570 12098 1602
rect 12130 1570 12166 1602
rect 12198 1570 12234 1602
rect 12266 1570 12302 1602
rect 12334 1570 12370 1602
rect 12402 1570 12438 1602
rect 12470 1570 12506 1602
rect 12538 1570 12574 1602
rect 12606 1570 12642 1602
rect 12674 1570 12710 1602
rect 12742 1570 12778 1602
rect 12810 1570 12846 1602
rect 12878 1570 12914 1602
rect 12946 1570 12982 1602
rect 13014 1570 13050 1602
rect 13082 1570 13118 1602
rect 13150 1570 13186 1602
rect 13218 1570 13254 1602
rect 13286 1570 13322 1602
rect 13354 1570 13390 1602
rect 13422 1570 13458 1602
rect 13490 1570 13526 1602
rect 13558 1570 13594 1602
rect 13626 1570 13662 1602
rect 13694 1570 13730 1602
rect 13762 1570 13798 1602
rect 13830 1570 13866 1602
rect 13898 1570 13934 1602
rect 13966 1570 14002 1602
rect 14034 1570 14070 1602
rect 14102 1570 14138 1602
rect 14170 1570 14206 1602
rect 14238 1570 14274 1602
rect 14306 1570 14342 1602
rect 14374 1570 14410 1602
rect 14442 1570 14478 1602
rect 14510 1570 14546 1602
rect 14578 1570 14614 1602
rect 14646 1570 14682 1602
rect 14714 1570 14750 1602
rect 14782 1570 14818 1602
rect 14850 1570 14886 1602
rect 14918 1570 14954 1602
rect 14986 1570 15022 1602
rect 15054 1570 15090 1602
rect 15122 1570 15158 1602
rect 15190 1570 15226 1602
rect 15258 1570 15294 1602
rect 15326 1570 15362 1602
rect 15394 1570 15430 1602
rect 15462 1570 15498 1602
rect 15530 1570 15566 1602
rect 15598 1570 15640 1602
rect 360 1566 7678 1570
rect 7718 1566 8282 1570
rect 8322 1566 15640 1570
rect 360 1552 15640 1566
rect 360 1516 428 1552
rect 360 1484 378 1516
rect 410 1484 428 1516
rect 15572 1516 15640 1552
rect 360 1448 428 1484
rect 360 1416 378 1448
rect 410 1416 428 1448
rect 360 1380 428 1416
rect 4027 1490 8194 1506
rect 4027 1474 7806 1490
rect 4027 1464 4069 1474
rect 4027 1398 4028 1464
rect 360 1348 378 1380
rect 410 1348 428 1380
rect 360 1312 428 1348
rect 360 1280 378 1312
rect 410 1280 428 1312
rect 3988 1342 4028 1398
rect 4068 1398 4069 1464
rect 7838 1474 8162 1490
rect 7677 1420 7719 1430
rect 4068 1342 4108 1398
rect 3988 1298 4108 1342
rect 360 1244 428 1280
rect 360 1212 378 1244
rect 410 1212 428 1244
rect 360 1176 428 1212
rect 360 1144 378 1176
rect 410 1144 428 1176
rect 360 1108 428 1144
rect 360 1076 378 1108
rect 410 1076 428 1108
rect 360 1040 428 1076
rect 360 1008 378 1040
rect 410 1008 428 1040
rect 360 972 428 1008
rect 360 940 378 972
rect 410 940 428 972
rect 360 904 428 940
rect 360 872 378 904
rect 410 872 428 904
rect 360 836 428 872
rect 360 804 378 836
rect 410 804 428 836
rect 360 768 428 804
rect 360 736 378 768
rect 410 736 428 768
rect 360 700 428 736
rect 360 668 378 700
rect 410 668 428 700
rect 360 632 428 668
rect 360 600 378 632
rect 410 600 428 632
rect 360 564 428 600
rect 360 532 378 564
rect 410 532 428 564
rect 7677 560 7678 1420
rect 7718 560 7719 1420
rect 7677 550 7719 560
rect 360 496 428 532
rect 360 464 378 496
rect 410 464 428 496
rect 7806 522 7838 1458
rect 7938 1420 8062 1430
rect 7938 560 7939 1420
rect 8061 560 8062 1420
rect 7938 550 8062 560
rect 7806 474 7838 490
rect 8162 522 8194 1458
rect 15572 1484 15590 1516
rect 15622 1484 15640 1516
rect 15572 1448 15640 1484
rect 8281 1420 8323 1430
rect 8281 560 8282 1420
rect 8322 560 8323 1420
rect 8281 550 8323 560
rect 15572 1416 15590 1448
rect 15622 1416 15640 1448
rect 15572 1380 15640 1416
rect 15572 1348 15590 1380
rect 15622 1348 15640 1380
rect 15572 1312 15640 1348
rect 15572 1280 15590 1312
rect 15622 1280 15640 1312
rect 15572 1244 15640 1280
rect 15572 1212 15590 1244
rect 15622 1212 15640 1244
rect 15572 1176 15640 1212
rect 15572 1144 15590 1176
rect 15622 1144 15640 1176
rect 15572 1108 15640 1144
rect 15572 1076 15590 1108
rect 15622 1076 15640 1108
rect 15572 1040 15640 1076
rect 15572 1008 15590 1040
rect 15622 1008 15640 1040
rect 15572 972 15640 1008
rect 15572 940 15590 972
rect 15622 940 15640 972
rect 15572 904 15640 940
rect 15572 872 15590 904
rect 15622 872 15640 904
rect 15572 836 15640 872
rect 15572 804 15590 836
rect 15622 804 15640 836
rect 15572 768 15640 804
rect 15572 736 15590 768
rect 15622 736 15640 768
rect 15572 700 15640 736
rect 15572 668 15590 700
rect 15622 668 15640 700
rect 15572 632 15640 668
rect 15572 600 15590 632
rect 15622 600 15640 632
rect 15572 564 15640 600
rect 8162 474 8194 490
rect 15572 532 15590 564
rect 15622 532 15640 564
rect 15572 496 15640 532
rect 360 428 428 464
rect 15572 464 15590 496
rect 15622 464 15640 496
rect 15572 428 15640 464
rect 360 414 15640 428
rect 360 410 7678 414
rect 7718 410 8282 414
rect 8322 410 15640 414
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7718 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8282 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 374 7678 378
rect 7718 374 8282 378
rect 8322 374 15640 378
rect 360 360 15640 374
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 15932 360 16000 396
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 7678 1602 7718 1606
rect 8282 1602 8322 1606
rect 7678 1570 7710 1602
rect 7710 1570 7718 1602
rect 8282 1570 8290 1602
rect 8290 1570 8322 1602
rect 7678 1566 7718 1570
rect 8282 1566 8322 1570
rect 4028 1342 4068 1464
rect 7678 1414 7718 1420
rect 7678 1382 7682 1414
rect 7682 1382 7714 1414
rect 7714 1382 7718 1414
rect 7678 1346 7718 1382
rect 7678 1314 7682 1346
rect 7682 1314 7714 1346
rect 7714 1314 7718 1346
rect 7678 1278 7718 1314
rect 7678 1246 7682 1278
rect 7682 1246 7714 1278
rect 7714 1246 7718 1278
rect 7678 1210 7718 1246
rect 7678 1178 7682 1210
rect 7682 1178 7714 1210
rect 7714 1178 7718 1210
rect 7678 1142 7718 1178
rect 7678 1110 7682 1142
rect 7682 1110 7714 1142
rect 7714 1110 7718 1142
rect 7678 1074 7718 1110
rect 7678 1042 7682 1074
rect 7682 1042 7714 1074
rect 7714 1042 7718 1074
rect 7678 1006 7718 1042
rect 7678 974 7682 1006
rect 7682 974 7714 1006
rect 7714 974 7718 1006
rect 7678 938 7718 974
rect 7678 906 7682 938
rect 7682 906 7714 938
rect 7714 906 7718 938
rect 7678 870 7718 906
rect 7678 838 7682 870
rect 7682 838 7714 870
rect 7714 838 7718 870
rect 7678 802 7718 838
rect 7678 770 7682 802
rect 7682 770 7714 802
rect 7714 770 7718 802
rect 7678 734 7718 770
rect 7678 702 7682 734
rect 7682 702 7714 734
rect 7714 702 7718 734
rect 7678 666 7718 702
rect 7678 634 7682 666
rect 7682 634 7714 666
rect 7714 634 7718 666
rect 7678 598 7718 634
rect 7678 566 7682 598
rect 7682 566 7714 598
rect 7714 566 7718 598
rect 7678 560 7718 566
rect 7939 1414 8061 1420
rect 7939 1382 7984 1414
rect 7984 1382 8016 1414
rect 8016 1382 8061 1414
rect 7939 1346 8061 1382
rect 7939 1314 7984 1346
rect 7984 1314 8016 1346
rect 8016 1314 8061 1346
rect 7939 1278 8061 1314
rect 7939 1246 7984 1278
rect 7984 1246 8016 1278
rect 8016 1246 8061 1278
rect 7939 1210 8061 1246
rect 7939 1178 7984 1210
rect 7984 1178 8016 1210
rect 8016 1178 8061 1210
rect 7939 1142 8061 1178
rect 7939 1110 7984 1142
rect 7984 1110 8016 1142
rect 8016 1110 8061 1142
rect 7939 1074 8061 1110
rect 7939 1042 7984 1074
rect 7984 1042 8016 1074
rect 8016 1042 8061 1074
rect 7939 1006 8061 1042
rect 7939 974 7984 1006
rect 7984 974 8016 1006
rect 8016 974 8061 1006
rect 7939 938 8061 974
rect 7939 906 7984 938
rect 7984 906 8016 938
rect 8016 906 8061 938
rect 7939 870 8061 906
rect 7939 838 7984 870
rect 7984 838 8016 870
rect 8016 838 8061 870
rect 7939 802 8061 838
rect 7939 770 7984 802
rect 7984 770 8016 802
rect 8016 770 8061 802
rect 7939 734 8061 770
rect 7939 702 7984 734
rect 7984 702 8016 734
rect 8016 702 8061 734
rect 7939 666 8061 702
rect 7939 634 7984 666
rect 7984 634 8016 666
rect 8016 634 8061 666
rect 7939 598 8061 634
rect 7939 566 7984 598
rect 7984 566 8016 598
rect 8016 566 8061 598
rect 7939 560 8061 566
rect 8282 1414 8322 1420
rect 8282 1382 8286 1414
rect 8286 1382 8318 1414
rect 8318 1382 8322 1414
rect 8282 1346 8322 1382
rect 8282 1314 8286 1346
rect 8286 1314 8318 1346
rect 8318 1314 8322 1346
rect 8282 1278 8322 1314
rect 8282 1246 8286 1278
rect 8286 1246 8318 1278
rect 8318 1246 8322 1278
rect 8282 1210 8322 1246
rect 8282 1178 8286 1210
rect 8286 1178 8318 1210
rect 8318 1178 8322 1210
rect 8282 1142 8322 1178
rect 8282 1110 8286 1142
rect 8286 1110 8318 1142
rect 8318 1110 8322 1142
rect 8282 1074 8322 1110
rect 8282 1042 8286 1074
rect 8286 1042 8318 1074
rect 8318 1042 8322 1074
rect 8282 1006 8322 1042
rect 8282 974 8286 1006
rect 8286 974 8318 1006
rect 8318 974 8322 1006
rect 8282 938 8322 974
rect 8282 906 8286 938
rect 8286 906 8318 938
rect 8318 906 8322 938
rect 8282 870 8322 906
rect 8282 838 8286 870
rect 8286 838 8318 870
rect 8318 838 8322 870
rect 8282 802 8322 838
rect 8282 770 8286 802
rect 8286 770 8318 802
rect 8318 770 8322 802
rect 8282 734 8322 770
rect 8282 702 8286 734
rect 8286 702 8318 734
rect 8318 702 8322 734
rect 8282 666 8322 702
rect 8282 634 8286 666
rect 8286 634 8318 666
rect 8318 634 8322 666
rect 8282 598 8322 634
rect 8282 566 8286 598
rect 8286 566 8318 598
rect 8318 566 8322 598
rect 8282 560 8322 566
rect 7678 410 7718 414
rect 8282 410 8322 414
rect 7678 378 7710 410
rect 7710 378 7718 410
rect 8282 378 8290 410
rect 8290 378 8322 410
rect 7678 374 7718 378
rect 8282 374 8322 378
<< metal2 >>
rect 4028 1464 4068 1980
rect 4028 1333 4068 1342
rect 7678 1953 7718 1980
rect 7939 1420 8061 1980
rect 7939 551 8061 560
rect 8282 1953 8322 1980
rect 7678 0 7718 27
rect 8282 0 8322 27
<< via2 >>
rect 7678 1606 7718 1953
rect 7678 1566 7718 1606
rect 7678 1420 7718 1566
rect 7678 560 7718 1420
rect 7678 414 7718 560
rect 8282 1606 8322 1953
rect 8282 1566 8322 1606
rect 8282 1420 8322 1566
rect 8282 560 8322 1420
rect 7678 374 7718 414
rect 7678 27 7718 374
rect 8282 414 8322 560
rect 8282 374 8322 414
rect 8282 27 8322 374
<< metal3 >>
rect 7678 1953 7718 1962
rect 7678 18 7718 27
rect 8282 1953 8322 1962
rect 8282 18 8322 27
<< labels >>
rlabel metal2 s 4028 1333 4068 1980 4 gate
port 3 nsew
rlabel metal2 s 7939 551 8061 1980 4 pad
port 2 nsew
rlabel comment s 394 394 394 394 4 sub!
flabel comment s 4048 1348 4048 1348 0 FreeSans 400 0 0 0 dant
flabel metal1 s 560 1560 834 1608 0 FreeSans 51 0 0 0 iovss
port 1 nsew
<< properties >>
string device primitive
string GDS_END 22786084
string GDS_FILE sg13g2_io.gds
string GDS_START 22710056
<< end >>
