magic
tech ihp-sg13g2
timestamp 1753041618
<< error_p >>
rect -18 3030 -13 3035
rect 13 3030 18 3035
rect 121 3030 126 3035
rect 152 3030 157 3035
rect 260 3030 265 3035
rect 291 3030 296 3035
rect 399 3030 404 3035
rect 430 3030 435 3035
rect 538 3030 543 3035
rect 569 3030 574 3035
rect 677 3030 682 3035
rect 708 3030 713 3035
rect 816 3030 821 3035
rect 847 3030 852 3035
rect 955 3030 960 3035
rect 986 3030 991 3035
rect 1094 3030 1099 3035
rect 1125 3030 1130 3035
rect 1233 3030 1238 3035
rect 1264 3030 1269 3035
rect 1372 3030 1377 3035
rect 1403 3030 1408 3035
rect 1511 3030 1516 3035
rect 1542 3030 1547 3035
rect 1650 3030 1655 3035
rect 1681 3030 1686 3035
rect 1789 3030 1794 3035
rect 1820 3030 1825 3035
rect 1928 3030 1933 3035
rect 1959 3030 1964 3035
rect -23 3025 23 3030
rect 116 3025 162 3030
rect 255 3025 301 3030
rect 394 3025 440 3030
rect 533 3025 579 3030
rect 672 3025 718 3030
rect 811 3025 857 3030
rect 950 3025 996 3030
rect 1089 3025 1135 3030
rect 1228 3025 1274 3030
rect 1367 3025 1413 3030
rect 1506 3025 1552 3030
rect 1645 3025 1691 3030
rect 1784 3025 1830 3030
rect 1923 3025 1969 3030
rect -18 3019 18 3025
rect 121 3019 157 3025
rect 260 3019 296 3025
rect 399 3019 435 3025
rect 538 3019 574 3025
rect 677 3019 713 3025
rect 816 3019 852 3025
rect 955 3019 991 3025
rect 1094 3019 1130 3025
rect 1233 3019 1269 3025
rect 1372 3019 1408 3025
rect 1511 3019 1547 3025
rect 1650 3019 1686 3025
rect 1789 3019 1825 3025
rect 1928 3019 1964 3025
rect -23 3014 23 3019
rect 116 3014 162 3019
rect 255 3014 301 3019
rect 394 3014 440 3019
rect 533 3014 579 3019
rect 672 3014 718 3019
rect 811 3014 857 3019
rect 950 3014 996 3019
rect 1089 3014 1135 3019
rect 1228 3014 1274 3019
rect 1367 3014 1413 3019
rect 1506 3014 1552 3019
rect 1645 3014 1691 3019
rect 1784 3014 1830 3019
rect 1923 3014 1969 3019
rect -18 3009 -13 3014
rect 13 3009 18 3014
rect 121 3009 126 3014
rect 152 3009 157 3014
rect 260 3009 265 3014
rect 291 3009 296 3014
rect 399 3009 404 3014
rect 430 3009 435 3014
rect 538 3009 543 3014
rect 569 3009 574 3014
rect 677 3009 682 3014
rect 708 3009 713 3014
rect 816 3009 821 3014
rect 847 3009 852 3014
rect 955 3009 960 3014
rect 986 3009 991 3014
rect 1094 3009 1099 3014
rect 1125 3009 1130 3014
rect 1233 3009 1238 3014
rect 1264 3009 1269 3014
rect 1372 3009 1377 3014
rect 1403 3009 1408 3014
rect 1511 3009 1516 3014
rect 1542 3009 1547 3014
rect 1650 3009 1655 3014
rect 1681 3009 1686 3014
rect 1789 3009 1794 3014
rect 1820 3009 1825 3014
rect 1928 3009 1933 3014
rect 1959 3009 1964 3014
rect -52 2993 -47 2998
rect -41 2993 -36 2998
rect 36 2993 41 2998
rect 47 2993 52 2998
rect 87 2993 92 2998
rect 98 2993 103 2998
rect 175 2993 180 2998
rect 186 2993 191 2998
rect 226 2993 231 2998
rect 237 2993 242 2998
rect 314 2993 319 2998
rect 325 2993 330 2998
rect 365 2993 370 2998
rect 376 2993 381 2998
rect 453 2993 458 2998
rect 464 2993 469 2998
rect 504 2993 509 2998
rect 515 2993 520 2998
rect 592 2993 597 2998
rect 603 2993 608 2998
rect 643 2993 648 2998
rect 654 2993 659 2998
rect 731 2993 736 2998
rect 742 2993 747 2998
rect 782 2993 787 2998
rect 793 2993 798 2998
rect 870 2993 875 2998
rect 881 2993 886 2998
rect 921 2993 926 2998
rect 932 2993 937 2998
rect 1009 2993 1014 2998
rect 1020 2993 1025 2998
rect 1060 2993 1065 2998
rect 1071 2993 1076 2998
rect 1148 2993 1153 2998
rect 1159 2993 1164 2998
rect 1199 2993 1204 2998
rect 1210 2993 1215 2998
rect 1287 2993 1292 2998
rect 1298 2993 1303 2998
rect 1338 2993 1343 2998
rect 1349 2993 1354 2998
rect 1426 2993 1431 2998
rect 1437 2993 1442 2998
rect 1477 2993 1482 2998
rect 1488 2993 1493 2998
rect 1565 2993 1570 2998
rect 1576 2993 1581 2998
rect 1616 2993 1621 2998
rect 1627 2993 1632 2998
rect 1704 2993 1709 2998
rect 1715 2993 1720 2998
rect 1755 2993 1760 2998
rect 1766 2993 1771 2998
rect 1843 2993 1848 2998
rect 1854 2993 1859 2998
rect 1894 2993 1899 2998
rect 1905 2993 1910 2998
rect 1982 2993 1987 2998
rect 1993 2993 1998 2998
rect -57 2988 -52 2993
rect -36 2988 -31 2993
rect 31 2988 36 2993
rect 52 2988 57 2993
rect 82 2988 87 2993
rect 103 2988 108 2993
rect 170 2988 175 2993
rect 191 2988 196 2993
rect 221 2988 226 2993
rect 242 2988 247 2993
rect 309 2988 314 2993
rect 330 2988 335 2993
rect 360 2988 365 2993
rect 381 2988 386 2993
rect 448 2988 453 2993
rect 469 2988 474 2993
rect 499 2988 504 2993
rect 520 2988 525 2993
rect 587 2988 592 2993
rect 608 2988 613 2993
rect 638 2988 643 2993
rect 659 2988 664 2993
rect 726 2988 731 2993
rect 747 2988 752 2993
rect 777 2988 782 2993
rect 798 2988 803 2993
rect 865 2988 870 2993
rect 886 2988 891 2993
rect 916 2988 921 2993
rect 937 2988 942 2993
rect 1004 2988 1009 2993
rect 1025 2988 1030 2993
rect 1055 2988 1060 2993
rect 1076 2988 1081 2993
rect 1143 2988 1148 2993
rect 1164 2988 1169 2993
rect 1194 2988 1199 2993
rect 1215 2988 1220 2993
rect 1282 2988 1287 2993
rect 1303 2988 1308 2993
rect 1333 2988 1338 2993
rect 1354 2988 1359 2993
rect 1421 2988 1426 2993
rect 1442 2988 1447 2993
rect 1472 2988 1477 2993
rect 1493 2988 1498 2993
rect 1560 2988 1565 2993
rect 1581 2988 1586 2993
rect 1611 2988 1616 2993
rect 1632 2988 1637 2993
rect 1699 2988 1704 2993
rect 1720 2988 1725 2993
rect 1750 2988 1755 2993
rect 1771 2988 1776 2993
rect 1838 2988 1843 2993
rect 1859 2988 1864 2993
rect 1889 2988 1894 2993
rect 1910 2988 1915 2993
rect 1977 2988 1982 2993
rect 1998 2988 2003 2993
rect -57 -2993 -52 -2988
rect -36 -2993 -31 -2988
rect 31 -2993 36 -2988
rect 52 -2993 57 -2988
rect 82 -2993 87 -2988
rect 103 -2993 108 -2988
rect 170 -2993 175 -2988
rect 191 -2993 196 -2988
rect 221 -2993 226 -2988
rect 242 -2993 247 -2988
rect 309 -2993 314 -2988
rect 330 -2993 335 -2988
rect 360 -2993 365 -2988
rect 381 -2993 386 -2988
rect 448 -2993 453 -2988
rect 469 -2993 474 -2988
rect 499 -2993 504 -2988
rect 520 -2993 525 -2988
rect 587 -2993 592 -2988
rect 608 -2993 613 -2988
rect 638 -2993 643 -2988
rect 659 -2993 664 -2988
rect 726 -2993 731 -2988
rect 747 -2993 752 -2988
rect 777 -2993 782 -2988
rect 798 -2993 803 -2988
rect 865 -2993 870 -2988
rect 886 -2993 891 -2988
rect 916 -2993 921 -2988
rect 937 -2993 942 -2988
rect 1004 -2993 1009 -2988
rect 1025 -2993 1030 -2988
rect 1055 -2993 1060 -2988
rect 1076 -2993 1081 -2988
rect 1143 -2993 1148 -2988
rect 1164 -2993 1169 -2988
rect 1194 -2993 1199 -2988
rect 1215 -2993 1220 -2988
rect 1282 -2993 1287 -2988
rect 1303 -2993 1308 -2988
rect 1333 -2993 1338 -2988
rect 1354 -2993 1359 -2988
rect 1421 -2993 1426 -2988
rect 1442 -2993 1447 -2988
rect 1472 -2993 1477 -2988
rect 1493 -2993 1498 -2988
rect 1560 -2993 1565 -2988
rect 1581 -2993 1586 -2988
rect 1611 -2993 1616 -2988
rect 1632 -2993 1637 -2988
rect 1699 -2993 1704 -2988
rect 1720 -2993 1725 -2988
rect 1750 -2993 1755 -2988
rect 1771 -2993 1776 -2988
rect 1838 -2993 1843 -2988
rect 1859 -2993 1864 -2988
rect 1889 -2993 1894 -2988
rect 1910 -2993 1915 -2988
rect 1977 -2993 1982 -2988
rect 1998 -2993 2003 -2988
rect -52 -2998 -47 -2993
rect -41 -2998 -36 -2993
rect 36 -2998 41 -2993
rect 47 -2998 52 -2993
rect 87 -2998 92 -2993
rect 98 -2998 103 -2993
rect 175 -2998 180 -2993
rect 186 -2998 191 -2993
rect 226 -2998 231 -2993
rect 237 -2998 242 -2993
rect 314 -2998 319 -2993
rect 325 -2998 330 -2993
rect 365 -2998 370 -2993
rect 376 -2998 381 -2993
rect 453 -2998 458 -2993
rect 464 -2998 469 -2993
rect 504 -2998 509 -2993
rect 515 -2998 520 -2993
rect 592 -2998 597 -2993
rect 603 -2998 608 -2993
rect 643 -2998 648 -2993
rect 654 -2998 659 -2993
rect 731 -2998 736 -2993
rect 742 -2998 747 -2993
rect 782 -2998 787 -2993
rect 793 -2998 798 -2993
rect 870 -2998 875 -2993
rect 881 -2998 886 -2993
rect 921 -2998 926 -2993
rect 932 -2998 937 -2993
rect 1009 -2998 1014 -2993
rect 1020 -2998 1025 -2993
rect 1060 -2998 1065 -2993
rect 1071 -2998 1076 -2993
rect 1148 -2998 1153 -2993
rect 1159 -2998 1164 -2993
rect 1199 -2998 1204 -2993
rect 1210 -2998 1215 -2993
rect 1287 -2998 1292 -2993
rect 1298 -2998 1303 -2993
rect 1338 -2998 1343 -2993
rect 1349 -2998 1354 -2993
rect 1426 -2998 1431 -2993
rect 1437 -2998 1442 -2993
rect 1477 -2998 1482 -2993
rect 1488 -2998 1493 -2993
rect 1565 -2998 1570 -2993
rect 1576 -2998 1581 -2993
rect 1616 -2998 1621 -2993
rect 1627 -2998 1632 -2993
rect 1704 -2998 1709 -2993
rect 1715 -2998 1720 -2993
rect 1755 -2998 1760 -2993
rect 1766 -2998 1771 -2993
rect 1843 -2998 1848 -2993
rect 1854 -2998 1859 -2993
rect 1894 -2998 1899 -2993
rect 1905 -2998 1910 -2993
rect 1982 -2998 1987 -2993
rect 1993 -2998 1998 -2993
rect -18 -3014 -13 -3009
rect 13 -3014 18 -3009
rect 121 -3014 126 -3009
rect 152 -3014 157 -3009
rect 260 -3014 265 -3009
rect 291 -3014 296 -3009
rect 399 -3014 404 -3009
rect 430 -3014 435 -3009
rect 538 -3014 543 -3009
rect 569 -3014 574 -3009
rect 677 -3014 682 -3009
rect 708 -3014 713 -3009
rect 816 -3014 821 -3009
rect 847 -3014 852 -3009
rect 955 -3014 960 -3009
rect 986 -3014 991 -3009
rect 1094 -3014 1099 -3009
rect 1125 -3014 1130 -3009
rect 1233 -3014 1238 -3009
rect 1264 -3014 1269 -3009
rect 1372 -3014 1377 -3009
rect 1403 -3014 1408 -3009
rect 1511 -3014 1516 -3009
rect 1542 -3014 1547 -3009
rect 1650 -3014 1655 -3009
rect 1681 -3014 1686 -3009
rect 1789 -3014 1794 -3009
rect 1820 -3014 1825 -3009
rect 1928 -3014 1933 -3009
rect 1959 -3014 1964 -3009
rect -23 -3019 23 -3014
rect 116 -3019 162 -3014
rect 255 -3019 301 -3014
rect 394 -3019 440 -3014
rect 533 -3019 579 -3014
rect 672 -3019 718 -3014
rect 811 -3019 857 -3014
rect 950 -3019 996 -3014
rect 1089 -3019 1135 -3014
rect 1228 -3019 1274 -3014
rect 1367 -3019 1413 -3014
rect 1506 -3019 1552 -3014
rect 1645 -3019 1691 -3014
rect 1784 -3019 1830 -3014
rect 1923 -3019 1969 -3014
rect -18 -3025 18 -3019
rect 121 -3025 157 -3019
rect 260 -3025 296 -3019
rect 399 -3025 435 -3019
rect 538 -3025 574 -3019
rect 677 -3025 713 -3019
rect 816 -3025 852 -3019
rect 955 -3025 991 -3019
rect 1094 -3025 1130 -3019
rect 1233 -3025 1269 -3019
rect 1372 -3025 1408 -3019
rect 1511 -3025 1547 -3019
rect 1650 -3025 1686 -3019
rect 1789 -3025 1825 -3019
rect 1928 -3025 1964 -3019
rect -23 -3030 23 -3025
rect 116 -3030 162 -3025
rect 255 -3030 301 -3025
rect 394 -3030 440 -3025
rect 533 -3030 579 -3025
rect 672 -3030 718 -3025
rect 811 -3030 857 -3025
rect 950 -3030 996 -3025
rect 1089 -3030 1135 -3025
rect 1228 -3030 1274 -3025
rect 1367 -3030 1413 -3025
rect 1506 -3030 1552 -3025
rect 1645 -3030 1691 -3025
rect 1784 -3030 1830 -3025
rect 1923 -3030 1969 -3025
rect -18 -3035 -13 -3030
rect 13 -3035 18 -3030
rect 121 -3035 126 -3030
rect 152 -3035 157 -3030
rect 260 -3035 265 -3030
rect 291 -3035 296 -3030
rect 399 -3035 404 -3030
rect 430 -3035 435 -3030
rect 538 -3035 543 -3030
rect 569 -3035 574 -3030
rect 677 -3035 682 -3030
rect 708 -3035 713 -3030
rect 816 -3035 821 -3030
rect 847 -3035 852 -3030
rect 955 -3035 960 -3030
rect 986 -3035 991 -3030
rect 1094 -3035 1099 -3030
rect 1125 -3035 1130 -3030
rect 1233 -3035 1238 -3030
rect 1264 -3035 1269 -3030
rect 1372 -3035 1377 -3030
rect 1403 -3035 1408 -3030
rect 1511 -3035 1516 -3030
rect 1542 -3035 1547 -3030
rect 1650 -3035 1655 -3030
rect 1681 -3035 1686 -3030
rect 1789 -3035 1794 -3030
rect 1820 -3035 1825 -3030
rect 1928 -3035 1933 -3030
rect 1959 -3035 1964 -3030
<< nwell >>
rect -259 -3173 2205 3173
<< hvpmos >>
rect -25 -3000 25 3000
rect 114 -3000 164 3000
rect 253 -3000 303 3000
rect 392 -3000 442 3000
rect 531 -3000 581 3000
rect 670 -3000 720 3000
rect 809 -3000 859 3000
rect 948 -3000 998 3000
rect 1087 -3000 1137 3000
rect 1226 -3000 1276 3000
rect 1365 -3000 1415 3000
rect 1504 -3000 1554 3000
rect 1643 -3000 1693 3000
rect 1782 -3000 1832 3000
rect 1921 -3000 1971 3000
<< hvpdiff >>
rect -59 2993 -25 3000
rect -59 -2993 -52 2993
rect -36 -2993 -25 2993
rect -59 -3000 -25 -2993
rect 25 2993 59 3000
rect 25 -2993 36 2993
rect 52 -2993 59 2993
rect 25 -3000 59 -2993
rect 80 2993 114 3000
rect 80 -2993 87 2993
rect 103 -2993 114 2993
rect 80 -3000 114 -2993
rect 164 2993 198 3000
rect 164 -2993 175 2993
rect 191 -2993 198 2993
rect 164 -3000 198 -2993
rect 219 2993 253 3000
rect 219 -2993 226 2993
rect 242 -2993 253 2993
rect 219 -3000 253 -2993
rect 303 2993 337 3000
rect 303 -2993 314 2993
rect 330 -2993 337 2993
rect 303 -3000 337 -2993
rect 358 2993 392 3000
rect 358 -2993 365 2993
rect 381 -2993 392 2993
rect 358 -3000 392 -2993
rect 442 2993 476 3000
rect 442 -2993 453 2993
rect 469 -2993 476 2993
rect 442 -3000 476 -2993
rect 497 2993 531 3000
rect 497 -2993 504 2993
rect 520 -2993 531 2993
rect 497 -3000 531 -2993
rect 581 2993 615 3000
rect 581 -2993 592 2993
rect 608 -2993 615 2993
rect 581 -3000 615 -2993
rect 636 2993 670 3000
rect 636 -2993 643 2993
rect 659 -2993 670 2993
rect 636 -3000 670 -2993
rect 720 2993 754 3000
rect 720 -2993 731 2993
rect 747 -2993 754 2993
rect 720 -3000 754 -2993
rect 775 2993 809 3000
rect 775 -2993 782 2993
rect 798 -2993 809 2993
rect 775 -3000 809 -2993
rect 859 2993 893 3000
rect 859 -2993 870 2993
rect 886 -2993 893 2993
rect 859 -3000 893 -2993
rect 914 2993 948 3000
rect 914 -2993 921 2993
rect 937 -2993 948 2993
rect 914 -3000 948 -2993
rect 998 2993 1032 3000
rect 998 -2993 1009 2993
rect 1025 -2993 1032 2993
rect 998 -3000 1032 -2993
rect 1053 2993 1087 3000
rect 1053 -2993 1060 2993
rect 1076 -2993 1087 2993
rect 1053 -3000 1087 -2993
rect 1137 2993 1171 3000
rect 1137 -2993 1148 2993
rect 1164 -2993 1171 2993
rect 1137 -3000 1171 -2993
rect 1192 2993 1226 3000
rect 1192 -2993 1199 2993
rect 1215 -2993 1226 2993
rect 1192 -3000 1226 -2993
rect 1276 2993 1310 3000
rect 1276 -2993 1287 2993
rect 1303 -2993 1310 2993
rect 1276 -3000 1310 -2993
rect 1331 2993 1365 3000
rect 1331 -2993 1338 2993
rect 1354 -2993 1365 2993
rect 1331 -3000 1365 -2993
rect 1415 2993 1449 3000
rect 1415 -2993 1426 2993
rect 1442 -2993 1449 2993
rect 1415 -3000 1449 -2993
rect 1470 2993 1504 3000
rect 1470 -2993 1477 2993
rect 1493 -2993 1504 2993
rect 1470 -3000 1504 -2993
rect 1554 2993 1588 3000
rect 1554 -2993 1565 2993
rect 1581 -2993 1588 2993
rect 1554 -3000 1588 -2993
rect 1609 2993 1643 3000
rect 1609 -2993 1616 2993
rect 1632 -2993 1643 2993
rect 1609 -3000 1643 -2993
rect 1693 2993 1727 3000
rect 1693 -2993 1704 2993
rect 1720 -2993 1727 2993
rect 1693 -3000 1727 -2993
rect 1748 2993 1782 3000
rect 1748 -2993 1755 2993
rect 1771 -2993 1782 2993
rect 1748 -3000 1782 -2993
rect 1832 2993 1866 3000
rect 1832 -2993 1843 2993
rect 1859 -2993 1866 2993
rect 1832 -3000 1866 -2993
rect 1887 2993 1921 3000
rect 1887 -2993 1894 2993
rect 1910 -2993 1921 2993
rect 1887 -3000 1921 -2993
rect 1971 2993 2005 3000
rect 1971 -2993 1982 2993
rect 1998 -2993 2005 2993
rect 1971 -3000 2005 -2993
<< hvpdiffc >>
rect -52 -2993 -36 2993
rect 36 -2993 52 2993
rect 87 -2993 103 2993
rect 175 -2993 191 2993
rect 226 -2993 242 2993
rect 314 -2993 330 2993
rect 365 -2993 381 2993
rect 453 -2993 469 2993
rect 504 -2993 520 2993
rect 592 -2993 608 2993
rect 643 -2993 659 2993
rect 731 -2993 747 2993
rect 782 -2993 798 2993
rect 870 -2993 886 2993
rect 921 -2993 937 2993
rect 1009 -2993 1025 2993
rect 1060 -2993 1076 2993
rect 1148 -2993 1164 2993
rect 1199 -2993 1215 2993
rect 1287 -2993 1303 2993
rect 1338 -2993 1354 2993
rect 1426 -2993 1442 2993
rect 1477 -2993 1493 2993
rect 1565 -2993 1581 2993
rect 1616 -2993 1632 2993
rect 1704 -2993 1720 2993
rect 1755 -2993 1771 2993
rect 1843 -2993 1859 2993
rect 1894 -2993 1910 2993
rect 1982 -2993 1998 2993
<< nsubdiff >>
rect -197 3104 2143 3111
rect -197 3088 -160 3104
rect 2106 3088 2143 3104
rect -197 3081 2143 3088
rect -197 3074 -167 3081
rect -197 -3074 -190 3074
rect -174 -3074 -167 3074
rect 2113 3074 2143 3081
rect -197 -3081 -167 -3074
rect 2113 -3074 2120 3074
rect 2136 -3074 2143 3074
rect 2113 -3081 2143 -3074
rect -197 -3088 2143 -3081
rect -197 -3104 -160 -3088
rect 2106 -3104 2143 -3088
rect -197 -3111 2143 -3104
<< nsubdiffcont >>
rect -160 3088 2106 3104
rect -190 -3074 -174 3074
rect 2120 -3074 2136 3074
rect -160 -3104 2106 -3088
<< poly >>
rect -25 3030 25 3037
rect -25 3014 -18 3030
rect 18 3014 25 3030
rect -25 3000 25 3014
rect 114 3030 164 3037
rect 114 3014 121 3030
rect 157 3014 164 3030
rect 114 3000 164 3014
rect 253 3030 303 3037
rect 253 3014 260 3030
rect 296 3014 303 3030
rect 253 3000 303 3014
rect 392 3030 442 3037
rect 392 3014 399 3030
rect 435 3014 442 3030
rect 392 3000 442 3014
rect 531 3030 581 3037
rect 531 3014 538 3030
rect 574 3014 581 3030
rect 531 3000 581 3014
rect 670 3030 720 3037
rect 670 3014 677 3030
rect 713 3014 720 3030
rect 670 3000 720 3014
rect 809 3030 859 3037
rect 809 3014 816 3030
rect 852 3014 859 3030
rect 809 3000 859 3014
rect 948 3030 998 3037
rect 948 3014 955 3030
rect 991 3014 998 3030
rect 948 3000 998 3014
rect 1087 3030 1137 3037
rect 1087 3014 1094 3030
rect 1130 3014 1137 3030
rect 1087 3000 1137 3014
rect 1226 3030 1276 3037
rect 1226 3014 1233 3030
rect 1269 3014 1276 3030
rect 1226 3000 1276 3014
rect 1365 3030 1415 3037
rect 1365 3014 1372 3030
rect 1408 3014 1415 3030
rect 1365 3000 1415 3014
rect 1504 3030 1554 3037
rect 1504 3014 1511 3030
rect 1547 3014 1554 3030
rect 1504 3000 1554 3014
rect 1643 3030 1693 3037
rect 1643 3014 1650 3030
rect 1686 3014 1693 3030
rect 1643 3000 1693 3014
rect 1782 3030 1832 3037
rect 1782 3014 1789 3030
rect 1825 3014 1832 3030
rect 1782 3000 1832 3014
rect 1921 3030 1971 3037
rect 1921 3014 1928 3030
rect 1964 3014 1971 3030
rect 1921 3000 1971 3014
rect -25 -3014 25 -3000
rect -25 -3030 -18 -3014
rect 18 -3030 25 -3014
rect -25 -3037 25 -3030
rect 114 -3014 164 -3000
rect 114 -3030 121 -3014
rect 157 -3030 164 -3014
rect 114 -3037 164 -3030
rect 253 -3014 303 -3000
rect 253 -3030 260 -3014
rect 296 -3030 303 -3014
rect 253 -3037 303 -3030
rect 392 -3014 442 -3000
rect 392 -3030 399 -3014
rect 435 -3030 442 -3014
rect 392 -3037 442 -3030
rect 531 -3014 581 -3000
rect 531 -3030 538 -3014
rect 574 -3030 581 -3014
rect 531 -3037 581 -3030
rect 670 -3014 720 -3000
rect 670 -3030 677 -3014
rect 713 -3030 720 -3014
rect 670 -3037 720 -3030
rect 809 -3014 859 -3000
rect 809 -3030 816 -3014
rect 852 -3030 859 -3014
rect 809 -3037 859 -3030
rect 948 -3014 998 -3000
rect 948 -3030 955 -3014
rect 991 -3030 998 -3014
rect 948 -3037 998 -3030
rect 1087 -3014 1137 -3000
rect 1087 -3030 1094 -3014
rect 1130 -3030 1137 -3014
rect 1087 -3037 1137 -3030
rect 1226 -3014 1276 -3000
rect 1226 -3030 1233 -3014
rect 1269 -3030 1276 -3014
rect 1226 -3037 1276 -3030
rect 1365 -3014 1415 -3000
rect 1365 -3030 1372 -3014
rect 1408 -3030 1415 -3014
rect 1365 -3037 1415 -3030
rect 1504 -3014 1554 -3000
rect 1504 -3030 1511 -3014
rect 1547 -3030 1554 -3014
rect 1504 -3037 1554 -3030
rect 1643 -3014 1693 -3000
rect 1643 -3030 1650 -3014
rect 1686 -3030 1693 -3014
rect 1643 -3037 1693 -3030
rect 1782 -3014 1832 -3000
rect 1782 -3030 1789 -3014
rect 1825 -3030 1832 -3014
rect 1782 -3037 1832 -3030
rect 1921 -3014 1971 -3000
rect 1921 -3030 1928 -3014
rect 1964 -3030 1971 -3014
rect 1921 -3037 1971 -3030
<< polycont >>
rect -18 3014 18 3030
rect 121 3014 157 3030
rect 260 3014 296 3030
rect 399 3014 435 3030
rect 538 3014 574 3030
rect 677 3014 713 3030
rect 816 3014 852 3030
rect 955 3014 991 3030
rect 1094 3014 1130 3030
rect 1233 3014 1269 3030
rect 1372 3014 1408 3030
rect 1511 3014 1547 3030
rect 1650 3014 1686 3030
rect 1789 3014 1825 3030
rect 1928 3014 1964 3030
rect -18 -3030 18 -3014
rect 121 -3030 157 -3014
rect 260 -3030 296 -3014
rect 399 -3030 435 -3014
rect 538 -3030 574 -3014
rect 677 -3030 713 -3014
rect 816 -3030 852 -3014
rect 955 -3030 991 -3014
rect 1094 -3030 1130 -3014
rect 1233 -3030 1269 -3014
rect 1372 -3030 1408 -3014
rect 1511 -3030 1547 -3014
rect 1650 -3030 1686 -3014
rect 1789 -3030 1825 -3014
rect 1928 -3030 1964 -3014
<< metal1 >>
rect -195 3104 2141 3109
rect -195 3088 -160 3104
rect 2106 3088 2141 3104
rect -195 3083 2141 3088
rect -195 3074 -169 3083
rect -195 -3074 -190 3074
rect -174 -3074 -169 3074
rect 2115 3074 2141 3083
rect -195 -3083 -169 -3074
rect 2115 -3074 2120 3074
rect 2136 -3074 2141 3074
rect 2115 -3083 2141 -3074
rect -195 -3088 2141 -3083
rect -195 -3104 -160 -3088
rect 2106 -3104 2141 -3088
rect -195 -3109 2141 -3104
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 60 l 0.5 nf 1 nx 15 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 2 glc 1 grc 1 gtc 1 gbc 1
<< end >>
