magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect -4 56 726 285
rect -26 -56 794 56
<< nmos >>
rect 90 149 116 259
rect 298 115 324 259
rect 400 115 426 259
rect 504 115 530 259
rect 606 115 632 259
<< pmos >>
rect 90 412 116 580
rect 298 412 324 636
rect 400 412 426 636
rect 504 412 530 636
rect 606 412 632 636
<< ndiff >>
rect 22 245 90 259
rect 22 213 36 245
rect 68 213 90 245
rect 22 149 90 213
rect 116 245 184 259
rect 116 213 138 245
rect 170 213 184 245
rect 116 149 184 213
rect 226 230 298 259
rect 226 198 241 230
rect 273 198 298 230
rect 226 162 298 198
rect 226 130 242 162
rect 274 130 298 162
rect 226 115 298 130
rect 324 161 400 259
rect 324 129 346 161
rect 378 129 400 161
rect 324 115 400 129
rect 426 233 504 259
rect 426 201 448 233
rect 480 201 504 233
rect 426 164 504 201
rect 426 132 448 164
rect 480 132 504 164
rect 426 115 504 132
rect 530 242 606 259
rect 530 210 552 242
rect 584 210 606 242
rect 530 115 606 210
rect 632 230 700 259
rect 632 198 654 230
rect 686 198 700 230
rect 632 162 700 198
rect 632 130 654 162
rect 686 130 700 162
rect 632 115 700 130
<< pdiff >>
rect 226 622 298 636
rect 226 590 240 622
rect 272 590 298 622
rect 22 566 90 580
rect 22 534 36 566
rect 68 534 90 566
rect 22 498 90 534
rect 22 466 36 498
rect 68 466 90 498
rect 22 412 90 466
rect 116 566 184 580
rect 116 534 138 566
rect 170 534 184 566
rect 116 498 184 534
rect 116 466 138 498
rect 170 466 184 498
rect 116 412 184 466
rect 226 554 298 590
rect 226 522 240 554
rect 272 522 298 554
rect 226 486 298 522
rect 226 454 240 486
rect 272 454 298 486
rect 226 412 298 454
rect 324 622 400 636
rect 324 590 346 622
rect 378 590 400 622
rect 324 554 400 590
rect 324 522 346 554
rect 378 522 400 554
rect 324 486 400 522
rect 324 454 346 486
rect 378 454 400 486
rect 324 412 400 454
rect 426 622 504 636
rect 426 590 448 622
rect 480 590 504 622
rect 426 554 504 590
rect 426 522 448 554
rect 480 522 504 554
rect 426 412 504 522
rect 530 622 606 636
rect 530 590 552 622
rect 584 590 606 622
rect 530 554 606 590
rect 530 522 552 554
rect 584 522 606 554
rect 530 486 606 522
rect 530 454 552 486
rect 584 454 606 486
rect 530 412 606 454
rect 632 622 702 636
rect 632 590 654 622
rect 686 590 702 622
rect 632 554 702 590
rect 632 522 654 554
rect 686 522 702 554
rect 632 486 702 522
rect 632 454 654 486
rect 686 454 702 486
rect 632 412 702 454
<< ndiffc >>
rect 36 213 68 245
rect 138 213 170 245
rect 241 198 273 230
rect 242 130 274 162
rect 346 129 378 161
rect 448 201 480 233
rect 448 132 480 164
rect 552 210 584 242
rect 654 198 686 230
rect 654 130 686 162
<< pdiffc >>
rect 240 590 272 622
rect 36 534 68 566
rect 36 466 68 498
rect 138 534 170 566
rect 138 466 170 498
rect 240 522 272 554
rect 240 454 272 486
rect 346 590 378 622
rect 346 522 378 554
rect 346 454 378 486
rect 448 590 480 622
rect 448 522 480 554
rect 552 590 584 622
rect 552 522 584 554
rect 552 454 584 486
rect 654 590 686 622
rect 654 522 686 554
rect 654 454 686 486
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 298 636 324 672
rect 400 636 426 672
rect 504 636 530 672
rect 606 636 632 672
rect 90 580 116 616
rect 90 366 116 412
rect 298 373 324 412
rect 66 352 126 366
rect 66 320 80 352
rect 112 320 126 352
rect 66 306 126 320
rect 238 359 324 373
rect 400 359 426 412
rect 504 373 530 412
rect 238 327 252 359
rect 284 327 426 359
rect 238 313 426 327
rect 462 359 530 373
rect 606 359 632 412
rect 462 327 476 359
rect 508 327 632 359
rect 462 313 632 327
rect 90 259 116 306
rect 298 259 324 313
rect 400 259 426 313
rect 504 259 530 313
rect 606 259 632 313
rect 90 113 116 149
rect 298 79 324 115
rect 400 79 426 115
rect 504 79 530 115
rect 606 79 632 115
<< polycont >>
rect 80 320 112 352
rect 252 327 284 359
rect 476 327 508 359
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 26 566 78 712
rect 230 622 282 712
rect 230 590 240 622
rect 272 590 282 622
rect 26 534 36 566
rect 68 534 78 566
rect 26 498 78 534
rect 26 466 36 498
rect 68 466 78 498
rect 26 456 78 466
rect 128 566 180 576
rect 128 534 138 566
rect 170 534 180 566
rect 128 498 180 534
rect 128 466 138 498
rect 170 468 180 498
rect 230 554 282 590
rect 230 522 240 554
rect 272 522 282 554
rect 230 486 282 522
rect 170 466 193 468
rect 128 442 193 466
rect 31 352 122 373
rect 31 320 80 352
rect 112 320 122 352
rect 31 295 122 320
rect 161 369 193 442
rect 230 454 240 486
rect 272 454 282 486
rect 230 425 282 454
rect 336 622 388 632
rect 336 590 346 622
rect 378 590 388 622
rect 336 554 388 590
rect 336 522 346 554
rect 378 522 388 554
rect 336 486 388 522
rect 438 622 490 712
rect 438 590 448 622
rect 480 590 490 622
rect 438 554 490 590
rect 438 522 448 554
rect 480 522 490 554
rect 438 512 490 522
rect 542 622 600 636
rect 542 590 552 622
rect 584 590 600 622
rect 542 554 600 590
rect 542 522 552 554
rect 584 522 600 554
rect 336 454 346 486
rect 378 472 388 486
rect 542 486 600 522
rect 542 472 552 486
rect 378 454 552 472
rect 584 454 600 486
rect 336 440 600 454
rect 644 622 696 712
rect 644 590 654 622
rect 686 590 696 622
rect 644 554 696 590
rect 644 522 654 554
rect 686 522 696 554
rect 644 486 696 522
rect 644 454 654 486
rect 686 454 696 486
rect 644 444 696 454
rect 161 359 294 369
rect 161 327 252 359
rect 284 327 294 359
rect 161 317 294 327
rect 432 359 518 369
rect 432 327 476 359
rect 508 327 518 359
rect 161 255 193 317
rect 432 307 518 327
rect 554 278 600 440
rect 26 245 78 255
rect 26 213 36 245
rect 68 213 78 245
rect 26 44 78 213
rect 128 245 193 255
rect 128 213 138 245
rect 170 213 193 245
rect 542 242 600 278
rect 128 203 193 213
rect 231 233 490 240
rect 231 230 448 233
rect 231 198 241 230
rect 273 207 448 230
rect 273 198 283 207
rect 231 162 283 198
rect 436 201 448 207
rect 480 201 490 233
rect 231 130 242 162
rect 274 130 283 162
rect 231 120 283 130
rect 336 161 388 171
rect 336 129 346 161
rect 378 129 388 161
rect 336 44 388 129
rect 436 164 490 201
rect 542 210 552 242
rect 584 210 600 242
rect 542 200 600 210
rect 640 230 696 240
rect 436 132 448 164
rect 480 152 490 164
rect 640 198 654 230
rect 686 198 696 230
rect 640 162 696 198
rect 640 152 654 162
rect 480 132 654 152
rect 436 130 654 132
rect 686 130 696 162
rect 436 106 696 130
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 31 295 122 373 0 FreeSans 400 0 0 0 A_N
port 2 nsew
flabel metal1 s 542 440 600 636 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 432 307 518 369 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 192274
string GDS_FILE 6_final.gds
string GDS_START 186666
<< end >>
