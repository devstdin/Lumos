magic
tech ihp-sg13g2
timestamp 1755542813
<< checkpaint >>
rect -1000 -1001 5225 3087
<< poly >>
rect 0 2079 100 2086
rect 0 2063 8 2079
rect 24 2063 42 2079
rect 58 2063 76 2079
rect 92 2063 100 2079
rect 0 2043 100 2063
rect 0 23 100 43
rect 0 7 8 23
rect 24 7 42 23
rect 58 7 76 23
rect 92 7 100 23
rect 0 0 100 7
rect 165 2079 265 2086
rect 165 2063 173 2079
rect 189 2063 207 2079
rect 223 2063 241 2079
rect 257 2063 265 2079
rect 165 2043 265 2063
rect 165 23 265 43
rect 165 7 173 23
rect 189 7 207 23
rect 223 7 241 23
rect 257 7 265 23
rect 165 0 265 7
rect 330 2079 430 2086
rect 330 2063 338 2079
rect 354 2063 372 2079
rect 388 2063 406 2079
rect 422 2063 430 2079
rect 330 2043 430 2063
rect 330 23 430 43
rect 330 7 338 23
rect 354 7 372 23
rect 388 7 406 23
rect 422 7 430 23
rect 330 0 430 7
rect 495 2079 595 2086
rect 495 2063 503 2079
rect 519 2063 537 2079
rect 553 2063 571 2079
rect 587 2063 595 2079
rect 495 2043 595 2063
rect 495 23 595 43
rect 495 7 503 23
rect 519 7 537 23
rect 553 7 571 23
rect 587 7 595 23
rect 495 0 595 7
rect 660 2079 760 2086
rect 660 2063 668 2079
rect 684 2063 702 2079
rect 718 2063 736 2079
rect 752 2063 760 2079
rect 660 2043 760 2063
rect 660 23 760 43
rect 660 7 668 23
rect 684 7 702 23
rect 718 7 736 23
rect 752 7 760 23
rect 660 0 760 7
rect 825 2079 925 2086
rect 825 2063 833 2079
rect 849 2063 867 2079
rect 883 2063 901 2079
rect 917 2063 925 2079
rect 825 2043 925 2063
rect 825 23 925 43
rect 825 7 833 23
rect 849 7 867 23
rect 883 7 901 23
rect 917 7 925 23
rect 825 0 925 7
rect 990 2079 1090 2086
rect 990 2063 998 2079
rect 1014 2063 1032 2079
rect 1048 2063 1066 2079
rect 1082 2063 1090 2079
rect 990 2043 1090 2063
rect 990 23 1090 43
rect 990 7 998 23
rect 1014 7 1032 23
rect 1048 7 1066 23
rect 1082 7 1090 23
rect 990 0 1090 7
rect 1155 2079 1255 2086
rect 1155 2063 1163 2079
rect 1179 2063 1197 2079
rect 1213 2063 1231 2079
rect 1247 2063 1255 2079
rect 1155 2043 1255 2063
rect 1155 23 1255 43
rect 1155 7 1163 23
rect 1179 7 1197 23
rect 1213 7 1231 23
rect 1247 7 1255 23
rect 1155 0 1255 7
rect 1320 2079 1420 2086
rect 1320 2063 1328 2079
rect 1344 2063 1362 2079
rect 1378 2063 1396 2079
rect 1412 2063 1420 2079
rect 1320 2043 1420 2063
rect 1320 23 1420 43
rect 1320 7 1328 23
rect 1344 7 1362 23
rect 1378 7 1396 23
rect 1412 7 1420 23
rect 1320 0 1420 7
rect 1485 2079 1585 2086
rect 1485 2063 1493 2079
rect 1509 2063 1527 2079
rect 1543 2063 1561 2079
rect 1577 2063 1585 2079
rect 1485 2043 1585 2063
rect 1485 23 1585 43
rect 1485 7 1493 23
rect 1509 7 1527 23
rect 1543 7 1561 23
rect 1577 7 1585 23
rect 1485 0 1585 7
rect 1650 2079 1750 2086
rect 1650 2063 1658 2079
rect 1674 2063 1692 2079
rect 1708 2063 1726 2079
rect 1742 2063 1750 2079
rect 1650 2043 1750 2063
rect 1650 23 1750 43
rect 1650 7 1658 23
rect 1674 7 1692 23
rect 1708 7 1726 23
rect 1742 7 1750 23
rect 1650 0 1750 7
rect 1815 2079 1915 2086
rect 1815 2063 1823 2079
rect 1839 2063 1857 2079
rect 1873 2063 1891 2079
rect 1907 2063 1915 2079
rect 1815 2043 1915 2063
rect 1815 23 1915 43
rect 1815 7 1823 23
rect 1839 7 1857 23
rect 1873 7 1891 23
rect 1907 7 1915 23
rect 1815 0 1915 7
rect 1980 2079 2080 2086
rect 1980 2063 1988 2079
rect 2004 2063 2022 2079
rect 2038 2063 2056 2079
rect 2072 2063 2080 2079
rect 1980 2043 2080 2063
rect 1980 23 2080 43
rect 1980 7 1988 23
rect 2004 7 2022 23
rect 2038 7 2056 23
rect 2072 7 2080 23
rect 1980 0 2080 7
rect 2145 2079 2245 2086
rect 2145 2063 2153 2079
rect 2169 2063 2187 2079
rect 2203 2063 2221 2079
rect 2237 2063 2245 2079
rect 2145 2043 2245 2063
rect 2145 23 2245 43
rect 2145 7 2153 23
rect 2169 7 2187 23
rect 2203 7 2221 23
rect 2237 7 2245 23
rect 2145 0 2245 7
rect 2310 2079 2410 2086
rect 2310 2063 2318 2079
rect 2334 2063 2352 2079
rect 2368 2063 2386 2079
rect 2402 2063 2410 2079
rect 2310 2043 2410 2063
rect 2310 23 2410 43
rect 2310 7 2318 23
rect 2334 7 2352 23
rect 2368 7 2386 23
rect 2402 7 2410 23
rect 2310 0 2410 7
rect 2475 2079 2575 2086
rect 2475 2063 2483 2079
rect 2499 2063 2517 2079
rect 2533 2063 2551 2079
rect 2567 2063 2575 2079
rect 2475 2043 2575 2063
rect 2475 23 2575 43
rect 2475 7 2483 23
rect 2499 7 2517 23
rect 2533 7 2551 23
rect 2567 7 2575 23
rect 2475 0 2575 7
rect 2640 2079 2740 2086
rect 2640 2063 2648 2079
rect 2664 2063 2682 2079
rect 2698 2063 2716 2079
rect 2732 2063 2740 2079
rect 2640 2043 2740 2063
rect 2640 23 2740 43
rect 2640 7 2648 23
rect 2664 7 2682 23
rect 2698 7 2716 23
rect 2732 7 2740 23
rect 2640 0 2740 7
rect 2805 2079 2905 2086
rect 2805 2063 2813 2079
rect 2829 2063 2847 2079
rect 2863 2063 2881 2079
rect 2897 2063 2905 2079
rect 2805 2043 2905 2063
rect 2805 23 2905 43
rect 2805 7 2813 23
rect 2829 7 2847 23
rect 2863 7 2881 23
rect 2897 7 2905 23
rect 2805 0 2905 7
rect 2970 2079 3070 2086
rect 2970 2063 2978 2079
rect 2994 2063 3012 2079
rect 3028 2063 3046 2079
rect 3062 2063 3070 2079
rect 2970 2043 3070 2063
rect 2970 23 3070 43
rect 2970 7 2978 23
rect 2994 7 3012 23
rect 3028 7 3046 23
rect 3062 7 3070 23
rect 2970 0 3070 7
rect 3135 2079 3235 2086
rect 3135 2063 3143 2079
rect 3159 2063 3177 2079
rect 3193 2063 3211 2079
rect 3227 2063 3235 2079
rect 3135 2043 3235 2063
rect 3135 23 3235 43
rect 3135 7 3143 23
rect 3159 7 3177 23
rect 3193 7 3211 23
rect 3227 7 3235 23
rect 3135 0 3235 7
rect 3300 2079 3400 2086
rect 3300 2063 3308 2079
rect 3324 2063 3342 2079
rect 3358 2063 3376 2079
rect 3392 2063 3400 2079
rect 3300 2043 3400 2063
rect 3300 23 3400 43
rect 3300 7 3308 23
rect 3324 7 3342 23
rect 3358 7 3376 23
rect 3392 7 3400 23
rect 3300 0 3400 7
rect 3465 2079 3565 2086
rect 3465 2063 3473 2079
rect 3489 2063 3507 2079
rect 3523 2063 3541 2079
rect 3557 2063 3565 2079
rect 3465 2043 3565 2063
rect 3465 23 3565 43
rect 3465 7 3473 23
rect 3489 7 3507 23
rect 3523 7 3541 23
rect 3557 7 3565 23
rect 3465 0 3565 7
rect 3630 2079 3730 2086
rect 3630 2063 3638 2079
rect 3654 2063 3672 2079
rect 3688 2063 3706 2079
rect 3722 2063 3730 2079
rect 3630 2043 3730 2063
rect 3630 23 3730 43
rect 3630 7 3638 23
rect 3654 7 3672 23
rect 3688 7 3706 23
rect 3722 7 3730 23
rect 3630 0 3730 7
rect 3795 2079 3895 2086
rect 3795 2063 3803 2079
rect 3819 2063 3837 2079
rect 3853 2063 3871 2079
rect 3887 2063 3895 2079
rect 3795 2043 3895 2063
rect 3795 23 3895 43
rect 3795 7 3803 23
rect 3819 7 3837 23
rect 3853 7 3871 23
rect 3887 7 3895 23
rect 3795 0 3895 7
rect 3960 2079 4060 2086
rect 3960 2063 3968 2079
rect 3984 2063 4002 2079
rect 4018 2063 4036 2079
rect 4052 2063 4060 2079
rect 3960 2043 4060 2063
rect 3960 23 4060 43
rect 3960 7 3968 23
rect 3984 7 4002 23
rect 4018 7 4036 23
rect 4052 7 4060 23
rect 3960 0 4060 7
rect 4125 2079 4225 2086
rect 4125 2063 4133 2079
rect 4149 2063 4167 2079
rect 4183 2063 4201 2079
rect 4217 2063 4225 2079
rect 4125 2043 4225 2063
rect 4125 23 4225 43
rect 4125 7 4133 23
rect 4149 7 4167 23
rect 4183 7 4201 23
rect 4217 7 4225 23
rect 4125 0 4225 7
<< polycont >>
rect 8 2063 24 2079
rect 42 2063 58 2079
rect 76 2063 92 2079
rect 8 7 24 23
rect 42 7 58 23
rect 76 7 92 23
rect 173 2063 189 2079
rect 207 2063 223 2079
rect 241 2063 257 2079
rect 173 7 189 23
rect 207 7 223 23
rect 241 7 257 23
rect 338 2063 354 2079
rect 372 2063 388 2079
rect 406 2063 422 2079
rect 338 7 354 23
rect 372 7 388 23
rect 406 7 422 23
rect 503 2063 519 2079
rect 537 2063 553 2079
rect 571 2063 587 2079
rect 503 7 519 23
rect 537 7 553 23
rect 571 7 587 23
rect 668 2063 684 2079
rect 702 2063 718 2079
rect 736 2063 752 2079
rect 668 7 684 23
rect 702 7 718 23
rect 736 7 752 23
rect 833 2063 849 2079
rect 867 2063 883 2079
rect 901 2063 917 2079
rect 833 7 849 23
rect 867 7 883 23
rect 901 7 917 23
rect 998 2063 1014 2079
rect 1032 2063 1048 2079
rect 1066 2063 1082 2079
rect 998 7 1014 23
rect 1032 7 1048 23
rect 1066 7 1082 23
rect 1163 2063 1179 2079
rect 1197 2063 1213 2079
rect 1231 2063 1247 2079
rect 1163 7 1179 23
rect 1197 7 1213 23
rect 1231 7 1247 23
rect 1328 2063 1344 2079
rect 1362 2063 1378 2079
rect 1396 2063 1412 2079
rect 1328 7 1344 23
rect 1362 7 1378 23
rect 1396 7 1412 23
rect 1493 2063 1509 2079
rect 1527 2063 1543 2079
rect 1561 2063 1577 2079
rect 1493 7 1509 23
rect 1527 7 1543 23
rect 1561 7 1577 23
rect 1658 2063 1674 2079
rect 1692 2063 1708 2079
rect 1726 2063 1742 2079
rect 1658 7 1674 23
rect 1692 7 1708 23
rect 1726 7 1742 23
rect 1823 2063 1839 2079
rect 1857 2063 1873 2079
rect 1891 2063 1907 2079
rect 1823 7 1839 23
rect 1857 7 1873 23
rect 1891 7 1907 23
rect 1988 2063 2004 2079
rect 2022 2063 2038 2079
rect 2056 2063 2072 2079
rect 1988 7 2004 23
rect 2022 7 2038 23
rect 2056 7 2072 23
rect 2153 2063 2169 2079
rect 2187 2063 2203 2079
rect 2221 2063 2237 2079
rect 2153 7 2169 23
rect 2187 7 2203 23
rect 2221 7 2237 23
rect 2318 2063 2334 2079
rect 2352 2063 2368 2079
rect 2386 2063 2402 2079
rect 2318 7 2334 23
rect 2352 7 2368 23
rect 2386 7 2402 23
rect 2483 2063 2499 2079
rect 2517 2063 2533 2079
rect 2551 2063 2567 2079
rect 2483 7 2499 23
rect 2517 7 2533 23
rect 2551 7 2567 23
rect 2648 2063 2664 2079
rect 2682 2063 2698 2079
rect 2716 2063 2732 2079
rect 2648 7 2664 23
rect 2682 7 2698 23
rect 2716 7 2732 23
rect 2813 2063 2829 2079
rect 2847 2063 2863 2079
rect 2881 2063 2897 2079
rect 2813 7 2829 23
rect 2847 7 2863 23
rect 2881 7 2897 23
rect 2978 2063 2994 2079
rect 3012 2063 3028 2079
rect 3046 2063 3062 2079
rect 2978 7 2994 23
rect 3012 7 3028 23
rect 3046 7 3062 23
rect 3143 2063 3159 2079
rect 3177 2063 3193 2079
rect 3211 2063 3227 2079
rect 3143 7 3159 23
rect 3177 7 3193 23
rect 3211 7 3227 23
rect 3308 2063 3324 2079
rect 3342 2063 3358 2079
rect 3376 2063 3392 2079
rect 3308 7 3324 23
rect 3342 7 3358 23
rect 3376 7 3392 23
rect 3473 2063 3489 2079
rect 3507 2063 3523 2079
rect 3541 2063 3557 2079
rect 3473 7 3489 23
rect 3507 7 3523 23
rect 3541 7 3557 23
rect 3638 2063 3654 2079
rect 3672 2063 3688 2079
rect 3706 2063 3722 2079
rect 3638 7 3654 23
rect 3672 7 3688 23
rect 3706 7 3722 23
rect 3803 2063 3819 2079
rect 3837 2063 3853 2079
rect 3871 2063 3887 2079
rect 3803 7 3819 23
rect 3837 7 3853 23
rect 3871 7 3887 23
rect 3968 2063 3984 2079
rect 4002 2063 4018 2079
rect 4036 2063 4052 2079
rect 3968 7 3984 23
rect 4002 7 4018 23
rect 4036 7 4052 23
rect 4133 2063 4149 2079
rect 4167 2063 4183 2079
rect 4201 2063 4217 2079
rect 4133 7 4149 23
rect 4167 7 4183 23
rect 4201 7 4217 23
<< ppolyres >>
rect 0 43 100 2043
rect 165 43 265 2043
rect 330 43 430 2043
rect 495 43 595 2043
rect 660 43 760 2043
rect 825 43 925 2043
rect 990 43 1090 2043
rect 1155 43 1255 2043
rect 1320 43 1420 2043
rect 1485 43 1585 2043
rect 1650 43 1750 2043
rect 1815 43 1915 2043
rect 1980 43 2080 2043
rect 2145 43 2245 2043
rect 2310 43 2410 2043
rect 2475 43 2575 2043
rect 2640 43 2740 2043
rect 2805 43 2905 2043
rect 2970 43 3070 2043
rect 3135 43 3235 2043
rect 3300 43 3400 2043
rect 3465 43 3565 2043
rect 3630 43 3730 2043
rect 3795 43 3895 2043
rect 3960 43 4060 2043
rect 4125 43 4225 2043
<< metal1 >>
rect 8 2079 257 2087
rect 24 2063 42 2079
rect 58 2063 76 2079
rect 92 2063 173 2079
rect 189 2063 207 2079
rect 223 2063 241 2079
rect 8 2055 257 2063
rect 338 2079 587 2087
rect 354 2063 372 2079
rect 388 2063 406 2079
rect 422 2063 503 2079
rect 519 2063 537 2079
rect 553 2063 571 2079
rect 338 2055 587 2063
rect 668 2079 917 2087
rect 684 2063 702 2079
rect 718 2063 736 2079
rect 752 2063 833 2079
rect 849 2063 867 2079
rect 883 2063 901 2079
rect 668 2055 917 2063
rect 998 2079 1247 2087
rect 1014 2063 1032 2079
rect 1048 2063 1066 2079
rect 1082 2063 1163 2079
rect 1179 2063 1197 2079
rect 1213 2063 1231 2079
rect 998 2055 1247 2063
rect 1328 2079 1577 2087
rect 1344 2063 1362 2079
rect 1378 2063 1396 2079
rect 1412 2063 1493 2079
rect 1509 2063 1527 2079
rect 1543 2063 1561 2079
rect 1328 2055 1577 2063
rect 1658 2079 1907 2087
rect 1674 2063 1692 2079
rect 1708 2063 1726 2079
rect 1742 2063 1823 2079
rect 1839 2063 1857 2079
rect 1873 2063 1891 2079
rect 1658 2055 1907 2063
rect 1988 2079 2237 2087
rect 2004 2063 2022 2079
rect 2038 2063 2056 2079
rect 2072 2063 2153 2079
rect 2169 2063 2187 2079
rect 2203 2063 2221 2079
rect 1988 2055 2237 2063
rect 2318 2079 2567 2087
rect 2334 2063 2352 2079
rect 2368 2063 2386 2079
rect 2402 2063 2483 2079
rect 2499 2063 2517 2079
rect 2533 2063 2551 2079
rect 2318 2055 2567 2063
rect 2648 2079 2897 2087
rect 2664 2063 2682 2079
rect 2698 2063 2716 2079
rect 2732 2063 2813 2079
rect 2829 2063 2847 2079
rect 2863 2063 2881 2079
rect 2648 2055 2897 2063
rect 2978 2079 3227 2087
rect 2994 2063 3012 2079
rect 3028 2063 3046 2079
rect 3062 2063 3143 2079
rect 3159 2063 3177 2079
rect 3193 2063 3211 2079
rect 2978 2055 3227 2063
rect 3308 2079 3557 2087
rect 3324 2063 3342 2079
rect 3358 2063 3376 2079
rect 3392 2063 3473 2079
rect 3489 2063 3507 2079
rect 3523 2063 3541 2079
rect 3308 2055 3557 2063
rect 3638 2079 3887 2087
rect 3654 2063 3672 2079
rect 3688 2063 3706 2079
rect 3722 2063 3803 2079
rect 3819 2063 3837 2079
rect 3853 2063 3871 2079
rect 3638 2055 3887 2063
rect 3968 2079 4217 2087
rect 3984 2063 4002 2079
rect 4018 2063 4036 2079
rect 4052 2063 4133 2079
rect 4149 2063 4167 2079
rect 4183 2063 4201 2079
rect 3968 2055 4217 2063
rect 8 23 92 31
rect 24 7 42 23
rect 58 7 76 23
rect 8 -1 92 7
rect 173 23 422 31
rect 189 7 207 23
rect 223 7 241 23
rect 257 7 338 23
rect 354 7 372 23
rect 388 7 406 23
rect 173 -1 422 7
rect 503 23 752 31
rect 519 7 537 23
rect 553 7 571 23
rect 587 7 668 23
rect 684 7 702 23
rect 718 7 736 23
rect 503 -1 752 7
rect 833 23 1082 31
rect 849 7 867 23
rect 883 7 901 23
rect 917 7 998 23
rect 1014 7 1032 23
rect 1048 7 1066 23
rect 833 -1 1082 7
rect 1163 23 1412 31
rect 1179 7 1197 23
rect 1213 7 1231 23
rect 1247 7 1328 23
rect 1344 7 1362 23
rect 1378 7 1396 23
rect 1163 -1 1412 7
rect 1493 23 1742 31
rect 1509 7 1527 23
rect 1543 7 1561 23
rect 1577 7 1658 23
rect 1674 7 1692 23
rect 1708 7 1726 23
rect 1493 -1 1742 7
rect 1823 23 2072 31
rect 1839 7 1857 23
rect 1873 7 1891 23
rect 1907 7 1988 23
rect 2004 7 2022 23
rect 2038 7 2056 23
rect 1823 -1 2072 7
rect 2153 23 2402 31
rect 2169 7 2187 23
rect 2203 7 2221 23
rect 2237 7 2318 23
rect 2334 7 2352 23
rect 2368 7 2386 23
rect 2153 -1 2402 7
rect 2483 23 2732 31
rect 2499 7 2517 23
rect 2533 7 2551 23
rect 2567 7 2648 23
rect 2664 7 2682 23
rect 2698 7 2716 23
rect 2483 -1 2732 7
rect 2813 23 3062 31
rect 2829 7 2847 23
rect 2863 7 2881 23
rect 2897 7 2978 23
rect 2994 7 3012 23
rect 3028 7 3046 23
rect 2813 -1 3062 7
rect 3143 23 3392 31
rect 3159 7 3177 23
rect 3193 7 3211 23
rect 3227 7 3308 23
rect 3324 7 3342 23
rect 3358 7 3376 23
rect 3143 -1 3392 7
rect 3473 23 3722 31
rect 3489 7 3507 23
rect 3523 7 3541 23
rect 3557 7 3638 23
rect 3654 7 3672 23
rect 3688 7 3706 23
rect 3473 -1 3722 7
rect 3803 23 4052 31
rect 3819 7 3837 23
rect 3853 7 3871 23
rect 3887 7 3968 23
rect 3984 7 4002 23
rect 4018 7 4036 23
rect 3803 -1 4052 7
rect 4133 23 4217 31
rect 4149 7 4167 23
rect 4183 7 4201 23
rect 4133 -1 4217 7
<< labels >>
rlabel comment s 3350 1043 3350 1043 4 rppd r=7.938k
rlabel comment s 710 1043 710 1043 4 rppd r=7.938k
rlabel comment s 3680 1043 3680 1043 4 rppd r=7.938k
rlabel comment s 1040 1043 1040 1043 4 rppd r=7.938k
rlabel comment s 3020 1043 3020 1043 4 rppd r=7.938k
rlabel comment s 50 1043 50 1043 4 rppd r=7.938k
rlabel comment s 2855 1043 2855 1043 4 rppd r=7.938k
rlabel comment s 380 1043 380 1043 4 rppd r=7.938k
rlabel comment s 2030 1043 2030 1043 4 rppd r=7.938k
rlabel comment s 2195 1043 2195 1043 4 rppd r=7.938k
rlabel comment s 2360 1043 2360 1043 4 rppd r=7.938k
rlabel comment s 3185 1043 3185 1043 4 rppd r=7.938k
rlabel comment s 1205 1043 1205 1043 4 rppd r=7.938k
rlabel comment s 875 1043 875 1043 4 rppd r=7.938k
rlabel comment s 3515 1043 3515 1043 4 rppd r=7.938k
rlabel comment s 3845 1043 3845 1043 4 rppd r=7.938k
rlabel comment s 4175 1043 4175 1043 4 rppd r=7.938k
rlabel comment s 215 1043 215 1043 4 rppd r=7.938k
rlabel comment s 1700 1043 1700 1043 4 rppd r=7.938k
rlabel comment s 1535 1043 1535 1043 4 rppd r=7.938k
rlabel comment s 4010 1043 4010 1043 4 rppd r=7.938k
rlabel comment s 2525 1043 2525 1043 4 rppd r=7.938k
rlabel comment s 1370 1043 1370 1043 4 rppd r=7.938k
rlabel comment s 1865 1043 1865 1043 4 rppd r=7.938k
rlabel comment s 2690 1043 2690 1043 4 rppd r=7.938k
rlabel comment s 545 1043 545 1043 4 rppd r=7.938k
rlabel metal1 s 4133 -1 4217 31 4 pin2
port 2 nsew
rlabel metal1 s 8 -1 92 31 4 pin1
port 1 nsew
<< properties >>
string device primitive
string GDS_END 548860
string GDS_FILE sg13g2_io.gds
string GDS_START 533780
<< end >>
