magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757523409
<< error_p >>
rect -67745 131856 135535 132116
rect -67745 131276 -67485 131856
rect -68585 131016 -67485 131276
rect -67453 131564 135243 131824
rect -68585 130436 -68325 131016
rect -67453 130984 -67193 131564
rect -69425 130176 -68325 130436
rect -68293 130724 -67193 130984
rect 134983 130984 135243 131564
rect 135275 131276 135535 131856
rect 135275 131016 136375 131276
rect 134983 130724 136083 130984
rect -69425 129596 -69165 130176
rect -68293 130144 -68033 130724
rect -70265 129336 -69165 129596
rect -69133 129884 -68033 130144
rect 135823 130144 136083 130724
rect 136115 130436 136375 131016
rect 136115 130176 137215 130436
rect 135823 129884 136923 130144
rect -70265 128756 -70005 129336
rect -69133 129304 -68873 129884
rect -71105 128496 -70005 128756
rect -69973 129044 -68873 129304
rect 136663 129304 136923 129884
rect 136955 129596 137215 130176
rect 136955 129336 138055 129596
rect 136663 129044 137763 129304
rect -71105 -58264 -70845 128496
rect -69973 128464 -69713 129044
rect -70813 128204 -69713 128464
rect 137503 128464 137763 129044
rect 137795 128756 138055 129336
rect 137795 128496 138895 128756
rect 137503 128204 138603 128464
rect -70813 -57972 -70553 128204
rect 138343 -57972 138603 128204
rect -70813 -58232 -69713 -57972
rect -71105 -58524 -70005 -58264
rect -70265 -59104 -70005 -58524
rect -69973 -58812 -69713 -58232
rect 137503 -58232 138603 -57972
rect 137503 -58812 137763 -58232
rect 138635 -58264 138895 128496
rect -69973 -59072 -68873 -58812
rect -70265 -59364 -69165 -59104
rect -69425 -59944 -69165 -59364
rect -69133 -59652 -68873 -59072
rect 136663 -59072 137763 -58812
rect 137795 -58524 138895 -58264
rect 136663 -59652 136923 -59072
rect 137795 -59104 138055 -58524
rect -69133 -59912 -68033 -59652
rect -69425 -60204 -68325 -59944
rect -68585 -60784 -68325 -60204
rect -68293 -60492 -68033 -59912
rect 135823 -59912 136923 -59652
rect 136955 -59364 138055 -59104
rect 135823 -60492 136083 -59912
rect 136955 -59944 137215 -59364
rect -68293 -60752 -67193 -60492
rect -68585 -61044 -67485 -60784
rect -67745 -61624 -67485 -61044
rect -67453 -61332 -67193 -60752
rect 134983 -60752 136083 -60492
rect 136115 -60204 137215 -59944
rect 134983 -61332 135243 -60752
rect 136115 -60784 136375 -60204
rect -67453 -61592 135243 -61332
rect 135275 -61044 136375 -60784
rect 135275 -61624 135535 -61044
rect -67745 -61884 135535 -61624
<< error_s >>
rect 103320 -22834 104381 -21414
rect 99075 -27884 99524 -26065
<< metal1 >>
rect -13105 125216 895 125217
rect 79078 60362 81602 60462
rect 79078 60062 79178 60362
rect 81502 60062 81602 60362
rect 79078 59651 81602 60062
rect 79191 59505 79310 59515
rect 79191 59333 79201 59505
rect 79300 59333 79310 59505
rect 79191 59323 79310 59333
rect 81370 59505 81489 59515
rect 81370 59333 81380 59505
rect 81479 59333 81489 59505
rect 81370 59323 81489 59333
rect 76856 56581 78306 56591
rect 76856 56201 77898 56581
rect 78296 56201 78306 56581
rect 76856 56191 78306 56201
rect 76844 55881 79502 55891
rect 76844 55501 79094 55881
rect 79492 55501 79502 55881
rect 76844 55491 79502 55501
rect -5432 -2570 -5032 -977
rect -5432 -2968 -5422 -2570
rect -5042 -2968 -5032 -2570
rect -5432 -2978 -5032 -2968
rect 6796 -2392 7596 -577
rect 6796 -2402 13997 -2392
rect 6796 -3182 13207 -2402
rect 13987 -3182 13997 -2402
rect 6796 -3192 13997 -3182
<< via1 >>
rect 79178 60062 81502 60362
rect 79201 59333 79300 59505
rect 81380 59333 81479 59505
rect 77898 56201 78296 56581
rect 79094 55501 79492 55881
rect -5422 -2968 -5042 -2570
rect 13207 -3182 13987 -2402
<< metal2 >>
rect -13105 125216 895 125217
rect 26895 74716 30589 79602
rect 30991 74716 34685 79602
rect 35085 74716 38779 79600
rect 26895 73816 38779 74716
rect 26895 72016 26995 73816
rect 38679 72016 38779 73816
rect 73524 72971 74266 75230
rect 26895 71916 38779 72016
rect 71788 72229 74266 72971
rect 71788 70944 72530 72229
rect 77888 66902 82133 67320
rect 77888 56581 78306 66902
rect 79078 60362 81602 60462
rect 79078 60062 79178 60362
rect 81502 60062 81602 60362
rect 79078 59962 81602 60062
rect 78580 59515 78972 59615
rect 78580 59323 78680 59515
rect 78872 59505 79310 59515
rect 78872 59333 79201 59505
rect 79300 59333 79310 59505
rect 78872 59323 79310 59333
rect 81370 59505 81489 59515
rect 81370 59333 81380 59505
rect 81479 59450 81489 59505
rect 81479 59392 81953 59450
rect 81479 59333 81489 59392
rect 81370 59323 81489 59333
rect 78580 59223 78972 59323
rect 77888 56201 77898 56581
rect 78296 56201 78306 56581
rect 77888 56191 78306 56201
rect 79084 58602 82133 59020
rect 79084 55881 79502 58602
rect 79084 55501 79094 55881
rect 79492 55501 79502 55881
rect 79084 55491 79502 55501
rect 77664 42909 81969 43309
rect 77664 41183 78064 42909
rect 77664 40172 81064 40572
rect 77664 39175 80064 39575
rect 77664 38173 79064 38573
rect -18582 27900 -10905 28000
rect -18582 24306 -12805 27900
rect -13705 23906 -12805 24306
rect -18583 20212 -12805 23906
rect -13705 19810 -12805 20212
rect -18582 16216 -12805 19810
rect -11005 16216 -10905 27900
rect -18582 16116 -10905 16216
rect 44922 -1733 47089 -1210
rect 77664 -1614 78064 37562
rect 13197 -2402 13997 -2392
rect -5432 -2570 -2375 -2560
rect -5432 -2968 -5422 -2570
rect -5042 -2968 -2375 -2570
rect -5432 -2978 -2375 -2968
rect -2793 -4942 -2375 -2978
rect 13197 -3182 13207 -2402
rect 13987 -3182 13997 -2402
rect 13197 -4998 13997 -3182
rect 32499 -3900 47089 -1733
rect 74172 -1624 78064 -1614
rect 74172 -2004 74182 -1624
rect 74580 -2004 78064 -1624
rect 74172 -2014 78064 -2004
rect 78664 -2902 79064 38173
rect 79664 3311 80064 39175
rect 80664 23310 81064 40172
rect 80664 22910 81963 23310
rect 79664 2911 81965 3311
rect 73202 -2912 79064 -2902
rect 73202 -3292 73212 -2912
rect 73610 -3292 79064 -2912
rect 73202 -3302 79064 -3292
rect 32499 -5017 34666 -3900
<< via2 >>
rect 26995 72016 38679 73816
rect 79178 60062 81502 60362
rect 78680 59323 78872 59515
rect -12805 16216 -11005 27900
rect 74182 -2004 74580 -1624
rect 73212 -3292 73610 -2912
<< metal3 >>
rect -13105 125216 895 125217
rect 26895 73816 38779 73916
rect 26895 72016 26995 73816
rect 38679 72016 38779 73816
rect 26895 71916 38779 72016
rect 79078 60362 81602 60462
rect 79078 60062 79178 60362
rect 81502 60062 81602 60362
rect 79078 59962 81602 60062
rect 78580 59515 78972 59615
rect 78580 59323 78680 59515
rect 78872 59323 78972 59515
rect 78580 59223 78972 59323
rect -12905 27900 -10905 28000
rect -12905 16216 -12805 27900
rect -11005 16216 -10905 27900
rect -12905 16116 -10905 16216
rect -12905 9516 -7905 9616
rect -12905 -3284 -12805 9516
rect -11005 5641 -7905 9516
rect -11005 5244 -10891 5641
rect -8914 5244 -7905 5641
rect -11005 991 -7905 5244
rect -11005 594 -10891 991
rect -8914 594 -7905 991
rect -11005 -3284 -7905 594
rect 74172 -1624 74590 -1614
rect 74172 -2004 74182 -1624
rect 74580 -2004 74590 -1624
rect -12905 -3384 -7905 -3284
rect 73202 -2912 73620 -2902
rect 73202 -3292 73212 -2912
rect 73610 -3292 73620 -2912
rect 73202 -4942 73620 -3292
rect 74172 -4942 74590 -2004
<< via3 >>
rect 26995 72016 38679 73816
rect 79178 60062 81502 60362
rect 78680 59323 78872 59515
rect -12805 16216 -11005 27900
rect -12805 -3284 -11005 9516
<< metal4 >>
rect -13105 125216 895 125217
rect 26895 73816 38779 73916
rect 26895 72016 26995 73816
rect 38679 72016 38779 73816
rect 26895 71916 38779 72016
rect 79078 60362 81602 60462
rect 79078 60062 79178 60362
rect 81502 60062 81602 60362
rect 79078 59962 81602 60062
rect 78580 59515 78972 59615
rect 78580 59323 78680 59515
rect 78872 59323 78972 59515
rect 78580 59223 78972 59323
rect -12905 27900 -7905 28000
rect -12905 16216 -12805 27900
rect -11005 24306 -7905 27900
rect -11005 23908 -10889 24306
rect -8911 23908 -7905 24306
rect -11005 20212 -7905 23908
rect -11005 19814 -10889 20212
rect -8911 19814 -7905 20212
rect -11005 16216 -7905 19814
rect -12905 16116 -7905 16216
rect -12905 9516 -10905 9616
rect -12905 -3284 -12805 9516
rect -11005 -3284 -10905 9516
rect -12905 -3384 -10905 -3284
<< via4 >>
rect 26995 72016 38679 73816
rect 79178 60062 81502 60362
rect 78680 59323 78872 59515
rect -12805 -3284 -11005 9516
<< metal5 >>
rect -13105 125216 895 125217
rect 26895 73816 38779 73916
rect 26895 72016 26995 73816
rect 38679 72016 38779 73816
rect 26895 71916 38779 72016
rect 47395 73816 60395 73916
rect 47395 72016 47495 73816
rect 60295 72016 60395 73816
rect 47395 71895 60395 72016
rect 47395 70837 51025 71895
rect 52025 70837 55698 71895
rect 56698 70837 60395 71895
rect 47395 69916 60395 70837
rect 79078 60362 81602 60462
rect 79078 60062 79178 60362
rect 81502 60062 81602 60362
rect 79078 59962 81602 60062
rect 75580 59515 78972 59615
rect 75580 59323 78680 59515
rect 78872 59323 78972 59515
rect 75580 59223 78972 59323
rect -12905 9516 -10905 9616
rect -12905 -3284 -12805 9516
rect -11005 -3284 -10905 9516
rect -12905 -3384 -10905 -3284
<< via5 >>
rect 26995 72016 38679 73816
rect 47495 72016 60295 73816
rect 79178 60062 81502 60362
rect -12805 -3284 -11005 9516
<< metal6 >>
rect -13105 125216 895 125217
rect 26895 73816 38779 73916
rect 26895 72016 26995 73816
rect 38679 72016 38779 73816
rect 26895 71913 38779 72016
rect 47395 73816 60395 73916
rect 47395 72016 47495 73816
rect 60295 72016 60395 73816
rect 47395 71916 60395 72016
rect 26895 70815 30273 71913
rect 31273 70815 34387 71913
rect 35387 70815 38779 71913
rect 26895 69916 38779 70815
rect 75578 60362 81602 60462
rect 75578 60062 79178 60362
rect 81502 60062 81602 60362
rect 75578 59962 81602 60062
rect -12905 9516 -10905 9616
rect -12905 -3284 -12805 9516
rect -11005 -3284 -10905 9516
rect -12905 -3384 -10905 -3284
<< via6 >>
rect 47495 72016 60295 73816
rect -12805 -3284 -11005 9516
<< metal7 >>
rect -13105 125216 895 125416
rect 6895 125216 20895 125416
rect 26895 125216 40895 125416
rect 46895 125216 60895 125416
rect 66895 125216 80895 125416
rect 47395 79790 60395 79874
rect 47395 73946 51025 79790
rect 52025 73946 55705 79790
rect 56705 73946 60395 79790
rect 47395 73816 60395 73946
rect 47395 72016 47495 73816
rect 60295 72016 60395 73816
rect 47395 71916 60395 72016
rect -64405 56116 -64205 70116
rect 131995 56116 132195 70116
rect -64405 36116 -64205 50116
rect 131995 36116 132195 50116
rect -64405 16116 -64205 30116
rect 131995 16116 132195 30116
rect -64405 -3884 -64205 10116
rect -18854 9516 -10905 9616
rect -18854 5944 -12805 9516
rect -18854 4950 -18805 5944
rect -12938 4950 -12805 5944
rect -18854 1279 -12805 4950
rect -18854 285 -18805 1279
rect -12938 285 -12805 1279
rect -18854 -3284 -12805 285
rect -11005 -3284 -10905 9516
rect -18854 -3384 -10905 -3284
rect 131995 -3884 132195 10116
rect -13105 -55184 895 -54984
rect 6895 -55184 20895 -54984
rect 26895 -55184 40895 -54984
rect 66896 -55184 80896 -54984
use core  core_0 .
timestamp 1757454070
transform 1 0 -3548 0 1 4450
box -7353 -5827 81612 68359
use padring  padring_0 .
timestamp 1756924281
transform 1 0 0 0 1 0
box -64405 -55184 132195 125416
use rhigh_NHH9UC  rhigh_NHH9UC_0
timestamp 1757266023
transform 0 1 80340 -1 0 59419
box -280 -1266 280 1266
use sealring  sealring_0 .
timestamp 1756676971
transform 1 0 0 0 1 0
box -72685 -63464 140475 133696
<< labels >>
flabel metal7 -64405 -3884 -64205 10116 0 FreeSans 8000 0 0 0 AVDD
port 0 nsew
flabel metal7 -64405 16116 -64205 30116 0 FreeSans 8000 0 0 0 VSS
port 1 nsew
flabel metal7 -64405 36116 -64205 50116 0 FreeSans 8000 0 0 0 IOAVDD
port 2 nsew
flabel metal7 -64405 56116 -64205 70116 0 FreeSans 8000 0 0 0 IOAVSS
port 3 nsew
flabel metal7 -13105 125216 895 125416 0 FreeSans 8000 0 0 0 IODVSS
port 4 nsew
flabel metal7 6895 125216 20895 125416 0 FreeSans 8000 0 0 0 IODVDD
port 5 nsew
flabel metal7 46895 125216 60895 125416 0 FreeSans 8000 0 0 0 DVDD
port 6 nsew
flabel metal7 66895 125216 80895 125416 0 FreeSans 8000 0 0 0 OSC
port 7 nsew
flabel metal7 131995 56116 132195 70116 0 FreeSans 8000 0 0 0 RESET
port 8 nsew
flabel metal7 131995 36116 132195 50116 0 FreeSans 8000 0 0 0 CS
port 9 nsew
flabel metal7 131995 16116 132195 30116 0 FreeSans 8000 0 0 0 SCLK
port 10 nsew
flabel metal7 131995 -3884 132195 10116 0 FreeSans 8000 0 0 0 DIN
port 11 nsew
flabel metal7 66896 -55184 80896 -54984 0 FreeSans 8000 0 0 0 DOUT
port 12 nsew
flabel metal7 26895 -55184 40895 -54984 0 FreeSans 8000 0 0 0 VLDO
port 13 nsew
flabel metal7 6895 -55184 20895 -54984 0 FreeSans 8000 0 0 0 FTOP
port 14 nsew
flabel metal7 -13105 -55184 895 -54984 0 FreeSans 8000 0 0 0 FPROG
port 15 nsew
<< end >>
