magic
tech ihp-sg13g2
magscale 1 2
timestamp 1749474908
<< metal1 >>
rect 3 16613 1559 17112
rect 1677 3009 2446 3452
rect 1677 2597 1885 3009
rect 2017 2958 2109 2968
rect 2017 2890 2027 2958
rect 2099 2890 2109 2958
rect 2017 2824 2109 2890
rect 208 2508 1885 2597
rect 208 78 577 2508
rect 739 2325 831 2508
rect 875 2325 1103 2377
rect 1147 2325 1375 2377
rect 739 213 967 265
rect 1011 213 1239 265
rect 1283 199 1375 265
rect 1283 136 1293 199
rect 1365 136 1375 199
rect 1283 126 1375 136
rect 1509 78 1885 2508
rect 2241 527 2446 3009
rect 2017 199 2109 264
rect 2017 136 2027 199
rect 2099 136 2109 199
rect 2017 126 2109 136
rect 2241 78 3959 527
rect 208 28 3959 78
<< via1 >>
rect 2027 2890 2099 2958
rect 1293 136 1365 199
rect 2027 136 2099 199
<< metal2 >>
rect 12248 16506 13538 17112
rect 3 6748 427 7176
rect 3 6247 427 6674
rect 3 5096 429 5478
rect 558 2968 758 3044
rect 558 2958 2109 2968
rect 0 2759 430 2957
rect 558 2890 2027 2958
rect 2099 2890 2109 2958
rect 558 2880 2109 2890
rect 0 2676 1729 2759
rect 0 2604 430 2676
rect 1646 209 1729 2676
rect 1283 199 2109 209
rect 1283 136 1293 199
rect 1365 136 2027 199
rect 2099 136 2109 199
rect 1283 126 2109 136
use ldoota  ldoota_0
timestamp 1749471858
transform 1 0 -3160 0 1 15008
box 3161 -15009 33091 2104
use rhigh_BJZ3BW  rhigh_BJZ3BW_0
timestamp 1749470838
transform 1 0 785 0 1 1295
box -230 -1266 774 1266
use rhigh_KA4Q3N  rhigh_KA4Q3N_0
timestamp 1749470838
transform 1 0 2063 0 1 1544
box -230 -1516 230 1516
<< labels >>
flabel metal2 0 2604 430 2957 0 FreeSans 800 0 0 0 FBOUT
port 0 nsew
flabel metal1 2403 28 3959 527 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel metal2 3 5096 429 5478 0 FreeSans 800 0 0 0 IB
port 5 nsew
flabel metal2 3 6247 427 6674 0 FreeSans 800 0 0 0 FBIN
port 7 nsew
flabel metal2 3 6748 427 7176 0 FreeSans 800 0 0 0 VREF
port 8 nsew
flabel metal1 3 16613 1559 17112 0 FreeSans 800 0 0 0 VDD
port 10 nsew
flabel metal2 12248 16506 13538 17112 0 FreeSans 800 0 0 0 VLDO
port 14 nsew
<< end >>
