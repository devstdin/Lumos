magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -924 2524 37600
<< isosubstrate >>
rect 44 23124 356 28034
rect 44 18112 356 22924
rect 44 13000 356 17912
<< nwell >>
rect -124 33246 524 33554
rect -124 29546 524 29854
rect -124 1076 524 12324
<< pwell >>
rect 144 31456 256 31524
rect 18 31344 382 31456
rect 144 31276 256 31344
rect 18 12974 382 28060
<< psubdiff >>
rect 116 31384 148 31416
rect 184 31384 216 31416
rect 252 31384 284 31416
rect 184 31316 216 31348
rect 184 27939 216 27971
rect 256 27939 288 27971
rect 112 27867 144 27899
rect 184 27867 216 27899
rect 256 27867 288 27899
rect 112 27795 144 27827
rect 184 27795 216 27827
rect 256 27795 288 27827
rect 112 27723 144 27755
rect 184 27723 216 27755
rect 256 27723 288 27755
rect 112 27651 144 27683
rect 184 27651 216 27683
rect 256 27651 288 27683
rect 112 27579 144 27611
rect 184 27579 216 27611
rect 256 27579 288 27611
rect 112 27507 144 27539
rect 184 27507 216 27539
rect 256 27507 288 27539
rect 112 27435 144 27467
rect 184 27435 216 27467
rect 256 27435 288 27467
rect 112 27363 144 27395
rect 184 27363 216 27395
rect 256 27363 288 27395
rect 112 27291 144 27323
rect 184 27291 216 27323
rect 256 27291 288 27323
rect 112 27219 144 27251
rect 184 27219 216 27251
rect 256 27219 288 27251
rect 112 27147 144 27179
rect 184 27147 216 27179
rect 256 27147 288 27179
rect 112 27075 144 27107
rect 184 27075 216 27107
rect 256 27075 288 27107
rect 112 27003 144 27035
rect 184 27003 216 27035
rect 256 27003 288 27035
rect 112 26931 144 26963
rect 184 26931 216 26963
rect 256 26931 288 26963
rect 112 26859 144 26891
rect 184 26859 216 26891
rect 256 26859 288 26891
rect 112 26787 144 26819
rect 184 26787 216 26819
rect 256 26787 288 26819
rect 112 26715 144 26747
rect 184 26715 216 26747
rect 256 26715 288 26747
rect 112 26643 144 26675
rect 184 26643 216 26675
rect 256 26643 288 26675
rect 112 26571 144 26603
rect 184 26571 216 26603
rect 256 26571 288 26603
rect 112 26499 144 26531
rect 184 26499 216 26531
rect 256 26499 288 26531
rect 112 26427 144 26459
rect 184 26427 216 26459
rect 256 26427 288 26459
rect 112 26355 144 26387
rect 184 26355 216 26387
rect 256 26355 288 26387
rect 112 26283 144 26315
rect 184 26283 216 26315
rect 256 26283 288 26315
rect 112 26211 144 26243
rect 184 26211 216 26243
rect 256 26211 288 26243
rect 112 26139 144 26171
rect 184 26139 216 26171
rect 256 26139 288 26171
rect 112 26067 144 26099
rect 184 26067 216 26099
rect 256 26067 288 26099
rect 112 25995 144 26027
rect 184 25995 216 26027
rect 256 25995 288 26027
rect 112 25923 144 25955
rect 184 25923 216 25955
rect 256 25923 288 25955
rect 112 25851 144 25883
rect 184 25851 216 25883
rect 256 25851 288 25883
rect 112 25779 144 25811
rect 184 25779 216 25811
rect 256 25779 288 25811
rect 112 25707 144 25739
rect 184 25707 216 25739
rect 256 25707 288 25739
rect 112 25635 144 25667
rect 184 25635 216 25667
rect 256 25635 288 25667
rect 112 25563 144 25595
rect 184 25563 216 25595
rect 256 25563 288 25595
rect 112 25491 144 25523
rect 184 25491 216 25523
rect 256 25491 288 25523
rect 112 25419 144 25451
rect 184 25419 216 25451
rect 256 25419 288 25451
rect 112 25347 144 25379
rect 184 25347 216 25379
rect 256 25347 288 25379
rect 112 25275 144 25307
rect 184 25275 216 25307
rect 256 25275 288 25307
rect 112 25203 144 25235
rect 184 25203 216 25235
rect 256 25203 288 25235
rect 112 25131 144 25163
rect 184 25131 216 25163
rect 256 25131 288 25163
rect 112 25059 144 25091
rect 184 25059 216 25091
rect 256 25059 288 25091
rect 112 24987 144 25019
rect 184 24987 216 25019
rect 256 24987 288 25019
rect 112 24915 144 24947
rect 184 24915 216 24947
rect 256 24915 288 24947
rect 112 24843 144 24875
rect 184 24843 216 24875
rect 256 24843 288 24875
rect 112 24771 144 24803
rect 184 24771 216 24803
rect 256 24771 288 24803
rect 112 24699 144 24731
rect 184 24699 216 24731
rect 256 24699 288 24731
rect 112 24627 144 24659
rect 184 24627 216 24659
rect 256 24627 288 24659
rect 112 24555 144 24587
rect 184 24555 216 24587
rect 256 24555 288 24587
rect 112 24483 144 24515
rect 184 24483 216 24515
rect 256 24483 288 24515
rect 112 24411 144 24443
rect 184 24411 216 24443
rect 256 24411 288 24443
rect 112 24339 144 24371
rect 184 24339 216 24371
rect 256 24339 288 24371
rect 112 24267 144 24299
rect 184 24267 216 24299
rect 256 24267 288 24299
rect 112 24195 144 24227
rect 184 24195 216 24227
rect 256 24195 288 24227
rect 112 24123 144 24155
rect 184 24123 216 24155
rect 256 24123 288 24155
rect 112 24051 144 24083
rect 184 24051 216 24083
rect 256 24051 288 24083
rect 112 23979 144 24011
rect 184 23979 216 24011
rect 256 23979 288 24011
rect 112 23907 144 23939
rect 184 23907 216 23939
rect 256 23907 288 23939
rect 112 23835 144 23867
rect 184 23835 216 23867
rect 256 23835 288 23867
rect 112 23763 144 23795
rect 184 23763 216 23795
rect 256 23763 288 23795
rect 112 23691 144 23723
rect 184 23691 216 23723
rect 256 23691 288 23723
rect 112 23619 144 23651
rect 184 23619 216 23651
rect 256 23619 288 23651
rect 112 23547 144 23579
rect 184 23547 216 23579
rect 256 23547 288 23579
rect 112 23475 144 23507
rect 184 23475 216 23507
rect 256 23475 288 23507
rect 112 23403 144 23435
rect 184 23403 216 23435
rect 256 23403 288 23435
rect 112 23331 144 23363
rect 184 23331 216 23363
rect 256 23331 288 23363
rect 112 23259 144 23291
rect 184 23259 216 23291
rect 256 23259 288 23291
rect 112 23187 144 23219
rect 184 23187 216 23219
rect 256 23187 288 23219
rect 184 22842 216 22874
rect 256 22842 288 22874
rect 112 22770 144 22802
rect 184 22770 216 22802
rect 256 22770 288 22802
rect 112 22698 144 22730
rect 184 22698 216 22730
rect 256 22698 288 22730
rect 112 22626 144 22658
rect 184 22626 216 22658
rect 256 22626 288 22658
rect 112 22554 144 22586
rect 184 22554 216 22586
rect 256 22554 288 22586
rect 112 22482 144 22514
rect 184 22482 216 22514
rect 256 22482 288 22514
rect 112 22410 144 22442
rect 184 22410 216 22442
rect 256 22410 288 22442
rect 112 22338 144 22370
rect 184 22338 216 22370
rect 256 22338 288 22370
rect 112 22266 144 22298
rect 184 22266 216 22298
rect 256 22266 288 22298
rect 112 22194 144 22226
rect 184 22194 216 22226
rect 256 22194 288 22226
rect 112 22122 144 22154
rect 184 22122 216 22154
rect 256 22122 288 22154
rect 112 22050 144 22082
rect 184 22050 216 22082
rect 256 22050 288 22082
rect 112 21978 144 22010
rect 184 21978 216 22010
rect 256 21978 288 22010
rect 112 21906 144 21938
rect 184 21906 216 21938
rect 256 21906 288 21938
rect 112 21834 144 21866
rect 184 21834 216 21866
rect 256 21834 288 21866
rect 112 21762 144 21794
rect 184 21762 216 21794
rect 256 21762 288 21794
rect 112 21690 144 21722
rect 184 21690 216 21722
rect 256 21690 288 21722
rect 112 21618 144 21650
rect 184 21618 216 21650
rect 256 21618 288 21650
rect 112 21546 144 21578
rect 184 21546 216 21578
rect 256 21546 288 21578
rect 112 21474 144 21506
rect 184 21474 216 21506
rect 256 21474 288 21506
rect 112 21402 144 21434
rect 184 21402 216 21434
rect 256 21402 288 21434
rect 112 21330 144 21362
rect 184 21330 216 21362
rect 256 21330 288 21362
rect 112 21258 144 21290
rect 184 21258 216 21290
rect 256 21258 288 21290
rect 112 21186 144 21218
rect 184 21186 216 21218
rect 256 21186 288 21218
rect 112 21114 144 21146
rect 184 21114 216 21146
rect 256 21114 288 21146
rect 112 21042 144 21074
rect 184 21042 216 21074
rect 256 21042 288 21074
rect 112 20970 144 21002
rect 184 20970 216 21002
rect 256 20970 288 21002
rect 112 20898 144 20930
rect 184 20898 216 20930
rect 256 20898 288 20930
rect 112 20826 144 20858
rect 184 20826 216 20858
rect 256 20826 288 20858
rect 112 20754 144 20786
rect 184 20754 216 20786
rect 256 20754 288 20786
rect 112 20682 144 20714
rect 184 20682 216 20714
rect 256 20682 288 20714
rect 112 20610 144 20642
rect 184 20610 216 20642
rect 256 20610 288 20642
rect 112 20538 144 20570
rect 184 20538 216 20570
rect 256 20538 288 20570
rect 112 20466 144 20498
rect 184 20466 216 20498
rect 256 20466 288 20498
rect 112 20394 144 20426
rect 184 20394 216 20426
rect 256 20394 288 20426
rect 112 20322 144 20354
rect 184 20322 216 20354
rect 256 20322 288 20354
rect 112 20250 144 20282
rect 184 20250 216 20282
rect 256 20250 288 20282
rect 112 20178 144 20210
rect 184 20178 216 20210
rect 256 20178 288 20210
rect 112 20106 144 20138
rect 184 20106 216 20138
rect 256 20106 288 20138
rect 112 20034 144 20066
rect 184 20034 216 20066
rect 256 20034 288 20066
rect 112 19962 144 19994
rect 184 19962 216 19994
rect 256 19962 288 19994
rect 112 19890 144 19922
rect 184 19890 216 19922
rect 256 19890 288 19922
rect 112 19818 144 19850
rect 184 19818 216 19850
rect 256 19818 288 19850
rect 112 19746 144 19778
rect 184 19746 216 19778
rect 256 19746 288 19778
rect 112 19674 144 19706
rect 184 19674 216 19706
rect 256 19674 288 19706
rect 112 19602 144 19634
rect 184 19602 216 19634
rect 256 19602 288 19634
rect 112 19530 144 19562
rect 184 19530 216 19562
rect 256 19530 288 19562
rect 112 19458 144 19490
rect 184 19458 216 19490
rect 256 19458 288 19490
rect 112 19386 144 19418
rect 184 19386 216 19418
rect 256 19386 288 19418
rect 112 19314 144 19346
rect 184 19314 216 19346
rect 256 19314 288 19346
rect 112 19242 144 19274
rect 184 19242 216 19274
rect 256 19242 288 19274
rect 112 19170 144 19202
rect 184 19170 216 19202
rect 256 19170 288 19202
rect 112 19098 144 19130
rect 184 19098 216 19130
rect 256 19098 288 19130
rect 112 19026 144 19058
rect 184 19026 216 19058
rect 256 19026 288 19058
rect 112 18954 144 18986
rect 184 18954 216 18986
rect 256 18954 288 18986
rect 112 18882 144 18914
rect 184 18882 216 18914
rect 256 18882 288 18914
rect 112 18810 144 18842
rect 184 18810 216 18842
rect 256 18810 288 18842
rect 112 18738 144 18770
rect 184 18738 216 18770
rect 256 18738 288 18770
rect 112 18666 144 18698
rect 184 18666 216 18698
rect 256 18666 288 18698
rect 112 18594 144 18626
rect 184 18594 216 18626
rect 256 18594 288 18626
rect 112 18522 144 18554
rect 184 18522 216 18554
rect 256 18522 288 18554
rect 112 18450 144 18482
rect 184 18450 216 18482
rect 256 18450 288 18482
rect 112 18378 144 18410
rect 184 18378 216 18410
rect 256 18378 288 18410
rect 112 18306 144 18338
rect 184 18306 216 18338
rect 256 18306 288 18338
rect 112 18234 144 18266
rect 184 18234 216 18266
rect 256 18234 288 18266
rect 112 18162 144 18194
rect 184 18162 216 18194
rect 256 18162 288 18194
rect 184 17816 216 17848
rect 256 17816 288 17848
rect 112 17744 144 17776
rect 184 17744 216 17776
rect 256 17744 288 17776
rect 112 17672 144 17704
rect 184 17672 216 17704
rect 256 17672 288 17704
rect 112 17600 144 17632
rect 184 17600 216 17632
rect 256 17600 288 17632
rect 112 17528 144 17560
rect 184 17528 216 17560
rect 256 17528 288 17560
rect 112 17456 144 17488
rect 184 17456 216 17488
rect 256 17456 288 17488
rect 112 17384 144 17416
rect 184 17384 216 17416
rect 256 17384 288 17416
rect 112 17312 144 17344
rect 184 17312 216 17344
rect 256 17312 288 17344
rect 112 17240 144 17272
rect 184 17240 216 17272
rect 256 17240 288 17272
rect 112 17168 144 17200
rect 184 17168 216 17200
rect 256 17168 288 17200
rect 112 17096 144 17128
rect 184 17096 216 17128
rect 256 17096 288 17128
rect 112 17024 144 17056
rect 184 17024 216 17056
rect 256 17024 288 17056
rect 112 16952 144 16984
rect 184 16952 216 16984
rect 256 16952 288 16984
rect 112 16880 144 16912
rect 184 16880 216 16912
rect 256 16880 288 16912
rect 112 16808 144 16840
rect 184 16808 216 16840
rect 256 16808 288 16840
rect 112 16736 144 16768
rect 184 16736 216 16768
rect 256 16736 288 16768
rect 112 16664 144 16696
rect 184 16664 216 16696
rect 256 16664 288 16696
rect 112 16592 144 16624
rect 184 16592 216 16624
rect 256 16592 288 16624
rect 112 16520 144 16552
rect 184 16520 216 16552
rect 256 16520 288 16552
rect 112 16448 144 16480
rect 184 16448 216 16480
rect 256 16448 288 16480
rect 112 16376 144 16408
rect 184 16376 216 16408
rect 256 16376 288 16408
rect 112 16304 144 16336
rect 184 16304 216 16336
rect 256 16304 288 16336
rect 112 16232 144 16264
rect 184 16232 216 16264
rect 256 16232 288 16264
rect 112 16160 144 16192
rect 184 16160 216 16192
rect 256 16160 288 16192
rect 112 16088 144 16120
rect 184 16088 216 16120
rect 256 16088 288 16120
rect 112 16016 144 16048
rect 184 16016 216 16048
rect 256 16016 288 16048
rect 112 15944 144 15976
rect 184 15944 216 15976
rect 256 15944 288 15976
rect 112 15872 144 15904
rect 184 15872 216 15904
rect 256 15872 288 15904
rect 112 15800 144 15832
rect 184 15800 216 15832
rect 256 15800 288 15832
rect 112 15728 144 15760
rect 184 15728 216 15760
rect 256 15728 288 15760
rect 112 15656 144 15688
rect 184 15656 216 15688
rect 256 15656 288 15688
rect 112 15584 144 15616
rect 184 15584 216 15616
rect 256 15584 288 15616
rect 112 15512 144 15544
rect 184 15512 216 15544
rect 256 15512 288 15544
rect 112 15440 144 15472
rect 184 15440 216 15472
rect 256 15440 288 15472
rect 112 15368 144 15400
rect 184 15368 216 15400
rect 256 15368 288 15400
rect 112 15296 144 15328
rect 184 15296 216 15328
rect 256 15296 288 15328
rect 112 15224 144 15256
rect 184 15224 216 15256
rect 256 15224 288 15256
rect 112 15152 144 15184
rect 184 15152 216 15184
rect 256 15152 288 15184
rect 112 15080 144 15112
rect 184 15080 216 15112
rect 256 15080 288 15112
rect 112 15008 144 15040
rect 184 15008 216 15040
rect 256 15008 288 15040
rect 112 14936 144 14968
rect 184 14936 216 14968
rect 256 14936 288 14968
rect 112 14864 144 14896
rect 184 14864 216 14896
rect 256 14864 288 14896
rect 112 14792 144 14824
rect 184 14792 216 14824
rect 256 14792 288 14824
rect 112 14720 144 14752
rect 184 14720 216 14752
rect 256 14720 288 14752
rect 112 14648 144 14680
rect 184 14648 216 14680
rect 256 14648 288 14680
rect 112 14576 144 14608
rect 184 14576 216 14608
rect 256 14576 288 14608
rect 112 14504 144 14536
rect 184 14504 216 14536
rect 256 14504 288 14536
rect 112 14432 144 14464
rect 184 14432 216 14464
rect 256 14432 288 14464
rect 112 14360 144 14392
rect 184 14360 216 14392
rect 256 14360 288 14392
rect 112 14288 144 14320
rect 184 14288 216 14320
rect 256 14288 288 14320
rect 112 14216 144 14248
rect 184 14216 216 14248
rect 256 14216 288 14248
rect 112 14144 144 14176
rect 184 14144 216 14176
rect 256 14144 288 14176
rect 112 14072 144 14104
rect 184 14072 216 14104
rect 256 14072 288 14104
rect 112 14000 144 14032
rect 184 14000 216 14032
rect 256 14000 288 14032
rect 112 13928 144 13960
rect 184 13928 216 13960
rect 256 13928 288 13960
rect 112 13856 144 13888
rect 184 13856 216 13888
rect 256 13856 288 13888
rect 112 13784 144 13816
rect 184 13784 216 13816
rect 256 13784 288 13816
rect 112 13712 144 13744
rect 184 13712 216 13744
rect 256 13712 288 13744
rect 112 13640 144 13672
rect 184 13640 216 13672
rect 256 13640 288 13672
rect 112 13568 144 13600
rect 184 13568 216 13600
rect 256 13568 288 13600
rect 112 13496 144 13528
rect 184 13496 216 13528
rect 256 13496 288 13528
rect 112 13424 144 13456
rect 184 13424 216 13456
rect 256 13424 288 13456
rect 112 13352 144 13384
rect 184 13352 216 13384
rect 256 13352 288 13384
rect 112 13280 144 13312
rect 184 13280 216 13312
rect 256 13280 288 13312
rect 112 13208 144 13240
rect 184 13208 216 13240
rect 256 13208 288 13240
rect 112 13136 144 13168
rect 184 13136 216 13168
rect 256 13136 288 13168
rect 112 13064 144 13096
rect 184 13064 216 13096
rect 256 13064 288 13096
rect 170 31484 230 31498
rect 170 31452 184 31484
rect 216 31452 230 31484
rect 170 31430 230 31452
rect 44 31416 356 31430
rect 44 31384 116 31416
rect 148 31384 184 31416
rect 216 31384 252 31416
rect 284 31384 356 31416
rect 44 31370 356 31384
rect 170 31348 230 31370
rect 170 31316 184 31348
rect 216 31316 230 31348
rect 170 31302 230 31316
rect 44 27971 356 28034
rect 44 27939 112 27971
rect 144 27939 184 27971
rect 216 27939 256 27971
rect 288 27939 356 27971
rect 44 27899 356 27939
rect 44 27867 112 27899
rect 144 27867 184 27899
rect 216 27867 256 27899
rect 288 27867 356 27899
rect 44 27827 356 27867
rect 44 27795 112 27827
rect 144 27795 184 27827
rect 216 27795 256 27827
rect 288 27795 356 27827
rect 44 27755 356 27795
rect 44 27723 112 27755
rect 144 27723 184 27755
rect 216 27723 256 27755
rect 288 27723 356 27755
rect 44 27683 356 27723
rect 44 27651 112 27683
rect 144 27651 184 27683
rect 216 27651 256 27683
rect 288 27651 356 27683
rect 44 27611 356 27651
rect 44 27579 112 27611
rect 144 27579 184 27611
rect 216 27579 256 27611
rect 288 27579 356 27611
rect 44 27539 356 27579
rect 44 27507 112 27539
rect 144 27507 184 27539
rect 216 27507 256 27539
rect 288 27507 356 27539
rect 44 27467 356 27507
rect 44 27435 112 27467
rect 144 27435 184 27467
rect 216 27435 256 27467
rect 288 27435 356 27467
rect 44 27395 356 27435
rect 44 27363 112 27395
rect 144 27363 184 27395
rect 216 27363 256 27395
rect 288 27363 356 27395
rect 44 27323 356 27363
rect 44 27291 112 27323
rect 144 27291 184 27323
rect 216 27291 256 27323
rect 288 27291 356 27323
rect 44 27251 356 27291
rect 44 27219 112 27251
rect 144 27219 184 27251
rect 216 27219 256 27251
rect 288 27219 356 27251
rect 44 27179 356 27219
rect 44 27147 112 27179
rect 144 27147 184 27179
rect 216 27147 256 27179
rect 288 27147 356 27179
rect 44 27107 356 27147
rect 44 27075 112 27107
rect 144 27075 184 27107
rect 216 27075 256 27107
rect 288 27075 356 27107
rect 44 27035 356 27075
rect 44 27003 112 27035
rect 144 27003 184 27035
rect 216 27003 256 27035
rect 288 27003 356 27035
rect 44 26963 356 27003
rect 44 26931 112 26963
rect 144 26931 184 26963
rect 216 26931 256 26963
rect 288 26931 356 26963
rect 44 26891 356 26931
rect 44 26859 112 26891
rect 144 26859 184 26891
rect 216 26859 256 26891
rect 288 26859 356 26891
rect 44 26819 356 26859
rect 44 26787 112 26819
rect 144 26787 184 26819
rect 216 26787 256 26819
rect 288 26787 356 26819
rect 44 26747 356 26787
rect 44 26715 112 26747
rect 144 26715 184 26747
rect 216 26715 256 26747
rect 288 26715 356 26747
rect 44 26675 356 26715
rect 44 26643 112 26675
rect 144 26643 184 26675
rect 216 26643 256 26675
rect 288 26643 356 26675
rect 44 26603 356 26643
rect 44 26571 112 26603
rect 144 26571 184 26603
rect 216 26571 256 26603
rect 288 26571 356 26603
rect 44 26531 356 26571
rect 44 26499 112 26531
rect 144 26499 184 26531
rect 216 26499 256 26531
rect 288 26499 356 26531
rect 44 26459 356 26499
rect 44 26427 112 26459
rect 144 26427 184 26459
rect 216 26427 256 26459
rect 288 26427 356 26459
rect 44 26387 356 26427
rect 44 26355 112 26387
rect 144 26355 184 26387
rect 216 26355 256 26387
rect 288 26355 356 26387
rect 44 26315 356 26355
rect 44 26283 112 26315
rect 144 26283 184 26315
rect 216 26283 256 26315
rect 288 26283 356 26315
rect 44 26243 356 26283
rect 44 26211 112 26243
rect 144 26211 184 26243
rect 216 26211 256 26243
rect 288 26211 356 26243
rect 44 26171 356 26211
rect 44 26139 112 26171
rect 144 26139 184 26171
rect 216 26139 256 26171
rect 288 26139 356 26171
rect 44 26099 356 26139
rect 44 26067 112 26099
rect 144 26067 184 26099
rect 216 26067 256 26099
rect 288 26067 356 26099
rect 44 26027 356 26067
rect 44 25995 112 26027
rect 144 25995 184 26027
rect 216 25995 256 26027
rect 288 25995 356 26027
rect 44 25955 356 25995
rect 44 25923 112 25955
rect 144 25923 184 25955
rect 216 25923 256 25955
rect 288 25923 356 25955
rect 44 25883 356 25923
rect 44 25851 112 25883
rect 144 25851 184 25883
rect 216 25851 256 25883
rect 288 25851 356 25883
rect 44 25811 356 25851
rect 44 25779 112 25811
rect 144 25779 184 25811
rect 216 25779 256 25811
rect 288 25779 356 25811
rect 44 25739 356 25779
rect 44 25707 112 25739
rect 144 25707 184 25739
rect 216 25707 256 25739
rect 288 25707 356 25739
rect 44 25667 356 25707
rect 44 25635 112 25667
rect 144 25635 184 25667
rect 216 25635 256 25667
rect 288 25635 356 25667
rect 44 25595 356 25635
rect 44 25563 112 25595
rect 144 25563 184 25595
rect 216 25563 256 25595
rect 288 25563 356 25595
rect 44 25523 356 25563
rect 44 25491 112 25523
rect 144 25491 184 25523
rect 216 25491 256 25523
rect 288 25491 356 25523
rect 44 25451 356 25491
rect 44 25419 112 25451
rect 144 25419 184 25451
rect 216 25419 256 25451
rect 288 25419 356 25451
rect 44 25379 356 25419
rect 44 25347 112 25379
rect 144 25347 184 25379
rect 216 25347 256 25379
rect 288 25347 356 25379
rect 44 25307 356 25347
rect 44 25275 112 25307
rect 144 25275 184 25307
rect 216 25275 256 25307
rect 288 25275 356 25307
rect 44 25235 356 25275
rect 44 25203 112 25235
rect 144 25203 184 25235
rect 216 25203 256 25235
rect 288 25203 356 25235
rect 44 25163 356 25203
rect 44 25131 112 25163
rect 144 25131 184 25163
rect 216 25131 256 25163
rect 288 25131 356 25163
rect 44 25091 356 25131
rect 44 25059 112 25091
rect 144 25059 184 25091
rect 216 25059 256 25091
rect 288 25059 356 25091
rect 44 25019 356 25059
rect 44 24987 112 25019
rect 144 24987 184 25019
rect 216 24987 256 25019
rect 288 24987 356 25019
rect 44 24947 356 24987
rect 44 24915 112 24947
rect 144 24915 184 24947
rect 216 24915 256 24947
rect 288 24915 356 24947
rect 44 24875 356 24915
rect 44 24843 112 24875
rect 144 24843 184 24875
rect 216 24843 256 24875
rect 288 24843 356 24875
rect 44 24803 356 24843
rect 44 24771 112 24803
rect 144 24771 184 24803
rect 216 24771 256 24803
rect 288 24771 356 24803
rect 44 24731 356 24771
rect 44 24699 112 24731
rect 144 24699 184 24731
rect 216 24699 256 24731
rect 288 24699 356 24731
rect 44 24659 356 24699
rect 44 24627 112 24659
rect 144 24627 184 24659
rect 216 24627 256 24659
rect 288 24627 356 24659
rect 44 24587 356 24627
rect 44 24555 112 24587
rect 144 24555 184 24587
rect 216 24555 256 24587
rect 288 24555 356 24587
rect 44 24515 356 24555
rect 44 24483 112 24515
rect 144 24483 184 24515
rect 216 24483 256 24515
rect 288 24483 356 24515
rect 44 24443 356 24483
rect 44 24411 112 24443
rect 144 24411 184 24443
rect 216 24411 256 24443
rect 288 24411 356 24443
rect 44 24371 356 24411
rect 44 24339 112 24371
rect 144 24339 184 24371
rect 216 24339 256 24371
rect 288 24339 356 24371
rect 44 24299 356 24339
rect 44 24267 112 24299
rect 144 24267 184 24299
rect 216 24267 256 24299
rect 288 24267 356 24299
rect 44 24227 356 24267
rect 44 24195 112 24227
rect 144 24195 184 24227
rect 216 24195 256 24227
rect 288 24195 356 24227
rect 44 24155 356 24195
rect 44 24123 112 24155
rect 144 24123 184 24155
rect 216 24123 256 24155
rect 288 24123 356 24155
rect 44 24083 356 24123
rect 44 24051 112 24083
rect 144 24051 184 24083
rect 216 24051 256 24083
rect 288 24051 356 24083
rect 44 24011 356 24051
rect 44 23979 112 24011
rect 144 23979 184 24011
rect 216 23979 256 24011
rect 288 23979 356 24011
rect 44 23939 356 23979
rect 44 23907 112 23939
rect 144 23907 184 23939
rect 216 23907 256 23939
rect 288 23907 356 23939
rect 44 23867 356 23907
rect 44 23835 112 23867
rect 144 23835 184 23867
rect 216 23835 256 23867
rect 288 23835 356 23867
rect 44 23795 356 23835
rect 44 23763 112 23795
rect 144 23763 184 23795
rect 216 23763 256 23795
rect 288 23763 356 23795
rect 44 23723 356 23763
rect 44 23691 112 23723
rect 144 23691 184 23723
rect 216 23691 256 23723
rect 288 23691 356 23723
rect 44 23651 356 23691
rect 44 23619 112 23651
rect 144 23619 184 23651
rect 216 23619 256 23651
rect 288 23619 356 23651
rect 44 23579 356 23619
rect 44 23547 112 23579
rect 144 23547 184 23579
rect 216 23547 256 23579
rect 288 23547 356 23579
rect 44 23507 356 23547
rect 44 23475 112 23507
rect 144 23475 184 23507
rect 216 23475 256 23507
rect 288 23475 356 23507
rect 44 23435 356 23475
rect 44 23403 112 23435
rect 144 23403 184 23435
rect 216 23403 256 23435
rect 288 23403 356 23435
rect 44 23363 356 23403
rect 44 23331 112 23363
rect 144 23331 184 23363
rect 216 23331 256 23363
rect 288 23331 356 23363
rect 44 23291 356 23331
rect 44 23259 112 23291
rect 144 23259 184 23291
rect 216 23259 256 23291
rect 288 23259 356 23291
rect 44 23219 356 23259
rect 44 23187 112 23219
rect 144 23187 184 23219
rect 216 23187 256 23219
rect 288 23187 356 23219
rect 44 23124 356 23187
rect 44 22874 356 22924
rect 44 22842 112 22874
rect 144 22842 184 22874
rect 216 22842 256 22874
rect 288 22842 356 22874
rect 44 22802 356 22842
rect 44 22770 112 22802
rect 144 22770 184 22802
rect 216 22770 256 22802
rect 288 22770 356 22802
rect 44 22730 356 22770
rect 44 22698 112 22730
rect 144 22698 184 22730
rect 216 22698 256 22730
rect 288 22698 356 22730
rect 44 22658 356 22698
rect 44 22626 112 22658
rect 144 22626 184 22658
rect 216 22626 256 22658
rect 288 22626 356 22658
rect 44 22586 356 22626
rect 44 22554 112 22586
rect 144 22554 184 22586
rect 216 22554 256 22586
rect 288 22554 356 22586
rect 44 22514 356 22554
rect 44 22482 112 22514
rect 144 22482 184 22514
rect 216 22482 256 22514
rect 288 22482 356 22514
rect 44 22442 356 22482
rect 44 22410 112 22442
rect 144 22410 184 22442
rect 216 22410 256 22442
rect 288 22410 356 22442
rect 44 22370 356 22410
rect 44 22338 112 22370
rect 144 22338 184 22370
rect 216 22338 256 22370
rect 288 22338 356 22370
rect 44 22298 356 22338
rect 44 22266 112 22298
rect 144 22266 184 22298
rect 216 22266 256 22298
rect 288 22266 356 22298
rect 44 22226 356 22266
rect 44 22194 112 22226
rect 144 22194 184 22226
rect 216 22194 256 22226
rect 288 22194 356 22226
rect 44 22154 356 22194
rect 44 22122 112 22154
rect 144 22122 184 22154
rect 216 22122 256 22154
rect 288 22122 356 22154
rect 44 22082 356 22122
rect 44 22050 112 22082
rect 144 22050 184 22082
rect 216 22050 256 22082
rect 288 22050 356 22082
rect 44 22010 356 22050
rect 44 21978 112 22010
rect 144 21978 184 22010
rect 216 21978 256 22010
rect 288 21978 356 22010
rect 44 21938 356 21978
rect 44 21906 112 21938
rect 144 21906 184 21938
rect 216 21906 256 21938
rect 288 21906 356 21938
rect 44 21866 356 21906
rect 44 21834 112 21866
rect 144 21834 184 21866
rect 216 21834 256 21866
rect 288 21834 356 21866
rect 44 21794 356 21834
rect 44 21762 112 21794
rect 144 21762 184 21794
rect 216 21762 256 21794
rect 288 21762 356 21794
rect 44 21722 356 21762
rect 44 21690 112 21722
rect 144 21690 184 21722
rect 216 21690 256 21722
rect 288 21690 356 21722
rect 44 21650 356 21690
rect 44 21618 112 21650
rect 144 21618 184 21650
rect 216 21618 256 21650
rect 288 21618 356 21650
rect 44 21578 356 21618
rect 44 21546 112 21578
rect 144 21546 184 21578
rect 216 21546 256 21578
rect 288 21546 356 21578
rect 44 21506 356 21546
rect 44 21474 112 21506
rect 144 21474 184 21506
rect 216 21474 256 21506
rect 288 21474 356 21506
rect 44 21434 356 21474
rect 44 21402 112 21434
rect 144 21402 184 21434
rect 216 21402 256 21434
rect 288 21402 356 21434
rect 44 21362 356 21402
rect 44 21330 112 21362
rect 144 21330 184 21362
rect 216 21330 256 21362
rect 288 21330 356 21362
rect 44 21290 356 21330
rect 44 21258 112 21290
rect 144 21258 184 21290
rect 216 21258 256 21290
rect 288 21258 356 21290
rect 44 21218 356 21258
rect 44 21186 112 21218
rect 144 21186 184 21218
rect 216 21186 256 21218
rect 288 21186 356 21218
rect 44 21146 356 21186
rect 44 21114 112 21146
rect 144 21114 184 21146
rect 216 21114 256 21146
rect 288 21114 356 21146
rect 44 21074 356 21114
rect 44 21042 112 21074
rect 144 21042 184 21074
rect 216 21042 256 21074
rect 288 21042 356 21074
rect 44 21002 356 21042
rect 44 20970 112 21002
rect 144 20970 184 21002
rect 216 20970 256 21002
rect 288 20970 356 21002
rect 44 20930 356 20970
rect 44 20898 112 20930
rect 144 20898 184 20930
rect 216 20898 256 20930
rect 288 20898 356 20930
rect 44 20858 356 20898
rect 44 20826 112 20858
rect 144 20826 184 20858
rect 216 20826 256 20858
rect 288 20826 356 20858
rect 44 20786 356 20826
rect 44 20754 112 20786
rect 144 20754 184 20786
rect 216 20754 256 20786
rect 288 20754 356 20786
rect 44 20714 356 20754
rect 44 20682 112 20714
rect 144 20682 184 20714
rect 216 20682 256 20714
rect 288 20682 356 20714
rect 44 20642 356 20682
rect 44 20610 112 20642
rect 144 20610 184 20642
rect 216 20610 256 20642
rect 288 20610 356 20642
rect 44 20570 356 20610
rect 44 20538 112 20570
rect 144 20538 184 20570
rect 216 20538 256 20570
rect 288 20538 356 20570
rect 44 20498 356 20538
rect 44 20466 112 20498
rect 144 20466 184 20498
rect 216 20466 256 20498
rect 288 20466 356 20498
rect 44 20426 356 20466
rect 44 20394 112 20426
rect 144 20394 184 20426
rect 216 20394 256 20426
rect 288 20394 356 20426
rect 44 20354 356 20394
rect 44 20322 112 20354
rect 144 20322 184 20354
rect 216 20322 256 20354
rect 288 20322 356 20354
rect 44 20282 356 20322
rect 44 20250 112 20282
rect 144 20250 184 20282
rect 216 20250 256 20282
rect 288 20250 356 20282
rect 44 20210 356 20250
rect 44 20178 112 20210
rect 144 20178 184 20210
rect 216 20178 256 20210
rect 288 20178 356 20210
rect 44 20138 356 20178
rect 44 20106 112 20138
rect 144 20106 184 20138
rect 216 20106 256 20138
rect 288 20106 356 20138
rect 44 20066 356 20106
rect 44 20034 112 20066
rect 144 20034 184 20066
rect 216 20034 256 20066
rect 288 20034 356 20066
rect 44 19994 356 20034
rect 44 19962 112 19994
rect 144 19962 184 19994
rect 216 19962 256 19994
rect 288 19962 356 19994
rect 44 19922 356 19962
rect 44 19890 112 19922
rect 144 19890 184 19922
rect 216 19890 256 19922
rect 288 19890 356 19922
rect 44 19850 356 19890
rect 44 19818 112 19850
rect 144 19818 184 19850
rect 216 19818 256 19850
rect 288 19818 356 19850
rect 44 19778 356 19818
rect 44 19746 112 19778
rect 144 19746 184 19778
rect 216 19746 256 19778
rect 288 19746 356 19778
rect 44 19706 356 19746
rect 44 19674 112 19706
rect 144 19674 184 19706
rect 216 19674 256 19706
rect 288 19674 356 19706
rect 44 19634 356 19674
rect 44 19602 112 19634
rect 144 19602 184 19634
rect 216 19602 256 19634
rect 288 19602 356 19634
rect 44 19562 356 19602
rect 44 19530 112 19562
rect 144 19530 184 19562
rect 216 19530 256 19562
rect 288 19530 356 19562
rect 44 19490 356 19530
rect 44 19458 112 19490
rect 144 19458 184 19490
rect 216 19458 256 19490
rect 288 19458 356 19490
rect 44 19418 356 19458
rect 44 19386 112 19418
rect 144 19386 184 19418
rect 216 19386 256 19418
rect 288 19386 356 19418
rect 44 19346 356 19386
rect 44 19314 112 19346
rect 144 19314 184 19346
rect 216 19314 256 19346
rect 288 19314 356 19346
rect 44 19274 356 19314
rect 44 19242 112 19274
rect 144 19242 184 19274
rect 216 19242 256 19274
rect 288 19242 356 19274
rect 44 19202 356 19242
rect 44 19170 112 19202
rect 144 19170 184 19202
rect 216 19170 256 19202
rect 288 19170 356 19202
rect 44 19130 356 19170
rect 44 19098 112 19130
rect 144 19098 184 19130
rect 216 19098 256 19130
rect 288 19098 356 19130
rect 44 19058 356 19098
rect 44 19026 112 19058
rect 144 19026 184 19058
rect 216 19026 256 19058
rect 288 19026 356 19058
rect 44 18986 356 19026
rect 44 18954 112 18986
rect 144 18954 184 18986
rect 216 18954 256 18986
rect 288 18954 356 18986
rect 44 18914 356 18954
rect 44 18882 112 18914
rect 144 18882 184 18914
rect 216 18882 256 18914
rect 288 18882 356 18914
rect 44 18842 356 18882
rect 44 18810 112 18842
rect 144 18810 184 18842
rect 216 18810 256 18842
rect 288 18810 356 18842
rect 44 18770 356 18810
rect 44 18738 112 18770
rect 144 18738 184 18770
rect 216 18738 256 18770
rect 288 18738 356 18770
rect 44 18698 356 18738
rect 44 18666 112 18698
rect 144 18666 184 18698
rect 216 18666 256 18698
rect 288 18666 356 18698
rect 44 18626 356 18666
rect 44 18594 112 18626
rect 144 18594 184 18626
rect 216 18594 256 18626
rect 288 18594 356 18626
rect 44 18554 356 18594
rect 44 18522 112 18554
rect 144 18522 184 18554
rect 216 18522 256 18554
rect 288 18522 356 18554
rect 44 18482 356 18522
rect 44 18450 112 18482
rect 144 18450 184 18482
rect 216 18450 256 18482
rect 288 18450 356 18482
rect 44 18410 356 18450
rect 44 18378 112 18410
rect 144 18378 184 18410
rect 216 18378 256 18410
rect 288 18378 356 18410
rect 44 18338 356 18378
rect 44 18306 112 18338
rect 144 18306 184 18338
rect 216 18306 256 18338
rect 288 18306 356 18338
rect 44 18266 356 18306
rect 44 18234 112 18266
rect 144 18234 184 18266
rect 216 18234 256 18266
rect 288 18234 356 18266
rect 44 18194 356 18234
rect 44 18162 112 18194
rect 144 18162 184 18194
rect 216 18162 256 18194
rect 288 18162 356 18194
rect 44 18112 356 18162
rect 44 17848 356 17912
rect 44 17816 112 17848
rect 144 17816 184 17848
rect 216 17816 256 17848
rect 288 17816 356 17848
rect 44 17776 356 17816
rect 44 17744 112 17776
rect 144 17744 184 17776
rect 216 17744 256 17776
rect 288 17744 356 17776
rect 44 17704 356 17744
rect 44 17672 112 17704
rect 144 17672 184 17704
rect 216 17672 256 17704
rect 288 17672 356 17704
rect 44 17632 356 17672
rect 44 17600 112 17632
rect 144 17600 184 17632
rect 216 17600 256 17632
rect 288 17600 356 17632
rect 44 17560 356 17600
rect 44 17528 112 17560
rect 144 17528 184 17560
rect 216 17528 256 17560
rect 288 17528 356 17560
rect 44 17488 356 17528
rect 44 17456 112 17488
rect 144 17456 184 17488
rect 216 17456 256 17488
rect 288 17456 356 17488
rect 44 17416 356 17456
rect 44 17384 112 17416
rect 144 17384 184 17416
rect 216 17384 256 17416
rect 288 17384 356 17416
rect 44 17344 356 17384
rect 44 17312 112 17344
rect 144 17312 184 17344
rect 216 17312 256 17344
rect 288 17312 356 17344
rect 44 17272 356 17312
rect 44 17240 112 17272
rect 144 17240 184 17272
rect 216 17240 256 17272
rect 288 17240 356 17272
rect 44 17200 356 17240
rect 44 17168 112 17200
rect 144 17168 184 17200
rect 216 17168 256 17200
rect 288 17168 356 17200
rect 44 17128 356 17168
rect 44 17096 112 17128
rect 144 17096 184 17128
rect 216 17096 256 17128
rect 288 17096 356 17128
rect 44 17056 356 17096
rect 44 17024 112 17056
rect 144 17024 184 17056
rect 216 17024 256 17056
rect 288 17024 356 17056
rect 44 16984 356 17024
rect 44 16952 112 16984
rect 144 16952 184 16984
rect 216 16952 256 16984
rect 288 16952 356 16984
rect 44 16912 356 16952
rect 44 16880 112 16912
rect 144 16880 184 16912
rect 216 16880 256 16912
rect 288 16880 356 16912
rect 44 16840 356 16880
rect 44 16808 112 16840
rect 144 16808 184 16840
rect 216 16808 256 16840
rect 288 16808 356 16840
rect 44 16768 356 16808
rect 44 16736 112 16768
rect 144 16736 184 16768
rect 216 16736 256 16768
rect 288 16736 356 16768
rect 44 16696 356 16736
rect 44 16664 112 16696
rect 144 16664 184 16696
rect 216 16664 256 16696
rect 288 16664 356 16696
rect 44 16624 356 16664
rect 44 16592 112 16624
rect 144 16592 184 16624
rect 216 16592 256 16624
rect 288 16592 356 16624
rect 44 16552 356 16592
rect 44 16520 112 16552
rect 144 16520 184 16552
rect 216 16520 256 16552
rect 288 16520 356 16552
rect 44 16480 356 16520
rect 44 16448 112 16480
rect 144 16448 184 16480
rect 216 16448 256 16480
rect 288 16448 356 16480
rect 44 16408 356 16448
rect 44 16376 112 16408
rect 144 16376 184 16408
rect 216 16376 256 16408
rect 288 16376 356 16408
rect 44 16336 356 16376
rect 44 16304 112 16336
rect 144 16304 184 16336
rect 216 16304 256 16336
rect 288 16304 356 16336
rect 44 16264 356 16304
rect 44 16232 112 16264
rect 144 16232 184 16264
rect 216 16232 256 16264
rect 288 16232 356 16264
rect 44 16192 356 16232
rect 44 16160 112 16192
rect 144 16160 184 16192
rect 216 16160 256 16192
rect 288 16160 356 16192
rect 44 16120 356 16160
rect 44 16088 112 16120
rect 144 16088 184 16120
rect 216 16088 256 16120
rect 288 16088 356 16120
rect 44 16048 356 16088
rect 44 16016 112 16048
rect 144 16016 184 16048
rect 216 16016 256 16048
rect 288 16016 356 16048
rect 44 15976 356 16016
rect 44 15944 112 15976
rect 144 15944 184 15976
rect 216 15944 256 15976
rect 288 15944 356 15976
rect 44 15904 356 15944
rect 44 15872 112 15904
rect 144 15872 184 15904
rect 216 15872 256 15904
rect 288 15872 356 15904
rect 44 15832 356 15872
rect 44 15800 112 15832
rect 144 15800 184 15832
rect 216 15800 256 15832
rect 288 15800 356 15832
rect 44 15760 356 15800
rect 44 15728 112 15760
rect 144 15728 184 15760
rect 216 15728 256 15760
rect 288 15728 356 15760
rect 44 15688 356 15728
rect 44 15656 112 15688
rect 144 15656 184 15688
rect 216 15656 256 15688
rect 288 15656 356 15688
rect 44 15616 356 15656
rect 44 15584 112 15616
rect 144 15584 184 15616
rect 216 15584 256 15616
rect 288 15584 356 15616
rect 44 15544 356 15584
rect 44 15512 112 15544
rect 144 15512 184 15544
rect 216 15512 256 15544
rect 288 15512 356 15544
rect 44 15472 356 15512
rect 44 15440 112 15472
rect 144 15440 184 15472
rect 216 15440 256 15472
rect 288 15440 356 15472
rect 44 15400 356 15440
rect 44 15368 112 15400
rect 144 15368 184 15400
rect 216 15368 256 15400
rect 288 15368 356 15400
rect 44 15328 356 15368
rect 44 15296 112 15328
rect 144 15296 184 15328
rect 216 15296 256 15328
rect 288 15296 356 15328
rect 44 15256 356 15296
rect 44 15224 112 15256
rect 144 15224 184 15256
rect 216 15224 256 15256
rect 288 15224 356 15256
rect 44 15184 356 15224
rect 44 15152 112 15184
rect 144 15152 184 15184
rect 216 15152 256 15184
rect 288 15152 356 15184
rect 44 15112 356 15152
rect 44 15080 112 15112
rect 144 15080 184 15112
rect 216 15080 256 15112
rect 288 15080 356 15112
rect 44 15040 356 15080
rect 44 15008 112 15040
rect 144 15008 184 15040
rect 216 15008 256 15040
rect 288 15008 356 15040
rect 44 14968 356 15008
rect 44 14936 112 14968
rect 144 14936 184 14968
rect 216 14936 256 14968
rect 288 14936 356 14968
rect 44 14896 356 14936
rect 44 14864 112 14896
rect 144 14864 184 14896
rect 216 14864 256 14896
rect 288 14864 356 14896
rect 44 14824 356 14864
rect 44 14792 112 14824
rect 144 14792 184 14824
rect 216 14792 256 14824
rect 288 14792 356 14824
rect 44 14752 356 14792
rect 44 14720 112 14752
rect 144 14720 184 14752
rect 216 14720 256 14752
rect 288 14720 356 14752
rect 44 14680 356 14720
rect 44 14648 112 14680
rect 144 14648 184 14680
rect 216 14648 256 14680
rect 288 14648 356 14680
rect 44 14608 356 14648
rect 44 14576 112 14608
rect 144 14576 184 14608
rect 216 14576 256 14608
rect 288 14576 356 14608
rect 44 14536 356 14576
rect 44 14504 112 14536
rect 144 14504 184 14536
rect 216 14504 256 14536
rect 288 14504 356 14536
rect 44 14464 356 14504
rect 44 14432 112 14464
rect 144 14432 184 14464
rect 216 14432 256 14464
rect 288 14432 356 14464
rect 44 14392 356 14432
rect 44 14360 112 14392
rect 144 14360 184 14392
rect 216 14360 256 14392
rect 288 14360 356 14392
rect 44 14320 356 14360
rect 44 14288 112 14320
rect 144 14288 184 14320
rect 216 14288 256 14320
rect 288 14288 356 14320
rect 44 14248 356 14288
rect 44 14216 112 14248
rect 144 14216 184 14248
rect 216 14216 256 14248
rect 288 14216 356 14248
rect 44 14176 356 14216
rect 44 14144 112 14176
rect 144 14144 184 14176
rect 216 14144 256 14176
rect 288 14144 356 14176
rect 44 14104 356 14144
rect 44 14072 112 14104
rect 144 14072 184 14104
rect 216 14072 256 14104
rect 288 14072 356 14104
rect 44 14032 356 14072
rect 44 14000 112 14032
rect 144 14000 184 14032
rect 216 14000 256 14032
rect 288 14000 356 14032
rect 44 13960 356 14000
rect 44 13928 112 13960
rect 144 13928 184 13960
rect 216 13928 256 13960
rect 288 13928 356 13960
rect 44 13888 356 13928
rect 44 13856 112 13888
rect 144 13856 184 13888
rect 216 13856 256 13888
rect 288 13856 356 13888
rect 44 13816 356 13856
rect 44 13784 112 13816
rect 144 13784 184 13816
rect 216 13784 256 13816
rect 288 13784 356 13816
rect 44 13744 356 13784
rect 44 13712 112 13744
rect 144 13712 184 13744
rect 216 13712 256 13744
rect 288 13712 356 13744
rect 44 13672 356 13712
rect 44 13640 112 13672
rect 144 13640 184 13672
rect 216 13640 256 13672
rect 288 13640 356 13672
rect 44 13600 356 13640
rect 44 13568 112 13600
rect 144 13568 184 13600
rect 216 13568 256 13600
rect 288 13568 356 13600
rect 44 13528 356 13568
rect 44 13496 112 13528
rect 144 13496 184 13528
rect 216 13496 256 13528
rect 288 13496 356 13528
rect 44 13456 356 13496
rect 44 13424 112 13456
rect 144 13424 184 13456
rect 216 13424 256 13456
rect 288 13424 356 13456
rect 44 13384 356 13424
rect 44 13352 112 13384
rect 144 13352 184 13384
rect 216 13352 256 13384
rect 288 13352 356 13384
rect 44 13312 356 13352
rect 44 13280 112 13312
rect 144 13280 184 13312
rect 216 13280 256 13312
rect 288 13280 356 13312
rect 44 13240 356 13280
rect 44 13208 112 13240
rect 144 13208 184 13240
rect 216 13208 256 13240
rect 288 13208 356 13240
rect 44 13168 356 13208
rect 44 13136 112 13168
rect 144 13136 184 13168
rect 216 13136 256 13168
rect 288 13136 356 13168
rect 44 13096 356 13136
rect 44 13064 112 13096
rect 144 13064 184 13096
rect 216 13064 256 13096
rect 288 13064 356 13096
rect 44 13000 356 13064
<< nsubdiff >>
rect 184 33384 216 33416
rect 256 33384 288 33416
rect 184 29684 216 29716
rect 256 29684 288 29716
rect 112 12112 144 12144
rect 184 12112 216 12144
rect 256 12112 288 12144
rect 328 12112 360 12144
rect 40 12040 72 12072
rect 112 12040 144 12072
rect 184 12040 216 12072
rect 256 12040 288 12072
rect 328 12040 360 12072
rect 40 11968 72 12000
rect 112 11968 144 12000
rect 184 11968 216 12000
rect 256 11968 288 12000
rect 328 11968 360 12000
rect 40 11896 72 11928
rect 112 11896 144 11928
rect 184 11896 216 11928
rect 256 11896 288 11928
rect 328 11896 360 11928
rect 40 11824 72 11856
rect 112 11824 144 11856
rect 184 11824 216 11856
rect 256 11824 288 11856
rect 328 11824 360 11856
rect 40 11752 72 11784
rect 112 11752 144 11784
rect 184 11752 216 11784
rect 256 11752 288 11784
rect 328 11752 360 11784
rect 40 11680 72 11712
rect 112 11680 144 11712
rect 184 11680 216 11712
rect 256 11680 288 11712
rect 328 11680 360 11712
rect 40 11608 72 11640
rect 112 11608 144 11640
rect 184 11608 216 11640
rect 256 11608 288 11640
rect 328 11608 360 11640
rect 40 11536 72 11568
rect 112 11536 144 11568
rect 184 11536 216 11568
rect 256 11536 288 11568
rect 328 11536 360 11568
rect 40 11464 72 11496
rect 112 11464 144 11496
rect 184 11464 216 11496
rect 256 11464 288 11496
rect 328 11464 360 11496
rect 40 11392 72 11424
rect 112 11392 144 11424
rect 184 11392 216 11424
rect 256 11392 288 11424
rect 328 11392 360 11424
rect 40 11320 72 11352
rect 112 11320 144 11352
rect 184 11320 216 11352
rect 256 11320 288 11352
rect 328 11320 360 11352
rect 40 11248 72 11280
rect 112 11248 144 11280
rect 184 11248 216 11280
rect 256 11248 288 11280
rect 328 11248 360 11280
rect 40 11176 72 11208
rect 112 11176 144 11208
rect 184 11176 216 11208
rect 256 11176 288 11208
rect 328 11176 360 11208
rect 40 11104 72 11136
rect 112 11104 144 11136
rect 184 11104 216 11136
rect 256 11104 288 11136
rect 328 11104 360 11136
rect 40 11032 72 11064
rect 112 11032 144 11064
rect 184 11032 216 11064
rect 256 11032 288 11064
rect 328 11032 360 11064
rect 40 10960 72 10992
rect 112 10960 144 10992
rect 184 10960 216 10992
rect 256 10960 288 10992
rect 328 10960 360 10992
rect 40 10888 72 10920
rect 112 10888 144 10920
rect 184 10888 216 10920
rect 256 10888 288 10920
rect 328 10888 360 10920
rect 40 10816 72 10848
rect 112 10816 144 10848
rect 184 10816 216 10848
rect 256 10816 288 10848
rect 328 10816 360 10848
rect 40 10744 72 10776
rect 112 10744 144 10776
rect 184 10744 216 10776
rect 256 10744 288 10776
rect 328 10744 360 10776
rect 40 10672 72 10704
rect 112 10672 144 10704
rect 184 10672 216 10704
rect 256 10672 288 10704
rect 328 10672 360 10704
rect 40 10600 72 10632
rect 112 10600 144 10632
rect 184 10600 216 10632
rect 256 10600 288 10632
rect 328 10600 360 10632
rect 40 10528 72 10560
rect 112 10528 144 10560
rect 184 10528 216 10560
rect 256 10528 288 10560
rect 328 10528 360 10560
rect 40 10456 72 10488
rect 112 10456 144 10488
rect 184 10456 216 10488
rect 256 10456 288 10488
rect 328 10456 360 10488
rect 40 10384 72 10416
rect 112 10384 144 10416
rect 184 10384 216 10416
rect 256 10384 288 10416
rect 328 10384 360 10416
rect 40 10312 72 10344
rect 112 10312 144 10344
rect 184 10312 216 10344
rect 256 10312 288 10344
rect 328 10312 360 10344
rect 40 10240 72 10272
rect 112 10240 144 10272
rect 184 10240 216 10272
rect 256 10240 288 10272
rect 328 10240 360 10272
rect 40 10168 72 10200
rect 112 10168 144 10200
rect 184 10168 216 10200
rect 256 10168 288 10200
rect 328 10168 360 10200
rect 40 10096 72 10128
rect 112 10096 144 10128
rect 184 10096 216 10128
rect 256 10096 288 10128
rect 328 10096 360 10128
rect 40 10024 72 10056
rect 112 10024 144 10056
rect 184 10024 216 10056
rect 256 10024 288 10056
rect 328 10024 360 10056
rect 40 9952 72 9984
rect 112 9952 144 9984
rect 184 9952 216 9984
rect 256 9952 288 9984
rect 328 9952 360 9984
rect 40 9880 72 9912
rect 112 9880 144 9912
rect 184 9880 216 9912
rect 256 9880 288 9912
rect 328 9880 360 9912
rect 40 9808 72 9840
rect 112 9808 144 9840
rect 184 9808 216 9840
rect 256 9808 288 9840
rect 328 9808 360 9840
rect 40 9736 72 9768
rect 112 9736 144 9768
rect 184 9736 216 9768
rect 256 9736 288 9768
rect 328 9736 360 9768
rect 40 9664 72 9696
rect 112 9664 144 9696
rect 184 9664 216 9696
rect 256 9664 288 9696
rect 328 9664 360 9696
rect 40 9592 72 9624
rect 112 9592 144 9624
rect 184 9592 216 9624
rect 256 9592 288 9624
rect 328 9592 360 9624
rect 40 9520 72 9552
rect 112 9520 144 9552
rect 184 9520 216 9552
rect 256 9520 288 9552
rect 328 9520 360 9552
rect 40 9448 72 9480
rect 112 9448 144 9480
rect 184 9448 216 9480
rect 256 9448 288 9480
rect 328 9448 360 9480
rect 40 9376 72 9408
rect 112 9376 144 9408
rect 184 9376 216 9408
rect 256 9376 288 9408
rect 328 9376 360 9408
rect 40 9304 72 9336
rect 112 9304 144 9336
rect 184 9304 216 9336
rect 256 9304 288 9336
rect 328 9304 360 9336
rect 40 9232 72 9264
rect 112 9232 144 9264
rect 184 9232 216 9264
rect 256 9232 288 9264
rect 328 9232 360 9264
rect 40 9160 72 9192
rect 112 9160 144 9192
rect 184 9160 216 9192
rect 256 9160 288 9192
rect 328 9160 360 9192
rect 40 9088 72 9120
rect 112 9088 144 9120
rect 184 9088 216 9120
rect 256 9088 288 9120
rect 328 9088 360 9120
rect 40 9016 72 9048
rect 112 9016 144 9048
rect 184 9016 216 9048
rect 256 9016 288 9048
rect 328 9016 360 9048
rect 40 8944 72 8976
rect 112 8944 144 8976
rect 184 8944 216 8976
rect 256 8944 288 8976
rect 328 8944 360 8976
rect 40 8872 72 8904
rect 112 8872 144 8904
rect 184 8872 216 8904
rect 256 8872 288 8904
rect 328 8872 360 8904
rect 40 8800 72 8832
rect 112 8800 144 8832
rect 184 8800 216 8832
rect 256 8800 288 8832
rect 328 8800 360 8832
rect 40 8728 72 8760
rect 112 8728 144 8760
rect 184 8728 216 8760
rect 256 8728 288 8760
rect 328 8728 360 8760
rect 40 8656 72 8688
rect 112 8656 144 8688
rect 184 8656 216 8688
rect 256 8656 288 8688
rect 328 8656 360 8688
rect 40 8584 72 8616
rect 112 8584 144 8616
rect 184 8584 216 8616
rect 256 8584 288 8616
rect 328 8584 360 8616
rect 40 8512 72 8544
rect 112 8512 144 8544
rect 184 8512 216 8544
rect 256 8512 288 8544
rect 328 8512 360 8544
rect 40 8440 72 8472
rect 112 8440 144 8472
rect 184 8440 216 8472
rect 256 8440 288 8472
rect 328 8440 360 8472
rect 40 8368 72 8400
rect 112 8368 144 8400
rect 184 8368 216 8400
rect 256 8368 288 8400
rect 328 8368 360 8400
rect 40 8296 72 8328
rect 112 8296 144 8328
rect 184 8296 216 8328
rect 256 8296 288 8328
rect 328 8296 360 8328
rect 40 8224 72 8256
rect 112 8224 144 8256
rect 184 8224 216 8256
rect 256 8224 288 8256
rect 328 8224 360 8256
rect 40 8152 72 8184
rect 112 8152 144 8184
rect 184 8152 216 8184
rect 256 8152 288 8184
rect 328 8152 360 8184
rect 40 8080 72 8112
rect 112 8080 144 8112
rect 184 8080 216 8112
rect 256 8080 288 8112
rect 328 8080 360 8112
rect 40 8008 72 8040
rect 112 8008 144 8040
rect 184 8008 216 8040
rect 256 8008 288 8040
rect 328 8008 360 8040
rect 40 7936 72 7968
rect 112 7936 144 7968
rect 184 7936 216 7968
rect 256 7936 288 7968
rect 328 7936 360 7968
rect 40 7864 72 7896
rect 112 7864 144 7896
rect 184 7864 216 7896
rect 256 7864 288 7896
rect 328 7864 360 7896
rect 40 7792 72 7824
rect 112 7792 144 7824
rect 184 7792 216 7824
rect 256 7792 288 7824
rect 328 7792 360 7824
rect 40 7720 72 7752
rect 112 7720 144 7752
rect 184 7720 216 7752
rect 256 7720 288 7752
rect 328 7720 360 7752
rect 40 7648 72 7680
rect 112 7648 144 7680
rect 184 7648 216 7680
rect 256 7648 288 7680
rect 328 7648 360 7680
rect 40 7576 72 7608
rect 112 7576 144 7608
rect 184 7576 216 7608
rect 256 7576 288 7608
rect 328 7576 360 7608
rect 40 7504 72 7536
rect 112 7504 144 7536
rect 184 7504 216 7536
rect 256 7504 288 7536
rect 328 7504 360 7536
rect 40 7432 72 7464
rect 112 7432 144 7464
rect 184 7432 216 7464
rect 256 7432 288 7464
rect 328 7432 360 7464
rect 40 7360 72 7392
rect 112 7360 144 7392
rect 184 7360 216 7392
rect 256 7360 288 7392
rect 328 7360 360 7392
rect 40 7288 72 7320
rect 112 7288 144 7320
rect 184 7288 216 7320
rect 256 7288 288 7320
rect 328 7288 360 7320
rect 40 7216 72 7248
rect 112 7216 144 7248
rect 184 7216 216 7248
rect 256 7216 288 7248
rect 328 7216 360 7248
rect 40 7144 72 7176
rect 112 7144 144 7176
rect 184 7144 216 7176
rect 256 7144 288 7176
rect 328 7144 360 7176
rect 40 7072 72 7104
rect 112 7072 144 7104
rect 184 7072 216 7104
rect 256 7072 288 7104
rect 328 7072 360 7104
rect 40 7000 72 7032
rect 112 7000 144 7032
rect 184 7000 216 7032
rect 256 7000 288 7032
rect 328 7000 360 7032
rect 40 6928 72 6960
rect 112 6928 144 6960
rect 184 6928 216 6960
rect 256 6928 288 6960
rect 328 6928 360 6960
rect 40 6856 72 6888
rect 112 6856 144 6888
rect 184 6856 216 6888
rect 256 6856 288 6888
rect 328 6856 360 6888
rect 112 6512 144 6544
rect 184 6512 216 6544
rect 256 6512 288 6544
rect 328 6512 360 6544
rect 40 6440 72 6472
rect 112 6440 144 6472
rect 184 6440 216 6472
rect 256 6440 288 6472
rect 328 6440 360 6472
rect 40 6368 72 6400
rect 112 6368 144 6400
rect 184 6368 216 6400
rect 256 6368 288 6400
rect 328 6368 360 6400
rect 40 6296 72 6328
rect 112 6296 144 6328
rect 184 6296 216 6328
rect 256 6296 288 6328
rect 328 6296 360 6328
rect 40 6224 72 6256
rect 112 6224 144 6256
rect 184 6224 216 6256
rect 256 6224 288 6256
rect 328 6224 360 6256
rect 40 6152 72 6184
rect 112 6152 144 6184
rect 184 6152 216 6184
rect 256 6152 288 6184
rect 328 6152 360 6184
rect 40 6080 72 6112
rect 112 6080 144 6112
rect 184 6080 216 6112
rect 256 6080 288 6112
rect 328 6080 360 6112
rect 40 6008 72 6040
rect 112 6008 144 6040
rect 184 6008 216 6040
rect 256 6008 288 6040
rect 328 6008 360 6040
rect 40 5936 72 5968
rect 112 5936 144 5968
rect 184 5936 216 5968
rect 256 5936 288 5968
rect 328 5936 360 5968
rect 40 5864 72 5896
rect 112 5864 144 5896
rect 184 5864 216 5896
rect 256 5864 288 5896
rect 328 5864 360 5896
rect 40 5792 72 5824
rect 112 5792 144 5824
rect 184 5792 216 5824
rect 256 5792 288 5824
rect 328 5792 360 5824
rect 40 5720 72 5752
rect 112 5720 144 5752
rect 184 5720 216 5752
rect 256 5720 288 5752
rect 328 5720 360 5752
rect 40 5648 72 5680
rect 112 5648 144 5680
rect 184 5648 216 5680
rect 256 5648 288 5680
rect 328 5648 360 5680
rect 40 5576 72 5608
rect 112 5576 144 5608
rect 184 5576 216 5608
rect 256 5576 288 5608
rect 328 5576 360 5608
rect 40 5504 72 5536
rect 112 5504 144 5536
rect 184 5504 216 5536
rect 256 5504 288 5536
rect 328 5504 360 5536
rect 40 5432 72 5464
rect 112 5432 144 5464
rect 184 5432 216 5464
rect 256 5432 288 5464
rect 328 5432 360 5464
rect 40 5360 72 5392
rect 112 5360 144 5392
rect 184 5360 216 5392
rect 256 5360 288 5392
rect 328 5360 360 5392
rect 40 5288 72 5320
rect 112 5288 144 5320
rect 184 5288 216 5320
rect 256 5288 288 5320
rect 328 5288 360 5320
rect 40 5216 72 5248
rect 112 5216 144 5248
rect 184 5216 216 5248
rect 256 5216 288 5248
rect 328 5216 360 5248
rect 40 5144 72 5176
rect 112 5144 144 5176
rect 184 5144 216 5176
rect 256 5144 288 5176
rect 328 5144 360 5176
rect 40 5072 72 5104
rect 112 5072 144 5104
rect 184 5072 216 5104
rect 256 5072 288 5104
rect 328 5072 360 5104
rect 40 5000 72 5032
rect 112 5000 144 5032
rect 184 5000 216 5032
rect 256 5000 288 5032
rect 328 5000 360 5032
rect 40 4928 72 4960
rect 112 4928 144 4960
rect 184 4928 216 4960
rect 256 4928 288 4960
rect 328 4928 360 4960
rect 40 4856 72 4888
rect 112 4856 144 4888
rect 184 4856 216 4888
rect 256 4856 288 4888
rect 328 4856 360 4888
rect 40 4784 72 4816
rect 112 4784 144 4816
rect 184 4784 216 4816
rect 256 4784 288 4816
rect 328 4784 360 4816
rect 40 4712 72 4744
rect 112 4712 144 4744
rect 184 4712 216 4744
rect 256 4712 288 4744
rect 328 4712 360 4744
rect 40 4640 72 4672
rect 112 4640 144 4672
rect 184 4640 216 4672
rect 256 4640 288 4672
rect 328 4640 360 4672
rect 40 4568 72 4600
rect 112 4568 144 4600
rect 184 4568 216 4600
rect 256 4568 288 4600
rect 328 4568 360 4600
rect 40 4496 72 4528
rect 112 4496 144 4528
rect 184 4496 216 4528
rect 256 4496 288 4528
rect 328 4496 360 4528
rect 40 4424 72 4456
rect 112 4424 144 4456
rect 184 4424 216 4456
rect 256 4424 288 4456
rect 328 4424 360 4456
rect 40 4352 72 4384
rect 112 4352 144 4384
rect 184 4352 216 4384
rect 256 4352 288 4384
rect 328 4352 360 4384
rect 40 4280 72 4312
rect 112 4280 144 4312
rect 184 4280 216 4312
rect 256 4280 288 4312
rect 328 4280 360 4312
rect 40 4208 72 4240
rect 112 4208 144 4240
rect 184 4208 216 4240
rect 256 4208 288 4240
rect 328 4208 360 4240
rect 40 4136 72 4168
rect 112 4136 144 4168
rect 184 4136 216 4168
rect 256 4136 288 4168
rect 328 4136 360 4168
rect 40 4064 72 4096
rect 112 4064 144 4096
rect 184 4064 216 4096
rect 256 4064 288 4096
rect 328 4064 360 4096
rect 40 3992 72 4024
rect 112 3992 144 4024
rect 184 3992 216 4024
rect 256 3992 288 4024
rect 328 3992 360 4024
rect 40 3920 72 3952
rect 112 3920 144 3952
rect 184 3920 216 3952
rect 256 3920 288 3952
rect 328 3920 360 3952
rect 40 3848 72 3880
rect 112 3848 144 3880
rect 184 3848 216 3880
rect 256 3848 288 3880
rect 328 3848 360 3880
rect 40 3776 72 3808
rect 112 3776 144 3808
rect 184 3776 216 3808
rect 256 3776 288 3808
rect 328 3776 360 3808
rect 40 3704 72 3736
rect 112 3704 144 3736
rect 184 3704 216 3736
rect 256 3704 288 3736
rect 328 3704 360 3736
rect 40 3632 72 3664
rect 112 3632 144 3664
rect 184 3632 216 3664
rect 256 3632 288 3664
rect 328 3632 360 3664
rect 40 3560 72 3592
rect 112 3560 144 3592
rect 184 3560 216 3592
rect 256 3560 288 3592
rect 328 3560 360 3592
rect 40 3488 72 3520
rect 112 3488 144 3520
rect 184 3488 216 3520
rect 256 3488 288 3520
rect 328 3488 360 3520
rect 40 3416 72 3448
rect 112 3416 144 3448
rect 184 3416 216 3448
rect 256 3416 288 3448
rect 328 3416 360 3448
rect 40 3344 72 3376
rect 112 3344 144 3376
rect 184 3344 216 3376
rect 256 3344 288 3376
rect 328 3344 360 3376
rect 40 3272 72 3304
rect 112 3272 144 3304
rect 184 3272 216 3304
rect 256 3272 288 3304
rect 328 3272 360 3304
rect 40 3200 72 3232
rect 112 3200 144 3232
rect 184 3200 216 3232
rect 256 3200 288 3232
rect 328 3200 360 3232
rect 40 3128 72 3160
rect 112 3128 144 3160
rect 184 3128 216 3160
rect 256 3128 288 3160
rect 328 3128 360 3160
rect 40 3056 72 3088
rect 112 3056 144 3088
rect 184 3056 216 3088
rect 256 3056 288 3088
rect 328 3056 360 3088
rect 40 2984 72 3016
rect 112 2984 144 3016
rect 184 2984 216 3016
rect 256 2984 288 3016
rect 328 2984 360 3016
rect 40 2912 72 2944
rect 112 2912 144 2944
rect 184 2912 216 2944
rect 256 2912 288 2944
rect 328 2912 360 2944
rect 40 2840 72 2872
rect 112 2840 144 2872
rect 184 2840 216 2872
rect 256 2840 288 2872
rect 328 2840 360 2872
rect 40 2768 72 2800
rect 112 2768 144 2800
rect 184 2768 216 2800
rect 256 2768 288 2800
rect 328 2768 360 2800
rect 40 2696 72 2728
rect 112 2696 144 2728
rect 184 2696 216 2728
rect 256 2696 288 2728
rect 328 2696 360 2728
rect 40 2624 72 2656
rect 112 2624 144 2656
rect 184 2624 216 2656
rect 256 2624 288 2656
rect 328 2624 360 2656
rect 40 2552 72 2584
rect 112 2552 144 2584
rect 184 2552 216 2584
rect 256 2552 288 2584
rect 328 2552 360 2584
rect 40 2480 72 2512
rect 112 2480 144 2512
rect 184 2480 216 2512
rect 256 2480 288 2512
rect 328 2480 360 2512
rect 40 2408 72 2440
rect 112 2408 144 2440
rect 184 2408 216 2440
rect 256 2408 288 2440
rect 328 2408 360 2440
rect 40 2336 72 2368
rect 112 2336 144 2368
rect 184 2336 216 2368
rect 256 2336 288 2368
rect 328 2336 360 2368
rect 40 2264 72 2296
rect 112 2264 144 2296
rect 184 2264 216 2296
rect 256 2264 288 2296
rect 328 2264 360 2296
rect 40 2192 72 2224
rect 112 2192 144 2224
rect 184 2192 216 2224
rect 256 2192 288 2224
rect 328 2192 360 2224
rect 40 2120 72 2152
rect 112 2120 144 2152
rect 184 2120 216 2152
rect 256 2120 288 2152
rect 328 2120 360 2152
rect 40 2048 72 2080
rect 112 2048 144 2080
rect 184 2048 216 2080
rect 256 2048 288 2080
rect 328 2048 360 2080
rect 40 1976 72 2008
rect 112 1976 144 2008
rect 184 1976 216 2008
rect 256 1976 288 2008
rect 328 1976 360 2008
rect 40 1904 72 1936
rect 112 1904 144 1936
rect 184 1904 216 1936
rect 256 1904 288 1936
rect 328 1904 360 1936
rect 40 1832 72 1864
rect 112 1832 144 1864
rect 184 1832 216 1864
rect 256 1832 288 1864
rect 328 1832 360 1864
rect 40 1760 72 1792
rect 112 1760 144 1792
rect 184 1760 216 1792
rect 256 1760 288 1792
rect 328 1760 360 1792
rect 40 1688 72 1720
rect 112 1688 144 1720
rect 184 1688 216 1720
rect 256 1688 288 1720
rect 328 1688 360 1720
rect 40 1616 72 1648
rect 112 1616 144 1648
rect 184 1616 216 1648
rect 256 1616 288 1648
rect 328 1616 360 1648
rect 40 1544 72 1576
rect 112 1544 144 1576
rect 184 1544 216 1576
rect 256 1544 288 1576
rect 328 1544 360 1576
rect 40 1472 72 1504
rect 112 1472 144 1504
rect 184 1472 216 1504
rect 256 1472 288 1504
rect 328 1472 360 1504
rect 40 1400 72 1432
rect 112 1400 144 1432
rect 184 1400 216 1432
rect 256 1400 288 1432
rect 328 1400 360 1432
rect 40 1328 72 1360
rect 112 1328 144 1360
rect 184 1328 216 1360
rect 256 1328 288 1360
rect 328 1328 360 1360
rect 40 1256 72 1288
rect 112 1256 144 1288
rect 184 1256 216 1288
rect 256 1256 288 1288
rect 328 1256 360 1288
rect 0 33416 400 33430
rect 0 33384 112 33416
rect 144 33384 184 33416
rect 216 33384 256 33416
rect 288 33384 400 33416
rect 0 33370 400 33384
rect 0 29716 400 29730
rect 0 29684 112 29716
rect 144 29684 184 29716
rect 216 29684 256 29716
rect 288 29684 400 29716
rect 0 29670 400 29684
rect 0 12144 400 12200
rect 0 12112 40 12144
rect 72 12112 112 12144
rect 144 12112 184 12144
rect 216 12112 256 12144
rect 288 12112 328 12144
rect 360 12112 400 12144
rect 0 12072 400 12112
rect 0 12040 40 12072
rect 72 12040 112 12072
rect 144 12040 184 12072
rect 216 12040 256 12072
rect 288 12040 328 12072
rect 360 12040 400 12072
rect 0 12000 400 12040
rect 0 11968 40 12000
rect 72 11968 112 12000
rect 144 11968 184 12000
rect 216 11968 256 12000
rect 288 11968 328 12000
rect 360 11968 400 12000
rect 0 11928 400 11968
rect 0 11896 40 11928
rect 72 11896 112 11928
rect 144 11896 184 11928
rect 216 11896 256 11928
rect 288 11896 328 11928
rect 360 11896 400 11928
rect 0 11856 400 11896
rect 0 11824 40 11856
rect 72 11824 112 11856
rect 144 11824 184 11856
rect 216 11824 256 11856
rect 288 11824 328 11856
rect 360 11824 400 11856
rect 0 11784 400 11824
rect 0 11752 40 11784
rect 72 11752 112 11784
rect 144 11752 184 11784
rect 216 11752 256 11784
rect 288 11752 328 11784
rect 360 11752 400 11784
rect 0 11712 400 11752
rect 0 11680 40 11712
rect 72 11680 112 11712
rect 144 11680 184 11712
rect 216 11680 256 11712
rect 288 11680 328 11712
rect 360 11680 400 11712
rect 0 11640 400 11680
rect 0 11608 40 11640
rect 72 11608 112 11640
rect 144 11608 184 11640
rect 216 11608 256 11640
rect 288 11608 328 11640
rect 360 11608 400 11640
rect 0 11568 400 11608
rect 0 11536 40 11568
rect 72 11536 112 11568
rect 144 11536 184 11568
rect 216 11536 256 11568
rect 288 11536 328 11568
rect 360 11536 400 11568
rect 0 11496 400 11536
rect 0 11464 40 11496
rect 72 11464 112 11496
rect 144 11464 184 11496
rect 216 11464 256 11496
rect 288 11464 328 11496
rect 360 11464 400 11496
rect 0 11424 400 11464
rect 0 11392 40 11424
rect 72 11392 112 11424
rect 144 11392 184 11424
rect 216 11392 256 11424
rect 288 11392 328 11424
rect 360 11392 400 11424
rect 0 11352 400 11392
rect 0 11320 40 11352
rect 72 11320 112 11352
rect 144 11320 184 11352
rect 216 11320 256 11352
rect 288 11320 328 11352
rect 360 11320 400 11352
rect 0 11280 400 11320
rect 0 11248 40 11280
rect 72 11248 112 11280
rect 144 11248 184 11280
rect 216 11248 256 11280
rect 288 11248 328 11280
rect 360 11248 400 11280
rect 0 11208 400 11248
rect 0 11176 40 11208
rect 72 11176 112 11208
rect 144 11176 184 11208
rect 216 11176 256 11208
rect 288 11176 328 11208
rect 360 11176 400 11208
rect 0 11136 400 11176
rect 0 11104 40 11136
rect 72 11104 112 11136
rect 144 11104 184 11136
rect 216 11104 256 11136
rect 288 11104 328 11136
rect 360 11104 400 11136
rect 0 11064 400 11104
rect 0 11032 40 11064
rect 72 11032 112 11064
rect 144 11032 184 11064
rect 216 11032 256 11064
rect 288 11032 328 11064
rect 360 11032 400 11064
rect 0 10992 400 11032
rect 0 10960 40 10992
rect 72 10960 112 10992
rect 144 10960 184 10992
rect 216 10960 256 10992
rect 288 10960 328 10992
rect 360 10960 400 10992
rect 0 10920 400 10960
rect 0 10888 40 10920
rect 72 10888 112 10920
rect 144 10888 184 10920
rect 216 10888 256 10920
rect 288 10888 328 10920
rect 360 10888 400 10920
rect 0 10848 400 10888
rect 0 10816 40 10848
rect 72 10816 112 10848
rect 144 10816 184 10848
rect 216 10816 256 10848
rect 288 10816 328 10848
rect 360 10816 400 10848
rect 0 10776 400 10816
rect 0 10744 40 10776
rect 72 10744 112 10776
rect 144 10744 184 10776
rect 216 10744 256 10776
rect 288 10744 328 10776
rect 360 10744 400 10776
rect 0 10704 400 10744
rect 0 10672 40 10704
rect 72 10672 112 10704
rect 144 10672 184 10704
rect 216 10672 256 10704
rect 288 10672 328 10704
rect 360 10672 400 10704
rect 0 10632 400 10672
rect 0 10600 40 10632
rect 72 10600 112 10632
rect 144 10600 184 10632
rect 216 10600 256 10632
rect 288 10600 328 10632
rect 360 10600 400 10632
rect 0 10560 400 10600
rect 0 10528 40 10560
rect 72 10528 112 10560
rect 144 10528 184 10560
rect 216 10528 256 10560
rect 288 10528 328 10560
rect 360 10528 400 10560
rect 0 10488 400 10528
rect 0 10456 40 10488
rect 72 10456 112 10488
rect 144 10456 184 10488
rect 216 10456 256 10488
rect 288 10456 328 10488
rect 360 10456 400 10488
rect 0 10416 400 10456
rect 0 10384 40 10416
rect 72 10384 112 10416
rect 144 10384 184 10416
rect 216 10384 256 10416
rect 288 10384 328 10416
rect 360 10384 400 10416
rect 0 10344 400 10384
rect 0 10312 40 10344
rect 72 10312 112 10344
rect 144 10312 184 10344
rect 216 10312 256 10344
rect 288 10312 328 10344
rect 360 10312 400 10344
rect 0 10272 400 10312
rect 0 10240 40 10272
rect 72 10240 112 10272
rect 144 10240 184 10272
rect 216 10240 256 10272
rect 288 10240 328 10272
rect 360 10240 400 10272
rect 0 10200 400 10240
rect 0 10168 40 10200
rect 72 10168 112 10200
rect 144 10168 184 10200
rect 216 10168 256 10200
rect 288 10168 328 10200
rect 360 10168 400 10200
rect 0 10128 400 10168
rect 0 10096 40 10128
rect 72 10096 112 10128
rect 144 10096 184 10128
rect 216 10096 256 10128
rect 288 10096 328 10128
rect 360 10096 400 10128
rect 0 10056 400 10096
rect 0 10024 40 10056
rect 72 10024 112 10056
rect 144 10024 184 10056
rect 216 10024 256 10056
rect 288 10024 328 10056
rect 360 10024 400 10056
rect 0 9984 400 10024
rect 0 9952 40 9984
rect 72 9952 112 9984
rect 144 9952 184 9984
rect 216 9952 256 9984
rect 288 9952 328 9984
rect 360 9952 400 9984
rect 0 9912 400 9952
rect 0 9880 40 9912
rect 72 9880 112 9912
rect 144 9880 184 9912
rect 216 9880 256 9912
rect 288 9880 328 9912
rect 360 9880 400 9912
rect 0 9840 400 9880
rect 0 9808 40 9840
rect 72 9808 112 9840
rect 144 9808 184 9840
rect 216 9808 256 9840
rect 288 9808 328 9840
rect 360 9808 400 9840
rect 0 9768 400 9808
rect 0 9736 40 9768
rect 72 9736 112 9768
rect 144 9736 184 9768
rect 216 9736 256 9768
rect 288 9736 328 9768
rect 360 9736 400 9768
rect 0 9696 400 9736
rect 0 9664 40 9696
rect 72 9664 112 9696
rect 144 9664 184 9696
rect 216 9664 256 9696
rect 288 9664 328 9696
rect 360 9664 400 9696
rect 0 9624 400 9664
rect 0 9592 40 9624
rect 72 9592 112 9624
rect 144 9592 184 9624
rect 216 9592 256 9624
rect 288 9592 328 9624
rect 360 9592 400 9624
rect 0 9552 400 9592
rect 0 9520 40 9552
rect 72 9520 112 9552
rect 144 9520 184 9552
rect 216 9520 256 9552
rect 288 9520 328 9552
rect 360 9520 400 9552
rect 0 9480 400 9520
rect 0 9448 40 9480
rect 72 9448 112 9480
rect 144 9448 184 9480
rect 216 9448 256 9480
rect 288 9448 328 9480
rect 360 9448 400 9480
rect 0 9408 400 9448
rect 0 9376 40 9408
rect 72 9376 112 9408
rect 144 9376 184 9408
rect 216 9376 256 9408
rect 288 9376 328 9408
rect 360 9376 400 9408
rect 0 9336 400 9376
rect 0 9304 40 9336
rect 72 9304 112 9336
rect 144 9304 184 9336
rect 216 9304 256 9336
rect 288 9304 328 9336
rect 360 9304 400 9336
rect 0 9264 400 9304
rect 0 9232 40 9264
rect 72 9232 112 9264
rect 144 9232 184 9264
rect 216 9232 256 9264
rect 288 9232 328 9264
rect 360 9232 400 9264
rect 0 9192 400 9232
rect 0 9160 40 9192
rect 72 9160 112 9192
rect 144 9160 184 9192
rect 216 9160 256 9192
rect 288 9160 328 9192
rect 360 9160 400 9192
rect 0 9120 400 9160
rect 0 9088 40 9120
rect 72 9088 112 9120
rect 144 9088 184 9120
rect 216 9088 256 9120
rect 288 9088 328 9120
rect 360 9088 400 9120
rect 0 9048 400 9088
rect 0 9016 40 9048
rect 72 9016 112 9048
rect 144 9016 184 9048
rect 216 9016 256 9048
rect 288 9016 328 9048
rect 360 9016 400 9048
rect 0 8976 400 9016
rect 0 8944 40 8976
rect 72 8944 112 8976
rect 144 8944 184 8976
rect 216 8944 256 8976
rect 288 8944 328 8976
rect 360 8944 400 8976
rect 0 8904 400 8944
rect 0 8872 40 8904
rect 72 8872 112 8904
rect 144 8872 184 8904
rect 216 8872 256 8904
rect 288 8872 328 8904
rect 360 8872 400 8904
rect 0 8832 400 8872
rect 0 8800 40 8832
rect 72 8800 112 8832
rect 144 8800 184 8832
rect 216 8800 256 8832
rect 288 8800 328 8832
rect 360 8800 400 8832
rect 0 8760 400 8800
rect 0 8728 40 8760
rect 72 8728 112 8760
rect 144 8728 184 8760
rect 216 8728 256 8760
rect 288 8728 328 8760
rect 360 8728 400 8760
rect 0 8688 400 8728
rect 0 8656 40 8688
rect 72 8656 112 8688
rect 144 8656 184 8688
rect 216 8656 256 8688
rect 288 8656 328 8688
rect 360 8656 400 8688
rect 0 8616 400 8656
rect 0 8584 40 8616
rect 72 8584 112 8616
rect 144 8584 184 8616
rect 216 8584 256 8616
rect 288 8584 328 8616
rect 360 8584 400 8616
rect 0 8544 400 8584
rect 0 8512 40 8544
rect 72 8512 112 8544
rect 144 8512 184 8544
rect 216 8512 256 8544
rect 288 8512 328 8544
rect 360 8512 400 8544
rect 0 8472 400 8512
rect 0 8440 40 8472
rect 72 8440 112 8472
rect 144 8440 184 8472
rect 216 8440 256 8472
rect 288 8440 328 8472
rect 360 8440 400 8472
rect 0 8400 400 8440
rect 0 8368 40 8400
rect 72 8368 112 8400
rect 144 8368 184 8400
rect 216 8368 256 8400
rect 288 8368 328 8400
rect 360 8368 400 8400
rect 0 8328 400 8368
rect 0 8296 40 8328
rect 72 8296 112 8328
rect 144 8296 184 8328
rect 216 8296 256 8328
rect 288 8296 328 8328
rect 360 8296 400 8328
rect 0 8256 400 8296
rect 0 8224 40 8256
rect 72 8224 112 8256
rect 144 8224 184 8256
rect 216 8224 256 8256
rect 288 8224 328 8256
rect 360 8224 400 8256
rect 0 8184 400 8224
rect 0 8152 40 8184
rect 72 8152 112 8184
rect 144 8152 184 8184
rect 216 8152 256 8184
rect 288 8152 328 8184
rect 360 8152 400 8184
rect 0 8112 400 8152
rect 0 8080 40 8112
rect 72 8080 112 8112
rect 144 8080 184 8112
rect 216 8080 256 8112
rect 288 8080 328 8112
rect 360 8080 400 8112
rect 0 8040 400 8080
rect 0 8008 40 8040
rect 72 8008 112 8040
rect 144 8008 184 8040
rect 216 8008 256 8040
rect 288 8008 328 8040
rect 360 8008 400 8040
rect 0 7968 400 8008
rect 0 7936 40 7968
rect 72 7936 112 7968
rect 144 7936 184 7968
rect 216 7936 256 7968
rect 288 7936 328 7968
rect 360 7936 400 7968
rect 0 7896 400 7936
rect 0 7864 40 7896
rect 72 7864 112 7896
rect 144 7864 184 7896
rect 216 7864 256 7896
rect 288 7864 328 7896
rect 360 7864 400 7896
rect 0 7824 400 7864
rect 0 7792 40 7824
rect 72 7792 112 7824
rect 144 7792 184 7824
rect 216 7792 256 7824
rect 288 7792 328 7824
rect 360 7792 400 7824
rect 0 7752 400 7792
rect 0 7720 40 7752
rect 72 7720 112 7752
rect 144 7720 184 7752
rect 216 7720 256 7752
rect 288 7720 328 7752
rect 360 7720 400 7752
rect 0 7680 400 7720
rect 0 7648 40 7680
rect 72 7648 112 7680
rect 144 7648 184 7680
rect 216 7648 256 7680
rect 288 7648 328 7680
rect 360 7648 400 7680
rect 0 7608 400 7648
rect 0 7576 40 7608
rect 72 7576 112 7608
rect 144 7576 184 7608
rect 216 7576 256 7608
rect 288 7576 328 7608
rect 360 7576 400 7608
rect 0 7536 400 7576
rect 0 7504 40 7536
rect 72 7504 112 7536
rect 144 7504 184 7536
rect 216 7504 256 7536
rect 288 7504 328 7536
rect 360 7504 400 7536
rect 0 7464 400 7504
rect 0 7432 40 7464
rect 72 7432 112 7464
rect 144 7432 184 7464
rect 216 7432 256 7464
rect 288 7432 328 7464
rect 360 7432 400 7464
rect 0 7392 400 7432
rect 0 7360 40 7392
rect 72 7360 112 7392
rect 144 7360 184 7392
rect 216 7360 256 7392
rect 288 7360 328 7392
rect 360 7360 400 7392
rect 0 7320 400 7360
rect 0 7288 40 7320
rect 72 7288 112 7320
rect 144 7288 184 7320
rect 216 7288 256 7320
rect 288 7288 328 7320
rect 360 7288 400 7320
rect 0 7248 400 7288
rect 0 7216 40 7248
rect 72 7216 112 7248
rect 144 7216 184 7248
rect 216 7216 256 7248
rect 288 7216 328 7248
rect 360 7216 400 7248
rect 0 7176 400 7216
rect 0 7144 40 7176
rect 72 7144 112 7176
rect 144 7144 184 7176
rect 216 7144 256 7176
rect 288 7144 328 7176
rect 360 7144 400 7176
rect 0 7104 400 7144
rect 0 7072 40 7104
rect 72 7072 112 7104
rect 144 7072 184 7104
rect 216 7072 256 7104
rect 288 7072 328 7104
rect 360 7072 400 7104
rect 0 7032 400 7072
rect 0 7000 40 7032
rect 72 7000 112 7032
rect 144 7000 184 7032
rect 216 7000 256 7032
rect 288 7000 328 7032
rect 360 7000 400 7032
rect 0 6960 400 7000
rect 0 6928 40 6960
rect 72 6928 112 6960
rect 144 6928 184 6960
rect 216 6928 256 6960
rect 288 6928 328 6960
rect 360 6928 400 6960
rect 0 6888 400 6928
rect 0 6856 40 6888
rect 72 6856 112 6888
rect 144 6856 184 6888
rect 216 6856 256 6888
rect 288 6856 328 6888
rect 360 6856 400 6888
rect 0 6800 400 6856
rect 0 6544 400 6600
rect 0 6512 40 6544
rect 72 6512 112 6544
rect 144 6512 184 6544
rect 216 6512 256 6544
rect 288 6512 328 6544
rect 360 6512 400 6544
rect 0 6472 400 6512
rect 0 6440 40 6472
rect 72 6440 112 6472
rect 144 6440 184 6472
rect 216 6440 256 6472
rect 288 6440 328 6472
rect 360 6440 400 6472
rect 0 6400 400 6440
rect 0 6368 40 6400
rect 72 6368 112 6400
rect 144 6368 184 6400
rect 216 6368 256 6400
rect 288 6368 328 6400
rect 360 6368 400 6400
rect 0 6328 400 6368
rect 0 6296 40 6328
rect 72 6296 112 6328
rect 144 6296 184 6328
rect 216 6296 256 6328
rect 288 6296 328 6328
rect 360 6296 400 6328
rect 0 6256 400 6296
rect 0 6224 40 6256
rect 72 6224 112 6256
rect 144 6224 184 6256
rect 216 6224 256 6256
rect 288 6224 328 6256
rect 360 6224 400 6256
rect 0 6184 400 6224
rect 0 6152 40 6184
rect 72 6152 112 6184
rect 144 6152 184 6184
rect 216 6152 256 6184
rect 288 6152 328 6184
rect 360 6152 400 6184
rect 0 6112 400 6152
rect 0 6080 40 6112
rect 72 6080 112 6112
rect 144 6080 184 6112
rect 216 6080 256 6112
rect 288 6080 328 6112
rect 360 6080 400 6112
rect 0 6040 400 6080
rect 0 6008 40 6040
rect 72 6008 112 6040
rect 144 6008 184 6040
rect 216 6008 256 6040
rect 288 6008 328 6040
rect 360 6008 400 6040
rect 0 5968 400 6008
rect 0 5936 40 5968
rect 72 5936 112 5968
rect 144 5936 184 5968
rect 216 5936 256 5968
rect 288 5936 328 5968
rect 360 5936 400 5968
rect 0 5896 400 5936
rect 0 5864 40 5896
rect 72 5864 112 5896
rect 144 5864 184 5896
rect 216 5864 256 5896
rect 288 5864 328 5896
rect 360 5864 400 5896
rect 0 5824 400 5864
rect 0 5792 40 5824
rect 72 5792 112 5824
rect 144 5792 184 5824
rect 216 5792 256 5824
rect 288 5792 328 5824
rect 360 5792 400 5824
rect 0 5752 400 5792
rect 0 5720 40 5752
rect 72 5720 112 5752
rect 144 5720 184 5752
rect 216 5720 256 5752
rect 288 5720 328 5752
rect 360 5720 400 5752
rect 0 5680 400 5720
rect 0 5648 40 5680
rect 72 5648 112 5680
rect 144 5648 184 5680
rect 216 5648 256 5680
rect 288 5648 328 5680
rect 360 5648 400 5680
rect 0 5608 400 5648
rect 0 5576 40 5608
rect 72 5576 112 5608
rect 144 5576 184 5608
rect 216 5576 256 5608
rect 288 5576 328 5608
rect 360 5576 400 5608
rect 0 5536 400 5576
rect 0 5504 40 5536
rect 72 5504 112 5536
rect 144 5504 184 5536
rect 216 5504 256 5536
rect 288 5504 328 5536
rect 360 5504 400 5536
rect 0 5464 400 5504
rect 0 5432 40 5464
rect 72 5432 112 5464
rect 144 5432 184 5464
rect 216 5432 256 5464
rect 288 5432 328 5464
rect 360 5432 400 5464
rect 0 5392 400 5432
rect 0 5360 40 5392
rect 72 5360 112 5392
rect 144 5360 184 5392
rect 216 5360 256 5392
rect 288 5360 328 5392
rect 360 5360 400 5392
rect 0 5320 400 5360
rect 0 5288 40 5320
rect 72 5288 112 5320
rect 144 5288 184 5320
rect 216 5288 256 5320
rect 288 5288 328 5320
rect 360 5288 400 5320
rect 0 5248 400 5288
rect 0 5216 40 5248
rect 72 5216 112 5248
rect 144 5216 184 5248
rect 216 5216 256 5248
rect 288 5216 328 5248
rect 360 5216 400 5248
rect 0 5176 400 5216
rect 0 5144 40 5176
rect 72 5144 112 5176
rect 144 5144 184 5176
rect 216 5144 256 5176
rect 288 5144 328 5176
rect 360 5144 400 5176
rect 0 5104 400 5144
rect 0 5072 40 5104
rect 72 5072 112 5104
rect 144 5072 184 5104
rect 216 5072 256 5104
rect 288 5072 328 5104
rect 360 5072 400 5104
rect 0 5032 400 5072
rect 0 5000 40 5032
rect 72 5000 112 5032
rect 144 5000 184 5032
rect 216 5000 256 5032
rect 288 5000 328 5032
rect 360 5000 400 5032
rect 0 4960 400 5000
rect 0 4928 40 4960
rect 72 4928 112 4960
rect 144 4928 184 4960
rect 216 4928 256 4960
rect 288 4928 328 4960
rect 360 4928 400 4960
rect 0 4888 400 4928
rect 0 4856 40 4888
rect 72 4856 112 4888
rect 144 4856 184 4888
rect 216 4856 256 4888
rect 288 4856 328 4888
rect 360 4856 400 4888
rect 0 4816 400 4856
rect 0 4784 40 4816
rect 72 4784 112 4816
rect 144 4784 184 4816
rect 216 4784 256 4816
rect 288 4784 328 4816
rect 360 4784 400 4816
rect 0 4744 400 4784
rect 0 4712 40 4744
rect 72 4712 112 4744
rect 144 4712 184 4744
rect 216 4712 256 4744
rect 288 4712 328 4744
rect 360 4712 400 4744
rect 0 4672 400 4712
rect 0 4640 40 4672
rect 72 4640 112 4672
rect 144 4640 184 4672
rect 216 4640 256 4672
rect 288 4640 328 4672
rect 360 4640 400 4672
rect 0 4600 400 4640
rect 0 4568 40 4600
rect 72 4568 112 4600
rect 144 4568 184 4600
rect 216 4568 256 4600
rect 288 4568 328 4600
rect 360 4568 400 4600
rect 0 4528 400 4568
rect 0 4496 40 4528
rect 72 4496 112 4528
rect 144 4496 184 4528
rect 216 4496 256 4528
rect 288 4496 328 4528
rect 360 4496 400 4528
rect 0 4456 400 4496
rect 0 4424 40 4456
rect 72 4424 112 4456
rect 144 4424 184 4456
rect 216 4424 256 4456
rect 288 4424 328 4456
rect 360 4424 400 4456
rect 0 4384 400 4424
rect 0 4352 40 4384
rect 72 4352 112 4384
rect 144 4352 184 4384
rect 216 4352 256 4384
rect 288 4352 328 4384
rect 360 4352 400 4384
rect 0 4312 400 4352
rect 0 4280 40 4312
rect 72 4280 112 4312
rect 144 4280 184 4312
rect 216 4280 256 4312
rect 288 4280 328 4312
rect 360 4280 400 4312
rect 0 4240 400 4280
rect 0 4208 40 4240
rect 72 4208 112 4240
rect 144 4208 184 4240
rect 216 4208 256 4240
rect 288 4208 328 4240
rect 360 4208 400 4240
rect 0 4168 400 4208
rect 0 4136 40 4168
rect 72 4136 112 4168
rect 144 4136 184 4168
rect 216 4136 256 4168
rect 288 4136 328 4168
rect 360 4136 400 4168
rect 0 4096 400 4136
rect 0 4064 40 4096
rect 72 4064 112 4096
rect 144 4064 184 4096
rect 216 4064 256 4096
rect 288 4064 328 4096
rect 360 4064 400 4096
rect 0 4024 400 4064
rect 0 3992 40 4024
rect 72 3992 112 4024
rect 144 3992 184 4024
rect 216 3992 256 4024
rect 288 3992 328 4024
rect 360 3992 400 4024
rect 0 3952 400 3992
rect 0 3920 40 3952
rect 72 3920 112 3952
rect 144 3920 184 3952
rect 216 3920 256 3952
rect 288 3920 328 3952
rect 360 3920 400 3952
rect 0 3880 400 3920
rect 0 3848 40 3880
rect 72 3848 112 3880
rect 144 3848 184 3880
rect 216 3848 256 3880
rect 288 3848 328 3880
rect 360 3848 400 3880
rect 0 3808 400 3848
rect 0 3776 40 3808
rect 72 3776 112 3808
rect 144 3776 184 3808
rect 216 3776 256 3808
rect 288 3776 328 3808
rect 360 3776 400 3808
rect 0 3736 400 3776
rect 0 3704 40 3736
rect 72 3704 112 3736
rect 144 3704 184 3736
rect 216 3704 256 3736
rect 288 3704 328 3736
rect 360 3704 400 3736
rect 0 3664 400 3704
rect 0 3632 40 3664
rect 72 3632 112 3664
rect 144 3632 184 3664
rect 216 3632 256 3664
rect 288 3632 328 3664
rect 360 3632 400 3664
rect 0 3592 400 3632
rect 0 3560 40 3592
rect 72 3560 112 3592
rect 144 3560 184 3592
rect 216 3560 256 3592
rect 288 3560 328 3592
rect 360 3560 400 3592
rect 0 3520 400 3560
rect 0 3488 40 3520
rect 72 3488 112 3520
rect 144 3488 184 3520
rect 216 3488 256 3520
rect 288 3488 328 3520
rect 360 3488 400 3520
rect 0 3448 400 3488
rect 0 3416 40 3448
rect 72 3416 112 3448
rect 144 3416 184 3448
rect 216 3416 256 3448
rect 288 3416 328 3448
rect 360 3416 400 3448
rect 0 3376 400 3416
rect 0 3344 40 3376
rect 72 3344 112 3376
rect 144 3344 184 3376
rect 216 3344 256 3376
rect 288 3344 328 3376
rect 360 3344 400 3376
rect 0 3304 400 3344
rect 0 3272 40 3304
rect 72 3272 112 3304
rect 144 3272 184 3304
rect 216 3272 256 3304
rect 288 3272 328 3304
rect 360 3272 400 3304
rect 0 3232 400 3272
rect 0 3200 40 3232
rect 72 3200 112 3232
rect 144 3200 184 3232
rect 216 3200 256 3232
rect 288 3200 328 3232
rect 360 3200 400 3232
rect 0 3160 400 3200
rect 0 3128 40 3160
rect 72 3128 112 3160
rect 144 3128 184 3160
rect 216 3128 256 3160
rect 288 3128 328 3160
rect 360 3128 400 3160
rect 0 3088 400 3128
rect 0 3056 40 3088
rect 72 3056 112 3088
rect 144 3056 184 3088
rect 216 3056 256 3088
rect 288 3056 328 3088
rect 360 3056 400 3088
rect 0 3016 400 3056
rect 0 2984 40 3016
rect 72 2984 112 3016
rect 144 2984 184 3016
rect 216 2984 256 3016
rect 288 2984 328 3016
rect 360 2984 400 3016
rect 0 2944 400 2984
rect 0 2912 40 2944
rect 72 2912 112 2944
rect 144 2912 184 2944
rect 216 2912 256 2944
rect 288 2912 328 2944
rect 360 2912 400 2944
rect 0 2872 400 2912
rect 0 2840 40 2872
rect 72 2840 112 2872
rect 144 2840 184 2872
rect 216 2840 256 2872
rect 288 2840 328 2872
rect 360 2840 400 2872
rect 0 2800 400 2840
rect 0 2768 40 2800
rect 72 2768 112 2800
rect 144 2768 184 2800
rect 216 2768 256 2800
rect 288 2768 328 2800
rect 360 2768 400 2800
rect 0 2728 400 2768
rect 0 2696 40 2728
rect 72 2696 112 2728
rect 144 2696 184 2728
rect 216 2696 256 2728
rect 288 2696 328 2728
rect 360 2696 400 2728
rect 0 2656 400 2696
rect 0 2624 40 2656
rect 72 2624 112 2656
rect 144 2624 184 2656
rect 216 2624 256 2656
rect 288 2624 328 2656
rect 360 2624 400 2656
rect 0 2584 400 2624
rect 0 2552 40 2584
rect 72 2552 112 2584
rect 144 2552 184 2584
rect 216 2552 256 2584
rect 288 2552 328 2584
rect 360 2552 400 2584
rect 0 2512 400 2552
rect 0 2480 40 2512
rect 72 2480 112 2512
rect 144 2480 184 2512
rect 216 2480 256 2512
rect 288 2480 328 2512
rect 360 2480 400 2512
rect 0 2440 400 2480
rect 0 2408 40 2440
rect 72 2408 112 2440
rect 144 2408 184 2440
rect 216 2408 256 2440
rect 288 2408 328 2440
rect 360 2408 400 2440
rect 0 2368 400 2408
rect 0 2336 40 2368
rect 72 2336 112 2368
rect 144 2336 184 2368
rect 216 2336 256 2368
rect 288 2336 328 2368
rect 360 2336 400 2368
rect 0 2296 400 2336
rect 0 2264 40 2296
rect 72 2264 112 2296
rect 144 2264 184 2296
rect 216 2264 256 2296
rect 288 2264 328 2296
rect 360 2264 400 2296
rect 0 2224 400 2264
rect 0 2192 40 2224
rect 72 2192 112 2224
rect 144 2192 184 2224
rect 216 2192 256 2224
rect 288 2192 328 2224
rect 360 2192 400 2224
rect 0 2152 400 2192
rect 0 2120 40 2152
rect 72 2120 112 2152
rect 144 2120 184 2152
rect 216 2120 256 2152
rect 288 2120 328 2152
rect 360 2120 400 2152
rect 0 2080 400 2120
rect 0 2048 40 2080
rect 72 2048 112 2080
rect 144 2048 184 2080
rect 216 2048 256 2080
rect 288 2048 328 2080
rect 360 2048 400 2080
rect 0 2008 400 2048
rect 0 1976 40 2008
rect 72 1976 112 2008
rect 144 1976 184 2008
rect 216 1976 256 2008
rect 288 1976 328 2008
rect 360 1976 400 2008
rect 0 1936 400 1976
rect 0 1904 40 1936
rect 72 1904 112 1936
rect 144 1904 184 1936
rect 216 1904 256 1936
rect 288 1904 328 1936
rect 360 1904 400 1936
rect 0 1864 400 1904
rect 0 1832 40 1864
rect 72 1832 112 1864
rect 144 1832 184 1864
rect 216 1832 256 1864
rect 288 1832 328 1864
rect 360 1832 400 1864
rect 0 1792 400 1832
rect 0 1760 40 1792
rect 72 1760 112 1792
rect 144 1760 184 1792
rect 216 1760 256 1792
rect 288 1760 328 1792
rect 360 1760 400 1792
rect 0 1720 400 1760
rect 0 1688 40 1720
rect 72 1688 112 1720
rect 144 1688 184 1720
rect 216 1688 256 1720
rect 288 1688 328 1720
rect 360 1688 400 1720
rect 0 1648 400 1688
rect 0 1616 40 1648
rect 72 1616 112 1648
rect 144 1616 184 1648
rect 216 1616 256 1648
rect 288 1616 328 1648
rect 360 1616 400 1648
rect 0 1576 400 1616
rect 0 1544 40 1576
rect 72 1544 112 1576
rect 144 1544 184 1576
rect 216 1544 256 1576
rect 288 1544 328 1576
rect 360 1544 400 1576
rect 0 1504 400 1544
rect 0 1472 40 1504
rect 72 1472 112 1504
rect 144 1472 184 1504
rect 216 1472 256 1504
rect 288 1472 328 1504
rect 360 1472 400 1504
rect 0 1432 400 1472
rect 0 1400 40 1432
rect 72 1400 112 1432
rect 144 1400 184 1432
rect 216 1400 256 1432
rect 288 1400 328 1432
rect 360 1400 400 1432
rect 0 1360 400 1400
rect 0 1328 40 1360
rect 72 1328 112 1360
rect 144 1328 184 1360
rect 216 1328 256 1360
rect 288 1328 328 1360
rect 360 1328 400 1360
rect 0 1288 400 1328
rect 0 1256 40 1288
rect 72 1256 112 1288
rect 144 1256 184 1288
rect 216 1256 256 1288
rect 288 1256 328 1288
rect 360 1256 400 1288
rect 0 1200 400 1256
<< psubdiffcont >>
rect 184 31452 216 31484
rect 112 27939 144 27971
rect 112 22842 144 22874
rect 112 17816 144 17848
<< nsubdiffcont >>
rect 112 33384 144 33416
rect 112 29684 144 29716
rect 40 12112 72 12144
rect 40 6512 72 6544
<< metal1 >>
rect 184 33384 216 33416
rect 256 33384 288 33416
rect 184 29684 216 29716
rect 256 29684 288 29716
rect 112 12112 144 12144
rect 184 12112 216 12144
rect 256 12112 288 12144
rect 328 12112 360 12144
rect 40 12040 72 12072
rect 112 12040 144 12072
rect 184 12040 216 12072
rect 256 12040 288 12072
rect 328 12040 360 12072
rect 40 11968 72 12000
rect 112 11968 144 12000
rect 184 11968 216 12000
rect 256 11968 288 12000
rect 328 11968 360 12000
rect 40 11896 72 11928
rect 112 11896 144 11928
rect 184 11896 216 11928
rect 256 11896 288 11928
rect 328 11896 360 11928
rect 40 11824 72 11856
rect 112 11824 144 11856
rect 184 11824 216 11856
rect 256 11824 288 11856
rect 328 11824 360 11856
rect 40 11752 72 11784
rect 112 11752 144 11784
rect 184 11752 216 11784
rect 256 11752 288 11784
rect 328 11752 360 11784
rect 40 11680 72 11712
rect 112 11680 144 11712
rect 184 11680 216 11712
rect 256 11680 288 11712
rect 328 11680 360 11712
rect 40 11608 72 11640
rect 112 11608 144 11640
rect 184 11608 216 11640
rect 256 11608 288 11640
rect 328 11608 360 11640
rect 40 11536 72 11568
rect 112 11536 144 11568
rect 184 11536 216 11568
rect 256 11536 288 11568
rect 328 11536 360 11568
rect 40 11464 72 11496
rect 112 11464 144 11496
rect 184 11464 216 11496
rect 256 11464 288 11496
rect 328 11464 360 11496
rect 40 11392 72 11424
rect 112 11392 144 11424
rect 184 11392 216 11424
rect 256 11392 288 11424
rect 328 11392 360 11424
rect 40 11320 72 11352
rect 112 11320 144 11352
rect 184 11320 216 11352
rect 256 11320 288 11352
rect 328 11320 360 11352
rect 40 11248 72 11280
rect 112 11248 144 11280
rect 184 11248 216 11280
rect 256 11248 288 11280
rect 328 11248 360 11280
rect 40 11176 72 11208
rect 112 11176 144 11208
rect 184 11176 216 11208
rect 256 11176 288 11208
rect 328 11176 360 11208
rect 40 11104 72 11136
rect 112 11104 144 11136
rect 184 11104 216 11136
rect 256 11104 288 11136
rect 328 11104 360 11136
rect 40 11032 72 11064
rect 112 11032 144 11064
rect 184 11032 216 11064
rect 256 11032 288 11064
rect 328 11032 360 11064
rect 40 10960 72 10992
rect 112 10960 144 10992
rect 184 10960 216 10992
rect 256 10960 288 10992
rect 328 10960 360 10992
rect 40 10888 72 10920
rect 112 10888 144 10920
rect 184 10888 216 10920
rect 256 10888 288 10920
rect 328 10888 360 10920
rect 40 10816 72 10848
rect 112 10816 144 10848
rect 184 10816 216 10848
rect 256 10816 288 10848
rect 328 10816 360 10848
rect 40 10744 72 10776
rect 112 10744 144 10776
rect 184 10744 216 10776
rect 256 10744 288 10776
rect 328 10744 360 10776
rect 40 10672 72 10704
rect 112 10672 144 10704
rect 184 10672 216 10704
rect 256 10672 288 10704
rect 328 10672 360 10704
rect 40 10600 72 10632
rect 112 10600 144 10632
rect 184 10600 216 10632
rect 256 10600 288 10632
rect 328 10600 360 10632
rect 40 10528 72 10560
rect 112 10528 144 10560
rect 184 10528 216 10560
rect 256 10528 288 10560
rect 328 10528 360 10560
rect 40 10456 72 10488
rect 112 10456 144 10488
rect 184 10456 216 10488
rect 256 10456 288 10488
rect 328 10456 360 10488
rect 40 10384 72 10416
rect 112 10384 144 10416
rect 184 10384 216 10416
rect 256 10384 288 10416
rect 328 10384 360 10416
rect 40 10312 72 10344
rect 112 10312 144 10344
rect 184 10312 216 10344
rect 256 10312 288 10344
rect 328 10312 360 10344
rect 40 10240 72 10272
rect 112 10240 144 10272
rect 184 10240 216 10272
rect 256 10240 288 10272
rect 328 10240 360 10272
rect 40 10168 72 10200
rect 112 10168 144 10200
rect 184 10168 216 10200
rect 256 10168 288 10200
rect 328 10168 360 10200
rect 40 10096 72 10128
rect 112 10096 144 10128
rect 184 10096 216 10128
rect 256 10096 288 10128
rect 328 10096 360 10128
rect 40 10024 72 10056
rect 112 10024 144 10056
rect 184 10024 216 10056
rect 256 10024 288 10056
rect 328 10024 360 10056
rect 40 9952 72 9984
rect 112 9952 144 9984
rect 184 9952 216 9984
rect 256 9952 288 9984
rect 328 9952 360 9984
rect 40 9880 72 9912
rect 112 9880 144 9912
rect 184 9880 216 9912
rect 256 9880 288 9912
rect 328 9880 360 9912
rect 40 9808 72 9840
rect 112 9808 144 9840
rect 184 9808 216 9840
rect 256 9808 288 9840
rect 328 9808 360 9840
rect 40 9736 72 9768
rect 112 9736 144 9768
rect 184 9736 216 9768
rect 256 9736 288 9768
rect 328 9736 360 9768
rect 40 9664 72 9696
rect 112 9664 144 9696
rect 184 9664 216 9696
rect 256 9664 288 9696
rect 328 9664 360 9696
rect 40 9592 72 9624
rect 112 9592 144 9624
rect 184 9592 216 9624
rect 256 9592 288 9624
rect 328 9592 360 9624
rect 40 9520 72 9552
rect 112 9520 144 9552
rect 184 9520 216 9552
rect 256 9520 288 9552
rect 328 9520 360 9552
rect 40 9448 72 9480
rect 112 9448 144 9480
rect 184 9448 216 9480
rect 256 9448 288 9480
rect 328 9448 360 9480
rect 40 9376 72 9408
rect 112 9376 144 9408
rect 184 9376 216 9408
rect 256 9376 288 9408
rect 328 9376 360 9408
rect 40 9304 72 9336
rect 112 9304 144 9336
rect 184 9304 216 9336
rect 256 9304 288 9336
rect 328 9304 360 9336
rect 40 9232 72 9264
rect 112 9232 144 9264
rect 184 9232 216 9264
rect 256 9232 288 9264
rect 328 9232 360 9264
rect 40 9160 72 9192
rect 112 9160 144 9192
rect 184 9160 216 9192
rect 256 9160 288 9192
rect 328 9160 360 9192
rect 40 9088 72 9120
rect 112 9088 144 9120
rect 184 9088 216 9120
rect 256 9088 288 9120
rect 328 9088 360 9120
rect 40 9016 72 9048
rect 112 9016 144 9048
rect 184 9016 216 9048
rect 256 9016 288 9048
rect 328 9016 360 9048
rect 40 8944 72 8976
rect 112 8944 144 8976
rect 184 8944 216 8976
rect 256 8944 288 8976
rect 328 8944 360 8976
rect 40 8872 72 8904
rect 112 8872 144 8904
rect 184 8872 216 8904
rect 256 8872 288 8904
rect 328 8872 360 8904
rect 40 8800 72 8832
rect 112 8800 144 8832
rect 184 8800 216 8832
rect 256 8800 288 8832
rect 328 8800 360 8832
rect 40 8728 72 8760
rect 112 8728 144 8760
rect 184 8728 216 8760
rect 256 8728 288 8760
rect 328 8728 360 8760
rect 40 8656 72 8688
rect 112 8656 144 8688
rect 184 8656 216 8688
rect 256 8656 288 8688
rect 328 8656 360 8688
rect 40 8584 72 8616
rect 112 8584 144 8616
rect 184 8584 216 8616
rect 256 8584 288 8616
rect 328 8584 360 8616
rect 40 8512 72 8544
rect 112 8512 144 8544
rect 184 8512 216 8544
rect 256 8512 288 8544
rect 328 8512 360 8544
rect 40 8440 72 8472
rect 112 8440 144 8472
rect 184 8440 216 8472
rect 256 8440 288 8472
rect 328 8440 360 8472
rect 40 8368 72 8400
rect 112 8368 144 8400
rect 184 8368 216 8400
rect 256 8368 288 8400
rect 328 8368 360 8400
rect 40 8296 72 8328
rect 112 8296 144 8328
rect 184 8296 216 8328
rect 256 8296 288 8328
rect 328 8296 360 8328
rect 40 8224 72 8256
rect 112 8224 144 8256
rect 184 8224 216 8256
rect 256 8224 288 8256
rect 328 8224 360 8256
rect 40 8152 72 8184
rect 112 8152 144 8184
rect 184 8152 216 8184
rect 256 8152 288 8184
rect 328 8152 360 8184
rect 40 8080 72 8112
rect 112 8080 144 8112
rect 184 8080 216 8112
rect 256 8080 288 8112
rect 328 8080 360 8112
rect 40 8008 72 8040
rect 112 8008 144 8040
rect 184 8008 216 8040
rect 256 8008 288 8040
rect 328 8008 360 8040
rect 40 7936 72 7968
rect 112 7936 144 7968
rect 184 7936 216 7968
rect 256 7936 288 7968
rect 328 7936 360 7968
rect 40 7864 72 7896
rect 112 7864 144 7896
rect 184 7864 216 7896
rect 256 7864 288 7896
rect 328 7864 360 7896
rect 40 7792 72 7824
rect 112 7792 144 7824
rect 184 7792 216 7824
rect 256 7792 288 7824
rect 328 7792 360 7824
rect 40 7720 72 7752
rect 112 7720 144 7752
rect 184 7720 216 7752
rect 256 7720 288 7752
rect 328 7720 360 7752
rect 40 7648 72 7680
rect 112 7648 144 7680
rect 184 7648 216 7680
rect 256 7648 288 7680
rect 328 7648 360 7680
rect 40 7576 72 7608
rect 112 7576 144 7608
rect 184 7576 216 7608
rect 256 7576 288 7608
rect 328 7576 360 7608
rect 40 7504 72 7536
rect 112 7504 144 7536
rect 184 7504 216 7536
rect 256 7504 288 7536
rect 328 7504 360 7536
rect 40 7432 72 7464
rect 112 7432 144 7464
rect 184 7432 216 7464
rect 256 7432 288 7464
rect 328 7432 360 7464
rect 40 7360 72 7392
rect 112 7360 144 7392
rect 184 7360 216 7392
rect 256 7360 288 7392
rect 328 7360 360 7392
rect 40 7288 72 7320
rect 112 7288 144 7320
rect 184 7288 216 7320
rect 256 7288 288 7320
rect 328 7288 360 7320
rect 40 7216 72 7248
rect 112 7216 144 7248
rect 184 7216 216 7248
rect 256 7216 288 7248
rect 328 7216 360 7248
rect 40 7144 72 7176
rect 112 7144 144 7176
rect 184 7144 216 7176
rect 256 7144 288 7176
rect 328 7144 360 7176
rect 40 7072 72 7104
rect 112 7072 144 7104
rect 184 7072 216 7104
rect 256 7072 288 7104
rect 328 7072 360 7104
rect 40 7000 72 7032
rect 112 7000 144 7032
rect 184 7000 216 7032
rect 256 7000 288 7032
rect 328 7000 360 7032
rect 40 6928 72 6960
rect 112 6928 144 6960
rect 184 6928 216 6960
rect 256 6928 288 6960
rect 328 6928 360 6960
rect 40 6856 72 6888
rect 112 6856 144 6888
rect 184 6856 216 6888
rect 256 6856 288 6888
rect 328 6856 360 6888
rect 112 6512 144 6544
rect 184 6512 216 6544
rect 256 6512 288 6544
rect 328 6512 360 6544
rect 40 6440 72 6472
rect 112 6440 144 6472
rect 184 6440 216 6472
rect 256 6440 288 6472
rect 328 6440 360 6472
rect 40 6368 72 6400
rect 112 6368 144 6400
rect 184 6368 216 6400
rect 256 6368 288 6400
rect 328 6368 360 6400
rect 40 6296 72 6328
rect 112 6296 144 6328
rect 184 6296 216 6328
rect 256 6296 288 6328
rect 328 6296 360 6328
rect 40 6224 72 6256
rect 112 6224 144 6256
rect 184 6224 216 6256
rect 256 6224 288 6256
rect 328 6224 360 6256
rect 40 6152 72 6184
rect 112 6152 144 6184
rect 184 6152 216 6184
rect 256 6152 288 6184
rect 328 6152 360 6184
rect 40 6080 72 6112
rect 112 6080 144 6112
rect 184 6080 216 6112
rect 256 6080 288 6112
rect 328 6080 360 6112
rect 40 6008 72 6040
rect 112 6008 144 6040
rect 184 6008 216 6040
rect 256 6008 288 6040
rect 328 6008 360 6040
rect 40 5936 72 5968
rect 112 5936 144 5968
rect 184 5936 216 5968
rect 256 5936 288 5968
rect 328 5936 360 5968
rect 40 5864 72 5896
rect 112 5864 144 5896
rect 184 5864 216 5896
rect 256 5864 288 5896
rect 328 5864 360 5896
rect 40 5792 72 5824
rect 112 5792 144 5824
rect 184 5792 216 5824
rect 256 5792 288 5824
rect 328 5792 360 5824
rect 40 5720 72 5752
rect 112 5720 144 5752
rect 184 5720 216 5752
rect 256 5720 288 5752
rect 328 5720 360 5752
rect 40 5648 72 5680
rect 112 5648 144 5680
rect 184 5648 216 5680
rect 256 5648 288 5680
rect 328 5648 360 5680
rect 40 5576 72 5608
rect 112 5576 144 5608
rect 184 5576 216 5608
rect 256 5576 288 5608
rect 328 5576 360 5608
rect 40 5504 72 5536
rect 112 5504 144 5536
rect 184 5504 216 5536
rect 256 5504 288 5536
rect 328 5504 360 5536
rect 40 5432 72 5464
rect 112 5432 144 5464
rect 184 5432 216 5464
rect 256 5432 288 5464
rect 328 5432 360 5464
rect 40 5360 72 5392
rect 112 5360 144 5392
rect 184 5360 216 5392
rect 256 5360 288 5392
rect 328 5360 360 5392
rect 40 5288 72 5320
rect 112 5288 144 5320
rect 184 5288 216 5320
rect 256 5288 288 5320
rect 328 5288 360 5320
rect 40 5216 72 5248
rect 112 5216 144 5248
rect 184 5216 216 5248
rect 256 5216 288 5248
rect 328 5216 360 5248
rect 40 5144 72 5176
rect 112 5144 144 5176
rect 184 5144 216 5176
rect 256 5144 288 5176
rect 328 5144 360 5176
rect 40 5072 72 5104
rect 112 5072 144 5104
rect 184 5072 216 5104
rect 256 5072 288 5104
rect 328 5072 360 5104
rect 40 5000 72 5032
rect 112 5000 144 5032
rect 184 5000 216 5032
rect 256 5000 288 5032
rect 328 5000 360 5032
rect 40 4928 72 4960
rect 112 4928 144 4960
rect 184 4928 216 4960
rect 256 4928 288 4960
rect 328 4928 360 4960
rect 40 4856 72 4888
rect 112 4856 144 4888
rect 184 4856 216 4888
rect 256 4856 288 4888
rect 328 4856 360 4888
rect 40 4784 72 4816
rect 112 4784 144 4816
rect 184 4784 216 4816
rect 256 4784 288 4816
rect 328 4784 360 4816
rect 40 4712 72 4744
rect 112 4712 144 4744
rect 184 4712 216 4744
rect 256 4712 288 4744
rect 328 4712 360 4744
rect 40 4640 72 4672
rect 112 4640 144 4672
rect 184 4640 216 4672
rect 256 4640 288 4672
rect 328 4640 360 4672
rect 40 4568 72 4600
rect 112 4568 144 4600
rect 184 4568 216 4600
rect 256 4568 288 4600
rect 328 4568 360 4600
rect 40 4496 72 4528
rect 112 4496 144 4528
rect 184 4496 216 4528
rect 256 4496 288 4528
rect 328 4496 360 4528
rect 40 4424 72 4456
rect 112 4424 144 4456
rect 184 4424 216 4456
rect 256 4424 288 4456
rect 328 4424 360 4456
rect 40 4352 72 4384
rect 112 4352 144 4384
rect 184 4352 216 4384
rect 256 4352 288 4384
rect 328 4352 360 4384
rect 40 4280 72 4312
rect 112 4280 144 4312
rect 184 4280 216 4312
rect 256 4280 288 4312
rect 328 4280 360 4312
rect 40 4208 72 4240
rect 112 4208 144 4240
rect 184 4208 216 4240
rect 256 4208 288 4240
rect 328 4208 360 4240
rect 40 4136 72 4168
rect 112 4136 144 4168
rect 184 4136 216 4168
rect 256 4136 288 4168
rect 328 4136 360 4168
rect 40 4064 72 4096
rect 112 4064 144 4096
rect 184 4064 216 4096
rect 256 4064 288 4096
rect 328 4064 360 4096
rect 40 3992 72 4024
rect 112 3992 144 4024
rect 184 3992 216 4024
rect 256 3992 288 4024
rect 328 3992 360 4024
rect 40 3920 72 3952
rect 112 3920 144 3952
rect 184 3920 216 3952
rect 256 3920 288 3952
rect 328 3920 360 3952
rect 40 3848 72 3880
rect 112 3848 144 3880
rect 184 3848 216 3880
rect 256 3848 288 3880
rect 328 3848 360 3880
rect 40 3776 72 3808
rect 112 3776 144 3808
rect 184 3776 216 3808
rect 256 3776 288 3808
rect 328 3776 360 3808
rect 40 3704 72 3736
rect 112 3704 144 3736
rect 184 3704 216 3736
rect 256 3704 288 3736
rect 328 3704 360 3736
rect 40 3632 72 3664
rect 112 3632 144 3664
rect 184 3632 216 3664
rect 256 3632 288 3664
rect 328 3632 360 3664
rect 40 3560 72 3592
rect 112 3560 144 3592
rect 184 3560 216 3592
rect 256 3560 288 3592
rect 328 3560 360 3592
rect 40 3488 72 3520
rect 112 3488 144 3520
rect 184 3488 216 3520
rect 256 3488 288 3520
rect 328 3488 360 3520
rect 40 3416 72 3448
rect 112 3416 144 3448
rect 184 3416 216 3448
rect 256 3416 288 3448
rect 328 3416 360 3448
rect 40 3344 72 3376
rect 112 3344 144 3376
rect 184 3344 216 3376
rect 256 3344 288 3376
rect 328 3344 360 3376
rect 40 3272 72 3304
rect 112 3272 144 3304
rect 184 3272 216 3304
rect 256 3272 288 3304
rect 328 3272 360 3304
rect 40 3200 72 3232
rect 112 3200 144 3232
rect 184 3200 216 3232
rect 256 3200 288 3232
rect 328 3200 360 3232
rect 40 3128 72 3160
rect 112 3128 144 3160
rect 184 3128 216 3160
rect 256 3128 288 3160
rect 328 3128 360 3160
rect 40 3056 72 3088
rect 112 3056 144 3088
rect 184 3056 216 3088
rect 256 3056 288 3088
rect 328 3056 360 3088
rect 40 2984 72 3016
rect 112 2984 144 3016
rect 184 2984 216 3016
rect 256 2984 288 3016
rect 328 2984 360 3016
rect 40 2912 72 2944
rect 112 2912 144 2944
rect 184 2912 216 2944
rect 256 2912 288 2944
rect 328 2912 360 2944
rect 40 2840 72 2872
rect 112 2840 144 2872
rect 184 2840 216 2872
rect 256 2840 288 2872
rect 328 2840 360 2872
rect 40 2768 72 2800
rect 112 2768 144 2800
rect 184 2768 216 2800
rect 256 2768 288 2800
rect 328 2768 360 2800
rect 40 2696 72 2728
rect 112 2696 144 2728
rect 184 2696 216 2728
rect 256 2696 288 2728
rect 328 2696 360 2728
rect 40 2624 72 2656
rect 112 2624 144 2656
rect 184 2624 216 2656
rect 256 2624 288 2656
rect 328 2624 360 2656
rect 40 2552 72 2584
rect 112 2552 144 2584
rect 184 2552 216 2584
rect 256 2552 288 2584
rect 328 2552 360 2584
rect 40 2480 72 2512
rect 112 2480 144 2512
rect 184 2480 216 2512
rect 256 2480 288 2512
rect 328 2480 360 2512
rect 40 2408 72 2440
rect 112 2408 144 2440
rect 184 2408 216 2440
rect 256 2408 288 2440
rect 328 2408 360 2440
rect 40 2336 72 2368
rect 112 2336 144 2368
rect 184 2336 216 2368
rect 256 2336 288 2368
rect 328 2336 360 2368
rect 40 2264 72 2296
rect 112 2264 144 2296
rect 184 2264 216 2296
rect 256 2264 288 2296
rect 328 2264 360 2296
rect 40 2192 72 2224
rect 112 2192 144 2224
rect 184 2192 216 2224
rect 256 2192 288 2224
rect 328 2192 360 2224
rect 40 2120 72 2152
rect 112 2120 144 2152
rect 184 2120 216 2152
rect 256 2120 288 2152
rect 328 2120 360 2152
rect 40 2048 72 2080
rect 112 2048 144 2080
rect 184 2048 216 2080
rect 256 2048 288 2080
rect 328 2048 360 2080
rect 40 1976 72 2008
rect 112 1976 144 2008
rect 184 1976 216 2008
rect 256 1976 288 2008
rect 328 1976 360 2008
rect 40 1904 72 1936
rect 112 1904 144 1936
rect 184 1904 216 1936
rect 256 1904 288 1936
rect 328 1904 360 1936
rect 40 1832 72 1864
rect 112 1832 144 1864
rect 184 1832 216 1864
rect 256 1832 288 1864
rect 328 1832 360 1864
rect 40 1760 72 1792
rect 112 1760 144 1792
rect 184 1760 216 1792
rect 256 1760 288 1792
rect 328 1760 360 1792
rect 40 1688 72 1720
rect 112 1688 144 1720
rect 184 1688 216 1720
rect 256 1688 288 1720
rect 328 1688 360 1720
rect 40 1616 72 1648
rect 112 1616 144 1648
rect 184 1616 216 1648
rect 256 1616 288 1648
rect 328 1616 360 1648
rect 40 1544 72 1576
rect 112 1544 144 1576
rect 184 1544 216 1576
rect 256 1544 288 1576
rect 328 1544 360 1576
rect 40 1472 72 1504
rect 112 1472 144 1504
rect 184 1472 216 1504
rect 256 1472 288 1504
rect 328 1472 360 1504
rect 40 1400 72 1432
rect 112 1400 144 1432
rect 184 1400 216 1432
rect 256 1400 288 1432
rect 328 1400 360 1432
rect 40 1328 72 1360
rect 112 1328 144 1360
rect 184 1328 216 1360
rect 256 1328 288 1360
rect 328 1328 360 1360
rect 40 1256 72 1288
rect 112 1256 144 1288
rect 184 1256 216 1288
rect 256 1256 288 1288
rect 328 1256 360 1288
rect 116 31384 148 31416
rect 184 31384 216 31416
rect 252 31384 284 31416
rect 184 31316 216 31348
rect 184 27939 216 27971
rect 256 27939 288 27971
rect 112 27867 144 27899
rect 184 27867 216 27899
rect 256 27867 288 27899
rect 112 27795 144 27827
rect 184 27795 216 27827
rect 256 27795 288 27827
rect 112 27723 144 27755
rect 184 27723 216 27755
rect 256 27723 288 27755
rect 112 27651 144 27683
rect 184 27651 216 27683
rect 256 27651 288 27683
rect 112 27579 144 27611
rect 184 27579 216 27611
rect 256 27579 288 27611
rect 112 27507 144 27539
rect 184 27507 216 27539
rect 256 27507 288 27539
rect 112 27435 144 27467
rect 184 27435 216 27467
rect 256 27435 288 27467
rect 112 27363 144 27395
rect 184 27363 216 27395
rect 256 27363 288 27395
rect 112 27291 144 27323
rect 184 27291 216 27323
rect 256 27291 288 27323
rect 112 27219 144 27251
rect 184 27219 216 27251
rect 256 27219 288 27251
rect 112 27147 144 27179
rect 184 27147 216 27179
rect 256 27147 288 27179
rect 112 27075 144 27107
rect 184 27075 216 27107
rect 256 27075 288 27107
rect 112 27003 144 27035
rect 184 27003 216 27035
rect 256 27003 288 27035
rect 112 26931 144 26963
rect 184 26931 216 26963
rect 256 26931 288 26963
rect 112 26859 144 26891
rect 184 26859 216 26891
rect 256 26859 288 26891
rect 112 26787 144 26819
rect 184 26787 216 26819
rect 256 26787 288 26819
rect 112 26715 144 26747
rect 184 26715 216 26747
rect 256 26715 288 26747
rect 112 26643 144 26675
rect 184 26643 216 26675
rect 256 26643 288 26675
rect 112 26571 144 26603
rect 184 26571 216 26603
rect 256 26571 288 26603
rect 112 26499 144 26531
rect 184 26499 216 26531
rect 256 26499 288 26531
rect 112 26427 144 26459
rect 184 26427 216 26459
rect 256 26427 288 26459
rect 112 26355 144 26387
rect 184 26355 216 26387
rect 256 26355 288 26387
rect 112 26283 144 26315
rect 184 26283 216 26315
rect 256 26283 288 26315
rect 112 26211 144 26243
rect 184 26211 216 26243
rect 256 26211 288 26243
rect 112 26139 144 26171
rect 184 26139 216 26171
rect 256 26139 288 26171
rect 112 26067 144 26099
rect 184 26067 216 26099
rect 256 26067 288 26099
rect 112 25995 144 26027
rect 184 25995 216 26027
rect 256 25995 288 26027
rect 112 25923 144 25955
rect 184 25923 216 25955
rect 256 25923 288 25955
rect 112 25851 144 25883
rect 184 25851 216 25883
rect 256 25851 288 25883
rect 112 25779 144 25811
rect 184 25779 216 25811
rect 256 25779 288 25811
rect 112 25707 144 25739
rect 184 25707 216 25739
rect 256 25707 288 25739
rect 112 25635 144 25667
rect 184 25635 216 25667
rect 256 25635 288 25667
rect 112 25563 144 25595
rect 184 25563 216 25595
rect 256 25563 288 25595
rect 112 25491 144 25523
rect 184 25491 216 25523
rect 256 25491 288 25523
rect 112 25419 144 25451
rect 184 25419 216 25451
rect 256 25419 288 25451
rect 112 25347 144 25379
rect 184 25347 216 25379
rect 256 25347 288 25379
rect 112 25275 144 25307
rect 184 25275 216 25307
rect 256 25275 288 25307
rect 112 25203 144 25235
rect 184 25203 216 25235
rect 256 25203 288 25235
rect 112 25131 144 25163
rect 184 25131 216 25163
rect 256 25131 288 25163
rect 112 25059 144 25091
rect 184 25059 216 25091
rect 256 25059 288 25091
rect 112 24987 144 25019
rect 184 24987 216 25019
rect 256 24987 288 25019
rect 112 24915 144 24947
rect 184 24915 216 24947
rect 256 24915 288 24947
rect 112 24843 144 24875
rect 184 24843 216 24875
rect 256 24843 288 24875
rect 112 24771 144 24803
rect 184 24771 216 24803
rect 256 24771 288 24803
rect 112 24699 144 24731
rect 184 24699 216 24731
rect 256 24699 288 24731
rect 112 24627 144 24659
rect 184 24627 216 24659
rect 256 24627 288 24659
rect 112 24555 144 24587
rect 184 24555 216 24587
rect 256 24555 288 24587
rect 112 24483 144 24515
rect 184 24483 216 24515
rect 256 24483 288 24515
rect 112 24411 144 24443
rect 184 24411 216 24443
rect 256 24411 288 24443
rect 112 24339 144 24371
rect 184 24339 216 24371
rect 256 24339 288 24371
rect 112 24267 144 24299
rect 184 24267 216 24299
rect 256 24267 288 24299
rect 112 24195 144 24227
rect 184 24195 216 24227
rect 256 24195 288 24227
rect 112 24123 144 24155
rect 184 24123 216 24155
rect 256 24123 288 24155
rect 112 24051 144 24083
rect 184 24051 216 24083
rect 256 24051 288 24083
rect 112 23979 144 24011
rect 184 23979 216 24011
rect 256 23979 288 24011
rect 112 23907 144 23939
rect 184 23907 216 23939
rect 256 23907 288 23939
rect 112 23835 144 23867
rect 184 23835 216 23867
rect 256 23835 288 23867
rect 112 23763 144 23795
rect 184 23763 216 23795
rect 256 23763 288 23795
rect 112 23691 144 23723
rect 184 23691 216 23723
rect 256 23691 288 23723
rect 112 23619 144 23651
rect 184 23619 216 23651
rect 256 23619 288 23651
rect 112 23547 144 23579
rect 184 23547 216 23579
rect 256 23547 288 23579
rect 112 23475 144 23507
rect 184 23475 216 23507
rect 256 23475 288 23507
rect 112 23403 144 23435
rect 184 23403 216 23435
rect 256 23403 288 23435
rect 112 23331 144 23363
rect 184 23331 216 23363
rect 256 23331 288 23363
rect 112 23259 144 23291
rect 184 23259 216 23291
rect 256 23259 288 23291
rect 112 23187 144 23219
rect 184 23187 216 23219
rect 256 23187 288 23219
rect 184 22842 216 22874
rect 256 22842 288 22874
rect 112 22770 144 22802
rect 184 22770 216 22802
rect 256 22770 288 22802
rect 112 22698 144 22730
rect 184 22698 216 22730
rect 256 22698 288 22730
rect 112 22626 144 22658
rect 184 22626 216 22658
rect 256 22626 288 22658
rect 112 22554 144 22586
rect 184 22554 216 22586
rect 256 22554 288 22586
rect 112 22482 144 22514
rect 184 22482 216 22514
rect 256 22482 288 22514
rect 112 22410 144 22442
rect 184 22410 216 22442
rect 256 22410 288 22442
rect 112 22338 144 22370
rect 184 22338 216 22370
rect 256 22338 288 22370
rect 112 22266 144 22298
rect 184 22266 216 22298
rect 256 22266 288 22298
rect 112 22194 144 22226
rect 184 22194 216 22226
rect 256 22194 288 22226
rect 112 22122 144 22154
rect 184 22122 216 22154
rect 256 22122 288 22154
rect 112 22050 144 22082
rect 184 22050 216 22082
rect 256 22050 288 22082
rect 112 21978 144 22010
rect 184 21978 216 22010
rect 256 21978 288 22010
rect 112 21906 144 21938
rect 184 21906 216 21938
rect 256 21906 288 21938
rect 112 21834 144 21866
rect 184 21834 216 21866
rect 256 21834 288 21866
rect 112 21762 144 21794
rect 184 21762 216 21794
rect 256 21762 288 21794
rect 112 21690 144 21722
rect 184 21690 216 21722
rect 256 21690 288 21722
rect 112 21618 144 21650
rect 184 21618 216 21650
rect 256 21618 288 21650
rect 112 21546 144 21578
rect 184 21546 216 21578
rect 256 21546 288 21578
rect 112 21474 144 21506
rect 184 21474 216 21506
rect 256 21474 288 21506
rect 112 21402 144 21434
rect 184 21402 216 21434
rect 256 21402 288 21434
rect 112 21330 144 21362
rect 184 21330 216 21362
rect 256 21330 288 21362
rect 112 21258 144 21290
rect 184 21258 216 21290
rect 256 21258 288 21290
rect 112 21186 144 21218
rect 184 21186 216 21218
rect 256 21186 288 21218
rect 112 21114 144 21146
rect 184 21114 216 21146
rect 256 21114 288 21146
rect 112 21042 144 21074
rect 184 21042 216 21074
rect 256 21042 288 21074
rect 112 20970 144 21002
rect 184 20970 216 21002
rect 256 20970 288 21002
rect 112 20898 144 20930
rect 184 20898 216 20930
rect 256 20898 288 20930
rect 112 20826 144 20858
rect 184 20826 216 20858
rect 256 20826 288 20858
rect 112 20754 144 20786
rect 184 20754 216 20786
rect 256 20754 288 20786
rect 112 20682 144 20714
rect 184 20682 216 20714
rect 256 20682 288 20714
rect 112 20610 144 20642
rect 184 20610 216 20642
rect 256 20610 288 20642
rect 112 20538 144 20570
rect 184 20538 216 20570
rect 256 20538 288 20570
rect 112 20466 144 20498
rect 184 20466 216 20498
rect 256 20466 288 20498
rect 112 20394 144 20426
rect 184 20394 216 20426
rect 256 20394 288 20426
rect 112 20322 144 20354
rect 184 20322 216 20354
rect 256 20322 288 20354
rect 112 20250 144 20282
rect 184 20250 216 20282
rect 256 20250 288 20282
rect 112 20178 144 20210
rect 184 20178 216 20210
rect 256 20178 288 20210
rect 112 20106 144 20138
rect 184 20106 216 20138
rect 256 20106 288 20138
rect 112 20034 144 20066
rect 184 20034 216 20066
rect 256 20034 288 20066
rect 112 19962 144 19994
rect 184 19962 216 19994
rect 256 19962 288 19994
rect 112 19890 144 19922
rect 184 19890 216 19922
rect 256 19890 288 19922
rect 112 19818 144 19850
rect 184 19818 216 19850
rect 256 19818 288 19850
rect 112 19746 144 19778
rect 184 19746 216 19778
rect 256 19746 288 19778
rect 112 19674 144 19706
rect 184 19674 216 19706
rect 256 19674 288 19706
rect 112 19602 144 19634
rect 184 19602 216 19634
rect 256 19602 288 19634
rect 112 19530 144 19562
rect 184 19530 216 19562
rect 256 19530 288 19562
rect 112 19458 144 19490
rect 184 19458 216 19490
rect 256 19458 288 19490
rect 112 19386 144 19418
rect 184 19386 216 19418
rect 256 19386 288 19418
rect 112 19314 144 19346
rect 184 19314 216 19346
rect 256 19314 288 19346
rect 112 19242 144 19274
rect 184 19242 216 19274
rect 256 19242 288 19274
rect 112 19170 144 19202
rect 184 19170 216 19202
rect 256 19170 288 19202
rect 112 19098 144 19130
rect 184 19098 216 19130
rect 256 19098 288 19130
rect 112 19026 144 19058
rect 184 19026 216 19058
rect 256 19026 288 19058
rect 112 18954 144 18986
rect 184 18954 216 18986
rect 256 18954 288 18986
rect 112 18882 144 18914
rect 184 18882 216 18914
rect 256 18882 288 18914
rect 112 18810 144 18842
rect 184 18810 216 18842
rect 256 18810 288 18842
rect 112 18738 144 18770
rect 184 18738 216 18770
rect 256 18738 288 18770
rect 112 18666 144 18698
rect 184 18666 216 18698
rect 256 18666 288 18698
rect 112 18594 144 18626
rect 184 18594 216 18626
rect 256 18594 288 18626
rect 112 18522 144 18554
rect 184 18522 216 18554
rect 256 18522 288 18554
rect 112 18450 144 18482
rect 184 18450 216 18482
rect 256 18450 288 18482
rect 112 18378 144 18410
rect 184 18378 216 18410
rect 256 18378 288 18410
rect 112 18306 144 18338
rect 184 18306 216 18338
rect 256 18306 288 18338
rect 112 18234 144 18266
rect 184 18234 216 18266
rect 256 18234 288 18266
rect 112 18162 144 18194
rect 184 18162 216 18194
rect 256 18162 288 18194
rect 184 17816 216 17848
rect 256 17816 288 17848
rect 112 17744 144 17776
rect 184 17744 216 17776
rect 256 17744 288 17776
rect 112 17672 144 17704
rect 184 17672 216 17704
rect 256 17672 288 17704
rect 112 17600 144 17632
rect 184 17600 216 17632
rect 256 17600 288 17632
rect 112 17528 144 17560
rect 184 17528 216 17560
rect 256 17528 288 17560
rect 112 17456 144 17488
rect 184 17456 216 17488
rect 256 17456 288 17488
rect 112 17384 144 17416
rect 184 17384 216 17416
rect 256 17384 288 17416
rect 112 17312 144 17344
rect 184 17312 216 17344
rect 256 17312 288 17344
rect 112 17240 144 17272
rect 184 17240 216 17272
rect 256 17240 288 17272
rect 112 17168 144 17200
rect 184 17168 216 17200
rect 256 17168 288 17200
rect 112 17096 144 17128
rect 184 17096 216 17128
rect 256 17096 288 17128
rect 112 17024 144 17056
rect 184 17024 216 17056
rect 256 17024 288 17056
rect 112 16952 144 16984
rect 184 16952 216 16984
rect 256 16952 288 16984
rect 112 16880 144 16912
rect 184 16880 216 16912
rect 256 16880 288 16912
rect 112 16808 144 16840
rect 184 16808 216 16840
rect 256 16808 288 16840
rect 112 16736 144 16768
rect 184 16736 216 16768
rect 256 16736 288 16768
rect 112 16664 144 16696
rect 184 16664 216 16696
rect 256 16664 288 16696
rect 112 16592 144 16624
rect 184 16592 216 16624
rect 256 16592 288 16624
rect 112 16520 144 16552
rect 184 16520 216 16552
rect 256 16520 288 16552
rect 112 16448 144 16480
rect 184 16448 216 16480
rect 256 16448 288 16480
rect 112 16376 144 16408
rect 184 16376 216 16408
rect 256 16376 288 16408
rect 112 16304 144 16336
rect 184 16304 216 16336
rect 256 16304 288 16336
rect 112 16232 144 16264
rect 184 16232 216 16264
rect 256 16232 288 16264
rect 112 16160 144 16192
rect 184 16160 216 16192
rect 256 16160 288 16192
rect 112 16088 144 16120
rect 184 16088 216 16120
rect 256 16088 288 16120
rect 112 16016 144 16048
rect 184 16016 216 16048
rect 256 16016 288 16048
rect 112 15944 144 15976
rect 184 15944 216 15976
rect 256 15944 288 15976
rect 112 15872 144 15904
rect 184 15872 216 15904
rect 256 15872 288 15904
rect 112 15800 144 15832
rect 184 15800 216 15832
rect 256 15800 288 15832
rect 112 15728 144 15760
rect 184 15728 216 15760
rect 256 15728 288 15760
rect 112 15656 144 15688
rect 184 15656 216 15688
rect 256 15656 288 15688
rect 112 15584 144 15616
rect 184 15584 216 15616
rect 256 15584 288 15616
rect 112 15512 144 15544
rect 184 15512 216 15544
rect 256 15512 288 15544
rect 112 15440 144 15472
rect 184 15440 216 15472
rect 256 15440 288 15472
rect 112 15368 144 15400
rect 184 15368 216 15400
rect 256 15368 288 15400
rect 112 15296 144 15328
rect 184 15296 216 15328
rect 256 15296 288 15328
rect 112 15224 144 15256
rect 184 15224 216 15256
rect 256 15224 288 15256
rect 112 15152 144 15184
rect 184 15152 216 15184
rect 256 15152 288 15184
rect 112 15080 144 15112
rect 184 15080 216 15112
rect 256 15080 288 15112
rect 112 15008 144 15040
rect 184 15008 216 15040
rect 256 15008 288 15040
rect 112 14936 144 14968
rect 184 14936 216 14968
rect 256 14936 288 14968
rect 112 14864 144 14896
rect 184 14864 216 14896
rect 256 14864 288 14896
rect 112 14792 144 14824
rect 184 14792 216 14824
rect 256 14792 288 14824
rect 112 14720 144 14752
rect 184 14720 216 14752
rect 256 14720 288 14752
rect 112 14648 144 14680
rect 184 14648 216 14680
rect 256 14648 288 14680
rect 112 14576 144 14608
rect 184 14576 216 14608
rect 256 14576 288 14608
rect 112 14504 144 14536
rect 184 14504 216 14536
rect 256 14504 288 14536
rect 112 14432 144 14464
rect 184 14432 216 14464
rect 256 14432 288 14464
rect 112 14360 144 14392
rect 184 14360 216 14392
rect 256 14360 288 14392
rect 112 14288 144 14320
rect 184 14288 216 14320
rect 256 14288 288 14320
rect 112 14216 144 14248
rect 184 14216 216 14248
rect 256 14216 288 14248
rect 112 14144 144 14176
rect 184 14144 216 14176
rect 256 14144 288 14176
rect 112 14072 144 14104
rect 184 14072 216 14104
rect 256 14072 288 14104
rect 112 14000 144 14032
rect 184 14000 216 14032
rect 256 14000 288 14032
rect 112 13928 144 13960
rect 184 13928 216 13960
rect 256 13928 288 13960
rect 112 13856 144 13888
rect 184 13856 216 13888
rect 256 13856 288 13888
rect 112 13784 144 13816
rect 184 13784 216 13816
rect 256 13784 288 13816
rect 112 13712 144 13744
rect 184 13712 216 13744
rect 256 13712 288 13744
rect 112 13640 144 13672
rect 184 13640 216 13672
rect 256 13640 288 13672
rect 112 13568 144 13600
rect 184 13568 216 13600
rect 256 13568 288 13600
rect 112 13496 144 13528
rect 184 13496 216 13528
rect 256 13496 288 13528
rect 112 13424 144 13456
rect 184 13424 216 13456
rect 256 13424 288 13456
rect 112 13352 144 13384
rect 184 13352 216 13384
rect 256 13352 288 13384
rect 112 13280 144 13312
rect 184 13280 216 13312
rect 256 13280 288 13312
rect 112 13208 144 13240
rect 184 13208 216 13240
rect 256 13208 288 13240
rect 112 13136 144 13168
rect 184 13136 216 13168
rect 256 13136 288 13168
rect 112 13064 144 13096
rect 184 13064 216 13096
rect 256 13064 288 13096
rect 0 33384 112 33416
rect 144 33384 184 33416
rect 216 33384 256 33416
rect 288 33384 400 33416
rect 184 31484 216 31498
rect 184 31416 216 31452
rect 0 31384 116 31416
rect 148 31384 184 31416
rect 216 31384 252 31416
rect 284 31384 400 31416
rect 184 31348 216 31384
rect 184 31302 216 31316
rect 0 29684 112 29716
rect 144 29684 184 29716
rect 216 29684 256 29716
rect 288 29684 400 29716
rect 0 27971 400 28034
rect 0 27939 112 27971
rect 144 27939 184 27971
rect 216 27939 256 27971
rect 288 27939 400 27971
rect 0 27899 400 27939
rect 0 27867 112 27899
rect 144 27867 184 27899
rect 216 27867 256 27899
rect 288 27867 400 27899
rect 0 27827 400 27867
rect 0 27795 112 27827
rect 144 27795 184 27827
rect 216 27795 256 27827
rect 288 27795 400 27827
rect 0 27755 400 27795
rect 0 27723 112 27755
rect 144 27723 184 27755
rect 216 27723 256 27755
rect 288 27723 400 27755
rect 0 27683 400 27723
rect 0 27651 112 27683
rect 144 27651 184 27683
rect 216 27651 256 27683
rect 288 27651 400 27683
rect 0 27611 400 27651
rect 0 27579 112 27611
rect 144 27579 184 27611
rect 216 27579 256 27611
rect 288 27579 400 27611
rect 0 27539 400 27579
rect 0 27507 112 27539
rect 144 27507 184 27539
rect 216 27507 256 27539
rect 288 27507 400 27539
rect 0 27467 400 27507
rect 0 27435 112 27467
rect 144 27435 184 27467
rect 216 27435 256 27467
rect 288 27435 400 27467
rect 0 27395 400 27435
rect 0 27363 112 27395
rect 144 27363 184 27395
rect 216 27363 256 27395
rect 288 27363 400 27395
rect 0 27323 400 27363
rect 0 27291 112 27323
rect 144 27291 184 27323
rect 216 27291 256 27323
rect 288 27291 400 27323
rect 0 27251 400 27291
rect 0 27219 112 27251
rect 144 27219 184 27251
rect 216 27219 256 27251
rect 288 27219 400 27251
rect 0 27179 400 27219
rect 0 27147 112 27179
rect 144 27147 184 27179
rect 216 27147 256 27179
rect 288 27147 400 27179
rect 0 27107 400 27147
rect 0 27075 112 27107
rect 144 27075 184 27107
rect 216 27075 256 27107
rect 288 27075 400 27107
rect 0 27035 400 27075
rect 0 27003 112 27035
rect 144 27003 184 27035
rect 216 27003 256 27035
rect 288 27003 400 27035
rect 0 26963 400 27003
rect 0 26931 112 26963
rect 144 26931 184 26963
rect 216 26931 256 26963
rect 288 26931 400 26963
rect 0 26891 400 26931
rect 0 26859 112 26891
rect 144 26859 184 26891
rect 216 26859 256 26891
rect 288 26859 400 26891
rect 0 26819 400 26859
rect 0 26787 112 26819
rect 144 26787 184 26819
rect 216 26787 256 26819
rect 288 26787 400 26819
rect 0 26747 400 26787
rect 0 26715 112 26747
rect 144 26715 184 26747
rect 216 26715 256 26747
rect 288 26715 400 26747
rect 0 26675 400 26715
rect 0 26643 112 26675
rect 144 26643 184 26675
rect 216 26643 256 26675
rect 288 26643 400 26675
rect 0 26603 400 26643
rect 0 26571 112 26603
rect 144 26571 184 26603
rect 216 26571 256 26603
rect 288 26571 400 26603
rect 0 26531 400 26571
rect 0 26499 112 26531
rect 144 26499 184 26531
rect 216 26499 256 26531
rect 288 26499 400 26531
rect 0 26459 400 26499
rect 0 26427 112 26459
rect 144 26427 184 26459
rect 216 26427 256 26459
rect 288 26427 400 26459
rect 0 26387 400 26427
rect 0 26355 112 26387
rect 144 26355 184 26387
rect 216 26355 256 26387
rect 288 26355 400 26387
rect 0 26315 400 26355
rect 0 26283 112 26315
rect 144 26283 184 26315
rect 216 26283 256 26315
rect 288 26283 400 26315
rect 0 26243 400 26283
rect 0 26211 112 26243
rect 144 26211 184 26243
rect 216 26211 256 26243
rect 288 26211 400 26243
rect 0 26171 400 26211
rect 0 26139 112 26171
rect 144 26139 184 26171
rect 216 26139 256 26171
rect 288 26139 400 26171
rect 0 26099 400 26139
rect 0 26067 112 26099
rect 144 26067 184 26099
rect 216 26067 256 26099
rect 288 26067 400 26099
rect 0 26027 400 26067
rect 0 25995 112 26027
rect 144 25995 184 26027
rect 216 25995 256 26027
rect 288 25995 400 26027
rect 0 25955 400 25995
rect 0 25923 112 25955
rect 144 25923 184 25955
rect 216 25923 256 25955
rect 288 25923 400 25955
rect 0 25883 400 25923
rect 0 25851 112 25883
rect 144 25851 184 25883
rect 216 25851 256 25883
rect 288 25851 400 25883
rect 0 25811 400 25851
rect 0 25779 112 25811
rect 144 25779 184 25811
rect 216 25779 256 25811
rect 288 25779 400 25811
rect 0 25739 400 25779
rect 0 25707 112 25739
rect 144 25707 184 25739
rect 216 25707 256 25739
rect 288 25707 400 25739
rect 0 25667 400 25707
rect 0 25635 112 25667
rect 144 25635 184 25667
rect 216 25635 256 25667
rect 288 25635 400 25667
rect 0 25595 400 25635
rect 0 25563 112 25595
rect 144 25563 184 25595
rect 216 25563 256 25595
rect 288 25563 400 25595
rect 0 25523 400 25563
rect 0 25491 112 25523
rect 144 25491 184 25523
rect 216 25491 256 25523
rect 288 25491 400 25523
rect 0 25451 400 25491
rect 0 25419 112 25451
rect 144 25419 184 25451
rect 216 25419 256 25451
rect 288 25419 400 25451
rect 0 25379 400 25419
rect 0 25347 112 25379
rect 144 25347 184 25379
rect 216 25347 256 25379
rect 288 25347 400 25379
rect 0 25307 400 25347
rect 0 25275 112 25307
rect 144 25275 184 25307
rect 216 25275 256 25307
rect 288 25275 400 25307
rect 0 25235 400 25275
rect 0 25203 112 25235
rect 144 25203 184 25235
rect 216 25203 256 25235
rect 288 25203 400 25235
rect 0 25163 400 25203
rect 0 25131 112 25163
rect 144 25131 184 25163
rect 216 25131 256 25163
rect 288 25131 400 25163
rect 0 25091 400 25131
rect 0 25059 112 25091
rect 144 25059 184 25091
rect 216 25059 256 25091
rect 288 25059 400 25091
rect 0 25019 400 25059
rect 0 24987 112 25019
rect 144 24987 184 25019
rect 216 24987 256 25019
rect 288 24987 400 25019
rect 0 24947 400 24987
rect 0 24915 112 24947
rect 144 24915 184 24947
rect 216 24915 256 24947
rect 288 24915 400 24947
rect 0 24875 400 24915
rect 0 24843 112 24875
rect 144 24843 184 24875
rect 216 24843 256 24875
rect 288 24843 400 24875
rect 0 24803 400 24843
rect 0 24771 112 24803
rect 144 24771 184 24803
rect 216 24771 256 24803
rect 288 24771 400 24803
rect 0 24731 400 24771
rect 0 24699 112 24731
rect 144 24699 184 24731
rect 216 24699 256 24731
rect 288 24699 400 24731
rect 0 24659 400 24699
rect 0 24627 112 24659
rect 144 24627 184 24659
rect 216 24627 256 24659
rect 288 24627 400 24659
rect 0 24587 400 24627
rect 0 24555 112 24587
rect 144 24555 184 24587
rect 216 24555 256 24587
rect 288 24555 400 24587
rect 0 24515 400 24555
rect 0 24483 112 24515
rect 144 24483 184 24515
rect 216 24483 256 24515
rect 288 24483 400 24515
rect 0 24443 400 24483
rect 0 24411 112 24443
rect 144 24411 184 24443
rect 216 24411 256 24443
rect 288 24411 400 24443
rect 0 24371 400 24411
rect 0 24339 112 24371
rect 144 24339 184 24371
rect 216 24339 256 24371
rect 288 24339 400 24371
rect 0 24299 400 24339
rect 0 24267 112 24299
rect 144 24267 184 24299
rect 216 24267 256 24299
rect 288 24267 400 24299
rect 0 24227 400 24267
rect 0 24195 112 24227
rect 144 24195 184 24227
rect 216 24195 256 24227
rect 288 24195 400 24227
rect 0 24155 400 24195
rect 0 24123 112 24155
rect 144 24123 184 24155
rect 216 24123 256 24155
rect 288 24123 400 24155
rect 0 24083 400 24123
rect 0 24051 112 24083
rect 144 24051 184 24083
rect 216 24051 256 24083
rect 288 24051 400 24083
rect 0 24011 400 24051
rect 0 23979 112 24011
rect 144 23979 184 24011
rect 216 23979 256 24011
rect 288 23979 400 24011
rect 0 23939 400 23979
rect 0 23907 112 23939
rect 144 23907 184 23939
rect 216 23907 256 23939
rect 288 23907 400 23939
rect 0 23867 400 23907
rect 0 23835 112 23867
rect 144 23835 184 23867
rect 216 23835 256 23867
rect 288 23835 400 23867
rect 0 23795 400 23835
rect 0 23763 112 23795
rect 144 23763 184 23795
rect 216 23763 256 23795
rect 288 23763 400 23795
rect 0 23723 400 23763
rect 0 23691 112 23723
rect 144 23691 184 23723
rect 216 23691 256 23723
rect 288 23691 400 23723
rect 0 23651 400 23691
rect 0 23619 112 23651
rect 144 23619 184 23651
rect 216 23619 256 23651
rect 288 23619 400 23651
rect 0 23579 400 23619
rect 0 23547 112 23579
rect 144 23547 184 23579
rect 216 23547 256 23579
rect 288 23547 400 23579
rect 0 23507 400 23547
rect 0 23475 112 23507
rect 144 23475 184 23507
rect 216 23475 256 23507
rect 288 23475 400 23507
rect 0 23435 400 23475
rect 0 23403 112 23435
rect 144 23403 184 23435
rect 216 23403 256 23435
rect 288 23403 400 23435
rect 0 23363 400 23403
rect 0 23331 112 23363
rect 144 23331 184 23363
rect 216 23331 256 23363
rect 288 23331 400 23363
rect 0 23291 400 23331
rect 0 23259 112 23291
rect 144 23259 184 23291
rect 216 23259 256 23291
rect 288 23259 400 23291
rect 0 23219 400 23259
rect 0 23187 112 23219
rect 144 23187 184 23219
rect 216 23187 256 23219
rect 288 23187 400 23219
rect 0 23124 400 23187
rect 0 22874 400 22924
rect 0 22842 112 22874
rect 144 22842 184 22874
rect 216 22842 256 22874
rect 288 22842 400 22874
rect 0 22802 400 22842
rect 0 22770 112 22802
rect 144 22770 184 22802
rect 216 22770 256 22802
rect 288 22770 400 22802
rect 0 22730 400 22770
rect 0 22698 112 22730
rect 144 22698 184 22730
rect 216 22698 256 22730
rect 288 22698 400 22730
rect 0 22658 400 22698
rect 0 22626 112 22658
rect 144 22626 184 22658
rect 216 22626 256 22658
rect 288 22626 400 22658
rect 0 22586 400 22626
rect 0 22554 112 22586
rect 144 22554 184 22586
rect 216 22554 256 22586
rect 288 22554 400 22586
rect 0 22514 400 22554
rect 0 22482 112 22514
rect 144 22482 184 22514
rect 216 22482 256 22514
rect 288 22482 400 22514
rect 0 22442 400 22482
rect 0 22410 112 22442
rect 144 22410 184 22442
rect 216 22410 256 22442
rect 288 22410 400 22442
rect 0 22370 400 22410
rect 0 22338 112 22370
rect 144 22338 184 22370
rect 216 22338 256 22370
rect 288 22338 400 22370
rect 0 22298 400 22338
rect 0 22266 112 22298
rect 144 22266 184 22298
rect 216 22266 256 22298
rect 288 22266 400 22298
rect 0 22226 400 22266
rect 0 22194 112 22226
rect 144 22194 184 22226
rect 216 22194 256 22226
rect 288 22194 400 22226
rect 0 22154 400 22194
rect 0 22122 112 22154
rect 144 22122 184 22154
rect 216 22122 256 22154
rect 288 22122 400 22154
rect 0 22082 400 22122
rect 0 22050 112 22082
rect 144 22050 184 22082
rect 216 22050 256 22082
rect 288 22050 400 22082
rect 0 22010 400 22050
rect 0 21978 112 22010
rect 144 21978 184 22010
rect 216 21978 256 22010
rect 288 21978 400 22010
rect 0 21938 400 21978
rect 0 21906 112 21938
rect 144 21906 184 21938
rect 216 21906 256 21938
rect 288 21906 400 21938
rect 0 21866 400 21906
rect 0 21834 112 21866
rect 144 21834 184 21866
rect 216 21834 256 21866
rect 288 21834 400 21866
rect 0 21794 400 21834
rect 0 21762 112 21794
rect 144 21762 184 21794
rect 216 21762 256 21794
rect 288 21762 400 21794
rect 0 21722 400 21762
rect 0 21690 112 21722
rect 144 21690 184 21722
rect 216 21690 256 21722
rect 288 21690 400 21722
rect 0 21650 400 21690
rect 0 21618 112 21650
rect 144 21618 184 21650
rect 216 21618 256 21650
rect 288 21618 400 21650
rect 0 21578 400 21618
rect 0 21546 112 21578
rect 144 21546 184 21578
rect 216 21546 256 21578
rect 288 21546 400 21578
rect 0 21506 400 21546
rect 0 21474 112 21506
rect 144 21474 184 21506
rect 216 21474 256 21506
rect 288 21474 400 21506
rect 0 21434 400 21474
rect 0 21402 112 21434
rect 144 21402 184 21434
rect 216 21402 256 21434
rect 288 21402 400 21434
rect 0 21362 400 21402
rect 0 21330 112 21362
rect 144 21330 184 21362
rect 216 21330 256 21362
rect 288 21330 400 21362
rect 0 21290 400 21330
rect 0 21258 112 21290
rect 144 21258 184 21290
rect 216 21258 256 21290
rect 288 21258 400 21290
rect 0 21218 400 21258
rect 0 21186 112 21218
rect 144 21186 184 21218
rect 216 21186 256 21218
rect 288 21186 400 21218
rect 0 21146 400 21186
rect 0 21114 112 21146
rect 144 21114 184 21146
rect 216 21114 256 21146
rect 288 21114 400 21146
rect 0 21074 400 21114
rect 0 21042 112 21074
rect 144 21042 184 21074
rect 216 21042 256 21074
rect 288 21042 400 21074
rect 0 21002 400 21042
rect 0 20970 112 21002
rect 144 20970 184 21002
rect 216 20970 256 21002
rect 288 20970 400 21002
rect 0 20930 400 20970
rect 0 20898 112 20930
rect 144 20898 184 20930
rect 216 20898 256 20930
rect 288 20898 400 20930
rect 0 20858 400 20898
rect 0 20826 112 20858
rect 144 20826 184 20858
rect 216 20826 256 20858
rect 288 20826 400 20858
rect 0 20786 400 20826
rect 0 20754 112 20786
rect 144 20754 184 20786
rect 216 20754 256 20786
rect 288 20754 400 20786
rect 0 20714 400 20754
rect 0 20682 112 20714
rect 144 20682 184 20714
rect 216 20682 256 20714
rect 288 20682 400 20714
rect 0 20642 400 20682
rect 0 20610 112 20642
rect 144 20610 184 20642
rect 216 20610 256 20642
rect 288 20610 400 20642
rect 0 20570 400 20610
rect 0 20538 112 20570
rect 144 20538 184 20570
rect 216 20538 256 20570
rect 288 20538 400 20570
rect 0 20498 400 20538
rect 0 20466 112 20498
rect 144 20466 184 20498
rect 216 20466 256 20498
rect 288 20466 400 20498
rect 0 20426 400 20466
rect 0 20394 112 20426
rect 144 20394 184 20426
rect 216 20394 256 20426
rect 288 20394 400 20426
rect 0 20354 400 20394
rect 0 20322 112 20354
rect 144 20322 184 20354
rect 216 20322 256 20354
rect 288 20322 400 20354
rect 0 20282 400 20322
rect 0 20250 112 20282
rect 144 20250 184 20282
rect 216 20250 256 20282
rect 288 20250 400 20282
rect 0 20210 400 20250
rect 0 20178 112 20210
rect 144 20178 184 20210
rect 216 20178 256 20210
rect 288 20178 400 20210
rect 0 20138 400 20178
rect 0 20106 112 20138
rect 144 20106 184 20138
rect 216 20106 256 20138
rect 288 20106 400 20138
rect 0 20066 400 20106
rect 0 20034 112 20066
rect 144 20034 184 20066
rect 216 20034 256 20066
rect 288 20034 400 20066
rect 0 19994 400 20034
rect 0 19962 112 19994
rect 144 19962 184 19994
rect 216 19962 256 19994
rect 288 19962 400 19994
rect 0 19922 400 19962
rect 0 19890 112 19922
rect 144 19890 184 19922
rect 216 19890 256 19922
rect 288 19890 400 19922
rect 0 19850 400 19890
rect 0 19818 112 19850
rect 144 19818 184 19850
rect 216 19818 256 19850
rect 288 19818 400 19850
rect 0 19778 400 19818
rect 0 19746 112 19778
rect 144 19746 184 19778
rect 216 19746 256 19778
rect 288 19746 400 19778
rect 0 19706 400 19746
rect 0 19674 112 19706
rect 144 19674 184 19706
rect 216 19674 256 19706
rect 288 19674 400 19706
rect 0 19634 400 19674
rect 0 19602 112 19634
rect 144 19602 184 19634
rect 216 19602 256 19634
rect 288 19602 400 19634
rect 0 19562 400 19602
rect 0 19530 112 19562
rect 144 19530 184 19562
rect 216 19530 256 19562
rect 288 19530 400 19562
rect 0 19490 400 19530
rect 0 19458 112 19490
rect 144 19458 184 19490
rect 216 19458 256 19490
rect 288 19458 400 19490
rect 0 19418 400 19458
rect 0 19386 112 19418
rect 144 19386 184 19418
rect 216 19386 256 19418
rect 288 19386 400 19418
rect 0 19346 400 19386
rect 0 19314 112 19346
rect 144 19314 184 19346
rect 216 19314 256 19346
rect 288 19314 400 19346
rect 0 19274 400 19314
rect 0 19242 112 19274
rect 144 19242 184 19274
rect 216 19242 256 19274
rect 288 19242 400 19274
rect 0 19202 400 19242
rect 0 19170 112 19202
rect 144 19170 184 19202
rect 216 19170 256 19202
rect 288 19170 400 19202
rect 0 19130 400 19170
rect 0 19098 112 19130
rect 144 19098 184 19130
rect 216 19098 256 19130
rect 288 19098 400 19130
rect 0 19058 400 19098
rect 0 19026 112 19058
rect 144 19026 184 19058
rect 216 19026 256 19058
rect 288 19026 400 19058
rect 0 18986 400 19026
rect 0 18954 112 18986
rect 144 18954 184 18986
rect 216 18954 256 18986
rect 288 18954 400 18986
rect 0 18914 400 18954
rect 0 18882 112 18914
rect 144 18882 184 18914
rect 216 18882 256 18914
rect 288 18882 400 18914
rect 0 18842 400 18882
rect 0 18810 112 18842
rect 144 18810 184 18842
rect 216 18810 256 18842
rect 288 18810 400 18842
rect 0 18770 400 18810
rect 0 18738 112 18770
rect 144 18738 184 18770
rect 216 18738 256 18770
rect 288 18738 400 18770
rect 0 18698 400 18738
rect 0 18666 112 18698
rect 144 18666 184 18698
rect 216 18666 256 18698
rect 288 18666 400 18698
rect 0 18626 400 18666
rect 0 18594 112 18626
rect 144 18594 184 18626
rect 216 18594 256 18626
rect 288 18594 400 18626
rect 0 18554 400 18594
rect 0 18522 112 18554
rect 144 18522 184 18554
rect 216 18522 256 18554
rect 288 18522 400 18554
rect 0 18482 400 18522
rect 0 18450 112 18482
rect 144 18450 184 18482
rect 216 18450 256 18482
rect 288 18450 400 18482
rect 0 18410 400 18450
rect 0 18378 112 18410
rect 144 18378 184 18410
rect 216 18378 256 18410
rect 288 18378 400 18410
rect 0 18338 400 18378
rect 0 18306 112 18338
rect 144 18306 184 18338
rect 216 18306 256 18338
rect 288 18306 400 18338
rect 0 18266 400 18306
rect 0 18234 112 18266
rect 144 18234 184 18266
rect 216 18234 256 18266
rect 288 18234 400 18266
rect 0 18194 400 18234
rect 0 18162 112 18194
rect 144 18162 184 18194
rect 216 18162 256 18194
rect 288 18162 400 18194
rect 0 18112 400 18162
rect 0 17848 400 17912
rect 0 17816 112 17848
rect 144 17816 184 17848
rect 216 17816 256 17848
rect 288 17816 400 17848
rect 0 17776 400 17816
rect 0 17744 112 17776
rect 144 17744 184 17776
rect 216 17744 256 17776
rect 288 17744 400 17776
rect 0 17704 400 17744
rect 0 17672 112 17704
rect 144 17672 184 17704
rect 216 17672 256 17704
rect 288 17672 400 17704
rect 0 17632 400 17672
rect 0 17600 112 17632
rect 144 17600 184 17632
rect 216 17600 256 17632
rect 288 17600 400 17632
rect 0 17560 400 17600
rect 0 17528 112 17560
rect 144 17528 184 17560
rect 216 17528 256 17560
rect 288 17528 400 17560
rect 0 17488 400 17528
rect 0 17456 112 17488
rect 144 17456 184 17488
rect 216 17456 256 17488
rect 288 17456 400 17488
rect 0 17416 400 17456
rect 0 17384 112 17416
rect 144 17384 184 17416
rect 216 17384 256 17416
rect 288 17384 400 17416
rect 0 17344 400 17384
rect 0 17312 112 17344
rect 144 17312 184 17344
rect 216 17312 256 17344
rect 288 17312 400 17344
rect 0 17272 400 17312
rect 0 17240 112 17272
rect 144 17240 184 17272
rect 216 17240 256 17272
rect 288 17240 400 17272
rect 0 17200 400 17240
rect 0 17168 112 17200
rect 144 17168 184 17200
rect 216 17168 256 17200
rect 288 17168 400 17200
rect 0 17128 400 17168
rect 0 17096 112 17128
rect 144 17096 184 17128
rect 216 17096 256 17128
rect 288 17096 400 17128
rect 0 17056 400 17096
rect 0 17024 112 17056
rect 144 17024 184 17056
rect 216 17024 256 17056
rect 288 17024 400 17056
rect 0 16984 400 17024
rect 0 16952 112 16984
rect 144 16952 184 16984
rect 216 16952 256 16984
rect 288 16952 400 16984
rect 0 16912 400 16952
rect 0 16880 112 16912
rect 144 16880 184 16912
rect 216 16880 256 16912
rect 288 16880 400 16912
rect 0 16840 400 16880
rect 0 16808 112 16840
rect 144 16808 184 16840
rect 216 16808 256 16840
rect 288 16808 400 16840
rect 0 16768 400 16808
rect 0 16736 112 16768
rect 144 16736 184 16768
rect 216 16736 256 16768
rect 288 16736 400 16768
rect 0 16696 400 16736
rect 0 16664 112 16696
rect 144 16664 184 16696
rect 216 16664 256 16696
rect 288 16664 400 16696
rect 0 16624 400 16664
rect 0 16592 112 16624
rect 144 16592 184 16624
rect 216 16592 256 16624
rect 288 16592 400 16624
rect 0 16552 400 16592
rect 0 16520 112 16552
rect 144 16520 184 16552
rect 216 16520 256 16552
rect 288 16520 400 16552
rect 0 16480 400 16520
rect 0 16448 112 16480
rect 144 16448 184 16480
rect 216 16448 256 16480
rect 288 16448 400 16480
rect 0 16408 400 16448
rect 0 16376 112 16408
rect 144 16376 184 16408
rect 216 16376 256 16408
rect 288 16376 400 16408
rect 0 16336 400 16376
rect 0 16304 112 16336
rect 144 16304 184 16336
rect 216 16304 256 16336
rect 288 16304 400 16336
rect 0 16264 400 16304
rect 0 16232 112 16264
rect 144 16232 184 16264
rect 216 16232 256 16264
rect 288 16232 400 16264
rect 0 16192 400 16232
rect 0 16160 112 16192
rect 144 16160 184 16192
rect 216 16160 256 16192
rect 288 16160 400 16192
rect 0 16120 400 16160
rect 0 16088 112 16120
rect 144 16088 184 16120
rect 216 16088 256 16120
rect 288 16088 400 16120
rect 0 16048 400 16088
rect 0 16016 112 16048
rect 144 16016 184 16048
rect 216 16016 256 16048
rect 288 16016 400 16048
rect 0 15976 400 16016
rect 0 15944 112 15976
rect 144 15944 184 15976
rect 216 15944 256 15976
rect 288 15944 400 15976
rect 0 15904 400 15944
rect 0 15872 112 15904
rect 144 15872 184 15904
rect 216 15872 256 15904
rect 288 15872 400 15904
rect 0 15832 400 15872
rect 0 15800 112 15832
rect 144 15800 184 15832
rect 216 15800 256 15832
rect 288 15800 400 15832
rect 0 15760 400 15800
rect 0 15728 112 15760
rect 144 15728 184 15760
rect 216 15728 256 15760
rect 288 15728 400 15760
rect 0 15688 400 15728
rect 0 15656 112 15688
rect 144 15656 184 15688
rect 216 15656 256 15688
rect 288 15656 400 15688
rect 0 15616 400 15656
rect 0 15584 112 15616
rect 144 15584 184 15616
rect 216 15584 256 15616
rect 288 15584 400 15616
rect 0 15544 400 15584
rect 0 15512 112 15544
rect 144 15512 184 15544
rect 216 15512 256 15544
rect 288 15512 400 15544
rect 0 15472 400 15512
rect 0 15440 112 15472
rect 144 15440 184 15472
rect 216 15440 256 15472
rect 288 15440 400 15472
rect 0 15400 400 15440
rect 0 15368 112 15400
rect 144 15368 184 15400
rect 216 15368 256 15400
rect 288 15368 400 15400
rect 0 15328 400 15368
rect 0 15296 112 15328
rect 144 15296 184 15328
rect 216 15296 256 15328
rect 288 15296 400 15328
rect 0 15256 400 15296
rect 0 15224 112 15256
rect 144 15224 184 15256
rect 216 15224 256 15256
rect 288 15224 400 15256
rect 0 15184 400 15224
rect 0 15152 112 15184
rect 144 15152 184 15184
rect 216 15152 256 15184
rect 288 15152 400 15184
rect 0 15112 400 15152
rect 0 15080 112 15112
rect 144 15080 184 15112
rect 216 15080 256 15112
rect 288 15080 400 15112
rect 0 15040 400 15080
rect 0 15008 112 15040
rect 144 15008 184 15040
rect 216 15008 256 15040
rect 288 15008 400 15040
rect 0 14968 400 15008
rect 0 14936 112 14968
rect 144 14936 184 14968
rect 216 14936 256 14968
rect 288 14936 400 14968
rect 0 14896 400 14936
rect 0 14864 112 14896
rect 144 14864 184 14896
rect 216 14864 256 14896
rect 288 14864 400 14896
rect 0 14824 400 14864
rect 0 14792 112 14824
rect 144 14792 184 14824
rect 216 14792 256 14824
rect 288 14792 400 14824
rect 0 14752 400 14792
rect 0 14720 112 14752
rect 144 14720 184 14752
rect 216 14720 256 14752
rect 288 14720 400 14752
rect 0 14680 400 14720
rect 0 14648 112 14680
rect 144 14648 184 14680
rect 216 14648 256 14680
rect 288 14648 400 14680
rect 0 14608 400 14648
rect 0 14576 112 14608
rect 144 14576 184 14608
rect 216 14576 256 14608
rect 288 14576 400 14608
rect 0 14536 400 14576
rect 0 14504 112 14536
rect 144 14504 184 14536
rect 216 14504 256 14536
rect 288 14504 400 14536
rect 0 14464 400 14504
rect 0 14432 112 14464
rect 144 14432 184 14464
rect 216 14432 256 14464
rect 288 14432 400 14464
rect 0 14392 400 14432
rect 0 14360 112 14392
rect 144 14360 184 14392
rect 216 14360 256 14392
rect 288 14360 400 14392
rect 0 14320 400 14360
rect 0 14288 112 14320
rect 144 14288 184 14320
rect 216 14288 256 14320
rect 288 14288 400 14320
rect 0 14248 400 14288
rect 0 14216 112 14248
rect 144 14216 184 14248
rect 216 14216 256 14248
rect 288 14216 400 14248
rect 0 14176 400 14216
rect 0 14144 112 14176
rect 144 14144 184 14176
rect 216 14144 256 14176
rect 288 14144 400 14176
rect 0 14104 400 14144
rect 0 14072 112 14104
rect 144 14072 184 14104
rect 216 14072 256 14104
rect 288 14072 400 14104
rect 0 14032 400 14072
rect 0 14000 112 14032
rect 144 14000 184 14032
rect 216 14000 256 14032
rect 288 14000 400 14032
rect 0 13960 400 14000
rect 0 13928 112 13960
rect 144 13928 184 13960
rect 216 13928 256 13960
rect 288 13928 400 13960
rect 0 13888 400 13928
rect 0 13856 112 13888
rect 144 13856 184 13888
rect 216 13856 256 13888
rect 288 13856 400 13888
rect 0 13816 400 13856
rect 0 13784 112 13816
rect 144 13784 184 13816
rect 216 13784 256 13816
rect 288 13784 400 13816
rect 0 13744 400 13784
rect 0 13712 112 13744
rect 144 13712 184 13744
rect 216 13712 256 13744
rect 288 13712 400 13744
rect 0 13672 400 13712
rect 0 13640 112 13672
rect 144 13640 184 13672
rect 216 13640 256 13672
rect 288 13640 400 13672
rect 0 13600 400 13640
rect 0 13568 112 13600
rect 144 13568 184 13600
rect 216 13568 256 13600
rect 288 13568 400 13600
rect 0 13528 400 13568
rect 0 13496 112 13528
rect 144 13496 184 13528
rect 216 13496 256 13528
rect 288 13496 400 13528
rect 0 13456 400 13496
rect 0 13424 112 13456
rect 144 13424 184 13456
rect 216 13424 256 13456
rect 288 13424 400 13456
rect 0 13384 400 13424
rect 0 13352 112 13384
rect 144 13352 184 13384
rect 216 13352 256 13384
rect 288 13352 400 13384
rect 0 13312 400 13352
rect 0 13280 112 13312
rect 144 13280 184 13312
rect 216 13280 256 13312
rect 288 13280 400 13312
rect 0 13240 400 13280
rect 0 13208 112 13240
rect 144 13208 184 13240
rect 216 13208 256 13240
rect 288 13208 400 13240
rect 0 13168 400 13208
rect 0 13136 112 13168
rect 144 13136 184 13168
rect 216 13136 256 13168
rect 288 13136 400 13168
rect 0 13096 400 13136
rect 0 13064 112 13096
rect 144 13064 184 13096
rect 216 13064 256 13096
rect 288 13064 400 13096
rect 0 13000 400 13064
rect 0 12144 400 12200
rect 0 12112 40 12144
rect 72 12112 112 12144
rect 144 12112 184 12144
rect 216 12112 256 12144
rect 288 12112 328 12144
rect 360 12112 400 12144
rect 0 12072 400 12112
rect 0 12040 40 12072
rect 72 12040 112 12072
rect 144 12040 184 12072
rect 216 12040 256 12072
rect 288 12040 328 12072
rect 360 12040 400 12072
rect 0 12000 400 12040
rect 0 11968 40 12000
rect 72 11968 112 12000
rect 144 11968 184 12000
rect 216 11968 256 12000
rect 288 11968 328 12000
rect 360 11968 400 12000
rect 0 11928 400 11968
rect 0 11896 40 11928
rect 72 11896 112 11928
rect 144 11896 184 11928
rect 216 11896 256 11928
rect 288 11896 328 11928
rect 360 11896 400 11928
rect 0 11856 400 11896
rect 0 11824 40 11856
rect 72 11824 112 11856
rect 144 11824 184 11856
rect 216 11824 256 11856
rect 288 11824 328 11856
rect 360 11824 400 11856
rect 0 11784 400 11824
rect 0 11752 40 11784
rect 72 11752 112 11784
rect 144 11752 184 11784
rect 216 11752 256 11784
rect 288 11752 328 11784
rect 360 11752 400 11784
rect 0 11712 400 11752
rect 0 11680 40 11712
rect 72 11680 112 11712
rect 144 11680 184 11712
rect 216 11680 256 11712
rect 288 11680 328 11712
rect 360 11680 400 11712
rect 0 11640 400 11680
rect 0 11608 40 11640
rect 72 11608 112 11640
rect 144 11608 184 11640
rect 216 11608 256 11640
rect 288 11608 328 11640
rect 360 11608 400 11640
rect 0 11568 400 11608
rect 0 11536 40 11568
rect 72 11536 112 11568
rect 144 11536 184 11568
rect 216 11536 256 11568
rect 288 11536 328 11568
rect 360 11536 400 11568
rect 0 11496 400 11536
rect 0 11464 40 11496
rect 72 11464 112 11496
rect 144 11464 184 11496
rect 216 11464 256 11496
rect 288 11464 328 11496
rect 360 11464 400 11496
rect 0 11424 400 11464
rect 0 11392 40 11424
rect 72 11392 112 11424
rect 144 11392 184 11424
rect 216 11392 256 11424
rect 288 11392 328 11424
rect 360 11392 400 11424
rect 0 11352 400 11392
rect 0 11320 40 11352
rect 72 11320 112 11352
rect 144 11320 184 11352
rect 216 11320 256 11352
rect 288 11320 328 11352
rect 360 11320 400 11352
rect 0 11280 400 11320
rect 0 11248 40 11280
rect 72 11248 112 11280
rect 144 11248 184 11280
rect 216 11248 256 11280
rect 288 11248 328 11280
rect 360 11248 400 11280
rect 0 11208 400 11248
rect 0 11176 40 11208
rect 72 11176 112 11208
rect 144 11176 184 11208
rect 216 11176 256 11208
rect 288 11176 328 11208
rect 360 11176 400 11208
rect 0 11136 400 11176
rect 0 11104 40 11136
rect 72 11104 112 11136
rect 144 11104 184 11136
rect 216 11104 256 11136
rect 288 11104 328 11136
rect 360 11104 400 11136
rect 0 11064 400 11104
rect 0 11032 40 11064
rect 72 11032 112 11064
rect 144 11032 184 11064
rect 216 11032 256 11064
rect 288 11032 328 11064
rect 360 11032 400 11064
rect 0 10992 400 11032
rect 0 10960 40 10992
rect 72 10960 112 10992
rect 144 10960 184 10992
rect 216 10960 256 10992
rect 288 10960 328 10992
rect 360 10960 400 10992
rect 0 10920 400 10960
rect 0 10888 40 10920
rect 72 10888 112 10920
rect 144 10888 184 10920
rect 216 10888 256 10920
rect 288 10888 328 10920
rect 360 10888 400 10920
rect 0 10848 400 10888
rect 0 10816 40 10848
rect 72 10816 112 10848
rect 144 10816 184 10848
rect 216 10816 256 10848
rect 288 10816 328 10848
rect 360 10816 400 10848
rect 0 10776 400 10816
rect 0 10744 40 10776
rect 72 10744 112 10776
rect 144 10744 184 10776
rect 216 10744 256 10776
rect 288 10744 328 10776
rect 360 10744 400 10776
rect 0 10704 400 10744
rect 0 10672 40 10704
rect 72 10672 112 10704
rect 144 10672 184 10704
rect 216 10672 256 10704
rect 288 10672 328 10704
rect 360 10672 400 10704
rect 0 10632 400 10672
rect 0 10600 40 10632
rect 72 10600 112 10632
rect 144 10600 184 10632
rect 216 10600 256 10632
rect 288 10600 328 10632
rect 360 10600 400 10632
rect 0 10560 400 10600
rect 0 10528 40 10560
rect 72 10528 112 10560
rect 144 10528 184 10560
rect 216 10528 256 10560
rect 288 10528 328 10560
rect 360 10528 400 10560
rect 0 10488 400 10528
rect 0 10456 40 10488
rect 72 10456 112 10488
rect 144 10456 184 10488
rect 216 10456 256 10488
rect 288 10456 328 10488
rect 360 10456 400 10488
rect 0 10416 400 10456
rect 0 10384 40 10416
rect 72 10384 112 10416
rect 144 10384 184 10416
rect 216 10384 256 10416
rect 288 10384 328 10416
rect 360 10384 400 10416
rect 0 10344 400 10384
rect 0 10312 40 10344
rect 72 10312 112 10344
rect 144 10312 184 10344
rect 216 10312 256 10344
rect 288 10312 328 10344
rect 360 10312 400 10344
rect 0 10272 400 10312
rect 0 10240 40 10272
rect 72 10240 112 10272
rect 144 10240 184 10272
rect 216 10240 256 10272
rect 288 10240 328 10272
rect 360 10240 400 10272
rect 0 10200 400 10240
rect 0 10168 40 10200
rect 72 10168 112 10200
rect 144 10168 184 10200
rect 216 10168 256 10200
rect 288 10168 328 10200
rect 360 10168 400 10200
rect 0 10128 400 10168
rect 0 10096 40 10128
rect 72 10096 112 10128
rect 144 10096 184 10128
rect 216 10096 256 10128
rect 288 10096 328 10128
rect 360 10096 400 10128
rect 0 10056 400 10096
rect 0 10024 40 10056
rect 72 10024 112 10056
rect 144 10024 184 10056
rect 216 10024 256 10056
rect 288 10024 328 10056
rect 360 10024 400 10056
rect 0 9984 400 10024
rect 0 9952 40 9984
rect 72 9952 112 9984
rect 144 9952 184 9984
rect 216 9952 256 9984
rect 288 9952 328 9984
rect 360 9952 400 9984
rect 0 9912 400 9952
rect 0 9880 40 9912
rect 72 9880 112 9912
rect 144 9880 184 9912
rect 216 9880 256 9912
rect 288 9880 328 9912
rect 360 9880 400 9912
rect 0 9840 400 9880
rect 0 9808 40 9840
rect 72 9808 112 9840
rect 144 9808 184 9840
rect 216 9808 256 9840
rect 288 9808 328 9840
rect 360 9808 400 9840
rect 0 9768 400 9808
rect 0 9736 40 9768
rect 72 9736 112 9768
rect 144 9736 184 9768
rect 216 9736 256 9768
rect 288 9736 328 9768
rect 360 9736 400 9768
rect 0 9696 400 9736
rect 0 9664 40 9696
rect 72 9664 112 9696
rect 144 9664 184 9696
rect 216 9664 256 9696
rect 288 9664 328 9696
rect 360 9664 400 9696
rect 0 9624 400 9664
rect 0 9592 40 9624
rect 72 9592 112 9624
rect 144 9592 184 9624
rect 216 9592 256 9624
rect 288 9592 328 9624
rect 360 9592 400 9624
rect 0 9552 400 9592
rect 0 9520 40 9552
rect 72 9520 112 9552
rect 144 9520 184 9552
rect 216 9520 256 9552
rect 288 9520 328 9552
rect 360 9520 400 9552
rect 0 9480 400 9520
rect 0 9448 40 9480
rect 72 9448 112 9480
rect 144 9448 184 9480
rect 216 9448 256 9480
rect 288 9448 328 9480
rect 360 9448 400 9480
rect 0 9408 400 9448
rect 0 9376 40 9408
rect 72 9376 112 9408
rect 144 9376 184 9408
rect 216 9376 256 9408
rect 288 9376 328 9408
rect 360 9376 400 9408
rect 0 9336 400 9376
rect 0 9304 40 9336
rect 72 9304 112 9336
rect 144 9304 184 9336
rect 216 9304 256 9336
rect 288 9304 328 9336
rect 360 9304 400 9336
rect 0 9264 400 9304
rect 0 9232 40 9264
rect 72 9232 112 9264
rect 144 9232 184 9264
rect 216 9232 256 9264
rect 288 9232 328 9264
rect 360 9232 400 9264
rect 0 9192 400 9232
rect 0 9160 40 9192
rect 72 9160 112 9192
rect 144 9160 184 9192
rect 216 9160 256 9192
rect 288 9160 328 9192
rect 360 9160 400 9192
rect 0 9120 400 9160
rect 0 9088 40 9120
rect 72 9088 112 9120
rect 144 9088 184 9120
rect 216 9088 256 9120
rect 288 9088 328 9120
rect 360 9088 400 9120
rect 0 9048 400 9088
rect 0 9016 40 9048
rect 72 9016 112 9048
rect 144 9016 184 9048
rect 216 9016 256 9048
rect 288 9016 328 9048
rect 360 9016 400 9048
rect 0 8976 400 9016
rect 0 8944 40 8976
rect 72 8944 112 8976
rect 144 8944 184 8976
rect 216 8944 256 8976
rect 288 8944 328 8976
rect 360 8944 400 8976
rect 0 8904 400 8944
rect 0 8872 40 8904
rect 72 8872 112 8904
rect 144 8872 184 8904
rect 216 8872 256 8904
rect 288 8872 328 8904
rect 360 8872 400 8904
rect 0 8832 400 8872
rect 0 8800 40 8832
rect 72 8800 112 8832
rect 144 8800 184 8832
rect 216 8800 256 8832
rect 288 8800 328 8832
rect 360 8800 400 8832
rect 0 8760 400 8800
rect 0 8728 40 8760
rect 72 8728 112 8760
rect 144 8728 184 8760
rect 216 8728 256 8760
rect 288 8728 328 8760
rect 360 8728 400 8760
rect 0 8688 400 8728
rect 0 8656 40 8688
rect 72 8656 112 8688
rect 144 8656 184 8688
rect 216 8656 256 8688
rect 288 8656 328 8688
rect 360 8656 400 8688
rect 0 8616 400 8656
rect 0 8584 40 8616
rect 72 8584 112 8616
rect 144 8584 184 8616
rect 216 8584 256 8616
rect 288 8584 328 8616
rect 360 8584 400 8616
rect 0 8544 400 8584
rect 0 8512 40 8544
rect 72 8512 112 8544
rect 144 8512 184 8544
rect 216 8512 256 8544
rect 288 8512 328 8544
rect 360 8512 400 8544
rect 0 8472 400 8512
rect 0 8440 40 8472
rect 72 8440 112 8472
rect 144 8440 184 8472
rect 216 8440 256 8472
rect 288 8440 328 8472
rect 360 8440 400 8472
rect 0 8400 400 8440
rect 0 8368 40 8400
rect 72 8368 112 8400
rect 144 8368 184 8400
rect 216 8368 256 8400
rect 288 8368 328 8400
rect 360 8368 400 8400
rect 0 8328 400 8368
rect 0 8296 40 8328
rect 72 8296 112 8328
rect 144 8296 184 8328
rect 216 8296 256 8328
rect 288 8296 328 8328
rect 360 8296 400 8328
rect 0 8256 400 8296
rect 0 8224 40 8256
rect 72 8224 112 8256
rect 144 8224 184 8256
rect 216 8224 256 8256
rect 288 8224 328 8256
rect 360 8224 400 8256
rect 0 8184 400 8224
rect 0 8152 40 8184
rect 72 8152 112 8184
rect 144 8152 184 8184
rect 216 8152 256 8184
rect 288 8152 328 8184
rect 360 8152 400 8184
rect 0 8112 400 8152
rect 0 8080 40 8112
rect 72 8080 112 8112
rect 144 8080 184 8112
rect 216 8080 256 8112
rect 288 8080 328 8112
rect 360 8080 400 8112
rect 0 8040 400 8080
rect 0 8008 40 8040
rect 72 8008 112 8040
rect 144 8008 184 8040
rect 216 8008 256 8040
rect 288 8008 328 8040
rect 360 8008 400 8040
rect 0 7968 400 8008
rect 0 7936 40 7968
rect 72 7936 112 7968
rect 144 7936 184 7968
rect 216 7936 256 7968
rect 288 7936 328 7968
rect 360 7936 400 7968
rect 0 7896 400 7936
rect 0 7864 40 7896
rect 72 7864 112 7896
rect 144 7864 184 7896
rect 216 7864 256 7896
rect 288 7864 328 7896
rect 360 7864 400 7896
rect 0 7824 400 7864
rect 0 7792 40 7824
rect 72 7792 112 7824
rect 144 7792 184 7824
rect 216 7792 256 7824
rect 288 7792 328 7824
rect 360 7792 400 7824
rect 0 7752 400 7792
rect 0 7720 40 7752
rect 72 7720 112 7752
rect 144 7720 184 7752
rect 216 7720 256 7752
rect 288 7720 328 7752
rect 360 7720 400 7752
rect 0 7680 400 7720
rect 0 7648 40 7680
rect 72 7648 112 7680
rect 144 7648 184 7680
rect 216 7648 256 7680
rect 288 7648 328 7680
rect 360 7648 400 7680
rect 0 7608 400 7648
rect 0 7576 40 7608
rect 72 7576 112 7608
rect 144 7576 184 7608
rect 216 7576 256 7608
rect 288 7576 328 7608
rect 360 7576 400 7608
rect 0 7536 400 7576
rect 0 7504 40 7536
rect 72 7504 112 7536
rect 144 7504 184 7536
rect 216 7504 256 7536
rect 288 7504 328 7536
rect 360 7504 400 7536
rect 0 7464 400 7504
rect 0 7432 40 7464
rect 72 7432 112 7464
rect 144 7432 184 7464
rect 216 7432 256 7464
rect 288 7432 328 7464
rect 360 7432 400 7464
rect 0 7392 400 7432
rect 0 7360 40 7392
rect 72 7360 112 7392
rect 144 7360 184 7392
rect 216 7360 256 7392
rect 288 7360 328 7392
rect 360 7360 400 7392
rect 0 7320 400 7360
rect 0 7288 40 7320
rect 72 7288 112 7320
rect 144 7288 184 7320
rect 216 7288 256 7320
rect 288 7288 328 7320
rect 360 7288 400 7320
rect 0 7248 400 7288
rect 0 7216 40 7248
rect 72 7216 112 7248
rect 144 7216 184 7248
rect 216 7216 256 7248
rect 288 7216 328 7248
rect 360 7216 400 7248
rect 0 7176 400 7216
rect 0 7144 40 7176
rect 72 7144 112 7176
rect 144 7144 184 7176
rect 216 7144 256 7176
rect 288 7144 328 7176
rect 360 7144 400 7176
rect 0 7104 400 7144
rect 0 7072 40 7104
rect 72 7072 112 7104
rect 144 7072 184 7104
rect 216 7072 256 7104
rect 288 7072 328 7104
rect 360 7072 400 7104
rect 0 7032 400 7072
rect 0 7000 40 7032
rect 72 7000 112 7032
rect 144 7000 184 7032
rect 216 7000 256 7032
rect 288 7000 328 7032
rect 360 7000 400 7032
rect 0 6960 400 7000
rect 0 6928 40 6960
rect 72 6928 112 6960
rect 144 6928 184 6960
rect 216 6928 256 6960
rect 288 6928 328 6960
rect 360 6928 400 6960
rect 0 6888 400 6928
rect 0 6856 40 6888
rect 72 6856 112 6888
rect 144 6856 184 6888
rect 216 6856 256 6888
rect 288 6856 328 6888
rect 360 6856 400 6888
rect 0 6800 400 6856
rect 0 6544 400 6600
rect 0 6512 40 6544
rect 72 6512 112 6544
rect 144 6512 184 6544
rect 216 6512 256 6544
rect 288 6512 328 6544
rect 360 6512 400 6544
rect 0 6472 400 6512
rect 0 6440 40 6472
rect 72 6440 112 6472
rect 144 6440 184 6472
rect 216 6440 256 6472
rect 288 6440 328 6472
rect 360 6440 400 6472
rect 0 6400 400 6440
rect 0 6368 40 6400
rect 72 6368 112 6400
rect 144 6368 184 6400
rect 216 6368 256 6400
rect 288 6368 328 6400
rect 360 6368 400 6400
rect 0 6328 400 6368
rect 0 6296 40 6328
rect 72 6296 112 6328
rect 144 6296 184 6328
rect 216 6296 256 6328
rect 288 6296 328 6328
rect 360 6296 400 6328
rect 0 6256 400 6296
rect 0 6224 40 6256
rect 72 6224 112 6256
rect 144 6224 184 6256
rect 216 6224 256 6256
rect 288 6224 328 6256
rect 360 6224 400 6256
rect 0 6184 400 6224
rect 0 6152 40 6184
rect 72 6152 112 6184
rect 144 6152 184 6184
rect 216 6152 256 6184
rect 288 6152 328 6184
rect 360 6152 400 6184
rect 0 6112 400 6152
rect 0 6080 40 6112
rect 72 6080 112 6112
rect 144 6080 184 6112
rect 216 6080 256 6112
rect 288 6080 328 6112
rect 360 6080 400 6112
rect 0 6040 400 6080
rect 0 6008 40 6040
rect 72 6008 112 6040
rect 144 6008 184 6040
rect 216 6008 256 6040
rect 288 6008 328 6040
rect 360 6008 400 6040
rect 0 5968 400 6008
rect 0 5936 40 5968
rect 72 5936 112 5968
rect 144 5936 184 5968
rect 216 5936 256 5968
rect 288 5936 328 5968
rect 360 5936 400 5968
rect 0 5896 400 5936
rect 0 5864 40 5896
rect 72 5864 112 5896
rect 144 5864 184 5896
rect 216 5864 256 5896
rect 288 5864 328 5896
rect 360 5864 400 5896
rect 0 5824 400 5864
rect 0 5792 40 5824
rect 72 5792 112 5824
rect 144 5792 184 5824
rect 216 5792 256 5824
rect 288 5792 328 5824
rect 360 5792 400 5824
rect 0 5752 400 5792
rect 0 5720 40 5752
rect 72 5720 112 5752
rect 144 5720 184 5752
rect 216 5720 256 5752
rect 288 5720 328 5752
rect 360 5720 400 5752
rect 0 5680 400 5720
rect 0 5648 40 5680
rect 72 5648 112 5680
rect 144 5648 184 5680
rect 216 5648 256 5680
rect 288 5648 328 5680
rect 360 5648 400 5680
rect 0 5608 400 5648
rect 0 5576 40 5608
rect 72 5576 112 5608
rect 144 5576 184 5608
rect 216 5576 256 5608
rect 288 5576 328 5608
rect 360 5576 400 5608
rect 0 5536 400 5576
rect 0 5504 40 5536
rect 72 5504 112 5536
rect 144 5504 184 5536
rect 216 5504 256 5536
rect 288 5504 328 5536
rect 360 5504 400 5536
rect 0 5464 400 5504
rect 0 5432 40 5464
rect 72 5432 112 5464
rect 144 5432 184 5464
rect 216 5432 256 5464
rect 288 5432 328 5464
rect 360 5432 400 5464
rect 0 5392 400 5432
rect 0 5360 40 5392
rect 72 5360 112 5392
rect 144 5360 184 5392
rect 216 5360 256 5392
rect 288 5360 328 5392
rect 360 5360 400 5392
rect 0 5320 400 5360
rect 0 5288 40 5320
rect 72 5288 112 5320
rect 144 5288 184 5320
rect 216 5288 256 5320
rect 288 5288 328 5320
rect 360 5288 400 5320
rect 0 5248 400 5288
rect 0 5216 40 5248
rect 72 5216 112 5248
rect 144 5216 184 5248
rect 216 5216 256 5248
rect 288 5216 328 5248
rect 360 5216 400 5248
rect 0 5176 400 5216
rect 0 5144 40 5176
rect 72 5144 112 5176
rect 144 5144 184 5176
rect 216 5144 256 5176
rect 288 5144 328 5176
rect 360 5144 400 5176
rect 0 5104 400 5144
rect 0 5072 40 5104
rect 72 5072 112 5104
rect 144 5072 184 5104
rect 216 5072 256 5104
rect 288 5072 328 5104
rect 360 5072 400 5104
rect 0 5032 400 5072
rect 0 5000 40 5032
rect 72 5000 112 5032
rect 144 5000 184 5032
rect 216 5000 256 5032
rect 288 5000 328 5032
rect 360 5000 400 5032
rect 0 4960 400 5000
rect 0 4928 40 4960
rect 72 4928 112 4960
rect 144 4928 184 4960
rect 216 4928 256 4960
rect 288 4928 328 4960
rect 360 4928 400 4960
rect 0 4888 400 4928
rect 0 4856 40 4888
rect 72 4856 112 4888
rect 144 4856 184 4888
rect 216 4856 256 4888
rect 288 4856 328 4888
rect 360 4856 400 4888
rect 0 4816 400 4856
rect 0 4784 40 4816
rect 72 4784 112 4816
rect 144 4784 184 4816
rect 216 4784 256 4816
rect 288 4784 328 4816
rect 360 4784 400 4816
rect 0 4744 400 4784
rect 0 4712 40 4744
rect 72 4712 112 4744
rect 144 4712 184 4744
rect 216 4712 256 4744
rect 288 4712 328 4744
rect 360 4712 400 4744
rect 0 4672 400 4712
rect 0 4640 40 4672
rect 72 4640 112 4672
rect 144 4640 184 4672
rect 216 4640 256 4672
rect 288 4640 328 4672
rect 360 4640 400 4672
rect 0 4600 400 4640
rect 0 4568 40 4600
rect 72 4568 112 4600
rect 144 4568 184 4600
rect 216 4568 256 4600
rect 288 4568 328 4600
rect 360 4568 400 4600
rect 0 4528 400 4568
rect 0 4496 40 4528
rect 72 4496 112 4528
rect 144 4496 184 4528
rect 216 4496 256 4528
rect 288 4496 328 4528
rect 360 4496 400 4528
rect 0 4456 400 4496
rect 0 4424 40 4456
rect 72 4424 112 4456
rect 144 4424 184 4456
rect 216 4424 256 4456
rect 288 4424 328 4456
rect 360 4424 400 4456
rect 0 4384 400 4424
rect 0 4352 40 4384
rect 72 4352 112 4384
rect 144 4352 184 4384
rect 216 4352 256 4384
rect 288 4352 328 4384
rect 360 4352 400 4384
rect 0 4312 400 4352
rect 0 4280 40 4312
rect 72 4280 112 4312
rect 144 4280 184 4312
rect 216 4280 256 4312
rect 288 4280 328 4312
rect 360 4280 400 4312
rect 0 4240 400 4280
rect 0 4208 40 4240
rect 72 4208 112 4240
rect 144 4208 184 4240
rect 216 4208 256 4240
rect 288 4208 328 4240
rect 360 4208 400 4240
rect 0 4168 400 4208
rect 0 4136 40 4168
rect 72 4136 112 4168
rect 144 4136 184 4168
rect 216 4136 256 4168
rect 288 4136 328 4168
rect 360 4136 400 4168
rect 0 4096 400 4136
rect 0 4064 40 4096
rect 72 4064 112 4096
rect 144 4064 184 4096
rect 216 4064 256 4096
rect 288 4064 328 4096
rect 360 4064 400 4096
rect 0 4024 400 4064
rect 0 3992 40 4024
rect 72 3992 112 4024
rect 144 3992 184 4024
rect 216 3992 256 4024
rect 288 3992 328 4024
rect 360 3992 400 4024
rect 0 3952 400 3992
rect 0 3920 40 3952
rect 72 3920 112 3952
rect 144 3920 184 3952
rect 216 3920 256 3952
rect 288 3920 328 3952
rect 360 3920 400 3952
rect 0 3880 400 3920
rect 0 3848 40 3880
rect 72 3848 112 3880
rect 144 3848 184 3880
rect 216 3848 256 3880
rect 288 3848 328 3880
rect 360 3848 400 3880
rect 0 3808 400 3848
rect 0 3776 40 3808
rect 72 3776 112 3808
rect 144 3776 184 3808
rect 216 3776 256 3808
rect 288 3776 328 3808
rect 360 3776 400 3808
rect 0 3736 400 3776
rect 0 3704 40 3736
rect 72 3704 112 3736
rect 144 3704 184 3736
rect 216 3704 256 3736
rect 288 3704 328 3736
rect 360 3704 400 3736
rect 0 3664 400 3704
rect 0 3632 40 3664
rect 72 3632 112 3664
rect 144 3632 184 3664
rect 216 3632 256 3664
rect 288 3632 328 3664
rect 360 3632 400 3664
rect 0 3592 400 3632
rect 0 3560 40 3592
rect 72 3560 112 3592
rect 144 3560 184 3592
rect 216 3560 256 3592
rect 288 3560 328 3592
rect 360 3560 400 3592
rect 0 3520 400 3560
rect 0 3488 40 3520
rect 72 3488 112 3520
rect 144 3488 184 3520
rect 216 3488 256 3520
rect 288 3488 328 3520
rect 360 3488 400 3520
rect 0 3448 400 3488
rect 0 3416 40 3448
rect 72 3416 112 3448
rect 144 3416 184 3448
rect 216 3416 256 3448
rect 288 3416 328 3448
rect 360 3416 400 3448
rect 0 3376 400 3416
rect 0 3344 40 3376
rect 72 3344 112 3376
rect 144 3344 184 3376
rect 216 3344 256 3376
rect 288 3344 328 3376
rect 360 3344 400 3376
rect 0 3304 400 3344
rect 0 3272 40 3304
rect 72 3272 112 3304
rect 144 3272 184 3304
rect 216 3272 256 3304
rect 288 3272 328 3304
rect 360 3272 400 3304
rect 0 3232 400 3272
rect 0 3200 40 3232
rect 72 3200 112 3232
rect 144 3200 184 3232
rect 216 3200 256 3232
rect 288 3200 328 3232
rect 360 3200 400 3232
rect 0 3160 400 3200
rect 0 3128 40 3160
rect 72 3128 112 3160
rect 144 3128 184 3160
rect 216 3128 256 3160
rect 288 3128 328 3160
rect 360 3128 400 3160
rect 0 3088 400 3128
rect 0 3056 40 3088
rect 72 3056 112 3088
rect 144 3056 184 3088
rect 216 3056 256 3088
rect 288 3056 328 3088
rect 360 3056 400 3088
rect 0 3016 400 3056
rect 0 2984 40 3016
rect 72 2984 112 3016
rect 144 2984 184 3016
rect 216 2984 256 3016
rect 288 2984 328 3016
rect 360 2984 400 3016
rect 0 2944 400 2984
rect 0 2912 40 2944
rect 72 2912 112 2944
rect 144 2912 184 2944
rect 216 2912 256 2944
rect 288 2912 328 2944
rect 360 2912 400 2944
rect 0 2872 400 2912
rect 0 2840 40 2872
rect 72 2840 112 2872
rect 144 2840 184 2872
rect 216 2840 256 2872
rect 288 2840 328 2872
rect 360 2840 400 2872
rect 0 2800 400 2840
rect 0 2768 40 2800
rect 72 2768 112 2800
rect 144 2768 184 2800
rect 216 2768 256 2800
rect 288 2768 328 2800
rect 360 2768 400 2800
rect 0 2728 400 2768
rect 0 2696 40 2728
rect 72 2696 112 2728
rect 144 2696 184 2728
rect 216 2696 256 2728
rect 288 2696 328 2728
rect 360 2696 400 2728
rect 0 2656 400 2696
rect 0 2624 40 2656
rect 72 2624 112 2656
rect 144 2624 184 2656
rect 216 2624 256 2656
rect 288 2624 328 2656
rect 360 2624 400 2656
rect 0 2584 400 2624
rect 0 2552 40 2584
rect 72 2552 112 2584
rect 144 2552 184 2584
rect 216 2552 256 2584
rect 288 2552 328 2584
rect 360 2552 400 2584
rect 0 2512 400 2552
rect 0 2480 40 2512
rect 72 2480 112 2512
rect 144 2480 184 2512
rect 216 2480 256 2512
rect 288 2480 328 2512
rect 360 2480 400 2512
rect 0 2440 400 2480
rect 0 2408 40 2440
rect 72 2408 112 2440
rect 144 2408 184 2440
rect 216 2408 256 2440
rect 288 2408 328 2440
rect 360 2408 400 2440
rect 0 2368 400 2408
rect 0 2336 40 2368
rect 72 2336 112 2368
rect 144 2336 184 2368
rect 216 2336 256 2368
rect 288 2336 328 2368
rect 360 2336 400 2368
rect 0 2296 400 2336
rect 0 2264 40 2296
rect 72 2264 112 2296
rect 144 2264 184 2296
rect 216 2264 256 2296
rect 288 2264 328 2296
rect 360 2264 400 2296
rect 0 2224 400 2264
rect 0 2192 40 2224
rect 72 2192 112 2224
rect 144 2192 184 2224
rect 216 2192 256 2224
rect 288 2192 328 2224
rect 360 2192 400 2224
rect 0 2152 400 2192
rect 0 2120 40 2152
rect 72 2120 112 2152
rect 144 2120 184 2152
rect 216 2120 256 2152
rect 288 2120 328 2152
rect 360 2120 400 2152
rect 0 2080 400 2120
rect 0 2048 40 2080
rect 72 2048 112 2080
rect 144 2048 184 2080
rect 216 2048 256 2080
rect 288 2048 328 2080
rect 360 2048 400 2080
rect 0 2008 400 2048
rect 0 1976 40 2008
rect 72 1976 112 2008
rect 144 1976 184 2008
rect 216 1976 256 2008
rect 288 1976 328 2008
rect 360 1976 400 2008
rect 0 1936 400 1976
rect 0 1904 40 1936
rect 72 1904 112 1936
rect 144 1904 184 1936
rect 216 1904 256 1936
rect 288 1904 328 1936
rect 360 1904 400 1936
rect 0 1864 400 1904
rect 0 1832 40 1864
rect 72 1832 112 1864
rect 144 1832 184 1864
rect 216 1832 256 1864
rect 288 1832 328 1864
rect 360 1832 400 1864
rect 0 1792 400 1832
rect 0 1760 40 1792
rect 72 1760 112 1792
rect 144 1760 184 1792
rect 216 1760 256 1792
rect 288 1760 328 1792
rect 360 1760 400 1792
rect 0 1720 400 1760
rect 0 1688 40 1720
rect 72 1688 112 1720
rect 144 1688 184 1720
rect 216 1688 256 1720
rect 288 1688 328 1720
rect 360 1688 400 1720
rect 0 1648 400 1688
rect 0 1616 40 1648
rect 72 1616 112 1648
rect 144 1616 184 1648
rect 216 1616 256 1648
rect 288 1616 328 1648
rect 360 1616 400 1648
rect 0 1576 400 1616
rect 0 1544 40 1576
rect 72 1544 112 1576
rect 144 1544 184 1576
rect 216 1544 256 1576
rect 288 1544 328 1576
rect 360 1544 400 1576
rect 0 1504 400 1544
rect 0 1472 40 1504
rect 72 1472 112 1504
rect 144 1472 184 1504
rect 216 1472 256 1504
rect 288 1472 328 1504
rect 360 1472 400 1504
rect 0 1432 400 1472
rect 0 1400 40 1432
rect 72 1400 112 1432
rect 144 1400 184 1432
rect 216 1400 256 1432
rect 288 1400 328 1432
rect 360 1400 400 1432
rect 0 1360 400 1400
rect 0 1328 40 1360
rect 72 1328 112 1360
rect 144 1328 184 1360
rect 216 1328 256 1360
rect 288 1328 328 1360
rect 360 1328 400 1360
rect 0 1288 400 1328
rect 0 1256 40 1288
rect 72 1256 112 1288
rect 144 1256 184 1288
rect 216 1256 256 1288
rect 288 1256 328 1288
rect 360 1256 400 1288
rect 0 1200 400 1256
<< metal3 >>
rect 0 32000 400 35600
rect 0 28000 400 31600
rect 0 25200 400 26800
rect 0 18700 400 23800
rect 0 13200 400 18300
rect 0 6900 400 12000
rect 0 1400 400 6500
<< metal4 >>
rect 0 32440 400 35600
rect 0 28000 400 31160
rect 0 25200 400 26800
rect 0 18700 400 23800
rect 0 13200 400 18300
rect 0 6900 400 12000
rect 0 1400 400 6500
<< metal5 >>
rect 0 32000 400 35600
rect 0 28000 400 31600
rect 0 25200 400 26800
rect 0 18700 400 23800
rect 0 13200 400 18300
rect 0 6900 400 12000
rect 0 1400 400 6500
<< metal6 >>
rect 0 32000 400 35600
rect 0 28000 400 31600
rect 0 25200 400 26800
rect 0 18700 400 23800
rect 0 13200 400 18300
rect 0 6900 400 12000
rect 0 1400 400 6500
<< metal7 >>
rect 0 25500 400 26500
rect 0 19000 400 23500
rect 0 13500 400 18000
rect 0 7200 400 11700
rect 0 1700 400 6200
<< labels >>
rlabel metal3 s 0 32000 400 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 400 31600 4 vss
port 1 nsew
rlabel metal3 s 0 13200 400 18300 4 iovdd
port 4 nsew
rlabel metal3 s 0 18700 400 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 6900 400 12000 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 400 6500 4 iovss
port 3 nsew
rlabel metal3 s 0 25200 400 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 400 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 400 35600 4 vss
port 1 nsew
rlabel metal4 s 0 13200 400 18300 4 iovdd
port 4 nsew
rlabel metal4 s 0 18700 400 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 6900 400 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 400 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 25200 400 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 400 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 400 35600 4 vss
port 1 nsew
rlabel metal5 s 0 13200 400 18300 4 iovdd
port 4 nsew
rlabel metal5 s 0 18700 400 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 6900 400 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 400 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 25200 400 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 400 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 400 35600 4 vss
port 1 nsew
rlabel metal6 s 0 13200 400 18300 4 iovdd
port 4 nsew
rlabel metal6 s 0 18700 400 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 6900 400 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 400 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 25200 400 26800 4 iovss
port 3 nsew
rlabel metal7 s 0 19000 400 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 13500 400 18000 4 iovdd
port 4 nsew
rlabel metal7 s 0 25500 400 26500 4 iovss
port 3 nsew
rlabel metal7 s 0 7200 400 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 1700 400 6200 4 iovss
port 3 nsew
flabel comment s 201 31406 201 31406 0 FreeSans 400 0 0 0 sub!
flabel comment s 144 17716 144 17716 0 FreeSans 400 0 0 0 sub!
flabel comment s 144 22746 144 22746 0 FreeSans 400 0 0 0 sub!
flabel comment s 144 27899 144 27899 0 FreeSans 400 0 0 0 sub!
flabel metal1 s 184 31394 228 31409 0 FreeSans 400 0 0 0 vss
port 1 nsew
flabel metal1 s 119 6535 243 6580 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 142 12096 256 12161 0 FreeSans 400 0 0 0 iovdd
port 4 nsew
flabel metal1 s 179 17776 271 17842 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 179 22786 271 22852 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 179 27929 271 27995 0 FreeSans 400 0 0 0 iovss
port 3 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 400 36000
string GDS_END 63578248
string GDS_FILE sg13g2_io.gds
string GDS_START 63482824
<< end >>
