magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2127 -6054 3768 4524
<< metal1 >>
rect 0 2161 1644 2400
rect 0 2121 9 2161
rect 49 2121 1644 2161
rect 0 2112 1644 2121
rect 270 2067 312 2076
rect 270 2027 271 2067
rect 311 2027 312 2067
rect 270 2018 312 2027
rect 750 2067 792 2076
rect 750 2027 751 2067
rect 791 2027 792 2067
rect 750 2018 792 2027
rect 880 1258 922 1267
rect 880 1218 881 1258
rect 921 1218 922 1258
rect 880 1209 922 1218
rect 1230 1258 1272 1267
rect 1230 1218 1231 1258
rect 1271 1218 1272 1258
rect 1230 1209 1272 1218
rect 400 1158 442 1167
rect 400 1118 401 1158
rect 441 1118 442 1158
rect 400 1109 442 1118
rect 1332 1158 1374 1167
rect 1332 1118 1333 1158
rect 1373 1118 1374 1158
rect 1332 1109 1374 1118
rect 478 373 520 382
rect 478 333 479 373
rect 519 333 520 373
rect 478 324 520 333
rect 958 373 1000 382
rect 958 333 959 373
rect 999 333 1000 373
rect 958 324 1000 333
rect 0 49 1644 288
rect 0 9 1595 49
rect 1635 9 1644 49
rect 0 0 1644 9
rect 8 -188 942 -179
rect 8 -228 9 -188
rect 49 -221 942 -188
rect 49 -228 50 -221
rect 8 -237 50 -228
rect 1594 -2159 1636 -2150
rect 1594 -2199 1595 -2159
rect 1635 -2199 1636 -2159
rect 1594 -2208 1636 -2199
rect 0 -3921 1644 -3879
<< via1 >>
rect 9 2121 49 2161
rect 271 2027 311 2067
rect 751 2027 791 2067
rect 881 1218 921 1258
rect 1231 1218 1271 1258
rect 401 1118 441 1158
rect 1333 1118 1373 1158
rect 479 333 519 373
rect 959 333 999 373
rect 1595 9 1635 49
rect 9 -228 49 -188
rect 1595 -2199 1635 -2159
<< metal2 >>
rect 9 2161 49 2170
rect 9 -188 49 2121
rect 271 2076 329 2400
rect 271 2067 791 2076
rect 311 2027 751 2067
rect 271 2018 791 2027
rect 881 1267 939 2400
rect 881 1258 1271 1267
rect 921 1218 1231 1258
rect 881 1209 1271 1218
rect 401 1158 1373 1167
rect 441 1118 1333 1158
rect 401 1109 1373 1118
rect 9 -237 49 -228
rect 475 373 519 382
rect 475 333 479 373
rect 475 324 519 333
rect 959 373 1217 382
rect 999 333 1217 373
rect 959 324 1217 333
rect 475 -2047 515 324
rect 1177 -2047 1217 324
rect 1595 49 1635 58
rect 1595 -2159 1635 9
rect 1595 -2208 1635 -2199
rect 876 -3696 916 -2408
rect 1578 -3696 1618 -2408
use sg13g2_io_inv_x1  sg13g2_io_inv_x1_0
timestamp 1755542813
transform 1 0 1200 0 1 0
box -124 -5 364 2524
use sg13g2_io_nand2_x1  sg13g2_io_nand2_x1_0
timestamp 1755542813
transform 1 0 720 0 1 0
box -124 -5 604 2524
use sg13g2_io_nor2_x1  sg13g2_io_nor2_x1_0
timestamp 1755542813
transform 1 0 240 0 1 0
box -124 -5 604 2524
use sg13g2_io_tie  sg13g2_io_tie_0
timestamp 1755542813
transform 1 0 0 0 1 0
box -124 -5 364 2524
use sg13g2_LevelUp  sg13g2_LevelUp_0
timestamp 1755542813
transform 1 0 240 0 1 -3900
box -124 -154 826 3854
use sg13g2_LevelUp  sg13g2_LevelUp_1
timestamp 1755542813
transform 1 0 942 0 1 -3900
box -124 -154 826 3854
<< labels >>
rlabel metal1 s 0 -3921 1644 -3879 4 iovdd
port 3 nsew
rlabel metal1 s 0 2112 1644 2400 4 vdd
port 1 nsew
rlabel metal1 s 0 0 1644 288 4 vss
port 2 nsew
flabel metal2 s 881 1209 939 2400 0 FreeSans 800 0 0 0 en
port 5 nsew
rlabel metal2 s 876 -3696 916 -2408 4 ngate
port 6 nsew
rlabel metal2 s 271 2018 329 2400 4 core
port 4 nsew
flabel metal2 s 1578 -3696 1618 -2408 0 FreeSans 800 0 0 0 pgate
port 7 nsew
<< properties >>
string device primitive
string GDS_END 22710006
string GDS_FILE sg13g2_io.gds
string GDS_START 22706728
<< end >>
