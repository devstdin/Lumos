magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752511086
<< nwell >>
rect -868 1612 -816 2172
rect 5 1728 49 1768
rect -407 1344 -121 1378
rect 550 1367 1370 2172
rect -707 134 -621 182
rect -407 -8 288 1344
<< metal1 >>
rect -868 2000 659 2129
rect -868 1688 -685 2000
rect -441 1888 -369 1940
rect -194 1908 279 1940
rect -653 1814 -473 1866
rect -421 1792 -389 1888
rect -194 1866 -157 1908
rect 207 1888 279 1908
rect -337 1864 -157 1866
rect -337 1816 -327 1864
rect -167 1816 -157 1864
rect -337 1814 -157 1816
rect -5 1863 175 1866
rect -5 1817 5 1863
rect 165 1817 175 1863
rect -5 1814 175 1817
rect 227 1792 259 1888
rect 311 1814 491 1866
rect -441 1772 -369 1792
rect -441 1768 59 1772
rect -441 1740 5 1768
rect -5 1728 5 1740
rect 49 1728 59 1768
rect 207 1740 279 1792
rect -5 1724 59 1728
rect 508 1688 659 2000
rect -868 1572 659 1688
rect -868 1274 334 1384
rect -868 49 -812 1274
rect -718 1235 -611 1238
rect -718 1189 -706 1235
rect -621 1189 -611 1235
rect -718 1186 -611 1189
rect 26 1235 133 1238
rect 26 1189 38 1235
rect 123 1189 133 1235
rect 26 1186 133 1189
rect -768 238 -662 1132
rect -612 1122 -556 1132
rect -612 248 -606 1122
rect -562 248 -556 1122
rect -612 238 -556 248
rect -24 238 82 1132
rect 132 1122 188 1132
rect 132 248 138 1122
rect 182 248 188 1122
rect 132 238 188 248
rect -718 182 -611 184
rect -718 134 -707 182
rect -621 134 -611 182
rect -718 132 -611 134
rect 26 182 133 184
rect 26 134 37 182
rect 123 134 133 182
rect 26 132 133 134
rect 283 49 334 1274
rect 552 1309 659 1572
rect 552 1195 1298 1309
rect 552 99 697 1195
rect 924 1091 996 1143
rect 727 287 898 1059
rect 944 255 976 1091
rect 1022 1049 1078 1059
rect 1022 297 1032 1049
rect 1072 297 1078 1049
rect 1022 287 1078 297
rect 924 245 996 255
rect 924 196 934 245
rect 986 196 996 245
rect 924 187 996 196
rect 1200 100 1298 1195
rect -868 -8 334 49
rect -868 -920 -811 -62
rect -417 -72 -118 -62
rect -417 -116 -407 -72
rect -367 -116 -170 -72
rect -128 -116 -118 -72
rect -417 -126 -118 -116
rect -718 -153 -611 -150
rect -718 -199 -704 -153
rect -621 -199 -611 -153
rect 26 -153 133 -150
rect -718 -202 -611 -199
rect -777 -778 -662 -256
rect -612 -265 -556 -256
rect -612 -768 -606 -265
rect -562 -768 -556 -265
rect -461 -276 -54 -186
rect 26 -199 40 -153
rect 123 -199 133 -153
rect 26 -202 133 -199
rect -329 -331 -257 -328
rect -329 -377 -319 -331
rect -267 -377 -257 -331
rect -329 -380 -257 -377
rect -175 -334 -119 -324
rect -612 -778 -556 -768
rect -462 -784 -355 -412
rect -309 -816 -277 -380
rect -175 -412 -170 -334
rect -231 -452 -170 -412
rect -125 -452 -119 -334
rect -231 -462 -119 -452
rect -231 -784 -175 -462
rect -33 -778 82 -256
rect 132 -265 188 -256
rect 132 -768 138 -265
rect 182 -768 188 -265
rect 283 -276 1297 -186
rect 924 -317 996 -312
rect 415 -331 487 -328
rect 415 -377 425 -331
rect 477 -377 487 -331
rect 415 -380 487 -377
rect 569 -334 625 -324
rect 132 -778 188 -768
rect 282 -784 389 -412
rect 435 -816 467 -380
rect 569 -412 574 -334
rect 513 -452 574 -412
rect 619 -452 625 -334
rect 924 -360 934 -317
rect 986 -360 996 -317
rect 924 -380 996 -360
rect 513 -462 625 -452
rect 513 -784 569 -462
rect 726 -784 898 -412
rect 944 -816 976 -380
rect 1022 -422 1078 -412
rect 1022 -774 1032 -422
rect 1072 -774 1078 -422
rect 1022 -784 1078 -774
rect -718 -835 -611 -832
rect -718 -881 -706 -835
rect -621 -881 -611 -835
rect -329 -868 -257 -816
rect 26 -835 133 -832
rect -718 -884 -611 -881
rect 26 -881 38 -835
rect 123 -881 133 -835
rect 415 -868 487 -816
rect 924 -868 996 -816
rect 26 -884 133 -881
rect 1200 -920 1297 -276
rect -868 -1043 1297 -920
<< via1 >>
rect -327 1816 -167 1864
rect 5 1817 165 1863
rect 5 1728 49 1768
rect -706 1189 -621 1235
rect 38 1189 123 1235
rect -606 248 -562 1122
rect 138 248 182 1122
rect -707 134 -621 182
rect 37 134 123 182
rect 1032 297 1072 1049
rect 934 196 986 245
rect -407 -116 -367 -72
rect -170 -116 -128 -72
rect -704 -199 -621 -153
rect -606 -768 -562 -265
rect 40 -199 123 -153
rect -319 -377 -267 -331
rect -170 -452 -125 -334
rect 138 -768 182 -265
rect 425 -377 477 -331
rect 574 -452 619 -334
rect 934 -360 986 -317
rect 1032 -774 1072 -422
rect -706 -881 -621 -835
rect 38 -881 123 -835
<< metal2 >>
rect -337 1864 -157 1866
rect -337 1816 -327 1864
rect -167 1816 -157 1864
rect -337 1814 -157 1816
rect -215 1670 -157 1814
rect -298 1614 -157 1670
rect -5 1863 175 1866
rect -5 1817 5 1863
rect 165 1817 175 1863
rect -5 1814 175 1817
rect -5 1768 59 1814
rect -5 1728 5 1768
rect 49 1728 59 1768
rect -5 1670 59 1728
rect -5 1614 479 1670
rect -820 1235 -611 1238
rect -820 1189 -706 1235
rect -621 1189 -611 1235
rect -820 1186 -611 1189
rect -820 184 -760 1186
rect -612 1122 -556 1132
rect -612 248 -606 1122
rect -562 289 -556 1122
rect -562 248 -510 289
rect -612 238 -510 248
rect -820 182 -611 184
rect -820 134 -707 182
rect -621 134 -611 182
rect -820 132 -611 134
rect -820 54 -760 132
rect -868 -132 -760 54
rect -820 -150 -760 -132
rect -556 -62 -510 238
rect -556 -72 -356 -62
rect -556 -116 -407 -72
rect -367 -116 -356 -72
rect -556 -126 -356 -116
rect -820 -153 -611 -150
rect -820 -199 -704 -153
rect -621 -199 -611 -153
rect -820 -202 -611 -199
rect -820 -832 -760 -202
rect -556 -256 -510 -126
rect -612 -265 -510 -256
rect -612 -768 -606 -265
rect -562 -328 -510 -265
rect -298 -220 -248 1614
rect -76 1235 133 1238
rect -76 1189 38 1235
rect 123 1189 133 1235
rect -76 1186 133 1189
rect -76 184 -16 1186
rect 132 1122 188 1132
rect 132 248 138 1122
rect 182 289 188 1122
rect 182 248 234 289
rect 132 238 234 248
rect -76 182 133 184
rect -76 134 37 182
rect 123 134 133 182
rect -76 132 133 134
rect -76 -62 -16 132
rect -180 -72 -16 -62
rect -180 -116 -170 -72
rect -128 -116 -16 -72
rect -180 -126 -16 -116
rect -76 -150 -16 -126
rect -76 -153 133 -150
rect -76 -199 40 -153
rect 123 -199 133 -153
rect -76 -202 133 -199
rect -298 -276 -119 -220
rect -562 -331 -257 -328
rect -562 -377 -319 -331
rect -267 -377 -257 -331
rect -562 -380 -257 -377
rect -175 -334 -119 -276
rect -562 -768 -556 -380
rect -175 -452 -170 -334
rect -125 -452 -119 -334
rect -175 -462 -119 -452
rect -612 -778 -556 -768
rect -76 -832 -16 -202
rect 188 -256 234 238
rect 132 -265 234 -256
rect 132 -768 138 -265
rect 182 -328 234 -265
rect 423 7 479 1614
rect 1022 1049 1135 1059
rect 1022 297 1032 1049
rect 1072 297 1135 1049
rect 1022 287 1135 297
rect 789 196 934 245
rect 986 196 996 245
rect 789 187 996 196
rect 789 7 850 187
rect 423 -65 850 7
rect 423 -220 479 -65
rect 423 -276 625 -220
rect 182 -331 487 -328
rect 182 -377 425 -331
rect 477 -377 487 -331
rect 182 -380 487 -377
rect 569 -334 625 -276
rect 182 -768 188 -380
rect 569 -452 574 -334
rect 619 -452 625 -334
rect 789 -312 850 -65
rect 1077 29 1135 287
rect 1077 -111 1301 29
rect 789 -317 996 -312
rect 789 -360 934 -317
rect 986 -360 996 -317
rect 789 -370 996 -360
rect 1077 -412 1135 -111
rect 569 -462 625 -452
rect 1022 -422 1135 -412
rect 132 -778 188 -768
rect 1022 -774 1032 -422
rect 1072 -774 1135 -422
rect 1022 -784 1135 -774
rect -820 -835 -611 -832
rect -820 -881 -706 -835
rect -621 -881 -611 -835
rect -820 -884 -611 -881
rect -76 -835 133 -832
rect -76 -881 38 -835
rect 123 -881 133 -835
rect -76 -884 133 -881
use hvnmos_S23XCS  hvnmos_S23XCS_0
timestamp 1752442741
transform 1 0 960 0 1 -598
box -286 -378 286 378
use hvnmos_SAXWCS  hvnmos_SAXWCS_0
timestamp 1752440150
transform 1 0 -293 0 1 -598
box -118 -378 118 378
use hvnmos_SAXWCS  hvnmos_SAXWCS_1
timestamp 1752440150
transform 1 0 451 0 1 -598
box -118 -378 118 378
use hvpmos_G6BEXS  hvpmos_G6BEXS_0
timestamp 1752441215
transform 1 0 -405 0 1 1840
box -416 -332 1064 332
use hvpmos_Q23XCS  hvpmos_Q23XCS_0
timestamp 1752442741
transform 1 0 960 0 1 673
box -410 -702 410 702
use lvnmos_5Y4P6Y  lvnmos_5Y4P6Y_0
timestamp 1752439852
transform 1 0 -637 0 1 -517
box -183 -459 183 459
use lvnmos_5Y4P6Y  lvnmos_5Y4P6Y_1
timestamp 1752439852
transform 1 0 107 0 1 -517
box -183 -459 183 459
use lvpmos_5A4K6Y  lvpmos_5A4K6Y_0
timestamp 1752439852
transform 1 0 -637 0 1 685
box -231 -693 231 693
use lvpmos_5A4K6Y  lvpmos_5A4K6Y_1
timestamp 1752439852
transform 1 0 107 0 1 685
box -231 -693 231 693
<< labels >>
flabel metal1 -868 1066 -821 1384 0 FreeSans 400 0 0 0 VDDL
port 1 nsew
flabel metal1 -868 -1043 -821 -725 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal2 -868 -132 -821 54 0 FreeSans 400 0 0 0 IN
port 3 nsew
flabel metal2 1253 -111 1301 29 0 FreeSans 400 0 0 0 OUT
port 4 nsew
flabel metal1 -868 1572 -751 2129 0 FreeSans 400 0 0 0 VDDH
port 0 nsew
<< end >>
