magic
tech ihp-sg13g2
magscale 1 2
timestamp 1748517704
<< error_p >>
rect -1586 14768 -1576 14778
rect 1576 14768 1586 14778
rect -1596 14758 -1586 14768
rect 1586 14758 1596 14768
rect -1596 14736 -1586 14746
rect 1586 14736 1596 14746
rect -1586 14726 -1576 14736
rect 1576 14726 1586 14736
rect -1654 14694 -1644 14704
rect -1632 14694 -1622 14704
rect 1622 14694 1632 14704
rect 1644 14694 1654 14704
rect -1664 14684 -1654 14694
rect -1622 14684 -1612 14694
rect 1612 14684 1622 14694
rect 1654 14684 1664 14694
rect -1664 13722 -1654 13732
rect -1622 13722 -1612 13732
rect 1612 13722 1622 13732
rect 1654 13722 1664 13732
rect -1654 13712 -1644 13722
rect -1632 13712 -1622 13722
rect 1622 13712 1632 13722
rect 1644 13712 1654 13722
rect -1586 13680 -1576 13690
rect 1576 13680 1586 13690
rect -1596 13670 -1586 13680
rect 1586 13670 1596 13680
rect -1596 13648 -1586 13658
rect 1586 13648 1596 13658
rect -1586 13638 -1576 13648
rect 1576 13638 1586 13648
rect -1586 13584 -1576 13594
rect 1576 13584 1586 13594
rect -1596 13574 -1586 13584
rect 1586 13574 1596 13584
rect -1596 13552 -1586 13562
rect 1586 13552 1596 13562
rect -1586 13542 -1576 13552
rect 1576 13542 1586 13552
rect -1654 13510 -1644 13520
rect -1632 13510 -1622 13520
rect 1622 13510 1632 13520
rect 1644 13510 1654 13520
rect -1664 13500 -1654 13510
rect -1622 13500 -1612 13510
rect 1612 13500 1622 13510
rect 1654 13500 1664 13510
rect -1664 12538 -1654 12548
rect -1622 12538 -1612 12548
rect 1612 12538 1622 12548
rect 1654 12538 1664 12548
rect -1654 12528 -1644 12538
rect -1632 12528 -1622 12538
rect 1622 12528 1632 12538
rect 1644 12528 1654 12538
rect -1586 12496 -1576 12506
rect 1576 12496 1586 12506
rect -1596 12486 -1586 12496
rect 1586 12486 1596 12496
rect -1596 12464 -1586 12474
rect 1586 12464 1596 12474
rect -1586 12454 -1576 12464
rect 1576 12454 1586 12464
rect -1586 12400 -1576 12410
rect 1576 12400 1586 12410
rect -1596 12390 -1586 12400
rect 1586 12390 1596 12400
rect -1596 12368 -1586 12378
rect 1586 12368 1596 12378
rect -1586 12358 -1576 12368
rect 1576 12358 1586 12368
rect -1654 12326 -1644 12336
rect -1632 12326 -1622 12336
rect 1622 12326 1632 12336
rect 1644 12326 1654 12336
rect -1664 12316 -1654 12326
rect -1622 12316 -1612 12326
rect 1612 12316 1622 12326
rect 1654 12316 1664 12326
rect -1664 11354 -1654 11364
rect -1622 11354 -1612 11364
rect 1612 11354 1622 11364
rect 1654 11354 1664 11364
rect -1654 11344 -1644 11354
rect -1632 11344 -1622 11354
rect 1622 11344 1632 11354
rect 1644 11344 1654 11354
rect -1586 11312 -1576 11322
rect 1576 11312 1586 11322
rect -1596 11302 -1586 11312
rect 1586 11302 1596 11312
rect -1596 11280 -1586 11290
rect 1586 11280 1596 11290
rect -1586 11270 -1576 11280
rect 1576 11270 1586 11280
rect -1586 11216 -1576 11226
rect 1576 11216 1586 11226
rect -1596 11206 -1586 11216
rect 1586 11206 1596 11216
rect -1596 11184 -1586 11194
rect 1586 11184 1596 11194
rect -1586 11174 -1576 11184
rect 1576 11174 1586 11184
rect -1654 11142 -1644 11152
rect -1632 11142 -1622 11152
rect 1622 11142 1632 11152
rect 1644 11142 1654 11152
rect -1664 11132 -1654 11142
rect -1622 11132 -1612 11142
rect 1612 11132 1622 11142
rect 1654 11132 1664 11142
rect -1664 10170 -1654 10180
rect -1622 10170 -1612 10180
rect 1612 10170 1622 10180
rect 1654 10170 1664 10180
rect -1654 10160 -1644 10170
rect -1632 10160 -1622 10170
rect 1622 10160 1632 10170
rect 1644 10160 1654 10170
rect -1586 10128 -1576 10138
rect 1576 10128 1586 10138
rect -1596 10118 -1586 10128
rect 1586 10118 1596 10128
rect -1596 10096 -1586 10106
rect 1586 10096 1596 10106
rect -1586 10086 -1576 10096
rect 1576 10086 1586 10096
rect -1586 10032 -1576 10042
rect 1576 10032 1586 10042
rect -1596 10022 -1586 10032
rect 1586 10022 1596 10032
rect -1596 10000 -1586 10010
rect 1586 10000 1596 10010
rect -1586 9990 -1576 10000
rect 1576 9990 1586 10000
rect -1654 9958 -1644 9968
rect -1632 9958 -1622 9968
rect 1622 9958 1632 9968
rect 1644 9958 1654 9968
rect -1664 9948 -1654 9958
rect -1622 9948 -1612 9958
rect 1612 9948 1622 9958
rect 1654 9948 1664 9958
rect -1664 8986 -1654 8996
rect -1622 8986 -1612 8996
rect 1612 8986 1622 8996
rect 1654 8986 1664 8996
rect -1654 8976 -1644 8986
rect -1632 8976 -1622 8986
rect 1622 8976 1632 8986
rect 1644 8976 1654 8986
rect -1586 8944 -1576 8954
rect 1576 8944 1586 8954
rect -1596 8934 -1586 8944
rect 1586 8934 1596 8944
rect -1596 8912 -1586 8922
rect 1586 8912 1596 8922
rect -1586 8902 -1576 8912
rect 1576 8902 1586 8912
rect -1586 8848 -1576 8858
rect 1576 8848 1586 8858
rect -1596 8838 -1586 8848
rect 1586 8838 1596 8848
rect -1596 8816 -1586 8826
rect 1586 8816 1596 8826
rect -1586 8806 -1576 8816
rect 1576 8806 1586 8816
rect -1654 8774 -1644 8784
rect -1632 8774 -1622 8784
rect 1622 8774 1632 8784
rect 1644 8774 1654 8784
rect -1664 8764 -1654 8774
rect -1622 8764 -1612 8774
rect 1612 8764 1622 8774
rect 1654 8764 1664 8774
rect -1664 7802 -1654 7812
rect -1622 7802 -1612 7812
rect 1612 7802 1622 7812
rect 1654 7802 1664 7812
rect -1654 7792 -1644 7802
rect -1632 7792 -1622 7802
rect 1622 7792 1632 7802
rect 1644 7792 1654 7802
rect -1586 7760 -1576 7770
rect 1576 7760 1586 7770
rect -1596 7750 -1586 7760
rect 1586 7750 1596 7760
rect -1596 7728 -1586 7738
rect 1586 7728 1596 7738
rect -1586 7718 -1576 7728
rect 1576 7718 1586 7728
rect -1586 7664 -1576 7674
rect 1576 7664 1586 7674
rect -1596 7654 -1586 7664
rect 1586 7654 1596 7664
rect -1596 7632 -1586 7642
rect 1586 7632 1596 7642
rect -1586 7622 -1576 7632
rect 1576 7622 1586 7632
rect -1654 7590 -1644 7600
rect -1632 7590 -1622 7600
rect 1622 7590 1632 7600
rect 1644 7590 1654 7600
rect -1664 7580 -1654 7590
rect -1622 7580 -1612 7590
rect 1612 7580 1622 7590
rect 1654 7580 1664 7590
rect -1664 6618 -1654 6628
rect -1622 6618 -1612 6628
rect 1612 6618 1622 6628
rect 1654 6618 1664 6628
rect -1654 6608 -1644 6618
rect -1632 6608 -1622 6618
rect 1622 6608 1632 6618
rect 1644 6608 1654 6618
rect -1586 6576 -1576 6586
rect 1576 6576 1586 6586
rect -1596 6566 -1586 6576
rect 1586 6566 1596 6576
rect -1596 6544 -1586 6554
rect 1586 6544 1596 6554
rect -1586 6534 -1576 6544
rect 1576 6534 1586 6544
rect -1586 6480 -1576 6490
rect 1576 6480 1586 6490
rect -1596 6470 -1586 6480
rect 1586 6470 1596 6480
rect -1596 6448 -1586 6458
rect 1586 6448 1596 6458
rect -1586 6438 -1576 6448
rect 1576 6438 1586 6448
rect -1654 6406 -1644 6416
rect -1632 6406 -1622 6416
rect 1622 6406 1632 6416
rect 1644 6406 1654 6416
rect -1664 6396 -1654 6406
rect -1622 6396 -1612 6406
rect 1612 6396 1622 6406
rect 1654 6396 1664 6406
rect -1664 5434 -1654 5444
rect -1622 5434 -1612 5444
rect 1612 5434 1622 5444
rect 1654 5434 1664 5444
rect -1654 5424 -1644 5434
rect -1632 5424 -1622 5434
rect 1622 5424 1632 5434
rect 1644 5424 1654 5434
rect -1586 5392 -1576 5402
rect 1576 5392 1586 5402
rect -1596 5382 -1586 5392
rect 1586 5382 1596 5392
rect -1596 5360 -1586 5370
rect 1586 5360 1596 5370
rect -1586 5350 -1576 5360
rect 1576 5350 1586 5360
rect -1586 5296 -1576 5306
rect 1576 5296 1586 5306
rect -1596 5286 -1586 5296
rect 1586 5286 1596 5296
rect -1596 5264 -1586 5274
rect 1586 5264 1596 5274
rect -1586 5254 -1576 5264
rect 1576 5254 1586 5264
rect -1654 5222 -1644 5232
rect -1632 5222 -1622 5232
rect 1622 5222 1632 5232
rect 1644 5222 1654 5232
rect -1664 5212 -1654 5222
rect -1622 5212 -1612 5222
rect 1612 5212 1622 5222
rect 1654 5212 1664 5222
rect -1664 4250 -1654 4260
rect -1622 4250 -1612 4260
rect 1612 4250 1622 4260
rect 1654 4250 1664 4260
rect -1654 4240 -1644 4250
rect -1632 4240 -1622 4250
rect 1622 4240 1632 4250
rect 1644 4240 1654 4250
rect -1586 4208 -1576 4218
rect 1576 4208 1586 4218
rect -1596 4198 -1586 4208
rect 1586 4198 1596 4208
rect -1596 4176 -1586 4186
rect 1586 4176 1596 4186
rect -1586 4166 -1576 4176
rect 1576 4166 1586 4176
rect -1586 4112 -1576 4122
rect 1576 4112 1586 4122
rect -1596 4102 -1586 4112
rect 1586 4102 1596 4112
rect -1596 4080 -1586 4090
rect 1586 4080 1596 4090
rect -1586 4070 -1576 4080
rect 1576 4070 1586 4080
rect -1654 4038 -1644 4048
rect -1632 4038 -1622 4048
rect 1622 4038 1632 4048
rect 1644 4038 1654 4048
rect -1664 4028 -1654 4038
rect -1622 4028 -1612 4038
rect 1612 4028 1622 4038
rect 1654 4028 1664 4038
rect -1664 3066 -1654 3076
rect -1622 3066 -1612 3076
rect 1612 3066 1622 3076
rect 1654 3066 1664 3076
rect -1654 3056 -1644 3066
rect -1632 3056 -1622 3066
rect 1622 3056 1632 3066
rect 1644 3056 1654 3066
rect -1586 3024 -1576 3034
rect 1576 3024 1586 3034
rect -1596 3014 -1586 3024
rect 1586 3014 1596 3024
rect -1596 2992 -1586 3002
rect 1586 2992 1596 3002
rect -1586 2982 -1576 2992
rect 1576 2982 1586 2992
rect -1586 2928 -1576 2938
rect 1576 2928 1586 2938
rect -1596 2918 -1586 2928
rect 1586 2918 1596 2928
rect -1596 2896 -1586 2906
rect 1586 2896 1596 2906
rect -1586 2886 -1576 2896
rect 1576 2886 1586 2896
rect -1654 2854 -1644 2864
rect -1632 2854 -1622 2864
rect 1622 2854 1632 2864
rect 1644 2854 1654 2864
rect -1664 2844 -1654 2854
rect -1622 2844 -1612 2854
rect 1612 2844 1622 2854
rect 1654 2844 1664 2854
rect -1664 1882 -1654 1892
rect -1622 1882 -1612 1892
rect 1612 1882 1622 1892
rect 1654 1882 1664 1892
rect -1654 1872 -1644 1882
rect -1632 1872 -1622 1882
rect 1622 1872 1632 1882
rect 1644 1872 1654 1882
rect -1586 1840 -1576 1850
rect 1576 1840 1586 1850
rect -1596 1830 -1586 1840
rect 1586 1830 1596 1840
rect -1596 1808 -1586 1818
rect 1586 1808 1596 1818
rect -1586 1798 -1576 1808
rect 1576 1798 1586 1808
rect -1586 1744 -1576 1754
rect 1576 1744 1586 1754
rect -1596 1734 -1586 1744
rect 1586 1734 1596 1744
rect -1596 1712 -1586 1722
rect 1586 1712 1596 1722
rect -1586 1702 -1576 1712
rect 1576 1702 1586 1712
rect -1654 1670 -1644 1680
rect -1632 1670 -1622 1680
rect 1622 1670 1632 1680
rect 1644 1670 1654 1680
rect -1664 1660 -1654 1670
rect -1622 1660 -1612 1670
rect 1612 1660 1622 1670
rect 1654 1660 1664 1670
rect -1664 698 -1654 708
rect -1622 698 -1612 708
rect 1612 698 1622 708
rect 1654 698 1664 708
rect -1654 688 -1644 698
rect -1632 688 -1622 698
rect 1622 688 1632 698
rect 1644 688 1654 698
rect -1586 656 -1576 666
rect 1576 656 1586 666
rect -1596 646 -1586 656
rect 1586 646 1596 656
rect -1596 624 -1586 634
rect 1586 624 1596 634
rect -1586 614 -1576 624
rect 1576 614 1586 624
rect -1586 560 -1576 570
rect 1576 560 1586 570
rect -1596 550 -1586 560
rect 1586 550 1596 560
rect -1596 528 -1586 538
rect 1586 528 1596 538
rect -1586 518 -1576 528
rect 1576 518 1586 528
rect -1654 486 -1644 496
rect -1632 486 -1622 496
rect 1622 486 1632 496
rect 1644 486 1654 496
rect -1664 476 -1654 486
rect -1622 476 -1612 486
rect 1612 476 1622 486
rect 1654 476 1664 486
rect -1664 -486 -1654 -476
rect -1622 -486 -1612 -476
rect 1612 -486 1622 -476
rect 1654 -486 1664 -476
rect -1654 -496 -1644 -486
rect -1632 -496 -1622 -486
rect 1622 -496 1632 -486
rect 1644 -496 1654 -486
rect -1586 -528 -1576 -518
rect 1576 -528 1586 -518
rect -1596 -538 -1586 -528
rect 1586 -538 1596 -528
rect -1596 -560 -1586 -550
rect 1586 -560 1596 -550
rect -1586 -570 -1576 -560
rect 1576 -570 1586 -560
<< hvnmos >>
rect -1600 13708 1600 14708
rect -1600 12524 1600 13524
rect -1600 11340 1600 12340
rect -1600 10156 1600 11156
rect -1600 8972 1600 9972
rect -1600 7788 1600 8788
rect -1600 6604 1600 7604
rect -1600 5420 1600 6420
rect -1600 4236 1600 5236
rect -1600 3052 1600 4052
rect -1600 1868 1600 2868
rect -1600 684 1600 1684
rect -1600 -500 1600 500
<< hvndiff >>
rect -1668 14694 -1600 14708
rect -1668 13722 -1654 14694
rect -1622 13722 -1600 14694
rect -1668 13708 -1600 13722
rect 1600 14694 1668 14708
rect 1600 13722 1622 14694
rect 1654 13722 1668 14694
rect 1600 13708 1668 13722
rect -1668 13510 -1600 13524
rect -1668 12538 -1654 13510
rect -1622 12538 -1600 13510
rect -1668 12524 -1600 12538
rect 1600 13510 1668 13524
rect 1600 12538 1622 13510
rect 1654 12538 1668 13510
rect 1600 12524 1668 12538
rect -1668 12326 -1600 12340
rect -1668 11354 -1654 12326
rect -1622 11354 -1600 12326
rect -1668 11340 -1600 11354
rect 1600 12326 1668 12340
rect 1600 11354 1622 12326
rect 1654 11354 1668 12326
rect 1600 11340 1668 11354
rect -1668 11142 -1600 11156
rect -1668 10170 -1654 11142
rect -1622 10170 -1600 11142
rect -1668 10156 -1600 10170
rect 1600 11142 1668 11156
rect 1600 10170 1622 11142
rect 1654 10170 1668 11142
rect 1600 10156 1668 10170
rect -1668 9958 -1600 9972
rect -1668 8986 -1654 9958
rect -1622 8986 -1600 9958
rect -1668 8972 -1600 8986
rect 1600 9958 1668 9972
rect 1600 8986 1622 9958
rect 1654 8986 1668 9958
rect 1600 8972 1668 8986
rect -1668 8774 -1600 8788
rect -1668 7802 -1654 8774
rect -1622 7802 -1600 8774
rect -1668 7788 -1600 7802
rect 1600 8774 1668 8788
rect 1600 7802 1622 8774
rect 1654 7802 1668 8774
rect 1600 7788 1668 7802
rect -1668 7590 -1600 7604
rect -1668 6618 -1654 7590
rect -1622 6618 -1600 7590
rect -1668 6604 -1600 6618
rect 1600 7590 1668 7604
rect 1600 6618 1622 7590
rect 1654 6618 1668 7590
rect 1600 6604 1668 6618
rect -1668 6406 -1600 6420
rect -1668 5434 -1654 6406
rect -1622 5434 -1600 6406
rect -1668 5420 -1600 5434
rect 1600 6406 1668 6420
rect 1600 5434 1622 6406
rect 1654 5434 1668 6406
rect 1600 5420 1668 5434
rect -1668 5222 -1600 5236
rect -1668 4250 -1654 5222
rect -1622 4250 -1600 5222
rect -1668 4236 -1600 4250
rect 1600 5222 1668 5236
rect 1600 4250 1622 5222
rect 1654 4250 1668 5222
rect 1600 4236 1668 4250
rect -1668 4038 -1600 4052
rect -1668 3066 -1654 4038
rect -1622 3066 -1600 4038
rect -1668 3052 -1600 3066
rect 1600 4038 1668 4052
rect 1600 3066 1622 4038
rect 1654 3066 1668 4038
rect 1600 3052 1668 3066
rect -1668 2854 -1600 2868
rect -1668 1882 -1654 2854
rect -1622 1882 -1600 2854
rect -1668 1868 -1600 1882
rect 1600 2854 1668 2868
rect 1600 1882 1622 2854
rect 1654 1882 1668 2854
rect 1600 1868 1668 1882
rect -1668 1670 -1600 1684
rect -1668 698 -1654 1670
rect -1622 698 -1600 1670
rect -1668 684 -1600 698
rect 1600 1670 1668 1684
rect 1600 698 1622 1670
rect 1654 698 1668 1670
rect 1600 684 1668 698
rect -1668 486 -1600 500
rect -1668 -486 -1654 486
rect -1622 -486 -1600 486
rect -1668 -500 -1600 -486
rect 1600 486 1668 500
rect 1600 -486 1622 486
rect 1654 -486 1668 486
rect 1600 -500 1668 -486
<< hvndiffc >>
rect -1654 13722 -1622 14694
rect 1622 13722 1654 14694
rect -1654 12538 -1622 13510
rect 1622 12538 1654 13510
rect -1654 11354 -1622 12326
rect 1622 11354 1654 12326
rect -1654 10170 -1622 11142
rect 1622 10170 1654 11142
rect -1654 8986 -1622 9958
rect 1622 8986 1654 9958
rect -1654 7802 -1622 8774
rect 1622 7802 1654 8774
rect -1654 6618 -1622 7590
rect 1622 6618 1654 7590
rect -1654 5434 -1622 6406
rect 1622 5434 1654 6406
rect -1654 4250 -1622 5222
rect 1622 4250 1654 5222
rect -1654 3066 -1622 4038
rect 1622 3066 1654 4038
rect -1654 1882 -1622 2854
rect 1622 1882 1654 2854
rect -1654 698 -1622 1670
rect 1622 698 1654 1670
rect -1654 -486 -1622 486
rect 1622 -486 1654 486
<< psubdiff >>
rect -1858 14881 1858 14895
rect -1858 14849 -1784 14881
rect 1784 14849 1858 14881
rect -1858 14835 1858 14849
rect -1858 14821 -1798 14835
rect -1858 -613 -1844 14821
rect -1812 -613 -1798 14821
rect 1798 14821 1858 14835
rect -1858 -627 -1798 -613
rect 1798 -613 1812 14821
rect 1844 -613 1858 14821
rect 1798 -627 1858 -613
rect -1858 -641 1858 -627
rect -1858 -673 -1784 -641
rect 1784 -673 1858 -641
rect -1858 -687 1858 -673
<< psubdiffcont >>
rect -1784 14849 1784 14881
rect -1844 -613 -1812 14821
rect 1812 -613 1844 14821
rect -1784 -673 1784 -641
<< poly >>
rect -1600 14768 1600 14782
rect -1600 14736 -1586 14768
rect 1586 14736 1600 14768
rect -1600 14708 1600 14736
rect -1600 13680 1600 13708
rect -1600 13648 -1586 13680
rect 1586 13648 1600 13680
rect -1600 13634 1600 13648
rect -1600 13584 1600 13598
rect -1600 13552 -1586 13584
rect 1586 13552 1600 13584
rect -1600 13524 1600 13552
rect -1600 12496 1600 12524
rect -1600 12464 -1586 12496
rect 1586 12464 1600 12496
rect -1600 12450 1600 12464
rect -1600 12400 1600 12414
rect -1600 12368 -1586 12400
rect 1586 12368 1600 12400
rect -1600 12340 1600 12368
rect -1600 11312 1600 11340
rect -1600 11280 -1586 11312
rect 1586 11280 1600 11312
rect -1600 11266 1600 11280
rect -1600 11216 1600 11230
rect -1600 11184 -1586 11216
rect 1586 11184 1600 11216
rect -1600 11156 1600 11184
rect -1600 10128 1600 10156
rect -1600 10096 -1586 10128
rect 1586 10096 1600 10128
rect -1600 10082 1600 10096
rect -1600 10032 1600 10046
rect -1600 10000 -1586 10032
rect 1586 10000 1600 10032
rect -1600 9972 1600 10000
rect -1600 8944 1600 8972
rect -1600 8912 -1586 8944
rect 1586 8912 1600 8944
rect -1600 8898 1600 8912
rect -1600 8848 1600 8862
rect -1600 8816 -1586 8848
rect 1586 8816 1600 8848
rect -1600 8788 1600 8816
rect -1600 7760 1600 7788
rect -1600 7728 -1586 7760
rect 1586 7728 1600 7760
rect -1600 7714 1600 7728
rect -1600 7664 1600 7678
rect -1600 7632 -1586 7664
rect 1586 7632 1600 7664
rect -1600 7604 1600 7632
rect -1600 6576 1600 6604
rect -1600 6544 -1586 6576
rect 1586 6544 1600 6576
rect -1600 6530 1600 6544
rect -1600 6480 1600 6494
rect -1600 6448 -1586 6480
rect 1586 6448 1600 6480
rect -1600 6420 1600 6448
rect -1600 5392 1600 5420
rect -1600 5360 -1586 5392
rect 1586 5360 1600 5392
rect -1600 5346 1600 5360
rect -1600 5296 1600 5310
rect -1600 5264 -1586 5296
rect 1586 5264 1600 5296
rect -1600 5236 1600 5264
rect -1600 4208 1600 4236
rect -1600 4176 -1586 4208
rect 1586 4176 1600 4208
rect -1600 4162 1600 4176
rect -1600 4112 1600 4126
rect -1600 4080 -1586 4112
rect 1586 4080 1600 4112
rect -1600 4052 1600 4080
rect -1600 3024 1600 3052
rect -1600 2992 -1586 3024
rect 1586 2992 1600 3024
rect -1600 2978 1600 2992
rect -1600 2928 1600 2942
rect -1600 2896 -1586 2928
rect 1586 2896 1600 2928
rect -1600 2868 1600 2896
rect -1600 1840 1600 1868
rect -1600 1808 -1586 1840
rect 1586 1808 1600 1840
rect -1600 1794 1600 1808
rect -1600 1744 1600 1758
rect -1600 1712 -1586 1744
rect 1586 1712 1600 1744
rect -1600 1684 1600 1712
rect -1600 656 1600 684
rect -1600 624 -1586 656
rect 1586 624 1600 656
rect -1600 610 1600 624
rect -1600 560 1600 574
rect -1600 528 -1586 560
rect 1586 528 1600 560
rect -1600 500 1600 528
rect -1600 -528 1600 -500
rect -1600 -560 -1586 -528
rect 1586 -560 1600 -528
rect -1600 -574 1600 -560
<< polycont >>
rect -1586 14736 1586 14768
rect -1586 13648 1586 13680
rect -1586 13552 1586 13584
rect -1586 12464 1586 12496
rect -1586 12368 1586 12400
rect -1586 11280 1586 11312
rect -1586 11184 1586 11216
rect -1586 10096 1586 10128
rect -1586 10000 1586 10032
rect -1586 8912 1586 8944
rect -1586 8816 1586 8848
rect -1586 7728 1586 7760
rect -1586 7632 1586 7664
rect -1586 6544 1586 6576
rect -1586 6448 1586 6480
rect -1586 5360 1586 5392
rect -1586 5264 1586 5296
rect -1586 4176 1586 4208
rect -1586 4080 1586 4112
rect -1586 2992 1586 3024
rect -1586 2896 1586 2928
rect -1586 1808 1586 1840
rect -1586 1712 1586 1744
rect -1586 624 1586 656
rect -1586 528 1586 560
rect -1586 -560 1586 -528
<< metal1 >>
rect -1854 14881 1854 14891
rect -1854 14849 -1784 14881
rect 1784 14849 1854 14881
rect -1854 14839 1854 14849
rect -1854 14821 -1802 14839
rect -1854 -613 -1844 14821
rect -1812 -613 -1802 14821
rect 1802 14821 1854 14839
rect -1854 -631 -1802 -613
rect 1802 -613 1812 14821
rect 1844 -613 1854 14821
rect 1802 -631 1854 -613
rect -1854 -641 1854 -631
rect -1854 -673 -1784 -641
rect 1784 -673 1854 -641
rect -1854 -683 1854 -673
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 5 l 16 nf 1 nx 1 dx 0.22 ny 13 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.2 glc 1 grc 1 gtc 1 gbc 1
<< end >>
