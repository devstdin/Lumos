magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 68 56 640 296
rect -26 -56 698 56
<< nmos >>
rect 162 160 188 270
rect 292 122 318 270
rect 394 122 420 270
rect 496 122 522 270
<< pmos >>
rect 184 412 210 580
rect 292 412 318 636
rect 394 412 420 636
rect 496 412 522 636
<< ndiff >>
rect 94 231 162 270
rect 94 199 108 231
rect 140 199 162 231
rect 94 160 162 199
rect 188 168 292 270
rect 188 160 227 168
rect 202 136 227 160
rect 259 136 292 168
rect 202 122 292 136
rect 318 122 394 270
rect 420 122 496 270
rect 522 236 614 270
rect 522 204 565 236
rect 597 204 614 236
rect 522 168 614 204
rect 522 136 565 168
rect 597 136 614 168
rect 522 122 614 136
<< pdiff >>
rect 224 622 292 636
rect 224 590 238 622
rect 270 590 292 622
rect 224 580 292 590
rect 116 566 184 580
rect 116 534 130 566
rect 162 534 184 566
rect 116 498 184 534
rect 116 466 130 498
rect 162 466 184 498
rect 116 412 184 466
rect 210 554 292 580
rect 210 522 238 554
rect 270 522 292 554
rect 210 486 292 522
rect 210 454 238 486
rect 270 454 292 486
rect 210 412 292 454
rect 318 622 394 636
rect 318 590 340 622
rect 372 590 394 622
rect 318 554 394 590
rect 318 522 340 554
rect 372 522 394 554
rect 318 486 394 522
rect 318 454 340 486
rect 372 454 394 486
rect 318 412 394 454
rect 420 622 496 636
rect 420 590 442 622
rect 474 590 496 622
rect 420 554 496 590
rect 420 522 442 554
rect 474 522 496 554
rect 420 412 496 522
rect 522 622 590 636
rect 522 590 544 622
rect 576 590 590 622
rect 522 554 590 590
rect 522 522 544 554
rect 576 522 590 554
rect 522 486 590 522
rect 522 454 544 486
rect 576 454 590 486
rect 522 412 590 454
<< ndiffc >>
rect 108 199 140 231
rect 227 136 259 168
rect 565 204 597 236
rect 565 136 597 168
<< pdiffc >>
rect 238 590 270 622
rect 130 534 162 566
rect 130 466 162 498
rect 238 522 270 554
rect 238 454 270 486
rect 340 590 372 622
rect 340 522 372 554
rect 340 454 372 486
rect 442 590 474 622
rect 442 522 474 554
rect 544 590 576 622
rect 544 522 576 554
rect 544 454 576 486
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 292 636 318 672
rect 394 636 420 672
rect 496 636 522 672
rect 184 580 210 616
rect 184 374 210 412
rect 292 374 318 412
rect 394 374 420 412
rect 496 374 522 412
rect 151 360 211 374
rect 151 328 165 360
rect 197 328 211 360
rect 151 314 211 328
rect 268 360 330 374
rect 268 328 282 360
rect 314 328 330 360
rect 268 314 330 328
rect 366 360 426 374
rect 366 328 380 360
rect 412 328 426 360
rect 366 314 426 328
rect 494 360 555 374
rect 494 328 509 360
rect 541 328 555 360
rect 494 314 555 328
rect 162 270 188 314
rect 292 270 318 314
rect 394 270 420 314
rect 496 270 522 314
rect 162 124 188 160
rect 292 86 318 122
rect 394 86 420 122
rect 496 86 522 122
<< polycont >>
rect 165 328 197 360
rect 282 328 314 360
rect 380 328 412 360
rect 509 328 541 360
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 228 622 280 712
rect 228 590 238 622
rect 270 590 280 622
rect 88 566 172 576
rect 88 534 130 566
rect 162 534 172 566
rect 88 498 172 534
rect 88 466 130 498
rect 162 466 172 498
rect 88 456 172 466
rect 228 554 280 590
rect 228 522 238 554
rect 270 522 280 554
rect 228 486 280 522
rect 88 246 122 456
rect 228 454 238 486
rect 270 454 280 486
rect 228 444 280 454
rect 330 622 382 632
rect 330 590 340 622
rect 372 590 382 622
rect 330 554 382 590
rect 330 522 340 554
rect 372 522 382 554
rect 330 486 382 522
rect 432 622 484 712
rect 432 590 442 622
rect 474 590 484 622
rect 432 554 484 590
rect 432 522 442 554
rect 474 522 484 554
rect 432 515 484 522
rect 534 622 626 632
rect 534 590 544 622
rect 576 590 626 622
rect 534 554 626 590
rect 534 522 544 554
rect 576 522 626 554
rect 330 454 340 486
rect 372 478 382 486
rect 534 486 626 522
rect 534 478 544 486
rect 372 454 544 478
rect 576 454 626 486
rect 330 440 626 454
rect 158 360 216 380
rect 158 328 165 360
rect 197 328 216 360
rect 158 295 216 328
rect 264 360 324 380
rect 264 328 282 360
rect 314 328 324 360
rect 264 295 324 328
rect 360 360 420 380
rect 360 328 380 360
rect 412 328 420 360
rect 360 295 420 328
rect 486 360 551 370
rect 486 328 509 360
rect 541 328 551 360
rect 486 318 551 328
rect 486 246 518 318
rect 592 246 626 440
rect 88 231 518 246
rect 88 199 108 231
rect 140 214 518 231
rect 555 236 626 246
rect 140 199 150 214
rect 88 189 150 199
rect 555 204 565 236
rect 597 204 626 236
rect 216 168 270 178
rect 216 136 227 168
rect 259 136 270 168
rect 216 44 270 136
rect 555 168 626 204
rect 555 136 565 168
rect 597 136 626 168
rect 555 126 626 136
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 158 295 216 380 0 FreeSans 400 0 0 0 A_N
port 2 nsew
flabel metal1 s 534 440 626 632 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 360 295 420 380 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel metal1 s 264 295 324 380 0 FreeSans 400 0 0 0 C
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 164924
string GDS_FILE 6_final.gds
string GDS_START 159126
<< end >>
