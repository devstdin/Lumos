magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2026 -2026 18026 9214
<< nwell >>
rect 3140 4750 12860 7214
<< pwell >>
rect -26 4372 16026 4492
rect -26 94 94 4372
rect 500 382 15500 4084
rect 15906 94 16026 4372
rect -26 -26 16026 94
<< hvnmos >>
rect 594 2258 2494 4058
rect 2570 2258 4470 4058
rect 4546 2258 6446 4058
rect 6522 2258 8422 4058
rect 8498 2258 10398 4058
rect 10474 2258 12374 4058
rect 12450 2258 14350 4058
rect 14426 2258 14526 4058
rect 14602 2258 14702 4058
rect 14778 2258 14878 4058
rect 14954 2258 15054 4058
rect 15130 2258 15230 4058
rect 15306 2258 15406 4058
rect 594 408 2494 2208
rect 2570 408 4470 2208
rect 4546 408 6446 2208
rect 6522 408 8422 2208
rect 8498 408 10398 2208
rect 10474 408 12374 2208
rect 12450 408 14350 2208
rect 14426 408 14526 2208
rect 14602 408 14702 2208
rect 14778 408 14878 2208
rect 14954 408 15054 2208
rect 15130 408 15230 2208
rect 15306 408 15406 2208
<< hvpmos >>
rect 3638 5282 3738 6682
rect 3814 5282 3914 6682
rect 3990 5282 4090 6682
rect 4166 5282 4266 6682
rect 4342 5282 4442 6682
rect 4518 5282 4618 6682
rect 4694 5282 4794 6682
rect 4870 5282 4970 6682
rect 5046 5282 5146 6682
rect 5222 5282 5322 6682
rect 5398 5282 5498 6682
rect 5574 5282 5674 6682
rect 5750 5282 5850 6682
rect 5926 5282 6026 6682
rect 6102 5282 6202 6682
rect 6278 5282 6378 6682
rect 6454 5282 6554 6682
rect 6630 5282 6730 6682
rect 6806 5282 6906 6682
rect 6982 5282 7082 6682
rect 7158 5282 7258 6682
rect 7334 5282 7434 6682
rect 7510 5282 7610 6682
rect 7686 5282 7786 6682
rect 7862 5282 7962 6682
rect 8038 5282 8138 6682
rect 8214 5282 8314 6682
rect 8390 5282 8490 6682
rect 8566 5282 8666 6682
rect 8742 5282 8842 6682
rect 8918 5282 9018 6682
rect 9094 5282 9194 6682
rect 9270 5282 9370 6682
rect 9446 5282 9546 6682
rect 9622 5282 9722 6682
rect 9798 5282 9898 6682
rect 9974 5282 10074 6682
rect 10150 5282 10250 6682
rect 10326 5282 10426 6682
rect 10502 5282 10602 6682
rect 10678 5282 10778 6682
rect 10854 5282 10954 6682
rect 11030 5282 11130 6682
rect 11206 5282 11306 6682
rect 11382 5282 11482 6682
rect 11558 5282 11658 6682
rect 11734 5282 11834 6682
rect 11910 5282 12010 6682
rect 12086 5282 12186 6682
rect 12262 5282 12362 6682
<< hvndiff >>
rect 526 4024 594 4058
rect 526 3992 540 4024
rect 572 3992 594 4024
rect 526 3956 594 3992
rect 526 3924 540 3956
rect 572 3924 594 3956
rect 526 3888 594 3924
rect 526 3856 540 3888
rect 572 3856 594 3888
rect 526 3820 594 3856
rect 526 3788 540 3820
rect 572 3788 594 3820
rect 526 3752 594 3788
rect 526 3720 540 3752
rect 572 3720 594 3752
rect 526 3684 594 3720
rect 526 3652 540 3684
rect 572 3652 594 3684
rect 526 3616 594 3652
rect 526 3584 540 3616
rect 572 3584 594 3616
rect 526 3548 594 3584
rect 526 3516 540 3548
rect 572 3516 594 3548
rect 526 3480 594 3516
rect 526 3448 540 3480
rect 572 3448 594 3480
rect 526 3412 594 3448
rect 526 3380 540 3412
rect 572 3380 594 3412
rect 526 3344 594 3380
rect 526 3312 540 3344
rect 572 3312 594 3344
rect 526 3276 594 3312
rect 526 3244 540 3276
rect 572 3244 594 3276
rect 526 3208 594 3244
rect 526 3176 540 3208
rect 572 3176 594 3208
rect 526 3140 594 3176
rect 526 3108 540 3140
rect 572 3108 594 3140
rect 526 3072 594 3108
rect 526 3040 540 3072
rect 572 3040 594 3072
rect 526 3004 594 3040
rect 526 2972 540 3004
rect 572 2972 594 3004
rect 526 2936 594 2972
rect 526 2904 540 2936
rect 572 2904 594 2936
rect 526 2868 594 2904
rect 526 2836 540 2868
rect 572 2836 594 2868
rect 526 2800 594 2836
rect 526 2768 540 2800
rect 572 2768 594 2800
rect 526 2732 594 2768
rect 526 2700 540 2732
rect 572 2700 594 2732
rect 526 2664 594 2700
rect 526 2632 540 2664
rect 572 2632 594 2664
rect 526 2596 594 2632
rect 526 2564 540 2596
rect 572 2564 594 2596
rect 526 2528 594 2564
rect 526 2496 540 2528
rect 572 2496 594 2528
rect 526 2460 594 2496
rect 526 2428 540 2460
rect 572 2428 594 2460
rect 526 2392 594 2428
rect 526 2360 540 2392
rect 572 2360 594 2392
rect 526 2324 594 2360
rect 526 2292 540 2324
rect 572 2292 594 2324
rect 526 2258 594 2292
rect 2494 4024 2570 4058
rect 2494 3992 2516 4024
rect 2548 3992 2570 4024
rect 2494 3956 2570 3992
rect 2494 3924 2516 3956
rect 2548 3924 2570 3956
rect 2494 3888 2570 3924
rect 2494 3856 2516 3888
rect 2548 3856 2570 3888
rect 2494 3820 2570 3856
rect 2494 3788 2516 3820
rect 2548 3788 2570 3820
rect 2494 3752 2570 3788
rect 2494 3720 2516 3752
rect 2548 3720 2570 3752
rect 2494 3684 2570 3720
rect 2494 3652 2516 3684
rect 2548 3652 2570 3684
rect 2494 3616 2570 3652
rect 2494 3584 2516 3616
rect 2548 3584 2570 3616
rect 2494 3548 2570 3584
rect 2494 3516 2516 3548
rect 2548 3516 2570 3548
rect 2494 3480 2570 3516
rect 2494 3448 2516 3480
rect 2548 3448 2570 3480
rect 2494 3412 2570 3448
rect 2494 3380 2516 3412
rect 2548 3380 2570 3412
rect 2494 3344 2570 3380
rect 2494 3312 2516 3344
rect 2548 3312 2570 3344
rect 2494 3276 2570 3312
rect 2494 3244 2516 3276
rect 2548 3244 2570 3276
rect 2494 3208 2570 3244
rect 2494 3176 2516 3208
rect 2548 3176 2570 3208
rect 2494 3140 2570 3176
rect 2494 3108 2516 3140
rect 2548 3108 2570 3140
rect 2494 3072 2570 3108
rect 2494 3040 2516 3072
rect 2548 3040 2570 3072
rect 2494 3004 2570 3040
rect 2494 2972 2516 3004
rect 2548 2972 2570 3004
rect 2494 2936 2570 2972
rect 2494 2904 2516 2936
rect 2548 2904 2570 2936
rect 2494 2868 2570 2904
rect 2494 2836 2516 2868
rect 2548 2836 2570 2868
rect 2494 2800 2570 2836
rect 2494 2768 2516 2800
rect 2548 2768 2570 2800
rect 2494 2732 2570 2768
rect 2494 2700 2516 2732
rect 2548 2700 2570 2732
rect 2494 2664 2570 2700
rect 2494 2632 2516 2664
rect 2548 2632 2570 2664
rect 2494 2596 2570 2632
rect 2494 2564 2516 2596
rect 2548 2564 2570 2596
rect 2494 2528 2570 2564
rect 2494 2496 2516 2528
rect 2548 2496 2570 2528
rect 2494 2460 2570 2496
rect 2494 2428 2516 2460
rect 2548 2428 2570 2460
rect 2494 2392 2570 2428
rect 2494 2360 2516 2392
rect 2548 2360 2570 2392
rect 2494 2324 2570 2360
rect 2494 2292 2516 2324
rect 2548 2292 2570 2324
rect 2494 2258 2570 2292
rect 4470 4024 4546 4058
rect 4470 3992 4492 4024
rect 4524 3992 4546 4024
rect 4470 3956 4546 3992
rect 4470 3924 4492 3956
rect 4524 3924 4546 3956
rect 4470 3888 4546 3924
rect 4470 3856 4492 3888
rect 4524 3856 4546 3888
rect 4470 3820 4546 3856
rect 4470 3788 4492 3820
rect 4524 3788 4546 3820
rect 4470 3752 4546 3788
rect 4470 3720 4492 3752
rect 4524 3720 4546 3752
rect 4470 3684 4546 3720
rect 4470 3652 4492 3684
rect 4524 3652 4546 3684
rect 4470 3616 4546 3652
rect 4470 3584 4492 3616
rect 4524 3584 4546 3616
rect 4470 3548 4546 3584
rect 4470 3516 4492 3548
rect 4524 3516 4546 3548
rect 4470 3480 4546 3516
rect 4470 3448 4492 3480
rect 4524 3448 4546 3480
rect 4470 3412 4546 3448
rect 4470 3380 4492 3412
rect 4524 3380 4546 3412
rect 4470 3344 4546 3380
rect 4470 3312 4492 3344
rect 4524 3312 4546 3344
rect 4470 3276 4546 3312
rect 4470 3244 4492 3276
rect 4524 3244 4546 3276
rect 4470 3208 4546 3244
rect 4470 3176 4492 3208
rect 4524 3176 4546 3208
rect 4470 3140 4546 3176
rect 4470 3108 4492 3140
rect 4524 3108 4546 3140
rect 4470 3072 4546 3108
rect 4470 3040 4492 3072
rect 4524 3040 4546 3072
rect 4470 3004 4546 3040
rect 4470 2972 4492 3004
rect 4524 2972 4546 3004
rect 4470 2936 4546 2972
rect 4470 2904 4492 2936
rect 4524 2904 4546 2936
rect 4470 2868 4546 2904
rect 4470 2836 4492 2868
rect 4524 2836 4546 2868
rect 4470 2800 4546 2836
rect 4470 2768 4492 2800
rect 4524 2768 4546 2800
rect 4470 2732 4546 2768
rect 4470 2700 4492 2732
rect 4524 2700 4546 2732
rect 4470 2664 4546 2700
rect 4470 2632 4492 2664
rect 4524 2632 4546 2664
rect 4470 2596 4546 2632
rect 4470 2564 4492 2596
rect 4524 2564 4546 2596
rect 4470 2528 4546 2564
rect 4470 2496 4492 2528
rect 4524 2496 4546 2528
rect 4470 2460 4546 2496
rect 4470 2428 4492 2460
rect 4524 2428 4546 2460
rect 4470 2392 4546 2428
rect 4470 2360 4492 2392
rect 4524 2360 4546 2392
rect 4470 2324 4546 2360
rect 4470 2292 4492 2324
rect 4524 2292 4546 2324
rect 4470 2258 4546 2292
rect 6446 4024 6522 4058
rect 6446 3992 6468 4024
rect 6500 3992 6522 4024
rect 6446 3956 6522 3992
rect 6446 3924 6468 3956
rect 6500 3924 6522 3956
rect 6446 3888 6522 3924
rect 6446 3856 6468 3888
rect 6500 3856 6522 3888
rect 6446 3820 6522 3856
rect 6446 3788 6468 3820
rect 6500 3788 6522 3820
rect 6446 3752 6522 3788
rect 6446 3720 6468 3752
rect 6500 3720 6522 3752
rect 6446 3684 6522 3720
rect 6446 3652 6468 3684
rect 6500 3652 6522 3684
rect 6446 3616 6522 3652
rect 6446 3584 6468 3616
rect 6500 3584 6522 3616
rect 6446 3548 6522 3584
rect 6446 3516 6468 3548
rect 6500 3516 6522 3548
rect 6446 3480 6522 3516
rect 6446 3448 6468 3480
rect 6500 3448 6522 3480
rect 6446 3412 6522 3448
rect 6446 3380 6468 3412
rect 6500 3380 6522 3412
rect 6446 3344 6522 3380
rect 6446 3312 6468 3344
rect 6500 3312 6522 3344
rect 6446 3276 6522 3312
rect 6446 3244 6468 3276
rect 6500 3244 6522 3276
rect 6446 3208 6522 3244
rect 6446 3176 6468 3208
rect 6500 3176 6522 3208
rect 6446 3140 6522 3176
rect 6446 3108 6468 3140
rect 6500 3108 6522 3140
rect 6446 3072 6522 3108
rect 6446 3040 6468 3072
rect 6500 3040 6522 3072
rect 6446 3004 6522 3040
rect 6446 2972 6468 3004
rect 6500 2972 6522 3004
rect 6446 2936 6522 2972
rect 6446 2904 6468 2936
rect 6500 2904 6522 2936
rect 6446 2868 6522 2904
rect 6446 2836 6468 2868
rect 6500 2836 6522 2868
rect 6446 2800 6522 2836
rect 6446 2768 6468 2800
rect 6500 2768 6522 2800
rect 6446 2732 6522 2768
rect 6446 2700 6468 2732
rect 6500 2700 6522 2732
rect 6446 2664 6522 2700
rect 6446 2632 6468 2664
rect 6500 2632 6522 2664
rect 6446 2596 6522 2632
rect 6446 2564 6468 2596
rect 6500 2564 6522 2596
rect 6446 2528 6522 2564
rect 6446 2496 6468 2528
rect 6500 2496 6522 2528
rect 6446 2460 6522 2496
rect 6446 2428 6468 2460
rect 6500 2428 6522 2460
rect 6446 2392 6522 2428
rect 6446 2360 6468 2392
rect 6500 2360 6522 2392
rect 6446 2324 6522 2360
rect 6446 2292 6468 2324
rect 6500 2292 6522 2324
rect 6446 2258 6522 2292
rect 8422 4024 8498 4058
rect 8422 3992 8444 4024
rect 8476 3992 8498 4024
rect 8422 3956 8498 3992
rect 8422 3924 8444 3956
rect 8476 3924 8498 3956
rect 8422 3888 8498 3924
rect 8422 3856 8444 3888
rect 8476 3856 8498 3888
rect 8422 3820 8498 3856
rect 8422 3788 8444 3820
rect 8476 3788 8498 3820
rect 8422 3752 8498 3788
rect 8422 3720 8444 3752
rect 8476 3720 8498 3752
rect 8422 3684 8498 3720
rect 8422 3652 8444 3684
rect 8476 3652 8498 3684
rect 8422 3616 8498 3652
rect 8422 3584 8444 3616
rect 8476 3584 8498 3616
rect 8422 3548 8498 3584
rect 8422 3516 8444 3548
rect 8476 3516 8498 3548
rect 8422 3480 8498 3516
rect 8422 3448 8444 3480
rect 8476 3448 8498 3480
rect 8422 3412 8498 3448
rect 8422 3380 8444 3412
rect 8476 3380 8498 3412
rect 8422 3344 8498 3380
rect 8422 3312 8444 3344
rect 8476 3312 8498 3344
rect 8422 3276 8498 3312
rect 8422 3244 8444 3276
rect 8476 3244 8498 3276
rect 8422 3208 8498 3244
rect 8422 3176 8444 3208
rect 8476 3176 8498 3208
rect 8422 3140 8498 3176
rect 8422 3108 8444 3140
rect 8476 3108 8498 3140
rect 8422 3072 8498 3108
rect 8422 3040 8444 3072
rect 8476 3040 8498 3072
rect 8422 3004 8498 3040
rect 8422 2972 8444 3004
rect 8476 2972 8498 3004
rect 8422 2936 8498 2972
rect 8422 2904 8444 2936
rect 8476 2904 8498 2936
rect 8422 2868 8498 2904
rect 8422 2836 8444 2868
rect 8476 2836 8498 2868
rect 8422 2800 8498 2836
rect 8422 2768 8444 2800
rect 8476 2768 8498 2800
rect 8422 2732 8498 2768
rect 8422 2700 8444 2732
rect 8476 2700 8498 2732
rect 8422 2664 8498 2700
rect 8422 2632 8444 2664
rect 8476 2632 8498 2664
rect 8422 2596 8498 2632
rect 8422 2564 8444 2596
rect 8476 2564 8498 2596
rect 8422 2528 8498 2564
rect 8422 2496 8444 2528
rect 8476 2496 8498 2528
rect 8422 2460 8498 2496
rect 8422 2428 8444 2460
rect 8476 2428 8498 2460
rect 8422 2392 8498 2428
rect 8422 2360 8444 2392
rect 8476 2360 8498 2392
rect 8422 2324 8498 2360
rect 8422 2292 8444 2324
rect 8476 2292 8498 2324
rect 8422 2258 8498 2292
rect 10398 4024 10474 4058
rect 10398 3992 10420 4024
rect 10452 3992 10474 4024
rect 10398 3956 10474 3992
rect 10398 3924 10420 3956
rect 10452 3924 10474 3956
rect 10398 3888 10474 3924
rect 10398 3856 10420 3888
rect 10452 3856 10474 3888
rect 10398 3820 10474 3856
rect 10398 3788 10420 3820
rect 10452 3788 10474 3820
rect 10398 3752 10474 3788
rect 10398 3720 10420 3752
rect 10452 3720 10474 3752
rect 10398 3684 10474 3720
rect 10398 3652 10420 3684
rect 10452 3652 10474 3684
rect 10398 3616 10474 3652
rect 10398 3584 10420 3616
rect 10452 3584 10474 3616
rect 10398 3548 10474 3584
rect 10398 3516 10420 3548
rect 10452 3516 10474 3548
rect 10398 3480 10474 3516
rect 10398 3448 10420 3480
rect 10452 3448 10474 3480
rect 10398 3412 10474 3448
rect 10398 3380 10420 3412
rect 10452 3380 10474 3412
rect 10398 3344 10474 3380
rect 10398 3312 10420 3344
rect 10452 3312 10474 3344
rect 10398 3276 10474 3312
rect 10398 3244 10420 3276
rect 10452 3244 10474 3276
rect 10398 3208 10474 3244
rect 10398 3176 10420 3208
rect 10452 3176 10474 3208
rect 10398 3140 10474 3176
rect 10398 3108 10420 3140
rect 10452 3108 10474 3140
rect 10398 3072 10474 3108
rect 10398 3040 10420 3072
rect 10452 3040 10474 3072
rect 10398 3004 10474 3040
rect 10398 2972 10420 3004
rect 10452 2972 10474 3004
rect 10398 2936 10474 2972
rect 10398 2904 10420 2936
rect 10452 2904 10474 2936
rect 10398 2868 10474 2904
rect 10398 2836 10420 2868
rect 10452 2836 10474 2868
rect 10398 2800 10474 2836
rect 10398 2768 10420 2800
rect 10452 2768 10474 2800
rect 10398 2732 10474 2768
rect 10398 2700 10420 2732
rect 10452 2700 10474 2732
rect 10398 2664 10474 2700
rect 10398 2632 10420 2664
rect 10452 2632 10474 2664
rect 10398 2596 10474 2632
rect 10398 2564 10420 2596
rect 10452 2564 10474 2596
rect 10398 2528 10474 2564
rect 10398 2496 10420 2528
rect 10452 2496 10474 2528
rect 10398 2460 10474 2496
rect 10398 2428 10420 2460
rect 10452 2428 10474 2460
rect 10398 2392 10474 2428
rect 10398 2360 10420 2392
rect 10452 2360 10474 2392
rect 10398 2324 10474 2360
rect 10398 2292 10420 2324
rect 10452 2292 10474 2324
rect 10398 2258 10474 2292
rect 12374 4024 12450 4058
rect 12374 3992 12396 4024
rect 12428 3992 12450 4024
rect 12374 3956 12450 3992
rect 12374 3924 12396 3956
rect 12428 3924 12450 3956
rect 12374 3888 12450 3924
rect 12374 3856 12396 3888
rect 12428 3856 12450 3888
rect 12374 3820 12450 3856
rect 12374 3788 12396 3820
rect 12428 3788 12450 3820
rect 12374 3752 12450 3788
rect 12374 3720 12396 3752
rect 12428 3720 12450 3752
rect 12374 3684 12450 3720
rect 12374 3652 12396 3684
rect 12428 3652 12450 3684
rect 12374 3616 12450 3652
rect 12374 3584 12396 3616
rect 12428 3584 12450 3616
rect 12374 3548 12450 3584
rect 12374 3516 12396 3548
rect 12428 3516 12450 3548
rect 12374 3480 12450 3516
rect 12374 3448 12396 3480
rect 12428 3448 12450 3480
rect 12374 3412 12450 3448
rect 12374 3380 12396 3412
rect 12428 3380 12450 3412
rect 12374 3344 12450 3380
rect 12374 3312 12396 3344
rect 12428 3312 12450 3344
rect 12374 3276 12450 3312
rect 12374 3244 12396 3276
rect 12428 3244 12450 3276
rect 12374 3208 12450 3244
rect 12374 3176 12396 3208
rect 12428 3176 12450 3208
rect 12374 3140 12450 3176
rect 12374 3108 12396 3140
rect 12428 3108 12450 3140
rect 12374 3072 12450 3108
rect 12374 3040 12396 3072
rect 12428 3040 12450 3072
rect 12374 3004 12450 3040
rect 12374 2972 12396 3004
rect 12428 2972 12450 3004
rect 12374 2936 12450 2972
rect 12374 2904 12396 2936
rect 12428 2904 12450 2936
rect 12374 2868 12450 2904
rect 12374 2836 12396 2868
rect 12428 2836 12450 2868
rect 12374 2800 12450 2836
rect 12374 2768 12396 2800
rect 12428 2768 12450 2800
rect 12374 2732 12450 2768
rect 12374 2700 12396 2732
rect 12428 2700 12450 2732
rect 12374 2664 12450 2700
rect 12374 2632 12396 2664
rect 12428 2632 12450 2664
rect 12374 2596 12450 2632
rect 12374 2564 12396 2596
rect 12428 2564 12450 2596
rect 12374 2528 12450 2564
rect 12374 2496 12396 2528
rect 12428 2496 12450 2528
rect 12374 2460 12450 2496
rect 12374 2428 12396 2460
rect 12428 2428 12450 2460
rect 12374 2392 12450 2428
rect 12374 2360 12396 2392
rect 12428 2360 12450 2392
rect 12374 2324 12450 2360
rect 12374 2292 12396 2324
rect 12428 2292 12450 2324
rect 12374 2258 12450 2292
rect 14350 4024 14426 4058
rect 14350 3992 14372 4024
rect 14404 3992 14426 4024
rect 14350 3956 14426 3992
rect 14350 3924 14372 3956
rect 14404 3924 14426 3956
rect 14350 3888 14426 3924
rect 14350 3856 14372 3888
rect 14404 3856 14426 3888
rect 14350 3820 14426 3856
rect 14350 3788 14372 3820
rect 14404 3788 14426 3820
rect 14350 3752 14426 3788
rect 14350 3720 14372 3752
rect 14404 3720 14426 3752
rect 14350 3684 14426 3720
rect 14350 3652 14372 3684
rect 14404 3652 14426 3684
rect 14350 3616 14426 3652
rect 14350 3584 14372 3616
rect 14404 3584 14426 3616
rect 14350 3548 14426 3584
rect 14350 3516 14372 3548
rect 14404 3516 14426 3548
rect 14350 3480 14426 3516
rect 14350 3448 14372 3480
rect 14404 3448 14426 3480
rect 14350 3412 14426 3448
rect 14350 3380 14372 3412
rect 14404 3380 14426 3412
rect 14350 3344 14426 3380
rect 14350 3312 14372 3344
rect 14404 3312 14426 3344
rect 14350 3276 14426 3312
rect 14350 3244 14372 3276
rect 14404 3244 14426 3276
rect 14350 3208 14426 3244
rect 14350 3176 14372 3208
rect 14404 3176 14426 3208
rect 14350 3140 14426 3176
rect 14350 3108 14372 3140
rect 14404 3108 14426 3140
rect 14350 3072 14426 3108
rect 14350 3040 14372 3072
rect 14404 3040 14426 3072
rect 14350 3004 14426 3040
rect 14350 2972 14372 3004
rect 14404 2972 14426 3004
rect 14350 2936 14426 2972
rect 14350 2904 14372 2936
rect 14404 2904 14426 2936
rect 14350 2868 14426 2904
rect 14350 2836 14372 2868
rect 14404 2836 14426 2868
rect 14350 2800 14426 2836
rect 14350 2768 14372 2800
rect 14404 2768 14426 2800
rect 14350 2732 14426 2768
rect 14350 2700 14372 2732
rect 14404 2700 14426 2732
rect 14350 2664 14426 2700
rect 14350 2632 14372 2664
rect 14404 2632 14426 2664
rect 14350 2596 14426 2632
rect 14350 2564 14372 2596
rect 14404 2564 14426 2596
rect 14350 2528 14426 2564
rect 14350 2496 14372 2528
rect 14404 2496 14426 2528
rect 14350 2460 14426 2496
rect 14350 2428 14372 2460
rect 14404 2428 14426 2460
rect 14350 2392 14426 2428
rect 14350 2360 14372 2392
rect 14404 2360 14426 2392
rect 14350 2324 14426 2360
rect 14350 2292 14372 2324
rect 14404 2292 14426 2324
rect 14350 2258 14426 2292
rect 14526 4024 14602 4058
rect 14526 3992 14548 4024
rect 14580 3992 14602 4024
rect 14526 3956 14602 3992
rect 14526 3924 14548 3956
rect 14580 3924 14602 3956
rect 14526 3888 14602 3924
rect 14526 3856 14548 3888
rect 14580 3856 14602 3888
rect 14526 3820 14602 3856
rect 14526 3788 14548 3820
rect 14580 3788 14602 3820
rect 14526 3752 14602 3788
rect 14526 3720 14548 3752
rect 14580 3720 14602 3752
rect 14526 3684 14602 3720
rect 14526 3652 14548 3684
rect 14580 3652 14602 3684
rect 14526 3616 14602 3652
rect 14526 3584 14548 3616
rect 14580 3584 14602 3616
rect 14526 3548 14602 3584
rect 14526 3516 14548 3548
rect 14580 3516 14602 3548
rect 14526 3480 14602 3516
rect 14526 3448 14548 3480
rect 14580 3448 14602 3480
rect 14526 3412 14602 3448
rect 14526 3380 14548 3412
rect 14580 3380 14602 3412
rect 14526 3344 14602 3380
rect 14526 3312 14548 3344
rect 14580 3312 14602 3344
rect 14526 3276 14602 3312
rect 14526 3244 14548 3276
rect 14580 3244 14602 3276
rect 14526 3208 14602 3244
rect 14526 3176 14548 3208
rect 14580 3176 14602 3208
rect 14526 3140 14602 3176
rect 14526 3108 14548 3140
rect 14580 3108 14602 3140
rect 14526 3072 14602 3108
rect 14526 3040 14548 3072
rect 14580 3040 14602 3072
rect 14526 3004 14602 3040
rect 14526 2972 14548 3004
rect 14580 2972 14602 3004
rect 14526 2936 14602 2972
rect 14526 2904 14548 2936
rect 14580 2904 14602 2936
rect 14526 2868 14602 2904
rect 14526 2836 14548 2868
rect 14580 2836 14602 2868
rect 14526 2800 14602 2836
rect 14526 2768 14548 2800
rect 14580 2768 14602 2800
rect 14526 2732 14602 2768
rect 14526 2700 14548 2732
rect 14580 2700 14602 2732
rect 14526 2664 14602 2700
rect 14526 2632 14548 2664
rect 14580 2632 14602 2664
rect 14526 2596 14602 2632
rect 14526 2564 14548 2596
rect 14580 2564 14602 2596
rect 14526 2528 14602 2564
rect 14526 2496 14548 2528
rect 14580 2496 14602 2528
rect 14526 2460 14602 2496
rect 14526 2428 14548 2460
rect 14580 2428 14602 2460
rect 14526 2392 14602 2428
rect 14526 2360 14548 2392
rect 14580 2360 14602 2392
rect 14526 2324 14602 2360
rect 14526 2292 14548 2324
rect 14580 2292 14602 2324
rect 14526 2258 14602 2292
rect 14702 4024 14778 4058
rect 14702 3992 14724 4024
rect 14756 3992 14778 4024
rect 14702 3956 14778 3992
rect 14702 3924 14724 3956
rect 14756 3924 14778 3956
rect 14702 3888 14778 3924
rect 14702 3856 14724 3888
rect 14756 3856 14778 3888
rect 14702 3820 14778 3856
rect 14702 3788 14724 3820
rect 14756 3788 14778 3820
rect 14702 3752 14778 3788
rect 14702 3720 14724 3752
rect 14756 3720 14778 3752
rect 14702 3684 14778 3720
rect 14702 3652 14724 3684
rect 14756 3652 14778 3684
rect 14702 3616 14778 3652
rect 14702 3584 14724 3616
rect 14756 3584 14778 3616
rect 14702 3548 14778 3584
rect 14702 3516 14724 3548
rect 14756 3516 14778 3548
rect 14702 3480 14778 3516
rect 14702 3448 14724 3480
rect 14756 3448 14778 3480
rect 14702 3412 14778 3448
rect 14702 3380 14724 3412
rect 14756 3380 14778 3412
rect 14702 3344 14778 3380
rect 14702 3312 14724 3344
rect 14756 3312 14778 3344
rect 14702 3276 14778 3312
rect 14702 3244 14724 3276
rect 14756 3244 14778 3276
rect 14702 3208 14778 3244
rect 14702 3176 14724 3208
rect 14756 3176 14778 3208
rect 14702 3140 14778 3176
rect 14702 3108 14724 3140
rect 14756 3108 14778 3140
rect 14702 3072 14778 3108
rect 14702 3040 14724 3072
rect 14756 3040 14778 3072
rect 14702 3004 14778 3040
rect 14702 2972 14724 3004
rect 14756 2972 14778 3004
rect 14702 2936 14778 2972
rect 14702 2904 14724 2936
rect 14756 2904 14778 2936
rect 14702 2868 14778 2904
rect 14702 2836 14724 2868
rect 14756 2836 14778 2868
rect 14702 2800 14778 2836
rect 14702 2768 14724 2800
rect 14756 2768 14778 2800
rect 14702 2732 14778 2768
rect 14702 2700 14724 2732
rect 14756 2700 14778 2732
rect 14702 2664 14778 2700
rect 14702 2632 14724 2664
rect 14756 2632 14778 2664
rect 14702 2596 14778 2632
rect 14702 2564 14724 2596
rect 14756 2564 14778 2596
rect 14702 2528 14778 2564
rect 14702 2496 14724 2528
rect 14756 2496 14778 2528
rect 14702 2460 14778 2496
rect 14702 2428 14724 2460
rect 14756 2428 14778 2460
rect 14702 2392 14778 2428
rect 14702 2360 14724 2392
rect 14756 2360 14778 2392
rect 14702 2324 14778 2360
rect 14702 2292 14724 2324
rect 14756 2292 14778 2324
rect 14702 2258 14778 2292
rect 14878 4024 14954 4058
rect 14878 3992 14900 4024
rect 14932 3992 14954 4024
rect 14878 3956 14954 3992
rect 14878 3924 14900 3956
rect 14932 3924 14954 3956
rect 14878 3888 14954 3924
rect 14878 3856 14900 3888
rect 14932 3856 14954 3888
rect 14878 3820 14954 3856
rect 14878 3788 14900 3820
rect 14932 3788 14954 3820
rect 14878 3752 14954 3788
rect 14878 3720 14900 3752
rect 14932 3720 14954 3752
rect 14878 3684 14954 3720
rect 14878 3652 14900 3684
rect 14932 3652 14954 3684
rect 14878 3616 14954 3652
rect 14878 3584 14900 3616
rect 14932 3584 14954 3616
rect 14878 3548 14954 3584
rect 14878 3516 14900 3548
rect 14932 3516 14954 3548
rect 14878 3480 14954 3516
rect 14878 3448 14900 3480
rect 14932 3448 14954 3480
rect 14878 3412 14954 3448
rect 14878 3380 14900 3412
rect 14932 3380 14954 3412
rect 14878 3344 14954 3380
rect 14878 3312 14900 3344
rect 14932 3312 14954 3344
rect 14878 3276 14954 3312
rect 14878 3244 14900 3276
rect 14932 3244 14954 3276
rect 14878 3208 14954 3244
rect 14878 3176 14900 3208
rect 14932 3176 14954 3208
rect 14878 3140 14954 3176
rect 14878 3108 14900 3140
rect 14932 3108 14954 3140
rect 14878 3072 14954 3108
rect 14878 3040 14900 3072
rect 14932 3040 14954 3072
rect 14878 3004 14954 3040
rect 14878 2972 14900 3004
rect 14932 2972 14954 3004
rect 14878 2936 14954 2972
rect 14878 2904 14900 2936
rect 14932 2904 14954 2936
rect 14878 2868 14954 2904
rect 14878 2836 14900 2868
rect 14932 2836 14954 2868
rect 14878 2800 14954 2836
rect 14878 2768 14900 2800
rect 14932 2768 14954 2800
rect 14878 2732 14954 2768
rect 14878 2700 14900 2732
rect 14932 2700 14954 2732
rect 14878 2664 14954 2700
rect 14878 2632 14900 2664
rect 14932 2632 14954 2664
rect 14878 2596 14954 2632
rect 14878 2564 14900 2596
rect 14932 2564 14954 2596
rect 14878 2528 14954 2564
rect 14878 2496 14900 2528
rect 14932 2496 14954 2528
rect 14878 2460 14954 2496
rect 14878 2428 14900 2460
rect 14932 2428 14954 2460
rect 14878 2392 14954 2428
rect 14878 2360 14900 2392
rect 14932 2360 14954 2392
rect 14878 2324 14954 2360
rect 14878 2292 14900 2324
rect 14932 2292 14954 2324
rect 14878 2258 14954 2292
rect 15054 4024 15130 4058
rect 15054 3992 15076 4024
rect 15108 3992 15130 4024
rect 15054 3956 15130 3992
rect 15054 3924 15076 3956
rect 15108 3924 15130 3956
rect 15054 3888 15130 3924
rect 15054 3856 15076 3888
rect 15108 3856 15130 3888
rect 15054 3820 15130 3856
rect 15054 3788 15076 3820
rect 15108 3788 15130 3820
rect 15054 3752 15130 3788
rect 15054 3720 15076 3752
rect 15108 3720 15130 3752
rect 15054 3684 15130 3720
rect 15054 3652 15076 3684
rect 15108 3652 15130 3684
rect 15054 3616 15130 3652
rect 15054 3584 15076 3616
rect 15108 3584 15130 3616
rect 15054 3548 15130 3584
rect 15054 3516 15076 3548
rect 15108 3516 15130 3548
rect 15054 3480 15130 3516
rect 15054 3448 15076 3480
rect 15108 3448 15130 3480
rect 15054 3412 15130 3448
rect 15054 3380 15076 3412
rect 15108 3380 15130 3412
rect 15054 3344 15130 3380
rect 15054 3312 15076 3344
rect 15108 3312 15130 3344
rect 15054 3276 15130 3312
rect 15054 3244 15076 3276
rect 15108 3244 15130 3276
rect 15054 3208 15130 3244
rect 15054 3176 15076 3208
rect 15108 3176 15130 3208
rect 15054 3140 15130 3176
rect 15054 3108 15076 3140
rect 15108 3108 15130 3140
rect 15054 3072 15130 3108
rect 15054 3040 15076 3072
rect 15108 3040 15130 3072
rect 15054 3004 15130 3040
rect 15054 2972 15076 3004
rect 15108 2972 15130 3004
rect 15054 2936 15130 2972
rect 15054 2904 15076 2936
rect 15108 2904 15130 2936
rect 15054 2868 15130 2904
rect 15054 2836 15076 2868
rect 15108 2836 15130 2868
rect 15054 2800 15130 2836
rect 15054 2768 15076 2800
rect 15108 2768 15130 2800
rect 15054 2732 15130 2768
rect 15054 2700 15076 2732
rect 15108 2700 15130 2732
rect 15054 2664 15130 2700
rect 15054 2632 15076 2664
rect 15108 2632 15130 2664
rect 15054 2596 15130 2632
rect 15054 2564 15076 2596
rect 15108 2564 15130 2596
rect 15054 2528 15130 2564
rect 15054 2496 15076 2528
rect 15108 2496 15130 2528
rect 15054 2460 15130 2496
rect 15054 2428 15076 2460
rect 15108 2428 15130 2460
rect 15054 2392 15130 2428
rect 15054 2360 15076 2392
rect 15108 2360 15130 2392
rect 15054 2324 15130 2360
rect 15054 2292 15076 2324
rect 15108 2292 15130 2324
rect 15054 2258 15130 2292
rect 15230 4024 15306 4058
rect 15230 3992 15252 4024
rect 15284 3992 15306 4024
rect 15230 3956 15306 3992
rect 15230 3924 15252 3956
rect 15284 3924 15306 3956
rect 15230 3888 15306 3924
rect 15230 3856 15252 3888
rect 15284 3856 15306 3888
rect 15230 3820 15306 3856
rect 15230 3788 15252 3820
rect 15284 3788 15306 3820
rect 15230 3752 15306 3788
rect 15230 3720 15252 3752
rect 15284 3720 15306 3752
rect 15230 3684 15306 3720
rect 15230 3652 15252 3684
rect 15284 3652 15306 3684
rect 15230 3616 15306 3652
rect 15230 3584 15252 3616
rect 15284 3584 15306 3616
rect 15230 3548 15306 3584
rect 15230 3516 15252 3548
rect 15284 3516 15306 3548
rect 15230 3480 15306 3516
rect 15230 3448 15252 3480
rect 15284 3448 15306 3480
rect 15230 3412 15306 3448
rect 15230 3380 15252 3412
rect 15284 3380 15306 3412
rect 15230 3344 15306 3380
rect 15230 3312 15252 3344
rect 15284 3312 15306 3344
rect 15230 3276 15306 3312
rect 15230 3244 15252 3276
rect 15284 3244 15306 3276
rect 15230 3208 15306 3244
rect 15230 3176 15252 3208
rect 15284 3176 15306 3208
rect 15230 3140 15306 3176
rect 15230 3108 15252 3140
rect 15284 3108 15306 3140
rect 15230 3072 15306 3108
rect 15230 3040 15252 3072
rect 15284 3040 15306 3072
rect 15230 3004 15306 3040
rect 15230 2972 15252 3004
rect 15284 2972 15306 3004
rect 15230 2936 15306 2972
rect 15230 2904 15252 2936
rect 15284 2904 15306 2936
rect 15230 2868 15306 2904
rect 15230 2836 15252 2868
rect 15284 2836 15306 2868
rect 15230 2800 15306 2836
rect 15230 2768 15252 2800
rect 15284 2768 15306 2800
rect 15230 2732 15306 2768
rect 15230 2700 15252 2732
rect 15284 2700 15306 2732
rect 15230 2664 15306 2700
rect 15230 2632 15252 2664
rect 15284 2632 15306 2664
rect 15230 2596 15306 2632
rect 15230 2564 15252 2596
rect 15284 2564 15306 2596
rect 15230 2528 15306 2564
rect 15230 2496 15252 2528
rect 15284 2496 15306 2528
rect 15230 2460 15306 2496
rect 15230 2428 15252 2460
rect 15284 2428 15306 2460
rect 15230 2392 15306 2428
rect 15230 2360 15252 2392
rect 15284 2360 15306 2392
rect 15230 2324 15306 2360
rect 15230 2292 15252 2324
rect 15284 2292 15306 2324
rect 15230 2258 15306 2292
rect 15406 4024 15474 4058
rect 15406 3992 15428 4024
rect 15460 3992 15474 4024
rect 15406 3956 15474 3992
rect 15406 3924 15428 3956
rect 15460 3924 15474 3956
rect 15406 3888 15474 3924
rect 15406 3856 15428 3888
rect 15460 3856 15474 3888
rect 15406 3820 15474 3856
rect 15406 3788 15428 3820
rect 15460 3788 15474 3820
rect 15406 3752 15474 3788
rect 15406 3720 15428 3752
rect 15460 3720 15474 3752
rect 15406 3684 15474 3720
rect 15406 3652 15428 3684
rect 15460 3652 15474 3684
rect 15406 3616 15474 3652
rect 15406 3584 15428 3616
rect 15460 3584 15474 3616
rect 15406 3548 15474 3584
rect 15406 3516 15428 3548
rect 15460 3516 15474 3548
rect 15406 3480 15474 3516
rect 15406 3448 15428 3480
rect 15460 3448 15474 3480
rect 15406 3412 15474 3448
rect 15406 3380 15428 3412
rect 15460 3380 15474 3412
rect 15406 3344 15474 3380
rect 15406 3312 15428 3344
rect 15460 3312 15474 3344
rect 15406 3276 15474 3312
rect 15406 3244 15428 3276
rect 15460 3244 15474 3276
rect 15406 3208 15474 3244
rect 15406 3176 15428 3208
rect 15460 3176 15474 3208
rect 15406 3140 15474 3176
rect 15406 3108 15428 3140
rect 15460 3108 15474 3140
rect 15406 3072 15474 3108
rect 15406 3040 15428 3072
rect 15460 3040 15474 3072
rect 15406 3004 15474 3040
rect 15406 2972 15428 3004
rect 15460 2972 15474 3004
rect 15406 2936 15474 2972
rect 15406 2904 15428 2936
rect 15460 2904 15474 2936
rect 15406 2868 15474 2904
rect 15406 2836 15428 2868
rect 15460 2836 15474 2868
rect 15406 2800 15474 2836
rect 15406 2768 15428 2800
rect 15460 2768 15474 2800
rect 15406 2732 15474 2768
rect 15406 2700 15428 2732
rect 15460 2700 15474 2732
rect 15406 2664 15474 2700
rect 15406 2632 15428 2664
rect 15460 2632 15474 2664
rect 15406 2596 15474 2632
rect 15406 2564 15428 2596
rect 15460 2564 15474 2596
rect 15406 2528 15474 2564
rect 15406 2496 15428 2528
rect 15460 2496 15474 2528
rect 15406 2460 15474 2496
rect 15406 2428 15428 2460
rect 15460 2428 15474 2460
rect 15406 2392 15474 2428
rect 15406 2360 15428 2392
rect 15460 2360 15474 2392
rect 15406 2324 15474 2360
rect 15406 2292 15428 2324
rect 15460 2292 15474 2324
rect 15406 2258 15474 2292
rect 526 2174 594 2208
rect 526 2142 540 2174
rect 572 2142 594 2174
rect 526 2106 594 2142
rect 526 2074 540 2106
rect 572 2074 594 2106
rect 526 2038 594 2074
rect 526 2006 540 2038
rect 572 2006 594 2038
rect 526 1970 594 2006
rect 526 1938 540 1970
rect 572 1938 594 1970
rect 526 1902 594 1938
rect 526 1870 540 1902
rect 572 1870 594 1902
rect 526 1834 594 1870
rect 526 1802 540 1834
rect 572 1802 594 1834
rect 526 1766 594 1802
rect 526 1734 540 1766
rect 572 1734 594 1766
rect 526 1698 594 1734
rect 526 1666 540 1698
rect 572 1666 594 1698
rect 526 1630 594 1666
rect 526 1598 540 1630
rect 572 1598 594 1630
rect 526 1562 594 1598
rect 526 1530 540 1562
rect 572 1530 594 1562
rect 526 1494 594 1530
rect 526 1462 540 1494
rect 572 1462 594 1494
rect 526 1426 594 1462
rect 526 1394 540 1426
rect 572 1394 594 1426
rect 526 1358 594 1394
rect 526 1326 540 1358
rect 572 1326 594 1358
rect 526 1290 594 1326
rect 526 1258 540 1290
rect 572 1258 594 1290
rect 526 1222 594 1258
rect 526 1190 540 1222
rect 572 1190 594 1222
rect 526 1154 594 1190
rect 526 1122 540 1154
rect 572 1122 594 1154
rect 526 1086 594 1122
rect 526 1054 540 1086
rect 572 1054 594 1086
rect 526 1018 594 1054
rect 526 986 540 1018
rect 572 986 594 1018
rect 526 950 594 986
rect 526 918 540 950
rect 572 918 594 950
rect 526 882 594 918
rect 526 850 540 882
rect 572 850 594 882
rect 526 814 594 850
rect 526 782 540 814
rect 572 782 594 814
rect 526 746 594 782
rect 526 714 540 746
rect 572 714 594 746
rect 526 678 594 714
rect 526 646 540 678
rect 572 646 594 678
rect 526 610 594 646
rect 526 578 540 610
rect 572 578 594 610
rect 526 542 594 578
rect 526 510 540 542
rect 572 510 594 542
rect 526 474 594 510
rect 526 442 540 474
rect 572 442 594 474
rect 526 408 594 442
rect 2494 2174 2570 2208
rect 2494 2142 2516 2174
rect 2548 2142 2570 2174
rect 2494 2106 2570 2142
rect 2494 2074 2516 2106
rect 2548 2074 2570 2106
rect 2494 2038 2570 2074
rect 2494 2006 2516 2038
rect 2548 2006 2570 2038
rect 2494 1970 2570 2006
rect 2494 1938 2516 1970
rect 2548 1938 2570 1970
rect 2494 1902 2570 1938
rect 2494 1870 2516 1902
rect 2548 1870 2570 1902
rect 2494 1834 2570 1870
rect 2494 1802 2516 1834
rect 2548 1802 2570 1834
rect 2494 1766 2570 1802
rect 2494 1734 2516 1766
rect 2548 1734 2570 1766
rect 2494 1698 2570 1734
rect 2494 1666 2516 1698
rect 2548 1666 2570 1698
rect 2494 1630 2570 1666
rect 2494 1598 2516 1630
rect 2548 1598 2570 1630
rect 2494 1562 2570 1598
rect 2494 1530 2516 1562
rect 2548 1530 2570 1562
rect 2494 1494 2570 1530
rect 2494 1462 2516 1494
rect 2548 1462 2570 1494
rect 2494 1426 2570 1462
rect 2494 1394 2516 1426
rect 2548 1394 2570 1426
rect 2494 1358 2570 1394
rect 2494 1326 2516 1358
rect 2548 1326 2570 1358
rect 2494 1290 2570 1326
rect 2494 1258 2516 1290
rect 2548 1258 2570 1290
rect 2494 1222 2570 1258
rect 2494 1190 2516 1222
rect 2548 1190 2570 1222
rect 2494 1154 2570 1190
rect 2494 1122 2516 1154
rect 2548 1122 2570 1154
rect 2494 1086 2570 1122
rect 2494 1054 2516 1086
rect 2548 1054 2570 1086
rect 2494 1018 2570 1054
rect 2494 986 2516 1018
rect 2548 986 2570 1018
rect 2494 950 2570 986
rect 2494 918 2516 950
rect 2548 918 2570 950
rect 2494 882 2570 918
rect 2494 850 2516 882
rect 2548 850 2570 882
rect 2494 814 2570 850
rect 2494 782 2516 814
rect 2548 782 2570 814
rect 2494 746 2570 782
rect 2494 714 2516 746
rect 2548 714 2570 746
rect 2494 678 2570 714
rect 2494 646 2516 678
rect 2548 646 2570 678
rect 2494 610 2570 646
rect 2494 578 2516 610
rect 2548 578 2570 610
rect 2494 542 2570 578
rect 2494 510 2516 542
rect 2548 510 2570 542
rect 2494 474 2570 510
rect 2494 442 2516 474
rect 2548 442 2570 474
rect 2494 408 2570 442
rect 4470 2174 4546 2208
rect 4470 2142 4492 2174
rect 4524 2142 4546 2174
rect 4470 2106 4546 2142
rect 4470 2074 4492 2106
rect 4524 2074 4546 2106
rect 4470 2038 4546 2074
rect 4470 2006 4492 2038
rect 4524 2006 4546 2038
rect 4470 1970 4546 2006
rect 4470 1938 4492 1970
rect 4524 1938 4546 1970
rect 4470 1902 4546 1938
rect 4470 1870 4492 1902
rect 4524 1870 4546 1902
rect 4470 1834 4546 1870
rect 4470 1802 4492 1834
rect 4524 1802 4546 1834
rect 4470 1766 4546 1802
rect 4470 1734 4492 1766
rect 4524 1734 4546 1766
rect 4470 1698 4546 1734
rect 4470 1666 4492 1698
rect 4524 1666 4546 1698
rect 4470 1630 4546 1666
rect 4470 1598 4492 1630
rect 4524 1598 4546 1630
rect 4470 1562 4546 1598
rect 4470 1530 4492 1562
rect 4524 1530 4546 1562
rect 4470 1494 4546 1530
rect 4470 1462 4492 1494
rect 4524 1462 4546 1494
rect 4470 1426 4546 1462
rect 4470 1394 4492 1426
rect 4524 1394 4546 1426
rect 4470 1358 4546 1394
rect 4470 1326 4492 1358
rect 4524 1326 4546 1358
rect 4470 1290 4546 1326
rect 4470 1258 4492 1290
rect 4524 1258 4546 1290
rect 4470 1222 4546 1258
rect 4470 1190 4492 1222
rect 4524 1190 4546 1222
rect 4470 1154 4546 1190
rect 4470 1122 4492 1154
rect 4524 1122 4546 1154
rect 4470 1086 4546 1122
rect 4470 1054 4492 1086
rect 4524 1054 4546 1086
rect 4470 1018 4546 1054
rect 4470 986 4492 1018
rect 4524 986 4546 1018
rect 4470 950 4546 986
rect 4470 918 4492 950
rect 4524 918 4546 950
rect 4470 882 4546 918
rect 4470 850 4492 882
rect 4524 850 4546 882
rect 4470 814 4546 850
rect 4470 782 4492 814
rect 4524 782 4546 814
rect 4470 746 4546 782
rect 4470 714 4492 746
rect 4524 714 4546 746
rect 4470 678 4546 714
rect 4470 646 4492 678
rect 4524 646 4546 678
rect 4470 610 4546 646
rect 4470 578 4492 610
rect 4524 578 4546 610
rect 4470 542 4546 578
rect 4470 510 4492 542
rect 4524 510 4546 542
rect 4470 474 4546 510
rect 4470 442 4492 474
rect 4524 442 4546 474
rect 4470 408 4546 442
rect 6446 2174 6522 2208
rect 6446 2142 6468 2174
rect 6500 2142 6522 2174
rect 6446 2106 6522 2142
rect 6446 2074 6468 2106
rect 6500 2074 6522 2106
rect 6446 2038 6522 2074
rect 6446 2006 6468 2038
rect 6500 2006 6522 2038
rect 6446 1970 6522 2006
rect 6446 1938 6468 1970
rect 6500 1938 6522 1970
rect 6446 1902 6522 1938
rect 6446 1870 6468 1902
rect 6500 1870 6522 1902
rect 6446 1834 6522 1870
rect 6446 1802 6468 1834
rect 6500 1802 6522 1834
rect 6446 1766 6522 1802
rect 6446 1734 6468 1766
rect 6500 1734 6522 1766
rect 6446 1698 6522 1734
rect 6446 1666 6468 1698
rect 6500 1666 6522 1698
rect 6446 1630 6522 1666
rect 6446 1598 6468 1630
rect 6500 1598 6522 1630
rect 6446 1562 6522 1598
rect 6446 1530 6468 1562
rect 6500 1530 6522 1562
rect 6446 1494 6522 1530
rect 6446 1462 6468 1494
rect 6500 1462 6522 1494
rect 6446 1426 6522 1462
rect 6446 1394 6468 1426
rect 6500 1394 6522 1426
rect 6446 1358 6522 1394
rect 6446 1326 6468 1358
rect 6500 1326 6522 1358
rect 6446 1290 6522 1326
rect 6446 1258 6468 1290
rect 6500 1258 6522 1290
rect 6446 1222 6522 1258
rect 6446 1190 6468 1222
rect 6500 1190 6522 1222
rect 6446 1154 6522 1190
rect 6446 1122 6468 1154
rect 6500 1122 6522 1154
rect 6446 1086 6522 1122
rect 6446 1054 6468 1086
rect 6500 1054 6522 1086
rect 6446 1018 6522 1054
rect 6446 986 6468 1018
rect 6500 986 6522 1018
rect 6446 950 6522 986
rect 6446 918 6468 950
rect 6500 918 6522 950
rect 6446 882 6522 918
rect 6446 850 6468 882
rect 6500 850 6522 882
rect 6446 814 6522 850
rect 6446 782 6468 814
rect 6500 782 6522 814
rect 6446 746 6522 782
rect 6446 714 6468 746
rect 6500 714 6522 746
rect 6446 678 6522 714
rect 6446 646 6468 678
rect 6500 646 6522 678
rect 6446 610 6522 646
rect 6446 578 6468 610
rect 6500 578 6522 610
rect 6446 542 6522 578
rect 6446 510 6468 542
rect 6500 510 6522 542
rect 6446 474 6522 510
rect 6446 442 6468 474
rect 6500 442 6522 474
rect 6446 408 6522 442
rect 8422 2174 8498 2208
rect 8422 2142 8444 2174
rect 8476 2142 8498 2174
rect 8422 2106 8498 2142
rect 8422 2074 8444 2106
rect 8476 2074 8498 2106
rect 8422 2038 8498 2074
rect 8422 2006 8444 2038
rect 8476 2006 8498 2038
rect 8422 1970 8498 2006
rect 8422 1938 8444 1970
rect 8476 1938 8498 1970
rect 8422 1902 8498 1938
rect 8422 1870 8444 1902
rect 8476 1870 8498 1902
rect 8422 1834 8498 1870
rect 8422 1802 8444 1834
rect 8476 1802 8498 1834
rect 8422 1766 8498 1802
rect 8422 1734 8444 1766
rect 8476 1734 8498 1766
rect 8422 1698 8498 1734
rect 8422 1666 8444 1698
rect 8476 1666 8498 1698
rect 8422 1630 8498 1666
rect 8422 1598 8444 1630
rect 8476 1598 8498 1630
rect 8422 1562 8498 1598
rect 8422 1530 8444 1562
rect 8476 1530 8498 1562
rect 8422 1494 8498 1530
rect 8422 1462 8444 1494
rect 8476 1462 8498 1494
rect 8422 1426 8498 1462
rect 8422 1394 8444 1426
rect 8476 1394 8498 1426
rect 8422 1358 8498 1394
rect 8422 1326 8444 1358
rect 8476 1326 8498 1358
rect 8422 1290 8498 1326
rect 8422 1258 8444 1290
rect 8476 1258 8498 1290
rect 8422 1222 8498 1258
rect 8422 1190 8444 1222
rect 8476 1190 8498 1222
rect 8422 1154 8498 1190
rect 8422 1122 8444 1154
rect 8476 1122 8498 1154
rect 8422 1086 8498 1122
rect 8422 1054 8444 1086
rect 8476 1054 8498 1086
rect 8422 1018 8498 1054
rect 8422 986 8444 1018
rect 8476 986 8498 1018
rect 8422 950 8498 986
rect 8422 918 8444 950
rect 8476 918 8498 950
rect 8422 882 8498 918
rect 8422 850 8444 882
rect 8476 850 8498 882
rect 8422 814 8498 850
rect 8422 782 8444 814
rect 8476 782 8498 814
rect 8422 746 8498 782
rect 8422 714 8444 746
rect 8476 714 8498 746
rect 8422 678 8498 714
rect 8422 646 8444 678
rect 8476 646 8498 678
rect 8422 610 8498 646
rect 8422 578 8444 610
rect 8476 578 8498 610
rect 8422 542 8498 578
rect 8422 510 8444 542
rect 8476 510 8498 542
rect 8422 474 8498 510
rect 8422 442 8444 474
rect 8476 442 8498 474
rect 8422 408 8498 442
rect 10398 2174 10474 2208
rect 10398 2142 10420 2174
rect 10452 2142 10474 2174
rect 10398 2106 10474 2142
rect 10398 2074 10420 2106
rect 10452 2074 10474 2106
rect 10398 2038 10474 2074
rect 10398 2006 10420 2038
rect 10452 2006 10474 2038
rect 10398 1970 10474 2006
rect 10398 1938 10420 1970
rect 10452 1938 10474 1970
rect 10398 1902 10474 1938
rect 10398 1870 10420 1902
rect 10452 1870 10474 1902
rect 10398 1834 10474 1870
rect 10398 1802 10420 1834
rect 10452 1802 10474 1834
rect 10398 1766 10474 1802
rect 10398 1734 10420 1766
rect 10452 1734 10474 1766
rect 10398 1698 10474 1734
rect 10398 1666 10420 1698
rect 10452 1666 10474 1698
rect 10398 1630 10474 1666
rect 10398 1598 10420 1630
rect 10452 1598 10474 1630
rect 10398 1562 10474 1598
rect 10398 1530 10420 1562
rect 10452 1530 10474 1562
rect 10398 1494 10474 1530
rect 10398 1462 10420 1494
rect 10452 1462 10474 1494
rect 10398 1426 10474 1462
rect 10398 1394 10420 1426
rect 10452 1394 10474 1426
rect 10398 1358 10474 1394
rect 10398 1326 10420 1358
rect 10452 1326 10474 1358
rect 10398 1290 10474 1326
rect 10398 1258 10420 1290
rect 10452 1258 10474 1290
rect 10398 1222 10474 1258
rect 10398 1190 10420 1222
rect 10452 1190 10474 1222
rect 10398 1154 10474 1190
rect 10398 1122 10420 1154
rect 10452 1122 10474 1154
rect 10398 1086 10474 1122
rect 10398 1054 10420 1086
rect 10452 1054 10474 1086
rect 10398 1018 10474 1054
rect 10398 986 10420 1018
rect 10452 986 10474 1018
rect 10398 950 10474 986
rect 10398 918 10420 950
rect 10452 918 10474 950
rect 10398 882 10474 918
rect 10398 850 10420 882
rect 10452 850 10474 882
rect 10398 814 10474 850
rect 10398 782 10420 814
rect 10452 782 10474 814
rect 10398 746 10474 782
rect 10398 714 10420 746
rect 10452 714 10474 746
rect 10398 678 10474 714
rect 10398 646 10420 678
rect 10452 646 10474 678
rect 10398 610 10474 646
rect 10398 578 10420 610
rect 10452 578 10474 610
rect 10398 542 10474 578
rect 10398 510 10420 542
rect 10452 510 10474 542
rect 10398 474 10474 510
rect 10398 442 10420 474
rect 10452 442 10474 474
rect 10398 408 10474 442
rect 12374 2174 12450 2208
rect 12374 2142 12396 2174
rect 12428 2142 12450 2174
rect 12374 2106 12450 2142
rect 12374 2074 12396 2106
rect 12428 2074 12450 2106
rect 12374 2038 12450 2074
rect 12374 2006 12396 2038
rect 12428 2006 12450 2038
rect 12374 1970 12450 2006
rect 12374 1938 12396 1970
rect 12428 1938 12450 1970
rect 12374 1902 12450 1938
rect 12374 1870 12396 1902
rect 12428 1870 12450 1902
rect 12374 1834 12450 1870
rect 12374 1802 12396 1834
rect 12428 1802 12450 1834
rect 12374 1766 12450 1802
rect 12374 1734 12396 1766
rect 12428 1734 12450 1766
rect 12374 1698 12450 1734
rect 12374 1666 12396 1698
rect 12428 1666 12450 1698
rect 12374 1630 12450 1666
rect 12374 1598 12396 1630
rect 12428 1598 12450 1630
rect 12374 1562 12450 1598
rect 12374 1530 12396 1562
rect 12428 1530 12450 1562
rect 12374 1494 12450 1530
rect 12374 1462 12396 1494
rect 12428 1462 12450 1494
rect 12374 1426 12450 1462
rect 12374 1394 12396 1426
rect 12428 1394 12450 1426
rect 12374 1358 12450 1394
rect 12374 1326 12396 1358
rect 12428 1326 12450 1358
rect 12374 1290 12450 1326
rect 12374 1258 12396 1290
rect 12428 1258 12450 1290
rect 12374 1222 12450 1258
rect 12374 1190 12396 1222
rect 12428 1190 12450 1222
rect 12374 1154 12450 1190
rect 12374 1122 12396 1154
rect 12428 1122 12450 1154
rect 12374 1086 12450 1122
rect 12374 1054 12396 1086
rect 12428 1054 12450 1086
rect 12374 1018 12450 1054
rect 12374 986 12396 1018
rect 12428 986 12450 1018
rect 12374 950 12450 986
rect 12374 918 12396 950
rect 12428 918 12450 950
rect 12374 882 12450 918
rect 12374 850 12396 882
rect 12428 850 12450 882
rect 12374 814 12450 850
rect 12374 782 12396 814
rect 12428 782 12450 814
rect 12374 746 12450 782
rect 12374 714 12396 746
rect 12428 714 12450 746
rect 12374 678 12450 714
rect 12374 646 12396 678
rect 12428 646 12450 678
rect 12374 610 12450 646
rect 12374 578 12396 610
rect 12428 578 12450 610
rect 12374 542 12450 578
rect 12374 510 12396 542
rect 12428 510 12450 542
rect 12374 474 12450 510
rect 12374 442 12396 474
rect 12428 442 12450 474
rect 12374 408 12450 442
rect 14350 2174 14426 2208
rect 14350 2142 14372 2174
rect 14404 2142 14426 2174
rect 14350 2106 14426 2142
rect 14350 2074 14372 2106
rect 14404 2074 14426 2106
rect 14350 2038 14426 2074
rect 14350 2006 14372 2038
rect 14404 2006 14426 2038
rect 14350 1970 14426 2006
rect 14350 1938 14372 1970
rect 14404 1938 14426 1970
rect 14350 1902 14426 1938
rect 14350 1870 14372 1902
rect 14404 1870 14426 1902
rect 14350 1834 14426 1870
rect 14350 1802 14372 1834
rect 14404 1802 14426 1834
rect 14350 1766 14426 1802
rect 14350 1734 14372 1766
rect 14404 1734 14426 1766
rect 14350 1698 14426 1734
rect 14350 1666 14372 1698
rect 14404 1666 14426 1698
rect 14350 1630 14426 1666
rect 14350 1598 14372 1630
rect 14404 1598 14426 1630
rect 14350 1562 14426 1598
rect 14350 1530 14372 1562
rect 14404 1530 14426 1562
rect 14350 1494 14426 1530
rect 14350 1462 14372 1494
rect 14404 1462 14426 1494
rect 14350 1426 14426 1462
rect 14350 1394 14372 1426
rect 14404 1394 14426 1426
rect 14350 1358 14426 1394
rect 14350 1326 14372 1358
rect 14404 1326 14426 1358
rect 14350 1290 14426 1326
rect 14350 1258 14372 1290
rect 14404 1258 14426 1290
rect 14350 1222 14426 1258
rect 14350 1190 14372 1222
rect 14404 1190 14426 1222
rect 14350 1154 14426 1190
rect 14350 1122 14372 1154
rect 14404 1122 14426 1154
rect 14350 1086 14426 1122
rect 14350 1054 14372 1086
rect 14404 1054 14426 1086
rect 14350 1018 14426 1054
rect 14350 986 14372 1018
rect 14404 986 14426 1018
rect 14350 950 14426 986
rect 14350 918 14372 950
rect 14404 918 14426 950
rect 14350 882 14426 918
rect 14350 850 14372 882
rect 14404 850 14426 882
rect 14350 814 14426 850
rect 14350 782 14372 814
rect 14404 782 14426 814
rect 14350 746 14426 782
rect 14350 714 14372 746
rect 14404 714 14426 746
rect 14350 678 14426 714
rect 14350 646 14372 678
rect 14404 646 14426 678
rect 14350 610 14426 646
rect 14350 578 14372 610
rect 14404 578 14426 610
rect 14350 542 14426 578
rect 14350 510 14372 542
rect 14404 510 14426 542
rect 14350 474 14426 510
rect 14350 442 14372 474
rect 14404 442 14426 474
rect 14350 408 14426 442
rect 14526 2174 14602 2208
rect 14526 2142 14548 2174
rect 14580 2142 14602 2174
rect 14526 2106 14602 2142
rect 14526 2074 14548 2106
rect 14580 2074 14602 2106
rect 14526 2038 14602 2074
rect 14526 2006 14548 2038
rect 14580 2006 14602 2038
rect 14526 1970 14602 2006
rect 14526 1938 14548 1970
rect 14580 1938 14602 1970
rect 14526 1902 14602 1938
rect 14526 1870 14548 1902
rect 14580 1870 14602 1902
rect 14526 1834 14602 1870
rect 14526 1802 14548 1834
rect 14580 1802 14602 1834
rect 14526 1766 14602 1802
rect 14526 1734 14548 1766
rect 14580 1734 14602 1766
rect 14526 1698 14602 1734
rect 14526 1666 14548 1698
rect 14580 1666 14602 1698
rect 14526 1630 14602 1666
rect 14526 1598 14548 1630
rect 14580 1598 14602 1630
rect 14526 1562 14602 1598
rect 14526 1530 14548 1562
rect 14580 1530 14602 1562
rect 14526 1494 14602 1530
rect 14526 1462 14548 1494
rect 14580 1462 14602 1494
rect 14526 1426 14602 1462
rect 14526 1394 14548 1426
rect 14580 1394 14602 1426
rect 14526 1358 14602 1394
rect 14526 1326 14548 1358
rect 14580 1326 14602 1358
rect 14526 1290 14602 1326
rect 14526 1258 14548 1290
rect 14580 1258 14602 1290
rect 14526 1222 14602 1258
rect 14526 1190 14548 1222
rect 14580 1190 14602 1222
rect 14526 1154 14602 1190
rect 14526 1122 14548 1154
rect 14580 1122 14602 1154
rect 14526 1086 14602 1122
rect 14526 1054 14548 1086
rect 14580 1054 14602 1086
rect 14526 1018 14602 1054
rect 14526 986 14548 1018
rect 14580 986 14602 1018
rect 14526 950 14602 986
rect 14526 918 14548 950
rect 14580 918 14602 950
rect 14526 882 14602 918
rect 14526 850 14548 882
rect 14580 850 14602 882
rect 14526 814 14602 850
rect 14526 782 14548 814
rect 14580 782 14602 814
rect 14526 746 14602 782
rect 14526 714 14548 746
rect 14580 714 14602 746
rect 14526 678 14602 714
rect 14526 646 14548 678
rect 14580 646 14602 678
rect 14526 610 14602 646
rect 14526 578 14548 610
rect 14580 578 14602 610
rect 14526 542 14602 578
rect 14526 510 14548 542
rect 14580 510 14602 542
rect 14526 474 14602 510
rect 14526 442 14548 474
rect 14580 442 14602 474
rect 14526 408 14602 442
rect 14702 2174 14778 2208
rect 14702 2142 14724 2174
rect 14756 2142 14778 2174
rect 14702 2106 14778 2142
rect 14702 2074 14724 2106
rect 14756 2074 14778 2106
rect 14702 2038 14778 2074
rect 14702 2006 14724 2038
rect 14756 2006 14778 2038
rect 14702 1970 14778 2006
rect 14702 1938 14724 1970
rect 14756 1938 14778 1970
rect 14702 1902 14778 1938
rect 14702 1870 14724 1902
rect 14756 1870 14778 1902
rect 14702 1834 14778 1870
rect 14702 1802 14724 1834
rect 14756 1802 14778 1834
rect 14702 1766 14778 1802
rect 14702 1734 14724 1766
rect 14756 1734 14778 1766
rect 14702 1698 14778 1734
rect 14702 1666 14724 1698
rect 14756 1666 14778 1698
rect 14702 1630 14778 1666
rect 14702 1598 14724 1630
rect 14756 1598 14778 1630
rect 14702 1562 14778 1598
rect 14702 1530 14724 1562
rect 14756 1530 14778 1562
rect 14702 1494 14778 1530
rect 14702 1462 14724 1494
rect 14756 1462 14778 1494
rect 14702 1426 14778 1462
rect 14702 1394 14724 1426
rect 14756 1394 14778 1426
rect 14702 1358 14778 1394
rect 14702 1326 14724 1358
rect 14756 1326 14778 1358
rect 14702 1290 14778 1326
rect 14702 1258 14724 1290
rect 14756 1258 14778 1290
rect 14702 1222 14778 1258
rect 14702 1190 14724 1222
rect 14756 1190 14778 1222
rect 14702 1154 14778 1190
rect 14702 1122 14724 1154
rect 14756 1122 14778 1154
rect 14702 1086 14778 1122
rect 14702 1054 14724 1086
rect 14756 1054 14778 1086
rect 14702 1018 14778 1054
rect 14702 986 14724 1018
rect 14756 986 14778 1018
rect 14702 950 14778 986
rect 14702 918 14724 950
rect 14756 918 14778 950
rect 14702 882 14778 918
rect 14702 850 14724 882
rect 14756 850 14778 882
rect 14702 814 14778 850
rect 14702 782 14724 814
rect 14756 782 14778 814
rect 14702 746 14778 782
rect 14702 714 14724 746
rect 14756 714 14778 746
rect 14702 678 14778 714
rect 14702 646 14724 678
rect 14756 646 14778 678
rect 14702 610 14778 646
rect 14702 578 14724 610
rect 14756 578 14778 610
rect 14702 542 14778 578
rect 14702 510 14724 542
rect 14756 510 14778 542
rect 14702 474 14778 510
rect 14702 442 14724 474
rect 14756 442 14778 474
rect 14702 408 14778 442
rect 14878 2174 14954 2208
rect 14878 2142 14900 2174
rect 14932 2142 14954 2174
rect 14878 2106 14954 2142
rect 14878 2074 14900 2106
rect 14932 2074 14954 2106
rect 14878 2038 14954 2074
rect 14878 2006 14900 2038
rect 14932 2006 14954 2038
rect 14878 1970 14954 2006
rect 14878 1938 14900 1970
rect 14932 1938 14954 1970
rect 14878 1902 14954 1938
rect 14878 1870 14900 1902
rect 14932 1870 14954 1902
rect 14878 1834 14954 1870
rect 14878 1802 14900 1834
rect 14932 1802 14954 1834
rect 14878 1766 14954 1802
rect 14878 1734 14900 1766
rect 14932 1734 14954 1766
rect 14878 1698 14954 1734
rect 14878 1666 14900 1698
rect 14932 1666 14954 1698
rect 14878 1630 14954 1666
rect 14878 1598 14900 1630
rect 14932 1598 14954 1630
rect 14878 1562 14954 1598
rect 14878 1530 14900 1562
rect 14932 1530 14954 1562
rect 14878 1494 14954 1530
rect 14878 1462 14900 1494
rect 14932 1462 14954 1494
rect 14878 1426 14954 1462
rect 14878 1394 14900 1426
rect 14932 1394 14954 1426
rect 14878 1358 14954 1394
rect 14878 1326 14900 1358
rect 14932 1326 14954 1358
rect 14878 1290 14954 1326
rect 14878 1258 14900 1290
rect 14932 1258 14954 1290
rect 14878 1222 14954 1258
rect 14878 1190 14900 1222
rect 14932 1190 14954 1222
rect 14878 1154 14954 1190
rect 14878 1122 14900 1154
rect 14932 1122 14954 1154
rect 14878 1086 14954 1122
rect 14878 1054 14900 1086
rect 14932 1054 14954 1086
rect 14878 1018 14954 1054
rect 14878 986 14900 1018
rect 14932 986 14954 1018
rect 14878 950 14954 986
rect 14878 918 14900 950
rect 14932 918 14954 950
rect 14878 882 14954 918
rect 14878 850 14900 882
rect 14932 850 14954 882
rect 14878 814 14954 850
rect 14878 782 14900 814
rect 14932 782 14954 814
rect 14878 746 14954 782
rect 14878 714 14900 746
rect 14932 714 14954 746
rect 14878 678 14954 714
rect 14878 646 14900 678
rect 14932 646 14954 678
rect 14878 610 14954 646
rect 14878 578 14900 610
rect 14932 578 14954 610
rect 14878 542 14954 578
rect 14878 510 14900 542
rect 14932 510 14954 542
rect 14878 474 14954 510
rect 14878 442 14900 474
rect 14932 442 14954 474
rect 14878 408 14954 442
rect 15054 2174 15130 2208
rect 15054 2142 15076 2174
rect 15108 2142 15130 2174
rect 15054 2106 15130 2142
rect 15054 2074 15076 2106
rect 15108 2074 15130 2106
rect 15054 2038 15130 2074
rect 15054 2006 15076 2038
rect 15108 2006 15130 2038
rect 15054 1970 15130 2006
rect 15054 1938 15076 1970
rect 15108 1938 15130 1970
rect 15054 1902 15130 1938
rect 15054 1870 15076 1902
rect 15108 1870 15130 1902
rect 15054 1834 15130 1870
rect 15054 1802 15076 1834
rect 15108 1802 15130 1834
rect 15054 1766 15130 1802
rect 15054 1734 15076 1766
rect 15108 1734 15130 1766
rect 15054 1698 15130 1734
rect 15054 1666 15076 1698
rect 15108 1666 15130 1698
rect 15054 1630 15130 1666
rect 15054 1598 15076 1630
rect 15108 1598 15130 1630
rect 15054 1562 15130 1598
rect 15054 1530 15076 1562
rect 15108 1530 15130 1562
rect 15054 1494 15130 1530
rect 15054 1462 15076 1494
rect 15108 1462 15130 1494
rect 15054 1426 15130 1462
rect 15054 1394 15076 1426
rect 15108 1394 15130 1426
rect 15054 1358 15130 1394
rect 15054 1326 15076 1358
rect 15108 1326 15130 1358
rect 15054 1290 15130 1326
rect 15054 1258 15076 1290
rect 15108 1258 15130 1290
rect 15054 1222 15130 1258
rect 15054 1190 15076 1222
rect 15108 1190 15130 1222
rect 15054 1154 15130 1190
rect 15054 1122 15076 1154
rect 15108 1122 15130 1154
rect 15054 1086 15130 1122
rect 15054 1054 15076 1086
rect 15108 1054 15130 1086
rect 15054 1018 15130 1054
rect 15054 986 15076 1018
rect 15108 986 15130 1018
rect 15054 950 15130 986
rect 15054 918 15076 950
rect 15108 918 15130 950
rect 15054 882 15130 918
rect 15054 850 15076 882
rect 15108 850 15130 882
rect 15054 814 15130 850
rect 15054 782 15076 814
rect 15108 782 15130 814
rect 15054 746 15130 782
rect 15054 714 15076 746
rect 15108 714 15130 746
rect 15054 678 15130 714
rect 15054 646 15076 678
rect 15108 646 15130 678
rect 15054 610 15130 646
rect 15054 578 15076 610
rect 15108 578 15130 610
rect 15054 542 15130 578
rect 15054 510 15076 542
rect 15108 510 15130 542
rect 15054 474 15130 510
rect 15054 442 15076 474
rect 15108 442 15130 474
rect 15054 408 15130 442
rect 15230 2174 15306 2208
rect 15230 2142 15252 2174
rect 15284 2142 15306 2174
rect 15230 2106 15306 2142
rect 15230 2074 15252 2106
rect 15284 2074 15306 2106
rect 15230 2038 15306 2074
rect 15230 2006 15252 2038
rect 15284 2006 15306 2038
rect 15230 1970 15306 2006
rect 15230 1938 15252 1970
rect 15284 1938 15306 1970
rect 15230 1902 15306 1938
rect 15230 1870 15252 1902
rect 15284 1870 15306 1902
rect 15230 1834 15306 1870
rect 15230 1802 15252 1834
rect 15284 1802 15306 1834
rect 15230 1766 15306 1802
rect 15230 1734 15252 1766
rect 15284 1734 15306 1766
rect 15230 1698 15306 1734
rect 15230 1666 15252 1698
rect 15284 1666 15306 1698
rect 15230 1630 15306 1666
rect 15230 1598 15252 1630
rect 15284 1598 15306 1630
rect 15230 1562 15306 1598
rect 15230 1530 15252 1562
rect 15284 1530 15306 1562
rect 15230 1494 15306 1530
rect 15230 1462 15252 1494
rect 15284 1462 15306 1494
rect 15230 1426 15306 1462
rect 15230 1394 15252 1426
rect 15284 1394 15306 1426
rect 15230 1358 15306 1394
rect 15230 1326 15252 1358
rect 15284 1326 15306 1358
rect 15230 1290 15306 1326
rect 15230 1258 15252 1290
rect 15284 1258 15306 1290
rect 15230 1222 15306 1258
rect 15230 1190 15252 1222
rect 15284 1190 15306 1222
rect 15230 1154 15306 1190
rect 15230 1122 15252 1154
rect 15284 1122 15306 1154
rect 15230 1086 15306 1122
rect 15230 1054 15252 1086
rect 15284 1054 15306 1086
rect 15230 1018 15306 1054
rect 15230 986 15252 1018
rect 15284 986 15306 1018
rect 15230 950 15306 986
rect 15230 918 15252 950
rect 15284 918 15306 950
rect 15230 882 15306 918
rect 15230 850 15252 882
rect 15284 850 15306 882
rect 15230 814 15306 850
rect 15230 782 15252 814
rect 15284 782 15306 814
rect 15230 746 15306 782
rect 15230 714 15252 746
rect 15284 714 15306 746
rect 15230 678 15306 714
rect 15230 646 15252 678
rect 15284 646 15306 678
rect 15230 610 15306 646
rect 15230 578 15252 610
rect 15284 578 15306 610
rect 15230 542 15306 578
rect 15230 510 15252 542
rect 15284 510 15306 542
rect 15230 474 15306 510
rect 15230 442 15252 474
rect 15284 442 15306 474
rect 15230 408 15306 442
rect 15406 2174 15474 2208
rect 15406 2142 15428 2174
rect 15460 2142 15474 2174
rect 15406 2106 15474 2142
rect 15406 2074 15428 2106
rect 15460 2074 15474 2106
rect 15406 2038 15474 2074
rect 15406 2006 15428 2038
rect 15460 2006 15474 2038
rect 15406 1970 15474 2006
rect 15406 1938 15428 1970
rect 15460 1938 15474 1970
rect 15406 1902 15474 1938
rect 15406 1870 15428 1902
rect 15460 1870 15474 1902
rect 15406 1834 15474 1870
rect 15406 1802 15428 1834
rect 15460 1802 15474 1834
rect 15406 1766 15474 1802
rect 15406 1734 15428 1766
rect 15460 1734 15474 1766
rect 15406 1698 15474 1734
rect 15406 1666 15428 1698
rect 15460 1666 15474 1698
rect 15406 1630 15474 1666
rect 15406 1598 15428 1630
rect 15460 1598 15474 1630
rect 15406 1562 15474 1598
rect 15406 1530 15428 1562
rect 15460 1530 15474 1562
rect 15406 1494 15474 1530
rect 15406 1462 15428 1494
rect 15460 1462 15474 1494
rect 15406 1426 15474 1462
rect 15406 1394 15428 1426
rect 15460 1394 15474 1426
rect 15406 1358 15474 1394
rect 15406 1326 15428 1358
rect 15460 1326 15474 1358
rect 15406 1290 15474 1326
rect 15406 1258 15428 1290
rect 15460 1258 15474 1290
rect 15406 1222 15474 1258
rect 15406 1190 15428 1222
rect 15460 1190 15474 1222
rect 15406 1154 15474 1190
rect 15406 1122 15428 1154
rect 15460 1122 15474 1154
rect 15406 1086 15474 1122
rect 15406 1054 15428 1086
rect 15460 1054 15474 1086
rect 15406 1018 15474 1054
rect 15406 986 15428 1018
rect 15460 986 15474 1018
rect 15406 950 15474 986
rect 15406 918 15428 950
rect 15460 918 15474 950
rect 15406 882 15474 918
rect 15406 850 15428 882
rect 15460 850 15474 882
rect 15406 814 15474 850
rect 15406 782 15428 814
rect 15460 782 15474 814
rect 15406 746 15474 782
rect 15406 714 15428 746
rect 15460 714 15474 746
rect 15406 678 15474 714
rect 15406 646 15428 678
rect 15460 646 15474 678
rect 15406 610 15474 646
rect 15406 578 15428 610
rect 15460 578 15474 610
rect 15406 542 15474 578
rect 15406 510 15428 542
rect 15460 510 15474 542
rect 15406 474 15474 510
rect 15406 442 15428 474
rect 15460 442 15474 474
rect 15406 408 15474 442
<< hvpdiff >>
rect 3570 6644 3638 6682
rect 3570 6612 3584 6644
rect 3616 6612 3638 6644
rect 3570 6576 3638 6612
rect 3570 6544 3584 6576
rect 3616 6544 3638 6576
rect 3570 6508 3638 6544
rect 3570 6476 3584 6508
rect 3616 6476 3638 6508
rect 3570 6440 3638 6476
rect 3570 6408 3584 6440
rect 3616 6408 3638 6440
rect 3570 6372 3638 6408
rect 3570 6340 3584 6372
rect 3616 6340 3638 6372
rect 3570 6304 3638 6340
rect 3570 6272 3584 6304
rect 3616 6272 3638 6304
rect 3570 6236 3638 6272
rect 3570 6204 3584 6236
rect 3616 6204 3638 6236
rect 3570 6168 3638 6204
rect 3570 6136 3584 6168
rect 3616 6136 3638 6168
rect 3570 6100 3638 6136
rect 3570 6068 3584 6100
rect 3616 6068 3638 6100
rect 3570 6032 3638 6068
rect 3570 6000 3584 6032
rect 3616 6000 3638 6032
rect 3570 5964 3638 6000
rect 3570 5932 3584 5964
rect 3616 5932 3638 5964
rect 3570 5896 3638 5932
rect 3570 5864 3584 5896
rect 3616 5864 3638 5896
rect 3570 5828 3638 5864
rect 3570 5796 3584 5828
rect 3616 5796 3638 5828
rect 3570 5760 3638 5796
rect 3570 5728 3584 5760
rect 3616 5728 3638 5760
rect 3570 5692 3638 5728
rect 3570 5660 3584 5692
rect 3616 5660 3638 5692
rect 3570 5624 3638 5660
rect 3570 5592 3584 5624
rect 3616 5592 3638 5624
rect 3570 5556 3638 5592
rect 3570 5524 3584 5556
rect 3616 5524 3638 5556
rect 3570 5488 3638 5524
rect 3570 5456 3584 5488
rect 3616 5456 3638 5488
rect 3570 5420 3638 5456
rect 3570 5388 3584 5420
rect 3616 5388 3638 5420
rect 3570 5352 3638 5388
rect 3570 5320 3584 5352
rect 3616 5320 3638 5352
rect 3570 5282 3638 5320
rect 3738 6644 3814 6682
rect 3738 6612 3760 6644
rect 3792 6612 3814 6644
rect 3738 6576 3814 6612
rect 3738 6544 3760 6576
rect 3792 6544 3814 6576
rect 3738 6508 3814 6544
rect 3738 6476 3760 6508
rect 3792 6476 3814 6508
rect 3738 6440 3814 6476
rect 3738 6408 3760 6440
rect 3792 6408 3814 6440
rect 3738 6372 3814 6408
rect 3738 6340 3760 6372
rect 3792 6340 3814 6372
rect 3738 6304 3814 6340
rect 3738 6272 3760 6304
rect 3792 6272 3814 6304
rect 3738 6236 3814 6272
rect 3738 6204 3760 6236
rect 3792 6204 3814 6236
rect 3738 6168 3814 6204
rect 3738 6136 3760 6168
rect 3792 6136 3814 6168
rect 3738 6100 3814 6136
rect 3738 6068 3760 6100
rect 3792 6068 3814 6100
rect 3738 6032 3814 6068
rect 3738 6000 3760 6032
rect 3792 6000 3814 6032
rect 3738 5964 3814 6000
rect 3738 5932 3760 5964
rect 3792 5932 3814 5964
rect 3738 5896 3814 5932
rect 3738 5864 3760 5896
rect 3792 5864 3814 5896
rect 3738 5828 3814 5864
rect 3738 5796 3760 5828
rect 3792 5796 3814 5828
rect 3738 5760 3814 5796
rect 3738 5728 3760 5760
rect 3792 5728 3814 5760
rect 3738 5692 3814 5728
rect 3738 5660 3760 5692
rect 3792 5660 3814 5692
rect 3738 5624 3814 5660
rect 3738 5592 3760 5624
rect 3792 5592 3814 5624
rect 3738 5556 3814 5592
rect 3738 5524 3760 5556
rect 3792 5524 3814 5556
rect 3738 5488 3814 5524
rect 3738 5456 3760 5488
rect 3792 5456 3814 5488
rect 3738 5420 3814 5456
rect 3738 5388 3760 5420
rect 3792 5388 3814 5420
rect 3738 5352 3814 5388
rect 3738 5320 3760 5352
rect 3792 5320 3814 5352
rect 3738 5282 3814 5320
rect 3914 6644 3990 6682
rect 3914 6612 3936 6644
rect 3968 6612 3990 6644
rect 3914 6576 3990 6612
rect 3914 6544 3936 6576
rect 3968 6544 3990 6576
rect 3914 6508 3990 6544
rect 3914 6476 3936 6508
rect 3968 6476 3990 6508
rect 3914 6440 3990 6476
rect 3914 6408 3936 6440
rect 3968 6408 3990 6440
rect 3914 6372 3990 6408
rect 3914 6340 3936 6372
rect 3968 6340 3990 6372
rect 3914 6304 3990 6340
rect 3914 6272 3936 6304
rect 3968 6272 3990 6304
rect 3914 6236 3990 6272
rect 3914 6204 3936 6236
rect 3968 6204 3990 6236
rect 3914 6168 3990 6204
rect 3914 6136 3936 6168
rect 3968 6136 3990 6168
rect 3914 6100 3990 6136
rect 3914 6068 3936 6100
rect 3968 6068 3990 6100
rect 3914 6032 3990 6068
rect 3914 6000 3936 6032
rect 3968 6000 3990 6032
rect 3914 5964 3990 6000
rect 3914 5932 3936 5964
rect 3968 5932 3990 5964
rect 3914 5896 3990 5932
rect 3914 5864 3936 5896
rect 3968 5864 3990 5896
rect 3914 5828 3990 5864
rect 3914 5796 3936 5828
rect 3968 5796 3990 5828
rect 3914 5760 3990 5796
rect 3914 5728 3936 5760
rect 3968 5728 3990 5760
rect 3914 5692 3990 5728
rect 3914 5660 3936 5692
rect 3968 5660 3990 5692
rect 3914 5624 3990 5660
rect 3914 5592 3936 5624
rect 3968 5592 3990 5624
rect 3914 5556 3990 5592
rect 3914 5524 3936 5556
rect 3968 5524 3990 5556
rect 3914 5488 3990 5524
rect 3914 5456 3936 5488
rect 3968 5456 3990 5488
rect 3914 5420 3990 5456
rect 3914 5388 3936 5420
rect 3968 5388 3990 5420
rect 3914 5352 3990 5388
rect 3914 5320 3936 5352
rect 3968 5320 3990 5352
rect 3914 5282 3990 5320
rect 4090 6644 4166 6682
rect 4090 6612 4112 6644
rect 4144 6612 4166 6644
rect 4090 6576 4166 6612
rect 4090 6544 4112 6576
rect 4144 6544 4166 6576
rect 4090 6508 4166 6544
rect 4090 6476 4112 6508
rect 4144 6476 4166 6508
rect 4090 6440 4166 6476
rect 4090 6408 4112 6440
rect 4144 6408 4166 6440
rect 4090 6372 4166 6408
rect 4090 6340 4112 6372
rect 4144 6340 4166 6372
rect 4090 6304 4166 6340
rect 4090 6272 4112 6304
rect 4144 6272 4166 6304
rect 4090 6236 4166 6272
rect 4090 6204 4112 6236
rect 4144 6204 4166 6236
rect 4090 6168 4166 6204
rect 4090 6136 4112 6168
rect 4144 6136 4166 6168
rect 4090 6100 4166 6136
rect 4090 6068 4112 6100
rect 4144 6068 4166 6100
rect 4090 6032 4166 6068
rect 4090 6000 4112 6032
rect 4144 6000 4166 6032
rect 4090 5964 4166 6000
rect 4090 5932 4112 5964
rect 4144 5932 4166 5964
rect 4090 5896 4166 5932
rect 4090 5864 4112 5896
rect 4144 5864 4166 5896
rect 4090 5828 4166 5864
rect 4090 5796 4112 5828
rect 4144 5796 4166 5828
rect 4090 5760 4166 5796
rect 4090 5728 4112 5760
rect 4144 5728 4166 5760
rect 4090 5692 4166 5728
rect 4090 5660 4112 5692
rect 4144 5660 4166 5692
rect 4090 5624 4166 5660
rect 4090 5592 4112 5624
rect 4144 5592 4166 5624
rect 4090 5556 4166 5592
rect 4090 5524 4112 5556
rect 4144 5524 4166 5556
rect 4090 5488 4166 5524
rect 4090 5456 4112 5488
rect 4144 5456 4166 5488
rect 4090 5420 4166 5456
rect 4090 5388 4112 5420
rect 4144 5388 4166 5420
rect 4090 5352 4166 5388
rect 4090 5320 4112 5352
rect 4144 5320 4166 5352
rect 4090 5282 4166 5320
rect 4266 6644 4342 6682
rect 4266 6612 4288 6644
rect 4320 6612 4342 6644
rect 4266 6576 4342 6612
rect 4266 6544 4288 6576
rect 4320 6544 4342 6576
rect 4266 6508 4342 6544
rect 4266 6476 4288 6508
rect 4320 6476 4342 6508
rect 4266 6440 4342 6476
rect 4266 6408 4288 6440
rect 4320 6408 4342 6440
rect 4266 6372 4342 6408
rect 4266 6340 4288 6372
rect 4320 6340 4342 6372
rect 4266 6304 4342 6340
rect 4266 6272 4288 6304
rect 4320 6272 4342 6304
rect 4266 6236 4342 6272
rect 4266 6204 4288 6236
rect 4320 6204 4342 6236
rect 4266 6168 4342 6204
rect 4266 6136 4288 6168
rect 4320 6136 4342 6168
rect 4266 6100 4342 6136
rect 4266 6068 4288 6100
rect 4320 6068 4342 6100
rect 4266 6032 4342 6068
rect 4266 6000 4288 6032
rect 4320 6000 4342 6032
rect 4266 5964 4342 6000
rect 4266 5932 4288 5964
rect 4320 5932 4342 5964
rect 4266 5896 4342 5932
rect 4266 5864 4288 5896
rect 4320 5864 4342 5896
rect 4266 5828 4342 5864
rect 4266 5796 4288 5828
rect 4320 5796 4342 5828
rect 4266 5760 4342 5796
rect 4266 5728 4288 5760
rect 4320 5728 4342 5760
rect 4266 5692 4342 5728
rect 4266 5660 4288 5692
rect 4320 5660 4342 5692
rect 4266 5624 4342 5660
rect 4266 5592 4288 5624
rect 4320 5592 4342 5624
rect 4266 5556 4342 5592
rect 4266 5524 4288 5556
rect 4320 5524 4342 5556
rect 4266 5488 4342 5524
rect 4266 5456 4288 5488
rect 4320 5456 4342 5488
rect 4266 5420 4342 5456
rect 4266 5388 4288 5420
rect 4320 5388 4342 5420
rect 4266 5352 4342 5388
rect 4266 5320 4288 5352
rect 4320 5320 4342 5352
rect 4266 5282 4342 5320
rect 4442 6644 4518 6682
rect 4442 6612 4464 6644
rect 4496 6612 4518 6644
rect 4442 6576 4518 6612
rect 4442 6544 4464 6576
rect 4496 6544 4518 6576
rect 4442 6508 4518 6544
rect 4442 6476 4464 6508
rect 4496 6476 4518 6508
rect 4442 6440 4518 6476
rect 4442 6408 4464 6440
rect 4496 6408 4518 6440
rect 4442 6372 4518 6408
rect 4442 6340 4464 6372
rect 4496 6340 4518 6372
rect 4442 6304 4518 6340
rect 4442 6272 4464 6304
rect 4496 6272 4518 6304
rect 4442 6236 4518 6272
rect 4442 6204 4464 6236
rect 4496 6204 4518 6236
rect 4442 6168 4518 6204
rect 4442 6136 4464 6168
rect 4496 6136 4518 6168
rect 4442 6100 4518 6136
rect 4442 6068 4464 6100
rect 4496 6068 4518 6100
rect 4442 6032 4518 6068
rect 4442 6000 4464 6032
rect 4496 6000 4518 6032
rect 4442 5964 4518 6000
rect 4442 5932 4464 5964
rect 4496 5932 4518 5964
rect 4442 5896 4518 5932
rect 4442 5864 4464 5896
rect 4496 5864 4518 5896
rect 4442 5828 4518 5864
rect 4442 5796 4464 5828
rect 4496 5796 4518 5828
rect 4442 5760 4518 5796
rect 4442 5728 4464 5760
rect 4496 5728 4518 5760
rect 4442 5692 4518 5728
rect 4442 5660 4464 5692
rect 4496 5660 4518 5692
rect 4442 5624 4518 5660
rect 4442 5592 4464 5624
rect 4496 5592 4518 5624
rect 4442 5556 4518 5592
rect 4442 5524 4464 5556
rect 4496 5524 4518 5556
rect 4442 5488 4518 5524
rect 4442 5456 4464 5488
rect 4496 5456 4518 5488
rect 4442 5420 4518 5456
rect 4442 5388 4464 5420
rect 4496 5388 4518 5420
rect 4442 5352 4518 5388
rect 4442 5320 4464 5352
rect 4496 5320 4518 5352
rect 4442 5282 4518 5320
rect 4618 6644 4694 6682
rect 4618 6612 4640 6644
rect 4672 6612 4694 6644
rect 4618 6576 4694 6612
rect 4618 6544 4640 6576
rect 4672 6544 4694 6576
rect 4618 6508 4694 6544
rect 4618 6476 4640 6508
rect 4672 6476 4694 6508
rect 4618 6440 4694 6476
rect 4618 6408 4640 6440
rect 4672 6408 4694 6440
rect 4618 6372 4694 6408
rect 4618 6340 4640 6372
rect 4672 6340 4694 6372
rect 4618 6304 4694 6340
rect 4618 6272 4640 6304
rect 4672 6272 4694 6304
rect 4618 6236 4694 6272
rect 4618 6204 4640 6236
rect 4672 6204 4694 6236
rect 4618 6168 4694 6204
rect 4618 6136 4640 6168
rect 4672 6136 4694 6168
rect 4618 6100 4694 6136
rect 4618 6068 4640 6100
rect 4672 6068 4694 6100
rect 4618 6032 4694 6068
rect 4618 6000 4640 6032
rect 4672 6000 4694 6032
rect 4618 5964 4694 6000
rect 4618 5932 4640 5964
rect 4672 5932 4694 5964
rect 4618 5896 4694 5932
rect 4618 5864 4640 5896
rect 4672 5864 4694 5896
rect 4618 5828 4694 5864
rect 4618 5796 4640 5828
rect 4672 5796 4694 5828
rect 4618 5760 4694 5796
rect 4618 5728 4640 5760
rect 4672 5728 4694 5760
rect 4618 5692 4694 5728
rect 4618 5660 4640 5692
rect 4672 5660 4694 5692
rect 4618 5624 4694 5660
rect 4618 5592 4640 5624
rect 4672 5592 4694 5624
rect 4618 5556 4694 5592
rect 4618 5524 4640 5556
rect 4672 5524 4694 5556
rect 4618 5488 4694 5524
rect 4618 5456 4640 5488
rect 4672 5456 4694 5488
rect 4618 5420 4694 5456
rect 4618 5388 4640 5420
rect 4672 5388 4694 5420
rect 4618 5352 4694 5388
rect 4618 5320 4640 5352
rect 4672 5320 4694 5352
rect 4618 5282 4694 5320
rect 4794 6644 4870 6682
rect 4794 6612 4816 6644
rect 4848 6612 4870 6644
rect 4794 6576 4870 6612
rect 4794 6544 4816 6576
rect 4848 6544 4870 6576
rect 4794 6508 4870 6544
rect 4794 6476 4816 6508
rect 4848 6476 4870 6508
rect 4794 6440 4870 6476
rect 4794 6408 4816 6440
rect 4848 6408 4870 6440
rect 4794 6372 4870 6408
rect 4794 6340 4816 6372
rect 4848 6340 4870 6372
rect 4794 6304 4870 6340
rect 4794 6272 4816 6304
rect 4848 6272 4870 6304
rect 4794 6236 4870 6272
rect 4794 6204 4816 6236
rect 4848 6204 4870 6236
rect 4794 6168 4870 6204
rect 4794 6136 4816 6168
rect 4848 6136 4870 6168
rect 4794 6100 4870 6136
rect 4794 6068 4816 6100
rect 4848 6068 4870 6100
rect 4794 6032 4870 6068
rect 4794 6000 4816 6032
rect 4848 6000 4870 6032
rect 4794 5964 4870 6000
rect 4794 5932 4816 5964
rect 4848 5932 4870 5964
rect 4794 5896 4870 5932
rect 4794 5864 4816 5896
rect 4848 5864 4870 5896
rect 4794 5828 4870 5864
rect 4794 5796 4816 5828
rect 4848 5796 4870 5828
rect 4794 5760 4870 5796
rect 4794 5728 4816 5760
rect 4848 5728 4870 5760
rect 4794 5692 4870 5728
rect 4794 5660 4816 5692
rect 4848 5660 4870 5692
rect 4794 5624 4870 5660
rect 4794 5592 4816 5624
rect 4848 5592 4870 5624
rect 4794 5556 4870 5592
rect 4794 5524 4816 5556
rect 4848 5524 4870 5556
rect 4794 5488 4870 5524
rect 4794 5456 4816 5488
rect 4848 5456 4870 5488
rect 4794 5420 4870 5456
rect 4794 5388 4816 5420
rect 4848 5388 4870 5420
rect 4794 5352 4870 5388
rect 4794 5320 4816 5352
rect 4848 5320 4870 5352
rect 4794 5282 4870 5320
rect 4970 6644 5046 6682
rect 4970 6612 4992 6644
rect 5024 6612 5046 6644
rect 4970 6576 5046 6612
rect 4970 6544 4992 6576
rect 5024 6544 5046 6576
rect 4970 6508 5046 6544
rect 4970 6476 4992 6508
rect 5024 6476 5046 6508
rect 4970 6440 5046 6476
rect 4970 6408 4992 6440
rect 5024 6408 5046 6440
rect 4970 6372 5046 6408
rect 4970 6340 4992 6372
rect 5024 6340 5046 6372
rect 4970 6304 5046 6340
rect 4970 6272 4992 6304
rect 5024 6272 5046 6304
rect 4970 6236 5046 6272
rect 4970 6204 4992 6236
rect 5024 6204 5046 6236
rect 4970 6168 5046 6204
rect 4970 6136 4992 6168
rect 5024 6136 5046 6168
rect 4970 6100 5046 6136
rect 4970 6068 4992 6100
rect 5024 6068 5046 6100
rect 4970 6032 5046 6068
rect 4970 6000 4992 6032
rect 5024 6000 5046 6032
rect 4970 5964 5046 6000
rect 4970 5932 4992 5964
rect 5024 5932 5046 5964
rect 4970 5896 5046 5932
rect 4970 5864 4992 5896
rect 5024 5864 5046 5896
rect 4970 5828 5046 5864
rect 4970 5796 4992 5828
rect 5024 5796 5046 5828
rect 4970 5760 5046 5796
rect 4970 5728 4992 5760
rect 5024 5728 5046 5760
rect 4970 5692 5046 5728
rect 4970 5660 4992 5692
rect 5024 5660 5046 5692
rect 4970 5624 5046 5660
rect 4970 5592 4992 5624
rect 5024 5592 5046 5624
rect 4970 5556 5046 5592
rect 4970 5524 4992 5556
rect 5024 5524 5046 5556
rect 4970 5488 5046 5524
rect 4970 5456 4992 5488
rect 5024 5456 5046 5488
rect 4970 5420 5046 5456
rect 4970 5388 4992 5420
rect 5024 5388 5046 5420
rect 4970 5352 5046 5388
rect 4970 5320 4992 5352
rect 5024 5320 5046 5352
rect 4970 5282 5046 5320
rect 5146 6644 5222 6682
rect 5146 6612 5168 6644
rect 5200 6612 5222 6644
rect 5146 6576 5222 6612
rect 5146 6544 5168 6576
rect 5200 6544 5222 6576
rect 5146 6508 5222 6544
rect 5146 6476 5168 6508
rect 5200 6476 5222 6508
rect 5146 6440 5222 6476
rect 5146 6408 5168 6440
rect 5200 6408 5222 6440
rect 5146 6372 5222 6408
rect 5146 6340 5168 6372
rect 5200 6340 5222 6372
rect 5146 6304 5222 6340
rect 5146 6272 5168 6304
rect 5200 6272 5222 6304
rect 5146 6236 5222 6272
rect 5146 6204 5168 6236
rect 5200 6204 5222 6236
rect 5146 6168 5222 6204
rect 5146 6136 5168 6168
rect 5200 6136 5222 6168
rect 5146 6100 5222 6136
rect 5146 6068 5168 6100
rect 5200 6068 5222 6100
rect 5146 6032 5222 6068
rect 5146 6000 5168 6032
rect 5200 6000 5222 6032
rect 5146 5964 5222 6000
rect 5146 5932 5168 5964
rect 5200 5932 5222 5964
rect 5146 5896 5222 5932
rect 5146 5864 5168 5896
rect 5200 5864 5222 5896
rect 5146 5828 5222 5864
rect 5146 5796 5168 5828
rect 5200 5796 5222 5828
rect 5146 5760 5222 5796
rect 5146 5728 5168 5760
rect 5200 5728 5222 5760
rect 5146 5692 5222 5728
rect 5146 5660 5168 5692
rect 5200 5660 5222 5692
rect 5146 5624 5222 5660
rect 5146 5592 5168 5624
rect 5200 5592 5222 5624
rect 5146 5556 5222 5592
rect 5146 5524 5168 5556
rect 5200 5524 5222 5556
rect 5146 5488 5222 5524
rect 5146 5456 5168 5488
rect 5200 5456 5222 5488
rect 5146 5420 5222 5456
rect 5146 5388 5168 5420
rect 5200 5388 5222 5420
rect 5146 5352 5222 5388
rect 5146 5320 5168 5352
rect 5200 5320 5222 5352
rect 5146 5282 5222 5320
rect 5322 6644 5398 6682
rect 5322 6612 5344 6644
rect 5376 6612 5398 6644
rect 5322 6576 5398 6612
rect 5322 6544 5344 6576
rect 5376 6544 5398 6576
rect 5322 6508 5398 6544
rect 5322 6476 5344 6508
rect 5376 6476 5398 6508
rect 5322 6440 5398 6476
rect 5322 6408 5344 6440
rect 5376 6408 5398 6440
rect 5322 6372 5398 6408
rect 5322 6340 5344 6372
rect 5376 6340 5398 6372
rect 5322 6304 5398 6340
rect 5322 6272 5344 6304
rect 5376 6272 5398 6304
rect 5322 6236 5398 6272
rect 5322 6204 5344 6236
rect 5376 6204 5398 6236
rect 5322 6168 5398 6204
rect 5322 6136 5344 6168
rect 5376 6136 5398 6168
rect 5322 6100 5398 6136
rect 5322 6068 5344 6100
rect 5376 6068 5398 6100
rect 5322 6032 5398 6068
rect 5322 6000 5344 6032
rect 5376 6000 5398 6032
rect 5322 5964 5398 6000
rect 5322 5932 5344 5964
rect 5376 5932 5398 5964
rect 5322 5896 5398 5932
rect 5322 5864 5344 5896
rect 5376 5864 5398 5896
rect 5322 5828 5398 5864
rect 5322 5796 5344 5828
rect 5376 5796 5398 5828
rect 5322 5760 5398 5796
rect 5322 5728 5344 5760
rect 5376 5728 5398 5760
rect 5322 5692 5398 5728
rect 5322 5660 5344 5692
rect 5376 5660 5398 5692
rect 5322 5624 5398 5660
rect 5322 5592 5344 5624
rect 5376 5592 5398 5624
rect 5322 5556 5398 5592
rect 5322 5524 5344 5556
rect 5376 5524 5398 5556
rect 5322 5488 5398 5524
rect 5322 5456 5344 5488
rect 5376 5456 5398 5488
rect 5322 5420 5398 5456
rect 5322 5388 5344 5420
rect 5376 5388 5398 5420
rect 5322 5352 5398 5388
rect 5322 5320 5344 5352
rect 5376 5320 5398 5352
rect 5322 5282 5398 5320
rect 5498 6644 5574 6682
rect 5498 6612 5520 6644
rect 5552 6612 5574 6644
rect 5498 6576 5574 6612
rect 5498 6544 5520 6576
rect 5552 6544 5574 6576
rect 5498 6508 5574 6544
rect 5498 6476 5520 6508
rect 5552 6476 5574 6508
rect 5498 6440 5574 6476
rect 5498 6408 5520 6440
rect 5552 6408 5574 6440
rect 5498 6372 5574 6408
rect 5498 6340 5520 6372
rect 5552 6340 5574 6372
rect 5498 6304 5574 6340
rect 5498 6272 5520 6304
rect 5552 6272 5574 6304
rect 5498 6236 5574 6272
rect 5498 6204 5520 6236
rect 5552 6204 5574 6236
rect 5498 6168 5574 6204
rect 5498 6136 5520 6168
rect 5552 6136 5574 6168
rect 5498 6100 5574 6136
rect 5498 6068 5520 6100
rect 5552 6068 5574 6100
rect 5498 6032 5574 6068
rect 5498 6000 5520 6032
rect 5552 6000 5574 6032
rect 5498 5964 5574 6000
rect 5498 5932 5520 5964
rect 5552 5932 5574 5964
rect 5498 5896 5574 5932
rect 5498 5864 5520 5896
rect 5552 5864 5574 5896
rect 5498 5828 5574 5864
rect 5498 5796 5520 5828
rect 5552 5796 5574 5828
rect 5498 5760 5574 5796
rect 5498 5728 5520 5760
rect 5552 5728 5574 5760
rect 5498 5692 5574 5728
rect 5498 5660 5520 5692
rect 5552 5660 5574 5692
rect 5498 5624 5574 5660
rect 5498 5592 5520 5624
rect 5552 5592 5574 5624
rect 5498 5556 5574 5592
rect 5498 5524 5520 5556
rect 5552 5524 5574 5556
rect 5498 5488 5574 5524
rect 5498 5456 5520 5488
rect 5552 5456 5574 5488
rect 5498 5420 5574 5456
rect 5498 5388 5520 5420
rect 5552 5388 5574 5420
rect 5498 5352 5574 5388
rect 5498 5320 5520 5352
rect 5552 5320 5574 5352
rect 5498 5282 5574 5320
rect 5674 6644 5750 6682
rect 5674 6612 5696 6644
rect 5728 6612 5750 6644
rect 5674 6576 5750 6612
rect 5674 6544 5696 6576
rect 5728 6544 5750 6576
rect 5674 6508 5750 6544
rect 5674 6476 5696 6508
rect 5728 6476 5750 6508
rect 5674 6440 5750 6476
rect 5674 6408 5696 6440
rect 5728 6408 5750 6440
rect 5674 6372 5750 6408
rect 5674 6340 5696 6372
rect 5728 6340 5750 6372
rect 5674 6304 5750 6340
rect 5674 6272 5696 6304
rect 5728 6272 5750 6304
rect 5674 6236 5750 6272
rect 5674 6204 5696 6236
rect 5728 6204 5750 6236
rect 5674 6168 5750 6204
rect 5674 6136 5696 6168
rect 5728 6136 5750 6168
rect 5674 6100 5750 6136
rect 5674 6068 5696 6100
rect 5728 6068 5750 6100
rect 5674 6032 5750 6068
rect 5674 6000 5696 6032
rect 5728 6000 5750 6032
rect 5674 5964 5750 6000
rect 5674 5932 5696 5964
rect 5728 5932 5750 5964
rect 5674 5896 5750 5932
rect 5674 5864 5696 5896
rect 5728 5864 5750 5896
rect 5674 5828 5750 5864
rect 5674 5796 5696 5828
rect 5728 5796 5750 5828
rect 5674 5760 5750 5796
rect 5674 5728 5696 5760
rect 5728 5728 5750 5760
rect 5674 5692 5750 5728
rect 5674 5660 5696 5692
rect 5728 5660 5750 5692
rect 5674 5624 5750 5660
rect 5674 5592 5696 5624
rect 5728 5592 5750 5624
rect 5674 5556 5750 5592
rect 5674 5524 5696 5556
rect 5728 5524 5750 5556
rect 5674 5488 5750 5524
rect 5674 5456 5696 5488
rect 5728 5456 5750 5488
rect 5674 5420 5750 5456
rect 5674 5388 5696 5420
rect 5728 5388 5750 5420
rect 5674 5352 5750 5388
rect 5674 5320 5696 5352
rect 5728 5320 5750 5352
rect 5674 5282 5750 5320
rect 5850 6644 5926 6682
rect 5850 6612 5872 6644
rect 5904 6612 5926 6644
rect 5850 6576 5926 6612
rect 5850 6544 5872 6576
rect 5904 6544 5926 6576
rect 5850 6508 5926 6544
rect 5850 6476 5872 6508
rect 5904 6476 5926 6508
rect 5850 6440 5926 6476
rect 5850 6408 5872 6440
rect 5904 6408 5926 6440
rect 5850 6372 5926 6408
rect 5850 6340 5872 6372
rect 5904 6340 5926 6372
rect 5850 6304 5926 6340
rect 5850 6272 5872 6304
rect 5904 6272 5926 6304
rect 5850 6236 5926 6272
rect 5850 6204 5872 6236
rect 5904 6204 5926 6236
rect 5850 6168 5926 6204
rect 5850 6136 5872 6168
rect 5904 6136 5926 6168
rect 5850 6100 5926 6136
rect 5850 6068 5872 6100
rect 5904 6068 5926 6100
rect 5850 6032 5926 6068
rect 5850 6000 5872 6032
rect 5904 6000 5926 6032
rect 5850 5964 5926 6000
rect 5850 5932 5872 5964
rect 5904 5932 5926 5964
rect 5850 5896 5926 5932
rect 5850 5864 5872 5896
rect 5904 5864 5926 5896
rect 5850 5828 5926 5864
rect 5850 5796 5872 5828
rect 5904 5796 5926 5828
rect 5850 5760 5926 5796
rect 5850 5728 5872 5760
rect 5904 5728 5926 5760
rect 5850 5692 5926 5728
rect 5850 5660 5872 5692
rect 5904 5660 5926 5692
rect 5850 5624 5926 5660
rect 5850 5592 5872 5624
rect 5904 5592 5926 5624
rect 5850 5556 5926 5592
rect 5850 5524 5872 5556
rect 5904 5524 5926 5556
rect 5850 5488 5926 5524
rect 5850 5456 5872 5488
rect 5904 5456 5926 5488
rect 5850 5420 5926 5456
rect 5850 5388 5872 5420
rect 5904 5388 5926 5420
rect 5850 5352 5926 5388
rect 5850 5320 5872 5352
rect 5904 5320 5926 5352
rect 5850 5282 5926 5320
rect 6026 6644 6102 6682
rect 6026 6612 6048 6644
rect 6080 6612 6102 6644
rect 6026 6576 6102 6612
rect 6026 6544 6048 6576
rect 6080 6544 6102 6576
rect 6026 6508 6102 6544
rect 6026 6476 6048 6508
rect 6080 6476 6102 6508
rect 6026 6440 6102 6476
rect 6026 6408 6048 6440
rect 6080 6408 6102 6440
rect 6026 6372 6102 6408
rect 6026 6340 6048 6372
rect 6080 6340 6102 6372
rect 6026 6304 6102 6340
rect 6026 6272 6048 6304
rect 6080 6272 6102 6304
rect 6026 6236 6102 6272
rect 6026 6204 6048 6236
rect 6080 6204 6102 6236
rect 6026 6168 6102 6204
rect 6026 6136 6048 6168
rect 6080 6136 6102 6168
rect 6026 6100 6102 6136
rect 6026 6068 6048 6100
rect 6080 6068 6102 6100
rect 6026 6032 6102 6068
rect 6026 6000 6048 6032
rect 6080 6000 6102 6032
rect 6026 5964 6102 6000
rect 6026 5932 6048 5964
rect 6080 5932 6102 5964
rect 6026 5896 6102 5932
rect 6026 5864 6048 5896
rect 6080 5864 6102 5896
rect 6026 5828 6102 5864
rect 6026 5796 6048 5828
rect 6080 5796 6102 5828
rect 6026 5760 6102 5796
rect 6026 5728 6048 5760
rect 6080 5728 6102 5760
rect 6026 5692 6102 5728
rect 6026 5660 6048 5692
rect 6080 5660 6102 5692
rect 6026 5624 6102 5660
rect 6026 5592 6048 5624
rect 6080 5592 6102 5624
rect 6026 5556 6102 5592
rect 6026 5524 6048 5556
rect 6080 5524 6102 5556
rect 6026 5488 6102 5524
rect 6026 5456 6048 5488
rect 6080 5456 6102 5488
rect 6026 5420 6102 5456
rect 6026 5388 6048 5420
rect 6080 5388 6102 5420
rect 6026 5352 6102 5388
rect 6026 5320 6048 5352
rect 6080 5320 6102 5352
rect 6026 5282 6102 5320
rect 6202 6644 6278 6682
rect 6202 6612 6224 6644
rect 6256 6612 6278 6644
rect 6202 6576 6278 6612
rect 6202 6544 6224 6576
rect 6256 6544 6278 6576
rect 6202 6508 6278 6544
rect 6202 6476 6224 6508
rect 6256 6476 6278 6508
rect 6202 6440 6278 6476
rect 6202 6408 6224 6440
rect 6256 6408 6278 6440
rect 6202 6372 6278 6408
rect 6202 6340 6224 6372
rect 6256 6340 6278 6372
rect 6202 6304 6278 6340
rect 6202 6272 6224 6304
rect 6256 6272 6278 6304
rect 6202 6236 6278 6272
rect 6202 6204 6224 6236
rect 6256 6204 6278 6236
rect 6202 6168 6278 6204
rect 6202 6136 6224 6168
rect 6256 6136 6278 6168
rect 6202 6100 6278 6136
rect 6202 6068 6224 6100
rect 6256 6068 6278 6100
rect 6202 6032 6278 6068
rect 6202 6000 6224 6032
rect 6256 6000 6278 6032
rect 6202 5964 6278 6000
rect 6202 5932 6224 5964
rect 6256 5932 6278 5964
rect 6202 5896 6278 5932
rect 6202 5864 6224 5896
rect 6256 5864 6278 5896
rect 6202 5828 6278 5864
rect 6202 5796 6224 5828
rect 6256 5796 6278 5828
rect 6202 5760 6278 5796
rect 6202 5728 6224 5760
rect 6256 5728 6278 5760
rect 6202 5692 6278 5728
rect 6202 5660 6224 5692
rect 6256 5660 6278 5692
rect 6202 5624 6278 5660
rect 6202 5592 6224 5624
rect 6256 5592 6278 5624
rect 6202 5556 6278 5592
rect 6202 5524 6224 5556
rect 6256 5524 6278 5556
rect 6202 5488 6278 5524
rect 6202 5456 6224 5488
rect 6256 5456 6278 5488
rect 6202 5420 6278 5456
rect 6202 5388 6224 5420
rect 6256 5388 6278 5420
rect 6202 5352 6278 5388
rect 6202 5320 6224 5352
rect 6256 5320 6278 5352
rect 6202 5282 6278 5320
rect 6378 6644 6454 6682
rect 6378 6612 6400 6644
rect 6432 6612 6454 6644
rect 6378 6576 6454 6612
rect 6378 6544 6400 6576
rect 6432 6544 6454 6576
rect 6378 6508 6454 6544
rect 6378 6476 6400 6508
rect 6432 6476 6454 6508
rect 6378 6440 6454 6476
rect 6378 6408 6400 6440
rect 6432 6408 6454 6440
rect 6378 6372 6454 6408
rect 6378 6340 6400 6372
rect 6432 6340 6454 6372
rect 6378 6304 6454 6340
rect 6378 6272 6400 6304
rect 6432 6272 6454 6304
rect 6378 6236 6454 6272
rect 6378 6204 6400 6236
rect 6432 6204 6454 6236
rect 6378 6168 6454 6204
rect 6378 6136 6400 6168
rect 6432 6136 6454 6168
rect 6378 6100 6454 6136
rect 6378 6068 6400 6100
rect 6432 6068 6454 6100
rect 6378 6032 6454 6068
rect 6378 6000 6400 6032
rect 6432 6000 6454 6032
rect 6378 5964 6454 6000
rect 6378 5932 6400 5964
rect 6432 5932 6454 5964
rect 6378 5896 6454 5932
rect 6378 5864 6400 5896
rect 6432 5864 6454 5896
rect 6378 5828 6454 5864
rect 6378 5796 6400 5828
rect 6432 5796 6454 5828
rect 6378 5760 6454 5796
rect 6378 5728 6400 5760
rect 6432 5728 6454 5760
rect 6378 5692 6454 5728
rect 6378 5660 6400 5692
rect 6432 5660 6454 5692
rect 6378 5624 6454 5660
rect 6378 5592 6400 5624
rect 6432 5592 6454 5624
rect 6378 5556 6454 5592
rect 6378 5524 6400 5556
rect 6432 5524 6454 5556
rect 6378 5488 6454 5524
rect 6378 5456 6400 5488
rect 6432 5456 6454 5488
rect 6378 5420 6454 5456
rect 6378 5388 6400 5420
rect 6432 5388 6454 5420
rect 6378 5352 6454 5388
rect 6378 5320 6400 5352
rect 6432 5320 6454 5352
rect 6378 5282 6454 5320
rect 6554 6644 6630 6682
rect 6554 6612 6576 6644
rect 6608 6612 6630 6644
rect 6554 6576 6630 6612
rect 6554 6544 6576 6576
rect 6608 6544 6630 6576
rect 6554 6508 6630 6544
rect 6554 6476 6576 6508
rect 6608 6476 6630 6508
rect 6554 6440 6630 6476
rect 6554 6408 6576 6440
rect 6608 6408 6630 6440
rect 6554 6372 6630 6408
rect 6554 6340 6576 6372
rect 6608 6340 6630 6372
rect 6554 6304 6630 6340
rect 6554 6272 6576 6304
rect 6608 6272 6630 6304
rect 6554 6236 6630 6272
rect 6554 6204 6576 6236
rect 6608 6204 6630 6236
rect 6554 6168 6630 6204
rect 6554 6136 6576 6168
rect 6608 6136 6630 6168
rect 6554 6100 6630 6136
rect 6554 6068 6576 6100
rect 6608 6068 6630 6100
rect 6554 6032 6630 6068
rect 6554 6000 6576 6032
rect 6608 6000 6630 6032
rect 6554 5964 6630 6000
rect 6554 5932 6576 5964
rect 6608 5932 6630 5964
rect 6554 5896 6630 5932
rect 6554 5864 6576 5896
rect 6608 5864 6630 5896
rect 6554 5828 6630 5864
rect 6554 5796 6576 5828
rect 6608 5796 6630 5828
rect 6554 5760 6630 5796
rect 6554 5728 6576 5760
rect 6608 5728 6630 5760
rect 6554 5692 6630 5728
rect 6554 5660 6576 5692
rect 6608 5660 6630 5692
rect 6554 5624 6630 5660
rect 6554 5592 6576 5624
rect 6608 5592 6630 5624
rect 6554 5556 6630 5592
rect 6554 5524 6576 5556
rect 6608 5524 6630 5556
rect 6554 5488 6630 5524
rect 6554 5456 6576 5488
rect 6608 5456 6630 5488
rect 6554 5420 6630 5456
rect 6554 5388 6576 5420
rect 6608 5388 6630 5420
rect 6554 5352 6630 5388
rect 6554 5320 6576 5352
rect 6608 5320 6630 5352
rect 6554 5282 6630 5320
rect 6730 6644 6806 6682
rect 6730 6612 6752 6644
rect 6784 6612 6806 6644
rect 6730 6576 6806 6612
rect 6730 6544 6752 6576
rect 6784 6544 6806 6576
rect 6730 6508 6806 6544
rect 6730 6476 6752 6508
rect 6784 6476 6806 6508
rect 6730 6440 6806 6476
rect 6730 6408 6752 6440
rect 6784 6408 6806 6440
rect 6730 6372 6806 6408
rect 6730 6340 6752 6372
rect 6784 6340 6806 6372
rect 6730 6304 6806 6340
rect 6730 6272 6752 6304
rect 6784 6272 6806 6304
rect 6730 6236 6806 6272
rect 6730 6204 6752 6236
rect 6784 6204 6806 6236
rect 6730 6168 6806 6204
rect 6730 6136 6752 6168
rect 6784 6136 6806 6168
rect 6730 6100 6806 6136
rect 6730 6068 6752 6100
rect 6784 6068 6806 6100
rect 6730 6032 6806 6068
rect 6730 6000 6752 6032
rect 6784 6000 6806 6032
rect 6730 5964 6806 6000
rect 6730 5932 6752 5964
rect 6784 5932 6806 5964
rect 6730 5896 6806 5932
rect 6730 5864 6752 5896
rect 6784 5864 6806 5896
rect 6730 5828 6806 5864
rect 6730 5796 6752 5828
rect 6784 5796 6806 5828
rect 6730 5760 6806 5796
rect 6730 5728 6752 5760
rect 6784 5728 6806 5760
rect 6730 5692 6806 5728
rect 6730 5660 6752 5692
rect 6784 5660 6806 5692
rect 6730 5624 6806 5660
rect 6730 5592 6752 5624
rect 6784 5592 6806 5624
rect 6730 5556 6806 5592
rect 6730 5524 6752 5556
rect 6784 5524 6806 5556
rect 6730 5488 6806 5524
rect 6730 5456 6752 5488
rect 6784 5456 6806 5488
rect 6730 5420 6806 5456
rect 6730 5388 6752 5420
rect 6784 5388 6806 5420
rect 6730 5352 6806 5388
rect 6730 5320 6752 5352
rect 6784 5320 6806 5352
rect 6730 5282 6806 5320
rect 6906 6644 6982 6682
rect 6906 6612 6928 6644
rect 6960 6612 6982 6644
rect 6906 6576 6982 6612
rect 6906 6544 6928 6576
rect 6960 6544 6982 6576
rect 6906 6508 6982 6544
rect 6906 6476 6928 6508
rect 6960 6476 6982 6508
rect 6906 6440 6982 6476
rect 6906 6408 6928 6440
rect 6960 6408 6982 6440
rect 6906 6372 6982 6408
rect 6906 6340 6928 6372
rect 6960 6340 6982 6372
rect 6906 6304 6982 6340
rect 6906 6272 6928 6304
rect 6960 6272 6982 6304
rect 6906 6236 6982 6272
rect 6906 6204 6928 6236
rect 6960 6204 6982 6236
rect 6906 6168 6982 6204
rect 6906 6136 6928 6168
rect 6960 6136 6982 6168
rect 6906 6100 6982 6136
rect 6906 6068 6928 6100
rect 6960 6068 6982 6100
rect 6906 6032 6982 6068
rect 6906 6000 6928 6032
rect 6960 6000 6982 6032
rect 6906 5964 6982 6000
rect 6906 5932 6928 5964
rect 6960 5932 6982 5964
rect 6906 5896 6982 5932
rect 6906 5864 6928 5896
rect 6960 5864 6982 5896
rect 6906 5828 6982 5864
rect 6906 5796 6928 5828
rect 6960 5796 6982 5828
rect 6906 5760 6982 5796
rect 6906 5728 6928 5760
rect 6960 5728 6982 5760
rect 6906 5692 6982 5728
rect 6906 5660 6928 5692
rect 6960 5660 6982 5692
rect 6906 5624 6982 5660
rect 6906 5592 6928 5624
rect 6960 5592 6982 5624
rect 6906 5556 6982 5592
rect 6906 5524 6928 5556
rect 6960 5524 6982 5556
rect 6906 5488 6982 5524
rect 6906 5456 6928 5488
rect 6960 5456 6982 5488
rect 6906 5420 6982 5456
rect 6906 5388 6928 5420
rect 6960 5388 6982 5420
rect 6906 5352 6982 5388
rect 6906 5320 6928 5352
rect 6960 5320 6982 5352
rect 6906 5282 6982 5320
rect 7082 6644 7158 6682
rect 7082 6612 7104 6644
rect 7136 6612 7158 6644
rect 7082 6576 7158 6612
rect 7082 6544 7104 6576
rect 7136 6544 7158 6576
rect 7082 6508 7158 6544
rect 7082 6476 7104 6508
rect 7136 6476 7158 6508
rect 7082 6440 7158 6476
rect 7082 6408 7104 6440
rect 7136 6408 7158 6440
rect 7082 6372 7158 6408
rect 7082 6340 7104 6372
rect 7136 6340 7158 6372
rect 7082 6304 7158 6340
rect 7082 6272 7104 6304
rect 7136 6272 7158 6304
rect 7082 6236 7158 6272
rect 7082 6204 7104 6236
rect 7136 6204 7158 6236
rect 7082 6168 7158 6204
rect 7082 6136 7104 6168
rect 7136 6136 7158 6168
rect 7082 6100 7158 6136
rect 7082 6068 7104 6100
rect 7136 6068 7158 6100
rect 7082 6032 7158 6068
rect 7082 6000 7104 6032
rect 7136 6000 7158 6032
rect 7082 5964 7158 6000
rect 7082 5932 7104 5964
rect 7136 5932 7158 5964
rect 7082 5896 7158 5932
rect 7082 5864 7104 5896
rect 7136 5864 7158 5896
rect 7082 5828 7158 5864
rect 7082 5796 7104 5828
rect 7136 5796 7158 5828
rect 7082 5760 7158 5796
rect 7082 5728 7104 5760
rect 7136 5728 7158 5760
rect 7082 5692 7158 5728
rect 7082 5660 7104 5692
rect 7136 5660 7158 5692
rect 7082 5624 7158 5660
rect 7082 5592 7104 5624
rect 7136 5592 7158 5624
rect 7082 5556 7158 5592
rect 7082 5524 7104 5556
rect 7136 5524 7158 5556
rect 7082 5488 7158 5524
rect 7082 5456 7104 5488
rect 7136 5456 7158 5488
rect 7082 5420 7158 5456
rect 7082 5388 7104 5420
rect 7136 5388 7158 5420
rect 7082 5352 7158 5388
rect 7082 5320 7104 5352
rect 7136 5320 7158 5352
rect 7082 5282 7158 5320
rect 7258 6644 7334 6682
rect 7258 6612 7280 6644
rect 7312 6612 7334 6644
rect 7258 6576 7334 6612
rect 7258 6544 7280 6576
rect 7312 6544 7334 6576
rect 7258 6508 7334 6544
rect 7258 6476 7280 6508
rect 7312 6476 7334 6508
rect 7258 6440 7334 6476
rect 7258 6408 7280 6440
rect 7312 6408 7334 6440
rect 7258 6372 7334 6408
rect 7258 6340 7280 6372
rect 7312 6340 7334 6372
rect 7258 6304 7334 6340
rect 7258 6272 7280 6304
rect 7312 6272 7334 6304
rect 7258 6236 7334 6272
rect 7258 6204 7280 6236
rect 7312 6204 7334 6236
rect 7258 6168 7334 6204
rect 7258 6136 7280 6168
rect 7312 6136 7334 6168
rect 7258 6100 7334 6136
rect 7258 6068 7280 6100
rect 7312 6068 7334 6100
rect 7258 6032 7334 6068
rect 7258 6000 7280 6032
rect 7312 6000 7334 6032
rect 7258 5964 7334 6000
rect 7258 5932 7280 5964
rect 7312 5932 7334 5964
rect 7258 5896 7334 5932
rect 7258 5864 7280 5896
rect 7312 5864 7334 5896
rect 7258 5828 7334 5864
rect 7258 5796 7280 5828
rect 7312 5796 7334 5828
rect 7258 5760 7334 5796
rect 7258 5728 7280 5760
rect 7312 5728 7334 5760
rect 7258 5692 7334 5728
rect 7258 5660 7280 5692
rect 7312 5660 7334 5692
rect 7258 5624 7334 5660
rect 7258 5592 7280 5624
rect 7312 5592 7334 5624
rect 7258 5556 7334 5592
rect 7258 5524 7280 5556
rect 7312 5524 7334 5556
rect 7258 5488 7334 5524
rect 7258 5456 7280 5488
rect 7312 5456 7334 5488
rect 7258 5420 7334 5456
rect 7258 5388 7280 5420
rect 7312 5388 7334 5420
rect 7258 5352 7334 5388
rect 7258 5320 7280 5352
rect 7312 5320 7334 5352
rect 7258 5282 7334 5320
rect 7434 6644 7510 6682
rect 7434 6612 7456 6644
rect 7488 6612 7510 6644
rect 7434 6576 7510 6612
rect 7434 6544 7456 6576
rect 7488 6544 7510 6576
rect 7434 6508 7510 6544
rect 7434 6476 7456 6508
rect 7488 6476 7510 6508
rect 7434 6440 7510 6476
rect 7434 6408 7456 6440
rect 7488 6408 7510 6440
rect 7434 6372 7510 6408
rect 7434 6340 7456 6372
rect 7488 6340 7510 6372
rect 7434 6304 7510 6340
rect 7434 6272 7456 6304
rect 7488 6272 7510 6304
rect 7434 6236 7510 6272
rect 7434 6204 7456 6236
rect 7488 6204 7510 6236
rect 7434 6168 7510 6204
rect 7434 6136 7456 6168
rect 7488 6136 7510 6168
rect 7434 6100 7510 6136
rect 7434 6068 7456 6100
rect 7488 6068 7510 6100
rect 7434 6032 7510 6068
rect 7434 6000 7456 6032
rect 7488 6000 7510 6032
rect 7434 5964 7510 6000
rect 7434 5932 7456 5964
rect 7488 5932 7510 5964
rect 7434 5896 7510 5932
rect 7434 5864 7456 5896
rect 7488 5864 7510 5896
rect 7434 5828 7510 5864
rect 7434 5796 7456 5828
rect 7488 5796 7510 5828
rect 7434 5760 7510 5796
rect 7434 5728 7456 5760
rect 7488 5728 7510 5760
rect 7434 5692 7510 5728
rect 7434 5660 7456 5692
rect 7488 5660 7510 5692
rect 7434 5624 7510 5660
rect 7434 5592 7456 5624
rect 7488 5592 7510 5624
rect 7434 5556 7510 5592
rect 7434 5524 7456 5556
rect 7488 5524 7510 5556
rect 7434 5488 7510 5524
rect 7434 5456 7456 5488
rect 7488 5456 7510 5488
rect 7434 5420 7510 5456
rect 7434 5388 7456 5420
rect 7488 5388 7510 5420
rect 7434 5352 7510 5388
rect 7434 5320 7456 5352
rect 7488 5320 7510 5352
rect 7434 5282 7510 5320
rect 7610 6644 7686 6682
rect 7610 6612 7632 6644
rect 7664 6612 7686 6644
rect 7610 6576 7686 6612
rect 7610 6544 7632 6576
rect 7664 6544 7686 6576
rect 7610 6508 7686 6544
rect 7610 6476 7632 6508
rect 7664 6476 7686 6508
rect 7610 6440 7686 6476
rect 7610 6408 7632 6440
rect 7664 6408 7686 6440
rect 7610 6372 7686 6408
rect 7610 6340 7632 6372
rect 7664 6340 7686 6372
rect 7610 6304 7686 6340
rect 7610 6272 7632 6304
rect 7664 6272 7686 6304
rect 7610 6236 7686 6272
rect 7610 6204 7632 6236
rect 7664 6204 7686 6236
rect 7610 6168 7686 6204
rect 7610 6136 7632 6168
rect 7664 6136 7686 6168
rect 7610 6100 7686 6136
rect 7610 6068 7632 6100
rect 7664 6068 7686 6100
rect 7610 6032 7686 6068
rect 7610 6000 7632 6032
rect 7664 6000 7686 6032
rect 7610 5964 7686 6000
rect 7610 5932 7632 5964
rect 7664 5932 7686 5964
rect 7610 5896 7686 5932
rect 7610 5864 7632 5896
rect 7664 5864 7686 5896
rect 7610 5828 7686 5864
rect 7610 5796 7632 5828
rect 7664 5796 7686 5828
rect 7610 5760 7686 5796
rect 7610 5728 7632 5760
rect 7664 5728 7686 5760
rect 7610 5692 7686 5728
rect 7610 5660 7632 5692
rect 7664 5660 7686 5692
rect 7610 5624 7686 5660
rect 7610 5592 7632 5624
rect 7664 5592 7686 5624
rect 7610 5556 7686 5592
rect 7610 5524 7632 5556
rect 7664 5524 7686 5556
rect 7610 5488 7686 5524
rect 7610 5456 7632 5488
rect 7664 5456 7686 5488
rect 7610 5420 7686 5456
rect 7610 5388 7632 5420
rect 7664 5388 7686 5420
rect 7610 5352 7686 5388
rect 7610 5320 7632 5352
rect 7664 5320 7686 5352
rect 7610 5282 7686 5320
rect 7786 6644 7862 6682
rect 7786 6612 7808 6644
rect 7840 6612 7862 6644
rect 7786 6576 7862 6612
rect 7786 6544 7808 6576
rect 7840 6544 7862 6576
rect 7786 6508 7862 6544
rect 7786 6476 7808 6508
rect 7840 6476 7862 6508
rect 7786 6440 7862 6476
rect 7786 6408 7808 6440
rect 7840 6408 7862 6440
rect 7786 6372 7862 6408
rect 7786 6340 7808 6372
rect 7840 6340 7862 6372
rect 7786 6304 7862 6340
rect 7786 6272 7808 6304
rect 7840 6272 7862 6304
rect 7786 6236 7862 6272
rect 7786 6204 7808 6236
rect 7840 6204 7862 6236
rect 7786 6168 7862 6204
rect 7786 6136 7808 6168
rect 7840 6136 7862 6168
rect 7786 6100 7862 6136
rect 7786 6068 7808 6100
rect 7840 6068 7862 6100
rect 7786 6032 7862 6068
rect 7786 6000 7808 6032
rect 7840 6000 7862 6032
rect 7786 5964 7862 6000
rect 7786 5932 7808 5964
rect 7840 5932 7862 5964
rect 7786 5896 7862 5932
rect 7786 5864 7808 5896
rect 7840 5864 7862 5896
rect 7786 5828 7862 5864
rect 7786 5796 7808 5828
rect 7840 5796 7862 5828
rect 7786 5760 7862 5796
rect 7786 5728 7808 5760
rect 7840 5728 7862 5760
rect 7786 5692 7862 5728
rect 7786 5660 7808 5692
rect 7840 5660 7862 5692
rect 7786 5624 7862 5660
rect 7786 5592 7808 5624
rect 7840 5592 7862 5624
rect 7786 5556 7862 5592
rect 7786 5524 7808 5556
rect 7840 5524 7862 5556
rect 7786 5488 7862 5524
rect 7786 5456 7808 5488
rect 7840 5456 7862 5488
rect 7786 5420 7862 5456
rect 7786 5388 7808 5420
rect 7840 5388 7862 5420
rect 7786 5352 7862 5388
rect 7786 5320 7808 5352
rect 7840 5320 7862 5352
rect 7786 5282 7862 5320
rect 7962 6644 8038 6682
rect 7962 6612 7984 6644
rect 8016 6612 8038 6644
rect 7962 6576 8038 6612
rect 7962 6544 7984 6576
rect 8016 6544 8038 6576
rect 7962 6508 8038 6544
rect 7962 6476 7984 6508
rect 8016 6476 8038 6508
rect 7962 6440 8038 6476
rect 7962 6408 7984 6440
rect 8016 6408 8038 6440
rect 7962 6372 8038 6408
rect 7962 6340 7984 6372
rect 8016 6340 8038 6372
rect 7962 6304 8038 6340
rect 7962 6272 7984 6304
rect 8016 6272 8038 6304
rect 7962 6236 8038 6272
rect 7962 6204 7984 6236
rect 8016 6204 8038 6236
rect 7962 6168 8038 6204
rect 7962 6136 7984 6168
rect 8016 6136 8038 6168
rect 7962 6100 8038 6136
rect 7962 6068 7984 6100
rect 8016 6068 8038 6100
rect 7962 6032 8038 6068
rect 7962 6000 7984 6032
rect 8016 6000 8038 6032
rect 7962 5964 8038 6000
rect 7962 5932 7984 5964
rect 8016 5932 8038 5964
rect 7962 5896 8038 5932
rect 7962 5864 7984 5896
rect 8016 5864 8038 5896
rect 7962 5828 8038 5864
rect 7962 5796 7984 5828
rect 8016 5796 8038 5828
rect 7962 5760 8038 5796
rect 7962 5728 7984 5760
rect 8016 5728 8038 5760
rect 7962 5692 8038 5728
rect 7962 5660 7984 5692
rect 8016 5660 8038 5692
rect 7962 5624 8038 5660
rect 7962 5592 7984 5624
rect 8016 5592 8038 5624
rect 7962 5556 8038 5592
rect 7962 5524 7984 5556
rect 8016 5524 8038 5556
rect 7962 5488 8038 5524
rect 7962 5456 7984 5488
rect 8016 5456 8038 5488
rect 7962 5420 8038 5456
rect 7962 5388 7984 5420
rect 8016 5388 8038 5420
rect 7962 5352 8038 5388
rect 7962 5320 7984 5352
rect 8016 5320 8038 5352
rect 7962 5282 8038 5320
rect 8138 6644 8214 6682
rect 8138 6612 8160 6644
rect 8192 6612 8214 6644
rect 8138 6576 8214 6612
rect 8138 6544 8160 6576
rect 8192 6544 8214 6576
rect 8138 6508 8214 6544
rect 8138 6476 8160 6508
rect 8192 6476 8214 6508
rect 8138 6440 8214 6476
rect 8138 6408 8160 6440
rect 8192 6408 8214 6440
rect 8138 6372 8214 6408
rect 8138 6340 8160 6372
rect 8192 6340 8214 6372
rect 8138 6304 8214 6340
rect 8138 6272 8160 6304
rect 8192 6272 8214 6304
rect 8138 6236 8214 6272
rect 8138 6204 8160 6236
rect 8192 6204 8214 6236
rect 8138 6168 8214 6204
rect 8138 6136 8160 6168
rect 8192 6136 8214 6168
rect 8138 6100 8214 6136
rect 8138 6068 8160 6100
rect 8192 6068 8214 6100
rect 8138 6032 8214 6068
rect 8138 6000 8160 6032
rect 8192 6000 8214 6032
rect 8138 5964 8214 6000
rect 8138 5932 8160 5964
rect 8192 5932 8214 5964
rect 8138 5896 8214 5932
rect 8138 5864 8160 5896
rect 8192 5864 8214 5896
rect 8138 5828 8214 5864
rect 8138 5796 8160 5828
rect 8192 5796 8214 5828
rect 8138 5760 8214 5796
rect 8138 5728 8160 5760
rect 8192 5728 8214 5760
rect 8138 5692 8214 5728
rect 8138 5660 8160 5692
rect 8192 5660 8214 5692
rect 8138 5624 8214 5660
rect 8138 5592 8160 5624
rect 8192 5592 8214 5624
rect 8138 5556 8214 5592
rect 8138 5524 8160 5556
rect 8192 5524 8214 5556
rect 8138 5488 8214 5524
rect 8138 5456 8160 5488
rect 8192 5456 8214 5488
rect 8138 5420 8214 5456
rect 8138 5388 8160 5420
rect 8192 5388 8214 5420
rect 8138 5352 8214 5388
rect 8138 5320 8160 5352
rect 8192 5320 8214 5352
rect 8138 5282 8214 5320
rect 8314 6644 8390 6682
rect 8314 6612 8336 6644
rect 8368 6612 8390 6644
rect 8314 6576 8390 6612
rect 8314 6544 8336 6576
rect 8368 6544 8390 6576
rect 8314 6508 8390 6544
rect 8314 6476 8336 6508
rect 8368 6476 8390 6508
rect 8314 6440 8390 6476
rect 8314 6408 8336 6440
rect 8368 6408 8390 6440
rect 8314 6372 8390 6408
rect 8314 6340 8336 6372
rect 8368 6340 8390 6372
rect 8314 6304 8390 6340
rect 8314 6272 8336 6304
rect 8368 6272 8390 6304
rect 8314 6236 8390 6272
rect 8314 6204 8336 6236
rect 8368 6204 8390 6236
rect 8314 6168 8390 6204
rect 8314 6136 8336 6168
rect 8368 6136 8390 6168
rect 8314 6100 8390 6136
rect 8314 6068 8336 6100
rect 8368 6068 8390 6100
rect 8314 6032 8390 6068
rect 8314 6000 8336 6032
rect 8368 6000 8390 6032
rect 8314 5964 8390 6000
rect 8314 5932 8336 5964
rect 8368 5932 8390 5964
rect 8314 5896 8390 5932
rect 8314 5864 8336 5896
rect 8368 5864 8390 5896
rect 8314 5828 8390 5864
rect 8314 5796 8336 5828
rect 8368 5796 8390 5828
rect 8314 5760 8390 5796
rect 8314 5728 8336 5760
rect 8368 5728 8390 5760
rect 8314 5692 8390 5728
rect 8314 5660 8336 5692
rect 8368 5660 8390 5692
rect 8314 5624 8390 5660
rect 8314 5592 8336 5624
rect 8368 5592 8390 5624
rect 8314 5556 8390 5592
rect 8314 5524 8336 5556
rect 8368 5524 8390 5556
rect 8314 5488 8390 5524
rect 8314 5456 8336 5488
rect 8368 5456 8390 5488
rect 8314 5420 8390 5456
rect 8314 5388 8336 5420
rect 8368 5388 8390 5420
rect 8314 5352 8390 5388
rect 8314 5320 8336 5352
rect 8368 5320 8390 5352
rect 8314 5282 8390 5320
rect 8490 6644 8566 6682
rect 8490 6612 8512 6644
rect 8544 6612 8566 6644
rect 8490 6576 8566 6612
rect 8490 6544 8512 6576
rect 8544 6544 8566 6576
rect 8490 6508 8566 6544
rect 8490 6476 8512 6508
rect 8544 6476 8566 6508
rect 8490 6440 8566 6476
rect 8490 6408 8512 6440
rect 8544 6408 8566 6440
rect 8490 6372 8566 6408
rect 8490 6340 8512 6372
rect 8544 6340 8566 6372
rect 8490 6304 8566 6340
rect 8490 6272 8512 6304
rect 8544 6272 8566 6304
rect 8490 6236 8566 6272
rect 8490 6204 8512 6236
rect 8544 6204 8566 6236
rect 8490 6168 8566 6204
rect 8490 6136 8512 6168
rect 8544 6136 8566 6168
rect 8490 6100 8566 6136
rect 8490 6068 8512 6100
rect 8544 6068 8566 6100
rect 8490 6032 8566 6068
rect 8490 6000 8512 6032
rect 8544 6000 8566 6032
rect 8490 5964 8566 6000
rect 8490 5932 8512 5964
rect 8544 5932 8566 5964
rect 8490 5896 8566 5932
rect 8490 5864 8512 5896
rect 8544 5864 8566 5896
rect 8490 5828 8566 5864
rect 8490 5796 8512 5828
rect 8544 5796 8566 5828
rect 8490 5760 8566 5796
rect 8490 5728 8512 5760
rect 8544 5728 8566 5760
rect 8490 5692 8566 5728
rect 8490 5660 8512 5692
rect 8544 5660 8566 5692
rect 8490 5624 8566 5660
rect 8490 5592 8512 5624
rect 8544 5592 8566 5624
rect 8490 5556 8566 5592
rect 8490 5524 8512 5556
rect 8544 5524 8566 5556
rect 8490 5488 8566 5524
rect 8490 5456 8512 5488
rect 8544 5456 8566 5488
rect 8490 5420 8566 5456
rect 8490 5388 8512 5420
rect 8544 5388 8566 5420
rect 8490 5352 8566 5388
rect 8490 5320 8512 5352
rect 8544 5320 8566 5352
rect 8490 5282 8566 5320
rect 8666 6644 8742 6682
rect 8666 6612 8688 6644
rect 8720 6612 8742 6644
rect 8666 6576 8742 6612
rect 8666 6544 8688 6576
rect 8720 6544 8742 6576
rect 8666 6508 8742 6544
rect 8666 6476 8688 6508
rect 8720 6476 8742 6508
rect 8666 6440 8742 6476
rect 8666 6408 8688 6440
rect 8720 6408 8742 6440
rect 8666 6372 8742 6408
rect 8666 6340 8688 6372
rect 8720 6340 8742 6372
rect 8666 6304 8742 6340
rect 8666 6272 8688 6304
rect 8720 6272 8742 6304
rect 8666 6236 8742 6272
rect 8666 6204 8688 6236
rect 8720 6204 8742 6236
rect 8666 6168 8742 6204
rect 8666 6136 8688 6168
rect 8720 6136 8742 6168
rect 8666 6100 8742 6136
rect 8666 6068 8688 6100
rect 8720 6068 8742 6100
rect 8666 6032 8742 6068
rect 8666 6000 8688 6032
rect 8720 6000 8742 6032
rect 8666 5964 8742 6000
rect 8666 5932 8688 5964
rect 8720 5932 8742 5964
rect 8666 5896 8742 5932
rect 8666 5864 8688 5896
rect 8720 5864 8742 5896
rect 8666 5828 8742 5864
rect 8666 5796 8688 5828
rect 8720 5796 8742 5828
rect 8666 5760 8742 5796
rect 8666 5728 8688 5760
rect 8720 5728 8742 5760
rect 8666 5692 8742 5728
rect 8666 5660 8688 5692
rect 8720 5660 8742 5692
rect 8666 5624 8742 5660
rect 8666 5592 8688 5624
rect 8720 5592 8742 5624
rect 8666 5556 8742 5592
rect 8666 5524 8688 5556
rect 8720 5524 8742 5556
rect 8666 5488 8742 5524
rect 8666 5456 8688 5488
rect 8720 5456 8742 5488
rect 8666 5420 8742 5456
rect 8666 5388 8688 5420
rect 8720 5388 8742 5420
rect 8666 5352 8742 5388
rect 8666 5320 8688 5352
rect 8720 5320 8742 5352
rect 8666 5282 8742 5320
rect 8842 6644 8918 6682
rect 8842 6612 8864 6644
rect 8896 6612 8918 6644
rect 8842 6576 8918 6612
rect 8842 6544 8864 6576
rect 8896 6544 8918 6576
rect 8842 6508 8918 6544
rect 8842 6476 8864 6508
rect 8896 6476 8918 6508
rect 8842 6440 8918 6476
rect 8842 6408 8864 6440
rect 8896 6408 8918 6440
rect 8842 6372 8918 6408
rect 8842 6340 8864 6372
rect 8896 6340 8918 6372
rect 8842 6304 8918 6340
rect 8842 6272 8864 6304
rect 8896 6272 8918 6304
rect 8842 6236 8918 6272
rect 8842 6204 8864 6236
rect 8896 6204 8918 6236
rect 8842 6168 8918 6204
rect 8842 6136 8864 6168
rect 8896 6136 8918 6168
rect 8842 6100 8918 6136
rect 8842 6068 8864 6100
rect 8896 6068 8918 6100
rect 8842 6032 8918 6068
rect 8842 6000 8864 6032
rect 8896 6000 8918 6032
rect 8842 5964 8918 6000
rect 8842 5932 8864 5964
rect 8896 5932 8918 5964
rect 8842 5896 8918 5932
rect 8842 5864 8864 5896
rect 8896 5864 8918 5896
rect 8842 5828 8918 5864
rect 8842 5796 8864 5828
rect 8896 5796 8918 5828
rect 8842 5760 8918 5796
rect 8842 5728 8864 5760
rect 8896 5728 8918 5760
rect 8842 5692 8918 5728
rect 8842 5660 8864 5692
rect 8896 5660 8918 5692
rect 8842 5624 8918 5660
rect 8842 5592 8864 5624
rect 8896 5592 8918 5624
rect 8842 5556 8918 5592
rect 8842 5524 8864 5556
rect 8896 5524 8918 5556
rect 8842 5488 8918 5524
rect 8842 5456 8864 5488
rect 8896 5456 8918 5488
rect 8842 5420 8918 5456
rect 8842 5388 8864 5420
rect 8896 5388 8918 5420
rect 8842 5352 8918 5388
rect 8842 5320 8864 5352
rect 8896 5320 8918 5352
rect 8842 5282 8918 5320
rect 9018 6644 9094 6682
rect 9018 6612 9040 6644
rect 9072 6612 9094 6644
rect 9018 6576 9094 6612
rect 9018 6544 9040 6576
rect 9072 6544 9094 6576
rect 9018 6508 9094 6544
rect 9018 6476 9040 6508
rect 9072 6476 9094 6508
rect 9018 6440 9094 6476
rect 9018 6408 9040 6440
rect 9072 6408 9094 6440
rect 9018 6372 9094 6408
rect 9018 6340 9040 6372
rect 9072 6340 9094 6372
rect 9018 6304 9094 6340
rect 9018 6272 9040 6304
rect 9072 6272 9094 6304
rect 9018 6236 9094 6272
rect 9018 6204 9040 6236
rect 9072 6204 9094 6236
rect 9018 6168 9094 6204
rect 9018 6136 9040 6168
rect 9072 6136 9094 6168
rect 9018 6100 9094 6136
rect 9018 6068 9040 6100
rect 9072 6068 9094 6100
rect 9018 6032 9094 6068
rect 9018 6000 9040 6032
rect 9072 6000 9094 6032
rect 9018 5964 9094 6000
rect 9018 5932 9040 5964
rect 9072 5932 9094 5964
rect 9018 5896 9094 5932
rect 9018 5864 9040 5896
rect 9072 5864 9094 5896
rect 9018 5828 9094 5864
rect 9018 5796 9040 5828
rect 9072 5796 9094 5828
rect 9018 5760 9094 5796
rect 9018 5728 9040 5760
rect 9072 5728 9094 5760
rect 9018 5692 9094 5728
rect 9018 5660 9040 5692
rect 9072 5660 9094 5692
rect 9018 5624 9094 5660
rect 9018 5592 9040 5624
rect 9072 5592 9094 5624
rect 9018 5556 9094 5592
rect 9018 5524 9040 5556
rect 9072 5524 9094 5556
rect 9018 5488 9094 5524
rect 9018 5456 9040 5488
rect 9072 5456 9094 5488
rect 9018 5420 9094 5456
rect 9018 5388 9040 5420
rect 9072 5388 9094 5420
rect 9018 5352 9094 5388
rect 9018 5320 9040 5352
rect 9072 5320 9094 5352
rect 9018 5282 9094 5320
rect 9194 6644 9270 6682
rect 9194 6612 9216 6644
rect 9248 6612 9270 6644
rect 9194 6576 9270 6612
rect 9194 6544 9216 6576
rect 9248 6544 9270 6576
rect 9194 6508 9270 6544
rect 9194 6476 9216 6508
rect 9248 6476 9270 6508
rect 9194 6440 9270 6476
rect 9194 6408 9216 6440
rect 9248 6408 9270 6440
rect 9194 6372 9270 6408
rect 9194 6340 9216 6372
rect 9248 6340 9270 6372
rect 9194 6304 9270 6340
rect 9194 6272 9216 6304
rect 9248 6272 9270 6304
rect 9194 6236 9270 6272
rect 9194 6204 9216 6236
rect 9248 6204 9270 6236
rect 9194 6168 9270 6204
rect 9194 6136 9216 6168
rect 9248 6136 9270 6168
rect 9194 6100 9270 6136
rect 9194 6068 9216 6100
rect 9248 6068 9270 6100
rect 9194 6032 9270 6068
rect 9194 6000 9216 6032
rect 9248 6000 9270 6032
rect 9194 5964 9270 6000
rect 9194 5932 9216 5964
rect 9248 5932 9270 5964
rect 9194 5896 9270 5932
rect 9194 5864 9216 5896
rect 9248 5864 9270 5896
rect 9194 5828 9270 5864
rect 9194 5796 9216 5828
rect 9248 5796 9270 5828
rect 9194 5760 9270 5796
rect 9194 5728 9216 5760
rect 9248 5728 9270 5760
rect 9194 5692 9270 5728
rect 9194 5660 9216 5692
rect 9248 5660 9270 5692
rect 9194 5624 9270 5660
rect 9194 5592 9216 5624
rect 9248 5592 9270 5624
rect 9194 5556 9270 5592
rect 9194 5524 9216 5556
rect 9248 5524 9270 5556
rect 9194 5488 9270 5524
rect 9194 5456 9216 5488
rect 9248 5456 9270 5488
rect 9194 5420 9270 5456
rect 9194 5388 9216 5420
rect 9248 5388 9270 5420
rect 9194 5352 9270 5388
rect 9194 5320 9216 5352
rect 9248 5320 9270 5352
rect 9194 5282 9270 5320
rect 9370 6644 9446 6682
rect 9370 6612 9392 6644
rect 9424 6612 9446 6644
rect 9370 6576 9446 6612
rect 9370 6544 9392 6576
rect 9424 6544 9446 6576
rect 9370 6508 9446 6544
rect 9370 6476 9392 6508
rect 9424 6476 9446 6508
rect 9370 6440 9446 6476
rect 9370 6408 9392 6440
rect 9424 6408 9446 6440
rect 9370 6372 9446 6408
rect 9370 6340 9392 6372
rect 9424 6340 9446 6372
rect 9370 6304 9446 6340
rect 9370 6272 9392 6304
rect 9424 6272 9446 6304
rect 9370 6236 9446 6272
rect 9370 6204 9392 6236
rect 9424 6204 9446 6236
rect 9370 6168 9446 6204
rect 9370 6136 9392 6168
rect 9424 6136 9446 6168
rect 9370 6100 9446 6136
rect 9370 6068 9392 6100
rect 9424 6068 9446 6100
rect 9370 6032 9446 6068
rect 9370 6000 9392 6032
rect 9424 6000 9446 6032
rect 9370 5964 9446 6000
rect 9370 5932 9392 5964
rect 9424 5932 9446 5964
rect 9370 5896 9446 5932
rect 9370 5864 9392 5896
rect 9424 5864 9446 5896
rect 9370 5828 9446 5864
rect 9370 5796 9392 5828
rect 9424 5796 9446 5828
rect 9370 5760 9446 5796
rect 9370 5728 9392 5760
rect 9424 5728 9446 5760
rect 9370 5692 9446 5728
rect 9370 5660 9392 5692
rect 9424 5660 9446 5692
rect 9370 5624 9446 5660
rect 9370 5592 9392 5624
rect 9424 5592 9446 5624
rect 9370 5556 9446 5592
rect 9370 5524 9392 5556
rect 9424 5524 9446 5556
rect 9370 5488 9446 5524
rect 9370 5456 9392 5488
rect 9424 5456 9446 5488
rect 9370 5420 9446 5456
rect 9370 5388 9392 5420
rect 9424 5388 9446 5420
rect 9370 5352 9446 5388
rect 9370 5320 9392 5352
rect 9424 5320 9446 5352
rect 9370 5282 9446 5320
rect 9546 6644 9622 6682
rect 9546 6612 9568 6644
rect 9600 6612 9622 6644
rect 9546 6576 9622 6612
rect 9546 6544 9568 6576
rect 9600 6544 9622 6576
rect 9546 6508 9622 6544
rect 9546 6476 9568 6508
rect 9600 6476 9622 6508
rect 9546 6440 9622 6476
rect 9546 6408 9568 6440
rect 9600 6408 9622 6440
rect 9546 6372 9622 6408
rect 9546 6340 9568 6372
rect 9600 6340 9622 6372
rect 9546 6304 9622 6340
rect 9546 6272 9568 6304
rect 9600 6272 9622 6304
rect 9546 6236 9622 6272
rect 9546 6204 9568 6236
rect 9600 6204 9622 6236
rect 9546 6168 9622 6204
rect 9546 6136 9568 6168
rect 9600 6136 9622 6168
rect 9546 6100 9622 6136
rect 9546 6068 9568 6100
rect 9600 6068 9622 6100
rect 9546 6032 9622 6068
rect 9546 6000 9568 6032
rect 9600 6000 9622 6032
rect 9546 5964 9622 6000
rect 9546 5932 9568 5964
rect 9600 5932 9622 5964
rect 9546 5896 9622 5932
rect 9546 5864 9568 5896
rect 9600 5864 9622 5896
rect 9546 5828 9622 5864
rect 9546 5796 9568 5828
rect 9600 5796 9622 5828
rect 9546 5760 9622 5796
rect 9546 5728 9568 5760
rect 9600 5728 9622 5760
rect 9546 5692 9622 5728
rect 9546 5660 9568 5692
rect 9600 5660 9622 5692
rect 9546 5624 9622 5660
rect 9546 5592 9568 5624
rect 9600 5592 9622 5624
rect 9546 5556 9622 5592
rect 9546 5524 9568 5556
rect 9600 5524 9622 5556
rect 9546 5488 9622 5524
rect 9546 5456 9568 5488
rect 9600 5456 9622 5488
rect 9546 5420 9622 5456
rect 9546 5388 9568 5420
rect 9600 5388 9622 5420
rect 9546 5352 9622 5388
rect 9546 5320 9568 5352
rect 9600 5320 9622 5352
rect 9546 5282 9622 5320
rect 9722 6644 9798 6682
rect 9722 6612 9744 6644
rect 9776 6612 9798 6644
rect 9722 6576 9798 6612
rect 9722 6544 9744 6576
rect 9776 6544 9798 6576
rect 9722 6508 9798 6544
rect 9722 6476 9744 6508
rect 9776 6476 9798 6508
rect 9722 6440 9798 6476
rect 9722 6408 9744 6440
rect 9776 6408 9798 6440
rect 9722 6372 9798 6408
rect 9722 6340 9744 6372
rect 9776 6340 9798 6372
rect 9722 6304 9798 6340
rect 9722 6272 9744 6304
rect 9776 6272 9798 6304
rect 9722 6236 9798 6272
rect 9722 6204 9744 6236
rect 9776 6204 9798 6236
rect 9722 6168 9798 6204
rect 9722 6136 9744 6168
rect 9776 6136 9798 6168
rect 9722 6100 9798 6136
rect 9722 6068 9744 6100
rect 9776 6068 9798 6100
rect 9722 6032 9798 6068
rect 9722 6000 9744 6032
rect 9776 6000 9798 6032
rect 9722 5964 9798 6000
rect 9722 5932 9744 5964
rect 9776 5932 9798 5964
rect 9722 5896 9798 5932
rect 9722 5864 9744 5896
rect 9776 5864 9798 5896
rect 9722 5828 9798 5864
rect 9722 5796 9744 5828
rect 9776 5796 9798 5828
rect 9722 5760 9798 5796
rect 9722 5728 9744 5760
rect 9776 5728 9798 5760
rect 9722 5692 9798 5728
rect 9722 5660 9744 5692
rect 9776 5660 9798 5692
rect 9722 5624 9798 5660
rect 9722 5592 9744 5624
rect 9776 5592 9798 5624
rect 9722 5556 9798 5592
rect 9722 5524 9744 5556
rect 9776 5524 9798 5556
rect 9722 5488 9798 5524
rect 9722 5456 9744 5488
rect 9776 5456 9798 5488
rect 9722 5420 9798 5456
rect 9722 5388 9744 5420
rect 9776 5388 9798 5420
rect 9722 5352 9798 5388
rect 9722 5320 9744 5352
rect 9776 5320 9798 5352
rect 9722 5282 9798 5320
rect 9898 6644 9974 6682
rect 9898 6612 9920 6644
rect 9952 6612 9974 6644
rect 9898 6576 9974 6612
rect 9898 6544 9920 6576
rect 9952 6544 9974 6576
rect 9898 6508 9974 6544
rect 9898 6476 9920 6508
rect 9952 6476 9974 6508
rect 9898 6440 9974 6476
rect 9898 6408 9920 6440
rect 9952 6408 9974 6440
rect 9898 6372 9974 6408
rect 9898 6340 9920 6372
rect 9952 6340 9974 6372
rect 9898 6304 9974 6340
rect 9898 6272 9920 6304
rect 9952 6272 9974 6304
rect 9898 6236 9974 6272
rect 9898 6204 9920 6236
rect 9952 6204 9974 6236
rect 9898 6168 9974 6204
rect 9898 6136 9920 6168
rect 9952 6136 9974 6168
rect 9898 6100 9974 6136
rect 9898 6068 9920 6100
rect 9952 6068 9974 6100
rect 9898 6032 9974 6068
rect 9898 6000 9920 6032
rect 9952 6000 9974 6032
rect 9898 5964 9974 6000
rect 9898 5932 9920 5964
rect 9952 5932 9974 5964
rect 9898 5896 9974 5932
rect 9898 5864 9920 5896
rect 9952 5864 9974 5896
rect 9898 5828 9974 5864
rect 9898 5796 9920 5828
rect 9952 5796 9974 5828
rect 9898 5760 9974 5796
rect 9898 5728 9920 5760
rect 9952 5728 9974 5760
rect 9898 5692 9974 5728
rect 9898 5660 9920 5692
rect 9952 5660 9974 5692
rect 9898 5624 9974 5660
rect 9898 5592 9920 5624
rect 9952 5592 9974 5624
rect 9898 5556 9974 5592
rect 9898 5524 9920 5556
rect 9952 5524 9974 5556
rect 9898 5488 9974 5524
rect 9898 5456 9920 5488
rect 9952 5456 9974 5488
rect 9898 5420 9974 5456
rect 9898 5388 9920 5420
rect 9952 5388 9974 5420
rect 9898 5352 9974 5388
rect 9898 5320 9920 5352
rect 9952 5320 9974 5352
rect 9898 5282 9974 5320
rect 10074 6644 10150 6682
rect 10074 6612 10096 6644
rect 10128 6612 10150 6644
rect 10074 6576 10150 6612
rect 10074 6544 10096 6576
rect 10128 6544 10150 6576
rect 10074 6508 10150 6544
rect 10074 6476 10096 6508
rect 10128 6476 10150 6508
rect 10074 6440 10150 6476
rect 10074 6408 10096 6440
rect 10128 6408 10150 6440
rect 10074 6372 10150 6408
rect 10074 6340 10096 6372
rect 10128 6340 10150 6372
rect 10074 6304 10150 6340
rect 10074 6272 10096 6304
rect 10128 6272 10150 6304
rect 10074 6236 10150 6272
rect 10074 6204 10096 6236
rect 10128 6204 10150 6236
rect 10074 6168 10150 6204
rect 10074 6136 10096 6168
rect 10128 6136 10150 6168
rect 10074 6100 10150 6136
rect 10074 6068 10096 6100
rect 10128 6068 10150 6100
rect 10074 6032 10150 6068
rect 10074 6000 10096 6032
rect 10128 6000 10150 6032
rect 10074 5964 10150 6000
rect 10074 5932 10096 5964
rect 10128 5932 10150 5964
rect 10074 5896 10150 5932
rect 10074 5864 10096 5896
rect 10128 5864 10150 5896
rect 10074 5828 10150 5864
rect 10074 5796 10096 5828
rect 10128 5796 10150 5828
rect 10074 5760 10150 5796
rect 10074 5728 10096 5760
rect 10128 5728 10150 5760
rect 10074 5692 10150 5728
rect 10074 5660 10096 5692
rect 10128 5660 10150 5692
rect 10074 5624 10150 5660
rect 10074 5592 10096 5624
rect 10128 5592 10150 5624
rect 10074 5556 10150 5592
rect 10074 5524 10096 5556
rect 10128 5524 10150 5556
rect 10074 5488 10150 5524
rect 10074 5456 10096 5488
rect 10128 5456 10150 5488
rect 10074 5420 10150 5456
rect 10074 5388 10096 5420
rect 10128 5388 10150 5420
rect 10074 5352 10150 5388
rect 10074 5320 10096 5352
rect 10128 5320 10150 5352
rect 10074 5282 10150 5320
rect 10250 6644 10326 6682
rect 10250 6612 10272 6644
rect 10304 6612 10326 6644
rect 10250 6576 10326 6612
rect 10250 6544 10272 6576
rect 10304 6544 10326 6576
rect 10250 6508 10326 6544
rect 10250 6476 10272 6508
rect 10304 6476 10326 6508
rect 10250 6440 10326 6476
rect 10250 6408 10272 6440
rect 10304 6408 10326 6440
rect 10250 6372 10326 6408
rect 10250 6340 10272 6372
rect 10304 6340 10326 6372
rect 10250 6304 10326 6340
rect 10250 6272 10272 6304
rect 10304 6272 10326 6304
rect 10250 6236 10326 6272
rect 10250 6204 10272 6236
rect 10304 6204 10326 6236
rect 10250 6168 10326 6204
rect 10250 6136 10272 6168
rect 10304 6136 10326 6168
rect 10250 6100 10326 6136
rect 10250 6068 10272 6100
rect 10304 6068 10326 6100
rect 10250 6032 10326 6068
rect 10250 6000 10272 6032
rect 10304 6000 10326 6032
rect 10250 5964 10326 6000
rect 10250 5932 10272 5964
rect 10304 5932 10326 5964
rect 10250 5896 10326 5932
rect 10250 5864 10272 5896
rect 10304 5864 10326 5896
rect 10250 5828 10326 5864
rect 10250 5796 10272 5828
rect 10304 5796 10326 5828
rect 10250 5760 10326 5796
rect 10250 5728 10272 5760
rect 10304 5728 10326 5760
rect 10250 5692 10326 5728
rect 10250 5660 10272 5692
rect 10304 5660 10326 5692
rect 10250 5624 10326 5660
rect 10250 5592 10272 5624
rect 10304 5592 10326 5624
rect 10250 5556 10326 5592
rect 10250 5524 10272 5556
rect 10304 5524 10326 5556
rect 10250 5488 10326 5524
rect 10250 5456 10272 5488
rect 10304 5456 10326 5488
rect 10250 5420 10326 5456
rect 10250 5388 10272 5420
rect 10304 5388 10326 5420
rect 10250 5352 10326 5388
rect 10250 5320 10272 5352
rect 10304 5320 10326 5352
rect 10250 5282 10326 5320
rect 10426 6644 10502 6682
rect 10426 6612 10448 6644
rect 10480 6612 10502 6644
rect 10426 6576 10502 6612
rect 10426 6544 10448 6576
rect 10480 6544 10502 6576
rect 10426 6508 10502 6544
rect 10426 6476 10448 6508
rect 10480 6476 10502 6508
rect 10426 6440 10502 6476
rect 10426 6408 10448 6440
rect 10480 6408 10502 6440
rect 10426 6372 10502 6408
rect 10426 6340 10448 6372
rect 10480 6340 10502 6372
rect 10426 6304 10502 6340
rect 10426 6272 10448 6304
rect 10480 6272 10502 6304
rect 10426 6236 10502 6272
rect 10426 6204 10448 6236
rect 10480 6204 10502 6236
rect 10426 6168 10502 6204
rect 10426 6136 10448 6168
rect 10480 6136 10502 6168
rect 10426 6100 10502 6136
rect 10426 6068 10448 6100
rect 10480 6068 10502 6100
rect 10426 6032 10502 6068
rect 10426 6000 10448 6032
rect 10480 6000 10502 6032
rect 10426 5964 10502 6000
rect 10426 5932 10448 5964
rect 10480 5932 10502 5964
rect 10426 5896 10502 5932
rect 10426 5864 10448 5896
rect 10480 5864 10502 5896
rect 10426 5828 10502 5864
rect 10426 5796 10448 5828
rect 10480 5796 10502 5828
rect 10426 5760 10502 5796
rect 10426 5728 10448 5760
rect 10480 5728 10502 5760
rect 10426 5692 10502 5728
rect 10426 5660 10448 5692
rect 10480 5660 10502 5692
rect 10426 5624 10502 5660
rect 10426 5592 10448 5624
rect 10480 5592 10502 5624
rect 10426 5556 10502 5592
rect 10426 5524 10448 5556
rect 10480 5524 10502 5556
rect 10426 5488 10502 5524
rect 10426 5456 10448 5488
rect 10480 5456 10502 5488
rect 10426 5420 10502 5456
rect 10426 5388 10448 5420
rect 10480 5388 10502 5420
rect 10426 5352 10502 5388
rect 10426 5320 10448 5352
rect 10480 5320 10502 5352
rect 10426 5282 10502 5320
rect 10602 6644 10678 6682
rect 10602 6612 10624 6644
rect 10656 6612 10678 6644
rect 10602 6576 10678 6612
rect 10602 6544 10624 6576
rect 10656 6544 10678 6576
rect 10602 6508 10678 6544
rect 10602 6476 10624 6508
rect 10656 6476 10678 6508
rect 10602 6440 10678 6476
rect 10602 6408 10624 6440
rect 10656 6408 10678 6440
rect 10602 6372 10678 6408
rect 10602 6340 10624 6372
rect 10656 6340 10678 6372
rect 10602 6304 10678 6340
rect 10602 6272 10624 6304
rect 10656 6272 10678 6304
rect 10602 6236 10678 6272
rect 10602 6204 10624 6236
rect 10656 6204 10678 6236
rect 10602 6168 10678 6204
rect 10602 6136 10624 6168
rect 10656 6136 10678 6168
rect 10602 6100 10678 6136
rect 10602 6068 10624 6100
rect 10656 6068 10678 6100
rect 10602 6032 10678 6068
rect 10602 6000 10624 6032
rect 10656 6000 10678 6032
rect 10602 5964 10678 6000
rect 10602 5932 10624 5964
rect 10656 5932 10678 5964
rect 10602 5896 10678 5932
rect 10602 5864 10624 5896
rect 10656 5864 10678 5896
rect 10602 5828 10678 5864
rect 10602 5796 10624 5828
rect 10656 5796 10678 5828
rect 10602 5760 10678 5796
rect 10602 5728 10624 5760
rect 10656 5728 10678 5760
rect 10602 5692 10678 5728
rect 10602 5660 10624 5692
rect 10656 5660 10678 5692
rect 10602 5624 10678 5660
rect 10602 5592 10624 5624
rect 10656 5592 10678 5624
rect 10602 5556 10678 5592
rect 10602 5524 10624 5556
rect 10656 5524 10678 5556
rect 10602 5488 10678 5524
rect 10602 5456 10624 5488
rect 10656 5456 10678 5488
rect 10602 5420 10678 5456
rect 10602 5388 10624 5420
rect 10656 5388 10678 5420
rect 10602 5352 10678 5388
rect 10602 5320 10624 5352
rect 10656 5320 10678 5352
rect 10602 5282 10678 5320
rect 10778 6644 10854 6682
rect 10778 6612 10800 6644
rect 10832 6612 10854 6644
rect 10778 6576 10854 6612
rect 10778 6544 10800 6576
rect 10832 6544 10854 6576
rect 10778 6508 10854 6544
rect 10778 6476 10800 6508
rect 10832 6476 10854 6508
rect 10778 6440 10854 6476
rect 10778 6408 10800 6440
rect 10832 6408 10854 6440
rect 10778 6372 10854 6408
rect 10778 6340 10800 6372
rect 10832 6340 10854 6372
rect 10778 6304 10854 6340
rect 10778 6272 10800 6304
rect 10832 6272 10854 6304
rect 10778 6236 10854 6272
rect 10778 6204 10800 6236
rect 10832 6204 10854 6236
rect 10778 6168 10854 6204
rect 10778 6136 10800 6168
rect 10832 6136 10854 6168
rect 10778 6100 10854 6136
rect 10778 6068 10800 6100
rect 10832 6068 10854 6100
rect 10778 6032 10854 6068
rect 10778 6000 10800 6032
rect 10832 6000 10854 6032
rect 10778 5964 10854 6000
rect 10778 5932 10800 5964
rect 10832 5932 10854 5964
rect 10778 5896 10854 5932
rect 10778 5864 10800 5896
rect 10832 5864 10854 5896
rect 10778 5828 10854 5864
rect 10778 5796 10800 5828
rect 10832 5796 10854 5828
rect 10778 5760 10854 5796
rect 10778 5728 10800 5760
rect 10832 5728 10854 5760
rect 10778 5692 10854 5728
rect 10778 5660 10800 5692
rect 10832 5660 10854 5692
rect 10778 5624 10854 5660
rect 10778 5592 10800 5624
rect 10832 5592 10854 5624
rect 10778 5556 10854 5592
rect 10778 5524 10800 5556
rect 10832 5524 10854 5556
rect 10778 5488 10854 5524
rect 10778 5456 10800 5488
rect 10832 5456 10854 5488
rect 10778 5420 10854 5456
rect 10778 5388 10800 5420
rect 10832 5388 10854 5420
rect 10778 5352 10854 5388
rect 10778 5320 10800 5352
rect 10832 5320 10854 5352
rect 10778 5282 10854 5320
rect 10954 6644 11030 6682
rect 10954 6612 10976 6644
rect 11008 6612 11030 6644
rect 10954 6576 11030 6612
rect 10954 6544 10976 6576
rect 11008 6544 11030 6576
rect 10954 6508 11030 6544
rect 10954 6476 10976 6508
rect 11008 6476 11030 6508
rect 10954 6440 11030 6476
rect 10954 6408 10976 6440
rect 11008 6408 11030 6440
rect 10954 6372 11030 6408
rect 10954 6340 10976 6372
rect 11008 6340 11030 6372
rect 10954 6304 11030 6340
rect 10954 6272 10976 6304
rect 11008 6272 11030 6304
rect 10954 6236 11030 6272
rect 10954 6204 10976 6236
rect 11008 6204 11030 6236
rect 10954 6168 11030 6204
rect 10954 6136 10976 6168
rect 11008 6136 11030 6168
rect 10954 6100 11030 6136
rect 10954 6068 10976 6100
rect 11008 6068 11030 6100
rect 10954 6032 11030 6068
rect 10954 6000 10976 6032
rect 11008 6000 11030 6032
rect 10954 5964 11030 6000
rect 10954 5932 10976 5964
rect 11008 5932 11030 5964
rect 10954 5896 11030 5932
rect 10954 5864 10976 5896
rect 11008 5864 11030 5896
rect 10954 5828 11030 5864
rect 10954 5796 10976 5828
rect 11008 5796 11030 5828
rect 10954 5760 11030 5796
rect 10954 5728 10976 5760
rect 11008 5728 11030 5760
rect 10954 5692 11030 5728
rect 10954 5660 10976 5692
rect 11008 5660 11030 5692
rect 10954 5624 11030 5660
rect 10954 5592 10976 5624
rect 11008 5592 11030 5624
rect 10954 5556 11030 5592
rect 10954 5524 10976 5556
rect 11008 5524 11030 5556
rect 10954 5488 11030 5524
rect 10954 5456 10976 5488
rect 11008 5456 11030 5488
rect 10954 5420 11030 5456
rect 10954 5388 10976 5420
rect 11008 5388 11030 5420
rect 10954 5352 11030 5388
rect 10954 5320 10976 5352
rect 11008 5320 11030 5352
rect 10954 5282 11030 5320
rect 11130 6644 11206 6682
rect 11130 6612 11152 6644
rect 11184 6612 11206 6644
rect 11130 6576 11206 6612
rect 11130 6544 11152 6576
rect 11184 6544 11206 6576
rect 11130 6508 11206 6544
rect 11130 6476 11152 6508
rect 11184 6476 11206 6508
rect 11130 6440 11206 6476
rect 11130 6408 11152 6440
rect 11184 6408 11206 6440
rect 11130 6372 11206 6408
rect 11130 6340 11152 6372
rect 11184 6340 11206 6372
rect 11130 6304 11206 6340
rect 11130 6272 11152 6304
rect 11184 6272 11206 6304
rect 11130 6236 11206 6272
rect 11130 6204 11152 6236
rect 11184 6204 11206 6236
rect 11130 6168 11206 6204
rect 11130 6136 11152 6168
rect 11184 6136 11206 6168
rect 11130 6100 11206 6136
rect 11130 6068 11152 6100
rect 11184 6068 11206 6100
rect 11130 6032 11206 6068
rect 11130 6000 11152 6032
rect 11184 6000 11206 6032
rect 11130 5964 11206 6000
rect 11130 5932 11152 5964
rect 11184 5932 11206 5964
rect 11130 5896 11206 5932
rect 11130 5864 11152 5896
rect 11184 5864 11206 5896
rect 11130 5828 11206 5864
rect 11130 5796 11152 5828
rect 11184 5796 11206 5828
rect 11130 5760 11206 5796
rect 11130 5728 11152 5760
rect 11184 5728 11206 5760
rect 11130 5692 11206 5728
rect 11130 5660 11152 5692
rect 11184 5660 11206 5692
rect 11130 5624 11206 5660
rect 11130 5592 11152 5624
rect 11184 5592 11206 5624
rect 11130 5556 11206 5592
rect 11130 5524 11152 5556
rect 11184 5524 11206 5556
rect 11130 5488 11206 5524
rect 11130 5456 11152 5488
rect 11184 5456 11206 5488
rect 11130 5420 11206 5456
rect 11130 5388 11152 5420
rect 11184 5388 11206 5420
rect 11130 5352 11206 5388
rect 11130 5320 11152 5352
rect 11184 5320 11206 5352
rect 11130 5282 11206 5320
rect 11306 6644 11382 6682
rect 11306 6612 11328 6644
rect 11360 6612 11382 6644
rect 11306 6576 11382 6612
rect 11306 6544 11328 6576
rect 11360 6544 11382 6576
rect 11306 6508 11382 6544
rect 11306 6476 11328 6508
rect 11360 6476 11382 6508
rect 11306 6440 11382 6476
rect 11306 6408 11328 6440
rect 11360 6408 11382 6440
rect 11306 6372 11382 6408
rect 11306 6340 11328 6372
rect 11360 6340 11382 6372
rect 11306 6304 11382 6340
rect 11306 6272 11328 6304
rect 11360 6272 11382 6304
rect 11306 6236 11382 6272
rect 11306 6204 11328 6236
rect 11360 6204 11382 6236
rect 11306 6168 11382 6204
rect 11306 6136 11328 6168
rect 11360 6136 11382 6168
rect 11306 6100 11382 6136
rect 11306 6068 11328 6100
rect 11360 6068 11382 6100
rect 11306 6032 11382 6068
rect 11306 6000 11328 6032
rect 11360 6000 11382 6032
rect 11306 5964 11382 6000
rect 11306 5932 11328 5964
rect 11360 5932 11382 5964
rect 11306 5896 11382 5932
rect 11306 5864 11328 5896
rect 11360 5864 11382 5896
rect 11306 5828 11382 5864
rect 11306 5796 11328 5828
rect 11360 5796 11382 5828
rect 11306 5760 11382 5796
rect 11306 5728 11328 5760
rect 11360 5728 11382 5760
rect 11306 5692 11382 5728
rect 11306 5660 11328 5692
rect 11360 5660 11382 5692
rect 11306 5624 11382 5660
rect 11306 5592 11328 5624
rect 11360 5592 11382 5624
rect 11306 5556 11382 5592
rect 11306 5524 11328 5556
rect 11360 5524 11382 5556
rect 11306 5488 11382 5524
rect 11306 5456 11328 5488
rect 11360 5456 11382 5488
rect 11306 5420 11382 5456
rect 11306 5388 11328 5420
rect 11360 5388 11382 5420
rect 11306 5352 11382 5388
rect 11306 5320 11328 5352
rect 11360 5320 11382 5352
rect 11306 5282 11382 5320
rect 11482 6644 11558 6682
rect 11482 6612 11504 6644
rect 11536 6612 11558 6644
rect 11482 6576 11558 6612
rect 11482 6544 11504 6576
rect 11536 6544 11558 6576
rect 11482 6508 11558 6544
rect 11482 6476 11504 6508
rect 11536 6476 11558 6508
rect 11482 6440 11558 6476
rect 11482 6408 11504 6440
rect 11536 6408 11558 6440
rect 11482 6372 11558 6408
rect 11482 6340 11504 6372
rect 11536 6340 11558 6372
rect 11482 6304 11558 6340
rect 11482 6272 11504 6304
rect 11536 6272 11558 6304
rect 11482 6236 11558 6272
rect 11482 6204 11504 6236
rect 11536 6204 11558 6236
rect 11482 6168 11558 6204
rect 11482 6136 11504 6168
rect 11536 6136 11558 6168
rect 11482 6100 11558 6136
rect 11482 6068 11504 6100
rect 11536 6068 11558 6100
rect 11482 6032 11558 6068
rect 11482 6000 11504 6032
rect 11536 6000 11558 6032
rect 11482 5964 11558 6000
rect 11482 5932 11504 5964
rect 11536 5932 11558 5964
rect 11482 5896 11558 5932
rect 11482 5864 11504 5896
rect 11536 5864 11558 5896
rect 11482 5828 11558 5864
rect 11482 5796 11504 5828
rect 11536 5796 11558 5828
rect 11482 5760 11558 5796
rect 11482 5728 11504 5760
rect 11536 5728 11558 5760
rect 11482 5692 11558 5728
rect 11482 5660 11504 5692
rect 11536 5660 11558 5692
rect 11482 5624 11558 5660
rect 11482 5592 11504 5624
rect 11536 5592 11558 5624
rect 11482 5556 11558 5592
rect 11482 5524 11504 5556
rect 11536 5524 11558 5556
rect 11482 5488 11558 5524
rect 11482 5456 11504 5488
rect 11536 5456 11558 5488
rect 11482 5420 11558 5456
rect 11482 5388 11504 5420
rect 11536 5388 11558 5420
rect 11482 5352 11558 5388
rect 11482 5320 11504 5352
rect 11536 5320 11558 5352
rect 11482 5282 11558 5320
rect 11658 6644 11734 6682
rect 11658 6612 11680 6644
rect 11712 6612 11734 6644
rect 11658 6576 11734 6612
rect 11658 6544 11680 6576
rect 11712 6544 11734 6576
rect 11658 6508 11734 6544
rect 11658 6476 11680 6508
rect 11712 6476 11734 6508
rect 11658 6440 11734 6476
rect 11658 6408 11680 6440
rect 11712 6408 11734 6440
rect 11658 6372 11734 6408
rect 11658 6340 11680 6372
rect 11712 6340 11734 6372
rect 11658 6304 11734 6340
rect 11658 6272 11680 6304
rect 11712 6272 11734 6304
rect 11658 6236 11734 6272
rect 11658 6204 11680 6236
rect 11712 6204 11734 6236
rect 11658 6168 11734 6204
rect 11658 6136 11680 6168
rect 11712 6136 11734 6168
rect 11658 6100 11734 6136
rect 11658 6068 11680 6100
rect 11712 6068 11734 6100
rect 11658 6032 11734 6068
rect 11658 6000 11680 6032
rect 11712 6000 11734 6032
rect 11658 5964 11734 6000
rect 11658 5932 11680 5964
rect 11712 5932 11734 5964
rect 11658 5896 11734 5932
rect 11658 5864 11680 5896
rect 11712 5864 11734 5896
rect 11658 5828 11734 5864
rect 11658 5796 11680 5828
rect 11712 5796 11734 5828
rect 11658 5760 11734 5796
rect 11658 5728 11680 5760
rect 11712 5728 11734 5760
rect 11658 5692 11734 5728
rect 11658 5660 11680 5692
rect 11712 5660 11734 5692
rect 11658 5624 11734 5660
rect 11658 5592 11680 5624
rect 11712 5592 11734 5624
rect 11658 5556 11734 5592
rect 11658 5524 11680 5556
rect 11712 5524 11734 5556
rect 11658 5488 11734 5524
rect 11658 5456 11680 5488
rect 11712 5456 11734 5488
rect 11658 5420 11734 5456
rect 11658 5388 11680 5420
rect 11712 5388 11734 5420
rect 11658 5352 11734 5388
rect 11658 5320 11680 5352
rect 11712 5320 11734 5352
rect 11658 5282 11734 5320
rect 11834 6644 11910 6682
rect 11834 6612 11856 6644
rect 11888 6612 11910 6644
rect 11834 6576 11910 6612
rect 11834 6544 11856 6576
rect 11888 6544 11910 6576
rect 11834 6508 11910 6544
rect 11834 6476 11856 6508
rect 11888 6476 11910 6508
rect 11834 6440 11910 6476
rect 11834 6408 11856 6440
rect 11888 6408 11910 6440
rect 11834 6372 11910 6408
rect 11834 6340 11856 6372
rect 11888 6340 11910 6372
rect 11834 6304 11910 6340
rect 11834 6272 11856 6304
rect 11888 6272 11910 6304
rect 11834 6236 11910 6272
rect 11834 6204 11856 6236
rect 11888 6204 11910 6236
rect 11834 6168 11910 6204
rect 11834 6136 11856 6168
rect 11888 6136 11910 6168
rect 11834 6100 11910 6136
rect 11834 6068 11856 6100
rect 11888 6068 11910 6100
rect 11834 6032 11910 6068
rect 11834 6000 11856 6032
rect 11888 6000 11910 6032
rect 11834 5964 11910 6000
rect 11834 5932 11856 5964
rect 11888 5932 11910 5964
rect 11834 5896 11910 5932
rect 11834 5864 11856 5896
rect 11888 5864 11910 5896
rect 11834 5828 11910 5864
rect 11834 5796 11856 5828
rect 11888 5796 11910 5828
rect 11834 5760 11910 5796
rect 11834 5728 11856 5760
rect 11888 5728 11910 5760
rect 11834 5692 11910 5728
rect 11834 5660 11856 5692
rect 11888 5660 11910 5692
rect 11834 5624 11910 5660
rect 11834 5592 11856 5624
rect 11888 5592 11910 5624
rect 11834 5556 11910 5592
rect 11834 5524 11856 5556
rect 11888 5524 11910 5556
rect 11834 5488 11910 5524
rect 11834 5456 11856 5488
rect 11888 5456 11910 5488
rect 11834 5420 11910 5456
rect 11834 5388 11856 5420
rect 11888 5388 11910 5420
rect 11834 5352 11910 5388
rect 11834 5320 11856 5352
rect 11888 5320 11910 5352
rect 11834 5282 11910 5320
rect 12010 6644 12086 6682
rect 12010 6612 12032 6644
rect 12064 6612 12086 6644
rect 12010 6576 12086 6612
rect 12010 6544 12032 6576
rect 12064 6544 12086 6576
rect 12010 6508 12086 6544
rect 12010 6476 12032 6508
rect 12064 6476 12086 6508
rect 12010 6440 12086 6476
rect 12010 6408 12032 6440
rect 12064 6408 12086 6440
rect 12010 6372 12086 6408
rect 12010 6340 12032 6372
rect 12064 6340 12086 6372
rect 12010 6304 12086 6340
rect 12010 6272 12032 6304
rect 12064 6272 12086 6304
rect 12010 6236 12086 6272
rect 12010 6204 12032 6236
rect 12064 6204 12086 6236
rect 12010 6168 12086 6204
rect 12010 6136 12032 6168
rect 12064 6136 12086 6168
rect 12010 6100 12086 6136
rect 12010 6068 12032 6100
rect 12064 6068 12086 6100
rect 12010 6032 12086 6068
rect 12010 6000 12032 6032
rect 12064 6000 12086 6032
rect 12010 5964 12086 6000
rect 12010 5932 12032 5964
rect 12064 5932 12086 5964
rect 12010 5896 12086 5932
rect 12010 5864 12032 5896
rect 12064 5864 12086 5896
rect 12010 5828 12086 5864
rect 12010 5796 12032 5828
rect 12064 5796 12086 5828
rect 12010 5760 12086 5796
rect 12010 5728 12032 5760
rect 12064 5728 12086 5760
rect 12010 5692 12086 5728
rect 12010 5660 12032 5692
rect 12064 5660 12086 5692
rect 12010 5624 12086 5660
rect 12010 5592 12032 5624
rect 12064 5592 12086 5624
rect 12010 5556 12086 5592
rect 12010 5524 12032 5556
rect 12064 5524 12086 5556
rect 12010 5488 12086 5524
rect 12010 5456 12032 5488
rect 12064 5456 12086 5488
rect 12010 5420 12086 5456
rect 12010 5388 12032 5420
rect 12064 5388 12086 5420
rect 12010 5352 12086 5388
rect 12010 5320 12032 5352
rect 12064 5320 12086 5352
rect 12010 5282 12086 5320
rect 12186 6644 12262 6682
rect 12186 6612 12208 6644
rect 12240 6612 12262 6644
rect 12186 6576 12262 6612
rect 12186 6544 12208 6576
rect 12240 6544 12262 6576
rect 12186 6508 12262 6544
rect 12186 6476 12208 6508
rect 12240 6476 12262 6508
rect 12186 6440 12262 6476
rect 12186 6408 12208 6440
rect 12240 6408 12262 6440
rect 12186 6372 12262 6408
rect 12186 6340 12208 6372
rect 12240 6340 12262 6372
rect 12186 6304 12262 6340
rect 12186 6272 12208 6304
rect 12240 6272 12262 6304
rect 12186 6236 12262 6272
rect 12186 6204 12208 6236
rect 12240 6204 12262 6236
rect 12186 6168 12262 6204
rect 12186 6136 12208 6168
rect 12240 6136 12262 6168
rect 12186 6100 12262 6136
rect 12186 6068 12208 6100
rect 12240 6068 12262 6100
rect 12186 6032 12262 6068
rect 12186 6000 12208 6032
rect 12240 6000 12262 6032
rect 12186 5964 12262 6000
rect 12186 5932 12208 5964
rect 12240 5932 12262 5964
rect 12186 5896 12262 5932
rect 12186 5864 12208 5896
rect 12240 5864 12262 5896
rect 12186 5828 12262 5864
rect 12186 5796 12208 5828
rect 12240 5796 12262 5828
rect 12186 5760 12262 5796
rect 12186 5728 12208 5760
rect 12240 5728 12262 5760
rect 12186 5692 12262 5728
rect 12186 5660 12208 5692
rect 12240 5660 12262 5692
rect 12186 5624 12262 5660
rect 12186 5592 12208 5624
rect 12240 5592 12262 5624
rect 12186 5556 12262 5592
rect 12186 5524 12208 5556
rect 12240 5524 12262 5556
rect 12186 5488 12262 5524
rect 12186 5456 12208 5488
rect 12240 5456 12262 5488
rect 12186 5420 12262 5456
rect 12186 5388 12208 5420
rect 12240 5388 12262 5420
rect 12186 5352 12262 5388
rect 12186 5320 12208 5352
rect 12240 5320 12262 5352
rect 12186 5282 12262 5320
rect 12362 6644 12430 6682
rect 12362 6612 12384 6644
rect 12416 6612 12430 6644
rect 12362 6576 12430 6612
rect 12362 6544 12384 6576
rect 12416 6544 12430 6576
rect 12362 6508 12430 6544
rect 12362 6476 12384 6508
rect 12416 6476 12430 6508
rect 12362 6440 12430 6476
rect 12362 6408 12384 6440
rect 12416 6408 12430 6440
rect 12362 6372 12430 6408
rect 12362 6340 12384 6372
rect 12416 6340 12430 6372
rect 12362 6304 12430 6340
rect 12362 6272 12384 6304
rect 12416 6272 12430 6304
rect 12362 6236 12430 6272
rect 12362 6204 12384 6236
rect 12416 6204 12430 6236
rect 12362 6168 12430 6204
rect 12362 6136 12384 6168
rect 12416 6136 12430 6168
rect 12362 6100 12430 6136
rect 12362 6068 12384 6100
rect 12416 6068 12430 6100
rect 12362 6032 12430 6068
rect 12362 6000 12384 6032
rect 12416 6000 12430 6032
rect 12362 5964 12430 6000
rect 12362 5932 12384 5964
rect 12416 5932 12430 5964
rect 12362 5896 12430 5932
rect 12362 5864 12384 5896
rect 12416 5864 12430 5896
rect 12362 5828 12430 5864
rect 12362 5796 12384 5828
rect 12416 5796 12430 5828
rect 12362 5760 12430 5796
rect 12362 5728 12384 5760
rect 12416 5728 12430 5760
rect 12362 5692 12430 5728
rect 12362 5660 12384 5692
rect 12416 5660 12430 5692
rect 12362 5624 12430 5660
rect 12362 5592 12384 5624
rect 12416 5592 12430 5624
rect 12362 5556 12430 5592
rect 12362 5524 12384 5556
rect 12416 5524 12430 5556
rect 12362 5488 12430 5524
rect 12362 5456 12384 5488
rect 12416 5456 12430 5488
rect 12362 5420 12430 5456
rect 12362 5388 12384 5420
rect 12416 5388 12430 5420
rect 12362 5352 12430 5388
rect 12362 5320 12384 5352
rect 12416 5320 12430 5352
rect 12362 5282 12430 5320
<< hvndiffc >>
rect 540 3992 572 4024
rect 540 3924 572 3956
rect 540 3856 572 3888
rect 540 3788 572 3820
rect 540 3720 572 3752
rect 540 3652 572 3684
rect 540 3584 572 3616
rect 540 3516 572 3548
rect 540 3448 572 3480
rect 540 3380 572 3412
rect 540 3312 572 3344
rect 540 3244 572 3276
rect 540 3176 572 3208
rect 540 3108 572 3140
rect 540 3040 572 3072
rect 540 2972 572 3004
rect 540 2904 572 2936
rect 540 2836 572 2868
rect 540 2768 572 2800
rect 540 2700 572 2732
rect 540 2632 572 2664
rect 540 2564 572 2596
rect 540 2496 572 2528
rect 540 2428 572 2460
rect 540 2360 572 2392
rect 540 2292 572 2324
rect 2516 3992 2548 4024
rect 2516 3924 2548 3956
rect 2516 3856 2548 3888
rect 2516 3788 2548 3820
rect 2516 3720 2548 3752
rect 2516 3652 2548 3684
rect 2516 3584 2548 3616
rect 2516 3516 2548 3548
rect 2516 3448 2548 3480
rect 2516 3380 2548 3412
rect 2516 3312 2548 3344
rect 2516 3244 2548 3276
rect 2516 3176 2548 3208
rect 2516 3108 2548 3140
rect 2516 3040 2548 3072
rect 2516 2972 2548 3004
rect 2516 2904 2548 2936
rect 2516 2836 2548 2868
rect 2516 2768 2548 2800
rect 2516 2700 2548 2732
rect 2516 2632 2548 2664
rect 2516 2564 2548 2596
rect 2516 2496 2548 2528
rect 2516 2428 2548 2460
rect 2516 2360 2548 2392
rect 2516 2292 2548 2324
rect 4492 3992 4524 4024
rect 4492 3924 4524 3956
rect 4492 3856 4524 3888
rect 4492 3788 4524 3820
rect 4492 3720 4524 3752
rect 4492 3652 4524 3684
rect 4492 3584 4524 3616
rect 4492 3516 4524 3548
rect 4492 3448 4524 3480
rect 4492 3380 4524 3412
rect 4492 3312 4524 3344
rect 4492 3244 4524 3276
rect 4492 3176 4524 3208
rect 4492 3108 4524 3140
rect 4492 3040 4524 3072
rect 4492 2972 4524 3004
rect 4492 2904 4524 2936
rect 4492 2836 4524 2868
rect 4492 2768 4524 2800
rect 4492 2700 4524 2732
rect 4492 2632 4524 2664
rect 4492 2564 4524 2596
rect 4492 2496 4524 2528
rect 4492 2428 4524 2460
rect 4492 2360 4524 2392
rect 4492 2292 4524 2324
rect 6468 3992 6500 4024
rect 6468 3924 6500 3956
rect 6468 3856 6500 3888
rect 6468 3788 6500 3820
rect 6468 3720 6500 3752
rect 6468 3652 6500 3684
rect 6468 3584 6500 3616
rect 6468 3516 6500 3548
rect 6468 3448 6500 3480
rect 6468 3380 6500 3412
rect 6468 3312 6500 3344
rect 6468 3244 6500 3276
rect 6468 3176 6500 3208
rect 6468 3108 6500 3140
rect 6468 3040 6500 3072
rect 6468 2972 6500 3004
rect 6468 2904 6500 2936
rect 6468 2836 6500 2868
rect 6468 2768 6500 2800
rect 6468 2700 6500 2732
rect 6468 2632 6500 2664
rect 6468 2564 6500 2596
rect 6468 2496 6500 2528
rect 6468 2428 6500 2460
rect 6468 2360 6500 2392
rect 6468 2292 6500 2324
rect 8444 3992 8476 4024
rect 8444 3924 8476 3956
rect 8444 3856 8476 3888
rect 8444 3788 8476 3820
rect 8444 3720 8476 3752
rect 8444 3652 8476 3684
rect 8444 3584 8476 3616
rect 8444 3516 8476 3548
rect 8444 3448 8476 3480
rect 8444 3380 8476 3412
rect 8444 3312 8476 3344
rect 8444 3244 8476 3276
rect 8444 3176 8476 3208
rect 8444 3108 8476 3140
rect 8444 3040 8476 3072
rect 8444 2972 8476 3004
rect 8444 2904 8476 2936
rect 8444 2836 8476 2868
rect 8444 2768 8476 2800
rect 8444 2700 8476 2732
rect 8444 2632 8476 2664
rect 8444 2564 8476 2596
rect 8444 2496 8476 2528
rect 8444 2428 8476 2460
rect 8444 2360 8476 2392
rect 8444 2292 8476 2324
rect 10420 3992 10452 4024
rect 10420 3924 10452 3956
rect 10420 3856 10452 3888
rect 10420 3788 10452 3820
rect 10420 3720 10452 3752
rect 10420 3652 10452 3684
rect 10420 3584 10452 3616
rect 10420 3516 10452 3548
rect 10420 3448 10452 3480
rect 10420 3380 10452 3412
rect 10420 3312 10452 3344
rect 10420 3244 10452 3276
rect 10420 3176 10452 3208
rect 10420 3108 10452 3140
rect 10420 3040 10452 3072
rect 10420 2972 10452 3004
rect 10420 2904 10452 2936
rect 10420 2836 10452 2868
rect 10420 2768 10452 2800
rect 10420 2700 10452 2732
rect 10420 2632 10452 2664
rect 10420 2564 10452 2596
rect 10420 2496 10452 2528
rect 10420 2428 10452 2460
rect 10420 2360 10452 2392
rect 10420 2292 10452 2324
rect 12396 3992 12428 4024
rect 12396 3924 12428 3956
rect 12396 3856 12428 3888
rect 12396 3788 12428 3820
rect 12396 3720 12428 3752
rect 12396 3652 12428 3684
rect 12396 3584 12428 3616
rect 12396 3516 12428 3548
rect 12396 3448 12428 3480
rect 12396 3380 12428 3412
rect 12396 3312 12428 3344
rect 12396 3244 12428 3276
rect 12396 3176 12428 3208
rect 12396 3108 12428 3140
rect 12396 3040 12428 3072
rect 12396 2972 12428 3004
rect 12396 2904 12428 2936
rect 12396 2836 12428 2868
rect 12396 2768 12428 2800
rect 12396 2700 12428 2732
rect 12396 2632 12428 2664
rect 12396 2564 12428 2596
rect 12396 2496 12428 2528
rect 12396 2428 12428 2460
rect 12396 2360 12428 2392
rect 12396 2292 12428 2324
rect 14372 3992 14404 4024
rect 14372 3924 14404 3956
rect 14372 3856 14404 3888
rect 14372 3788 14404 3820
rect 14372 3720 14404 3752
rect 14372 3652 14404 3684
rect 14372 3584 14404 3616
rect 14372 3516 14404 3548
rect 14372 3448 14404 3480
rect 14372 3380 14404 3412
rect 14372 3312 14404 3344
rect 14372 3244 14404 3276
rect 14372 3176 14404 3208
rect 14372 3108 14404 3140
rect 14372 3040 14404 3072
rect 14372 2972 14404 3004
rect 14372 2904 14404 2936
rect 14372 2836 14404 2868
rect 14372 2768 14404 2800
rect 14372 2700 14404 2732
rect 14372 2632 14404 2664
rect 14372 2564 14404 2596
rect 14372 2496 14404 2528
rect 14372 2428 14404 2460
rect 14372 2360 14404 2392
rect 14372 2292 14404 2324
rect 14548 3992 14580 4024
rect 14548 3924 14580 3956
rect 14548 3856 14580 3888
rect 14548 3788 14580 3820
rect 14548 3720 14580 3752
rect 14548 3652 14580 3684
rect 14548 3584 14580 3616
rect 14548 3516 14580 3548
rect 14548 3448 14580 3480
rect 14548 3380 14580 3412
rect 14548 3312 14580 3344
rect 14548 3244 14580 3276
rect 14548 3176 14580 3208
rect 14548 3108 14580 3140
rect 14548 3040 14580 3072
rect 14548 2972 14580 3004
rect 14548 2904 14580 2936
rect 14548 2836 14580 2868
rect 14548 2768 14580 2800
rect 14548 2700 14580 2732
rect 14548 2632 14580 2664
rect 14548 2564 14580 2596
rect 14548 2496 14580 2528
rect 14548 2428 14580 2460
rect 14548 2360 14580 2392
rect 14548 2292 14580 2324
rect 14724 3992 14756 4024
rect 14724 3924 14756 3956
rect 14724 3856 14756 3888
rect 14724 3788 14756 3820
rect 14724 3720 14756 3752
rect 14724 3652 14756 3684
rect 14724 3584 14756 3616
rect 14724 3516 14756 3548
rect 14724 3448 14756 3480
rect 14724 3380 14756 3412
rect 14724 3312 14756 3344
rect 14724 3244 14756 3276
rect 14724 3176 14756 3208
rect 14724 3108 14756 3140
rect 14724 3040 14756 3072
rect 14724 2972 14756 3004
rect 14724 2904 14756 2936
rect 14724 2836 14756 2868
rect 14724 2768 14756 2800
rect 14724 2700 14756 2732
rect 14724 2632 14756 2664
rect 14724 2564 14756 2596
rect 14724 2496 14756 2528
rect 14724 2428 14756 2460
rect 14724 2360 14756 2392
rect 14724 2292 14756 2324
rect 14900 3992 14932 4024
rect 14900 3924 14932 3956
rect 14900 3856 14932 3888
rect 14900 3788 14932 3820
rect 14900 3720 14932 3752
rect 14900 3652 14932 3684
rect 14900 3584 14932 3616
rect 14900 3516 14932 3548
rect 14900 3448 14932 3480
rect 14900 3380 14932 3412
rect 14900 3312 14932 3344
rect 14900 3244 14932 3276
rect 14900 3176 14932 3208
rect 14900 3108 14932 3140
rect 14900 3040 14932 3072
rect 14900 2972 14932 3004
rect 14900 2904 14932 2936
rect 14900 2836 14932 2868
rect 14900 2768 14932 2800
rect 14900 2700 14932 2732
rect 14900 2632 14932 2664
rect 14900 2564 14932 2596
rect 14900 2496 14932 2528
rect 14900 2428 14932 2460
rect 14900 2360 14932 2392
rect 14900 2292 14932 2324
rect 15076 3992 15108 4024
rect 15076 3924 15108 3956
rect 15076 3856 15108 3888
rect 15076 3788 15108 3820
rect 15076 3720 15108 3752
rect 15076 3652 15108 3684
rect 15076 3584 15108 3616
rect 15076 3516 15108 3548
rect 15076 3448 15108 3480
rect 15076 3380 15108 3412
rect 15076 3312 15108 3344
rect 15076 3244 15108 3276
rect 15076 3176 15108 3208
rect 15076 3108 15108 3140
rect 15076 3040 15108 3072
rect 15076 2972 15108 3004
rect 15076 2904 15108 2936
rect 15076 2836 15108 2868
rect 15076 2768 15108 2800
rect 15076 2700 15108 2732
rect 15076 2632 15108 2664
rect 15076 2564 15108 2596
rect 15076 2496 15108 2528
rect 15076 2428 15108 2460
rect 15076 2360 15108 2392
rect 15076 2292 15108 2324
rect 15252 3992 15284 4024
rect 15252 3924 15284 3956
rect 15252 3856 15284 3888
rect 15252 3788 15284 3820
rect 15252 3720 15284 3752
rect 15252 3652 15284 3684
rect 15252 3584 15284 3616
rect 15252 3516 15284 3548
rect 15252 3448 15284 3480
rect 15252 3380 15284 3412
rect 15252 3312 15284 3344
rect 15252 3244 15284 3276
rect 15252 3176 15284 3208
rect 15252 3108 15284 3140
rect 15252 3040 15284 3072
rect 15252 2972 15284 3004
rect 15252 2904 15284 2936
rect 15252 2836 15284 2868
rect 15252 2768 15284 2800
rect 15252 2700 15284 2732
rect 15252 2632 15284 2664
rect 15252 2564 15284 2596
rect 15252 2496 15284 2528
rect 15252 2428 15284 2460
rect 15252 2360 15284 2392
rect 15252 2292 15284 2324
rect 15428 3992 15460 4024
rect 15428 3924 15460 3956
rect 15428 3856 15460 3888
rect 15428 3788 15460 3820
rect 15428 3720 15460 3752
rect 15428 3652 15460 3684
rect 15428 3584 15460 3616
rect 15428 3516 15460 3548
rect 15428 3448 15460 3480
rect 15428 3380 15460 3412
rect 15428 3312 15460 3344
rect 15428 3244 15460 3276
rect 15428 3176 15460 3208
rect 15428 3108 15460 3140
rect 15428 3040 15460 3072
rect 15428 2972 15460 3004
rect 15428 2904 15460 2936
rect 15428 2836 15460 2868
rect 15428 2768 15460 2800
rect 15428 2700 15460 2732
rect 15428 2632 15460 2664
rect 15428 2564 15460 2596
rect 15428 2496 15460 2528
rect 15428 2428 15460 2460
rect 15428 2360 15460 2392
rect 15428 2292 15460 2324
rect 540 2142 572 2174
rect 540 2074 572 2106
rect 540 2006 572 2038
rect 540 1938 572 1970
rect 540 1870 572 1902
rect 540 1802 572 1834
rect 540 1734 572 1766
rect 540 1666 572 1698
rect 540 1598 572 1630
rect 540 1530 572 1562
rect 540 1462 572 1494
rect 540 1394 572 1426
rect 540 1326 572 1358
rect 540 1258 572 1290
rect 540 1190 572 1222
rect 540 1122 572 1154
rect 540 1054 572 1086
rect 540 986 572 1018
rect 540 918 572 950
rect 540 850 572 882
rect 540 782 572 814
rect 540 714 572 746
rect 540 646 572 678
rect 540 578 572 610
rect 540 510 572 542
rect 540 442 572 474
rect 2516 2142 2548 2174
rect 2516 2074 2548 2106
rect 2516 2006 2548 2038
rect 2516 1938 2548 1970
rect 2516 1870 2548 1902
rect 2516 1802 2548 1834
rect 2516 1734 2548 1766
rect 2516 1666 2548 1698
rect 2516 1598 2548 1630
rect 2516 1530 2548 1562
rect 2516 1462 2548 1494
rect 2516 1394 2548 1426
rect 2516 1326 2548 1358
rect 2516 1258 2548 1290
rect 2516 1190 2548 1222
rect 2516 1122 2548 1154
rect 2516 1054 2548 1086
rect 2516 986 2548 1018
rect 2516 918 2548 950
rect 2516 850 2548 882
rect 2516 782 2548 814
rect 2516 714 2548 746
rect 2516 646 2548 678
rect 2516 578 2548 610
rect 2516 510 2548 542
rect 2516 442 2548 474
rect 4492 2142 4524 2174
rect 4492 2074 4524 2106
rect 4492 2006 4524 2038
rect 4492 1938 4524 1970
rect 4492 1870 4524 1902
rect 4492 1802 4524 1834
rect 4492 1734 4524 1766
rect 4492 1666 4524 1698
rect 4492 1598 4524 1630
rect 4492 1530 4524 1562
rect 4492 1462 4524 1494
rect 4492 1394 4524 1426
rect 4492 1326 4524 1358
rect 4492 1258 4524 1290
rect 4492 1190 4524 1222
rect 4492 1122 4524 1154
rect 4492 1054 4524 1086
rect 4492 986 4524 1018
rect 4492 918 4524 950
rect 4492 850 4524 882
rect 4492 782 4524 814
rect 4492 714 4524 746
rect 4492 646 4524 678
rect 4492 578 4524 610
rect 4492 510 4524 542
rect 4492 442 4524 474
rect 6468 2142 6500 2174
rect 6468 2074 6500 2106
rect 6468 2006 6500 2038
rect 6468 1938 6500 1970
rect 6468 1870 6500 1902
rect 6468 1802 6500 1834
rect 6468 1734 6500 1766
rect 6468 1666 6500 1698
rect 6468 1598 6500 1630
rect 6468 1530 6500 1562
rect 6468 1462 6500 1494
rect 6468 1394 6500 1426
rect 6468 1326 6500 1358
rect 6468 1258 6500 1290
rect 6468 1190 6500 1222
rect 6468 1122 6500 1154
rect 6468 1054 6500 1086
rect 6468 986 6500 1018
rect 6468 918 6500 950
rect 6468 850 6500 882
rect 6468 782 6500 814
rect 6468 714 6500 746
rect 6468 646 6500 678
rect 6468 578 6500 610
rect 6468 510 6500 542
rect 6468 442 6500 474
rect 8444 2142 8476 2174
rect 8444 2074 8476 2106
rect 8444 2006 8476 2038
rect 8444 1938 8476 1970
rect 8444 1870 8476 1902
rect 8444 1802 8476 1834
rect 8444 1734 8476 1766
rect 8444 1666 8476 1698
rect 8444 1598 8476 1630
rect 8444 1530 8476 1562
rect 8444 1462 8476 1494
rect 8444 1394 8476 1426
rect 8444 1326 8476 1358
rect 8444 1258 8476 1290
rect 8444 1190 8476 1222
rect 8444 1122 8476 1154
rect 8444 1054 8476 1086
rect 8444 986 8476 1018
rect 8444 918 8476 950
rect 8444 850 8476 882
rect 8444 782 8476 814
rect 8444 714 8476 746
rect 8444 646 8476 678
rect 8444 578 8476 610
rect 8444 510 8476 542
rect 8444 442 8476 474
rect 10420 2142 10452 2174
rect 10420 2074 10452 2106
rect 10420 2006 10452 2038
rect 10420 1938 10452 1970
rect 10420 1870 10452 1902
rect 10420 1802 10452 1834
rect 10420 1734 10452 1766
rect 10420 1666 10452 1698
rect 10420 1598 10452 1630
rect 10420 1530 10452 1562
rect 10420 1462 10452 1494
rect 10420 1394 10452 1426
rect 10420 1326 10452 1358
rect 10420 1258 10452 1290
rect 10420 1190 10452 1222
rect 10420 1122 10452 1154
rect 10420 1054 10452 1086
rect 10420 986 10452 1018
rect 10420 918 10452 950
rect 10420 850 10452 882
rect 10420 782 10452 814
rect 10420 714 10452 746
rect 10420 646 10452 678
rect 10420 578 10452 610
rect 10420 510 10452 542
rect 10420 442 10452 474
rect 12396 2142 12428 2174
rect 12396 2074 12428 2106
rect 12396 2006 12428 2038
rect 12396 1938 12428 1970
rect 12396 1870 12428 1902
rect 12396 1802 12428 1834
rect 12396 1734 12428 1766
rect 12396 1666 12428 1698
rect 12396 1598 12428 1630
rect 12396 1530 12428 1562
rect 12396 1462 12428 1494
rect 12396 1394 12428 1426
rect 12396 1326 12428 1358
rect 12396 1258 12428 1290
rect 12396 1190 12428 1222
rect 12396 1122 12428 1154
rect 12396 1054 12428 1086
rect 12396 986 12428 1018
rect 12396 918 12428 950
rect 12396 850 12428 882
rect 12396 782 12428 814
rect 12396 714 12428 746
rect 12396 646 12428 678
rect 12396 578 12428 610
rect 12396 510 12428 542
rect 12396 442 12428 474
rect 14372 2142 14404 2174
rect 14372 2074 14404 2106
rect 14372 2006 14404 2038
rect 14372 1938 14404 1970
rect 14372 1870 14404 1902
rect 14372 1802 14404 1834
rect 14372 1734 14404 1766
rect 14372 1666 14404 1698
rect 14372 1598 14404 1630
rect 14372 1530 14404 1562
rect 14372 1462 14404 1494
rect 14372 1394 14404 1426
rect 14372 1326 14404 1358
rect 14372 1258 14404 1290
rect 14372 1190 14404 1222
rect 14372 1122 14404 1154
rect 14372 1054 14404 1086
rect 14372 986 14404 1018
rect 14372 918 14404 950
rect 14372 850 14404 882
rect 14372 782 14404 814
rect 14372 714 14404 746
rect 14372 646 14404 678
rect 14372 578 14404 610
rect 14372 510 14404 542
rect 14372 442 14404 474
rect 14548 2142 14580 2174
rect 14548 2074 14580 2106
rect 14548 2006 14580 2038
rect 14548 1938 14580 1970
rect 14548 1870 14580 1902
rect 14548 1802 14580 1834
rect 14548 1734 14580 1766
rect 14548 1666 14580 1698
rect 14548 1598 14580 1630
rect 14548 1530 14580 1562
rect 14548 1462 14580 1494
rect 14548 1394 14580 1426
rect 14548 1326 14580 1358
rect 14548 1258 14580 1290
rect 14548 1190 14580 1222
rect 14548 1122 14580 1154
rect 14548 1054 14580 1086
rect 14548 986 14580 1018
rect 14548 918 14580 950
rect 14548 850 14580 882
rect 14548 782 14580 814
rect 14548 714 14580 746
rect 14548 646 14580 678
rect 14548 578 14580 610
rect 14548 510 14580 542
rect 14548 442 14580 474
rect 14724 2142 14756 2174
rect 14724 2074 14756 2106
rect 14724 2006 14756 2038
rect 14724 1938 14756 1970
rect 14724 1870 14756 1902
rect 14724 1802 14756 1834
rect 14724 1734 14756 1766
rect 14724 1666 14756 1698
rect 14724 1598 14756 1630
rect 14724 1530 14756 1562
rect 14724 1462 14756 1494
rect 14724 1394 14756 1426
rect 14724 1326 14756 1358
rect 14724 1258 14756 1290
rect 14724 1190 14756 1222
rect 14724 1122 14756 1154
rect 14724 1054 14756 1086
rect 14724 986 14756 1018
rect 14724 918 14756 950
rect 14724 850 14756 882
rect 14724 782 14756 814
rect 14724 714 14756 746
rect 14724 646 14756 678
rect 14724 578 14756 610
rect 14724 510 14756 542
rect 14724 442 14756 474
rect 14900 2142 14932 2174
rect 14900 2074 14932 2106
rect 14900 2006 14932 2038
rect 14900 1938 14932 1970
rect 14900 1870 14932 1902
rect 14900 1802 14932 1834
rect 14900 1734 14932 1766
rect 14900 1666 14932 1698
rect 14900 1598 14932 1630
rect 14900 1530 14932 1562
rect 14900 1462 14932 1494
rect 14900 1394 14932 1426
rect 14900 1326 14932 1358
rect 14900 1258 14932 1290
rect 14900 1190 14932 1222
rect 14900 1122 14932 1154
rect 14900 1054 14932 1086
rect 14900 986 14932 1018
rect 14900 918 14932 950
rect 14900 850 14932 882
rect 14900 782 14932 814
rect 14900 714 14932 746
rect 14900 646 14932 678
rect 14900 578 14932 610
rect 14900 510 14932 542
rect 14900 442 14932 474
rect 15076 2142 15108 2174
rect 15076 2074 15108 2106
rect 15076 2006 15108 2038
rect 15076 1938 15108 1970
rect 15076 1870 15108 1902
rect 15076 1802 15108 1834
rect 15076 1734 15108 1766
rect 15076 1666 15108 1698
rect 15076 1598 15108 1630
rect 15076 1530 15108 1562
rect 15076 1462 15108 1494
rect 15076 1394 15108 1426
rect 15076 1326 15108 1358
rect 15076 1258 15108 1290
rect 15076 1190 15108 1222
rect 15076 1122 15108 1154
rect 15076 1054 15108 1086
rect 15076 986 15108 1018
rect 15076 918 15108 950
rect 15076 850 15108 882
rect 15076 782 15108 814
rect 15076 714 15108 746
rect 15076 646 15108 678
rect 15076 578 15108 610
rect 15076 510 15108 542
rect 15076 442 15108 474
rect 15252 2142 15284 2174
rect 15252 2074 15284 2106
rect 15252 2006 15284 2038
rect 15252 1938 15284 1970
rect 15252 1870 15284 1902
rect 15252 1802 15284 1834
rect 15252 1734 15284 1766
rect 15252 1666 15284 1698
rect 15252 1598 15284 1630
rect 15252 1530 15284 1562
rect 15252 1462 15284 1494
rect 15252 1394 15284 1426
rect 15252 1326 15284 1358
rect 15252 1258 15284 1290
rect 15252 1190 15284 1222
rect 15252 1122 15284 1154
rect 15252 1054 15284 1086
rect 15252 986 15284 1018
rect 15252 918 15284 950
rect 15252 850 15284 882
rect 15252 782 15284 814
rect 15252 714 15284 746
rect 15252 646 15284 678
rect 15252 578 15284 610
rect 15252 510 15284 542
rect 15252 442 15284 474
rect 15428 2142 15460 2174
rect 15428 2074 15460 2106
rect 15428 2006 15460 2038
rect 15428 1938 15460 1970
rect 15428 1870 15460 1902
rect 15428 1802 15460 1834
rect 15428 1734 15460 1766
rect 15428 1666 15460 1698
rect 15428 1598 15460 1630
rect 15428 1530 15460 1562
rect 15428 1462 15460 1494
rect 15428 1394 15460 1426
rect 15428 1326 15460 1358
rect 15428 1258 15460 1290
rect 15428 1190 15460 1222
rect 15428 1122 15460 1154
rect 15428 1054 15460 1086
rect 15428 986 15460 1018
rect 15428 918 15460 950
rect 15428 850 15460 882
rect 15428 782 15460 814
rect 15428 714 15460 746
rect 15428 646 15460 678
rect 15428 578 15460 610
rect 15428 510 15460 542
rect 15428 442 15460 474
<< hvpdiffc >>
rect 3584 6612 3616 6644
rect 3584 6544 3616 6576
rect 3584 6476 3616 6508
rect 3584 6408 3616 6440
rect 3584 6340 3616 6372
rect 3584 6272 3616 6304
rect 3584 6204 3616 6236
rect 3584 6136 3616 6168
rect 3584 6068 3616 6100
rect 3584 6000 3616 6032
rect 3584 5932 3616 5964
rect 3584 5864 3616 5896
rect 3584 5796 3616 5828
rect 3584 5728 3616 5760
rect 3584 5660 3616 5692
rect 3584 5592 3616 5624
rect 3584 5524 3616 5556
rect 3584 5456 3616 5488
rect 3584 5388 3616 5420
rect 3584 5320 3616 5352
rect 3760 6612 3792 6644
rect 3760 6544 3792 6576
rect 3760 6476 3792 6508
rect 3760 6408 3792 6440
rect 3760 6340 3792 6372
rect 3760 6272 3792 6304
rect 3760 6204 3792 6236
rect 3760 6136 3792 6168
rect 3760 6068 3792 6100
rect 3760 6000 3792 6032
rect 3760 5932 3792 5964
rect 3760 5864 3792 5896
rect 3760 5796 3792 5828
rect 3760 5728 3792 5760
rect 3760 5660 3792 5692
rect 3760 5592 3792 5624
rect 3760 5524 3792 5556
rect 3760 5456 3792 5488
rect 3760 5388 3792 5420
rect 3760 5320 3792 5352
rect 3936 6612 3968 6644
rect 3936 6544 3968 6576
rect 3936 6476 3968 6508
rect 3936 6408 3968 6440
rect 3936 6340 3968 6372
rect 3936 6272 3968 6304
rect 3936 6204 3968 6236
rect 3936 6136 3968 6168
rect 3936 6068 3968 6100
rect 3936 6000 3968 6032
rect 3936 5932 3968 5964
rect 3936 5864 3968 5896
rect 3936 5796 3968 5828
rect 3936 5728 3968 5760
rect 3936 5660 3968 5692
rect 3936 5592 3968 5624
rect 3936 5524 3968 5556
rect 3936 5456 3968 5488
rect 3936 5388 3968 5420
rect 3936 5320 3968 5352
rect 4112 6612 4144 6644
rect 4112 6544 4144 6576
rect 4112 6476 4144 6508
rect 4112 6408 4144 6440
rect 4112 6340 4144 6372
rect 4112 6272 4144 6304
rect 4112 6204 4144 6236
rect 4112 6136 4144 6168
rect 4112 6068 4144 6100
rect 4112 6000 4144 6032
rect 4112 5932 4144 5964
rect 4112 5864 4144 5896
rect 4112 5796 4144 5828
rect 4112 5728 4144 5760
rect 4112 5660 4144 5692
rect 4112 5592 4144 5624
rect 4112 5524 4144 5556
rect 4112 5456 4144 5488
rect 4112 5388 4144 5420
rect 4112 5320 4144 5352
rect 4288 6612 4320 6644
rect 4288 6544 4320 6576
rect 4288 6476 4320 6508
rect 4288 6408 4320 6440
rect 4288 6340 4320 6372
rect 4288 6272 4320 6304
rect 4288 6204 4320 6236
rect 4288 6136 4320 6168
rect 4288 6068 4320 6100
rect 4288 6000 4320 6032
rect 4288 5932 4320 5964
rect 4288 5864 4320 5896
rect 4288 5796 4320 5828
rect 4288 5728 4320 5760
rect 4288 5660 4320 5692
rect 4288 5592 4320 5624
rect 4288 5524 4320 5556
rect 4288 5456 4320 5488
rect 4288 5388 4320 5420
rect 4288 5320 4320 5352
rect 4464 6612 4496 6644
rect 4464 6544 4496 6576
rect 4464 6476 4496 6508
rect 4464 6408 4496 6440
rect 4464 6340 4496 6372
rect 4464 6272 4496 6304
rect 4464 6204 4496 6236
rect 4464 6136 4496 6168
rect 4464 6068 4496 6100
rect 4464 6000 4496 6032
rect 4464 5932 4496 5964
rect 4464 5864 4496 5896
rect 4464 5796 4496 5828
rect 4464 5728 4496 5760
rect 4464 5660 4496 5692
rect 4464 5592 4496 5624
rect 4464 5524 4496 5556
rect 4464 5456 4496 5488
rect 4464 5388 4496 5420
rect 4464 5320 4496 5352
rect 4640 6612 4672 6644
rect 4640 6544 4672 6576
rect 4640 6476 4672 6508
rect 4640 6408 4672 6440
rect 4640 6340 4672 6372
rect 4640 6272 4672 6304
rect 4640 6204 4672 6236
rect 4640 6136 4672 6168
rect 4640 6068 4672 6100
rect 4640 6000 4672 6032
rect 4640 5932 4672 5964
rect 4640 5864 4672 5896
rect 4640 5796 4672 5828
rect 4640 5728 4672 5760
rect 4640 5660 4672 5692
rect 4640 5592 4672 5624
rect 4640 5524 4672 5556
rect 4640 5456 4672 5488
rect 4640 5388 4672 5420
rect 4640 5320 4672 5352
rect 4816 6612 4848 6644
rect 4816 6544 4848 6576
rect 4816 6476 4848 6508
rect 4816 6408 4848 6440
rect 4816 6340 4848 6372
rect 4816 6272 4848 6304
rect 4816 6204 4848 6236
rect 4816 6136 4848 6168
rect 4816 6068 4848 6100
rect 4816 6000 4848 6032
rect 4816 5932 4848 5964
rect 4816 5864 4848 5896
rect 4816 5796 4848 5828
rect 4816 5728 4848 5760
rect 4816 5660 4848 5692
rect 4816 5592 4848 5624
rect 4816 5524 4848 5556
rect 4816 5456 4848 5488
rect 4816 5388 4848 5420
rect 4816 5320 4848 5352
rect 4992 6612 5024 6644
rect 4992 6544 5024 6576
rect 4992 6476 5024 6508
rect 4992 6408 5024 6440
rect 4992 6340 5024 6372
rect 4992 6272 5024 6304
rect 4992 6204 5024 6236
rect 4992 6136 5024 6168
rect 4992 6068 5024 6100
rect 4992 6000 5024 6032
rect 4992 5932 5024 5964
rect 4992 5864 5024 5896
rect 4992 5796 5024 5828
rect 4992 5728 5024 5760
rect 4992 5660 5024 5692
rect 4992 5592 5024 5624
rect 4992 5524 5024 5556
rect 4992 5456 5024 5488
rect 4992 5388 5024 5420
rect 4992 5320 5024 5352
rect 5168 6612 5200 6644
rect 5168 6544 5200 6576
rect 5168 6476 5200 6508
rect 5168 6408 5200 6440
rect 5168 6340 5200 6372
rect 5168 6272 5200 6304
rect 5168 6204 5200 6236
rect 5168 6136 5200 6168
rect 5168 6068 5200 6100
rect 5168 6000 5200 6032
rect 5168 5932 5200 5964
rect 5168 5864 5200 5896
rect 5168 5796 5200 5828
rect 5168 5728 5200 5760
rect 5168 5660 5200 5692
rect 5168 5592 5200 5624
rect 5168 5524 5200 5556
rect 5168 5456 5200 5488
rect 5168 5388 5200 5420
rect 5168 5320 5200 5352
rect 5344 6612 5376 6644
rect 5344 6544 5376 6576
rect 5344 6476 5376 6508
rect 5344 6408 5376 6440
rect 5344 6340 5376 6372
rect 5344 6272 5376 6304
rect 5344 6204 5376 6236
rect 5344 6136 5376 6168
rect 5344 6068 5376 6100
rect 5344 6000 5376 6032
rect 5344 5932 5376 5964
rect 5344 5864 5376 5896
rect 5344 5796 5376 5828
rect 5344 5728 5376 5760
rect 5344 5660 5376 5692
rect 5344 5592 5376 5624
rect 5344 5524 5376 5556
rect 5344 5456 5376 5488
rect 5344 5388 5376 5420
rect 5344 5320 5376 5352
rect 5520 6612 5552 6644
rect 5520 6544 5552 6576
rect 5520 6476 5552 6508
rect 5520 6408 5552 6440
rect 5520 6340 5552 6372
rect 5520 6272 5552 6304
rect 5520 6204 5552 6236
rect 5520 6136 5552 6168
rect 5520 6068 5552 6100
rect 5520 6000 5552 6032
rect 5520 5932 5552 5964
rect 5520 5864 5552 5896
rect 5520 5796 5552 5828
rect 5520 5728 5552 5760
rect 5520 5660 5552 5692
rect 5520 5592 5552 5624
rect 5520 5524 5552 5556
rect 5520 5456 5552 5488
rect 5520 5388 5552 5420
rect 5520 5320 5552 5352
rect 5696 6612 5728 6644
rect 5696 6544 5728 6576
rect 5696 6476 5728 6508
rect 5696 6408 5728 6440
rect 5696 6340 5728 6372
rect 5696 6272 5728 6304
rect 5696 6204 5728 6236
rect 5696 6136 5728 6168
rect 5696 6068 5728 6100
rect 5696 6000 5728 6032
rect 5696 5932 5728 5964
rect 5696 5864 5728 5896
rect 5696 5796 5728 5828
rect 5696 5728 5728 5760
rect 5696 5660 5728 5692
rect 5696 5592 5728 5624
rect 5696 5524 5728 5556
rect 5696 5456 5728 5488
rect 5696 5388 5728 5420
rect 5696 5320 5728 5352
rect 5872 6612 5904 6644
rect 5872 6544 5904 6576
rect 5872 6476 5904 6508
rect 5872 6408 5904 6440
rect 5872 6340 5904 6372
rect 5872 6272 5904 6304
rect 5872 6204 5904 6236
rect 5872 6136 5904 6168
rect 5872 6068 5904 6100
rect 5872 6000 5904 6032
rect 5872 5932 5904 5964
rect 5872 5864 5904 5896
rect 5872 5796 5904 5828
rect 5872 5728 5904 5760
rect 5872 5660 5904 5692
rect 5872 5592 5904 5624
rect 5872 5524 5904 5556
rect 5872 5456 5904 5488
rect 5872 5388 5904 5420
rect 5872 5320 5904 5352
rect 6048 6612 6080 6644
rect 6048 6544 6080 6576
rect 6048 6476 6080 6508
rect 6048 6408 6080 6440
rect 6048 6340 6080 6372
rect 6048 6272 6080 6304
rect 6048 6204 6080 6236
rect 6048 6136 6080 6168
rect 6048 6068 6080 6100
rect 6048 6000 6080 6032
rect 6048 5932 6080 5964
rect 6048 5864 6080 5896
rect 6048 5796 6080 5828
rect 6048 5728 6080 5760
rect 6048 5660 6080 5692
rect 6048 5592 6080 5624
rect 6048 5524 6080 5556
rect 6048 5456 6080 5488
rect 6048 5388 6080 5420
rect 6048 5320 6080 5352
rect 6224 6612 6256 6644
rect 6224 6544 6256 6576
rect 6224 6476 6256 6508
rect 6224 6408 6256 6440
rect 6224 6340 6256 6372
rect 6224 6272 6256 6304
rect 6224 6204 6256 6236
rect 6224 6136 6256 6168
rect 6224 6068 6256 6100
rect 6224 6000 6256 6032
rect 6224 5932 6256 5964
rect 6224 5864 6256 5896
rect 6224 5796 6256 5828
rect 6224 5728 6256 5760
rect 6224 5660 6256 5692
rect 6224 5592 6256 5624
rect 6224 5524 6256 5556
rect 6224 5456 6256 5488
rect 6224 5388 6256 5420
rect 6224 5320 6256 5352
rect 6400 6612 6432 6644
rect 6400 6544 6432 6576
rect 6400 6476 6432 6508
rect 6400 6408 6432 6440
rect 6400 6340 6432 6372
rect 6400 6272 6432 6304
rect 6400 6204 6432 6236
rect 6400 6136 6432 6168
rect 6400 6068 6432 6100
rect 6400 6000 6432 6032
rect 6400 5932 6432 5964
rect 6400 5864 6432 5896
rect 6400 5796 6432 5828
rect 6400 5728 6432 5760
rect 6400 5660 6432 5692
rect 6400 5592 6432 5624
rect 6400 5524 6432 5556
rect 6400 5456 6432 5488
rect 6400 5388 6432 5420
rect 6400 5320 6432 5352
rect 6576 6612 6608 6644
rect 6576 6544 6608 6576
rect 6576 6476 6608 6508
rect 6576 6408 6608 6440
rect 6576 6340 6608 6372
rect 6576 6272 6608 6304
rect 6576 6204 6608 6236
rect 6576 6136 6608 6168
rect 6576 6068 6608 6100
rect 6576 6000 6608 6032
rect 6576 5932 6608 5964
rect 6576 5864 6608 5896
rect 6576 5796 6608 5828
rect 6576 5728 6608 5760
rect 6576 5660 6608 5692
rect 6576 5592 6608 5624
rect 6576 5524 6608 5556
rect 6576 5456 6608 5488
rect 6576 5388 6608 5420
rect 6576 5320 6608 5352
rect 6752 6612 6784 6644
rect 6752 6544 6784 6576
rect 6752 6476 6784 6508
rect 6752 6408 6784 6440
rect 6752 6340 6784 6372
rect 6752 6272 6784 6304
rect 6752 6204 6784 6236
rect 6752 6136 6784 6168
rect 6752 6068 6784 6100
rect 6752 6000 6784 6032
rect 6752 5932 6784 5964
rect 6752 5864 6784 5896
rect 6752 5796 6784 5828
rect 6752 5728 6784 5760
rect 6752 5660 6784 5692
rect 6752 5592 6784 5624
rect 6752 5524 6784 5556
rect 6752 5456 6784 5488
rect 6752 5388 6784 5420
rect 6752 5320 6784 5352
rect 6928 6612 6960 6644
rect 6928 6544 6960 6576
rect 6928 6476 6960 6508
rect 6928 6408 6960 6440
rect 6928 6340 6960 6372
rect 6928 6272 6960 6304
rect 6928 6204 6960 6236
rect 6928 6136 6960 6168
rect 6928 6068 6960 6100
rect 6928 6000 6960 6032
rect 6928 5932 6960 5964
rect 6928 5864 6960 5896
rect 6928 5796 6960 5828
rect 6928 5728 6960 5760
rect 6928 5660 6960 5692
rect 6928 5592 6960 5624
rect 6928 5524 6960 5556
rect 6928 5456 6960 5488
rect 6928 5388 6960 5420
rect 6928 5320 6960 5352
rect 7104 6612 7136 6644
rect 7104 6544 7136 6576
rect 7104 6476 7136 6508
rect 7104 6408 7136 6440
rect 7104 6340 7136 6372
rect 7104 6272 7136 6304
rect 7104 6204 7136 6236
rect 7104 6136 7136 6168
rect 7104 6068 7136 6100
rect 7104 6000 7136 6032
rect 7104 5932 7136 5964
rect 7104 5864 7136 5896
rect 7104 5796 7136 5828
rect 7104 5728 7136 5760
rect 7104 5660 7136 5692
rect 7104 5592 7136 5624
rect 7104 5524 7136 5556
rect 7104 5456 7136 5488
rect 7104 5388 7136 5420
rect 7104 5320 7136 5352
rect 7280 6612 7312 6644
rect 7280 6544 7312 6576
rect 7280 6476 7312 6508
rect 7280 6408 7312 6440
rect 7280 6340 7312 6372
rect 7280 6272 7312 6304
rect 7280 6204 7312 6236
rect 7280 6136 7312 6168
rect 7280 6068 7312 6100
rect 7280 6000 7312 6032
rect 7280 5932 7312 5964
rect 7280 5864 7312 5896
rect 7280 5796 7312 5828
rect 7280 5728 7312 5760
rect 7280 5660 7312 5692
rect 7280 5592 7312 5624
rect 7280 5524 7312 5556
rect 7280 5456 7312 5488
rect 7280 5388 7312 5420
rect 7280 5320 7312 5352
rect 7456 6612 7488 6644
rect 7456 6544 7488 6576
rect 7456 6476 7488 6508
rect 7456 6408 7488 6440
rect 7456 6340 7488 6372
rect 7456 6272 7488 6304
rect 7456 6204 7488 6236
rect 7456 6136 7488 6168
rect 7456 6068 7488 6100
rect 7456 6000 7488 6032
rect 7456 5932 7488 5964
rect 7456 5864 7488 5896
rect 7456 5796 7488 5828
rect 7456 5728 7488 5760
rect 7456 5660 7488 5692
rect 7456 5592 7488 5624
rect 7456 5524 7488 5556
rect 7456 5456 7488 5488
rect 7456 5388 7488 5420
rect 7456 5320 7488 5352
rect 7632 6612 7664 6644
rect 7632 6544 7664 6576
rect 7632 6476 7664 6508
rect 7632 6408 7664 6440
rect 7632 6340 7664 6372
rect 7632 6272 7664 6304
rect 7632 6204 7664 6236
rect 7632 6136 7664 6168
rect 7632 6068 7664 6100
rect 7632 6000 7664 6032
rect 7632 5932 7664 5964
rect 7632 5864 7664 5896
rect 7632 5796 7664 5828
rect 7632 5728 7664 5760
rect 7632 5660 7664 5692
rect 7632 5592 7664 5624
rect 7632 5524 7664 5556
rect 7632 5456 7664 5488
rect 7632 5388 7664 5420
rect 7632 5320 7664 5352
rect 7808 6612 7840 6644
rect 7808 6544 7840 6576
rect 7808 6476 7840 6508
rect 7808 6408 7840 6440
rect 7808 6340 7840 6372
rect 7808 6272 7840 6304
rect 7808 6204 7840 6236
rect 7808 6136 7840 6168
rect 7808 6068 7840 6100
rect 7808 6000 7840 6032
rect 7808 5932 7840 5964
rect 7808 5864 7840 5896
rect 7808 5796 7840 5828
rect 7808 5728 7840 5760
rect 7808 5660 7840 5692
rect 7808 5592 7840 5624
rect 7808 5524 7840 5556
rect 7808 5456 7840 5488
rect 7808 5388 7840 5420
rect 7808 5320 7840 5352
rect 7984 6612 8016 6644
rect 7984 6544 8016 6576
rect 7984 6476 8016 6508
rect 7984 6408 8016 6440
rect 7984 6340 8016 6372
rect 7984 6272 8016 6304
rect 7984 6204 8016 6236
rect 7984 6136 8016 6168
rect 7984 6068 8016 6100
rect 7984 6000 8016 6032
rect 7984 5932 8016 5964
rect 7984 5864 8016 5896
rect 7984 5796 8016 5828
rect 7984 5728 8016 5760
rect 7984 5660 8016 5692
rect 7984 5592 8016 5624
rect 7984 5524 8016 5556
rect 7984 5456 8016 5488
rect 7984 5388 8016 5420
rect 7984 5320 8016 5352
rect 8160 6612 8192 6644
rect 8160 6544 8192 6576
rect 8160 6476 8192 6508
rect 8160 6408 8192 6440
rect 8160 6340 8192 6372
rect 8160 6272 8192 6304
rect 8160 6204 8192 6236
rect 8160 6136 8192 6168
rect 8160 6068 8192 6100
rect 8160 6000 8192 6032
rect 8160 5932 8192 5964
rect 8160 5864 8192 5896
rect 8160 5796 8192 5828
rect 8160 5728 8192 5760
rect 8160 5660 8192 5692
rect 8160 5592 8192 5624
rect 8160 5524 8192 5556
rect 8160 5456 8192 5488
rect 8160 5388 8192 5420
rect 8160 5320 8192 5352
rect 8336 6612 8368 6644
rect 8336 6544 8368 6576
rect 8336 6476 8368 6508
rect 8336 6408 8368 6440
rect 8336 6340 8368 6372
rect 8336 6272 8368 6304
rect 8336 6204 8368 6236
rect 8336 6136 8368 6168
rect 8336 6068 8368 6100
rect 8336 6000 8368 6032
rect 8336 5932 8368 5964
rect 8336 5864 8368 5896
rect 8336 5796 8368 5828
rect 8336 5728 8368 5760
rect 8336 5660 8368 5692
rect 8336 5592 8368 5624
rect 8336 5524 8368 5556
rect 8336 5456 8368 5488
rect 8336 5388 8368 5420
rect 8336 5320 8368 5352
rect 8512 6612 8544 6644
rect 8512 6544 8544 6576
rect 8512 6476 8544 6508
rect 8512 6408 8544 6440
rect 8512 6340 8544 6372
rect 8512 6272 8544 6304
rect 8512 6204 8544 6236
rect 8512 6136 8544 6168
rect 8512 6068 8544 6100
rect 8512 6000 8544 6032
rect 8512 5932 8544 5964
rect 8512 5864 8544 5896
rect 8512 5796 8544 5828
rect 8512 5728 8544 5760
rect 8512 5660 8544 5692
rect 8512 5592 8544 5624
rect 8512 5524 8544 5556
rect 8512 5456 8544 5488
rect 8512 5388 8544 5420
rect 8512 5320 8544 5352
rect 8688 6612 8720 6644
rect 8688 6544 8720 6576
rect 8688 6476 8720 6508
rect 8688 6408 8720 6440
rect 8688 6340 8720 6372
rect 8688 6272 8720 6304
rect 8688 6204 8720 6236
rect 8688 6136 8720 6168
rect 8688 6068 8720 6100
rect 8688 6000 8720 6032
rect 8688 5932 8720 5964
rect 8688 5864 8720 5896
rect 8688 5796 8720 5828
rect 8688 5728 8720 5760
rect 8688 5660 8720 5692
rect 8688 5592 8720 5624
rect 8688 5524 8720 5556
rect 8688 5456 8720 5488
rect 8688 5388 8720 5420
rect 8688 5320 8720 5352
rect 8864 6612 8896 6644
rect 8864 6544 8896 6576
rect 8864 6476 8896 6508
rect 8864 6408 8896 6440
rect 8864 6340 8896 6372
rect 8864 6272 8896 6304
rect 8864 6204 8896 6236
rect 8864 6136 8896 6168
rect 8864 6068 8896 6100
rect 8864 6000 8896 6032
rect 8864 5932 8896 5964
rect 8864 5864 8896 5896
rect 8864 5796 8896 5828
rect 8864 5728 8896 5760
rect 8864 5660 8896 5692
rect 8864 5592 8896 5624
rect 8864 5524 8896 5556
rect 8864 5456 8896 5488
rect 8864 5388 8896 5420
rect 8864 5320 8896 5352
rect 9040 6612 9072 6644
rect 9040 6544 9072 6576
rect 9040 6476 9072 6508
rect 9040 6408 9072 6440
rect 9040 6340 9072 6372
rect 9040 6272 9072 6304
rect 9040 6204 9072 6236
rect 9040 6136 9072 6168
rect 9040 6068 9072 6100
rect 9040 6000 9072 6032
rect 9040 5932 9072 5964
rect 9040 5864 9072 5896
rect 9040 5796 9072 5828
rect 9040 5728 9072 5760
rect 9040 5660 9072 5692
rect 9040 5592 9072 5624
rect 9040 5524 9072 5556
rect 9040 5456 9072 5488
rect 9040 5388 9072 5420
rect 9040 5320 9072 5352
rect 9216 6612 9248 6644
rect 9216 6544 9248 6576
rect 9216 6476 9248 6508
rect 9216 6408 9248 6440
rect 9216 6340 9248 6372
rect 9216 6272 9248 6304
rect 9216 6204 9248 6236
rect 9216 6136 9248 6168
rect 9216 6068 9248 6100
rect 9216 6000 9248 6032
rect 9216 5932 9248 5964
rect 9216 5864 9248 5896
rect 9216 5796 9248 5828
rect 9216 5728 9248 5760
rect 9216 5660 9248 5692
rect 9216 5592 9248 5624
rect 9216 5524 9248 5556
rect 9216 5456 9248 5488
rect 9216 5388 9248 5420
rect 9216 5320 9248 5352
rect 9392 6612 9424 6644
rect 9392 6544 9424 6576
rect 9392 6476 9424 6508
rect 9392 6408 9424 6440
rect 9392 6340 9424 6372
rect 9392 6272 9424 6304
rect 9392 6204 9424 6236
rect 9392 6136 9424 6168
rect 9392 6068 9424 6100
rect 9392 6000 9424 6032
rect 9392 5932 9424 5964
rect 9392 5864 9424 5896
rect 9392 5796 9424 5828
rect 9392 5728 9424 5760
rect 9392 5660 9424 5692
rect 9392 5592 9424 5624
rect 9392 5524 9424 5556
rect 9392 5456 9424 5488
rect 9392 5388 9424 5420
rect 9392 5320 9424 5352
rect 9568 6612 9600 6644
rect 9568 6544 9600 6576
rect 9568 6476 9600 6508
rect 9568 6408 9600 6440
rect 9568 6340 9600 6372
rect 9568 6272 9600 6304
rect 9568 6204 9600 6236
rect 9568 6136 9600 6168
rect 9568 6068 9600 6100
rect 9568 6000 9600 6032
rect 9568 5932 9600 5964
rect 9568 5864 9600 5896
rect 9568 5796 9600 5828
rect 9568 5728 9600 5760
rect 9568 5660 9600 5692
rect 9568 5592 9600 5624
rect 9568 5524 9600 5556
rect 9568 5456 9600 5488
rect 9568 5388 9600 5420
rect 9568 5320 9600 5352
rect 9744 6612 9776 6644
rect 9744 6544 9776 6576
rect 9744 6476 9776 6508
rect 9744 6408 9776 6440
rect 9744 6340 9776 6372
rect 9744 6272 9776 6304
rect 9744 6204 9776 6236
rect 9744 6136 9776 6168
rect 9744 6068 9776 6100
rect 9744 6000 9776 6032
rect 9744 5932 9776 5964
rect 9744 5864 9776 5896
rect 9744 5796 9776 5828
rect 9744 5728 9776 5760
rect 9744 5660 9776 5692
rect 9744 5592 9776 5624
rect 9744 5524 9776 5556
rect 9744 5456 9776 5488
rect 9744 5388 9776 5420
rect 9744 5320 9776 5352
rect 9920 6612 9952 6644
rect 9920 6544 9952 6576
rect 9920 6476 9952 6508
rect 9920 6408 9952 6440
rect 9920 6340 9952 6372
rect 9920 6272 9952 6304
rect 9920 6204 9952 6236
rect 9920 6136 9952 6168
rect 9920 6068 9952 6100
rect 9920 6000 9952 6032
rect 9920 5932 9952 5964
rect 9920 5864 9952 5896
rect 9920 5796 9952 5828
rect 9920 5728 9952 5760
rect 9920 5660 9952 5692
rect 9920 5592 9952 5624
rect 9920 5524 9952 5556
rect 9920 5456 9952 5488
rect 9920 5388 9952 5420
rect 9920 5320 9952 5352
rect 10096 6612 10128 6644
rect 10096 6544 10128 6576
rect 10096 6476 10128 6508
rect 10096 6408 10128 6440
rect 10096 6340 10128 6372
rect 10096 6272 10128 6304
rect 10096 6204 10128 6236
rect 10096 6136 10128 6168
rect 10096 6068 10128 6100
rect 10096 6000 10128 6032
rect 10096 5932 10128 5964
rect 10096 5864 10128 5896
rect 10096 5796 10128 5828
rect 10096 5728 10128 5760
rect 10096 5660 10128 5692
rect 10096 5592 10128 5624
rect 10096 5524 10128 5556
rect 10096 5456 10128 5488
rect 10096 5388 10128 5420
rect 10096 5320 10128 5352
rect 10272 6612 10304 6644
rect 10272 6544 10304 6576
rect 10272 6476 10304 6508
rect 10272 6408 10304 6440
rect 10272 6340 10304 6372
rect 10272 6272 10304 6304
rect 10272 6204 10304 6236
rect 10272 6136 10304 6168
rect 10272 6068 10304 6100
rect 10272 6000 10304 6032
rect 10272 5932 10304 5964
rect 10272 5864 10304 5896
rect 10272 5796 10304 5828
rect 10272 5728 10304 5760
rect 10272 5660 10304 5692
rect 10272 5592 10304 5624
rect 10272 5524 10304 5556
rect 10272 5456 10304 5488
rect 10272 5388 10304 5420
rect 10272 5320 10304 5352
rect 10448 6612 10480 6644
rect 10448 6544 10480 6576
rect 10448 6476 10480 6508
rect 10448 6408 10480 6440
rect 10448 6340 10480 6372
rect 10448 6272 10480 6304
rect 10448 6204 10480 6236
rect 10448 6136 10480 6168
rect 10448 6068 10480 6100
rect 10448 6000 10480 6032
rect 10448 5932 10480 5964
rect 10448 5864 10480 5896
rect 10448 5796 10480 5828
rect 10448 5728 10480 5760
rect 10448 5660 10480 5692
rect 10448 5592 10480 5624
rect 10448 5524 10480 5556
rect 10448 5456 10480 5488
rect 10448 5388 10480 5420
rect 10448 5320 10480 5352
rect 10624 6612 10656 6644
rect 10624 6544 10656 6576
rect 10624 6476 10656 6508
rect 10624 6408 10656 6440
rect 10624 6340 10656 6372
rect 10624 6272 10656 6304
rect 10624 6204 10656 6236
rect 10624 6136 10656 6168
rect 10624 6068 10656 6100
rect 10624 6000 10656 6032
rect 10624 5932 10656 5964
rect 10624 5864 10656 5896
rect 10624 5796 10656 5828
rect 10624 5728 10656 5760
rect 10624 5660 10656 5692
rect 10624 5592 10656 5624
rect 10624 5524 10656 5556
rect 10624 5456 10656 5488
rect 10624 5388 10656 5420
rect 10624 5320 10656 5352
rect 10800 6612 10832 6644
rect 10800 6544 10832 6576
rect 10800 6476 10832 6508
rect 10800 6408 10832 6440
rect 10800 6340 10832 6372
rect 10800 6272 10832 6304
rect 10800 6204 10832 6236
rect 10800 6136 10832 6168
rect 10800 6068 10832 6100
rect 10800 6000 10832 6032
rect 10800 5932 10832 5964
rect 10800 5864 10832 5896
rect 10800 5796 10832 5828
rect 10800 5728 10832 5760
rect 10800 5660 10832 5692
rect 10800 5592 10832 5624
rect 10800 5524 10832 5556
rect 10800 5456 10832 5488
rect 10800 5388 10832 5420
rect 10800 5320 10832 5352
rect 10976 6612 11008 6644
rect 10976 6544 11008 6576
rect 10976 6476 11008 6508
rect 10976 6408 11008 6440
rect 10976 6340 11008 6372
rect 10976 6272 11008 6304
rect 10976 6204 11008 6236
rect 10976 6136 11008 6168
rect 10976 6068 11008 6100
rect 10976 6000 11008 6032
rect 10976 5932 11008 5964
rect 10976 5864 11008 5896
rect 10976 5796 11008 5828
rect 10976 5728 11008 5760
rect 10976 5660 11008 5692
rect 10976 5592 11008 5624
rect 10976 5524 11008 5556
rect 10976 5456 11008 5488
rect 10976 5388 11008 5420
rect 10976 5320 11008 5352
rect 11152 6612 11184 6644
rect 11152 6544 11184 6576
rect 11152 6476 11184 6508
rect 11152 6408 11184 6440
rect 11152 6340 11184 6372
rect 11152 6272 11184 6304
rect 11152 6204 11184 6236
rect 11152 6136 11184 6168
rect 11152 6068 11184 6100
rect 11152 6000 11184 6032
rect 11152 5932 11184 5964
rect 11152 5864 11184 5896
rect 11152 5796 11184 5828
rect 11152 5728 11184 5760
rect 11152 5660 11184 5692
rect 11152 5592 11184 5624
rect 11152 5524 11184 5556
rect 11152 5456 11184 5488
rect 11152 5388 11184 5420
rect 11152 5320 11184 5352
rect 11328 6612 11360 6644
rect 11328 6544 11360 6576
rect 11328 6476 11360 6508
rect 11328 6408 11360 6440
rect 11328 6340 11360 6372
rect 11328 6272 11360 6304
rect 11328 6204 11360 6236
rect 11328 6136 11360 6168
rect 11328 6068 11360 6100
rect 11328 6000 11360 6032
rect 11328 5932 11360 5964
rect 11328 5864 11360 5896
rect 11328 5796 11360 5828
rect 11328 5728 11360 5760
rect 11328 5660 11360 5692
rect 11328 5592 11360 5624
rect 11328 5524 11360 5556
rect 11328 5456 11360 5488
rect 11328 5388 11360 5420
rect 11328 5320 11360 5352
rect 11504 6612 11536 6644
rect 11504 6544 11536 6576
rect 11504 6476 11536 6508
rect 11504 6408 11536 6440
rect 11504 6340 11536 6372
rect 11504 6272 11536 6304
rect 11504 6204 11536 6236
rect 11504 6136 11536 6168
rect 11504 6068 11536 6100
rect 11504 6000 11536 6032
rect 11504 5932 11536 5964
rect 11504 5864 11536 5896
rect 11504 5796 11536 5828
rect 11504 5728 11536 5760
rect 11504 5660 11536 5692
rect 11504 5592 11536 5624
rect 11504 5524 11536 5556
rect 11504 5456 11536 5488
rect 11504 5388 11536 5420
rect 11504 5320 11536 5352
rect 11680 6612 11712 6644
rect 11680 6544 11712 6576
rect 11680 6476 11712 6508
rect 11680 6408 11712 6440
rect 11680 6340 11712 6372
rect 11680 6272 11712 6304
rect 11680 6204 11712 6236
rect 11680 6136 11712 6168
rect 11680 6068 11712 6100
rect 11680 6000 11712 6032
rect 11680 5932 11712 5964
rect 11680 5864 11712 5896
rect 11680 5796 11712 5828
rect 11680 5728 11712 5760
rect 11680 5660 11712 5692
rect 11680 5592 11712 5624
rect 11680 5524 11712 5556
rect 11680 5456 11712 5488
rect 11680 5388 11712 5420
rect 11680 5320 11712 5352
rect 11856 6612 11888 6644
rect 11856 6544 11888 6576
rect 11856 6476 11888 6508
rect 11856 6408 11888 6440
rect 11856 6340 11888 6372
rect 11856 6272 11888 6304
rect 11856 6204 11888 6236
rect 11856 6136 11888 6168
rect 11856 6068 11888 6100
rect 11856 6000 11888 6032
rect 11856 5932 11888 5964
rect 11856 5864 11888 5896
rect 11856 5796 11888 5828
rect 11856 5728 11888 5760
rect 11856 5660 11888 5692
rect 11856 5592 11888 5624
rect 11856 5524 11888 5556
rect 11856 5456 11888 5488
rect 11856 5388 11888 5420
rect 11856 5320 11888 5352
rect 12032 6612 12064 6644
rect 12032 6544 12064 6576
rect 12032 6476 12064 6508
rect 12032 6408 12064 6440
rect 12032 6340 12064 6372
rect 12032 6272 12064 6304
rect 12032 6204 12064 6236
rect 12032 6136 12064 6168
rect 12032 6068 12064 6100
rect 12032 6000 12064 6032
rect 12032 5932 12064 5964
rect 12032 5864 12064 5896
rect 12032 5796 12064 5828
rect 12032 5728 12064 5760
rect 12032 5660 12064 5692
rect 12032 5592 12064 5624
rect 12032 5524 12064 5556
rect 12032 5456 12064 5488
rect 12032 5388 12064 5420
rect 12032 5320 12064 5352
rect 12208 6612 12240 6644
rect 12208 6544 12240 6576
rect 12208 6476 12240 6508
rect 12208 6408 12240 6440
rect 12208 6340 12240 6372
rect 12208 6272 12240 6304
rect 12208 6204 12240 6236
rect 12208 6136 12240 6168
rect 12208 6068 12240 6100
rect 12208 6000 12240 6032
rect 12208 5932 12240 5964
rect 12208 5864 12240 5896
rect 12208 5796 12240 5828
rect 12208 5728 12240 5760
rect 12208 5660 12240 5692
rect 12208 5592 12240 5624
rect 12208 5524 12240 5556
rect 12208 5456 12240 5488
rect 12208 5388 12240 5420
rect 12208 5320 12240 5352
rect 12384 6612 12416 6644
rect 12384 6544 12416 6576
rect 12384 6476 12416 6508
rect 12384 6408 12416 6440
rect 12384 6340 12416 6372
rect 12384 6272 12416 6304
rect 12384 6204 12416 6236
rect 12384 6136 12416 6168
rect 12384 6068 12416 6100
rect 12384 6000 12416 6032
rect 12384 5932 12416 5964
rect 12384 5864 12416 5896
rect 12384 5796 12416 5828
rect 12384 5728 12416 5760
rect 12384 5660 12416 5692
rect 12384 5592 12416 5624
rect 12384 5524 12416 5556
rect 12384 5456 12416 5488
rect 12384 5388 12416 5420
rect 12384 5320 12416 5352
<< psubdiff >>
rect 0 4448 16000 4466
rect 0 4416 28 4448
rect 60 4416 96 4448
rect 128 4416 164 4448
rect 196 4416 232 4448
rect 264 4416 300 4448
rect 332 4416 368 4448
rect 400 4416 436 4448
rect 468 4416 504 4448
rect 536 4416 572 4448
rect 604 4416 640 4448
rect 672 4416 708 4448
rect 740 4416 776 4448
rect 808 4416 844 4448
rect 876 4416 912 4448
rect 944 4416 980 4448
rect 1012 4416 1048 4448
rect 1080 4416 1116 4448
rect 1148 4416 1184 4448
rect 1216 4416 1252 4448
rect 1284 4416 1320 4448
rect 1352 4416 1388 4448
rect 1420 4416 1456 4448
rect 1488 4416 1524 4448
rect 1556 4416 1592 4448
rect 1624 4416 1660 4448
rect 1692 4416 1728 4448
rect 1760 4416 1796 4448
rect 1828 4416 1864 4448
rect 1896 4416 1932 4448
rect 1964 4416 2000 4448
rect 2032 4416 2068 4448
rect 2100 4416 2136 4448
rect 2168 4416 2204 4448
rect 2236 4416 2272 4448
rect 2304 4416 2340 4448
rect 2372 4416 2408 4448
rect 2440 4416 2476 4448
rect 2508 4416 2544 4448
rect 2576 4416 2612 4448
rect 2644 4416 2680 4448
rect 2712 4416 2748 4448
rect 2780 4416 2816 4448
rect 2848 4416 2884 4448
rect 2916 4416 2952 4448
rect 2984 4416 3020 4448
rect 3052 4416 3088 4448
rect 3120 4416 3156 4448
rect 3188 4416 3224 4448
rect 3256 4416 3292 4448
rect 3324 4416 3360 4448
rect 3392 4416 3428 4448
rect 3460 4416 3496 4448
rect 3528 4416 3564 4448
rect 3596 4416 3632 4448
rect 3664 4416 3700 4448
rect 3732 4416 3768 4448
rect 3800 4416 3836 4448
rect 3868 4416 3904 4448
rect 3936 4416 3972 4448
rect 4004 4416 4040 4448
rect 4072 4416 4108 4448
rect 4140 4416 4176 4448
rect 4208 4416 4244 4448
rect 4276 4416 4312 4448
rect 4344 4416 4380 4448
rect 4412 4416 4448 4448
rect 4480 4416 4516 4448
rect 4548 4416 4584 4448
rect 4616 4416 4652 4448
rect 4684 4416 4720 4448
rect 4752 4416 4788 4448
rect 4820 4416 4856 4448
rect 4888 4416 4924 4448
rect 4956 4416 4992 4448
rect 5024 4416 5060 4448
rect 5092 4416 5128 4448
rect 5160 4416 5196 4448
rect 5228 4416 5264 4448
rect 5296 4416 5332 4448
rect 5364 4416 5400 4448
rect 5432 4416 5468 4448
rect 5500 4416 5536 4448
rect 5568 4416 5604 4448
rect 5636 4416 5672 4448
rect 5704 4416 5740 4448
rect 5772 4416 5808 4448
rect 5840 4416 5876 4448
rect 5908 4416 5944 4448
rect 5976 4416 6012 4448
rect 6044 4416 6080 4448
rect 6112 4416 6148 4448
rect 6180 4416 6216 4448
rect 6248 4416 6284 4448
rect 6316 4416 6352 4448
rect 6384 4416 6420 4448
rect 6452 4416 6488 4448
rect 6520 4416 6556 4448
rect 6588 4416 6624 4448
rect 6656 4416 6692 4448
rect 6724 4416 6760 4448
rect 6792 4416 6828 4448
rect 6860 4416 6896 4448
rect 6928 4416 6964 4448
rect 6996 4416 7032 4448
rect 7064 4416 7100 4448
rect 7132 4416 7168 4448
rect 7200 4416 7236 4448
rect 7268 4416 7304 4448
rect 7336 4416 7372 4448
rect 7404 4416 7440 4448
rect 7472 4416 7508 4448
rect 7540 4416 7576 4448
rect 7608 4416 7644 4448
rect 7676 4416 7712 4448
rect 7744 4416 7780 4448
rect 7812 4416 7848 4448
rect 7880 4416 7916 4448
rect 7948 4416 7984 4448
rect 8016 4416 8052 4448
rect 8084 4416 8120 4448
rect 8152 4416 8188 4448
rect 8220 4416 8256 4448
rect 8288 4416 8324 4448
rect 8356 4416 8392 4448
rect 8424 4416 8460 4448
rect 8492 4416 8528 4448
rect 8560 4416 8596 4448
rect 8628 4416 8664 4448
rect 8696 4416 8732 4448
rect 8764 4416 8800 4448
rect 8832 4416 8868 4448
rect 8900 4416 8936 4448
rect 8968 4416 9004 4448
rect 9036 4416 9072 4448
rect 9104 4416 9140 4448
rect 9172 4416 9208 4448
rect 9240 4416 9276 4448
rect 9308 4416 9344 4448
rect 9376 4416 9412 4448
rect 9444 4416 9480 4448
rect 9512 4416 9548 4448
rect 9580 4416 9616 4448
rect 9648 4416 9684 4448
rect 9716 4416 9752 4448
rect 9784 4416 9820 4448
rect 9852 4416 9888 4448
rect 9920 4416 9956 4448
rect 9988 4416 10024 4448
rect 10056 4416 10092 4448
rect 10124 4416 10160 4448
rect 10192 4416 10228 4448
rect 10260 4416 10296 4448
rect 10328 4416 10364 4448
rect 10396 4416 10432 4448
rect 10464 4416 10500 4448
rect 10532 4416 10568 4448
rect 10600 4416 10636 4448
rect 10668 4416 10704 4448
rect 10736 4416 10772 4448
rect 10804 4416 10840 4448
rect 10872 4416 10908 4448
rect 10940 4416 10976 4448
rect 11008 4416 11044 4448
rect 11076 4416 11112 4448
rect 11144 4416 11180 4448
rect 11212 4416 11248 4448
rect 11280 4416 11316 4448
rect 11348 4416 11384 4448
rect 11416 4416 11452 4448
rect 11484 4416 11520 4448
rect 11552 4416 11588 4448
rect 11620 4416 11656 4448
rect 11688 4416 11724 4448
rect 11756 4416 11792 4448
rect 11824 4416 11860 4448
rect 11892 4416 11928 4448
rect 11960 4416 11996 4448
rect 12028 4416 12064 4448
rect 12096 4416 12132 4448
rect 12164 4416 12200 4448
rect 12232 4416 12268 4448
rect 12300 4416 12336 4448
rect 12368 4416 12404 4448
rect 12436 4416 12472 4448
rect 12504 4416 12540 4448
rect 12572 4416 12608 4448
rect 12640 4416 12676 4448
rect 12708 4416 12744 4448
rect 12776 4416 12812 4448
rect 12844 4416 12880 4448
rect 12912 4416 12948 4448
rect 12980 4416 13016 4448
rect 13048 4416 13084 4448
rect 13116 4416 13152 4448
rect 13184 4416 13220 4448
rect 13252 4416 13288 4448
rect 13320 4416 13356 4448
rect 13388 4416 13424 4448
rect 13456 4416 13492 4448
rect 13524 4416 13560 4448
rect 13592 4416 13628 4448
rect 13660 4416 13696 4448
rect 13728 4416 13764 4448
rect 13796 4416 13832 4448
rect 13864 4416 13900 4448
rect 13932 4416 13968 4448
rect 14000 4416 14036 4448
rect 14068 4416 14104 4448
rect 14136 4416 14172 4448
rect 14204 4416 14240 4448
rect 14272 4416 14308 4448
rect 14340 4416 14376 4448
rect 14408 4416 14444 4448
rect 14476 4416 14512 4448
rect 14544 4416 14580 4448
rect 14612 4416 14648 4448
rect 14680 4416 14716 4448
rect 14748 4416 14784 4448
rect 14816 4416 14852 4448
rect 14884 4416 14920 4448
rect 14952 4416 14988 4448
rect 15020 4416 15056 4448
rect 15088 4416 15124 4448
rect 15156 4416 15192 4448
rect 15224 4416 15260 4448
rect 15292 4416 15328 4448
rect 15360 4416 15396 4448
rect 15428 4416 15464 4448
rect 15496 4416 15532 4448
rect 15564 4416 15600 4448
rect 15632 4416 15668 4448
rect 15700 4416 15736 4448
rect 15768 4416 15804 4448
rect 15836 4416 15872 4448
rect 15904 4416 15940 4448
rect 15972 4416 16000 4448
rect 0 4398 16000 4416
rect 0 4357 68 4398
rect 0 4325 18 4357
rect 50 4325 68 4357
rect 0 4289 68 4325
rect 0 4257 18 4289
rect 50 4257 68 4289
rect 0 4221 68 4257
rect 0 4189 18 4221
rect 50 4189 68 4221
rect 0 4153 68 4189
rect 0 4121 18 4153
rect 50 4121 68 4153
rect 0 4085 68 4121
rect 15932 4357 16000 4398
rect 15932 4325 15950 4357
rect 15982 4325 16000 4357
rect 15932 4289 16000 4325
rect 15932 4257 15950 4289
rect 15982 4257 16000 4289
rect 15932 4221 16000 4257
rect 15932 4189 15950 4221
rect 15982 4189 16000 4221
rect 15932 4153 16000 4189
rect 15932 4121 15950 4153
rect 15982 4121 16000 4153
rect 0 4053 18 4085
rect 50 4053 68 4085
rect 15932 4085 16000 4121
rect 0 4017 68 4053
rect 0 3985 18 4017
rect 50 3985 68 4017
rect 0 3949 68 3985
rect 0 3917 18 3949
rect 50 3917 68 3949
rect 0 3881 68 3917
rect 0 3849 18 3881
rect 50 3849 68 3881
rect 0 3813 68 3849
rect 0 3781 18 3813
rect 50 3781 68 3813
rect 0 3745 68 3781
rect 0 3713 18 3745
rect 50 3713 68 3745
rect 0 3677 68 3713
rect 0 3645 18 3677
rect 50 3645 68 3677
rect 0 3609 68 3645
rect 0 3577 18 3609
rect 50 3577 68 3609
rect 0 3541 68 3577
rect 0 3509 18 3541
rect 50 3509 68 3541
rect 0 3473 68 3509
rect 0 3441 18 3473
rect 50 3441 68 3473
rect 0 3405 68 3441
rect 0 3373 18 3405
rect 50 3373 68 3405
rect 0 3337 68 3373
rect 0 3305 18 3337
rect 50 3305 68 3337
rect 0 3269 68 3305
rect 0 3237 18 3269
rect 50 3237 68 3269
rect 0 3201 68 3237
rect 0 3169 18 3201
rect 50 3169 68 3201
rect 0 3133 68 3169
rect 0 3101 18 3133
rect 50 3101 68 3133
rect 0 3065 68 3101
rect 0 3033 18 3065
rect 50 3033 68 3065
rect 0 2997 68 3033
rect 0 2965 18 2997
rect 50 2965 68 2997
rect 0 2929 68 2965
rect 0 2897 18 2929
rect 50 2897 68 2929
rect 0 2861 68 2897
rect 0 2829 18 2861
rect 50 2829 68 2861
rect 0 2793 68 2829
rect 0 2761 18 2793
rect 50 2761 68 2793
rect 0 2725 68 2761
rect 0 2693 18 2725
rect 50 2693 68 2725
rect 0 2657 68 2693
rect 0 2625 18 2657
rect 50 2625 68 2657
rect 0 2589 68 2625
rect 0 2557 18 2589
rect 50 2557 68 2589
rect 0 2521 68 2557
rect 0 2489 18 2521
rect 50 2489 68 2521
rect 0 2453 68 2489
rect 0 2421 18 2453
rect 50 2421 68 2453
rect 0 2385 68 2421
rect 0 2353 18 2385
rect 50 2353 68 2385
rect 0 2317 68 2353
rect 0 2285 18 2317
rect 50 2285 68 2317
rect 0 2249 68 2285
rect 15932 4053 15950 4085
rect 15982 4053 16000 4085
rect 15932 4017 16000 4053
rect 15932 3985 15950 4017
rect 15982 3985 16000 4017
rect 15932 3949 16000 3985
rect 15932 3917 15950 3949
rect 15982 3917 16000 3949
rect 15932 3881 16000 3917
rect 15932 3849 15950 3881
rect 15982 3849 16000 3881
rect 15932 3813 16000 3849
rect 15932 3781 15950 3813
rect 15982 3781 16000 3813
rect 15932 3745 16000 3781
rect 15932 3713 15950 3745
rect 15982 3713 16000 3745
rect 15932 3677 16000 3713
rect 15932 3645 15950 3677
rect 15982 3645 16000 3677
rect 15932 3609 16000 3645
rect 15932 3577 15950 3609
rect 15982 3577 16000 3609
rect 15932 3541 16000 3577
rect 15932 3509 15950 3541
rect 15982 3509 16000 3541
rect 15932 3473 16000 3509
rect 15932 3441 15950 3473
rect 15982 3441 16000 3473
rect 15932 3405 16000 3441
rect 15932 3373 15950 3405
rect 15982 3373 16000 3405
rect 15932 3337 16000 3373
rect 15932 3305 15950 3337
rect 15982 3305 16000 3337
rect 15932 3269 16000 3305
rect 15932 3237 15950 3269
rect 15982 3237 16000 3269
rect 15932 3201 16000 3237
rect 15932 3169 15950 3201
rect 15982 3169 16000 3201
rect 15932 3133 16000 3169
rect 15932 3101 15950 3133
rect 15982 3101 16000 3133
rect 15932 3065 16000 3101
rect 15932 3033 15950 3065
rect 15982 3033 16000 3065
rect 15932 2997 16000 3033
rect 15932 2965 15950 2997
rect 15982 2965 16000 2997
rect 15932 2929 16000 2965
rect 15932 2897 15950 2929
rect 15982 2897 16000 2929
rect 15932 2861 16000 2897
rect 15932 2829 15950 2861
rect 15982 2829 16000 2861
rect 15932 2793 16000 2829
rect 15932 2761 15950 2793
rect 15982 2761 16000 2793
rect 15932 2725 16000 2761
rect 15932 2693 15950 2725
rect 15982 2693 16000 2725
rect 15932 2657 16000 2693
rect 15932 2625 15950 2657
rect 15982 2625 16000 2657
rect 15932 2589 16000 2625
rect 15932 2557 15950 2589
rect 15982 2557 16000 2589
rect 15932 2521 16000 2557
rect 15932 2489 15950 2521
rect 15982 2489 16000 2521
rect 15932 2453 16000 2489
rect 15932 2421 15950 2453
rect 15982 2421 16000 2453
rect 15932 2385 16000 2421
rect 15932 2353 15950 2385
rect 15982 2353 16000 2385
rect 15932 2317 16000 2353
rect 15932 2285 15950 2317
rect 15982 2285 16000 2317
rect 0 2217 18 2249
rect 50 2217 68 2249
rect 0 2181 68 2217
rect 15932 2249 16000 2285
rect 15932 2217 15950 2249
rect 15982 2217 16000 2249
rect 0 2149 18 2181
rect 50 2149 68 2181
rect 0 2113 68 2149
rect 0 2081 18 2113
rect 50 2081 68 2113
rect 0 2045 68 2081
rect 0 2013 18 2045
rect 50 2013 68 2045
rect 0 1977 68 2013
rect 0 1945 18 1977
rect 50 1945 68 1977
rect 0 1909 68 1945
rect 0 1877 18 1909
rect 50 1877 68 1909
rect 0 1841 68 1877
rect 0 1809 18 1841
rect 50 1809 68 1841
rect 0 1773 68 1809
rect 0 1741 18 1773
rect 50 1741 68 1773
rect 0 1705 68 1741
rect 0 1673 18 1705
rect 50 1673 68 1705
rect 0 1637 68 1673
rect 0 1605 18 1637
rect 50 1605 68 1637
rect 0 1569 68 1605
rect 0 1537 18 1569
rect 50 1537 68 1569
rect 0 1501 68 1537
rect 0 1469 18 1501
rect 50 1469 68 1501
rect 0 1433 68 1469
rect 0 1401 18 1433
rect 50 1401 68 1433
rect 0 1365 68 1401
rect 0 1333 18 1365
rect 50 1333 68 1365
rect 0 1297 68 1333
rect 0 1265 18 1297
rect 50 1265 68 1297
rect 0 1229 68 1265
rect 0 1197 18 1229
rect 50 1197 68 1229
rect 0 1161 68 1197
rect 0 1129 18 1161
rect 50 1129 68 1161
rect 0 1093 68 1129
rect 0 1061 18 1093
rect 50 1061 68 1093
rect 0 1025 68 1061
rect 0 993 18 1025
rect 50 993 68 1025
rect 0 957 68 993
rect 0 925 18 957
rect 50 925 68 957
rect 0 889 68 925
rect 0 857 18 889
rect 50 857 68 889
rect 0 821 68 857
rect 0 789 18 821
rect 50 789 68 821
rect 0 753 68 789
rect 0 721 18 753
rect 50 721 68 753
rect 0 685 68 721
rect 0 653 18 685
rect 50 653 68 685
rect 0 617 68 653
rect 0 585 18 617
rect 50 585 68 617
rect 0 549 68 585
rect 0 517 18 549
rect 50 517 68 549
rect 0 481 68 517
rect 0 449 18 481
rect 50 449 68 481
rect 0 413 68 449
rect 0 381 18 413
rect 50 381 68 413
rect 15932 2181 16000 2217
rect 15932 2149 15950 2181
rect 15982 2149 16000 2181
rect 15932 2113 16000 2149
rect 15932 2081 15950 2113
rect 15982 2081 16000 2113
rect 15932 2045 16000 2081
rect 15932 2013 15950 2045
rect 15982 2013 16000 2045
rect 15932 1977 16000 2013
rect 15932 1945 15950 1977
rect 15982 1945 16000 1977
rect 15932 1909 16000 1945
rect 15932 1877 15950 1909
rect 15982 1877 16000 1909
rect 15932 1841 16000 1877
rect 15932 1809 15950 1841
rect 15982 1809 16000 1841
rect 15932 1773 16000 1809
rect 15932 1741 15950 1773
rect 15982 1741 16000 1773
rect 15932 1705 16000 1741
rect 15932 1673 15950 1705
rect 15982 1673 16000 1705
rect 15932 1637 16000 1673
rect 15932 1605 15950 1637
rect 15982 1605 16000 1637
rect 15932 1569 16000 1605
rect 15932 1537 15950 1569
rect 15982 1537 16000 1569
rect 15932 1501 16000 1537
rect 15932 1469 15950 1501
rect 15982 1469 16000 1501
rect 15932 1433 16000 1469
rect 15932 1401 15950 1433
rect 15982 1401 16000 1433
rect 15932 1365 16000 1401
rect 15932 1333 15950 1365
rect 15982 1333 16000 1365
rect 15932 1297 16000 1333
rect 15932 1265 15950 1297
rect 15982 1265 16000 1297
rect 15932 1229 16000 1265
rect 15932 1197 15950 1229
rect 15982 1197 16000 1229
rect 15932 1161 16000 1197
rect 15932 1129 15950 1161
rect 15982 1129 16000 1161
rect 15932 1093 16000 1129
rect 15932 1061 15950 1093
rect 15982 1061 16000 1093
rect 15932 1025 16000 1061
rect 15932 993 15950 1025
rect 15982 993 16000 1025
rect 15932 957 16000 993
rect 15932 925 15950 957
rect 15982 925 16000 957
rect 15932 889 16000 925
rect 15932 857 15950 889
rect 15982 857 16000 889
rect 15932 821 16000 857
rect 15932 789 15950 821
rect 15982 789 16000 821
rect 15932 753 16000 789
rect 15932 721 15950 753
rect 15982 721 16000 753
rect 15932 685 16000 721
rect 15932 653 15950 685
rect 15982 653 16000 685
rect 15932 617 16000 653
rect 15932 585 15950 617
rect 15982 585 16000 617
rect 15932 549 16000 585
rect 15932 517 15950 549
rect 15982 517 16000 549
rect 15932 481 16000 517
rect 15932 449 15950 481
rect 15982 449 16000 481
rect 15932 413 16000 449
rect 0 345 68 381
rect 0 313 18 345
rect 50 313 68 345
rect 15932 381 15950 413
rect 15982 381 16000 413
rect 15932 345 16000 381
rect 0 277 68 313
rect 0 245 18 277
rect 50 245 68 277
rect 0 209 68 245
rect 0 177 18 209
rect 50 177 68 209
rect 0 141 68 177
rect 0 109 18 141
rect 50 109 68 141
rect 0 68 68 109
rect 15932 313 15950 345
rect 15982 313 16000 345
rect 15932 277 16000 313
rect 15932 245 15950 277
rect 15982 245 16000 277
rect 15932 209 16000 245
rect 15932 177 15950 209
rect 15982 177 16000 209
rect 15932 141 16000 177
rect 15932 109 15950 141
rect 15982 109 16000 141
rect 15932 68 16000 109
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< nsubdiff >>
rect 3264 7072 12736 7090
rect 3264 7040 3292 7072
rect 3324 7040 3360 7072
rect 3392 7040 3428 7072
rect 3460 7040 3496 7072
rect 3528 7040 3564 7072
rect 3596 7040 3632 7072
rect 3664 7040 3700 7072
rect 3732 7040 3768 7072
rect 3800 7040 3836 7072
rect 3868 7040 3904 7072
rect 3936 7040 3972 7072
rect 4004 7040 4040 7072
rect 4072 7040 4108 7072
rect 4140 7040 4176 7072
rect 4208 7040 4244 7072
rect 4276 7040 4312 7072
rect 4344 7040 4380 7072
rect 4412 7040 4448 7072
rect 4480 7040 4516 7072
rect 4548 7040 4584 7072
rect 4616 7040 4652 7072
rect 4684 7040 4720 7072
rect 4752 7040 4788 7072
rect 4820 7040 4856 7072
rect 4888 7040 4924 7072
rect 4956 7040 4992 7072
rect 5024 7040 5060 7072
rect 5092 7040 5128 7072
rect 5160 7040 5196 7072
rect 5228 7040 5264 7072
rect 5296 7040 5332 7072
rect 5364 7040 5400 7072
rect 5432 7040 5468 7072
rect 5500 7040 5536 7072
rect 5568 7040 5604 7072
rect 5636 7040 5672 7072
rect 5704 7040 5740 7072
rect 5772 7040 5808 7072
rect 5840 7040 5876 7072
rect 5908 7040 5944 7072
rect 5976 7040 6012 7072
rect 6044 7040 6080 7072
rect 6112 7040 6148 7072
rect 6180 7040 6216 7072
rect 6248 7040 6284 7072
rect 6316 7040 6352 7072
rect 6384 7040 6420 7072
rect 6452 7040 6488 7072
rect 6520 7040 6556 7072
rect 6588 7040 6624 7072
rect 6656 7040 6692 7072
rect 6724 7040 6760 7072
rect 6792 7040 6828 7072
rect 6860 7040 6896 7072
rect 6928 7040 6964 7072
rect 6996 7040 7032 7072
rect 7064 7040 7100 7072
rect 7132 7040 7168 7072
rect 7200 7040 7236 7072
rect 7268 7040 7304 7072
rect 7336 7040 7372 7072
rect 7404 7040 7440 7072
rect 7472 7040 7508 7072
rect 7540 7040 7576 7072
rect 7608 7040 7644 7072
rect 7676 7040 7712 7072
rect 7744 7040 7780 7072
rect 7812 7040 7848 7072
rect 7880 7040 7916 7072
rect 7948 7040 7984 7072
rect 8016 7040 8052 7072
rect 8084 7040 8120 7072
rect 8152 7040 8188 7072
rect 8220 7040 8256 7072
rect 8288 7040 8324 7072
rect 8356 7040 8392 7072
rect 8424 7040 8460 7072
rect 8492 7040 8528 7072
rect 8560 7040 8596 7072
rect 8628 7040 8664 7072
rect 8696 7040 8732 7072
rect 8764 7040 8800 7072
rect 8832 7040 8868 7072
rect 8900 7040 8936 7072
rect 8968 7040 9004 7072
rect 9036 7040 9072 7072
rect 9104 7040 9140 7072
rect 9172 7040 9208 7072
rect 9240 7040 9276 7072
rect 9308 7040 9344 7072
rect 9376 7040 9412 7072
rect 9444 7040 9480 7072
rect 9512 7040 9548 7072
rect 9580 7040 9616 7072
rect 9648 7040 9684 7072
rect 9716 7040 9752 7072
rect 9784 7040 9820 7072
rect 9852 7040 9888 7072
rect 9920 7040 9956 7072
rect 9988 7040 10024 7072
rect 10056 7040 10092 7072
rect 10124 7040 10160 7072
rect 10192 7040 10228 7072
rect 10260 7040 10296 7072
rect 10328 7040 10364 7072
rect 10396 7040 10432 7072
rect 10464 7040 10500 7072
rect 10532 7040 10568 7072
rect 10600 7040 10636 7072
rect 10668 7040 10704 7072
rect 10736 7040 10772 7072
rect 10804 7040 10840 7072
rect 10872 7040 10908 7072
rect 10940 7040 10976 7072
rect 11008 7040 11044 7072
rect 11076 7040 11112 7072
rect 11144 7040 11180 7072
rect 11212 7040 11248 7072
rect 11280 7040 11316 7072
rect 11348 7040 11384 7072
rect 11416 7040 11452 7072
rect 11484 7040 11520 7072
rect 11552 7040 11588 7072
rect 11620 7040 11656 7072
rect 11688 7040 11724 7072
rect 11756 7040 11792 7072
rect 11824 7040 11860 7072
rect 11892 7040 11928 7072
rect 11960 7040 11996 7072
rect 12028 7040 12064 7072
rect 12096 7040 12132 7072
rect 12164 7040 12200 7072
rect 12232 7040 12268 7072
rect 12300 7040 12336 7072
rect 12368 7040 12404 7072
rect 12436 7040 12472 7072
rect 12504 7040 12540 7072
rect 12572 7040 12608 7072
rect 12640 7040 12676 7072
rect 12708 7040 12736 7072
rect 3264 7022 12736 7040
rect 3264 6984 3332 7022
rect 3264 6952 3282 6984
rect 3314 6952 3332 6984
rect 3264 6916 3332 6952
rect 3264 6884 3282 6916
rect 3314 6884 3332 6916
rect 3264 6848 3332 6884
rect 3264 6816 3282 6848
rect 3314 6816 3332 6848
rect 3264 6780 3332 6816
rect 3264 6748 3282 6780
rect 3314 6748 3332 6780
rect 12668 6984 12736 7022
rect 12668 6952 12686 6984
rect 12718 6952 12736 6984
rect 12668 6916 12736 6952
rect 12668 6884 12686 6916
rect 12718 6884 12736 6916
rect 12668 6848 12736 6884
rect 12668 6816 12686 6848
rect 12718 6816 12736 6848
rect 12668 6780 12736 6816
rect 3264 6712 3332 6748
rect 3264 6680 3282 6712
rect 3314 6680 3332 6712
rect 12668 6748 12686 6780
rect 12718 6748 12736 6780
rect 12668 6712 12736 6748
rect 3264 6644 3332 6680
rect 3264 6612 3282 6644
rect 3314 6612 3332 6644
rect 3264 6576 3332 6612
rect 3264 6544 3282 6576
rect 3314 6544 3332 6576
rect 3264 6508 3332 6544
rect 3264 6476 3282 6508
rect 3314 6476 3332 6508
rect 3264 6440 3332 6476
rect 3264 6408 3282 6440
rect 3314 6408 3332 6440
rect 3264 6372 3332 6408
rect 3264 6340 3282 6372
rect 3314 6340 3332 6372
rect 3264 6304 3332 6340
rect 3264 6272 3282 6304
rect 3314 6272 3332 6304
rect 3264 6236 3332 6272
rect 3264 6204 3282 6236
rect 3314 6204 3332 6236
rect 3264 6168 3332 6204
rect 3264 6136 3282 6168
rect 3314 6136 3332 6168
rect 3264 6100 3332 6136
rect 3264 6068 3282 6100
rect 3314 6068 3332 6100
rect 3264 6032 3332 6068
rect 3264 6000 3282 6032
rect 3314 6000 3332 6032
rect 3264 5964 3332 6000
rect 3264 5932 3282 5964
rect 3314 5932 3332 5964
rect 3264 5896 3332 5932
rect 3264 5864 3282 5896
rect 3314 5864 3332 5896
rect 3264 5828 3332 5864
rect 3264 5796 3282 5828
rect 3314 5796 3332 5828
rect 3264 5760 3332 5796
rect 3264 5728 3282 5760
rect 3314 5728 3332 5760
rect 3264 5692 3332 5728
rect 3264 5660 3282 5692
rect 3314 5660 3332 5692
rect 3264 5624 3332 5660
rect 3264 5592 3282 5624
rect 3314 5592 3332 5624
rect 3264 5556 3332 5592
rect 3264 5524 3282 5556
rect 3314 5524 3332 5556
rect 3264 5488 3332 5524
rect 3264 5456 3282 5488
rect 3314 5456 3332 5488
rect 3264 5420 3332 5456
rect 3264 5388 3282 5420
rect 3314 5388 3332 5420
rect 3264 5352 3332 5388
rect 3264 5320 3282 5352
rect 3314 5320 3332 5352
rect 3264 5284 3332 5320
rect 3264 5252 3282 5284
rect 3314 5252 3332 5284
rect 12668 6680 12686 6712
rect 12718 6680 12736 6712
rect 12668 6644 12736 6680
rect 12668 6612 12686 6644
rect 12718 6612 12736 6644
rect 12668 6576 12736 6612
rect 12668 6544 12686 6576
rect 12718 6544 12736 6576
rect 12668 6508 12736 6544
rect 12668 6476 12686 6508
rect 12718 6476 12736 6508
rect 12668 6440 12736 6476
rect 12668 6408 12686 6440
rect 12718 6408 12736 6440
rect 12668 6372 12736 6408
rect 12668 6340 12686 6372
rect 12718 6340 12736 6372
rect 12668 6304 12736 6340
rect 12668 6272 12686 6304
rect 12718 6272 12736 6304
rect 12668 6236 12736 6272
rect 12668 6204 12686 6236
rect 12718 6204 12736 6236
rect 12668 6168 12736 6204
rect 12668 6136 12686 6168
rect 12718 6136 12736 6168
rect 12668 6100 12736 6136
rect 12668 6068 12686 6100
rect 12718 6068 12736 6100
rect 12668 6032 12736 6068
rect 12668 6000 12686 6032
rect 12718 6000 12736 6032
rect 12668 5964 12736 6000
rect 12668 5932 12686 5964
rect 12718 5932 12736 5964
rect 12668 5896 12736 5932
rect 12668 5864 12686 5896
rect 12718 5864 12736 5896
rect 12668 5828 12736 5864
rect 12668 5796 12686 5828
rect 12718 5796 12736 5828
rect 12668 5760 12736 5796
rect 12668 5728 12686 5760
rect 12718 5728 12736 5760
rect 12668 5692 12736 5728
rect 12668 5660 12686 5692
rect 12718 5660 12736 5692
rect 12668 5624 12736 5660
rect 12668 5592 12686 5624
rect 12718 5592 12736 5624
rect 12668 5556 12736 5592
rect 12668 5524 12686 5556
rect 12718 5524 12736 5556
rect 12668 5488 12736 5524
rect 12668 5456 12686 5488
rect 12718 5456 12736 5488
rect 12668 5420 12736 5456
rect 12668 5388 12686 5420
rect 12718 5388 12736 5420
rect 12668 5352 12736 5388
rect 12668 5320 12686 5352
rect 12718 5320 12736 5352
rect 12668 5284 12736 5320
rect 3264 5216 3332 5252
rect 12668 5252 12686 5284
rect 12718 5252 12736 5284
rect 3264 5184 3282 5216
rect 3314 5184 3332 5216
rect 3264 5148 3332 5184
rect 3264 5116 3282 5148
rect 3314 5116 3332 5148
rect 3264 5080 3332 5116
rect 3264 5048 3282 5080
rect 3314 5048 3332 5080
rect 3264 5012 3332 5048
rect 3264 4980 3282 5012
rect 3314 4980 3332 5012
rect 3264 4942 3332 4980
rect 12668 5216 12736 5252
rect 12668 5184 12686 5216
rect 12718 5184 12736 5216
rect 12668 5148 12736 5184
rect 12668 5116 12686 5148
rect 12718 5116 12736 5148
rect 12668 5080 12736 5116
rect 12668 5048 12686 5080
rect 12718 5048 12736 5080
rect 12668 5012 12736 5048
rect 12668 4980 12686 5012
rect 12718 4980 12736 5012
rect 12668 4942 12736 4980
rect 3264 4924 12736 4942
rect 3264 4892 3292 4924
rect 3324 4892 3360 4924
rect 3392 4892 3428 4924
rect 3460 4892 3496 4924
rect 3528 4892 3564 4924
rect 3596 4892 3632 4924
rect 3664 4892 3700 4924
rect 3732 4892 3768 4924
rect 3800 4892 3836 4924
rect 3868 4892 3904 4924
rect 3936 4892 3972 4924
rect 4004 4892 4040 4924
rect 4072 4892 4108 4924
rect 4140 4892 4176 4924
rect 4208 4892 4244 4924
rect 4276 4892 4312 4924
rect 4344 4892 4380 4924
rect 4412 4892 4448 4924
rect 4480 4892 4516 4924
rect 4548 4892 4584 4924
rect 4616 4892 4652 4924
rect 4684 4892 4720 4924
rect 4752 4892 4788 4924
rect 4820 4892 4856 4924
rect 4888 4892 4924 4924
rect 4956 4892 4992 4924
rect 5024 4892 5060 4924
rect 5092 4892 5128 4924
rect 5160 4892 5196 4924
rect 5228 4892 5264 4924
rect 5296 4892 5332 4924
rect 5364 4892 5400 4924
rect 5432 4892 5468 4924
rect 5500 4892 5536 4924
rect 5568 4892 5604 4924
rect 5636 4892 5672 4924
rect 5704 4892 5740 4924
rect 5772 4892 5808 4924
rect 5840 4892 5876 4924
rect 5908 4892 5944 4924
rect 5976 4892 6012 4924
rect 6044 4892 6080 4924
rect 6112 4892 6148 4924
rect 6180 4892 6216 4924
rect 6248 4892 6284 4924
rect 6316 4892 6352 4924
rect 6384 4892 6420 4924
rect 6452 4892 6488 4924
rect 6520 4892 6556 4924
rect 6588 4892 6624 4924
rect 6656 4892 6692 4924
rect 6724 4892 6760 4924
rect 6792 4892 6828 4924
rect 6860 4892 6896 4924
rect 6928 4892 6964 4924
rect 6996 4892 7032 4924
rect 7064 4892 7100 4924
rect 7132 4892 7168 4924
rect 7200 4892 7236 4924
rect 7268 4892 7304 4924
rect 7336 4892 7372 4924
rect 7404 4892 7440 4924
rect 7472 4892 7508 4924
rect 7540 4892 7576 4924
rect 7608 4892 7644 4924
rect 7676 4892 7712 4924
rect 7744 4892 7780 4924
rect 7812 4892 7848 4924
rect 7880 4892 7916 4924
rect 7948 4892 7984 4924
rect 8016 4892 8052 4924
rect 8084 4892 8120 4924
rect 8152 4892 8188 4924
rect 8220 4892 8256 4924
rect 8288 4892 8324 4924
rect 8356 4892 8392 4924
rect 8424 4892 8460 4924
rect 8492 4892 8528 4924
rect 8560 4892 8596 4924
rect 8628 4892 8664 4924
rect 8696 4892 8732 4924
rect 8764 4892 8800 4924
rect 8832 4892 8868 4924
rect 8900 4892 8936 4924
rect 8968 4892 9004 4924
rect 9036 4892 9072 4924
rect 9104 4892 9140 4924
rect 9172 4892 9208 4924
rect 9240 4892 9276 4924
rect 9308 4892 9344 4924
rect 9376 4892 9412 4924
rect 9444 4892 9480 4924
rect 9512 4892 9548 4924
rect 9580 4892 9616 4924
rect 9648 4892 9684 4924
rect 9716 4892 9752 4924
rect 9784 4892 9820 4924
rect 9852 4892 9888 4924
rect 9920 4892 9956 4924
rect 9988 4892 10024 4924
rect 10056 4892 10092 4924
rect 10124 4892 10160 4924
rect 10192 4892 10228 4924
rect 10260 4892 10296 4924
rect 10328 4892 10364 4924
rect 10396 4892 10432 4924
rect 10464 4892 10500 4924
rect 10532 4892 10568 4924
rect 10600 4892 10636 4924
rect 10668 4892 10704 4924
rect 10736 4892 10772 4924
rect 10804 4892 10840 4924
rect 10872 4892 10908 4924
rect 10940 4892 10976 4924
rect 11008 4892 11044 4924
rect 11076 4892 11112 4924
rect 11144 4892 11180 4924
rect 11212 4892 11248 4924
rect 11280 4892 11316 4924
rect 11348 4892 11384 4924
rect 11416 4892 11452 4924
rect 11484 4892 11520 4924
rect 11552 4892 11588 4924
rect 11620 4892 11656 4924
rect 11688 4892 11724 4924
rect 11756 4892 11792 4924
rect 11824 4892 11860 4924
rect 11892 4892 11928 4924
rect 11960 4892 11996 4924
rect 12028 4892 12064 4924
rect 12096 4892 12132 4924
rect 12164 4892 12200 4924
rect 12232 4892 12268 4924
rect 12300 4892 12336 4924
rect 12368 4892 12404 4924
rect 12436 4892 12472 4924
rect 12504 4892 12540 4924
rect 12572 4892 12608 4924
rect 12640 4892 12676 4924
rect 12708 4892 12736 4924
rect 3264 4874 12736 4892
<< psubdiffcont >>
rect 28 4416 60 4448
rect 96 4416 128 4448
rect 164 4416 196 4448
rect 232 4416 264 4448
rect 300 4416 332 4448
rect 368 4416 400 4448
rect 436 4416 468 4448
rect 504 4416 536 4448
rect 572 4416 604 4448
rect 640 4416 672 4448
rect 708 4416 740 4448
rect 776 4416 808 4448
rect 844 4416 876 4448
rect 912 4416 944 4448
rect 980 4416 1012 4448
rect 1048 4416 1080 4448
rect 1116 4416 1148 4448
rect 1184 4416 1216 4448
rect 1252 4416 1284 4448
rect 1320 4416 1352 4448
rect 1388 4416 1420 4448
rect 1456 4416 1488 4448
rect 1524 4416 1556 4448
rect 1592 4416 1624 4448
rect 1660 4416 1692 4448
rect 1728 4416 1760 4448
rect 1796 4416 1828 4448
rect 1864 4416 1896 4448
rect 1932 4416 1964 4448
rect 2000 4416 2032 4448
rect 2068 4416 2100 4448
rect 2136 4416 2168 4448
rect 2204 4416 2236 4448
rect 2272 4416 2304 4448
rect 2340 4416 2372 4448
rect 2408 4416 2440 4448
rect 2476 4416 2508 4448
rect 2544 4416 2576 4448
rect 2612 4416 2644 4448
rect 2680 4416 2712 4448
rect 2748 4416 2780 4448
rect 2816 4416 2848 4448
rect 2884 4416 2916 4448
rect 2952 4416 2984 4448
rect 3020 4416 3052 4448
rect 3088 4416 3120 4448
rect 3156 4416 3188 4448
rect 3224 4416 3256 4448
rect 3292 4416 3324 4448
rect 3360 4416 3392 4448
rect 3428 4416 3460 4448
rect 3496 4416 3528 4448
rect 3564 4416 3596 4448
rect 3632 4416 3664 4448
rect 3700 4416 3732 4448
rect 3768 4416 3800 4448
rect 3836 4416 3868 4448
rect 3904 4416 3936 4448
rect 3972 4416 4004 4448
rect 4040 4416 4072 4448
rect 4108 4416 4140 4448
rect 4176 4416 4208 4448
rect 4244 4416 4276 4448
rect 4312 4416 4344 4448
rect 4380 4416 4412 4448
rect 4448 4416 4480 4448
rect 4516 4416 4548 4448
rect 4584 4416 4616 4448
rect 4652 4416 4684 4448
rect 4720 4416 4752 4448
rect 4788 4416 4820 4448
rect 4856 4416 4888 4448
rect 4924 4416 4956 4448
rect 4992 4416 5024 4448
rect 5060 4416 5092 4448
rect 5128 4416 5160 4448
rect 5196 4416 5228 4448
rect 5264 4416 5296 4448
rect 5332 4416 5364 4448
rect 5400 4416 5432 4448
rect 5468 4416 5500 4448
rect 5536 4416 5568 4448
rect 5604 4416 5636 4448
rect 5672 4416 5704 4448
rect 5740 4416 5772 4448
rect 5808 4416 5840 4448
rect 5876 4416 5908 4448
rect 5944 4416 5976 4448
rect 6012 4416 6044 4448
rect 6080 4416 6112 4448
rect 6148 4416 6180 4448
rect 6216 4416 6248 4448
rect 6284 4416 6316 4448
rect 6352 4416 6384 4448
rect 6420 4416 6452 4448
rect 6488 4416 6520 4448
rect 6556 4416 6588 4448
rect 6624 4416 6656 4448
rect 6692 4416 6724 4448
rect 6760 4416 6792 4448
rect 6828 4416 6860 4448
rect 6896 4416 6928 4448
rect 6964 4416 6996 4448
rect 7032 4416 7064 4448
rect 7100 4416 7132 4448
rect 7168 4416 7200 4448
rect 7236 4416 7268 4448
rect 7304 4416 7336 4448
rect 7372 4416 7404 4448
rect 7440 4416 7472 4448
rect 7508 4416 7540 4448
rect 7576 4416 7608 4448
rect 7644 4416 7676 4448
rect 7712 4416 7744 4448
rect 7780 4416 7812 4448
rect 7848 4416 7880 4448
rect 7916 4416 7948 4448
rect 7984 4416 8016 4448
rect 8052 4416 8084 4448
rect 8120 4416 8152 4448
rect 8188 4416 8220 4448
rect 8256 4416 8288 4448
rect 8324 4416 8356 4448
rect 8392 4416 8424 4448
rect 8460 4416 8492 4448
rect 8528 4416 8560 4448
rect 8596 4416 8628 4448
rect 8664 4416 8696 4448
rect 8732 4416 8764 4448
rect 8800 4416 8832 4448
rect 8868 4416 8900 4448
rect 8936 4416 8968 4448
rect 9004 4416 9036 4448
rect 9072 4416 9104 4448
rect 9140 4416 9172 4448
rect 9208 4416 9240 4448
rect 9276 4416 9308 4448
rect 9344 4416 9376 4448
rect 9412 4416 9444 4448
rect 9480 4416 9512 4448
rect 9548 4416 9580 4448
rect 9616 4416 9648 4448
rect 9684 4416 9716 4448
rect 9752 4416 9784 4448
rect 9820 4416 9852 4448
rect 9888 4416 9920 4448
rect 9956 4416 9988 4448
rect 10024 4416 10056 4448
rect 10092 4416 10124 4448
rect 10160 4416 10192 4448
rect 10228 4416 10260 4448
rect 10296 4416 10328 4448
rect 10364 4416 10396 4448
rect 10432 4416 10464 4448
rect 10500 4416 10532 4448
rect 10568 4416 10600 4448
rect 10636 4416 10668 4448
rect 10704 4416 10736 4448
rect 10772 4416 10804 4448
rect 10840 4416 10872 4448
rect 10908 4416 10940 4448
rect 10976 4416 11008 4448
rect 11044 4416 11076 4448
rect 11112 4416 11144 4448
rect 11180 4416 11212 4448
rect 11248 4416 11280 4448
rect 11316 4416 11348 4448
rect 11384 4416 11416 4448
rect 11452 4416 11484 4448
rect 11520 4416 11552 4448
rect 11588 4416 11620 4448
rect 11656 4416 11688 4448
rect 11724 4416 11756 4448
rect 11792 4416 11824 4448
rect 11860 4416 11892 4448
rect 11928 4416 11960 4448
rect 11996 4416 12028 4448
rect 12064 4416 12096 4448
rect 12132 4416 12164 4448
rect 12200 4416 12232 4448
rect 12268 4416 12300 4448
rect 12336 4416 12368 4448
rect 12404 4416 12436 4448
rect 12472 4416 12504 4448
rect 12540 4416 12572 4448
rect 12608 4416 12640 4448
rect 12676 4416 12708 4448
rect 12744 4416 12776 4448
rect 12812 4416 12844 4448
rect 12880 4416 12912 4448
rect 12948 4416 12980 4448
rect 13016 4416 13048 4448
rect 13084 4416 13116 4448
rect 13152 4416 13184 4448
rect 13220 4416 13252 4448
rect 13288 4416 13320 4448
rect 13356 4416 13388 4448
rect 13424 4416 13456 4448
rect 13492 4416 13524 4448
rect 13560 4416 13592 4448
rect 13628 4416 13660 4448
rect 13696 4416 13728 4448
rect 13764 4416 13796 4448
rect 13832 4416 13864 4448
rect 13900 4416 13932 4448
rect 13968 4416 14000 4448
rect 14036 4416 14068 4448
rect 14104 4416 14136 4448
rect 14172 4416 14204 4448
rect 14240 4416 14272 4448
rect 14308 4416 14340 4448
rect 14376 4416 14408 4448
rect 14444 4416 14476 4448
rect 14512 4416 14544 4448
rect 14580 4416 14612 4448
rect 14648 4416 14680 4448
rect 14716 4416 14748 4448
rect 14784 4416 14816 4448
rect 14852 4416 14884 4448
rect 14920 4416 14952 4448
rect 14988 4416 15020 4448
rect 15056 4416 15088 4448
rect 15124 4416 15156 4448
rect 15192 4416 15224 4448
rect 15260 4416 15292 4448
rect 15328 4416 15360 4448
rect 15396 4416 15428 4448
rect 15464 4416 15496 4448
rect 15532 4416 15564 4448
rect 15600 4416 15632 4448
rect 15668 4416 15700 4448
rect 15736 4416 15768 4448
rect 15804 4416 15836 4448
rect 15872 4416 15904 4448
rect 15940 4416 15972 4448
rect 18 4325 50 4357
rect 18 4257 50 4289
rect 18 4189 50 4221
rect 18 4121 50 4153
rect 15950 4325 15982 4357
rect 15950 4257 15982 4289
rect 15950 4189 15982 4221
rect 15950 4121 15982 4153
rect 18 4053 50 4085
rect 18 3985 50 4017
rect 18 3917 50 3949
rect 18 3849 50 3881
rect 18 3781 50 3813
rect 18 3713 50 3745
rect 18 3645 50 3677
rect 18 3577 50 3609
rect 18 3509 50 3541
rect 18 3441 50 3473
rect 18 3373 50 3405
rect 18 3305 50 3337
rect 18 3237 50 3269
rect 18 3169 50 3201
rect 18 3101 50 3133
rect 18 3033 50 3065
rect 18 2965 50 2997
rect 18 2897 50 2929
rect 18 2829 50 2861
rect 18 2761 50 2793
rect 18 2693 50 2725
rect 18 2625 50 2657
rect 18 2557 50 2589
rect 18 2489 50 2521
rect 18 2421 50 2453
rect 18 2353 50 2385
rect 18 2285 50 2317
rect 15950 4053 15982 4085
rect 15950 3985 15982 4017
rect 15950 3917 15982 3949
rect 15950 3849 15982 3881
rect 15950 3781 15982 3813
rect 15950 3713 15982 3745
rect 15950 3645 15982 3677
rect 15950 3577 15982 3609
rect 15950 3509 15982 3541
rect 15950 3441 15982 3473
rect 15950 3373 15982 3405
rect 15950 3305 15982 3337
rect 15950 3237 15982 3269
rect 15950 3169 15982 3201
rect 15950 3101 15982 3133
rect 15950 3033 15982 3065
rect 15950 2965 15982 2997
rect 15950 2897 15982 2929
rect 15950 2829 15982 2861
rect 15950 2761 15982 2793
rect 15950 2693 15982 2725
rect 15950 2625 15982 2657
rect 15950 2557 15982 2589
rect 15950 2489 15982 2521
rect 15950 2421 15982 2453
rect 15950 2353 15982 2385
rect 15950 2285 15982 2317
rect 18 2217 50 2249
rect 15950 2217 15982 2249
rect 18 2149 50 2181
rect 18 2081 50 2113
rect 18 2013 50 2045
rect 18 1945 50 1977
rect 18 1877 50 1909
rect 18 1809 50 1841
rect 18 1741 50 1773
rect 18 1673 50 1705
rect 18 1605 50 1637
rect 18 1537 50 1569
rect 18 1469 50 1501
rect 18 1401 50 1433
rect 18 1333 50 1365
rect 18 1265 50 1297
rect 18 1197 50 1229
rect 18 1129 50 1161
rect 18 1061 50 1093
rect 18 993 50 1025
rect 18 925 50 957
rect 18 857 50 889
rect 18 789 50 821
rect 18 721 50 753
rect 18 653 50 685
rect 18 585 50 617
rect 18 517 50 549
rect 18 449 50 481
rect 18 381 50 413
rect 15950 2149 15982 2181
rect 15950 2081 15982 2113
rect 15950 2013 15982 2045
rect 15950 1945 15982 1977
rect 15950 1877 15982 1909
rect 15950 1809 15982 1841
rect 15950 1741 15982 1773
rect 15950 1673 15982 1705
rect 15950 1605 15982 1637
rect 15950 1537 15982 1569
rect 15950 1469 15982 1501
rect 15950 1401 15982 1433
rect 15950 1333 15982 1365
rect 15950 1265 15982 1297
rect 15950 1197 15982 1229
rect 15950 1129 15982 1161
rect 15950 1061 15982 1093
rect 15950 993 15982 1025
rect 15950 925 15982 957
rect 15950 857 15982 889
rect 15950 789 15982 821
rect 15950 721 15982 753
rect 15950 653 15982 685
rect 15950 585 15982 617
rect 15950 517 15982 549
rect 15950 449 15982 481
rect 18 313 50 345
rect 15950 381 15982 413
rect 18 245 50 277
rect 18 177 50 209
rect 18 109 50 141
rect 15950 313 15982 345
rect 15950 245 15982 277
rect 15950 177 15982 209
rect 15950 109 15982 141
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< nsubdiffcont >>
rect 3292 7040 3324 7072
rect 3360 7040 3392 7072
rect 3428 7040 3460 7072
rect 3496 7040 3528 7072
rect 3564 7040 3596 7072
rect 3632 7040 3664 7072
rect 3700 7040 3732 7072
rect 3768 7040 3800 7072
rect 3836 7040 3868 7072
rect 3904 7040 3936 7072
rect 3972 7040 4004 7072
rect 4040 7040 4072 7072
rect 4108 7040 4140 7072
rect 4176 7040 4208 7072
rect 4244 7040 4276 7072
rect 4312 7040 4344 7072
rect 4380 7040 4412 7072
rect 4448 7040 4480 7072
rect 4516 7040 4548 7072
rect 4584 7040 4616 7072
rect 4652 7040 4684 7072
rect 4720 7040 4752 7072
rect 4788 7040 4820 7072
rect 4856 7040 4888 7072
rect 4924 7040 4956 7072
rect 4992 7040 5024 7072
rect 5060 7040 5092 7072
rect 5128 7040 5160 7072
rect 5196 7040 5228 7072
rect 5264 7040 5296 7072
rect 5332 7040 5364 7072
rect 5400 7040 5432 7072
rect 5468 7040 5500 7072
rect 5536 7040 5568 7072
rect 5604 7040 5636 7072
rect 5672 7040 5704 7072
rect 5740 7040 5772 7072
rect 5808 7040 5840 7072
rect 5876 7040 5908 7072
rect 5944 7040 5976 7072
rect 6012 7040 6044 7072
rect 6080 7040 6112 7072
rect 6148 7040 6180 7072
rect 6216 7040 6248 7072
rect 6284 7040 6316 7072
rect 6352 7040 6384 7072
rect 6420 7040 6452 7072
rect 6488 7040 6520 7072
rect 6556 7040 6588 7072
rect 6624 7040 6656 7072
rect 6692 7040 6724 7072
rect 6760 7040 6792 7072
rect 6828 7040 6860 7072
rect 6896 7040 6928 7072
rect 6964 7040 6996 7072
rect 7032 7040 7064 7072
rect 7100 7040 7132 7072
rect 7168 7040 7200 7072
rect 7236 7040 7268 7072
rect 7304 7040 7336 7072
rect 7372 7040 7404 7072
rect 7440 7040 7472 7072
rect 7508 7040 7540 7072
rect 7576 7040 7608 7072
rect 7644 7040 7676 7072
rect 7712 7040 7744 7072
rect 7780 7040 7812 7072
rect 7848 7040 7880 7072
rect 7916 7040 7948 7072
rect 7984 7040 8016 7072
rect 8052 7040 8084 7072
rect 8120 7040 8152 7072
rect 8188 7040 8220 7072
rect 8256 7040 8288 7072
rect 8324 7040 8356 7072
rect 8392 7040 8424 7072
rect 8460 7040 8492 7072
rect 8528 7040 8560 7072
rect 8596 7040 8628 7072
rect 8664 7040 8696 7072
rect 8732 7040 8764 7072
rect 8800 7040 8832 7072
rect 8868 7040 8900 7072
rect 8936 7040 8968 7072
rect 9004 7040 9036 7072
rect 9072 7040 9104 7072
rect 9140 7040 9172 7072
rect 9208 7040 9240 7072
rect 9276 7040 9308 7072
rect 9344 7040 9376 7072
rect 9412 7040 9444 7072
rect 9480 7040 9512 7072
rect 9548 7040 9580 7072
rect 9616 7040 9648 7072
rect 9684 7040 9716 7072
rect 9752 7040 9784 7072
rect 9820 7040 9852 7072
rect 9888 7040 9920 7072
rect 9956 7040 9988 7072
rect 10024 7040 10056 7072
rect 10092 7040 10124 7072
rect 10160 7040 10192 7072
rect 10228 7040 10260 7072
rect 10296 7040 10328 7072
rect 10364 7040 10396 7072
rect 10432 7040 10464 7072
rect 10500 7040 10532 7072
rect 10568 7040 10600 7072
rect 10636 7040 10668 7072
rect 10704 7040 10736 7072
rect 10772 7040 10804 7072
rect 10840 7040 10872 7072
rect 10908 7040 10940 7072
rect 10976 7040 11008 7072
rect 11044 7040 11076 7072
rect 11112 7040 11144 7072
rect 11180 7040 11212 7072
rect 11248 7040 11280 7072
rect 11316 7040 11348 7072
rect 11384 7040 11416 7072
rect 11452 7040 11484 7072
rect 11520 7040 11552 7072
rect 11588 7040 11620 7072
rect 11656 7040 11688 7072
rect 11724 7040 11756 7072
rect 11792 7040 11824 7072
rect 11860 7040 11892 7072
rect 11928 7040 11960 7072
rect 11996 7040 12028 7072
rect 12064 7040 12096 7072
rect 12132 7040 12164 7072
rect 12200 7040 12232 7072
rect 12268 7040 12300 7072
rect 12336 7040 12368 7072
rect 12404 7040 12436 7072
rect 12472 7040 12504 7072
rect 12540 7040 12572 7072
rect 12608 7040 12640 7072
rect 12676 7040 12708 7072
rect 3282 6952 3314 6984
rect 3282 6884 3314 6916
rect 3282 6816 3314 6848
rect 3282 6748 3314 6780
rect 12686 6952 12718 6984
rect 12686 6884 12718 6916
rect 12686 6816 12718 6848
rect 3282 6680 3314 6712
rect 12686 6748 12718 6780
rect 3282 6612 3314 6644
rect 3282 6544 3314 6576
rect 3282 6476 3314 6508
rect 3282 6408 3314 6440
rect 3282 6340 3314 6372
rect 3282 6272 3314 6304
rect 3282 6204 3314 6236
rect 3282 6136 3314 6168
rect 3282 6068 3314 6100
rect 3282 6000 3314 6032
rect 3282 5932 3314 5964
rect 3282 5864 3314 5896
rect 3282 5796 3314 5828
rect 3282 5728 3314 5760
rect 3282 5660 3314 5692
rect 3282 5592 3314 5624
rect 3282 5524 3314 5556
rect 3282 5456 3314 5488
rect 3282 5388 3314 5420
rect 3282 5320 3314 5352
rect 3282 5252 3314 5284
rect 12686 6680 12718 6712
rect 12686 6612 12718 6644
rect 12686 6544 12718 6576
rect 12686 6476 12718 6508
rect 12686 6408 12718 6440
rect 12686 6340 12718 6372
rect 12686 6272 12718 6304
rect 12686 6204 12718 6236
rect 12686 6136 12718 6168
rect 12686 6068 12718 6100
rect 12686 6000 12718 6032
rect 12686 5932 12718 5964
rect 12686 5864 12718 5896
rect 12686 5796 12718 5828
rect 12686 5728 12718 5760
rect 12686 5660 12718 5692
rect 12686 5592 12718 5624
rect 12686 5524 12718 5556
rect 12686 5456 12718 5488
rect 12686 5388 12718 5420
rect 12686 5320 12718 5352
rect 12686 5252 12718 5284
rect 3282 5184 3314 5216
rect 3282 5116 3314 5148
rect 3282 5048 3314 5080
rect 3282 4980 3314 5012
rect 12686 5184 12718 5216
rect 12686 5116 12718 5148
rect 12686 5048 12718 5080
rect 12686 4980 12718 5012
rect 3292 4892 3324 4924
rect 3360 4892 3392 4924
rect 3428 4892 3460 4924
rect 3496 4892 3528 4924
rect 3564 4892 3596 4924
rect 3632 4892 3664 4924
rect 3700 4892 3732 4924
rect 3768 4892 3800 4924
rect 3836 4892 3868 4924
rect 3904 4892 3936 4924
rect 3972 4892 4004 4924
rect 4040 4892 4072 4924
rect 4108 4892 4140 4924
rect 4176 4892 4208 4924
rect 4244 4892 4276 4924
rect 4312 4892 4344 4924
rect 4380 4892 4412 4924
rect 4448 4892 4480 4924
rect 4516 4892 4548 4924
rect 4584 4892 4616 4924
rect 4652 4892 4684 4924
rect 4720 4892 4752 4924
rect 4788 4892 4820 4924
rect 4856 4892 4888 4924
rect 4924 4892 4956 4924
rect 4992 4892 5024 4924
rect 5060 4892 5092 4924
rect 5128 4892 5160 4924
rect 5196 4892 5228 4924
rect 5264 4892 5296 4924
rect 5332 4892 5364 4924
rect 5400 4892 5432 4924
rect 5468 4892 5500 4924
rect 5536 4892 5568 4924
rect 5604 4892 5636 4924
rect 5672 4892 5704 4924
rect 5740 4892 5772 4924
rect 5808 4892 5840 4924
rect 5876 4892 5908 4924
rect 5944 4892 5976 4924
rect 6012 4892 6044 4924
rect 6080 4892 6112 4924
rect 6148 4892 6180 4924
rect 6216 4892 6248 4924
rect 6284 4892 6316 4924
rect 6352 4892 6384 4924
rect 6420 4892 6452 4924
rect 6488 4892 6520 4924
rect 6556 4892 6588 4924
rect 6624 4892 6656 4924
rect 6692 4892 6724 4924
rect 6760 4892 6792 4924
rect 6828 4892 6860 4924
rect 6896 4892 6928 4924
rect 6964 4892 6996 4924
rect 7032 4892 7064 4924
rect 7100 4892 7132 4924
rect 7168 4892 7200 4924
rect 7236 4892 7268 4924
rect 7304 4892 7336 4924
rect 7372 4892 7404 4924
rect 7440 4892 7472 4924
rect 7508 4892 7540 4924
rect 7576 4892 7608 4924
rect 7644 4892 7676 4924
rect 7712 4892 7744 4924
rect 7780 4892 7812 4924
rect 7848 4892 7880 4924
rect 7916 4892 7948 4924
rect 7984 4892 8016 4924
rect 8052 4892 8084 4924
rect 8120 4892 8152 4924
rect 8188 4892 8220 4924
rect 8256 4892 8288 4924
rect 8324 4892 8356 4924
rect 8392 4892 8424 4924
rect 8460 4892 8492 4924
rect 8528 4892 8560 4924
rect 8596 4892 8628 4924
rect 8664 4892 8696 4924
rect 8732 4892 8764 4924
rect 8800 4892 8832 4924
rect 8868 4892 8900 4924
rect 8936 4892 8968 4924
rect 9004 4892 9036 4924
rect 9072 4892 9104 4924
rect 9140 4892 9172 4924
rect 9208 4892 9240 4924
rect 9276 4892 9308 4924
rect 9344 4892 9376 4924
rect 9412 4892 9444 4924
rect 9480 4892 9512 4924
rect 9548 4892 9580 4924
rect 9616 4892 9648 4924
rect 9684 4892 9716 4924
rect 9752 4892 9784 4924
rect 9820 4892 9852 4924
rect 9888 4892 9920 4924
rect 9956 4892 9988 4924
rect 10024 4892 10056 4924
rect 10092 4892 10124 4924
rect 10160 4892 10192 4924
rect 10228 4892 10260 4924
rect 10296 4892 10328 4924
rect 10364 4892 10396 4924
rect 10432 4892 10464 4924
rect 10500 4892 10532 4924
rect 10568 4892 10600 4924
rect 10636 4892 10668 4924
rect 10704 4892 10736 4924
rect 10772 4892 10804 4924
rect 10840 4892 10872 4924
rect 10908 4892 10940 4924
rect 10976 4892 11008 4924
rect 11044 4892 11076 4924
rect 11112 4892 11144 4924
rect 11180 4892 11212 4924
rect 11248 4892 11280 4924
rect 11316 4892 11348 4924
rect 11384 4892 11416 4924
rect 11452 4892 11484 4924
rect 11520 4892 11552 4924
rect 11588 4892 11620 4924
rect 11656 4892 11688 4924
rect 11724 4892 11756 4924
rect 11792 4892 11824 4924
rect 11860 4892 11892 4924
rect 11928 4892 11960 4924
rect 11996 4892 12028 4924
rect 12064 4892 12096 4924
rect 12132 4892 12164 4924
rect 12200 4892 12232 4924
rect 12268 4892 12300 4924
rect 12336 4892 12368 4924
rect 12404 4892 12436 4924
rect 12472 4892 12504 4924
rect 12540 4892 12572 4924
rect 12608 4892 12640 4924
rect 12676 4892 12708 4924
<< poly >>
rect 3638 6742 12362 6756
rect 3638 6710 3666 6742
rect 3698 6710 3734 6742
rect 3766 6710 3802 6742
rect 3834 6710 3870 6742
rect 3902 6710 3938 6742
rect 3970 6710 4006 6742
rect 4038 6710 4074 6742
rect 4106 6710 4142 6742
rect 4174 6710 4210 6742
rect 4242 6710 4278 6742
rect 4310 6710 4346 6742
rect 4378 6710 4414 6742
rect 4446 6710 4482 6742
rect 4514 6710 4550 6742
rect 4582 6710 4618 6742
rect 4650 6710 4686 6742
rect 4718 6710 4754 6742
rect 4786 6710 4822 6742
rect 4854 6710 4890 6742
rect 4922 6710 4958 6742
rect 4990 6710 5026 6742
rect 5058 6710 5094 6742
rect 5126 6710 5162 6742
rect 5194 6710 5230 6742
rect 5262 6710 5298 6742
rect 5330 6710 5366 6742
rect 5398 6710 5434 6742
rect 5466 6710 5502 6742
rect 5534 6710 5570 6742
rect 5602 6710 5638 6742
rect 5670 6710 5706 6742
rect 5738 6710 5774 6742
rect 5806 6710 5842 6742
rect 5874 6710 5910 6742
rect 5942 6710 5978 6742
rect 6010 6710 6046 6742
rect 6078 6710 6114 6742
rect 6146 6710 6182 6742
rect 6214 6710 6250 6742
rect 6282 6710 6318 6742
rect 6350 6710 6386 6742
rect 6418 6710 6454 6742
rect 6486 6710 6522 6742
rect 6554 6710 6590 6742
rect 6622 6710 6658 6742
rect 6690 6710 6726 6742
rect 6758 6710 6794 6742
rect 6826 6710 6862 6742
rect 6894 6710 6930 6742
rect 6962 6710 6998 6742
rect 7030 6710 7066 6742
rect 7098 6710 7134 6742
rect 7166 6710 7202 6742
rect 7234 6710 7270 6742
rect 7302 6710 7338 6742
rect 7370 6710 7406 6742
rect 7438 6710 7474 6742
rect 7506 6710 7542 6742
rect 7574 6710 7610 6742
rect 7642 6710 7678 6742
rect 7710 6710 7746 6742
rect 7778 6710 7814 6742
rect 7846 6710 7882 6742
rect 7914 6710 7950 6742
rect 7982 6710 8018 6742
rect 8050 6710 8086 6742
rect 8118 6710 8154 6742
rect 8186 6710 8222 6742
rect 8254 6710 8290 6742
rect 8322 6710 8358 6742
rect 8390 6710 8426 6742
rect 8458 6710 8494 6742
rect 8526 6710 8562 6742
rect 8594 6710 8630 6742
rect 8662 6710 8698 6742
rect 8730 6710 8766 6742
rect 8798 6710 8834 6742
rect 8866 6710 8902 6742
rect 8934 6710 8970 6742
rect 9002 6710 9038 6742
rect 9070 6710 9106 6742
rect 9138 6710 9174 6742
rect 9206 6710 9242 6742
rect 9274 6710 9310 6742
rect 9342 6710 9378 6742
rect 9410 6710 9446 6742
rect 9478 6710 9514 6742
rect 9546 6710 9582 6742
rect 9614 6710 9650 6742
rect 9682 6710 9718 6742
rect 9750 6710 9786 6742
rect 9818 6710 9854 6742
rect 9886 6710 9922 6742
rect 9954 6710 9990 6742
rect 10022 6710 10058 6742
rect 10090 6710 10126 6742
rect 10158 6710 10194 6742
rect 10226 6710 10262 6742
rect 10294 6710 10330 6742
rect 10362 6710 10398 6742
rect 10430 6710 10466 6742
rect 10498 6710 10534 6742
rect 10566 6710 10602 6742
rect 10634 6710 10670 6742
rect 10702 6710 10738 6742
rect 10770 6710 10806 6742
rect 10838 6710 10874 6742
rect 10906 6710 10942 6742
rect 10974 6710 11010 6742
rect 11042 6710 11078 6742
rect 11110 6710 11146 6742
rect 11178 6710 11214 6742
rect 11246 6710 11282 6742
rect 11314 6710 11350 6742
rect 11382 6710 11418 6742
rect 11450 6710 11486 6742
rect 11518 6710 11554 6742
rect 11586 6710 11622 6742
rect 11654 6710 11690 6742
rect 11722 6710 11758 6742
rect 11790 6710 11826 6742
rect 11858 6710 11894 6742
rect 11926 6710 11962 6742
rect 11994 6710 12030 6742
rect 12062 6710 12098 6742
rect 12130 6710 12166 6742
rect 12198 6710 12234 6742
rect 12266 6710 12302 6742
rect 12334 6710 12362 6742
rect 3638 6696 12362 6710
rect 3638 6682 3738 6696
rect 3814 6682 3914 6696
rect 3990 6682 4090 6696
rect 4166 6682 4266 6696
rect 4342 6682 4442 6696
rect 4518 6682 4618 6696
rect 4694 6682 4794 6696
rect 4870 6682 4970 6696
rect 5046 6682 5146 6696
rect 5222 6682 5322 6696
rect 5398 6682 5498 6696
rect 5574 6682 5674 6696
rect 5750 6682 5850 6696
rect 5926 6682 6026 6696
rect 6102 6682 6202 6696
rect 6278 6682 6378 6696
rect 6454 6682 6554 6696
rect 6630 6682 6730 6696
rect 6806 6682 6906 6696
rect 6982 6682 7082 6696
rect 7158 6682 7258 6696
rect 7334 6682 7434 6696
rect 7510 6682 7610 6696
rect 7686 6682 7786 6696
rect 7862 6682 7962 6696
rect 8038 6682 8138 6696
rect 8214 6682 8314 6696
rect 8390 6682 8490 6696
rect 8566 6682 8666 6696
rect 8742 6682 8842 6696
rect 8918 6682 9018 6696
rect 9094 6682 9194 6696
rect 9270 6682 9370 6696
rect 9446 6682 9546 6696
rect 9622 6682 9722 6696
rect 9798 6682 9898 6696
rect 9974 6682 10074 6696
rect 10150 6682 10250 6696
rect 10326 6682 10426 6696
rect 10502 6682 10602 6696
rect 10678 6682 10778 6696
rect 10854 6682 10954 6696
rect 11030 6682 11130 6696
rect 11206 6682 11306 6696
rect 11382 6682 11482 6696
rect 11558 6682 11658 6696
rect 11734 6682 11834 6696
rect 11910 6682 12010 6696
rect 12086 6682 12186 6696
rect 12262 6682 12362 6696
rect 3638 5246 3738 5282
rect 3814 5246 3914 5282
rect 3990 5246 4090 5282
rect 4166 5246 4266 5282
rect 4342 5246 4442 5282
rect 4518 5246 4618 5282
rect 4694 5246 4794 5282
rect 4870 5246 4970 5282
rect 5046 5246 5146 5282
rect 5222 5246 5322 5282
rect 5398 5246 5498 5282
rect 5574 5246 5674 5282
rect 5750 5246 5850 5282
rect 5926 5246 6026 5282
rect 6102 5246 6202 5282
rect 6278 5246 6378 5282
rect 6454 5246 6554 5282
rect 6630 5246 6730 5282
rect 6806 5246 6906 5282
rect 6982 5246 7082 5282
rect 7158 5246 7258 5282
rect 7334 5246 7434 5282
rect 7510 5246 7610 5282
rect 7686 5246 7786 5282
rect 7862 5246 7962 5282
rect 8038 5246 8138 5282
rect 8214 5246 8314 5282
rect 8390 5246 8490 5282
rect 8566 5246 8666 5282
rect 8742 5246 8842 5282
rect 8918 5246 9018 5282
rect 9094 5246 9194 5282
rect 9270 5246 9370 5282
rect 9446 5246 9546 5282
rect 9622 5246 9722 5282
rect 9798 5246 9898 5282
rect 9974 5246 10074 5282
rect 10150 5246 10250 5282
rect 10326 5246 10426 5282
rect 10502 5246 10602 5282
rect 10678 5246 10778 5282
rect 10854 5246 10954 5282
rect 11030 5246 11130 5282
rect 11206 5246 11306 5282
rect 11382 5246 11482 5282
rect 11558 5246 11658 5282
rect 11734 5246 11834 5282
rect 11910 5246 12010 5282
rect 12086 5246 12186 5282
rect 12262 5246 12362 5282
rect 594 4058 2494 4094
rect 2570 4058 4470 4094
rect 4546 4058 6446 4094
rect 6522 4058 8422 4094
rect 8498 4058 10398 4094
rect 10474 4058 12374 4094
rect 12450 4058 14350 4094
rect 14426 4058 14526 4094
rect 14602 4058 14702 4094
rect 14778 4058 14878 4094
rect 14954 4058 15054 4094
rect 15130 4058 15230 4094
rect 15306 4058 15406 4094
rect 594 2208 2494 2258
rect 2570 2208 4470 2258
rect 4546 2208 6446 2258
rect 6522 2208 8422 2258
rect 8498 2208 10398 2258
rect 10474 2208 12374 2258
rect 12450 2208 14350 2258
rect 14426 2208 14526 2258
rect 14602 2208 14702 2258
rect 14778 2208 14878 2258
rect 14954 2208 15054 2258
rect 15130 2208 15230 2258
rect 15306 2208 15406 2258
rect 594 394 2494 408
rect 2570 394 4470 408
rect 4546 394 6446 408
rect 6522 394 8422 408
rect 8498 394 10398 408
rect 10474 394 12374 408
rect 12450 394 14350 408
rect 14426 394 14526 408
rect 14602 394 14702 408
rect 14778 394 14878 408
rect 14954 394 15054 408
rect 15130 394 15230 408
rect 15306 394 15406 408
rect 594 380 15406 394
rect 594 348 640 380
rect 672 348 708 380
rect 740 348 776 380
rect 808 348 844 380
rect 876 348 912 380
rect 944 348 980 380
rect 1012 348 1048 380
rect 1080 348 1116 380
rect 1148 348 1184 380
rect 1216 348 1252 380
rect 1284 348 1320 380
rect 1352 348 1388 380
rect 1420 348 1456 380
rect 1488 348 1524 380
rect 1556 348 1592 380
rect 1624 348 1660 380
rect 1692 348 1728 380
rect 1760 348 1796 380
rect 1828 348 1864 380
rect 1896 348 1932 380
rect 1964 348 2000 380
rect 2032 348 2068 380
rect 2100 348 2136 380
rect 2168 348 2204 380
rect 2236 348 2272 380
rect 2304 348 2340 380
rect 2372 348 2408 380
rect 2440 348 2476 380
rect 2508 348 2544 380
rect 2576 348 2612 380
rect 2644 348 2680 380
rect 2712 348 2748 380
rect 2780 348 2816 380
rect 2848 348 2884 380
rect 2916 348 2952 380
rect 2984 348 3020 380
rect 3052 348 3088 380
rect 3120 348 3156 380
rect 3188 348 3224 380
rect 3256 348 3292 380
rect 3324 348 3360 380
rect 3392 348 3428 380
rect 3460 348 3496 380
rect 3528 348 3564 380
rect 3596 348 3632 380
rect 3664 348 3700 380
rect 3732 348 3768 380
rect 3800 348 3836 380
rect 3868 348 3904 380
rect 3936 348 3972 380
rect 4004 348 4040 380
rect 4072 348 4108 380
rect 4140 348 4176 380
rect 4208 348 4244 380
rect 4276 348 4312 380
rect 4344 348 4380 380
rect 4412 348 4448 380
rect 4480 348 4516 380
rect 4548 348 4584 380
rect 4616 348 4652 380
rect 4684 348 4720 380
rect 4752 348 4788 380
rect 4820 348 4856 380
rect 4888 348 4924 380
rect 4956 348 4992 380
rect 5024 348 5060 380
rect 5092 348 5128 380
rect 5160 348 5196 380
rect 5228 348 5264 380
rect 5296 348 5332 380
rect 5364 348 5400 380
rect 5432 348 5468 380
rect 5500 348 5536 380
rect 5568 348 5604 380
rect 5636 348 5672 380
rect 5704 348 5740 380
rect 5772 348 5808 380
rect 5840 348 5876 380
rect 5908 348 5944 380
rect 5976 348 6012 380
rect 6044 348 6080 380
rect 6112 348 6148 380
rect 6180 348 6216 380
rect 6248 348 6284 380
rect 6316 348 6352 380
rect 6384 348 6420 380
rect 6452 348 6488 380
rect 6520 348 6556 380
rect 6588 348 6624 380
rect 6656 348 6692 380
rect 6724 348 6760 380
rect 6792 348 6828 380
rect 6860 348 6896 380
rect 6928 348 6964 380
rect 6996 348 7032 380
rect 7064 348 7100 380
rect 7132 348 7168 380
rect 7200 348 7236 380
rect 7268 348 7304 380
rect 7336 348 7372 380
rect 7404 348 7440 380
rect 7472 348 7508 380
rect 7540 348 7576 380
rect 7608 348 7644 380
rect 7676 348 7712 380
rect 7744 348 7780 380
rect 7812 348 7848 380
rect 7880 348 7916 380
rect 7948 348 7984 380
rect 8016 348 8052 380
rect 8084 348 8120 380
rect 8152 348 8188 380
rect 8220 348 8256 380
rect 8288 348 8324 380
rect 8356 348 8392 380
rect 8424 348 8460 380
rect 8492 348 8528 380
rect 8560 348 8596 380
rect 8628 348 8664 380
rect 8696 348 8732 380
rect 8764 348 8800 380
rect 8832 348 8868 380
rect 8900 348 8936 380
rect 8968 348 9004 380
rect 9036 348 9072 380
rect 9104 348 9140 380
rect 9172 348 9208 380
rect 9240 348 9276 380
rect 9308 348 9344 380
rect 9376 348 9412 380
rect 9444 348 9480 380
rect 9512 348 9548 380
rect 9580 348 9616 380
rect 9648 348 9684 380
rect 9716 348 9752 380
rect 9784 348 9820 380
rect 9852 348 9888 380
rect 9920 348 9956 380
rect 9988 348 10024 380
rect 10056 348 10092 380
rect 10124 348 10160 380
rect 10192 348 10228 380
rect 10260 348 10296 380
rect 10328 348 10364 380
rect 10396 348 10432 380
rect 10464 348 10500 380
rect 10532 348 10568 380
rect 10600 348 10636 380
rect 10668 348 10704 380
rect 10736 348 10772 380
rect 10804 348 10840 380
rect 10872 348 10908 380
rect 10940 348 10976 380
rect 11008 348 11044 380
rect 11076 348 11112 380
rect 11144 348 11180 380
rect 11212 348 11248 380
rect 11280 348 11316 380
rect 11348 348 11384 380
rect 11416 348 11452 380
rect 11484 348 11520 380
rect 11552 348 11588 380
rect 11620 348 11656 380
rect 11688 348 11724 380
rect 11756 348 11792 380
rect 11824 348 11860 380
rect 11892 348 11928 380
rect 11960 348 11996 380
rect 12028 348 12064 380
rect 12096 348 12132 380
rect 12164 348 12200 380
rect 12232 348 12268 380
rect 12300 348 12336 380
rect 12368 348 12404 380
rect 12436 348 12472 380
rect 12504 348 12540 380
rect 12572 348 12608 380
rect 12640 348 12676 380
rect 12708 348 12744 380
rect 12776 348 12812 380
rect 12844 348 12880 380
rect 12912 348 12948 380
rect 12980 348 13016 380
rect 13048 348 13084 380
rect 13116 348 13152 380
rect 13184 348 13220 380
rect 13252 348 13288 380
rect 13320 348 13356 380
rect 13388 348 13424 380
rect 13456 348 13492 380
rect 13524 348 13560 380
rect 13592 348 13628 380
rect 13660 348 13696 380
rect 13728 348 13764 380
rect 13796 348 13832 380
rect 13864 348 13900 380
rect 13932 348 13968 380
rect 14000 348 14036 380
rect 14068 348 14104 380
rect 14136 348 14172 380
rect 14204 348 14240 380
rect 14272 348 14308 380
rect 14340 348 14376 380
rect 14408 348 14444 380
rect 14476 348 14512 380
rect 14544 348 14580 380
rect 14612 348 14648 380
rect 14680 348 14716 380
rect 14748 348 14784 380
rect 14816 348 14852 380
rect 14884 348 14920 380
rect 14952 348 14988 380
rect 15020 348 15056 380
rect 15088 348 15124 380
rect 15156 348 15192 380
rect 15224 348 15260 380
rect 15292 348 15328 380
rect 15360 348 15406 380
rect 594 334 15406 348
<< polycont >>
rect 3666 6710 3698 6742
rect 3734 6710 3766 6742
rect 3802 6710 3834 6742
rect 3870 6710 3902 6742
rect 3938 6710 3970 6742
rect 4006 6710 4038 6742
rect 4074 6710 4106 6742
rect 4142 6710 4174 6742
rect 4210 6710 4242 6742
rect 4278 6710 4310 6742
rect 4346 6710 4378 6742
rect 4414 6710 4446 6742
rect 4482 6710 4514 6742
rect 4550 6710 4582 6742
rect 4618 6710 4650 6742
rect 4686 6710 4718 6742
rect 4754 6710 4786 6742
rect 4822 6710 4854 6742
rect 4890 6710 4922 6742
rect 4958 6710 4990 6742
rect 5026 6710 5058 6742
rect 5094 6710 5126 6742
rect 5162 6710 5194 6742
rect 5230 6710 5262 6742
rect 5298 6710 5330 6742
rect 5366 6710 5398 6742
rect 5434 6710 5466 6742
rect 5502 6710 5534 6742
rect 5570 6710 5602 6742
rect 5638 6710 5670 6742
rect 5706 6710 5738 6742
rect 5774 6710 5806 6742
rect 5842 6710 5874 6742
rect 5910 6710 5942 6742
rect 5978 6710 6010 6742
rect 6046 6710 6078 6742
rect 6114 6710 6146 6742
rect 6182 6710 6214 6742
rect 6250 6710 6282 6742
rect 6318 6710 6350 6742
rect 6386 6710 6418 6742
rect 6454 6710 6486 6742
rect 6522 6710 6554 6742
rect 6590 6710 6622 6742
rect 6658 6710 6690 6742
rect 6726 6710 6758 6742
rect 6794 6710 6826 6742
rect 6862 6710 6894 6742
rect 6930 6710 6962 6742
rect 6998 6710 7030 6742
rect 7066 6710 7098 6742
rect 7134 6710 7166 6742
rect 7202 6710 7234 6742
rect 7270 6710 7302 6742
rect 7338 6710 7370 6742
rect 7406 6710 7438 6742
rect 7474 6710 7506 6742
rect 7542 6710 7574 6742
rect 7610 6710 7642 6742
rect 7678 6710 7710 6742
rect 7746 6710 7778 6742
rect 7814 6710 7846 6742
rect 7882 6710 7914 6742
rect 7950 6710 7982 6742
rect 8018 6710 8050 6742
rect 8086 6710 8118 6742
rect 8154 6710 8186 6742
rect 8222 6710 8254 6742
rect 8290 6710 8322 6742
rect 8358 6710 8390 6742
rect 8426 6710 8458 6742
rect 8494 6710 8526 6742
rect 8562 6710 8594 6742
rect 8630 6710 8662 6742
rect 8698 6710 8730 6742
rect 8766 6710 8798 6742
rect 8834 6710 8866 6742
rect 8902 6710 8934 6742
rect 8970 6710 9002 6742
rect 9038 6710 9070 6742
rect 9106 6710 9138 6742
rect 9174 6710 9206 6742
rect 9242 6710 9274 6742
rect 9310 6710 9342 6742
rect 9378 6710 9410 6742
rect 9446 6710 9478 6742
rect 9514 6710 9546 6742
rect 9582 6710 9614 6742
rect 9650 6710 9682 6742
rect 9718 6710 9750 6742
rect 9786 6710 9818 6742
rect 9854 6710 9886 6742
rect 9922 6710 9954 6742
rect 9990 6710 10022 6742
rect 10058 6710 10090 6742
rect 10126 6710 10158 6742
rect 10194 6710 10226 6742
rect 10262 6710 10294 6742
rect 10330 6710 10362 6742
rect 10398 6710 10430 6742
rect 10466 6710 10498 6742
rect 10534 6710 10566 6742
rect 10602 6710 10634 6742
rect 10670 6710 10702 6742
rect 10738 6710 10770 6742
rect 10806 6710 10838 6742
rect 10874 6710 10906 6742
rect 10942 6710 10974 6742
rect 11010 6710 11042 6742
rect 11078 6710 11110 6742
rect 11146 6710 11178 6742
rect 11214 6710 11246 6742
rect 11282 6710 11314 6742
rect 11350 6710 11382 6742
rect 11418 6710 11450 6742
rect 11486 6710 11518 6742
rect 11554 6710 11586 6742
rect 11622 6710 11654 6742
rect 11690 6710 11722 6742
rect 11758 6710 11790 6742
rect 11826 6710 11858 6742
rect 11894 6710 11926 6742
rect 11962 6710 11994 6742
rect 12030 6710 12062 6742
rect 12098 6710 12130 6742
rect 12166 6710 12198 6742
rect 12234 6710 12266 6742
rect 12302 6710 12334 6742
rect 640 348 672 380
rect 708 348 740 380
rect 776 348 808 380
rect 844 348 876 380
rect 912 348 944 380
rect 980 348 1012 380
rect 1048 348 1080 380
rect 1116 348 1148 380
rect 1184 348 1216 380
rect 1252 348 1284 380
rect 1320 348 1352 380
rect 1388 348 1420 380
rect 1456 348 1488 380
rect 1524 348 1556 380
rect 1592 348 1624 380
rect 1660 348 1692 380
rect 1728 348 1760 380
rect 1796 348 1828 380
rect 1864 348 1896 380
rect 1932 348 1964 380
rect 2000 348 2032 380
rect 2068 348 2100 380
rect 2136 348 2168 380
rect 2204 348 2236 380
rect 2272 348 2304 380
rect 2340 348 2372 380
rect 2408 348 2440 380
rect 2476 348 2508 380
rect 2544 348 2576 380
rect 2612 348 2644 380
rect 2680 348 2712 380
rect 2748 348 2780 380
rect 2816 348 2848 380
rect 2884 348 2916 380
rect 2952 348 2984 380
rect 3020 348 3052 380
rect 3088 348 3120 380
rect 3156 348 3188 380
rect 3224 348 3256 380
rect 3292 348 3324 380
rect 3360 348 3392 380
rect 3428 348 3460 380
rect 3496 348 3528 380
rect 3564 348 3596 380
rect 3632 348 3664 380
rect 3700 348 3732 380
rect 3768 348 3800 380
rect 3836 348 3868 380
rect 3904 348 3936 380
rect 3972 348 4004 380
rect 4040 348 4072 380
rect 4108 348 4140 380
rect 4176 348 4208 380
rect 4244 348 4276 380
rect 4312 348 4344 380
rect 4380 348 4412 380
rect 4448 348 4480 380
rect 4516 348 4548 380
rect 4584 348 4616 380
rect 4652 348 4684 380
rect 4720 348 4752 380
rect 4788 348 4820 380
rect 4856 348 4888 380
rect 4924 348 4956 380
rect 4992 348 5024 380
rect 5060 348 5092 380
rect 5128 348 5160 380
rect 5196 348 5228 380
rect 5264 348 5296 380
rect 5332 348 5364 380
rect 5400 348 5432 380
rect 5468 348 5500 380
rect 5536 348 5568 380
rect 5604 348 5636 380
rect 5672 348 5704 380
rect 5740 348 5772 380
rect 5808 348 5840 380
rect 5876 348 5908 380
rect 5944 348 5976 380
rect 6012 348 6044 380
rect 6080 348 6112 380
rect 6148 348 6180 380
rect 6216 348 6248 380
rect 6284 348 6316 380
rect 6352 348 6384 380
rect 6420 348 6452 380
rect 6488 348 6520 380
rect 6556 348 6588 380
rect 6624 348 6656 380
rect 6692 348 6724 380
rect 6760 348 6792 380
rect 6828 348 6860 380
rect 6896 348 6928 380
rect 6964 348 6996 380
rect 7032 348 7064 380
rect 7100 348 7132 380
rect 7168 348 7200 380
rect 7236 348 7268 380
rect 7304 348 7336 380
rect 7372 348 7404 380
rect 7440 348 7472 380
rect 7508 348 7540 380
rect 7576 348 7608 380
rect 7644 348 7676 380
rect 7712 348 7744 380
rect 7780 348 7812 380
rect 7848 348 7880 380
rect 7916 348 7948 380
rect 7984 348 8016 380
rect 8052 348 8084 380
rect 8120 348 8152 380
rect 8188 348 8220 380
rect 8256 348 8288 380
rect 8324 348 8356 380
rect 8392 348 8424 380
rect 8460 348 8492 380
rect 8528 348 8560 380
rect 8596 348 8628 380
rect 8664 348 8696 380
rect 8732 348 8764 380
rect 8800 348 8832 380
rect 8868 348 8900 380
rect 8936 348 8968 380
rect 9004 348 9036 380
rect 9072 348 9104 380
rect 9140 348 9172 380
rect 9208 348 9240 380
rect 9276 348 9308 380
rect 9344 348 9376 380
rect 9412 348 9444 380
rect 9480 348 9512 380
rect 9548 348 9580 380
rect 9616 348 9648 380
rect 9684 348 9716 380
rect 9752 348 9784 380
rect 9820 348 9852 380
rect 9888 348 9920 380
rect 9956 348 9988 380
rect 10024 348 10056 380
rect 10092 348 10124 380
rect 10160 348 10192 380
rect 10228 348 10260 380
rect 10296 348 10328 380
rect 10364 348 10396 380
rect 10432 348 10464 380
rect 10500 348 10532 380
rect 10568 348 10600 380
rect 10636 348 10668 380
rect 10704 348 10736 380
rect 10772 348 10804 380
rect 10840 348 10872 380
rect 10908 348 10940 380
rect 10976 348 11008 380
rect 11044 348 11076 380
rect 11112 348 11144 380
rect 11180 348 11212 380
rect 11248 348 11280 380
rect 11316 348 11348 380
rect 11384 348 11416 380
rect 11452 348 11484 380
rect 11520 348 11552 380
rect 11588 348 11620 380
rect 11656 348 11688 380
rect 11724 348 11756 380
rect 11792 348 11824 380
rect 11860 348 11892 380
rect 11928 348 11960 380
rect 11996 348 12028 380
rect 12064 348 12096 380
rect 12132 348 12164 380
rect 12200 348 12232 380
rect 12268 348 12300 380
rect 12336 348 12368 380
rect 12404 348 12436 380
rect 12472 348 12504 380
rect 12540 348 12572 380
rect 12608 348 12640 380
rect 12676 348 12708 380
rect 12744 348 12776 380
rect 12812 348 12844 380
rect 12880 348 12912 380
rect 12948 348 12980 380
rect 13016 348 13048 380
rect 13084 348 13116 380
rect 13152 348 13184 380
rect 13220 348 13252 380
rect 13288 348 13320 380
rect 13356 348 13388 380
rect 13424 348 13456 380
rect 13492 348 13524 380
rect 13560 348 13592 380
rect 13628 348 13660 380
rect 13696 348 13728 380
rect 13764 348 13796 380
rect 13832 348 13864 380
rect 13900 348 13932 380
rect 13968 348 14000 380
rect 14036 348 14068 380
rect 14104 348 14136 380
rect 14172 348 14204 380
rect 14240 348 14272 380
rect 14308 348 14340 380
rect 14376 348 14408 380
rect 14444 348 14476 380
rect 14512 348 14544 380
rect 14580 348 14612 380
rect 14648 348 14680 380
rect 14716 348 14748 380
rect 14784 348 14816 380
rect 14852 348 14884 380
rect 14920 348 14952 380
rect 14988 348 15020 380
rect 15056 348 15088 380
rect 15124 348 15156 380
rect 15192 348 15224 380
rect 15260 348 15292 380
rect 15328 348 15360 380
<< metal1 >>
rect 3264 7072 12736 7090
rect 3264 7040 3292 7072
rect 3324 7040 3360 7072
rect 3392 7040 3428 7072
rect 3460 7040 3496 7072
rect 3528 7040 3564 7072
rect 3596 7040 3632 7072
rect 3664 7040 3700 7072
rect 3732 7040 3768 7072
rect 3800 7040 3836 7072
rect 3868 7040 3904 7072
rect 3936 7040 3972 7072
rect 4004 7040 4040 7072
rect 4072 7040 4108 7072
rect 4140 7040 4176 7072
rect 4208 7040 4244 7072
rect 4276 7040 4312 7072
rect 4344 7040 4380 7072
rect 4412 7040 4448 7072
rect 4480 7040 4516 7072
rect 4548 7040 4584 7072
rect 4616 7040 4652 7072
rect 4684 7040 4720 7072
rect 4752 7040 4788 7072
rect 4820 7040 4856 7072
rect 4888 7040 4924 7072
rect 4956 7040 4992 7072
rect 5024 7040 5060 7072
rect 5092 7040 5128 7072
rect 5160 7040 5196 7072
rect 5228 7040 5264 7072
rect 5296 7040 5332 7072
rect 5364 7040 5400 7072
rect 5432 7040 5468 7072
rect 5500 7040 5536 7072
rect 5568 7040 5604 7072
rect 5636 7040 5672 7072
rect 5704 7040 5740 7072
rect 5772 7040 5808 7072
rect 5840 7040 5876 7072
rect 5908 7040 5944 7072
rect 5976 7040 6012 7072
rect 6044 7040 6080 7072
rect 6112 7040 6148 7072
rect 6180 7040 6216 7072
rect 6248 7040 6284 7072
rect 6316 7040 6352 7072
rect 6384 7040 6420 7072
rect 6452 7040 6488 7072
rect 6520 7040 6556 7072
rect 6588 7040 6624 7072
rect 6656 7040 6692 7072
rect 6724 7040 6760 7072
rect 6792 7040 6828 7072
rect 6860 7040 6896 7072
rect 6928 7040 6964 7072
rect 6996 7040 7032 7072
rect 7064 7040 7100 7072
rect 7132 7040 7168 7072
rect 7200 7040 7236 7072
rect 7268 7040 7304 7072
rect 7336 7040 7372 7072
rect 7404 7040 7440 7072
rect 7472 7040 7508 7072
rect 7540 7040 7576 7072
rect 7608 7040 7644 7072
rect 7676 7040 7712 7072
rect 7744 7040 7780 7072
rect 7812 7040 7848 7072
rect 7880 7040 7916 7072
rect 7948 7040 7984 7072
rect 8016 7040 8052 7072
rect 8084 7040 8120 7072
rect 8152 7040 8188 7072
rect 8220 7040 8256 7072
rect 8288 7040 8324 7072
rect 8356 7040 8392 7072
rect 8424 7040 8460 7072
rect 8492 7040 8528 7072
rect 8560 7040 8596 7072
rect 8628 7040 8664 7072
rect 8696 7040 8732 7072
rect 8764 7040 8800 7072
rect 8832 7040 8868 7072
rect 8900 7040 8936 7072
rect 8968 7040 9004 7072
rect 9036 7040 9072 7072
rect 9104 7040 9140 7072
rect 9172 7040 9208 7072
rect 9240 7040 9276 7072
rect 9308 7040 9344 7072
rect 9376 7040 9412 7072
rect 9444 7040 9480 7072
rect 9512 7040 9548 7072
rect 9580 7040 9616 7072
rect 9648 7040 9684 7072
rect 9716 7040 9752 7072
rect 9784 7040 9820 7072
rect 9852 7040 9888 7072
rect 9920 7040 9956 7072
rect 9988 7040 10024 7072
rect 10056 7040 10092 7072
rect 10124 7040 10160 7072
rect 10192 7040 10228 7072
rect 10260 7040 10296 7072
rect 10328 7040 10364 7072
rect 10396 7040 10432 7072
rect 10464 7040 10500 7072
rect 10532 7040 10568 7072
rect 10600 7040 10636 7072
rect 10668 7040 10704 7072
rect 10736 7040 10772 7072
rect 10804 7040 10840 7072
rect 10872 7040 10908 7072
rect 10940 7040 10976 7072
rect 11008 7040 11044 7072
rect 11076 7040 11112 7072
rect 11144 7040 11180 7072
rect 11212 7040 11248 7072
rect 11280 7040 11316 7072
rect 11348 7040 11384 7072
rect 11416 7040 11452 7072
rect 11484 7040 11520 7072
rect 11552 7040 11588 7072
rect 11620 7040 11656 7072
rect 11688 7040 11724 7072
rect 11756 7040 11792 7072
rect 11824 7040 11860 7072
rect 11892 7040 11928 7072
rect 11960 7040 11996 7072
rect 12028 7040 12064 7072
rect 12096 7040 12132 7072
rect 12164 7040 12200 7072
rect 12232 7040 12268 7072
rect 12300 7040 12336 7072
rect 12368 7040 12404 7072
rect 12436 7040 12472 7072
rect 12504 7040 12540 7072
rect 12572 7040 12608 7072
rect 12640 7040 12676 7072
rect 12708 7040 12736 7072
rect 3264 7022 12736 7040
rect 3264 6984 3332 7022
rect 3264 6952 3282 6984
rect 3314 6952 3332 6984
rect 3264 6916 3332 6952
rect 3264 6884 3282 6916
rect 3314 6884 3332 6916
rect 3264 6848 3332 6884
rect 3264 6816 3282 6848
rect 3314 6816 3332 6848
rect 3264 6780 3332 6816
rect 12668 6984 12736 7022
rect 12668 6952 12686 6984
rect 12718 6952 12736 6984
rect 12668 6916 12736 6952
rect 12668 6884 12686 6916
rect 12718 6884 12736 6916
rect 12668 6848 12736 6884
rect 12668 6816 12686 6848
rect 12718 6816 12736 6848
rect 3264 6748 3282 6780
rect 3314 6748 3332 6780
rect 3264 6712 3332 6748
rect 3264 6680 3282 6712
rect 3314 6680 3332 6712
rect 3638 6784 12362 6785
rect 3638 6744 3675 6784
rect 12325 6744 12362 6784
rect 3638 6742 12362 6744
rect 3638 6710 3666 6742
rect 3698 6710 3734 6742
rect 3766 6710 3802 6742
rect 3834 6710 3870 6742
rect 3902 6710 3938 6742
rect 3970 6710 4006 6742
rect 4038 6710 4074 6742
rect 4106 6710 4142 6742
rect 4174 6710 4210 6742
rect 4242 6710 4278 6742
rect 4310 6710 4346 6742
rect 4378 6710 4414 6742
rect 4446 6710 4482 6742
rect 4514 6710 4550 6742
rect 4582 6710 4618 6742
rect 4650 6710 4686 6742
rect 4718 6710 4754 6742
rect 4786 6710 4822 6742
rect 4854 6710 4890 6742
rect 4922 6710 4958 6742
rect 4990 6710 5026 6742
rect 5058 6710 5094 6742
rect 5126 6710 5162 6742
rect 5194 6710 5230 6742
rect 5262 6710 5298 6742
rect 5330 6710 5366 6742
rect 5398 6710 5434 6742
rect 5466 6710 5502 6742
rect 5534 6710 5570 6742
rect 5602 6710 5638 6742
rect 5670 6710 5706 6742
rect 5738 6710 5774 6742
rect 5806 6710 5842 6742
rect 5874 6710 5910 6742
rect 5942 6710 5978 6742
rect 6010 6710 6046 6742
rect 6078 6710 6114 6742
rect 6146 6710 6182 6742
rect 6214 6710 6250 6742
rect 6282 6710 6318 6742
rect 6350 6710 6386 6742
rect 6418 6710 6454 6742
rect 6486 6710 6522 6742
rect 6554 6710 6590 6742
rect 6622 6710 6658 6742
rect 6690 6710 6726 6742
rect 6758 6710 6794 6742
rect 6826 6710 6862 6742
rect 6894 6710 6930 6742
rect 6962 6710 6998 6742
rect 7030 6710 7066 6742
rect 7098 6710 7134 6742
rect 7166 6710 7202 6742
rect 7234 6710 7270 6742
rect 7302 6710 7338 6742
rect 7370 6710 7406 6742
rect 7438 6710 7474 6742
rect 7506 6710 7542 6742
rect 7574 6710 7610 6742
rect 7642 6710 7678 6742
rect 7710 6710 7746 6742
rect 7778 6710 7814 6742
rect 7846 6710 7882 6742
rect 7914 6710 7950 6742
rect 7982 6710 8018 6742
rect 8050 6710 8086 6742
rect 8118 6710 8154 6742
rect 8186 6710 8222 6742
rect 8254 6710 8290 6742
rect 8322 6710 8358 6742
rect 8390 6710 8426 6742
rect 8458 6710 8494 6742
rect 8526 6710 8562 6742
rect 8594 6710 8630 6742
rect 8662 6710 8698 6742
rect 8730 6710 8766 6742
rect 8798 6710 8834 6742
rect 8866 6710 8902 6742
rect 8934 6710 8970 6742
rect 9002 6710 9038 6742
rect 9070 6710 9106 6742
rect 9138 6710 9174 6742
rect 9206 6710 9242 6742
rect 9274 6710 9310 6742
rect 9342 6710 9378 6742
rect 9410 6710 9446 6742
rect 9478 6710 9514 6742
rect 9546 6710 9582 6742
rect 9614 6710 9650 6742
rect 9682 6710 9718 6742
rect 9750 6710 9786 6742
rect 9818 6710 9854 6742
rect 9886 6710 9922 6742
rect 9954 6710 9990 6742
rect 10022 6710 10058 6742
rect 10090 6710 10126 6742
rect 10158 6710 10194 6742
rect 10226 6710 10262 6742
rect 10294 6710 10330 6742
rect 10362 6710 10398 6742
rect 10430 6710 10466 6742
rect 10498 6710 10534 6742
rect 10566 6710 10602 6742
rect 10634 6710 10670 6742
rect 10702 6710 10738 6742
rect 10770 6710 10806 6742
rect 10838 6710 10874 6742
rect 10906 6710 10942 6742
rect 10974 6710 11010 6742
rect 11042 6710 11078 6742
rect 11110 6710 11146 6742
rect 11178 6710 11214 6742
rect 11246 6710 11282 6742
rect 11314 6710 11350 6742
rect 11382 6710 11418 6742
rect 11450 6710 11486 6742
rect 11518 6710 11554 6742
rect 11586 6710 11622 6742
rect 11654 6710 11690 6742
rect 11722 6710 11758 6742
rect 11790 6710 11826 6742
rect 11858 6710 11894 6742
rect 11926 6710 11962 6742
rect 11994 6710 12030 6742
rect 12062 6710 12098 6742
rect 12130 6710 12166 6742
rect 12198 6710 12234 6742
rect 12266 6710 12302 6742
rect 12334 6710 12362 6742
rect 12668 6780 12736 6816
rect 12668 6748 12686 6780
rect 12718 6748 12736 6780
rect 12668 6712 12736 6748
rect 3264 6644 3332 6680
rect 12668 6680 12686 6712
rect 12718 6680 12736 6712
rect 3264 6612 3282 6644
rect 3314 6612 3332 6644
rect 3264 6576 3332 6612
rect 3264 6544 3282 6576
rect 3314 6544 3332 6576
rect 3264 6508 3332 6544
rect 3264 6476 3282 6508
rect 3314 6476 3332 6508
rect 3264 6440 3332 6476
rect 3264 6408 3282 6440
rect 3314 6408 3332 6440
rect 3264 6372 3332 6408
rect 3264 6340 3282 6372
rect 3314 6340 3332 6372
rect 3264 6304 3332 6340
rect 3264 6272 3282 6304
rect 3314 6272 3332 6304
rect 3264 6236 3332 6272
rect 3264 6204 3282 6236
rect 3314 6204 3332 6236
rect 3264 6168 3332 6204
rect 3264 6136 3282 6168
rect 3314 6136 3332 6168
rect 3264 6100 3332 6136
rect 3264 6068 3282 6100
rect 3314 6068 3332 6100
rect 3264 6032 3332 6068
rect 3264 6000 3282 6032
rect 3314 6000 3332 6032
rect 3264 5964 3332 6000
rect 3264 5932 3282 5964
rect 3314 5932 3332 5964
rect 3264 5896 3332 5932
rect 3264 5864 3282 5896
rect 3314 5864 3332 5896
rect 3264 5828 3332 5864
rect 3264 5796 3282 5828
rect 3314 5796 3332 5828
rect 3264 5760 3332 5796
rect 3264 5728 3282 5760
rect 3314 5728 3332 5760
rect 3264 5692 3332 5728
rect 3264 5660 3282 5692
rect 3314 5660 3332 5692
rect 3264 5624 3332 5660
rect 3264 5592 3282 5624
rect 3314 5592 3332 5624
rect 3264 5556 3332 5592
rect 3264 5524 3282 5556
rect 3314 5524 3332 5556
rect 3264 5488 3332 5524
rect 3264 5456 3282 5488
rect 3314 5456 3332 5488
rect 3264 5420 3332 5456
rect 3264 5388 3282 5420
rect 3314 5388 3332 5420
rect 3264 5352 3332 5388
rect 3264 5320 3282 5352
rect 3314 5320 3332 5352
rect 3264 5284 3332 5320
rect 3264 5252 3282 5284
rect 3314 5252 3332 5284
rect 3264 5216 3332 5252
rect 3264 5184 3282 5216
rect 3314 5184 3332 5216
rect 3264 5148 3332 5184
rect 3264 5116 3282 5148
rect 3314 5116 3332 5148
rect 3264 5080 3332 5116
rect 3264 5048 3282 5080
rect 3314 5048 3332 5080
rect 3264 5012 3332 5048
rect 3264 4980 3282 5012
rect 3314 4980 3332 5012
rect 3264 4942 3332 4980
rect 3584 6644 3616 6660
rect 3584 6576 3616 6612
rect 3584 6508 3616 6544
rect 3584 6440 3616 6476
rect 3584 6372 3616 6408
rect 3584 6304 3616 6340
rect 3584 6236 3616 6272
rect 3584 6168 3616 6204
rect 3584 6100 3616 6136
rect 3584 6032 3616 6068
rect 3584 5964 3616 6000
rect 3584 5896 3616 5932
rect 3584 5828 3616 5864
rect 3584 5760 3616 5796
rect 3584 5692 3616 5728
rect 3584 5624 3616 5660
rect 3584 5556 3616 5592
rect 3584 5488 3616 5524
rect 3584 5420 3616 5456
rect 3584 5352 3616 5388
rect 3584 4942 3616 5320
rect 3755 6644 3797 6660
rect 3755 6617 3760 6644
rect 3792 6617 3797 6644
rect 3755 5347 3756 6617
rect 3796 5347 3797 6617
rect 3755 5320 3760 5347
rect 3792 5320 3797 5347
rect 3755 5304 3797 5320
rect 3936 6644 3968 6660
rect 3936 6576 3968 6612
rect 3936 6508 3968 6544
rect 3936 6440 3968 6476
rect 3936 6372 3968 6408
rect 3936 6304 3968 6340
rect 3936 6236 3968 6272
rect 3936 6168 3968 6204
rect 3936 6100 3968 6136
rect 3936 6032 3968 6068
rect 3936 5964 3968 6000
rect 3936 5896 3968 5932
rect 3936 5828 3968 5864
rect 3936 5760 3968 5796
rect 3936 5692 3968 5728
rect 3936 5624 3968 5660
rect 3936 5556 3968 5592
rect 3936 5488 3968 5524
rect 3936 5420 3968 5456
rect 3936 5352 3968 5388
rect 3936 4942 3968 5320
rect 4107 6644 4149 6660
rect 4107 6617 4112 6644
rect 4144 6617 4149 6644
rect 4107 5347 4108 6617
rect 4148 5347 4149 6617
rect 4107 5320 4112 5347
rect 4144 5320 4149 5347
rect 4107 5304 4149 5320
rect 4288 6644 4320 6660
rect 4288 6576 4320 6612
rect 4288 6508 4320 6544
rect 4288 6440 4320 6476
rect 4288 6372 4320 6408
rect 4288 6304 4320 6340
rect 4288 6236 4320 6272
rect 4288 6168 4320 6204
rect 4288 6100 4320 6136
rect 4288 6032 4320 6068
rect 4288 5964 4320 6000
rect 4288 5896 4320 5932
rect 4288 5828 4320 5864
rect 4288 5760 4320 5796
rect 4288 5692 4320 5728
rect 4288 5624 4320 5660
rect 4288 5556 4320 5592
rect 4288 5488 4320 5524
rect 4288 5420 4320 5456
rect 4288 5352 4320 5388
rect 4288 4942 4320 5320
rect 4459 6644 4501 6660
rect 4459 6617 4464 6644
rect 4496 6617 4501 6644
rect 4459 5347 4460 6617
rect 4500 5347 4501 6617
rect 4459 5320 4464 5347
rect 4496 5320 4501 5347
rect 4459 5304 4501 5320
rect 4640 6644 4672 6660
rect 4640 6576 4672 6612
rect 4640 6508 4672 6544
rect 4640 6440 4672 6476
rect 4640 6372 4672 6408
rect 4640 6304 4672 6340
rect 4640 6236 4672 6272
rect 4640 6168 4672 6204
rect 4640 6100 4672 6136
rect 4640 6032 4672 6068
rect 4640 5964 4672 6000
rect 4640 5896 4672 5932
rect 4640 5828 4672 5864
rect 4640 5760 4672 5796
rect 4640 5692 4672 5728
rect 4640 5624 4672 5660
rect 4640 5556 4672 5592
rect 4640 5488 4672 5524
rect 4640 5420 4672 5456
rect 4640 5352 4672 5388
rect 4640 4942 4672 5320
rect 4811 6644 4853 6660
rect 4811 6617 4816 6644
rect 4848 6617 4853 6644
rect 4811 5347 4812 6617
rect 4852 5347 4853 6617
rect 4811 5320 4816 5347
rect 4848 5320 4853 5347
rect 4811 5304 4853 5320
rect 4992 6644 5024 6660
rect 4992 6576 5024 6612
rect 4992 6508 5024 6544
rect 4992 6440 5024 6476
rect 4992 6372 5024 6408
rect 4992 6304 5024 6340
rect 4992 6236 5024 6272
rect 4992 6168 5024 6204
rect 4992 6100 5024 6136
rect 4992 6032 5024 6068
rect 4992 5964 5024 6000
rect 4992 5896 5024 5932
rect 4992 5828 5024 5864
rect 4992 5760 5024 5796
rect 4992 5692 5024 5728
rect 4992 5624 5024 5660
rect 4992 5556 5024 5592
rect 4992 5488 5024 5524
rect 4992 5420 5024 5456
rect 4992 5352 5024 5388
rect 4992 4942 5024 5320
rect 5163 6644 5205 6660
rect 5163 6617 5168 6644
rect 5200 6617 5205 6644
rect 5163 5347 5164 6617
rect 5204 5347 5205 6617
rect 5163 5320 5168 5347
rect 5200 5320 5205 5347
rect 5163 5304 5205 5320
rect 5344 6644 5376 6660
rect 5344 6576 5376 6612
rect 5344 6508 5376 6544
rect 5344 6440 5376 6476
rect 5344 6372 5376 6408
rect 5344 6304 5376 6340
rect 5344 6236 5376 6272
rect 5344 6168 5376 6204
rect 5344 6100 5376 6136
rect 5344 6032 5376 6068
rect 5344 5964 5376 6000
rect 5344 5896 5376 5932
rect 5344 5828 5376 5864
rect 5344 5760 5376 5796
rect 5344 5692 5376 5728
rect 5344 5624 5376 5660
rect 5344 5556 5376 5592
rect 5344 5488 5376 5524
rect 5344 5420 5376 5456
rect 5344 5352 5376 5388
rect 5344 4942 5376 5320
rect 5515 6644 5557 6660
rect 5515 6617 5520 6644
rect 5552 6617 5557 6644
rect 5515 5347 5516 6617
rect 5556 5347 5557 6617
rect 5515 5320 5520 5347
rect 5552 5320 5557 5347
rect 5515 5304 5557 5320
rect 5696 6644 5728 6660
rect 5696 6576 5728 6612
rect 5696 6508 5728 6544
rect 5696 6440 5728 6476
rect 5696 6372 5728 6408
rect 5696 6304 5728 6340
rect 5696 6236 5728 6272
rect 5696 6168 5728 6204
rect 5696 6100 5728 6136
rect 5696 6032 5728 6068
rect 5696 5964 5728 6000
rect 5696 5896 5728 5932
rect 5696 5828 5728 5864
rect 5696 5760 5728 5796
rect 5696 5692 5728 5728
rect 5696 5624 5728 5660
rect 5696 5556 5728 5592
rect 5696 5488 5728 5524
rect 5696 5420 5728 5456
rect 5696 5352 5728 5388
rect 5696 4942 5728 5320
rect 5867 6644 5909 6660
rect 5867 6617 5872 6644
rect 5904 6617 5909 6644
rect 5867 5347 5868 6617
rect 5908 5347 5909 6617
rect 5867 5320 5872 5347
rect 5904 5320 5909 5347
rect 5867 5304 5909 5320
rect 6048 6644 6080 6660
rect 6048 6576 6080 6612
rect 6048 6508 6080 6544
rect 6048 6440 6080 6476
rect 6048 6372 6080 6408
rect 6048 6304 6080 6340
rect 6048 6236 6080 6272
rect 6048 6168 6080 6204
rect 6048 6100 6080 6136
rect 6048 6032 6080 6068
rect 6048 5964 6080 6000
rect 6048 5896 6080 5932
rect 6048 5828 6080 5864
rect 6048 5760 6080 5796
rect 6048 5692 6080 5728
rect 6048 5624 6080 5660
rect 6048 5556 6080 5592
rect 6048 5488 6080 5524
rect 6048 5420 6080 5456
rect 6048 5352 6080 5388
rect 6048 4942 6080 5320
rect 6219 6644 6261 6660
rect 6219 6617 6224 6644
rect 6256 6617 6261 6644
rect 6219 5347 6220 6617
rect 6260 5347 6261 6617
rect 6219 5320 6224 5347
rect 6256 5320 6261 5347
rect 6219 5304 6261 5320
rect 6400 6644 6432 6660
rect 6400 6576 6432 6612
rect 6400 6508 6432 6544
rect 6400 6440 6432 6476
rect 6400 6372 6432 6408
rect 6400 6304 6432 6340
rect 6400 6236 6432 6272
rect 6400 6168 6432 6204
rect 6400 6100 6432 6136
rect 6400 6032 6432 6068
rect 6400 5964 6432 6000
rect 6400 5896 6432 5932
rect 6400 5828 6432 5864
rect 6400 5760 6432 5796
rect 6400 5692 6432 5728
rect 6400 5624 6432 5660
rect 6400 5556 6432 5592
rect 6400 5488 6432 5524
rect 6400 5420 6432 5456
rect 6400 5352 6432 5388
rect 6400 4942 6432 5320
rect 6571 6644 6613 6660
rect 6571 6617 6576 6644
rect 6608 6617 6613 6644
rect 6571 5347 6572 6617
rect 6612 5347 6613 6617
rect 6571 5320 6576 5347
rect 6608 5320 6613 5347
rect 6571 5304 6613 5320
rect 6752 6644 6784 6660
rect 6752 6576 6784 6612
rect 6752 6508 6784 6544
rect 6752 6440 6784 6476
rect 6752 6372 6784 6408
rect 6752 6304 6784 6340
rect 6752 6236 6784 6272
rect 6752 6168 6784 6204
rect 6752 6100 6784 6136
rect 6752 6032 6784 6068
rect 6752 5964 6784 6000
rect 6752 5896 6784 5932
rect 6752 5828 6784 5864
rect 6752 5760 6784 5796
rect 6752 5692 6784 5728
rect 6752 5624 6784 5660
rect 6752 5556 6784 5592
rect 6752 5488 6784 5524
rect 6752 5420 6784 5456
rect 6752 5352 6784 5388
rect 6752 4942 6784 5320
rect 6923 6644 6965 6660
rect 6923 6617 6928 6644
rect 6960 6617 6965 6644
rect 6923 5347 6924 6617
rect 6964 5347 6965 6617
rect 6923 5320 6928 5347
rect 6960 5320 6965 5347
rect 6923 5304 6965 5320
rect 7104 6644 7136 6660
rect 7104 6576 7136 6612
rect 7104 6508 7136 6544
rect 7104 6440 7136 6476
rect 7104 6372 7136 6408
rect 7104 6304 7136 6340
rect 7104 6236 7136 6272
rect 7104 6168 7136 6204
rect 7104 6100 7136 6136
rect 7104 6032 7136 6068
rect 7104 5964 7136 6000
rect 7104 5896 7136 5932
rect 7104 5828 7136 5864
rect 7104 5760 7136 5796
rect 7104 5692 7136 5728
rect 7104 5624 7136 5660
rect 7104 5556 7136 5592
rect 7104 5488 7136 5524
rect 7104 5420 7136 5456
rect 7104 5352 7136 5388
rect 7104 4942 7136 5320
rect 7275 6644 7317 6660
rect 7275 6617 7280 6644
rect 7312 6617 7317 6644
rect 7275 5347 7276 6617
rect 7316 5347 7317 6617
rect 7275 5320 7280 5347
rect 7312 5320 7317 5347
rect 7275 5304 7317 5320
rect 7456 6644 7488 6660
rect 7456 6576 7488 6612
rect 7456 6508 7488 6544
rect 7456 6440 7488 6476
rect 7456 6372 7488 6408
rect 7456 6304 7488 6340
rect 7456 6236 7488 6272
rect 7456 6168 7488 6204
rect 7456 6100 7488 6136
rect 7456 6032 7488 6068
rect 7456 5964 7488 6000
rect 7456 5896 7488 5932
rect 7456 5828 7488 5864
rect 7456 5760 7488 5796
rect 7456 5692 7488 5728
rect 7456 5624 7488 5660
rect 7456 5556 7488 5592
rect 7456 5488 7488 5524
rect 7456 5420 7488 5456
rect 7456 5352 7488 5388
rect 7456 4942 7488 5320
rect 7627 6644 7669 6660
rect 7627 6617 7632 6644
rect 7664 6617 7669 6644
rect 7627 5347 7628 6617
rect 7668 5347 7669 6617
rect 7627 5320 7632 5347
rect 7664 5320 7669 5347
rect 7627 5304 7669 5320
rect 7808 6644 7840 6660
rect 7808 6576 7840 6612
rect 7808 6508 7840 6544
rect 7808 6440 7840 6476
rect 7808 6372 7840 6408
rect 7808 6304 7840 6340
rect 7808 6236 7840 6272
rect 7808 6168 7840 6204
rect 7808 6100 7840 6136
rect 7808 6032 7840 6068
rect 7808 5964 7840 6000
rect 7808 5896 7840 5932
rect 7808 5828 7840 5864
rect 7808 5760 7840 5796
rect 7808 5692 7840 5728
rect 7808 5624 7840 5660
rect 7808 5556 7840 5592
rect 7808 5488 7840 5524
rect 7808 5420 7840 5456
rect 7808 5352 7840 5388
rect 7808 4942 7840 5320
rect 7979 6644 8021 6660
rect 7979 6617 7984 6644
rect 8016 6617 8021 6644
rect 7979 5347 7980 6617
rect 8020 5347 8021 6617
rect 7979 5320 7984 5347
rect 8016 5320 8021 5347
rect 7979 5304 8021 5320
rect 8160 6644 8192 6660
rect 8160 6576 8192 6612
rect 8160 6508 8192 6544
rect 8160 6440 8192 6476
rect 8160 6372 8192 6408
rect 8160 6304 8192 6340
rect 8160 6236 8192 6272
rect 8160 6168 8192 6204
rect 8160 6100 8192 6136
rect 8160 6032 8192 6068
rect 8160 5964 8192 6000
rect 8160 5896 8192 5932
rect 8160 5828 8192 5864
rect 8160 5760 8192 5796
rect 8160 5692 8192 5728
rect 8160 5624 8192 5660
rect 8160 5556 8192 5592
rect 8160 5488 8192 5524
rect 8160 5420 8192 5456
rect 8160 5352 8192 5388
rect 8160 4942 8192 5320
rect 8331 6644 8373 6660
rect 8331 6617 8336 6644
rect 8368 6617 8373 6644
rect 8331 5347 8332 6617
rect 8372 5347 8373 6617
rect 8331 5320 8336 5347
rect 8368 5320 8373 5347
rect 8331 5304 8373 5320
rect 8512 6644 8544 6660
rect 8512 6576 8544 6612
rect 8512 6508 8544 6544
rect 8512 6440 8544 6476
rect 8512 6372 8544 6408
rect 8512 6304 8544 6340
rect 8512 6236 8544 6272
rect 8512 6168 8544 6204
rect 8512 6100 8544 6136
rect 8512 6032 8544 6068
rect 8512 5964 8544 6000
rect 8512 5896 8544 5932
rect 8512 5828 8544 5864
rect 8512 5760 8544 5796
rect 8512 5692 8544 5728
rect 8512 5624 8544 5660
rect 8512 5556 8544 5592
rect 8512 5488 8544 5524
rect 8512 5420 8544 5456
rect 8512 5352 8544 5388
rect 8512 4942 8544 5320
rect 8683 6644 8725 6660
rect 8683 6617 8688 6644
rect 8720 6617 8725 6644
rect 8683 5347 8684 6617
rect 8724 5347 8725 6617
rect 8683 5320 8688 5347
rect 8720 5320 8725 5347
rect 8683 5304 8725 5320
rect 8864 6644 8896 6660
rect 8864 6576 8896 6612
rect 8864 6508 8896 6544
rect 8864 6440 8896 6476
rect 8864 6372 8896 6408
rect 8864 6304 8896 6340
rect 8864 6236 8896 6272
rect 8864 6168 8896 6204
rect 8864 6100 8896 6136
rect 8864 6032 8896 6068
rect 8864 5964 8896 6000
rect 8864 5896 8896 5932
rect 8864 5828 8896 5864
rect 8864 5760 8896 5796
rect 8864 5692 8896 5728
rect 8864 5624 8896 5660
rect 8864 5556 8896 5592
rect 8864 5488 8896 5524
rect 8864 5420 8896 5456
rect 8864 5352 8896 5388
rect 8864 4942 8896 5320
rect 9035 6644 9077 6660
rect 9035 6617 9040 6644
rect 9072 6617 9077 6644
rect 9035 5347 9036 6617
rect 9076 5347 9077 6617
rect 9035 5320 9040 5347
rect 9072 5320 9077 5347
rect 9035 5304 9077 5320
rect 9216 6644 9248 6660
rect 9216 6576 9248 6612
rect 9216 6508 9248 6544
rect 9216 6440 9248 6476
rect 9216 6372 9248 6408
rect 9216 6304 9248 6340
rect 9216 6236 9248 6272
rect 9216 6168 9248 6204
rect 9216 6100 9248 6136
rect 9216 6032 9248 6068
rect 9216 5964 9248 6000
rect 9216 5896 9248 5932
rect 9216 5828 9248 5864
rect 9216 5760 9248 5796
rect 9216 5692 9248 5728
rect 9216 5624 9248 5660
rect 9216 5556 9248 5592
rect 9216 5488 9248 5524
rect 9216 5420 9248 5456
rect 9216 5352 9248 5388
rect 9216 4942 9248 5320
rect 9387 6644 9429 6660
rect 9387 6617 9392 6644
rect 9424 6617 9429 6644
rect 9387 5347 9388 6617
rect 9428 5347 9429 6617
rect 9387 5320 9392 5347
rect 9424 5320 9429 5347
rect 9387 5304 9429 5320
rect 9568 6644 9600 6660
rect 9568 6576 9600 6612
rect 9568 6508 9600 6544
rect 9568 6440 9600 6476
rect 9568 6372 9600 6408
rect 9568 6304 9600 6340
rect 9568 6236 9600 6272
rect 9568 6168 9600 6204
rect 9568 6100 9600 6136
rect 9568 6032 9600 6068
rect 9568 5964 9600 6000
rect 9568 5896 9600 5932
rect 9568 5828 9600 5864
rect 9568 5760 9600 5796
rect 9568 5692 9600 5728
rect 9568 5624 9600 5660
rect 9568 5556 9600 5592
rect 9568 5488 9600 5524
rect 9568 5420 9600 5456
rect 9568 5352 9600 5388
rect 9568 4942 9600 5320
rect 9739 6644 9781 6660
rect 9739 6617 9744 6644
rect 9776 6617 9781 6644
rect 9739 5347 9740 6617
rect 9780 5347 9781 6617
rect 9739 5320 9744 5347
rect 9776 5320 9781 5347
rect 9739 5304 9781 5320
rect 9920 6644 9952 6660
rect 9920 6576 9952 6612
rect 9920 6508 9952 6544
rect 9920 6440 9952 6476
rect 9920 6372 9952 6408
rect 9920 6304 9952 6340
rect 9920 6236 9952 6272
rect 9920 6168 9952 6204
rect 9920 6100 9952 6136
rect 9920 6032 9952 6068
rect 9920 5964 9952 6000
rect 9920 5896 9952 5932
rect 9920 5828 9952 5864
rect 9920 5760 9952 5796
rect 9920 5692 9952 5728
rect 9920 5624 9952 5660
rect 9920 5556 9952 5592
rect 9920 5488 9952 5524
rect 9920 5420 9952 5456
rect 9920 5352 9952 5388
rect 9920 4942 9952 5320
rect 10091 6644 10133 6660
rect 10091 6617 10096 6644
rect 10128 6617 10133 6644
rect 10091 5347 10092 6617
rect 10132 5347 10133 6617
rect 10091 5320 10096 5347
rect 10128 5320 10133 5347
rect 10091 5304 10133 5320
rect 10272 6644 10304 6660
rect 10272 6576 10304 6612
rect 10272 6508 10304 6544
rect 10272 6440 10304 6476
rect 10272 6372 10304 6408
rect 10272 6304 10304 6340
rect 10272 6236 10304 6272
rect 10272 6168 10304 6204
rect 10272 6100 10304 6136
rect 10272 6032 10304 6068
rect 10272 5964 10304 6000
rect 10272 5896 10304 5932
rect 10272 5828 10304 5864
rect 10272 5760 10304 5796
rect 10272 5692 10304 5728
rect 10272 5624 10304 5660
rect 10272 5556 10304 5592
rect 10272 5488 10304 5524
rect 10272 5420 10304 5456
rect 10272 5352 10304 5388
rect 10272 4942 10304 5320
rect 10443 6644 10485 6660
rect 10443 6617 10448 6644
rect 10480 6617 10485 6644
rect 10443 5347 10444 6617
rect 10484 5347 10485 6617
rect 10443 5320 10448 5347
rect 10480 5320 10485 5347
rect 10443 5304 10485 5320
rect 10624 6644 10656 6660
rect 10624 6576 10656 6612
rect 10624 6508 10656 6544
rect 10624 6440 10656 6476
rect 10624 6372 10656 6408
rect 10624 6304 10656 6340
rect 10624 6236 10656 6272
rect 10624 6168 10656 6204
rect 10624 6100 10656 6136
rect 10624 6032 10656 6068
rect 10624 5964 10656 6000
rect 10624 5896 10656 5932
rect 10624 5828 10656 5864
rect 10624 5760 10656 5796
rect 10624 5692 10656 5728
rect 10624 5624 10656 5660
rect 10624 5556 10656 5592
rect 10624 5488 10656 5524
rect 10624 5420 10656 5456
rect 10624 5352 10656 5388
rect 10624 4942 10656 5320
rect 10795 6644 10837 6660
rect 10795 6617 10800 6644
rect 10832 6617 10837 6644
rect 10795 5347 10796 6617
rect 10836 5347 10837 6617
rect 10795 5320 10800 5347
rect 10832 5320 10837 5347
rect 10795 5304 10837 5320
rect 10976 6644 11008 6660
rect 10976 6576 11008 6612
rect 10976 6508 11008 6544
rect 10976 6440 11008 6476
rect 10976 6372 11008 6408
rect 10976 6304 11008 6340
rect 10976 6236 11008 6272
rect 10976 6168 11008 6204
rect 10976 6100 11008 6136
rect 10976 6032 11008 6068
rect 10976 5964 11008 6000
rect 10976 5896 11008 5932
rect 10976 5828 11008 5864
rect 10976 5760 11008 5796
rect 10976 5692 11008 5728
rect 10976 5624 11008 5660
rect 10976 5556 11008 5592
rect 10976 5488 11008 5524
rect 10976 5420 11008 5456
rect 10976 5352 11008 5388
rect 10976 4942 11008 5320
rect 11147 6644 11189 6660
rect 11147 6617 11152 6644
rect 11184 6617 11189 6644
rect 11147 5347 11148 6617
rect 11188 5347 11189 6617
rect 11147 5320 11152 5347
rect 11184 5320 11189 5347
rect 11147 5304 11189 5320
rect 11328 6644 11360 6660
rect 11328 6576 11360 6612
rect 11328 6508 11360 6544
rect 11328 6440 11360 6476
rect 11328 6372 11360 6408
rect 11328 6304 11360 6340
rect 11328 6236 11360 6272
rect 11328 6168 11360 6204
rect 11328 6100 11360 6136
rect 11328 6032 11360 6068
rect 11328 5964 11360 6000
rect 11328 5896 11360 5932
rect 11328 5828 11360 5864
rect 11328 5760 11360 5796
rect 11328 5692 11360 5728
rect 11328 5624 11360 5660
rect 11328 5556 11360 5592
rect 11328 5488 11360 5524
rect 11328 5420 11360 5456
rect 11328 5352 11360 5388
rect 11328 4942 11360 5320
rect 11499 6644 11541 6660
rect 11499 6617 11504 6644
rect 11536 6617 11541 6644
rect 11499 5347 11500 6617
rect 11540 5347 11541 6617
rect 11499 5320 11504 5347
rect 11536 5320 11541 5347
rect 11499 5304 11541 5320
rect 11680 6644 11712 6660
rect 11680 6576 11712 6612
rect 11680 6508 11712 6544
rect 11680 6440 11712 6476
rect 11680 6372 11712 6408
rect 11680 6304 11712 6340
rect 11680 6236 11712 6272
rect 11680 6168 11712 6204
rect 11680 6100 11712 6136
rect 11680 6032 11712 6068
rect 11680 5964 11712 6000
rect 11680 5896 11712 5932
rect 11680 5828 11712 5864
rect 11680 5760 11712 5796
rect 11680 5692 11712 5728
rect 11680 5624 11712 5660
rect 11680 5556 11712 5592
rect 11680 5488 11712 5524
rect 11680 5420 11712 5456
rect 11680 5352 11712 5388
rect 11680 4942 11712 5320
rect 11851 6644 11893 6660
rect 11851 6617 11856 6644
rect 11888 6617 11893 6644
rect 11851 5347 11852 6617
rect 11892 5347 11893 6617
rect 11851 5320 11856 5347
rect 11888 5320 11893 5347
rect 11851 5304 11893 5320
rect 12032 6644 12064 6660
rect 12032 6576 12064 6612
rect 12032 6508 12064 6544
rect 12032 6440 12064 6476
rect 12032 6372 12064 6408
rect 12032 6304 12064 6340
rect 12032 6236 12064 6272
rect 12032 6168 12064 6204
rect 12032 6100 12064 6136
rect 12032 6032 12064 6068
rect 12032 5964 12064 6000
rect 12032 5896 12064 5932
rect 12032 5828 12064 5864
rect 12032 5760 12064 5796
rect 12032 5692 12064 5728
rect 12032 5624 12064 5660
rect 12032 5556 12064 5592
rect 12032 5488 12064 5524
rect 12032 5420 12064 5456
rect 12032 5352 12064 5388
rect 12032 4942 12064 5320
rect 12203 6644 12245 6660
rect 12203 6617 12208 6644
rect 12240 6617 12245 6644
rect 12203 5347 12204 6617
rect 12244 5347 12245 6617
rect 12203 5320 12208 5347
rect 12240 5320 12245 5347
rect 12203 5304 12245 5320
rect 12384 6644 12416 6660
rect 12384 6576 12416 6612
rect 12384 6508 12416 6544
rect 12384 6440 12416 6476
rect 12384 6372 12416 6408
rect 12384 6304 12416 6340
rect 12384 6236 12416 6272
rect 12384 6168 12416 6204
rect 12384 6100 12416 6136
rect 12384 6032 12416 6068
rect 12384 5964 12416 6000
rect 12384 5896 12416 5932
rect 12384 5828 12416 5864
rect 12384 5760 12416 5796
rect 12384 5692 12416 5728
rect 12384 5624 12416 5660
rect 12384 5556 12416 5592
rect 12384 5488 12416 5524
rect 12384 5420 12416 5456
rect 12384 5352 12416 5388
rect 12384 4942 12416 5320
rect 12668 6644 12736 6680
rect 12668 6612 12686 6644
rect 12718 6612 12736 6644
rect 12668 6576 12736 6612
rect 12668 6544 12686 6576
rect 12718 6544 12736 6576
rect 12668 6508 12736 6544
rect 12668 6476 12686 6508
rect 12718 6476 12736 6508
rect 12668 6440 12736 6476
rect 12668 6408 12686 6440
rect 12718 6408 12736 6440
rect 12668 6372 12736 6408
rect 12668 6340 12686 6372
rect 12718 6340 12736 6372
rect 12668 6304 12736 6340
rect 12668 6272 12686 6304
rect 12718 6272 12736 6304
rect 12668 6236 12736 6272
rect 12668 6204 12686 6236
rect 12718 6204 12736 6236
rect 12668 6168 12736 6204
rect 12668 6136 12686 6168
rect 12718 6136 12736 6168
rect 12668 6100 12736 6136
rect 12668 6068 12686 6100
rect 12718 6068 12736 6100
rect 12668 6032 12736 6068
rect 12668 6000 12686 6032
rect 12718 6000 12736 6032
rect 12668 5964 12736 6000
rect 12668 5932 12686 5964
rect 12718 5932 12736 5964
rect 12668 5896 12736 5932
rect 12668 5864 12686 5896
rect 12718 5864 12736 5896
rect 12668 5828 12736 5864
rect 12668 5796 12686 5828
rect 12718 5796 12736 5828
rect 12668 5760 12736 5796
rect 12668 5728 12686 5760
rect 12718 5728 12736 5760
rect 12668 5692 12736 5728
rect 12668 5660 12686 5692
rect 12718 5660 12736 5692
rect 12668 5624 12736 5660
rect 12668 5592 12686 5624
rect 12718 5592 12736 5624
rect 12668 5556 12736 5592
rect 12668 5524 12686 5556
rect 12718 5524 12736 5556
rect 12668 5488 12736 5524
rect 12668 5456 12686 5488
rect 12718 5456 12736 5488
rect 12668 5420 12736 5456
rect 12668 5388 12686 5420
rect 12718 5388 12736 5420
rect 12668 5352 12736 5388
rect 12668 5320 12686 5352
rect 12718 5320 12736 5352
rect 12668 5284 12736 5320
rect 12668 5252 12686 5284
rect 12718 5252 12736 5284
rect 12668 5216 12736 5252
rect 12668 5184 12686 5216
rect 12718 5184 12736 5216
rect 12668 5148 12736 5184
rect 12668 5116 12686 5148
rect 12718 5116 12736 5148
rect 12668 5080 12736 5116
rect 12668 5048 12686 5080
rect 12718 5048 12736 5080
rect 12668 5012 12736 5048
rect 12668 4980 12686 5012
rect 12718 4980 12736 5012
rect 12668 4942 12736 4980
rect 3264 4924 12736 4942
rect 3264 4892 3292 4924
rect 3324 4892 3360 4924
rect 3392 4892 3428 4924
rect 3460 4892 3496 4924
rect 3528 4892 3564 4924
rect 3596 4892 3632 4924
rect 3664 4892 3700 4924
rect 3732 4892 3768 4924
rect 3800 4892 3836 4924
rect 3868 4892 3904 4924
rect 3936 4892 3972 4924
rect 4004 4892 4040 4924
rect 4072 4892 4108 4924
rect 4140 4892 4176 4924
rect 4208 4892 4244 4924
rect 4276 4892 4312 4924
rect 4344 4892 4380 4924
rect 4412 4892 4448 4924
rect 4480 4892 4516 4924
rect 4548 4892 4584 4924
rect 4616 4892 4652 4924
rect 4684 4892 4720 4924
rect 4752 4892 4788 4924
rect 4820 4892 4856 4924
rect 4888 4892 4924 4924
rect 4956 4892 4992 4924
rect 5024 4892 5060 4924
rect 5092 4892 5128 4924
rect 5160 4892 5196 4924
rect 5228 4892 5264 4924
rect 5296 4892 5332 4924
rect 5364 4892 5400 4924
rect 5432 4892 5468 4924
rect 5500 4892 5536 4924
rect 5568 4892 5604 4924
rect 5636 4892 5672 4924
rect 5704 4892 5740 4924
rect 5772 4892 5808 4924
rect 5840 4892 5876 4924
rect 5908 4892 5944 4924
rect 5976 4892 6012 4924
rect 6044 4892 6080 4924
rect 6112 4892 6148 4924
rect 6180 4892 6216 4924
rect 6248 4892 6284 4924
rect 6316 4892 6352 4924
rect 6384 4892 6420 4924
rect 6452 4892 6488 4924
rect 6520 4892 6556 4924
rect 6588 4892 6624 4924
rect 6656 4892 6692 4924
rect 6724 4892 6760 4924
rect 6792 4892 6828 4924
rect 6860 4892 6896 4924
rect 6928 4892 6964 4924
rect 6996 4892 7032 4924
rect 7064 4892 7100 4924
rect 7132 4892 7168 4924
rect 7200 4892 7236 4924
rect 7268 4892 7304 4924
rect 7336 4892 7372 4924
rect 7404 4892 7440 4924
rect 7472 4892 7508 4924
rect 7540 4892 7576 4924
rect 7608 4892 7644 4924
rect 7676 4892 7712 4924
rect 7744 4892 7780 4924
rect 7812 4892 7848 4924
rect 7880 4892 7916 4924
rect 7948 4892 7984 4924
rect 8016 4892 8052 4924
rect 8084 4892 8120 4924
rect 8152 4892 8188 4924
rect 8220 4892 8256 4924
rect 8288 4892 8324 4924
rect 8356 4892 8392 4924
rect 8424 4892 8460 4924
rect 8492 4892 8528 4924
rect 8560 4892 8596 4924
rect 8628 4892 8664 4924
rect 8696 4892 8732 4924
rect 8764 4892 8800 4924
rect 8832 4892 8868 4924
rect 8900 4892 8936 4924
rect 8968 4892 9004 4924
rect 9036 4892 9072 4924
rect 9104 4892 9140 4924
rect 9172 4892 9208 4924
rect 9240 4892 9276 4924
rect 9308 4892 9344 4924
rect 9376 4892 9412 4924
rect 9444 4892 9480 4924
rect 9512 4892 9548 4924
rect 9580 4892 9616 4924
rect 9648 4892 9684 4924
rect 9716 4892 9752 4924
rect 9784 4892 9820 4924
rect 9852 4892 9888 4924
rect 9920 4892 9956 4924
rect 9988 4892 10024 4924
rect 10056 4892 10092 4924
rect 10124 4892 10160 4924
rect 10192 4892 10228 4924
rect 10260 4892 10296 4924
rect 10328 4892 10364 4924
rect 10396 4892 10432 4924
rect 10464 4892 10500 4924
rect 10532 4892 10568 4924
rect 10600 4892 10636 4924
rect 10668 4892 10704 4924
rect 10736 4892 10772 4924
rect 10804 4892 10840 4924
rect 10872 4892 10908 4924
rect 10940 4892 10976 4924
rect 11008 4892 11044 4924
rect 11076 4892 11112 4924
rect 11144 4892 11180 4924
rect 11212 4892 11248 4924
rect 11280 4892 11316 4924
rect 11348 4892 11384 4924
rect 11416 4892 11452 4924
rect 11484 4892 11520 4924
rect 11552 4892 11588 4924
rect 11620 4892 11656 4924
rect 11688 4892 11724 4924
rect 11756 4892 11792 4924
rect 11824 4892 11860 4924
rect 11892 4892 11928 4924
rect 11960 4892 11996 4924
rect 12028 4892 12064 4924
rect 12096 4892 12132 4924
rect 12164 4892 12200 4924
rect 12232 4892 12268 4924
rect 12300 4892 12336 4924
rect 12368 4892 12404 4924
rect 12436 4892 12472 4924
rect 12504 4892 12540 4924
rect 12572 4892 12608 4924
rect 12640 4892 12676 4924
rect 12708 4892 12736 4924
rect 3264 4874 12736 4892
rect 0 4448 16000 4466
rect 0 4416 28 4448
rect 60 4416 96 4448
rect 128 4416 164 4448
rect 196 4416 232 4448
rect 264 4416 300 4448
rect 332 4416 368 4448
rect 400 4416 436 4448
rect 468 4416 504 4448
rect 536 4416 572 4448
rect 604 4416 640 4448
rect 672 4416 708 4448
rect 740 4416 776 4448
rect 808 4416 844 4448
rect 876 4416 912 4448
rect 944 4416 980 4448
rect 1012 4416 1048 4448
rect 1080 4416 1116 4448
rect 1148 4416 1184 4448
rect 1216 4416 1252 4448
rect 1284 4416 1320 4448
rect 1352 4416 1388 4448
rect 1420 4416 1456 4448
rect 1488 4416 1524 4448
rect 1556 4416 1592 4448
rect 1624 4416 1660 4448
rect 1692 4416 1728 4448
rect 1760 4416 1796 4448
rect 1828 4416 1864 4448
rect 1896 4416 1932 4448
rect 1964 4416 2000 4448
rect 2032 4416 2068 4448
rect 2100 4416 2136 4448
rect 2168 4416 2204 4448
rect 2236 4416 2272 4448
rect 2304 4416 2340 4448
rect 2372 4416 2408 4448
rect 2440 4416 2476 4448
rect 2508 4416 2544 4448
rect 2576 4416 2612 4448
rect 2644 4416 2680 4448
rect 2712 4416 2748 4448
rect 2780 4416 2816 4448
rect 2848 4416 2884 4448
rect 2916 4416 2952 4448
rect 2984 4416 3020 4448
rect 3052 4416 3088 4448
rect 3120 4416 3156 4448
rect 3188 4416 3224 4448
rect 3256 4416 3292 4448
rect 3324 4416 3360 4448
rect 3392 4416 3428 4448
rect 3460 4416 3496 4448
rect 3528 4416 3564 4448
rect 3596 4416 3632 4448
rect 3664 4416 3700 4448
rect 3732 4416 3768 4448
rect 3800 4416 3836 4448
rect 3868 4416 3904 4448
rect 3936 4416 3972 4448
rect 4004 4416 4040 4448
rect 4072 4416 4108 4448
rect 4140 4416 4176 4448
rect 4208 4416 4244 4448
rect 4276 4416 4312 4448
rect 4344 4416 4380 4448
rect 4412 4416 4448 4448
rect 4480 4416 4516 4448
rect 4548 4416 4584 4448
rect 4616 4416 4652 4448
rect 4684 4416 4720 4448
rect 4752 4416 4788 4448
rect 4820 4416 4856 4448
rect 4888 4416 4924 4448
rect 4956 4416 4992 4448
rect 5024 4416 5060 4448
rect 5092 4416 5128 4448
rect 5160 4416 5196 4448
rect 5228 4416 5264 4448
rect 5296 4416 5332 4448
rect 5364 4416 5400 4448
rect 5432 4416 5468 4448
rect 5500 4416 5536 4448
rect 5568 4416 5604 4448
rect 5636 4416 5672 4448
rect 5704 4416 5740 4448
rect 5772 4416 5808 4448
rect 5840 4416 5876 4448
rect 5908 4416 5944 4448
rect 5976 4416 6012 4448
rect 6044 4416 6080 4448
rect 6112 4416 6148 4448
rect 6180 4416 6216 4448
rect 6248 4416 6284 4448
rect 6316 4416 6352 4448
rect 6384 4416 6420 4448
rect 6452 4416 6488 4448
rect 6520 4416 6556 4448
rect 6588 4416 6624 4448
rect 6656 4416 6692 4448
rect 6724 4416 6760 4448
rect 6792 4416 6828 4448
rect 6860 4416 6896 4448
rect 6928 4416 6964 4448
rect 6996 4416 7032 4448
rect 7064 4416 7100 4448
rect 7132 4416 7168 4448
rect 7200 4416 7236 4448
rect 7268 4416 7304 4448
rect 7336 4416 7372 4448
rect 7404 4416 7440 4448
rect 7472 4416 7508 4448
rect 7540 4416 7576 4448
rect 7608 4416 7644 4448
rect 7676 4416 7712 4448
rect 7744 4416 7780 4448
rect 7812 4416 7848 4448
rect 7880 4416 7916 4448
rect 7948 4416 7984 4448
rect 8016 4416 8052 4448
rect 8084 4416 8120 4448
rect 8152 4416 8188 4448
rect 8220 4416 8256 4448
rect 8288 4416 8324 4448
rect 8356 4416 8392 4448
rect 8424 4416 8460 4448
rect 8492 4416 8528 4448
rect 8560 4416 8596 4448
rect 8628 4416 8664 4448
rect 8696 4416 8732 4448
rect 8764 4416 8800 4448
rect 8832 4416 8868 4448
rect 8900 4416 8936 4448
rect 8968 4416 9004 4448
rect 9036 4416 9072 4448
rect 9104 4416 9140 4448
rect 9172 4416 9208 4448
rect 9240 4416 9276 4448
rect 9308 4416 9344 4448
rect 9376 4416 9412 4448
rect 9444 4416 9480 4448
rect 9512 4416 9548 4448
rect 9580 4416 9616 4448
rect 9648 4416 9684 4448
rect 9716 4416 9752 4448
rect 9784 4416 9820 4448
rect 9852 4416 9888 4448
rect 9920 4416 9956 4448
rect 9988 4416 10024 4448
rect 10056 4416 10092 4448
rect 10124 4416 10160 4448
rect 10192 4416 10228 4448
rect 10260 4416 10296 4448
rect 10328 4416 10364 4448
rect 10396 4416 10432 4448
rect 10464 4416 10500 4448
rect 10532 4416 10568 4448
rect 10600 4416 10636 4448
rect 10668 4416 10704 4448
rect 10736 4416 10772 4448
rect 10804 4416 10840 4448
rect 10872 4416 10908 4448
rect 10940 4416 10976 4448
rect 11008 4416 11044 4448
rect 11076 4416 11112 4448
rect 11144 4416 11180 4448
rect 11212 4416 11248 4448
rect 11280 4416 11316 4448
rect 11348 4416 11384 4448
rect 11416 4416 11452 4448
rect 11484 4416 11520 4448
rect 11552 4416 11588 4448
rect 11620 4416 11656 4448
rect 11688 4416 11724 4448
rect 11756 4416 11792 4448
rect 11824 4416 11860 4448
rect 11892 4416 11928 4448
rect 11960 4416 11996 4448
rect 12028 4416 12064 4448
rect 12096 4416 12132 4448
rect 12164 4416 12200 4448
rect 12232 4416 12268 4448
rect 12300 4416 12336 4448
rect 12368 4416 12404 4448
rect 12436 4416 12472 4448
rect 12504 4416 12540 4448
rect 12572 4416 12608 4448
rect 12640 4416 12676 4448
rect 12708 4416 12744 4448
rect 12776 4416 12812 4448
rect 12844 4416 12880 4448
rect 12912 4416 12948 4448
rect 12980 4416 13016 4448
rect 13048 4416 13084 4448
rect 13116 4416 13152 4448
rect 13184 4416 13220 4448
rect 13252 4416 13288 4448
rect 13320 4416 13356 4448
rect 13388 4416 13424 4448
rect 13456 4416 13492 4448
rect 13524 4416 13560 4448
rect 13592 4416 13628 4448
rect 13660 4416 13696 4448
rect 13728 4416 13764 4448
rect 13796 4416 13832 4448
rect 13864 4416 13900 4448
rect 13932 4416 13968 4448
rect 14000 4416 14036 4448
rect 14068 4416 14104 4448
rect 14136 4416 14172 4448
rect 14204 4416 14240 4448
rect 14272 4416 14308 4448
rect 14340 4416 14376 4448
rect 14408 4416 14444 4448
rect 14476 4416 14512 4448
rect 14544 4416 14580 4448
rect 14612 4416 14648 4448
rect 14680 4416 14716 4448
rect 14748 4416 14784 4448
rect 14816 4416 14852 4448
rect 14884 4416 14920 4448
rect 14952 4416 14988 4448
rect 15020 4416 15056 4448
rect 15088 4416 15124 4448
rect 15156 4416 15192 4448
rect 15224 4416 15260 4448
rect 15292 4416 15328 4448
rect 15360 4416 15396 4448
rect 15428 4416 15464 4448
rect 15496 4416 15532 4448
rect 15564 4416 15600 4448
rect 15632 4416 15668 4448
rect 15700 4416 15736 4448
rect 15768 4416 15804 4448
rect 15836 4416 15872 4448
rect 15904 4416 15940 4448
rect 15972 4416 16000 4448
rect 0 4398 16000 4416
rect 0 4357 68 4398
rect 0 4325 18 4357
rect 50 4325 68 4357
rect 0 4289 68 4325
rect 0 4257 18 4289
rect 50 4257 68 4289
rect 0 4221 68 4257
rect 0 4189 18 4221
rect 50 4189 68 4221
rect 0 4153 68 4189
rect 0 4121 18 4153
rect 50 4121 68 4153
rect 0 4085 68 4121
rect 0 4053 18 4085
rect 50 4053 68 4085
rect 0 4017 68 4053
rect 0 3985 18 4017
rect 50 3985 68 4017
rect 0 3949 68 3985
rect 0 3917 18 3949
rect 50 3917 68 3949
rect 0 3881 68 3917
rect 0 3849 18 3881
rect 50 3849 68 3881
rect 0 3813 68 3849
rect 0 3781 18 3813
rect 50 3781 68 3813
rect 0 3745 68 3781
rect 0 3713 18 3745
rect 50 3713 68 3745
rect 0 3677 68 3713
rect 0 3645 18 3677
rect 50 3645 68 3677
rect 0 3609 68 3645
rect 0 3577 18 3609
rect 50 3577 68 3609
rect 0 3541 68 3577
rect 0 3509 18 3541
rect 50 3509 68 3541
rect 0 3473 68 3509
rect 0 3441 18 3473
rect 50 3441 68 3473
rect 0 3405 68 3441
rect 0 3373 18 3405
rect 50 3373 68 3405
rect 0 3337 68 3373
rect 0 3305 18 3337
rect 50 3305 68 3337
rect 0 3269 68 3305
rect 0 3237 18 3269
rect 50 3237 68 3269
rect 0 3201 68 3237
rect 0 3169 18 3201
rect 50 3169 68 3201
rect 0 3133 68 3169
rect 0 3101 18 3133
rect 50 3101 68 3133
rect 0 3065 68 3101
rect 0 3033 18 3065
rect 50 3033 68 3065
rect 0 2997 68 3033
rect 0 2965 18 2997
rect 50 2965 68 2997
rect 0 2929 68 2965
rect 0 2897 18 2929
rect 50 2897 68 2929
rect 0 2861 68 2897
rect 0 2829 18 2861
rect 50 2829 68 2861
rect 0 2793 68 2829
rect 0 2761 18 2793
rect 50 2761 68 2793
rect 0 2725 68 2761
rect 0 2693 18 2725
rect 50 2693 68 2725
rect 0 2657 68 2693
rect 0 2625 18 2657
rect 50 2625 68 2657
rect 0 2589 68 2625
rect 0 2557 18 2589
rect 50 2557 68 2589
rect 0 2521 68 2557
rect 0 2489 18 2521
rect 50 2489 68 2521
rect 0 2453 68 2489
rect 0 2421 18 2453
rect 50 2421 68 2453
rect 0 2385 68 2421
rect 0 2353 18 2385
rect 50 2353 68 2385
rect 0 2317 68 2353
rect 0 2285 18 2317
rect 50 2285 68 2317
rect 0 2249 68 2285
rect 0 2217 18 2249
rect 50 2217 68 2249
rect 0 2181 68 2217
rect 0 2149 18 2181
rect 50 2149 68 2181
rect 0 2113 68 2149
rect 0 2081 18 2113
rect 50 2081 68 2113
rect 0 2045 68 2081
rect 0 2013 18 2045
rect 50 2013 68 2045
rect 0 1977 68 2013
rect 0 1945 18 1977
rect 50 1945 68 1977
rect 0 1909 68 1945
rect 0 1877 18 1909
rect 50 1877 68 1909
rect 0 1841 68 1877
rect 0 1809 18 1841
rect 50 1809 68 1841
rect 0 1773 68 1809
rect 0 1741 18 1773
rect 50 1741 68 1773
rect 0 1705 68 1741
rect 0 1673 18 1705
rect 50 1673 68 1705
rect 0 1637 68 1673
rect 0 1605 18 1637
rect 50 1605 68 1637
rect 0 1569 68 1605
rect 0 1537 18 1569
rect 50 1537 68 1569
rect 0 1501 68 1537
rect 0 1469 18 1501
rect 50 1469 68 1501
rect 0 1433 68 1469
rect 0 1401 18 1433
rect 50 1401 68 1433
rect 0 1365 68 1401
rect 0 1333 18 1365
rect 50 1333 68 1365
rect 0 1297 68 1333
rect 0 1265 18 1297
rect 50 1265 68 1297
rect 0 1229 68 1265
rect 0 1197 18 1229
rect 50 1197 68 1229
rect 0 1161 68 1197
rect 0 1129 18 1161
rect 50 1129 68 1161
rect 0 1093 68 1129
rect 0 1061 18 1093
rect 50 1061 68 1093
rect 0 1025 68 1061
rect 0 993 18 1025
rect 50 993 68 1025
rect 0 957 68 993
rect 0 925 18 957
rect 50 925 68 957
rect 0 889 68 925
rect 0 857 18 889
rect 50 857 68 889
rect 0 821 68 857
rect 0 789 18 821
rect 50 789 68 821
rect 0 753 68 789
rect 0 721 18 753
rect 50 721 68 753
rect 0 685 68 721
rect 0 653 18 685
rect 50 653 68 685
rect 0 617 68 653
rect 0 585 18 617
rect 50 585 68 617
rect 0 549 68 585
rect 0 517 18 549
rect 50 517 68 549
rect 0 481 68 517
rect 0 449 18 481
rect 50 449 68 481
rect 0 413 68 449
rect 540 4024 572 4398
rect 540 3956 572 3992
rect 540 3888 572 3924
rect 540 3820 572 3856
rect 540 3752 572 3788
rect 540 3684 572 3720
rect 540 3616 572 3652
rect 540 3548 572 3584
rect 540 3480 572 3516
rect 540 3412 572 3448
rect 540 3344 572 3380
rect 540 3276 572 3312
rect 540 3208 572 3244
rect 540 3140 572 3176
rect 540 3072 572 3108
rect 540 3004 572 3040
rect 540 2936 572 2972
rect 540 2868 572 2904
rect 540 2800 572 2836
rect 540 2732 572 2768
rect 540 2664 572 2700
rect 540 2596 572 2632
rect 540 2528 572 2564
rect 540 2460 572 2496
rect 540 2392 572 2428
rect 540 2324 572 2360
rect 540 2174 572 2292
rect 540 2106 572 2142
rect 540 2038 572 2074
rect 540 1970 572 2006
rect 540 1902 572 1938
rect 540 1834 572 1870
rect 540 1766 572 1802
rect 540 1698 572 1734
rect 540 1630 572 1666
rect 540 1562 572 1598
rect 540 1494 572 1530
rect 540 1426 572 1462
rect 540 1358 572 1394
rect 540 1290 572 1326
rect 540 1222 572 1258
rect 540 1154 572 1190
rect 540 1086 572 1122
rect 540 1018 572 1054
rect 540 950 572 986
rect 540 882 572 918
rect 540 814 572 850
rect 540 746 572 782
rect 540 678 572 714
rect 540 610 572 646
rect 540 542 572 578
rect 540 474 572 510
rect 540 426 572 442
rect 2516 4024 2548 4398
rect 2516 3956 2548 3992
rect 2516 3888 2548 3924
rect 2516 3820 2548 3856
rect 2516 3752 2548 3788
rect 2516 3684 2548 3720
rect 2516 3616 2548 3652
rect 2516 3548 2548 3584
rect 2516 3480 2548 3516
rect 2516 3412 2548 3448
rect 2516 3344 2548 3380
rect 2516 3276 2548 3312
rect 2516 3208 2548 3244
rect 2516 3140 2548 3176
rect 2516 3072 2548 3108
rect 2516 3004 2548 3040
rect 2516 2936 2548 2972
rect 2516 2868 2548 2904
rect 2516 2800 2548 2836
rect 2516 2732 2548 2768
rect 2516 2664 2548 2700
rect 2516 2596 2548 2632
rect 2516 2528 2548 2564
rect 2516 2460 2548 2496
rect 2516 2392 2548 2428
rect 2516 2324 2548 2360
rect 2516 2174 2548 2292
rect 2516 2106 2548 2142
rect 2516 2038 2548 2074
rect 2516 1970 2548 2006
rect 2516 1902 2548 1938
rect 2516 1834 2548 1870
rect 2516 1766 2548 1802
rect 2516 1698 2548 1734
rect 2516 1630 2548 1666
rect 2516 1562 2548 1598
rect 2516 1494 2548 1530
rect 2516 1426 2548 1462
rect 2516 1358 2548 1394
rect 2516 1290 2548 1326
rect 2516 1222 2548 1258
rect 2516 1154 2548 1190
rect 2516 1086 2548 1122
rect 2516 1018 2548 1054
rect 2516 950 2548 986
rect 2516 882 2548 918
rect 2516 814 2548 850
rect 2516 746 2548 782
rect 2516 678 2548 714
rect 2516 610 2548 646
rect 2516 542 2548 578
rect 2516 474 2548 510
rect 2516 426 2548 442
rect 4492 4024 4524 4398
rect 4492 3956 4524 3992
rect 4492 3888 4524 3924
rect 4492 3820 4524 3856
rect 4492 3752 4524 3788
rect 4492 3684 4524 3720
rect 4492 3616 4524 3652
rect 4492 3548 4524 3584
rect 4492 3480 4524 3516
rect 4492 3412 4524 3448
rect 4492 3344 4524 3380
rect 4492 3276 4524 3312
rect 4492 3208 4524 3244
rect 4492 3140 4524 3176
rect 4492 3072 4524 3108
rect 4492 3004 4524 3040
rect 4492 2936 4524 2972
rect 4492 2868 4524 2904
rect 4492 2800 4524 2836
rect 4492 2732 4524 2768
rect 4492 2664 4524 2700
rect 4492 2596 4524 2632
rect 4492 2528 4524 2564
rect 4492 2460 4524 2496
rect 4492 2392 4524 2428
rect 4492 2324 4524 2360
rect 4492 2174 4524 2292
rect 4492 2106 4524 2142
rect 4492 2038 4524 2074
rect 4492 1970 4524 2006
rect 4492 1902 4524 1938
rect 4492 1834 4524 1870
rect 4492 1766 4524 1802
rect 4492 1698 4524 1734
rect 4492 1630 4524 1666
rect 4492 1562 4524 1598
rect 4492 1494 4524 1530
rect 4492 1426 4524 1462
rect 4492 1358 4524 1394
rect 4492 1290 4524 1326
rect 4492 1222 4524 1258
rect 4492 1154 4524 1190
rect 4492 1086 4524 1122
rect 4492 1018 4524 1054
rect 4492 950 4524 986
rect 4492 882 4524 918
rect 4492 814 4524 850
rect 4492 746 4524 782
rect 4492 678 4524 714
rect 4492 610 4524 646
rect 4492 542 4524 578
rect 4492 474 4524 510
rect 4492 426 4524 442
rect 6468 4024 6500 4398
rect 6468 3956 6500 3992
rect 6468 3888 6500 3924
rect 6468 3820 6500 3856
rect 6468 3752 6500 3788
rect 6468 3684 6500 3720
rect 6468 3616 6500 3652
rect 6468 3548 6500 3584
rect 6468 3480 6500 3516
rect 6468 3412 6500 3448
rect 6468 3344 6500 3380
rect 6468 3276 6500 3312
rect 6468 3208 6500 3244
rect 6468 3140 6500 3176
rect 6468 3072 6500 3108
rect 6468 3004 6500 3040
rect 6468 2936 6500 2972
rect 6468 2868 6500 2904
rect 6468 2800 6500 2836
rect 6468 2732 6500 2768
rect 6468 2664 6500 2700
rect 6468 2596 6500 2632
rect 6468 2528 6500 2564
rect 6468 2460 6500 2496
rect 6468 2392 6500 2428
rect 6468 2324 6500 2360
rect 6468 2174 6500 2292
rect 6468 2106 6500 2142
rect 6468 2038 6500 2074
rect 6468 1970 6500 2006
rect 6468 1902 6500 1938
rect 6468 1834 6500 1870
rect 6468 1766 6500 1802
rect 6468 1698 6500 1734
rect 6468 1630 6500 1666
rect 6468 1562 6500 1598
rect 6468 1494 6500 1530
rect 6468 1426 6500 1462
rect 6468 1358 6500 1394
rect 6468 1290 6500 1326
rect 6468 1222 6500 1258
rect 6468 1154 6500 1190
rect 6468 1086 6500 1122
rect 6468 1018 6500 1054
rect 6468 950 6500 986
rect 6468 882 6500 918
rect 6468 814 6500 850
rect 6468 746 6500 782
rect 6468 678 6500 714
rect 6468 610 6500 646
rect 6468 542 6500 578
rect 6468 474 6500 510
rect 6468 426 6500 442
rect 8444 4024 8476 4398
rect 8444 3956 8476 3992
rect 8444 3888 8476 3924
rect 8444 3820 8476 3856
rect 8444 3752 8476 3788
rect 8444 3684 8476 3720
rect 8444 3616 8476 3652
rect 8444 3548 8476 3584
rect 8444 3480 8476 3516
rect 8444 3412 8476 3448
rect 8444 3344 8476 3380
rect 8444 3276 8476 3312
rect 8444 3208 8476 3244
rect 8444 3140 8476 3176
rect 8444 3072 8476 3108
rect 8444 3004 8476 3040
rect 8444 2936 8476 2972
rect 8444 2868 8476 2904
rect 8444 2800 8476 2836
rect 8444 2732 8476 2768
rect 8444 2664 8476 2700
rect 8444 2596 8476 2632
rect 8444 2528 8476 2564
rect 8444 2460 8476 2496
rect 8444 2392 8476 2428
rect 8444 2324 8476 2360
rect 8444 2174 8476 2292
rect 8444 2106 8476 2142
rect 8444 2038 8476 2074
rect 8444 1970 8476 2006
rect 8444 1902 8476 1938
rect 8444 1834 8476 1870
rect 8444 1766 8476 1802
rect 8444 1698 8476 1734
rect 8444 1630 8476 1666
rect 8444 1562 8476 1598
rect 8444 1494 8476 1530
rect 8444 1426 8476 1462
rect 8444 1358 8476 1394
rect 8444 1290 8476 1326
rect 8444 1222 8476 1258
rect 8444 1154 8476 1190
rect 8444 1086 8476 1122
rect 8444 1018 8476 1054
rect 8444 950 8476 986
rect 8444 882 8476 918
rect 8444 814 8476 850
rect 8444 746 8476 782
rect 8444 678 8476 714
rect 8444 610 8476 646
rect 8444 542 8476 578
rect 8444 474 8476 510
rect 8444 426 8476 442
rect 10420 4024 10452 4398
rect 10420 3956 10452 3992
rect 10420 3888 10452 3924
rect 10420 3820 10452 3856
rect 10420 3752 10452 3788
rect 10420 3684 10452 3720
rect 10420 3616 10452 3652
rect 10420 3548 10452 3584
rect 10420 3480 10452 3516
rect 10420 3412 10452 3448
rect 10420 3344 10452 3380
rect 10420 3276 10452 3312
rect 10420 3208 10452 3244
rect 10420 3140 10452 3176
rect 10420 3072 10452 3108
rect 10420 3004 10452 3040
rect 10420 2936 10452 2972
rect 10420 2868 10452 2904
rect 10420 2800 10452 2836
rect 10420 2732 10452 2768
rect 10420 2664 10452 2700
rect 10420 2596 10452 2632
rect 10420 2528 10452 2564
rect 10420 2460 10452 2496
rect 10420 2392 10452 2428
rect 10420 2324 10452 2360
rect 10420 2174 10452 2292
rect 10420 2106 10452 2142
rect 10420 2038 10452 2074
rect 10420 1970 10452 2006
rect 10420 1902 10452 1938
rect 10420 1834 10452 1870
rect 10420 1766 10452 1802
rect 10420 1698 10452 1734
rect 10420 1630 10452 1666
rect 10420 1562 10452 1598
rect 10420 1494 10452 1530
rect 10420 1426 10452 1462
rect 10420 1358 10452 1394
rect 10420 1290 10452 1326
rect 10420 1222 10452 1258
rect 10420 1154 10452 1190
rect 10420 1086 10452 1122
rect 10420 1018 10452 1054
rect 10420 950 10452 986
rect 10420 882 10452 918
rect 10420 814 10452 850
rect 10420 746 10452 782
rect 10420 678 10452 714
rect 10420 610 10452 646
rect 10420 542 10452 578
rect 10420 474 10452 510
rect 10420 426 10452 442
rect 12396 4024 12428 4398
rect 12396 3956 12428 3992
rect 12396 3888 12428 3924
rect 12396 3820 12428 3856
rect 12396 3752 12428 3788
rect 12396 3684 12428 3720
rect 12396 3616 12428 3652
rect 12396 3548 12428 3584
rect 12396 3480 12428 3516
rect 12396 3412 12428 3448
rect 12396 3344 12428 3380
rect 12396 3276 12428 3312
rect 12396 3208 12428 3244
rect 12396 3140 12428 3176
rect 12396 3072 12428 3108
rect 12396 3004 12428 3040
rect 12396 2936 12428 2972
rect 12396 2868 12428 2904
rect 12396 2800 12428 2836
rect 12396 2732 12428 2768
rect 12396 2664 12428 2700
rect 12396 2596 12428 2632
rect 12396 2528 12428 2564
rect 12396 2460 12428 2496
rect 12396 2392 12428 2428
rect 12396 2324 12428 2360
rect 12396 2174 12428 2292
rect 12396 2106 12428 2142
rect 12396 2038 12428 2074
rect 12396 1970 12428 2006
rect 12396 1902 12428 1938
rect 12396 1834 12428 1870
rect 12396 1766 12428 1802
rect 12396 1698 12428 1734
rect 12396 1630 12428 1666
rect 12396 1562 12428 1598
rect 12396 1494 12428 1530
rect 12396 1426 12428 1462
rect 12396 1358 12428 1394
rect 12396 1290 12428 1326
rect 12396 1222 12428 1258
rect 12396 1154 12428 1190
rect 12396 1086 12428 1122
rect 12396 1018 12428 1054
rect 12396 950 12428 986
rect 12396 882 12428 918
rect 12396 814 12428 850
rect 12396 746 12428 782
rect 12396 678 12428 714
rect 12396 610 12428 646
rect 12396 542 12428 578
rect 12396 474 12428 510
rect 12396 426 12428 442
rect 14372 4024 14404 4398
rect 14372 3956 14404 3992
rect 14372 3888 14404 3924
rect 14372 3820 14404 3856
rect 14372 3752 14404 3788
rect 14372 3684 14404 3720
rect 14372 3616 14404 3652
rect 14372 3548 14404 3584
rect 14372 3480 14404 3516
rect 14372 3412 14404 3448
rect 14372 3344 14404 3380
rect 14372 3276 14404 3312
rect 14372 3208 14404 3244
rect 14372 3140 14404 3176
rect 14372 3072 14404 3108
rect 14372 3004 14404 3040
rect 14372 2936 14404 2972
rect 14372 2868 14404 2904
rect 14372 2800 14404 2836
rect 14372 2732 14404 2768
rect 14372 2664 14404 2700
rect 14372 2596 14404 2632
rect 14372 2528 14404 2564
rect 14372 2460 14404 2496
rect 14372 2392 14404 2428
rect 14372 2324 14404 2360
rect 14372 2174 14404 2292
rect 14543 4024 14585 4040
rect 14543 3998 14548 4024
rect 14580 3998 14585 4024
rect 14543 2318 14544 3998
rect 14584 2318 14585 3998
rect 14543 2292 14548 2318
rect 14580 2292 14585 2318
rect 14543 2276 14585 2292
rect 14724 4024 14756 4398
rect 14724 3956 14756 3992
rect 14724 3888 14756 3924
rect 14724 3820 14756 3856
rect 14724 3752 14756 3788
rect 14724 3684 14756 3720
rect 14724 3616 14756 3652
rect 14724 3548 14756 3584
rect 14724 3480 14756 3516
rect 14724 3412 14756 3448
rect 14724 3344 14756 3380
rect 14724 3276 14756 3312
rect 14724 3208 14756 3244
rect 14724 3140 14756 3176
rect 14724 3072 14756 3108
rect 14724 3004 14756 3040
rect 14724 2936 14756 2972
rect 14724 2868 14756 2904
rect 14724 2800 14756 2836
rect 14724 2732 14756 2768
rect 14724 2664 14756 2700
rect 14724 2596 14756 2632
rect 14724 2528 14756 2564
rect 14724 2460 14756 2496
rect 14724 2392 14756 2428
rect 14724 2324 14756 2360
rect 14372 2106 14404 2142
rect 14372 2038 14404 2074
rect 14372 1970 14404 2006
rect 14372 1902 14404 1938
rect 14372 1834 14404 1870
rect 14372 1766 14404 1802
rect 14372 1698 14404 1734
rect 14372 1630 14404 1666
rect 14372 1562 14404 1598
rect 14372 1494 14404 1530
rect 14372 1426 14404 1462
rect 14372 1358 14404 1394
rect 14372 1290 14404 1326
rect 14372 1222 14404 1258
rect 14372 1154 14404 1190
rect 14372 1086 14404 1122
rect 14372 1018 14404 1054
rect 14372 950 14404 986
rect 14372 882 14404 918
rect 14372 814 14404 850
rect 14372 746 14404 782
rect 14372 678 14404 714
rect 14372 610 14404 646
rect 14372 542 14404 578
rect 14372 474 14404 510
rect 14372 426 14404 442
rect 14543 2174 14585 2190
rect 14543 2148 14548 2174
rect 14580 2148 14585 2174
rect 14543 468 14544 2148
rect 14584 468 14585 2148
rect 14543 442 14548 468
rect 14580 442 14585 468
rect 14543 426 14585 442
rect 14724 2174 14756 2292
rect 14895 4024 14937 4040
rect 14895 3998 14900 4024
rect 14932 3998 14937 4024
rect 14895 2318 14896 3998
rect 14936 2318 14937 3998
rect 14895 2292 14900 2318
rect 14932 2292 14937 2318
rect 14895 2276 14937 2292
rect 15076 4024 15108 4398
rect 15076 3956 15108 3992
rect 15076 3888 15108 3924
rect 15076 3820 15108 3856
rect 15076 3752 15108 3788
rect 15076 3684 15108 3720
rect 15076 3616 15108 3652
rect 15076 3548 15108 3584
rect 15076 3480 15108 3516
rect 15076 3412 15108 3448
rect 15076 3344 15108 3380
rect 15076 3276 15108 3312
rect 15076 3208 15108 3244
rect 15076 3140 15108 3176
rect 15076 3072 15108 3108
rect 15076 3004 15108 3040
rect 15076 2936 15108 2972
rect 15076 2868 15108 2904
rect 15076 2800 15108 2836
rect 15076 2732 15108 2768
rect 15076 2664 15108 2700
rect 15076 2596 15108 2632
rect 15076 2528 15108 2564
rect 15076 2460 15108 2496
rect 15076 2392 15108 2428
rect 15076 2324 15108 2360
rect 14724 2106 14756 2142
rect 14724 2038 14756 2074
rect 14724 1970 14756 2006
rect 14724 1902 14756 1938
rect 14724 1834 14756 1870
rect 14724 1766 14756 1802
rect 14724 1698 14756 1734
rect 14724 1630 14756 1666
rect 14724 1562 14756 1598
rect 14724 1494 14756 1530
rect 14724 1426 14756 1462
rect 14724 1358 14756 1394
rect 14724 1290 14756 1326
rect 14724 1222 14756 1258
rect 14724 1154 14756 1190
rect 14724 1086 14756 1122
rect 14724 1018 14756 1054
rect 14724 950 14756 986
rect 14724 882 14756 918
rect 14724 814 14756 850
rect 14724 746 14756 782
rect 14724 678 14756 714
rect 14724 610 14756 646
rect 14724 542 14756 578
rect 14724 474 14756 510
rect 14724 426 14756 442
rect 14895 2174 14937 2190
rect 14895 2148 14900 2174
rect 14932 2148 14937 2174
rect 14895 468 14896 2148
rect 14936 468 14937 2148
rect 14895 442 14900 468
rect 14932 442 14937 468
rect 14895 426 14937 442
rect 15076 2174 15108 2292
rect 15247 4024 15289 4040
rect 15247 3998 15252 4024
rect 15284 3998 15289 4024
rect 15247 2318 15248 3998
rect 15288 2318 15289 3998
rect 15247 2292 15252 2318
rect 15284 2292 15289 2318
rect 15247 2276 15289 2292
rect 15428 4024 15460 4398
rect 15428 3956 15460 3992
rect 15428 3888 15460 3924
rect 15428 3820 15460 3856
rect 15428 3752 15460 3788
rect 15428 3684 15460 3720
rect 15428 3616 15460 3652
rect 15428 3548 15460 3584
rect 15428 3480 15460 3516
rect 15428 3412 15460 3448
rect 15428 3344 15460 3380
rect 15428 3276 15460 3312
rect 15428 3208 15460 3244
rect 15428 3140 15460 3176
rect 15428 3072 15460 3108
rect 15428 3004 15460 3040
rect 15428 2936 15460 2972
rect 15428 2868 15460 2904
rect 15428 2800 15460 2836
rect 15428 2732 15460 2768
rect 15428 2664 15460 2700
rect 15428 2596 15460 2632
rect 15428 2528 15460 2564
rect 15428 2460 15460 2496
rect 15428 2392 15460 2428
rect 15428 2324 15460 2360
rect 15076 2106 15108 2142
rect 15076 2038 15108 2074
rect 15076 1970 15108 2006
rect 15076 1902 15108 1938
rect 15076 1834 15108 1870
rect 15076 1766 15108 1802
rect 15076 1698 15108 1734
rect 15076 1630 15108 1666
rect 15076 1562 15108 1598
rect 15076 1494 15108 1530
rect 15076 1426 15108 1462
rect 15076 1358 15108 1394
rect 15076 1290 15108 1326
rect 15076 1222 15108 1258
rect 15076 1154 15108 1190
rect 15076 1086 15108 1122
rect 15076 1018 15108 1054
rect 15076 950 15108 986
rect 15076 882 15108 918
rect 15076 814 15108 850
rect 15076 746 15108 782
rect 15076 678 15108 714
rect 15076 610 15108 646
rect 15076 542 15108 578
rect 15076 474 15108 510
rect 15076 426 15108 442
rect 15247 2174 15289 2190
rect 15247 2148 15252 2174
rect 15284 2148 15289 2174
rect 15247 468 15248 2148
rect 15288 468 15289 2148
rect 15247 442 15252 468
rect 15284 442 15289 468
rect 15247 426 15289 442
rect 15428 2174 15460 2292
rect 15428 2106 15460 2142
rect 15428 2038 15460 2074
rect 15428 1970 15460 2006
rect 15428 1902 15460 1938
rect 15428 1834 15460 1870
rect 15428 1766 15460 1802
rect 15428 1698 15460 1734
rect 15428 1630 15460 1666
rect 15428 1562 15460 1598
rect 15428 1494 15460 1530
rect 15428 1426 15460 1462
rect 15428 1358 15460 1394
rect 15428 1290 15460 1326
rect 15428 1222 15460 1258
rect 15428 1154 15460 1190
rect 15428 1086 15460 1122
rect 15428 1018 15460 1054
rect 15428 950 15460 986
rect 15428 882 15460 918
rect 15428 814 15460 850
rect 15428 746 15460 782
rect 15428 678 15460 714
rect 15428 610 15460 646
rect 15428 542 15460 578
rect 15428 474 15460 510
rect 15428 426 15460 442
rect 15932 4357 16000 4398
rect 15932 4325 15950 4357
rect 15982 4325 16000 4357
rect 15932 4289 16000 4325
rect 15932 4257 15950 4289
rect 15982 4257 16000 4289
rect 15932 4221 16000 4257
rect 15932 4189 15950 4221
rect 15982 4189 16000 4221
rect 15932 4153 16000 4189
rect 15932 4121 15950 4153
rect 15982 4121 16000 4153
rect 15932 4085 16000 4121
rect 15932 4053 15950 4085
rect 15982 4053 16000 4085
rect 15932 4017 16000 4053
rect 15932 3985 15950 4017
rect 15982 3985 16000 4017
rect 15932 3949 16000 3985
rect 15932 3917 15950 3949
rect 15982 3917 16000 3949
rect 15932 3881 16000 3917
rect 15932 3849 15950 3881
rect 15982 3849 16000 3881
rect 15932 3813 16000 3849
rect 15932 3781 15950 3813
rect 15982 3781 16000 3813
rect 15932 3745 16000 3781
rect 15932 3713 15950 3745
rect 15982 3713 16000 3745
rect 15932 3677 16000 3713
rect 15932 3645 15950 3677
rect 15982 3645 16000 3677
rect 15932 3609 16000 3645
rect 15932 3577 15950 3609
rect 15982 3577 16000 3609
rect 15932 3541 16000 3577
rect 15932 3509 15950 3541
rect 15982 3509 16000 3541
rect 15932 3473 16000 3509
rect 15932 3441 15950 3473
rect 15982 3441 16000 3473
rect 15932 3405 16000 3441
rect 15932 3373 15950 3405
rect 15982 3373 16000 3405
rect 15932 3337 16000 3373
rect 15932 3305 15950 3337
rect 15982 3305 16000 3337
rect 15932 3269 16000 3305
rect 15932 3237 15950 3269
rect 15982 3237 16000 3269
rect 15932 3201 16000 3237
rect 15932 3169 15950 3201
rect 15982 3169 16000 3201
rect 15932 3133 16000 3169
rect 15932 3101 15950 3133
rect 15982 3101 16000 3133
rect 15932 3065 16000 3101
rect 15932 3033 15950 3065
rect 15982 3033 16000 3065
rect 15932 2997 16000 3033
rect 15932 2965 15950 2997
rect 15982 2965 16000 2997
rect 15932 2929 16000 2965
rect 15932 2897 15950 2929
rect 15982 2897 16000 2929
rect 15932 2861 16000 2897
rect 15932 2829 15950 2861
rect 15982 2829 16000 2861
rect 15932 2793 16000 2829
rect 15932 2761 15950 2793
rect 15982 2761 16000 2793
rect 15932 2725 16000 2761
rect 15932 2693 15950 2725
rect 15982 2693 16000 2725
rect 15932 2657 16000 2693
rect 15932 2625 15950 2657
rect 15982 2625 16000 2657
rect 15932 2589 16000 2625
rect 15932 2557 15950 2589
rect 15982 2557 16000 2589
rect 15932 2521 16000 2557
rect 15932 2489 15950 2521
rect 15982 2489 16000 2521
rect 15932 2453 16000 2489
rect 15932 2421 15950 2453
rect 15982 2421 16000 2453
rect 15932 2385 16000 2421
rect 15932 2353 15950 2385
rect 15982 2353 16000 2385
rect 15932 2317 16000 2353
rect 15932 2285 15950 2317
rect 15982 2285 16000 2317
rect 15932 2249 16000 2285
rect 15932 2217 15950 2249
rect 15982 2217 16000 2249
rect 15932 2181 16000 2217
rect 15932 2149 15950 2181
rect 15982 2149 16000 2181
rect 15932 2113 16000 2149
rect 15932 2081 15950 2113
rect 15982 2081 16000 2113
rect 15932 2045 16000 2081
rect 15932 2013 15950 2045
rect 15982 2013 16000 2045
rect 15932 1977 16000 2013
rect 15932 1945 15950 1977
rect 15982 1945 16000 1977
rect 15932 1909 16000 1945
rect 15932 1877 15950 1909
rect 15982 1877 16000 1909
rect 15932 1841 16000 1877
rect 15932 1809 15950 1841
rect 15982 1809 16000 1841
rect 15932 1773 16000 1809
rect 15932 1741 15950 1773
rect 15982 1741 16000 1773
rect 15932 1705 16000 1741
rect 15932 1673 15950 1705
rect 15982 1673 16000 1705
rect 15932 1637 16000 1673
rect 15932 1605 15950 1637
rect 15982 1605 16000 1637
rect 15932 1569 16000 1605
rect 15932 1537 15950 1569
rect 15982 1537 16000 1569
rect 15932 1501 16000 1537
rect 15932 1469 15950 1501
rect 15982 1469 16000 1501
rect 15932 1433 16000 1469
rect 15932 1401 15950 1433
rect 15982 1401 16000 1433
rect 15932 1365 16000 1401
rect 15932 1333 15950 1365
rect 15982 1333 16000 1365
rect 15932 1297 16000 1333
rect 15932 1265 15950 1297
rect 15982 1265 16000 1297
rect 15932 1229 16000 1265
rect 15932 1197 15950 1229
rect 15982 1197 16000 1229
rect 15932 1161 16000 1197
rect 15932 1129 15950 1161
rect 15982 1129 16000 1161
rect 15932 1093 16000 1129
rect 15932 1061 15950 1093
rect 15982 1061 16000 1093
rect 15932 1025 16000 1061
rect 15932 993 15950 1025
rect 15982 993 16000 1025
rect 15932 957 16000 993
rect 15932 925 15950 957
rect 15982 925 16000 957
rect 15932 889 16000 925
rect 15932 857 15950 889
rect 15982 857 16000 889
rect 15932 821 16000 857
rect 15932 789 15950 821
rect 15982 789 16000 821
rect 15932 753 16000 789
rect 15932 721 15950 753
rect 15982 721 16000 753
rect 15932 685 16000 721
rect 15932 653 15950 685
rect 15982 653 16000 685
rect 15932 617 16000 653
rect 15932 585 15950 617
rect 15982 585 16000 617
rect 15932 549 16000 585
rect 15932 517 15950 549
rect 15982 517 16000 549
rect 15932 481 16000 517
rect 15932 449 15950 481
rect 15982 449 16000 481
rect 0 381 18 413
rect 50 381 68 413
rect 0 345 68 381
rect 15932 413 16000 449
rect 15932 381 15950 413
rect 15982 381 16000 413
rect 0 313 18 345
rect 50 313 68 345
rect 0 277 68 313
rect 594 348 640 380
rect 672 348 708 380
rect 740 348 776 380
rect 808 348 844 380
rect 876 348 912 380
rect 944 348 980 380
rect 1012 348 1048 380
rect 1080 348 1116 380
rect 1148 348 1184 380
rect 1216 348 1252 380
rect 1284 348 1320 380
rect 1352 348 1388 380
rect 1420 348 1456 380
rect 1488 348 1524 380
rect 1556 348 1592 380
rect 1624 348 1660 380
rect 1692 348 1728 380
rect 1760 348 1796 380
rect 1828 348 1864 380
rect 1896 348 1932 380
rect 1964 348 2000 380
rect 2032 348 2068 380
rect 2100 348 2136 380
rect 2168 348 2204 380
rect 2236 348 2272 380
rect 2304 348 2340 380
rect 2372 348 2408 380
rect 2440 348 2476 380
rect 2508 348 2544 380
rect 2576 348 2612 380
rect 2644 348 2680 380
rect 2712 348 2748 380
rect 2780 348 2816 380
rect 2848 348 2884 380
rect 2916 348 2952 380
rect 2984 348 3020 380
rect 3052 348 3088 380
rect 3120 348 3156 380
rect 3188 348 3224 380
rect 3256 348 3292 380
rect 3324 348 3360 380
rect 3392 348 3428 380
rect 3460 348 3496 380
rect 3528 348 3564 380
rect 3596 348 3632 380
rect 3664 348 3700 380
rect 3732 348 3768 380
rect 3800 348 3836 380
rect 3868 348 3904 380
rect 3936 348 3972 380
rect 4004 348 4040 380
rect 4072 348 4108 380
rect 4140 348 4176 380
rect 4208 348 4244 380
rect 4276 348 4312 380
rect 4344 348 4380 380
rect 4412 348 4448 380
rect 4480 348 4516 380
rect 4548 348 4584 380
rect 4616 348 4652 380
rect 4684 348 4720 380
rect 4752 348 4788 380
rect 4820 348 4856 380
rect 4888 348 4924 380
rect 4956 348 4992 380
rect 5024 348 5060 380
rect 5092 348 5128 380
rect 5160 348 5196 380
rect 5228 348 5264 380
rect 5296 348 5332 380
rect 5364 348 5400 380
rect 5432 348 5468 380
rect 5500 348 5536 380
rect 5568 348 5604 380
rect 5636 348 5672 380
rect 5704 348 5740 380
rect 5772 348 5808 380
rect 5840 348 5876 380
rect 5908 348 5944 380
rect 5976 348 6012 380
rect 6044 348 6080 380
rect 6112 348 6148 380
rect 6180 348 6216 380
rect 6248 348 6284 380
rect 6316 348 6352 380
rect 6384 348 6420 380
rect 6452 348 6488 380
rect 6520 348 6556 380
rect 6588 348 6624 380
rect 6656 348 6692 380
rect 6724 348 6760 380
rect 6792 348 6828 380
rect 6860 348 6896 380
rect 6928 348 6964 380
rect 6996 348 7032 380
rect 7064 348 7100 380
rect 7132 348 7168 380
rect 7200 348 7236 380
rect 7268 348 7304 380
rect 7336 348 7372 380
rect 7404 348 7440 380
rect 7472 348 7508 380
rect 7540 348 7576 380
rect 7608 348 7644 380
rect 7676 348 7712 380
rect 7744 348 7780 380
rect 7812 348 7848 380
rect 7880 348 7916 380
rect 7948 348 7984 380
rect 8016 348 8052 380
rect 8084 348 8120 380
rect 8152 348 8188 380
rect 8220 348 8256 380
rect 8288 348 8324 380
rect 8356 348 8392 380
rect 8424 348 8460 380
rect 8492 348 8528 380
rect 8560 348 8596 380
rect 8628 348 8664 380
rect 8696 348 8732 380
rect 8764 348 8800 380
rect 8832 348 8868 380
rect 8900 348 8936 380
rect 8968 348 9004 380
rect 9036 348 9072 380
rect 9104 348 9140 380
rect 9172 348 9208 380
rect 9240 348 9276 380
rect 9308 348 9344 380
rect 9376 348 9412 380
rect 9444 348 9480 380
rect 9512 348 9548 380
rect 9580 348 9616 380
rect 9648 348 9684 380
rect 9716 348 9752 380
rect 9784 348 9820 380
rect 9852 348 9888 380
rect 9920 348 9956 380
rect 9988 348 10024 380
rect 10056 348 10092 380
rect 10124 348 10160 380
rect 10192 348 10228 380
rect 10260 348 10296 380
rect 10328 348 10364 380
rect 10396 348 10432 380
rect 10464 348 10500 380
rect 10532 348 10568 380
rect 10600 348 10636 380
rect 10668 348 10704 380
rect 10736 348 10772 380
rect 10804 348 10840 380
rect 10872 348 10908 380
rect 10940 348 10976 380
rect 11008 348 11044 380
rect 11076 348 11112 380
rect 11144 348 11180 380
rect 11212 348 11248 380
rect 11280 348 11316 380
rect 11348 348 11384 380
rect 11416 348 11452 380
rect 11484 348 11520 380
rect 11552 348 11588 380
rect 11620 348 11656 380
rect 11688 348 11724 380
rect 11756 348 11792 380
rect 11824 348 11860 380
rect 11892 348 11928 380
rect 11960 348 11996 380
rect 12028 348 12064 380
rect 12096 348 12132 380
rect 12164 348 12200 380
rect 12232 348 12268 380
rect 12300 348 12336 380
rect 12368 348 12404 380
rect 12436 348 12472 380
rect 12504 348 12540 380
rect 12572 348 12608 380
rect 12640 348 12676 380
rect 12708 348 12744 380
rect 12776 348 12812 380
rect 12844 348 12880 380
rect 12912 348 12948 380
rect 12980 348 13016 380
rect 13048 348 13084 380
rect 13116 348 13152 380
rect 13184 348 13220 380
rect 13252 348 13288 380
rect 13320 348 13356 380
rect 13388 348 13424 380
rect 13456 348 13492 380
rect 13524 348 13560 380
rect 13592 348 13628 380
rect 13660 348 13696 380
rect 13728 348 13764 380
rect 13796 348 13832 380
rect 13864 348 13900 380
rect 13932 348 13968 380
rect 14000 348 14036 380
rect 14068 348 14104 380
rect 14136 348 14172 380
rect 14204 348 14240 380
rect 14272 348 14308 380
rect 14340 348 14376 380
rect 14408 348 14444 380
rect 14476 348 14512 380
rect 14544 348 14580 380
rect 14612 348 14648 380
rect 14680 348 14716 380
rect 14748 348 14784 380
rect 14816 348 14852 380
rect 14884 348 14920 380
rect 14952 348 14988 380
rect 15020 348 15056 380
rect 15088 348 15124 380
rect 15156 348 15192 380
rect 15224 348 15260 380
rect 15292 348 15328 380
rect 15360 348 15406 380
rect 594 342 15406 348
rect 594 302 641 342
rect 15359 302 15406 342
rect 594 301 15406 302
rect 15932 345 16000 381
rect 15932 313 15950 345
rect 15982 313 16000 345
rect 0 245 18 277
rect 50 245 68 277
rect 0 209 68 245
rect 0 177 18 209
rect 50 177 68 209
rect 0 141 68 177
rect 0 109 18 141
rect 50 109 68 141
rect 0 68 68 109
rect 15932 277 16000 313
rect 15932 245 15950 277
rect 15982 245 16000 277
rect 15932 209 16000 245
rect 15932 177 15950 209
rect 15982 177 16000 209
rect 15932 141 16000 177
rect 15932 109 15950 141
rect 15982 109 16000 141
rect 15932 68 16000 109
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 3675 6744 12325 6784
rect 3756 6612 3760 6617
rect 3760 6612 3792 6617
rect 3792 6612 3796 6617
rect 3756 6576 3796 6612
rect 3756 6544 3760 6576
rect 3760 6544 3792 6576
rect 3792 6544 3796 6576
rect 3756 6508 3796 6544
rect 3756 6476 3760 6508
rect 3760 6476 3792 6508
rect 3792 6476 3796 6508
rect 3756 6440 3796 6476
rect 3756 6408 3760 6440
rect 3760 6408 3792 6440
rect 3792 6408 3796 6440
rect 3756 6372 3796 6408
rect 3756 6340 3760 6372
rect 3760 6340 3792 6372
rect 3792 6340 3796 6372
rect 3756 6304 3796 6340
rect 3756 6272 3760 6304
rect 3760 6272 3792 6304
rect 3792 6272 3796 6304
rect 3756 6236 3796 6272
rect 3756 6204 3760 6236
rect 3760 6204 3792 6236
rect 3792 6204 3796 6236
rect 3756 6168 3796 6204
rect 3756 6136 3760 6168
rect 3760 6136 3792 6168
rect 3792 6136 3796 6168
rect 3756 6100 3796 6136
rect 3756 6068 3760 6100
rect 3760 6068 3792 6100
rect 3792 6068 3796 6100
rect 3756 6032 3796 6068
rect 3756 6000 3760 6032
rect 3760 6000 3792 6032
rect 3792 6000 3796 6032
rect 3756 5964 3796 6000
rect 3756 5932 3760 5964
rect 3760 5932 3792 5964
rect 3792 5932 3796 5964
rect 3756 5896 3796 5932
rect 3756 5864 3760 5896
rect 3760 5864 3792 5896
rect 3792 5864 3796 5896
rect 3756 5828 3796 5864
rect 3756 5796 3760 5828
rect 3760 5796 3792 5828
rect 3792 5796 3796 5828
rect 3756 5760 3796 5796
rect 3756 5728 3760 5760
rect 3760 5728 3792 5760
rect 3792 5728 3796 5760
rect 3756 5692 3796 5728
rect 3756 5660 3760 5692
rect 3760 5660 3792 5692
rect 3792 5660 3796 5692
rect 3756 5624 3796 5660
rect 3756 5592 3760 5624
rect 3760 5592 3792 5624
rect 3792 5592 3796 5624
rect 3756 5556 3796 5592
rect 3756 5524 3760 5556
rect 3760 5524 3792 5556
rect 3792 5524 3796 5556
rect 3756 5488 3796 5524
rect 3756 5456 3760 5488
rect 3760 5456 3792 5488
rect 3792 5456 3796 5488
rect 3756 5420 3796 5456
rect 3756 5388 3760 5420
rect 3760 5388 3792 5420
rect 3792 5388 3796 5420
rect 3756 5352 3796 5388
rect 3756 5347 3760 5352
rect 3760 5347 3792 5352
rect 3792 5347 3796 5352
rect 4108 6612 4112 6617
rect 4112 6612 4144 6617
rect 4144 6612 4148 6617
rect 4108 6576 4148 6612
rect 4108 6544 4112 6576
rect 4112 6544 4144 6576
rect 4144 6544 4148 6576
rect 4108 6508 4148 6544
rect 4108 6476 4112 6508
rect 4112 6476 4144 6508
rect 4144 6476 4148 6508
rect 4108 6440 4148 6476
rect 4108 6408 4112 6440
rect 4112 6408 4144 6440
rect 4144 6408 4148 6440
rect 4108 6372 4148 6408
rect 4108 6340 4112 6372
rect 4112 6340 4144 6372
rect 4144 6340 4148 6372
rect 4108 6304 4148 6340
rect 4108 6272 4112 6304
rect 4112 6272 4144 6304
rect 4144 6272 4148 6304
rect 4108 6236 4148 6272
rect 4108 6204 4112 6236
rect 4112 6204 4144 6236
rect 4144 6204 4148 6236
rect 4108 6168 4148 6204
rect 4108 6136 4112 6168
rect 4112 6136 4144 6168
rect 4144 6136 4148 6168
rect 4108 6100 4148 6136
rect 4108 6068 4112 6100
rect 4112 6068 4144 6100
rect 4144 6068 4148 6100
rect 4108 6032 4148 6068
rect 4108 6000 4112 6032
rect 4112 6000 4144 6032
rect 4144 6000 4148 6032
rect 4108 5964 4148 6000
rect 4108 5932 4112 5964
rect 4112 5932 4144 5964
rect 4144 5932 4148 5964
rect 4108 5896 4148 5932
rect 4108 5864 4112 5896
rect 4112 5864 4144 5896
rect 4144 5864 4148 5896
rect 4108 5828 4148 5864
rect 4108 5796 4112 5828
rect 4112 5796 4144 5828
rect 4144 5796 4148 5828
rect 4108 5760 4148 5796
rect 4108 5728 4112 5760
rect 4112 5728 4144 5760
rect 4144 5728 4148 5760
rect 4108 5692 4148 5728
rect 4108 5660 4112 5692
rect 4112 5660 4144 5692
rect 4144 5660 4148 5692
rect 4108 5624 4148 5660
rect 4108 5592 4112 5624
rect 4112 5592 4144 5624
rect 4144 5592 4148 5624
rect 4108 5556 4148 5592
rect 4108 5524 4112 5556
rect 4112 5524 4144 5556
rect 4144 5524 4148 5556
rect 4108 5488 4148 5524
rect 4108 5456 4112 5488
rect 4112 5456 4144 5488
rect 4144 5456 4148 5488
rect 4108 5420 4148 5456
rect 4108 5388 4112 5420
rect 4112 5388 4144 5420
rect 4144 5388 4148 5420
rect 4108 5352 4148 5388
rect 4108 5347 4112 5352
rect 4112 5347 4144 5352
rect 4144 5347 4148 5352
rect 4460 6612 4464 6617
rect 4464 6612 4496 6617
rect 4496 6612 4500 6617
rect 4460 6576 4500 6612
rect 4460 6544 4464 6576
rect 4464 6544 4496 6576
rect 4496 6544 4500 6576
rect 4460 6508 4500 6544
rect 4460 6476 4464 6508
rect 4464 6476 4496 6508
rect 4496 6476 4500 6508
rect 4460 6440 4500 6476
rect 4460 6408 4464 6440
rect 4464 6408 4496 6440
rect 4496 6408 4500 6440
rect 4460 6372 4500 6408
rect 4460 6340 4464 6372
rect 4464 6340 4496 6372
rect 4496 6340 4500 6372
rect 4460 6304 4500 6340
rect 4460 6272 4464 6304
rect 4464 6272 4496 6304
rect 4496 6272 4500 6304
rect 4460 6236 4500 6272
rect 4460 6204 4464 6236
rect 4464 6204 4496 6236
rect 4496 6204 4500 6236
rect 4460 6168 4500 6204
rect 4460 6136 4464 6168
rect 4464 6136 4496 6168
rect 4496 6136 4500 6168
rect 4460 6100 4500 6136
rect 4460 6068 4464 6100
rect 4464 6068 4496 6100
rect 4496 6068 4500 6100
rect 4460 6032 4500 6068
rect 4460 6000 4464 6032
rect 4464 6000 4496 6032
rect 4496 6000 4500 6032
rect 4460 5964 4500 6000
rect 4460 5932 4464 5964
rect 4464 5932 4496 5964
rect 4496 5932 4500 5964
rect 4460 5896 4500 5932
rect 4460 5864 4464 5896
rect 4464 5864 4496 5896
rect 4496 5864 4500 5896
rect 4460 5828 4500 5864
rect 4460 5796 4464 5828
rect 4464 5796 4496 5828
rect 4496 5796 4500 5828
rect 4460 5760 4500 5796
rect 4460 5728 4464 5760
rect 4464 5728 4496 5760
rect 4496 5728 4500 5760
rect 4460 5692 4500 5728
rect 4460 5660 4464 5692
rect 4464 5660 4496 5692
rect 4496 5660 4500 5692
rect 4460 5624 4500 5660
rect 4460 5592 4464 5624
rect 4464 5592 4496 5624
rect 4496 5592 4500 5624
rect 4460 5556 4500 5592
rect 4460 5524 4464 5556
rect 4464 5524 4496 5556
rect 4496 5524 4500 5556
rect 4460 5488 4500 5524
rect 4460 5456 4464 5488
rect 4464 5456 4496 5488
rect 4496 5456 4500 5488
rect 4460 5420 4500 5456
rect 4460 5388 4464 5420
rect 4464 5388 4496 5420
rect 4496 5388 4500 5420
rect 4460 5352 4500 5388
rect 4460 5347 4464 5352
rect 4464 5347 4496 5352
rect 4496 5347 4500 5352
rect 4812 6612 4816 6617
rect 4816 6612 4848 6617
rect 4848 6612 4852 6617
rect 4812 6576 4852 6612
rect 4812 6544 4816 6576
rect 4816 6544 4848 6576
rect 4848 6544 4852 6576
rect 4812 6508 4852 6544
rect 4812 6476 4816 6508
rect 4816 6476 4848 6508
rect 4848 6476 4852 6508
rect 4812 6440 4852 6476
rect 4812 6408 4816 6440
rect 4816 6408 4848 6440
rect 4848 6408 4852 6440
rect 4812 6372 4852 6408
rect 4812 6340 4816 6372
rect 4816 6340 4848 6372
rect 4848 6340 4852 6372
rect 4812 6304 4852 6340
rect 4812 6272 4816 6304
rect 4816 6272 4848 6304
rect 4848 6272 4852 6304
rect 4812 6236 4852 6272
rect 4812 6204 4816 6236
rect 4816 6204 4848 6236
rect 4848 6204 4852 6236
rect 4812 6168 4852 6204
rect 4812 6136 4816 6168
rect 4816 6136 4848 6168
rect 4848 6136 4852 6168
rect 4812 6100 4852 6136
rect 4812 6068 4816 6100
rect 4816 6068 4848 6100
rect 4848 6068 4852 6100
rect 4812 6032 4852 6068
rect 4812 6000 4816 6032
rect 4816 6000 4848 6032
rect 4848 6000 4852 6032
rect 4812 5964 4852 6000
rect 4812 5932 4816 5964
rect 4816 5932 4848 5964
rect 4848 5932 4852 5964
rect 4812 5896 4852 5932
rect 4812 5864 4816 5896
rect 4816 5864 4848 5896
rect 4848 5864 4852 5896
rect 4812 5828 4852 5864
rect 4812 5796 4816 5828
rect 4816 5796 4848 5828
rect 4848 5796 4852 5828
rect 4812 5760 4852 5796
rect 4812 5728 4816 5760
rect 4816 5728 4848 5760
rect 4848 5728 4852 5760
rect 4812 5692 4852 5728
rect 4812 5660 4816 5692
rect 4816 5660 4848 5692
rect 4848 5660 4852 5692
rect 4812 5624 4852 5660
rect 4812 5592 4816 5624
rect 4816 5592 4848 5624
rect 4848 5592 4852 5624
rect 4812 5556 4852 5592
rect 4812 5524 4816 5556
rect 4816 5524 4848 5556
rect 4848 5524 4852 5556
rect 4812 5488 4852 5524
rect 4812 5456 4816 5488
rect 4816 5456 4848 5488
rect 4848 5456 4852 5488
rect 4812 5420 4852 5456
rect 4812 5388 4816 5420
rect 4816 5388 4848 5420
rect 4848 5388 4852 5420
rect 4812 5352 4852 5388
rect 4812 5347 4816 5352
rect 4816 5347 4848 5352
rect 4848 5347 4852 5352
rect 5164 6612 5168 6617
rect 5168 6612 5200 6617
rect 5200 6612 5204 6617
rect 5164 6576 5204 6612
rect 5164 6544 5168 6576
rect 5168 6544 5200 6576
rect 5200 6544 5204 6576
rect 5164 6508 5204 6544
rect 5164 6476 5168 6508
rect 5168 6476 5200 6508
rect 5200 6476 5204 6508
rect 5164 6440 5204 6476
rect 5164 6408 5168 6440
rect 5168 6408 5200 6440
rect 5200 6408 5204 6440
rect 5164 6372 5204 6408
rect 5164 6340 5168 6372
rect 5168 6340 5200 6372
rect 5200 6340 5204 6372
rect 5164 6304 5204 6340
rect 5164 6272 5168 6304
rect 5168 6272 5200 6304
rect 5200 6272 5204 6304
rect 5164 6236 5204 6272
rect 5164 6204 5168 6236
rect 5168 6204 5200 6236
rect 5200 6204 5204 6236
rect 5164 6168 5204 6204
rect 5164 6136 5168 6168
rect 5168 6136 5200 6168
rect 5200 6136 5204 6168
rect 5164 6100 5204 6136
rect 5164 6068 5168 6100
rect 5168 6068 5200 6100
rect 5200 6068 5204 6100
rect 5164 6032 5204 6068
rect 5164 6000 5168 6032
rect 5168 6000 5200 6032
rect 5200 6000 5204 6032
rect 5164 5964 5204 6000
rect 5164 5932 5168 5964
rect 5168 5932 5200 5964
rect 5200 5932 5204 5964
rect 5164 5896 5204 5932
rect 5164 5864 5168 5896
rect 5168 5864 5200 5896
rect 5200 5864 5204 5896
rect 5164 5828 5204 5864
rect 5164 5796 5168 5828
rect 5168 5796 5200 5828
rect 5200 5796 5204 5828
rect 5164 5760 5204 5796
rect 5164 5728 5168 5760
rect 5168 5728 5200 5760
rect 5200 5728 5204 5760
rect 5164 5692 5204 5728
rect 5164 5660 5168 5692
rect 5168 5660 5200 5692
rect 5200 5660 5204 5692
rect 5164 5624 5204 5660
rect 5164 5592 5168 5624
rect 5168 5592 5200 5624
rect 5200 5592 5204 5624
rect 5164 5556 5204 5592
rect 5164 5524 5168 5556
rect 5168 5524 5200 5556
rect 5200 5524 5204 5556
rect 5164 5488 5204 5524
rect 5164 5456 5168 5488
rect 5168 5456 5200 5488
rect 5200 5456 5204 5488
rect 5164 5420 5204 5456
rect 5164 5388 5168 5420
rect 5168 5388 5200 5420
rect 5200 5388 5204 5420
rect 5164 5352 5204 5388
rect 5164 5347 5168 5352
rect 5168 5347 5200 5352
rect 5200 5347 5204 5352
rect 5516 6612 5520 6617
rect 5520 6612 5552 6617
rect 5552 6612 5556 6617
rect 5516 6576 5556 6612
rect 5516 6544 5520 6576
rect 5520 6544 5552 6576
rect 5552 6544 5556 6576
rect 5516 6508 5556 6544
rect 5516 6476 5520 6508
rect 5520 6476 5552 6508
rect 5552 6476 5556 6508
rect 5516 6440 5556 6476
rect 5516 6408 5520 6440
rect 5520 6408 5552 6440
rect 5552 6408 5556 6440
rect 5516 6372 5556 6408
rect 5516 6340 5520 6372
rect 5520 6340 5552 6372
rect 5552 6340 5556 6372
rect 5516 6304 5556 6340
rect 5516 6272 5520 6304
rect 5520 6272 5552 6304
rect 5552 6272 5556 6304
rect 5516 6236 5556 6272
rect 5516 6204 5520 6236
rect 5520 6204 5552 6236
rect 5552 6204 5556 6236
rect 5516 6168 5556 6204
rect 5516 6136 5520 6168
rect 5520 6136 5552 6168
rect 5552 6136 5556 6168
rect 5516 6100 5556 6136
rect 5516 6068 5520 6100
rect 5520 6068 5552 6100
rect 5552 6068 5556 6100
rect 5516 6032 5556 6068
rect 5516 6000 5520 6032
rect 5520 6000 5552 6032
rect 5552 6000 5556 6032
rect 5516 5964 5556 6000
rect 5516 5932 5520 5964
rect 5520 5932 5552 5964
rect 5552 5932 5556 5964
rect 5516 5896 5556 5932
rect 5516 5864 5520 5896
rect 5520 5864 5552 5896
rect 5552 5864 5556 5896
rect 5516 5828 5556 5864
rect 5516 5796 5520 5828
rect 5520 5796 5552 5828
rect 5552 5796 5556 5828
rect 5516 5760 5556 5796
rect 5516 5728 5520 5760
rect 5520 5728 5552 5760
rect 5552 5728 5556 5760
rect 5516 5692 5556 5728
rect 5516 5660 5520 5692
rect 5520 5660 5552 5692
rect 5552 5660 5556 5692
rect 5516 5624 5556 5660
rect 5516 5592 5520 5624
rect 5520 5592 5552 5624
rect 5552 5592 5556 5624
rect 5516 5556 5556 5592
rect 5516 5524 5520 5556
rect 5520 5524 5552 5556
rect 5552 5524 5556 5556
rect 5516 5488 5556 5524
rect 5516 5456 5520 5488
rect 5520 5456 5552 5488
rect 5552 5456 5556 5488
rect 5516 5420 5556 5456
rect 5516 5388 5520 5420
rect 5520 5388 5552 5420
rect 5552 5388 5556 5420
rect 5516 5352 5556 5388
rect 5516 5347 5520 5352
rect 5520 5347 5552 5352
rect 5552 5347 5556 5352
rect 5868 6612 5872 6617
rect 5872 6612 5904 6617
rect 5904 6612 5908 6617
rect 5868 6576 5908 6612
rect 5868 6544 5872 6576
rect 5872 6544 5904 6576
rect 5904 6544 5908 6576
rect 5868 6508 5908 6544
rect 5868 6476 5872 6508
rect 5872 6476 5904 6508
rect 5904 6476 5908 6508
rect 5868 6440 5908 6476
rect 5868 6408 5872 6440
rect 5872 6408 5904 6440
rect 5904 6408 5908 6440
rect 5868 6372 5908 6408
rect 5868 6340 5872 6372
rect 5872 6340 5904 6372
rect 5904 6340 5908 6372
rect 5868 6304 5908 6340
rect 5868 6272 5872 6304
rect 5872 6272 5904 6304
rect 5904 6272 5908 6304
rect 5868 6236 5908 6272
rect 5868 6204 5872 6236
rect 5872 6204 5904 6236
rect 5904 6204 5908 6236
rect 5868 6168 5908 6204
rect 5868 6136 5872 6168
rect 5872 6136 5904 6168
rect 5904 6136 5908 6168
rect 5868 6100 5908 6136
rect 5868 6068 5872 6100
rect 5872 6068 5904 6100
rect 5904 6068 5908 6100
rect 5868 6032 5908 6068
rect 5868 6000 5872 6032
rect 5872 6000 5904 6032
rect 5904 6000 5908 6032
rect 5868 5964 5908 6000
rect 5868 5932 5872 5964
rect 5872 5932 5904 5964
rect 5904 5932 5908 5964
rect 5868 5896 5908 5932
rect 5868 5864 5872 5896
rect 5872 5864 5904 5896
rect 5904 5864 5908 5896
rect 5868 5828 5908 5864
rect 5868 5796 5872 5828
rect 5872 5796 5904 5828
rect 5904 5796 5908 5828
rect 5868 5760 5908 5796
rect 5868 5728 5872 5760
rect 5872 5728 5904 5760
rect 5904 5728 5908 5760
rect 5868 5692 5908 5728
rect 5868 5660 5872 5692
rect 5872 5660 5904 5692
rect 5904 5660 5908 5692
rect 5868 5624 5908 5660
rect 5868 5592 5872 5624
rect 5872 5592 5904 5624
rect 5904 5592 5908 5624
rect 5868 5556 5908 5592
rect 5868 5524 5872 5556
rect 5872 5524 5904 5556
rect 5904 5524 5908 5556
rect 5868 5488 5908 5524
rect 5868 5456 5872 5488
rect 5872 5456 5904 5488
rect 5904 5456 5908 5488
rect 5868 5420 5908 5456
rect 5868 5388 5872 5420
rect 5872 5388 5904 5420
rect 5904 5388 5908 5420
rect 5868 5352 5908 5388
rect 5868 5347 5872 5352
rect 5872 5347 5904 5352
rect 5904 5347 5908 5352
rect 6220 6612 6224 6617
rect 6224 6612 6256 6617
rect 6256 6612 6260 6617
rect 6220 6576 6260 6612
rect 6220 6544 6224 6576
rect 6224 6544 6256 6576
rect 6256 6544 6260 6576
rect 6220 6508 6260 6544
rect 6220 6476 6224 6508
rect 6224 6476 6256 6508
rect 6256 6476 6260 6508
rect 6220 6440 6260 6476
rect 6220 6408 6224 6440
rect 6224 6408 6256 6440
rect 6256 6408 6260 6440
rect 6220 6372 6260 6408
rect 6220 6340 6224 6372
rect 6224 6340 6256 6372
rect 6256 6340 6260 6372
rect 6220 6304 6260 6340
rect 6220 6272 6224 6304
rect 6224 6272 6256 6304
rect 6256 6272 6260 6304
rect 6220 6236 6260 6272
rect 6220 6204 6224 6236
rect 6224 6204 6256 6236
rect 6256 6204 6260 6236
rect 6220 6168 6260 6204
rect 6220 6136 6224 6168
rect 6224 6136 6256 6168
rect 6256 6136 6260 6168
rect 6220 6100 6260 6136
rect 6220 6068 6224 6100
rect 6224 6068 6256 6100
rect 6256 6068 6260 6100
rect 6220 6032 6260 6068
rect 6220 6000 6224 6032
rect 6224 6000 6256 6032
rect 6256 6000 6260 6032
rect 6220 5964 6260 6000
rect 6220 5932 6224 5964
rect 6224 5932 6256 5964
rect 6256 5932 6260 5964
rect 6220 5896 6260 5932
rect 6220 5864 6224 5896
rect 6224 5864 6256 5896
rect 6256 5864 6260 5896
rect 6220 5828 6260 5864
rect 6220 5796 6224 5828
rect 6224 5796 6256 5828
rect 6256 5796 6260 5828
rect 6220 5760 6260 5796
rect 6220 5728 6224 5760
rect 6224 5728 6256 5760
rect 6256 5728 6260 5760
rect 6220 5692 6260 5728
rect 6220 5660 6224 5692
rect 6224 5660 6256 5692
rect 6256 5660 6260 5692
rect 6220 5624 6260 5660
rect 6220 5592 6224 5624
rect 6224 5592 6256 5624
rect 6256 5592 6260 5624
rect 6220 5556 6260 5592
rect 6220 5524 6224 5556
rect 6224 5524 6256 5556
rect 6256 5524 6260 5556
rect 6220 5488 6260 5524
rect 6220 5456 6224 5488
rect 6224 5456 6256 5488
rect 6256 5456 6260 5488
rect 6220 5420 6260 5456
rect 6220 5388 6224 5420
rect 6224 5388 6256 5420
rect 6256 5388 6260 5420
rect 6220 5352 6260 5388
rect 6220 5347 6224 5352
rect 6224 5347 6256 5352
rect 6256 5347 6260 5352
rect 6572 6612 6576 6617
rect 6576 6612 6608 6617
rect 6608 6612 6612 6617
rect 6572 6576 6612 6612
rect 6572 6544 6576 6576
rect 6576 6544 6608 6576
rect 6608 6544 6612 6576
rect 6572 6508 6612 6544
rect 6572 6476 6576 6508
rect 6576 6476 6608 6508
rect 6608 6476 6612 6508
rect 6572 6440 6612 6476
rect 6572 6408 6576 6440
rect 6576 6408 6608 6440
rect 6608 6408 6612 6440
rect 6572 6372 6612 6408
rect 6572 6340 6576 6372
rect 6576 6340 6608 6372
rect 6608 6340 6612 6372
rect 6572 6304 6612 6340
rect 6572 6272 6576 6304
rect 6576 6272 6608 6304
rect 6608 6272 6612 6304
rect 6572 6236 6612 6272
rect 6572 6204 6576 6236
rect 6576 6204 6608 6236
rect 6608 6204 6612 6236
rect 6572 6168 6612 6204
rect 6572 6136 6576 6168
rect 6576 6136 6608 6168
rect 6608 6136 6612 6168
rect 6572 6100 6612 6136
rect 6572 6068 6576 6100
rect 6576 6068 6608 6100
rect 6608 6068 6612 6100
rect 6572 6032 6612 6068
rect 6572 6000 6576 6032
rect 6576 6000 6608 6032
rect 6608 6000 6612 6032
rect 6572 5964 6612 6000
rect 6572 5932 6576 5964
rect 6576 5932 6608 5964
rect 6608 5932 6612 5964
rect 6572 5896 6612 5932
rect 6572 5864 6576 5896
rect 6576 5864 6608 5896
rect 6608 5864 6612 5896
rect 6572 5828 6612 5864
rect 6572 5796 6576 5828
rect 6576 5796 6608 5828
rect 6608 5796 6612 5828
rect 6572 5760 6612 5796
rect 6572 5728 6576 5760
rect 6576 5728 6608 5760
rect 6608 5728 6612 5760
rect 6572 5692 6612 5728
rect 6572 5660 6576 5692
rect 6576 5660 6608 5692
rect 6608 5660 6612 5692
rect 6572 5624 6612 5660
rect 6572 5592 6576 5624
rect 6576 5592 6608 5624
rect 6608 5592 6612 5624
rect 6572 5556 6612 5592
rect 6572 5524 6576 5556
rect 6576 5524 6608 5556
rect 6608 5524 6612 5556
rect 6572 5488 6612 5524
rect 6572 5456 6576 5488
rect 6576 5456 6608 5488
rect 6608 5456 6612 5488
rect 6572 5420 6612 5456
rect 6572 5388 6576 5420
rect 6576 5388 6608 5420
rect 6608 5388 6612 5420
rect 6572 5352 6612 5388
rect 6572 5347 6576 5352
rect 6576 5347 6608 5352
rect 6608 5347 6612 5352
rect 6924 6612 6928 6617
rect 6928 6612 6960 6617
rect 6960 6612 6964 6617
rect 6924 6576 6964 6612
rect 6924 6544 6928 6576
rect 6928 6544 6960 6576
rect 6960 6544 6964 6576
rect 6924 6508 6964 6544
rect 6924 6476 6928 6508
rect 6928 6476 6960 6508
rect 6960 6476 6964 6508
rect 6924 6440 6964 6476
rect 6924 6408 6928 6440
rect 6928 6408 6960 6440
rect 6960 6408 6964 6440
rect 6924 6372 6964 6408
rect 6924 6340 6928 6372
rect 6928 6340 6960 6372
rect 6960 6340 6964 6372
rect 6924 6304 6964 6340
rect 6924 6272 6928 6304
rect 6928 6272 6960 6304
rect 6960 6272 6964 6304
rect 6924 6236 6964 6272
rect 6924 6204 6928 6236
rect 6928 6204 6960 6236
rect 6960 6204 6964 6236
rect 6924 6168 6964 6204
rect 6924 6136 6928 6168
rect 6928 6136 6960 6168
rect 6960 6136 6964 6168
rect 6924 6100 6964 6136
rect 6924 6068 6928 6100
rect 6928 6068 6960 6100
rect 6960 6068 6964 6100
rect 6924 6032 6964 6068
rect 6924 6000 6928 6032
rect 6928 6000 6960 6032
rect 6960 6000 6964 6032
rect 6924 5964 6964 6000
rect 6924 5932 6928 5964
rect 6928 5932 6960 5964
rect 6960 5932 6964 5964
rect 6924 5896 6964 5932
rect 6924 5864 6928 5896
rect 6928 5864 6960 5896
rect 6960 5864 6964 5896
rect 6924 5828 6964 5864
rect 6924 5796 6928 5828
rect 6928 5796 6960 5828
rect 6960 5796 6964 5828
rect 6924 5760 6964 5796
rect 6924 5728 6928 5760
rect 6928 5728 6960 5760
rect 6960 5728 6964 5760
rect 6924 5692 6964 5728
rect 6924 5660 6928 5692
rect 6928 5660 6960 5692
rect 6960 5660 6964 5692
rect 6924 5624 6964 5660
rect 6924 5592 6928 5624
rect 6928 5592 6960 5624
rect 6960 5592 6964 5624
rect 6924 5556 6964 5592
rect 6924 5524 6928 5556
rect 6928 5524 6960 5556
rect 6960 5524 6964 5556
rect 6924 5488 6964 5524
rect 6924 5456 6928 5488
rect 6928 5456 6960 5488
rect 6960 5456 6964 5488
rect 6924 5420 6964 5456
rect 6924 5388 6928 5420
rect 6928 5388 6960 5420
rect 6960 5388 6964 5420
rect 6924 5352 6964 5388
rect 6924 5347 6928 5352
rect 6928 5347 6960 5352
rect 6960 5347 6964 5352
rect 7276 6612 7280 6617
rect 7280 6612 7312 6617
rect 7312 6612 7316 6617
rect 7276 6576 7316 6612
rect 7276 6544 7280 6576
rect 7280 6544 7312 6576
rect 7312 6544 7316 6576
rect 7276 6508 7316 6544
rect 7276 6476 7280 6508
rect 7280 6476 7312 6508
rect 7312 6476 7316 6508
rect 7276 6440 7316 6476
rect 7276 6408 7280 6440
rect 7280 6408 7312 6440
rect 7312 6408 7316 6440
rect 7276 6372 7316 6408
rect 7276 6340 7280 6372
rect 7280 6340 7312 6372
rect 7312 6340 7316 6372
rect 7276 6304 7316 6340
rect 7276 6272 7280 6304
rect 7280 6272 7312 6304
rect 7312 6272 7316 6304
rect 7276 6236 7316 6272
rect 7276 6204 7280 6236
rect 7280 6204 7312 6236
rect 7312 6204 7316 6236
rect 7276 6168 7316 6204
rect 7276 6136 7280 6168
rect 7280 6136 7312 6168
rect 7312 6136 7316 6168
rect 7276 6100 7316 6136
rect 7276 6068 7280 6100
rect 7280 6068 7312 6100
rect 7312 6068 7316 6100
rect 7276 6032 7316 6068
rect 7276 6000 7280 6032
rect 7280 6000 7312 6032
rect 7312 6000 7316 6032
rect 7276 5964 7316 6000
rect 7276 5932 7280 5964
rect 7280 5932 7312 5964
rect 7312 5932 7316 5964
rect 7276 5896 7316 5932
rect 7276 5864 7280 5896
rect 7280 5864 7312 5896
rect 7312 5864 7316 5896
rect 7276 5828 7316 5864
rect 7276 5796 7280 5828
rect 7280 5796 7312 5828
rect 7312 5796 7316 5828
rect 7276 5760 7316 5796
rect 7276 5728 7280 5760
rect 7280 5728 7312 5760
rect 7312 5728 7316 5760
rect 7276 5692 7316 5728
rect 7276 5660 7280 5692
rect 7280 5660 7312 5692
rect 7312 5660 7316 5692
rect 7276 5624 7316 5660
rect 7276 5592 7280 5624
rect 7280 5592 7312 5624
rect 7312 5592 7316 5624
rect 7276 5556 7316 5592
rect 7276 5524 7280 5556
rect 7280 5524 7312 5556
rect 7312 5524 7316 5556
rect 7276 5488 7316 5524
rect 7276 5456 7280 5488
rect 7280 5456 7312 5488
rect 7312 5456 7316 5488
rect 7276 5420 7316 5456
rect 7276 5388 7280 5420
rect 7280 5388 7312 5420
rect 7312 5388 7316 5420
rect 7276 5352 7316 5388
rect 7276 5347 7280 5352
rect 7280 5347 7312 5352
rect 7312 5347 7316 5352
rect 7628 6612 7632 6617
rect 7632 6612 7664 6617
rect 7664 6612 7668 6617
rect 7628 6576 7668 6612
rect 7628 6544 7632 6576
rect 7632 6544 7664 6576
rect 7664 6544 7668 6576
rect 7628 6508 7668 6544
rect 7628 6476 7632 6508
rect 7632 6476 7664 6508
rect 7664 6476 7668 6508
rect 7628 6440 7668 6476
rect 7628 6408 7632 6440
rect 7632 6408 7664 6440
rect 7664 6408 7668 6440
rect 7628 6372 7668 6408
rect 7628 6340 7632 6372
rect 7632 6340 7664 6372
rect 7664 6340 7668 6372
rect 7628 6304 7668 6340
rect 7628 6272 7632 6304
rect 7632 6272 7664 6304
rect 7664 6272 7668 6304
rect 7628 6236 7668 6272
rect 7628 6204 7632 6236
rect 7632 6204 7664 6236
rect 7664 6204 7668 6236
rect 7628 6168 7668 6204
rect 7628 6136 7632 6168
rect 7632 6136 7664 6168
rect 7664 6136 7668 6168
rect 7628 6100 7668 6136
rect 7628 6068 7632 6100
rect 7632 6068 7664 6100
rect 7664 6068 7668 6100
rect 7628 6032 7668 6068
rect 7628 6000 7632 6032
rect 7632 6000 7664 6032
rect 7664 6000 7668 6032
rect 7628 5964 7668 6000
rect 7628 5932 7632 5964
rect 7632 5932 7664 5964
rect 7664 5932 7668 5964
rect 7628 5896 7668 5932
rect 7628 5864 7632 5896
rect 7632 5864 7664 5896
rect 7664 5864 7668 5896
rect 7628 5828 7668 5864
rect 7628 5796 7632 5828
rect 7632 5796 7664 5828
rect 7664 5796 7668 5828
rect 7628 5760 7668 5796
rect 7628 5728 7632 5760
rect 7632 5728 7664 5760
rect 7664 5728 7668 5760
rect 7628 5692 7668 5728
rect 7628 5660 7632 5692
rect 7632 5660 7664 5692
rect 7664 5660 7668 5692
rect 7628 5624 7668 5660
rect 7628 5592 7632 5624
rect 7632 5592 7664 5624
rect 7664 5592 7668 5624
rect 7628 5556 7668 5592
rect 7628 5524 7632 5556
rect 7632 5524 7664 5556
rect 7664 5524 7668 5556
rect 7628 5488 7668 5524
rect 7628 5456 7632 5488
rect 7632 5456 7664 5488
rect 7664 5456 7668 5488
rect 7628 5420 7668 5456
rect 7628 5388 7632 5420
rect 7632 5388 7664 5420
rect 7664 5388 7668 5420
rect 7628 5352 7668 5388
rect 7628 5347 7632 5352
rect 7632 5347 7664 5352
rect 7664 5347 7668 5352
rect 7980 6612 7984 6617
rect 7984 6612 8016 6617
rect 8016 6612 8020 6617
rect 7980 6576 8020 6612
rect 7980 6544 7984 6576
rect 7984 6544 8016 6576
rect 8016 6544 8020 6576
rect 7980 6508 8020 6544
rect 7980 6476 7984 6508
rect 7984 6476 8016 6508
rect 8016 6476 8020 6508
rect 7980 6440 8020 6476
rect 7980 6408 7984 6440
rect 7984 6408 8016 6440
rect 8016 6408 8020 6440
rect 7980 6372 8020 6408
rect 7980 6340 7984 6372
rect 7984 6340 8016 6372
rect 8016 6340 8020 6372
rect 7980 6304 8020 6340
rect 7980 6272 7984 6304
rect 7984 6272 8016 6304
rect 8016 6272 8020 6304
rect 7980 6236 8020 6272
rect 7980 6204 7984 6236
rect 7984 6204 8016 6236
rect 8016 6204 8020 6236
rect 7980 6168 8020 6204
rect 7980 6136 7984 6168
rect 7984 6136 8016 6168
rect 8016 6136 8020 6168
rect 7980 6100 8020 6136
rect 7980 6068 7984 6100
rect 7984 6068 8016 6100
rect 8016 6068 8020 6100
rect 7980 6032 8020 6068
rect 7980 6000 7984 6032
rect 7984 6000 8016 6032
rect 8016 6000 8020 6032
rect 7980 5964 8020 6000
rect 7980 5932 7984 5964
rect 7984 5932 8016 5964
rect 8016 5932 8020 5964
rect 7980 5896 8020 5932
rect 7980 5864 7984 5896
rect 7984 5864 8016 5896
rect 8016 5864 8020 5896
rect 7980 5828 8020 5864
rect 7980 5796 7984 5828
rect 7984 5796 8016 5828
rect 8016 5796 8020 5828
rect 7980 5760 8020 5796
rect 7980 5728 7984 5760
rect 7984 5728 8016 5760
rect 8016 5728 8020 5760
rect 7980 5692 8020 5728
rect 7980 5660 7984 5692
rect 7984 5660 8016 5692
rect 8016 5660 8020 5692
rect 7980 5624 8020 5660
rect 7980 5592 7984 5624
rect 7984 5592 8016 5624
rect 8016 5592 8020 5624
rect 7980 5556 8020 5592
rect 7980 5524 7984 5556
rect 7984 5524 8016 5556
rect 8016 5524 8020 5556
rect 7980 5488 8020 5524
rect 7980 5456 7984 5488
rect 7984 5456 8016 5488
rect 8016 5456 8020 5488
rect 7980 5420 8020 5456
rect 7980 5388 7984 5420
rect 7984 5388 8016 5420
rect 8016 5388 8020 5420
rect 7980 5352 8020 5388
rect 7980 5347 7984 5352
rect 7984 5347 8016 5352
rect 8016 5347 8020 5352
rect 8332 6612 8336 6617
rect 8336 6612 8368 6617
rect 8368 6612 8372 6617
rect 8332 6576 8372 6612
rect 8332 6544 8336 6576
rect 8336 6544 8368 6576
rect 8368 6544 8372 6576
rect 8332 6508 8372 6544
rect 8332 6476 8336 6508
rect 8336 6476 8368 6508
rect 8368 6476 8372 6508
rect 8332 6440 8372 6476
rect 8332 6408 8336 6440
rect 8336 6408 8368 6440
rect 8368 6408 8372 6440
rect 8332 6372 8372 6408
rect 8332 6340 8336 6372
rect 8336 6340 8368 6372
rect 8368 6340 8372 6372
rect 8332 6304 8372 6340
rect 8332 6272 8336 6304
rect 8336 6272 8368 6304
rect 8368 6272 8372 6304
rect 8332 6236 8372 6272
rect 8332 6204 8336 6236
rect 8336 6204 8368 6236
rect 8368 6204 8372 6236
rect 8332 6168 8372 6204
rect 8332 6136 8336 6168
rect 8336 6136 8368 6168
rect 8368 6136 8372 6168
rect 8332 6100 8372 6136
rect 8332 6068 8336 6100
rect 8336 6068 8368 6100
rect 8368 6068 8372 6100
rect 8332 6032 8372 6068
rect 8332 6000 8336 6032
rect 8336 6000 8368 6032
rect 8368 6000 8372 6032
rect 8332 5964 8372 6000
rect 8332 5932 8336 5964
rect 8336 5932 8368 5964
rect 8368 5932 8372 5964
rect 8332 5896 8372 5932
rect 8332 5864 8336 5896
rect 8336 5864 8368 5896
rect 8368 5864 8372 5896
rect 8332 5828 8372 5864
rect 8332 5796 8336 5828
rect 8336 5796 8368 5828
rect 8368 5796 8372 5828
rect 8332 5760 8372 5796
rect 8332 5728 8336 5760
rect 8336 5728 8368 5760
rect 8368 5728 8372 5760
rect 8332 5692 8372 5728
rect 8332 5660 8336 5692
rect 8336 5660 8368 5692
rect 8368 5660 8372 5692
rect 8332 5624 8372 5660
rect 8332 5592 8336 5624
rect 8336 5592 8368 5624
rect 8368 5592 8372 5624
rect 8332 5556 8372 5592
rect 8332 5524 8336 5556
rect 8336 5524 8368 5556
rect 8368 5524 8372 5556
rect 8332 5488 8372 5524
rect 8332 5456 8336 5488
rect 8336 5456 8368 5488
rect 8368 5456 8372 5488
rect 8332 5420 8372 5456
rect 8332 5388 8336 5420
rect 8336 5388 8368 5420
rect 8368 5388 8372 5420
rect 8332 5352 8372 5388
rect 8332 5347 8336 5352
rect 8336 5347 8368 5352
rect 8368 5347 8372 5352
rect 8684 6612 8688 6617
rect 8688 6612 8720 6617
rect 8720 6612 8724 6617
rect 8684 6576 8724 6612
rect 8684 6544 8688 6576
rect 8688 6544 8720 6576
rect 8720 6544 8724 6576
rect 8684 6508 8724 6544
rect 8684 6476 8688 6508
rect 8688 6476 8720 6508
rect 8720 6476 8724 6508
rect 8684 6440 8724 6476
rect 8684 6408 8688 6440
rect 8688 6408 8720 6440
rect 8720 6408 8724 6440
rect 8684 6372 8724 6408
rect 8684 6340 8688 6372
rect 8688 6340 8720 6372
rect 8720 6340 8724 6372
rect 8684 6304 8724 6340
rect 8684 6272 8688 6304
rect 8688 6272 8720 6304
rect 8720 6272 8724 6304
rect 8684 6236 8724 6272
rect 8684 6204 8688 6236
rect 8688 6204 8720 6236
rect 8720 6204 8724 6236
rect 8684 6168 8724 6204
rect 8684 6136 8688 6168
rect 8688 6136 8720 6168
rect 8720 6136 8724 6168
rect 8684 6100 8724 6136
rect 8684 6068 8688 6100
rect 8688 6068 8720 6100
rect 8720 6068 8724 6100
rect 8684 6032 8724 6068
rect 8684 6000 8688 6032
rect 8688 6000 8720 6032
rect 8720 6000 8724 6032
rect 8684 5964 8724 6000
rect 8684 5932 8688 5964
rect 8688 5932 8720 5964
rect 8720 5932 8724 5964
rect 8684 5896 8724 5932
rect 8684 5864 8688 5896
rect 8688 5864 8720 5896
rect 8720 5864 8724 5896
rect 8684 5828 8724 5864
rect 8684 5796 8688 5828
rect 8688 5796 8720 5828
rect 8720 5796 8724 5828
rect 8684 5760 8724 5796
rect 8684 5728 8688 5760
rect 8688 5728 8720 5760
rect 8720 5728 8724 5760
rect 8684 5692 8724 5728
rect 8684 5660 8688 5692
rect 8688 5660 8720 5692
rect 8720 5660 8724 5692
rect 8684 5624 8724 5660
rect 8684 5592 8688 5624
rect 8688 5592 8720 5624
rect 8720 5592 8724 5624
rect 8684 5556 8724 5592
rect 8684 5524 8688 5556
rect 8688 5524 8720 5556
rect 8720 5524 8724 5556
rect 8684 5488 8724 5524
rect 8684 5456 8688 5488
rect 8688 5456 8720 5488
rect 8720 5456 8724 5488
rect 8684 5420 8724 5456
rect 8684 5388 8688 5420
rect 8688 5388 8720 5420
rect 8720 5388 8724 5420
rect 8684 5352 8724 5388
rect 8684 5347 8688 5352
rect 8688 5347 8720 5352
rect 8720 5347 8724 5352
rect 9036 6612 9040 6617
rect 9040 6612 9072 6617
rect 9072 6612 9076 6617
rect 9036 6576 9076 6612
rect 9036 6544 9040 6576
rect 9040 6544 9072 6576
rect 9072 6544 9076 6576
rect 9036 6508 9076 6544
rect 9036 6476 9040 6508
rect 9040 6476 9072 6508
rect 9072 6476 9076 6508
rect 9036 6440 9076 6476
rect 9036 6408 9040 6440
rect 9040 6408 9072 6440
rect 9072 6408 9076 6440
rect 9036 6372 9076 6408
rect 9036 6340 9040 6372
rect 9040 6340 9072 6372
rect 9072 6340 9076 6372
rect 9036 6304 9076 6340
rect 9036 6272 9040 6304
rect 9040 6272 9072 6304
rect 9072 6272 9076 6304
rect 9036 6236 9076 6272
rect 9036 6204 9040 6236
rect 9040 6204 9072 6236
rect 9072 6204 9076 6236
rect 9036 6168 9076 6204
rect 9036 6136 9040 6168
rect 9040 6136 9072 6168
rect 9072 6136 9076 6168
rect 9036 6100 9076 6136
rect 9036 6068 9040 6100
rect 9040 6068 9072 6100
rect 9072 6068 9076 6100
rect 9036 6032 9076 6068
rect 9036 6000 9040 6032
rect 9040 6000 9072 6032
rect 9072 6000 9076 6032
rect 9036 5964 9076 6000
rect 9036 5932 9040 5964
rect 9040 5932 9072 5964
rect 9072 5932 9076 5964
rect 9036 5896 9076 5932
rect 9036 5864 9040 5896
rect 9040 5864 9072 5896
rect 9072 5864 9076 5896
rect 9036 5828 9076 5864
rect 9036 5796 9040 5828
rect 9040 5796 9072 5828
rect 9072 5796 9076 5828
rect 9036 5760 9076 5796
rect 9036 5728 9040 5760
rect 9040 5728 9072 5760
rect 9072 5728 9076 5760
rect 9036 5692 9076 5728
rect 9036 5660 9040 5692
rect 9040 5660 9072 5692
rect 9072 5660 9076 5692
rect 9036 5624 9076 5660
rect 9036 5592 9040 5624
rect 9040 5592 9072 5624
rect 9072 5592 9076 5624
rect 9036 5556 9076 5592
rect 9036 5524 9040 5556
rect 9040 5524 9072 5556
rect 9072 5524 9076 5556
rect 9036 5488 9076 5524
rect 9036 5456 9040 5488
rect 9040 5456 9072 5488
rect 9072 5456 9076 5488
rect 9036 5420 9076 5456
rect 9036 5388 9040 5420
rect 9040 5388 9072 5420
rect 9072 5388 9076 5420
rect 9036 5352 9076 5388
rect 9036 5347 9040 5352
rect 9040 5347 9072 5352
rect 9072 5347 9076 5352
rect 9388 6612 9392 6617
rect 9392 6612 9424 6617
rect 9424 6612 9428 6617
rect 9388 6576 9428 6612
rect 9388 6544 9392 6576
rect 9392 6544 9424 6576
rect 9424 6544 9428 6576
rect 9388 6508 9428 6544
rect 9388 6476 9392 6508
rect 9392 6476 9424 6508
rect 9424 6476 9428 6508
rect 9388 6440 9428 6476
rect 9388 6408 9392 6440
rect 9392 6408 9424 6440
rect 9424 6408 9428 6440
rect 9388 6372 9428 6408
rect 9388 6340 9392 6372
rect 9392 6340 9424 6372
rect 9424 6340 9428 6372
rect 9388 6304 9428 6340
rect 9388 6272 9392 6304
rect 9392 6272 9424 6304
rect 9424 6272 9428 6304
rect 9388 6236 9428 6272
rect 9388 6204 9392 6236
rect 9392 6204 9424 6236
rect 9424 6204 9428 6236
rect 9388 6168 9428 6204
rect 9388 6136 9392 6168
rect 9392 6136 9424 6168
rect 9424 6136 9428 6168
rect 9388 6100 9428 6136
rect 9388 6068 9392 6100
rect 9392 6068 9424 6100
rect 9424 6068 9428 6100
rect 9388 6032 9428 6068
rect 9388 6000 9392 6032
rect 9392 6000 9424 6032
rect 9424 6000 9428 6032
rect 9388 5964 9428 6000
rect 9388 5932 9392 5964
rect 9392 5932 9424 5964
rect 9424 5932 9428 5964
rect 9388 5896 9428 5932
rect 9388 5864 9392 5896
rect 9392 5864 9424 5896
rect 9424 5864 9428 5896
rect 9388 5828 9428 5864
rect 9388 5796 9392 5828
rect 9392 5796 9424 5828
rect 9424 5796 9428 5828
rect 9388 5760 9428 5796
rect 9388 5728 9392 5760
rect 9392 5728 9424 5760
rect 9424 5728 9428 5760
rect 9388 5692 9428 5728
rect 9388 5660 9392 5692
rect 9392 5660 9424 5692
rect 9424 5660 9428 5692
rect 9388 5624 9428 5660
rect 9388 5592 9392 5624
rect 9392 5592 9424 5624
rect 9424 5592 9428 5624
rect 9388 5556 9428 5592
rect 9388 5524 9392 5556
rect 9392 5524 9424 5556
rect 9424 5524 9428 5556
rect 9388 5488 9428 5524
rect 9388 5456 9392 5488
rect 9392 5456 9424 5488
rect 9424 5456 9428 5488
rect 9388 5420 9428 5456
rect 9388 5388 9392 5420
rect 9392 5388 9424 5420
rect 9424 5388 9428 5420
rect 9388 5352 9428 5388
rect 9388 5347 9392 5352
rect 9392 5347 9424 5352
rect 9424 5347 9428 5352
rect 9740 6612 9744 6617
rect 9744 6612 9776 6617
rect 9776 6612 9780 6617
rect 9740 6576 9780 6612
rect 9740 6544 9744 6576
rect 9744 6544 9776 6576
rect 9776 6544 9780 6576
rect 9740 6508 9780 6544
rect 9740 6476 9744 6508
rect 9744 6476 9776 6508
rect 9776 6476 9780 6508
rect 9740 6440 9780 6476
rect 9740 6408 9744 6440
rect 9744 6408 9776 6440
rect 9776 6408 9780 6440
rect 9740 6372 9780 6408
rect 9740 6340 9744 6372
rect 9744 6340 9776 6372
rect 9776 6340 9780 6372
rect 9740 6304 9780 6340
rect 9740 6272 9744 6304
rect 9744 6272 9776 6304
rect 9776 6272 9780 6304
rect 9740 6236 9780 6272
rect 9740 6204 9744 6236
rect 9744 6204 9776 6236
rect 9776 6204 9780 6236
rect 9740 6168 9780 6204
rect 9740 6136 9744 6168
rect 9744 6136 9776 6168
rect 9776 6136 9780 6168
rect 9740 6100 9780 6136
rect 9740 6068 9744 6100
rect 9744 6068 9776 6100
rect 9776 6068 9780 6100
rect 9740 6032 9780 6068
rect 9740 6000 9744 6032
rect 9744 6000 9776 6032
rect 9776 6000 9780 6032
rect 9740 5964 9780 6000
rect 9740 5932 9744 5964
rect 9744 5932 9776 5964
rect 9776 5932 9780 5964
rect 9740 5896 9780 5932
rect 9740 5864 9744 5896
rect 9744 5864 9776 5896
rect 9776 5864 9780 5896
rect 9740 5828 9780 5864
rect 9740 5796 9744 5828
rect 9744 5796 9776 5828
rect 9776 5796 9780 5828
rect 9740 5760 9780 5796
rect 9740 5728 9744 5760
rect 9744 5728 9776 5760
rect 9776 5728 9780 5760
rect 9740 5692 9780 5728
rect 9740 5660 9744 5692
rect 9744 5660 9776 5692
rect 9776 5660 9780 5692
rect 9740 5624 9780 5660
rect 9740 5592 9744 5624
rect 9744 5592 9776 5624
rect 9776 5592 9780 5624
rect 9740 5556 9780 5592
rect 9740 5524 9744 5556
rect 9744 5524 9776 5556
rect 9776 5524 9780 5556
rect 9740 5488 9780 5524
rect 9740 5456 9744 5488
rect 9744 5456 9776 5488
rect 9776 5456 9780 5488
rect 9740 5420 9780 5456
rect 9740 5388 9744 5420
rect 9744 5388 9776 5420
rect 9776 5388 9780 5420
rect 9740 5352 9780 5388
rect 9740 5347 9744 5352
rect 9744 5347 9776 5352
rect 9776 5347 9780 5352
rect 10092 6612 10096 6617
rect 10096 6612 10128 6617
rect 10128 6612 10132 6617
rect 10092 6576 10132 6612
rect 10092 6544 10096 6576
rect 10096 6544 10128 6576
rect 10128 6544 10132 6576
rect 10092 6508 10132 6544
rect 10092 6476 10096 6508
rect 10096 6476 10128 6508
rect 10128 6476 10132 6508
rect 10092 6440 10132 6476
rect 10092 6408 10096 6440
rect 10096 6408 10128 6440
rect 10128 6408 10132 6440
rect 10092 6372 10132 6408
rect 10092 6340 10096 6372
rect 10096 6340 10128 6372
rect 10128 6340 10132 6372
rect 10092 6304 10132 6340
rect 10092 6272 10096 6304
rect 10096 6272 10128 6304
rect 10128 6272 10132 6304
rect 10092 6236 10132 6272
rect 10092 6204 10096 6236
rect 10096 6204 10128 6236
rect 10128 6204 10132 6236
rect 10092 6168 10132 6204
rect 10092 6136 10096 6168
rect 10096 6136 10128 6168
rect 10128 6136 10132 6168
rect 10092 6100 10132 6136
rect 10092 6068 10096 6100
rect 10096 6068 10128 6100
rect 10128 6068 10132 6100
rect 10092 6032 10132 6068
rect 10092 6000 10096 6032
rect 10096 6000 10128 6032
rect 10128 6000 10132 6032
rect 10092 5964 10132 6000
rect 10092 5932 10096 5964
rect 10096 5932 10128 5964
rect 10128 5932 10132 5964
rect 10092 5896 10132 5932
rect 10092 5864 10096 5896
rect 10096 5864 10128 5896
rect 10128 5864 10132 5896
rect 10092 5828 10132 5864
rect 10092 5796 10096 5828
rect 10096 5796 10128 5828
rect 10128 5796 10132 5828
rect 10092 5760 10132 5796
rect 10092 5728 10096 5760
rect 10096 5728 10128 5760
rect 10128 5728 10132 5760
rect 10092 5692 10132 5728
rect 10092 5660 10096 5692
rect 10096 5660 10128 5692
rect 10128 5660 10132 5692
rect 10092 5624 10132 5660
rect 10092 5592 10096 5624
rect 10096 5592 10128 5624
rect 10128 5592 10132 5624
rect 10092 5556 10132 5592
rect 10092 5524 10096 5556
rect 10096 5524 10128 5556
rect 10128 5524 10132 5556
rect 10092 5488 10132 5524
rect 10092 5456 10096 5488
rect 10096 5456 10128 5488
rect 10128 5456 10132 5488
rect 10092 5420 10132 5456
rect 10092 5388 10096 5420
rect 10096 5388 10128 5420
rect 10128 5388 10132 5420
rect 10092 5352 10132 5388
rect 10092 5347 10096 5352
rect 10096 5347 10128 5352
rect 10128 5347 10132 5352
rect 10444 6612 10448 6617
rect 10448 6612 10480 6617
rect 10480 6612 10484 6617
rect 10444 6576 10484 6612
rect 10444 6544 10448 6576
rect 10448 6544 10480 6576
rect 10480 6544 10484 6576
rect 10444 6508 10484 6544
rect 10444 6476 10448 6508
rect 10448 6476 10480 6508
rect 10480 6476 10484 6508
rect 10444 6440 10484 6476
rect 10444 6408 10448 6440
rect 10448 6408 10480 6440
rect 10480 6408 10484 6440
rect 10444 6372 10484 6408
rect 10444 6340 10448 6372
rect 10448 6340 10480 6372
rect 10480 6340 10484 6372
rect 10444 6304 10484 6340
rect 10444 6272 10448 6304
rect 10448 6272 10480 6304
rect 10480 6272 10484 6304
rect 10444 6236 10484 6272
rect 10444 6204 10448 6236
rect 10448 6204 10480 6236
rect 10480 6204 10484 6236
rect 10444 6168 10484 6204
rect 10444 6136 10448 6168
rect 10448 6136 10480 6168
rect 10480 6136 10484 6168
rect 10444 6100 10484 6136
rect 10444 6068 10448 6100
rect 10448 6068 10480 6100
rect 10480 6068 10484 6100
rect 10444 6032 10484 6068
rect 10444 6000 10448 6032
rect 10448 6000 10480 6032
rect 10480 6000 10484 6032
rect 10444 5964 10484 6000
rect 10444 5932 10448 5964
rect 10448 5932 10480 5964
rect 10480 5932 10484 5964
rect 10444 5896 10484 5932
rect 10444 5864 10448 5896
rect 10448 5864 10480 5896
rect 10480 5864 10484 5896
rect 10444 5828 10484 5864
rect 10444 5796 10448 5828
rect 10448 5796 10480 5828
rect 10480 5796 10484 5828
rect 10444 5760 10484 5796
rect 10444 5728 10448 5760
rect 10448 5728 10480 5760
rect 10480 5728 10484 5760
rect 10444 5692 10484 5728
rect 10444 5660 10448 5692
rect 10448 5660 10480 5692
rect 10480 5660 10484 5692
rect 10444 5624 10484 5660
rect 10444 5592 10448 5624
rect 10448 5592 10480 5624
rect 10480 5592 10484 5624
rect 10444 5556 10484 5592
rect 10444 5524 10448 5556
rect 10448 5524 10480 5556
rect 10480 5524 10484 5556
rect 10444 5488 10484 5524
rect 10444 5456 10448 5488
rect 10448 5456 10480 5488
rect 10480 5456 10484 5488
rect 10444 5420 10484 5456
rect 10444 5388 10448 5420
rect 10448 5388 10480 5420
rect 10480 5388 10484 5420
rect 10444 5352 10484 5388
rect 10444 5347 10448 5352
rect 10448 5347 10480 5352
rect 10480 5347 10484 5352
rect 10796 6612 10800 6617
rect 10800 6612 10832 6617
rect 10832 6612 10836 6617
rect 10796 6576 10836 6612
rect 10796 6544 10800 6576
rect 10800 6544 10832 6576
rect 10832 6544 10836 6576
rect 10796 6508 10836 6544
rect 10796 6476 10800 6508
rect 10800 6476 10832 6508
rect 10832 6476 10836 6508
rect 10796 6440 10836 6476
rect 10796 6408 10800 6440
rect 10800 6408 10832 6440
rect 10832 6408 10836 6440
rect 10796 6372 10836 6408
rect 10796 6340 10800 6372
rect 10800 6340 10832 6372
rect 10832 6340 10836 6372
rect 10796 6304 10836 6340
rect 10796 6272 10800 6304
rect 10800 6272 10832 6304
rect 10832 6272 10836 6304
rect 10796 6236 10836 6272
rect 10796 6204 10800 6236
rect 10800 6204 10832 6236
rect 10832 6204 10836 6236
rect 10796 6168 10836 6204
rect 10796 6136 10800 6168
rect 10800 6136 10832 6168
rect 10832 6136 10836 6168
rect 10796 6100 10836 6136
rect 10796 6068 10800 6100
rect 10800 6068 10832 6100
rect 10832 6068 10836 6100
rect 10796 6032 10836 6068
rect 10796 6000 10800 6032
rect 10800 6000 10832 6032
rect 10832 6000 10836 6032
rect 10796 5964 10836 6000
rect 10796 5932 10800 5964
rect 10800 5932 10832 5964
rect 10832 5932 10836 5964
rect 10796 5896 10836 5932
rect 10796 5864 10800 5896
rect 10800 5864 10832 5896
rect 10832 5864 10836 5896
rect 10796 5828 10836 5864
rect 10796 5796 10800 5828
rect 10800 5796 10832 5828
rect 10832 5796 10836 5828
rect 10796 5760 10836 5796
rect 10796 5728 10800 5760
rect 10800 5728 10832 5760
rect 10832 5728 10836 5760
rect 10796 5692 10836 5728
rect 10796 5660 10800 5692
rect 10800 5660 10832 5692
rect 10832 5660 10836 5692
rect 10796 5624 10836 5660
rect 10796 5592 10800 5624
rect 10800 5592 10832 5624
rect 10832 5592 10836 5624
rect 10796 5556 10836 5592
rect 10796 5524 10800 5556
rect 10800 5524 10832 5556
rect 10832 5524 10836 5556
rect 10796 5488 10836 5524
rect 10796 5456 10800 5488
rect 10800 5456 10832 5488
rect 10832 5456 10836 5488
rect 10796 5420 10836 5456
rect 10796 5388 10800 5420
rect 10800 5388 10832 5420
rect 10832 5388 10836 5420
rect 10796 5352 10836 5388
rect 10796 5347 10800 5352
rect 10800 5347 10832 5352
rect 10832 5347 10836 5352
rect 11148 6612 11152 6617
rect 11152 6612 11184 6617
rect 11184 6612 11188 6617
rect 11148 6576 11188 6612
rect 11148 6544 11152 6576
rect 11152 6544 11184 6576
rect 11184 6544 11188 6576
rect 11148 6508 11188 6544
rect 11148 6476 11152 6508
rect 11152 6476 11184 6508
rect 11184 6476 11188 6508
rect 11148 6440 11188 6476
rect 11148 6408 11152 6440
rect 11152 6408 11184 6440
rect 11184 6408 11188 6440
rect 11148 6372 11188 6408
rect 11148 6340 11152 6372
rect 11152 6340 11184 6372
rect 11184 6340 11188 6372
rect 11148 6304 11188 6340
rect 11148 6272 11152 6304
rect 11152 6272 11184 6304
rect 11184 6272 11188 6304
rect 11148 6236 11188 6272
rect 11148 6204 11152 6236
rect 11152 6204 11184 6236
rect 11184 6204 11188 6236
rect 11148 6168 11188 6204
rect 11148 6136 11152 6168
rect 11152 6136 11184 6168
rect 11184 6136 11188 6168
rect 11148 6100 11188 6136
rect 11148 6068 11152 6100
rect 11152 6068 11184 6100
rect 11184 6068 11188 6100
rect 11148 6032 11188 6068
rect 11148 6000 11152 6032
rect 11152 6000 11184 6032
rect 11184 6000 11188 6032
rect 11148 5964 11188 6000
rect 11148 5932 11152 5964
rect 11152 5932 11184 5964
rect 11184 5932 11188 5964
rect 11148 5896 11188 5932
rect 11148 5864 11152 5896
rect 11152 5864 11184 5896
rect 11184 5864 11188 5896
rect 11148 5828 11188 5864
rect 11148 5796 11152 5828
rect 11152 5796 11184 5828
rect 11184 5796 11188 5828
rect 11148 5760 11188 5796
rect 11148 5728 11152 5760
rect 11152 5728 11184 5760
rect 11184 5728 11188 5760
rect 11148 5692 11188 5728
rect 11148 5660 11152 5692
rect 11152 5660 11184 5692
rect 11184 5660 11188 5692
rect 11148 5624 11188 5660
rect 11148 5592 11152 5624
rect 11152 5592 11184 5624
rect 11184 5592 11188 5624
rect 11148 5556 11188 5592
rect 11148 5524 11152 5556
rect 11152 5524 11184 5556
rect 11184 5524 11188 5556
rect 11148 5488 11188 5524
rect 11148 5456 11152 5488
rect 11152 5456 11184 5488
rect 11184 5456 11188 5488
rect 11148 5420 11188 5456
rect 11148 5388 11152 5420
rect 11152 5388 11184 5420
rect 11184 5388 11188 5420
rect 11148 5352 11188 5388
rect 11148 5347 11152 5352
rect 11152 5347 11184 5352
rect 11184 5347 11188 5352
rect 11500 6612 11504 6617
rect 11504 6612 11536 6617
rect 11536 6612 11540 6617
rect 11500 6576 11540 6612
rect 11500 6544 11504 6576
rect 11504 6544 11536 6576
rect 11536 6544 11540 6576
rect 11500 6508 11540 6544
rect 11500 6476 11504 6508
rect 11504 6476 11536 6508
rect 11536 6476 11540 6508
rect 11500 6440 11540 6476
rect 11500 6408 11504 6440
rect 11504 6408 11536 6440
rect 11536 6408 11540 6440
rect 11500 6372 11540 6408
rect 11500 6340 11504 6372
rect 11504 6340 11536 6372
rect 11536 6340 11540 6372
rect 11500 6304 11540 6340
rect 11500 6272 11504 6304
rect 11504 6272 11536 6304
rect 11536 6272 11540 6304
rect 11500 6236 11540 6272
rect 11500 6204 11504 6236
rect 11504 6204 11536 6236
rect 11536 6204 11540 6236
rect 11500 6168 11540 6204
rect 11500 6136 11504 6168
rect 11504 6136 11536 6168
rect 11536 6136 11540 6168
rect 11500 6100 11540 6136
rect 11500 6068 11504 6100
rect 11504 6068 11536 6100
rect 11536 6068 11540 6100
rect 11500 6032 11540 6068
rect 11500 6000 11504 6032
rect 11504 6000 11536 6032
rect 11536 6000 11540 6032
rect 11500 5964 11540 6000
rect 11500 5932 11504 5964
rect 11504 5932 11536 5964
rect 11536 5932 11540 5964
rect 11500 5896 11540 5932
rect 11500 5864 11504 5896
rect 11504 5864 11536 5896
rect 11536 5864 11540 5896
rect 11500 5828 11540 5864
rect 11500 5796 11504 5828
rect 11504 5796 11536 5828
rect 11536 5796 11540 5828
rect 11500 5760 11540 5796
rect 11500 5728 11504 5760
rect 11504 5728 11536 5760
rect 11536 5728 11540 5760
rect 11500 5692 11540 5728
rect 11500 5660 11504 5692
rect 11504 5660 11536 5692
rect 11536 5660 11540 5692
rect 11500 5624 11540 5660
rect 11500 5592 11504 5624
rect 11504 5592 11536 5624
rect 11536 5592 11540 5624
rect 11500 5556 11540 5592
rect 11500 5524 11504 5556
rect 11504 5524 11536 5556
rect 11536 5524 11540 5556
rect 11500 5488 11540 5524
rect 11500 5456 11504 5488
rect 11504 5456 11536 5488
rect 11536 5456 11540 5488
rect 11500 5420 11540 5456
rect 11500 5388 11504 5420
rect 11504 5388 11536 5420
rect 11536 5388 11540 5420
rect 11500 5352 11540 5388
rect 11500 5347 11504 5352
rect 11504 5347 11536 5352
rect 11536 5347 11540 5352
rect 11852 6612 11856 6617
rect 11856 6612 11888 6617
rect 11888 6612 11892 6617
rect 11852 6576 11892 6612
rect 11852 6544 11856 6576
rect 11856 6544 11888 6576
rect 11888 6544 11892 6576
rect 11852 6508 11892 6544
rect 11852 6476 11856 6508
rect 11856 6476 11888 6508
rect 11888 6476 11892 6508
rect 11852 6440 11892 6476
rect 11852 6408 11856 6440
rect 11856 6408 11888 6440
rect 11888 6408 11892 6440
rect 11852 6372 11892 6408
rect 11852 6340 11856 6372
rect 11856 6340 11888 6372
rect 11888 6340 11892 6372
rect 11852 6304 11892 6340
rect 11852 6272 11856 6304
rect 11856 6272 11888 6304
rect 11888 6272 11892 6304
rect 11852 6236 11892 6272
rect 11852 6204 11856 6236
rect 11856 6204 11888 6236
rect 11888 6204 11892 6236
rect 11852 6168 11892 6204
rect 11852 6136 11856 6168
rect 11856 6136 11888 6168
rect 11888 6136 11892 6168
rect 11852 6100 11892 6136
rect 11852 6068 11856 6100
rect 11856 6068 11888 6100
rect 11888 6068 11892 6100
rect 11852 6032 11892 6068
rect 11852 6000 11856 6032
rect 11856 6000 11888 6032
rect 11888 6000 11892 6032
rect 11852 5964 11892 6000
rect 11852 5932 11856 5964
rect 11856 5932 11888 5964
rect 11888 5932 11892 5964
rect 11852 5896 11892 5932
rect 11852 5864 11856 5896
rect 11856 5864 11888 5896
rect 11888 5864 11892 5896
rect 11852 5828 11892 5864
rect 11852 5796 11856 5828
rect 11856 5796 11888 5828
rect 11888 5796 11892 5828
rect 11852 5760 11892 5796
rect 11852 5728 11856 5760
rect 11856 5728 11888 5760
rect 11888 5728 11892 5760
rect 11852 5692 11892 5728
rect 11852 5660 11856 5692
rect 11856 5660 11888 5692
rect 11888 5660 11892 5692
rect 11852 5624 11892 5660
rect 11852 5592 11856 5624
rect 11856 5592 11888 5624
rect 11888 5592 11892 5624
rect 11852 5556 11892 5592
rect 11852 5524 11856 5556
rect 11856 5524 11888 5556
rect 11888 5524 11892 5556
rect 11852 5488 11892 5524
rect 11852 5456 11856 5488
rect 11856 5456 11888 5488
rect 11888 5456 11892 5488
rect 11852 5420 11892 5456
rect 11852 5388 11856 5420
rect 11856 5388 11888 5420
rect 11888 5388 11892 5420
rect 11852 5352 11892 5388
rect 11852 5347 11856 5352
rect 11856 5347 11888 5352
rect 11888 5347 11892 5352
rect 12204 6612 12208 6617
rect 12208 6612 12240 6617
rect 12240 6612 12244 6617
rect 12204 6576 12244 6612
rect 12204 6544 12208 6576
rect 12208 6544 12240 6576
rect 12240 6544 12244 6576
rect 12204 6508 12244 6544
rect 12204 6476 12208 6508
rect 12208 6476 12240 6508
rect 12240 6476 12244 6508
rect 12204 6440 12244 6476
rect 12204 6408 12208 6440
rect 12208 6408 12240 6440
rect 12240 6408 12244 6440
rect 12204 6372 12244 6408
rect 12204 6340 12208 6372
rect 12208 6340 12240 6372
rect 12240 6340 12244 6372
rect 12204 6304 12244 6340
rect 12204 6272 12208 6304
rect 12208 6272 12240 6304
rect 12240 6272 12244 6304
rect 12204 6236 12244 6272
rect 12204 6204 12208 6236
rect 12208 6204 12240 6236
rect 12240 6204 12244 6236
rect 12204 6168 12244 6204
rect 12204 6136 12208 6168
rect 12208 6136 12240 6168
rect 12240 6136 12244 6168
rect 12204 6100 12244 6136
rect 12204 6068 12208 6100
rect 12208 6068 12240 6100
rect 12240 6068 12244 6100
rect 12204 6032 12244 6068
rect 12204 6000 12208 6032
rect 12208 6000 12240 6032
rect 12240 6000 12244 6032
rect 12204 5964 12244 6000
rect 12204 5932 12208 5964
rect 12208 5932 12240 5964
rect 12240 5932 12244 5964
rect 12204 5896 12244 5932
rect 12204 5864 12208 5896
rect 12208 5864 12240 5896
rect 12240 5864 12244 5896
rect 12204 5828 12244 5864
rect 12204 5796 12208 5828
rect 12208 5796 12240 5828
rect 12240 5796 12244 5828
rect 12204 5760 12244 5796
rect 12204 5728 12208 5760
rect 12208 5728 12240 5760
rect 12240 5728 12244 5760
rect 12204 5692 12244 5728
rect 12204 5660 12208 5692
rect 12208 5660 12240 5692
rect 12240 5660 12244 5692
rect 12204 5624 12244 5660
rect 12204 5592 12208 5624
rect 12208 5592 12240 5624
rect 12240 5592 12244 5624
rect 12204 5556 12244 5592
rect 12204 5524 12208 5556
rect 12208 5524 12240 5556
rect 12240 5524 12244 5556
rect 12204 5488 12244 5524
rect 12204 5456 12208 5488
rect 12208 5456 12240 5488
rect 12240 5456 12244 5488
rect 12204 5420 12244 5456
rect 12204 5388 12208 5420
rect 12208 5388 12240 5420
rect 12240 5388 12244 5420
rect 12204 5352 12244 5388
rect 12204 5347 12208 5352
rect 12208 5347 12240 5352
rect 12240 5347 12244 5352
rect 14544 3992 14548 3998
rect 14548 3992 14580 3998
rect 14580 3992 14584 3998
rect 14544 3956 14584 3992
rect 14544 3924 14548 3956
rect 14548 3924 14580 3956
rect 14580 3924 14584 3956
rect 14544 3888 14584 3924
rect 14544 3856 14548 3888
rect 14548 3856 14580 3888
rect 14580 3856 14584 3888
rect 14544 3820 14584 3856
rect 14544 3788 14548 3820
rect 14548 3788 14580 3820
rect 14580 3788 14584 3820
rect 14544 3752 14584 3788
rect 14544 3720 14548 3752
rect 14548 3720 14580 3752
rect 14580 3720 14584 3752
rect 14544 3684 14584 3720
rect 14544 3652 14548 3684
rect 14548 3652 14580 3684
rect 14580 3652 14584 3684
rect 14544 3616 14584 3652
rect 14544 3584 14548 3616
rect 14548 3584 14580 3616
rect 14580 3584 14584 3616
rect 14544 3548 14584 3584
rect 14544 3516 14548 3548
rect 14548 3516 14580 3548
rect 14580 3516 14584 3548
rect 14544 3480 14584 3516
rect 14544 3448 14548 3480
rect 14548 3448 14580 3480
rect 14580 3448 14584 3480
rect 14544 3412 14584 3448
rect 14544 3380 14548 3412
rect 14548 3380 14580 3412
rect 14580 3380 14584 3412
rect 14544 3344 14584 3380
rect 14544 3312 14548 3344
rect 14548 3312 14580 3344
rect 14580 3312 14584 3344
rect 14544 3276 14584 3312
rect 14544 3244 14548 3276
rect 14548 3244 14580 3276
rect 14580 3244 14584 3276
rect 14544 3208 14584 3244
rect 14544 3176 14548 3208
rect 14548 3176 14580 3208
rect 14580 3176 14584 3208
rect 14544 3140 14584 3176
rect 14544 3108 14548 3140
rect 14548 3108 14580 3140
rect 14580 3108 14584 3140
rect 14544 3072 14584 3108
rect 14544 3040 14548 3072
rect 14548 3040 14580 3072
rect 14580 3040 14584 3072
rect 14544 3004 14584 3040
rect 14544 2972 14548 3004
rect 14548 2972 14580 3004
rect 14580 2972 14584 3004
rect 14544 2936 14584 2972
rect 14544 2904 14548 2936
rect 14548 2904 14580 2936
rect 14580 2904 14584 2936
rect 14544 2868 14584 2904
rect 14544 2836 14548 2868
rect 14548 2836 14580 2868
rect 14580 2836 14584 2868
rect 14544 2800 14584 2836
rect 14544 2768 14548 2800
rect 14548 2768 14580 2800
rect 14580 2768 14584 2800
rect 14544 2732 14584 2768
rect 14544 2700 14548 2732
rect 14548 2700 14580 2732
rect 14580 2700 14584 2732
rect 14544 2664 14584 2700
rect 14544 2632 14548 2664
rect 14548 2632 14580 2664
rect 14580 2632 14584 2664
rect 14544 2596 14584 2632
rect 14544 2564 14548 2596
rect 14548 2564 14580 2596
rect 14580 2564 14584 2596
rect 14544 2528 14584 2564
rect 14544 2496 14548 2528
rect 14548 2496 14580 2528
rect 14580 2496 14584 2528
rect 14544 2460 14584 2496
rect 14544 2428 14548 2460
rect 14548 2428 14580 2460
rect 14580 2428 14584 2460
rect 14544 2392 14584 2428
rect 14544 2360 14548 2392
rect 14548 2360 14580 2392
rect 14580 2360 14584 2392
rect 14544 2324 14584 2360
rect 14544 2318 14548 2324
rect 14548 2318 14580 2324
rect 14580 2318 14584 2324
rect 14544 2142 14548 2148
rect 14548 2142 14580 2148
rect 14580 2142 14584 2148
rect 14544 2106 14584 2142
rect 14544 2074 14548 2106
rect 14548 2074 14580 2106
rect 14580 2074 14584 2106
rect 14544 2038 14584 2074
rect 14544 2006 14548 2038
rect 14548 2006 14580 2038
rect 14580 2006 14584 2038
rect 14544 1970 14584 2006
rect 14544 1938 14548 1970
rect 14548 1938 14580 1970
rect 14580 1938 14584 1970
rect 14544 1902 14584 1938
rect 14544 1870 14548 1902
rect 14548 1870 14580 1902
rect 14580 1870 14584 1902
rect 14544 1834 14584 1870
rect 14544 1802 14548 1834
rect 14548 1802 14580 1834
rect 14580 1802 14584 1834
rect 14544 1766 14584 1802
rect 14544 1734 14548 1766
rect 14548 1734 14580 1766
rect 14580 1734 14584 1766
rect 14544 1698 14584 1734
rect 14544 1666 14548 1698
rect 14548 1666 14580 1698
rect 14580 1666 14584 1698
rect 14544 1630 14584 1666
rect 14544 1598 14548 1630
rect 14548 1598 14580 1630
rect 14580 1598 14584 1630
rect 14544 1562 14584 1598
rect 14544 1530 14548 1562
rect 14548 1530 14580 1562
rect 14580 1530 14584 1562
rect 14544 1494 14584 1530
rect 14544 1462 14548 1494
rect 14548 1462 14580 1494
rect 14580 1462 14584 1494
rect 14544 1426 14584 1462
rect 14544 1394 14548 1426
rect 14548 1394 14580 1426
rect 14580 1394 14584 1426
rect 14544 1358 14584 1394
rect 14544 1326 14548 1358
rect 14548 1326 14580 1358
rect 14580 1326 14584 1358
rect 14544 1290 14584 1326
rect 14544 1258 14548 1290
rect 14548 1258 14580 1290
rect 14580 1258 14584 1290
rect 14544 1222 14584 1258
rect 14544 1190 14548 1222
rect 14548 1190 14580 1222
rect 14580 1190 14584 1222
rect 14544 1154 14584 1190
rect 14544 1122 14548 1154
rect 14548 1122 14580 1154
rect 14580 1122 14584 1154
rect 14544 1086 14584 1122
rect 14544 1054 14548 1086
rect 14548 1054 14580 1086
rect 14580 1054 14584 1086
rect 14544 1018 14584 1054
rect 14544 986 14548 1018
rect 14548 986 14580 1018
rect 14580 986 14584 1018
rect 14544 950 14584 986
rect 14544 918 14548 950
rect 14548 918 14580 950
rect 14580 918 14584 950
rect 14544 882 14584 918
rect 14544 850 14548 882
rect 14548 850 14580 882
rect 14580 850 14584 882
rect 14544 814 14584 850
rect 14544 782 14548 814
rect 14548 782 14580 814
rect 14580 782 14584 814
rect 14544 746 14584 782
rect 14544 714 14548 746
rect 14548 714 14580 746
rect 14580 714 14584 746
rect 14544 678 14584 714
rect 14544 646 14548 678
rect 14548 646 14580 678
rect 14580 646 14584 678
rect 14544 610 14584 646
rect 14544 578 14548 610
rect 14548 578 14580 610
rect 14580 578 14584 610
rect 14544 542 14584 578
rect 14544 510 14548 542
rect 14548 510 14580 542
rect 14580 510 14584 542
rect 14544 474 14584 510
rect 14544 468 14548 474
rect 14548 468 14580 474
rect 14580 468 14584 474
rect 14896 3992 14900 3998
rect 14900 3992 14932 3998
rect 14932 3992 14936 3998
rect 14896 3956 14936 3992
rect 14896 3924 14900 3956
rect 14900 3924 14932 3956
rect 14932 3924 14936 3956
rect 14896 3888 14936 3924
rect 14896 3856 14900 3888
rect 14900 3856 14932 3888
rect 14932 3856 14936 3888
rect 14896 3820 14936 3856
rect 14896 3788 14900 3820
rect 14900 3788 14932 3820
rect 14932 3788 14936 3820
rect 14896 3752 14936 3788
rect 14896 3720 14900 3752
rect 14900 3720 14932 3752
rect 14932 3720 14936 3752
rect 14896 3684 14936 3720
rect 14896 3652 14900 3684
rect 14900 3652 14932 3684
rect 14932 3652 14936 3684
rect 14896 3616 14936 3652
rect 14896 3584 14900 3616
rect 14900 3584 14932 3616
rect 14932 3584 14936 3616
rect 14896 3548 14936 3584
rect 14896 3516 14900 3548
rect 14900 3516 14932 3548
rect 14932 3516 14936 3548
rect 14896 3480 14936 3516
rect 14896 3448 14900 3480
rect 14900 3448 14932 3480
rect 14932 3448 14936 3480
rect 14896 3412 14936 3448
rect 14896 3380 14900 3412
rect 14900 3380 14932 3412
rect 14932 3380 14936 3412
rect 14896 3344 14936 3380
rect 14896 3312 14900 3344
rect 14900 3312 14932 3344
rect 14932 3312 14936 3344
rect 14896 3276 14936 3312
rect 14896 3244 14900 3276
rect 14900 3244 14932 3276
rect 14932 3244 14936 3276
rect 14896 3208 14936 3244
rect 14896 3176 14900 3208
rect 14900 3176 14932 3208
rect 14932 3176 14936 3208
rect 14896 3140 14936 3176
rect 14896 3108 14900 3140
rect 14900 3108 14932 3140
rect 14932 3108 14936 3140
rect 14896 3072 14936 3108
rect 14896 3040 14900 3072
rect 14900 3040 14932 3072
rect 14932 3040 14936 3072
rect 14896 3004 14936 3040
rect 14896 2972 14900 3004
rect 14900 2972 14932 3004
rect 14932 2972 14936 3004
rect 14896 2936 14936 2972
rect 14896 2904 14900 2936
rect 14900 2904 14932 2936
rect 14932 2904 14936 2936
rect 14896 2868 14936 2904
rect 14896 2836 14900 2868
rect 14900 2836 14932 2868
rect 14932 2836 14936 2868
rect 14896 2800 14936 2836
rect 14896 2768 14900 2800
rect 14900 2768 14932 2800
rect 14932 2768 14936 2800
rect 14896 2732 14936 2768
rect 14896 2700 14900 2732
rect 14900 2700 14932 2732
rect 14932 2700 14936 2732
rect 14896 2664 14936 2700
rect 14896 2632 14900 2664
rect 14900 2632 14932 2664
rect 14932 2632 14936 2664
rect 14896 2596 14936 2632
rect 14896 2564 14900 2596
rect 14900 2564 14932 2596
rect 14932 2564 14936 2596
rect 14896 2528 14936 2564
rect 14896 2496 14900 2528
rect 14900 2496 14932 2528
rect 14932 2496 14936 2528
rect 14896 2460 14936 2496
rect 14896 2428 14900 2460
rect 14900 2428 14932 2460
rect 14932 2428 14936 2460
rect 14896 2392 14936 2428
rect 14896 2360 14900 2392
rect 14900 2360 14932 2392
rect 14932 2360 14936 2392
rect 14896 2324 14936 2360
rect 14896 2318 14900 2324
rect 14900 2318 14932 2324
rect 14932 2318 14936 2324
rect 14896 2142 14900 2148
rect 14900 2142 14932 2148
rect 14932 2142 14936 2148
rect 14896 2106 14936 2142
rect 14896 2074 14900 2106
rect 14900 2074 14932 2106
rect 14932 2074 14936 2106
rect 14896 2038 14936 2074
rect 14896 2006 14900 2038
rect 14900 2006 14932 2038
rect 14932 2006 14936 2038
rect 14896 1970 14936 2006
rect 14896 1938 14900 1970
rect 14900 1938 14932 1970
rect 14932 1938 14936 1970
rect 14896 1902 14936 1938
rect 14896 1870 14900 1902
rect 14900 1870 14932 1902
rect 14932 1870 14936 1902
rect 14896 1834 14936 1870
rect 14896 1802 14900 1834
rect 14900 1802 14932 1834
rect 14932 1802 14936 1834
rect 14896 1766 14936 1802
rect 14896 1734 14900 1766
rect 14900 1734 14932 1766
rect 14932 1734 14936 1766
rect 14896 1698 14936 1734
rect 14896 1666 14900 1698
rect 14900 1666 14932 1698
rect 14932 1666 14936 1698
rect 14896 1630 14936 1666
rect 14896 1598 14900 1630
rect 14900 1598 14932 1630
rect 14932 1598 14936 1630
rect 14896 1562 14936 1598
rect 14896 1530 14900 1562
rect 14900 1530 14932 1562
rect 14932 1530 14936 1562
rect 14896 1494 14936 1530
rect 14896 1462 14900 1494
rect 14900 1462 14932 1494
rect 14932 1462 14936 1494
rect 14896 1426 14936 1462
rect 14896 1394 14900 1426
rect 14900 1394 14932 1426
rect 14932 1394 14936 1426
rect 14896 1358 14936 1394
rect 14896 1326 14900 1358
rect 14900 1326 14932 1358
rect 14932 1326 14936 1358
rect 14896 1290 14936 1326
rect 14896 1258 14900 1290
rect 14900 1258 14932 1290
rect 14932 1258 14936 1290
rect 14896 1222 14936 1258
rect 14896 1190 14900 1222
rect 14900 1190 14932 1222
rect 14932 1190 14936 1222
rect 14896 1154 14936 1190
rect 14896 1122 14900 1154
rect 14900 1122 14932 1154
rect 14932 1122 14936 1154
rect 14896 1086 14936 1122
rect 14896 1054 14900 1086
rect 14900 1054 14932 1086
rect 14932 1054 14936 1086
rect 14896 1018 14936 1054
rect 14896 986 14900 1018
rect 14900 986 14932 1018
rect 14932 986 14936 1018
rect 14896 950 14936 986
rect 14896 918 14900 950
rect 14900 918 14932 950
rect 14932 918 14936 950
rect 14896 882 14936 918
rect 14896 850 14900 882
rect 14900 850 14932 882
rect 14932 850 14936 882
rect 14896 814 14936 850
rect 14896 782 14900 814
rect 14900 782 14932 814
rect 14932 782 14936 814
rect 14896 746 14936 782
rect 14896 714 14900 746
rect 14900 714 14932 746
rect 14932 714 14936 746
rect 14896 678 14936 714
rect 14896 646 14900 678
rect 14900 646 14932 678
rect 14932 646 14936 678
rect 14896 610 14936 646
rect 14896 578 14900 610
rect 14900 578 14932 610
rect 14932 578 14936 610
rect 14896 542 14936 578
rect 14896 510 14900 542
rect 14900 510 14932 542
rect 14932 510 14936 542
rect 14896 474 14936 510
rect 14896 468 14900 474
rect 14900 468 14932 474
rect 14932 468 14936 474
rect 15248 3992 15252 3998
rect 15252 3992 15284 3998
rect 15284 3992 15288 3998
rect 15248 3956 15288 3992
rect 15248 3924 15252 3956
rect 15252 3924 15284 3956
rect 15284 3924 15288 3956
rect 15248 3888 15288 3924
rect 15248 3856 15252 3888
rect 15252 3856 15284 3888
rect 15284 3856 15288 3888
rect 15248 3820 15288 3856
rect 15248 3788 15252 3820
rect 15252 3788 15284 3820
rect 15284 3788 15288 3820
rect 15248 3752 15288 3788
rect 15248 3720 15252 3752
rect 15252 3720 15284 3752
rect 15284 3720 15288 3752
rect 15248 3684 15288 3720
rect 15248 3652 15252 3684
rect 15252 3652 15284 3684
rect 15284 3652 15288 3684
rect 15248 3616 15288 3652
rect 15248 3584 15252 3616
rect 15252 3584 15284 3616
rect 15284 3584 15288 3616
rect 15248 3548 15288 3584
rect 15248 3516 15252 3548
rect 15252 3516 15284 3548
rect 15284 3516 15288 3548
rect 15248 3480 15288 3516
rect 15248 3448 15252 3480
rect 15252 3448 15284 3480
rect 15284 3448 15288 3480
rect 15248 3412 15288 3448
rect 15248 3380 15252 3412
rect 15252 3380 15284 3412
rect 15284 3380 15288 3412
rect 15248 3344 15288 3380
rect 15248 3312 15252 3344
rect 15252 3312 15284 3344
rect 15284 3312 15288 3344
rect 15248 3276 15288 3312
rect 15248 3244 15252 3276
rect 15252 3244 15284 3276
rect 15284 3244 15288 3276
rect 15248 3208 15288 3244
rect 15248 3176 15252 3208
rect 15252 3176 15284 3208
rect 15284 3176 15288 3208
rect 15248 3140 15288 3176
rect 15248 3108 15252 3140
rect 15252 3108 15284 3140
rect 15284 3108 15288 3140
rect 15248 3072 15288 3108
rect 15248 3040 15252 3072
rect 15252 3040 15284 3072
rect 15284 3040 15288 3072
rect 15248 3004 15288 3040
rect 15248 2972 15252 3004
rect 15252 2972 15284 3004
rect 15284 2972 15288 3004
rect 15248 2936 15288 2972
rect 15248 2904 15252 2936
rect 15252 2904 15284 2936
rect 15284 2904 15288 2936
rect 15248 2868 15288 2904
rect 15248 2836 15252 2868
rect 15252 2836 15284 2868
rect 15284 2836 15288 2868
rect 15248 2800 15288 2836
rect 15248 2768 15252 2800
rect 15252 2768 15284 2800
rect 15284 2768 15288 2800
rect 15248 2732 15288 2768
rect 15248 2700 15252 2732
rect 15252 2700 15284 2732
rect 15284 2700 15288 2732
rect 15248 2664 15288 2700
rect 15248 2632 15252 2664
rect 15252 2632 15284 2664
rect 15284 2632 15288 2664
rect 15248 2596 15288 2632
rect 15248 2564 15252 2596
rect 15252 2564 15284 2596
rect 15284 2564 15288 2596
rect 15248 2528 15288 2564
rect 15248 2496 15252 2528
rect 15252 2496 15284 2528
rect 15284 2496 15288 2528
rect 15248 2460 15288 2496
rect 15248 2428 15252 2460
rect 15252 2428 15284 2460
rect 15284 2428 15288 2460
rect 15248 2392 15288 2428
rect 15248 2360 15252 2392
rect 15252 2360 15284 2392
rect 15284 2360 15288 2392
rect 15248 2324 15288 2360
rect 15248 2318 15252 2324
rect 15252 2318 15284 2324
rect 15284 2318 15288 2324
rect 15248 2142 15252 2148
rect 15252 2142 15284 2148
rect 15284 2142 15288 2148
rect 15248 2106 15288 2142
rect 15248 2074 15252 2106
rect 15252 2074 15284 2106
rect 15284 2074 15288 2106
rect 15248 2038 15288 2074
rect 15248 2006 15252 2038
rect 15252 2006 15284 2038
rect 15284 2006 15288 2038
rect 15248 1970 15288 2006
rect 15248 1938 15252 1970
rect 15252 1938 15284 1970
rect 15284 1938 15288 1970
rect 15248 1902 15288 1938
rect 15248 1870 15252 1902
rect 15252 1870 15284 1902
rect 15284 1870 15288 1902
rect 15248 1834 15288 1870
rect 15248 1802 15252 1834
rect 15252 1802 15284 1834
rect 15284 1802 15288 1834
rect 15248 1766 15288 1802
rect 15248 1734 15252 1766
rect 15252 1734 15284 1766
rect 15284 1734 15288 1766
rect 15248 1698 15288 1734
rect 15248 1666 15252 1698
rect 15252 1666 15284 1698
rect 15284 1666 15288 1698
rect 15248 1630 15288 1666
rect 15248 1598 15252 1630
rect 15252 1598 15284 1630
rect 15284 1598 15288 1630
rect 15248 1562 15288 1598
rect 15248 1530 15252 1562
rect 15252 1530 15284 1562
rect 15284 1530 15288 1562
rect 15248 1494 15288 1530
rect 15248 1462 15252 1494
rect 15252 1462 15284 1494
rect 15284 1462 15288 1494
rect 15248 1426 15288 1462
rect 15248 1394 15252 1426
rect 15252 1394 15284 1426
rect 15284 1394 15288 1426
rect 15248 1358 15288 1394
rect 15248 1326 15252 1358
rect 15252 1326 15284 1358
rect 15284 1326 15288 1358
rect 15248 1290 15288 1326
rect 15248 1258 15252 1290
rect 15252 1258 15284 1290
rect 15284 1258 15288 1290
rect 15248 1222 15288 1258
rect 15248 1190 15252 1222
rect 15252 1190 15284 1222
rect 15284 1190 15288 1222
rect 15248 1154 15288 1190
rect 15248 1122 15252 1154
rect 15252 1122 15284 1154
rect 15284 1122 15288 1154
rect 15248 1086 15288 1122
rect 15248 1054 15252 1086
rect 15252 1054 15284 1086
rect 15284 1054 15288 1086
rect 15248 1018 15288 1054
rect 15248 986 15252 1018
rect 15252 986 15284 1018
rect 15284 986 15288 1018
rect 15248 950 15288 986
rect 15248 918 15252 950
rect 15252 918 15284 950
rect 15284 918 15288 950
rect 15248 882 15288 918
rect 15248 850 15252 882
rect 15252 850 15284 882
rect 15284 850 15288 882
rect 15248 814 15288 850
rect 15248 782 15252 814
rect 15252 782 15284 814
rect 15284 782 15288 814
rect 15248 746 15288 782
rect 15248 714 15252 746
rect 15252 714 15284 746
rect 15284 714 15288 746
rect 15248 678 15288 714
rect 15248 646 15252 678
rect 15252 646 15284 678
rect 15284 646 15288 678
rect 15248 610 15288 646
rect 15248 578 15252 610
rect 15252 578 15284 610
rect 15284 578 15288 610
rect 15248 542 15288 578
rect 15248 510 15252 542
rect 15252 510 15284 542
rect 15284 510 15288 542
rect 15248 474 15288 510
rect 15248 468 15252 474
rect 15252 468 15284 474
rect 15284 468 15288 474
rect 641 302 15359 342
<< metal2 >>
rect 594 6744 3675 6784
rect 12325 6744 12362 6784
rect 594 342 3630 6744
rect 3756 6617 15288 6660
rect 3796 5347 4108 6617
rect 4148 5347 4460 6617
rect 4500 5347 4812 6617
rect 4852 5347 5164 6617
rect 5204 5347 5516 6617
rect 5556 5347 5868 6617
rect 5908 5347 6220 6617
rect 6260 5347 6572 6617
rect 6612 5347 6924 6617
rect 6964 5347 7276 6617
rect 7316 5347 7628 6617
rect 7668 5347 7980 6617
rect 8020 5347 8332 6617
rect 8372 5347 8684 6617
rect 8724 5347 9036 6617
rect 9076 5347 9388 6617
rect 9428 5347 9740 6617
rect 9780 5347 10092 6617
rect 10132 5347 10444 6617
rect 10484 5347 10796 6617
rect 10836 5347 11148 6617
rect 11188 5347 11500 6617
rect 11540 5347 11852 6617
rect 11892 5347 12204 6617
rect 12244 5347 15288 6617
rect 3756 5304 15288 5347
rect 14544 3998 15288 5304
rect 14584 2318 14896 3998
rect 14936 2318 15248 3998
rect 14544 2148 15288 2318
rect 14584 468 14896 2148
rect 14936 468 15248 2148
rect 14544 426 15288 468
rect 594 302 641 342
rect 15359 302 15406 342
<< labels >>
flabel metal1 s 18 4406 228 4456 0 FreeSans 51 0 0 0 iovss
port 9 nsew
rlabel metal1 s 3264 7022 12736 7090 4 supply
port 1 nsew
rlabel metal2 s 14544 426 15288 6660 4 out
port 3 nsew
rlabel metal2 s 594 302 3630 6784 4 in
port 2 nsew
rlabel comment s 34 34 34 34 4 sub!
<< properties >>
string device primitive
string GDS_END 806518
string GDS_FILE sg13g2_io.gds
string GDS_START 548914
<< end >>
