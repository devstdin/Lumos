magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757368577
<< poly >>
rect -224 326 56 362
rect -224 294 -199 326
rect -167 294 -131 326
rect -99 294 -63 326
rect -31 294 56 326
rect -224 258 56 294
rect -224 226 -199 258
rect -167 226 -131 258
rect -99 226 -63 258
rect -31 226 56 258
rect -224 190 56 226
rect -224 158 -199 190
rect -167 158 -131 190
rect -99 158 -63 190
rect -31 188 56 190
rect 256 326 536 362
rect 256 294 342 326
rect 374 294 410 326
rect 442 294 478 326
rect 510 294 536 326
rect 256 258 536 294
rect 256 226 342 258
rect 374 226 410 258
rect 442 226 478 258
rect 510 226 536 258
rect 256 190 536 226
rect 256 188 342 190
rect -31 160 107 188
rect 205 160 342 188
rect -31 158 56 160
rect -224 122 56 158
rect -224 90 -199 122
rect -167 90 -131 122
rect -99 90 -63 122
rect -31 90 56 122
rect -224 54 56 90
rect -224 22 -199 54
rect -167 22 -131 54
rect -99 22 -63 54
rect -31 22 56 54
rect -224 -14 56 22
rect 256 158 342 160
rect 374 158 410 190
rect 442 158 478 190
rect 510 158 536 190
rect 256 122 536 158
rect 256 90 342 122
rect 374 90 410 122
rect 442 90 478 122
rect 510 90 536 122
rect 256 54 536 90
rect 256 22 342 54
rect 374 22 410 54
rect 442 22 478 54
rect 510 22 536 54
rect 256 -14 536 22
<< polycont >>
rect -199 294 -167 326
rect -131 294 -99 326
rect -63 294 -31 326
rect -199 226 -167 258
rect -131 226 -99 258
rect -63 226 -31 258
rect -199 158 -167 190
rect -131 158 -99 190
rect -63 158 -31 190
rect 342 294 374 326
rect 410 294 442 326
rect 478 294 510 326
rect 342 226 374 258
rect 410 226 442 258
rect 478 226 510 258
rect -199 90 -167 122
rect -131 90 -99 122
rect -63 90 -31 122
rect -199 22 -167 54
rect -131 22 -99 54
rect -63 22 -31 54
rect 342 158 374 190
rect 410 158 442 190
rect 478 158 510 190
rect 342 90 374 122
rect 410 90 442 122
rect 478 90 510 122
rect 342 22 374 54
rect 410 22 442 54
rect 478 22 510 54
<< metal1 >>
rect -586 1403 -5 1441
rect -586 1363 -556 1403
rect -516 1363 -460 1403
rect -420 1363 -364 1403
rect -324 1363 -268 1403
rect -228 1363 -172 1403
rect -132 1363 -76 1403
rect -36 1363 -5 1403
rect -586 1307 -5 1363
rect -586 1267 -556 1307
rect -516 1267 -460 1307
rect -420 1267 -364 1307
rect -324 1267 -268 1307
rect -228 1267 -172 1307
rect -132 1267 -76 1307
rect -36 1267 -5 1307
rect -586 1211 -5 1267
rect -586 1171 -556 1211
rect -516 1171 -460 1211
rect -420 1171 -364 1211
rect -324 1171 -268 1211
rect -228 1171 -172 1211
rect -132 1171 -76 1211
rect -36 1171 -5 1211
rect -586 1115 -5 1171
rect -586 1075 -556 1115
rect -516 1075 -460 1115
rect -420 1075 -364 1115
rect -324 1075 -268 1115
rect -228 1075 -172 1115
rect -132 1075 -76 1115
rect -36 1075 -5 1115
rect -586 1019 -5 1075
rect -586 979 -556 1019
rect -516 979 -460 1019
rect -420 979 -364 1019
rect -324 979 -268 1019
rect -228 979 -172 1019
rect -132 979 -76 1019
rect -36 979 -5 1019
rect -586 923 -5 979
rect -586 883 -556 923
rect -516 883 -460 923
rect -420 883 -364 923
rect -324 883 -268 923
rect -228 883 -172 923
rect -132 883 -76 923
rect -36 883 -5 923
rect -586 827 -5 883
rect -586 787 -556 827
rect -516 787 -460 827
rect -420 787 -364 827
rect -324 787 -268 827
rect -228 787 -172 827
rect -132 787 -76 827
rect -36 787 -5 827
rect -586 731 -5 787
rect -586 691 -556 731
rect -516 691 -460 731
rect -420 691 -364 731
rect -324 691 -268 731
rect -228 691 -172 731
rect -132 691 -76 731
rect -36 691 -5 731
rect -586 635 -5 691
rect -586 595 -556 635
rect -516 595 -460 635
rect -420 595 -364 635
rect -324 595 -268 635
rect -228 595 -172 635
rect -132 595 -76 635
rect -36 595 -5 635
rect -586 539 -5 595
rect -586 499 -556 539
rect -516 499 -460 539
rect -420 499 -364 539
rect -324 499 -268 539
rect -228 499 -172 539
rect -132 499 -76 539
rect -36 499 -5 539
rect -586 443 -5 499
rect -586 403 -556 443
rect -516 403 -460 443
rect -420 403 -364 443
rect -324 403 -268 443
rect -228 403 -172 443
rect -132 403 -76 443
rect -36 403 -5 443
rect -586 347 -5 403
rect -586 307 -556 347
rect -516 307 -460 347
rect -420 307 -364 347
rect -324 307 -268 347
rect -228 326 -172 347
rect -132 326 -76 347
rect -36 326 -5 347
rect -228 307 -199 326
rect -132 307 -131 326
rect -586 294 -199 307
rect -167 294 -131 307
rect -99 307 -76 326
rect -99 294 -63 307
rect -31 294 -5 326
rect -586 258 -5 294
rect -586 251 -199 258
rect -167 251 -131 258
rect -586 211 -556 251
rect -516 211 -460 251
rect -420 211 -364 251
rect -324 211 -268 251
rect -228 226 -199 251
rect -132 226 -131 251
rect -99 251 -63 258
rect -99 226 -76 251
rect -31 226 -5 258
rect -228 211 -172 226
rect -132 211 -76 226
rect -36 211 -5 226
rect -586 190 -5 211
rect -586 158 -199 190
rect -167 158 -131 190
rect -99 158 -63 190
rect -31 158 -5 190
rect -586 155 -5 158
rect -586 115 -556 155
rect -516 115 -460 155
rect -420 115 -364 155
rect -324 115 -268 155
rect -228 122 -172 155
rect -132 122 -76 155
rect -36 122 -5 155
rect -228 115 -199 122
rect -132 115 -131 122
rect -586 90 -199 115
rect -167 90 -131 115
rect -99 115 -76 122
rect -99 90 -63 115
rect -31 90 -5 122
rect -586 59 -5 90
rect -586 19 -556 59
rect -516 19 -460 59
rect -420 19 -364 59
rect -324 19 -268 59
rect -228 54 -172 59
rect -132 54 -76 59
rect -36 54 -5 59
rect -228 22 -199 54
rect -132 22 -131 54
rect -99 22 -76 54
rect -31 22 -5 54
rect -228 19 -172 22
rect -132 19 -76 22
rect -36 19 -5 22
rect -586 -37 -5 19
rect -586 -77 -556 -37
rect -516 -77 -460 -37
rect -420 -77 -364 -37
rect -324 -77 -268 -37
rect -228 -77 -172 -37
rect -132 -77 -76 -37
rect -36 -77 -5 -37
rect -586 -133 -5 -77
rect -586 -173 -556 -133
rect -516 -173 -460 -133
rect -420 -173 -364 -133
rect -324 -173 -268 -133
rect -228 -173 -172 -133
rect -132 -173 -76 -133
rect -36 -173 -5 -133
rect -586 -229 -5 -173
rect -586 -269 -556 -229
rect -516 -269 -460 -229
rect -420 -269 -364 -229
rect -324 -269 -268 -229
rect -228 -269 -172 -229
rect -132 -269 -76 -229
rect -36 -269 -5 -229
rect 317 586 657 622
rect 317 546 371 586
rect 411 546 467 586
rect 507 546 563 586
rect 603 546 657 586
rect 317 490 657 546
rect 317 450 371 490
rect 411 450 467 490
rect 507 450 563 490
rect 603 450 657 490
rect 317 394 657 450
rect 317 354 371 394
rect 411 354 467 394
rect 507 354 563 394
rect 603 354 657 394
rect 317 326 657 354
rect 317 294 342 326
rect 374 298 410 326
rect 442 298 478 326
rect 510 298 657 326
rect 442 294 467 298
rect 510 294 563 298
rect 317 258 371 294
rect 411 258 467 294
rect 507 258 563 294
rect 603 258 657 298
rect 317 226 342 258
rect 374 226 410 258
rect 442 226 478 258
rect 510 226 657 258
rect 317 202 657 226
rect 317 190 371 202
rect 411 190 467 202
rect 507 190 563 202
rect 317 158 342 190
rect 442 162 467 190
rect 510 162 563 190
rect 603 162 657 202
rect 374 158 410 162
rect 442 158 478 162
rect 510 158 657 162
rect 317 122 657 158
rect 317 90 342 122
rect 374 106 410 122
rect 442 106 478 122
rect 510 106 657 122
rect 442 90 467 106
rect 510 90 563 106
rect 317 66 371 90
rect 411 66 467 90
rect 507 66 563 90
rect 603 66 657 106
rect 317 54 657 66
rect 317 22 342 54
rect 374 22 410 54
rect 442 22 478 54
rect 510 22 657 54
rect 317 10 657 22
rect 317 -30 371 10
rect 411 -30 467 10
rect 507 -30 563 10
rect 603 -30 657 10
rect 317 -86 657 -30
rect 317 -126 371 -86
rect 411 -126 467 -86
rect 507 -126 563 -86
rect 603 -126 657 -86
rect 317 -182 657 -126
rect 317 -222 371 -182
rect 411 -222 467 -182
rect 507 -222 563 -182
rect 603 -222 657 -182
rect 317 -258 657 -222
rect -586 -325 -5 -269
rect -586 -365 -556 -325
rect -516 -365 -460 -325
rect -420 -365 -364 -325
rect -324 -365 -268 -325
rect -228 -365 -172 -325
rect -132 -365 -76 -325
rect -36 -365 -5 -325
rect -586 -421 -5 -365
rect -586 -461 -556 -421
rect -516 -461 -460 -421
rect -420 -461 -364 -421
rect -324 -461 -268 -421
rect -228 -461 -172 -421
rect -132 -461 -76 -421
rect -36 -461 -5 -421
rect -586 -517 -5 -461
rect -586 -557 -556 -517
rect -516 -557 -460 -517
rect -420 -557 -364 -517
rect -324 -557 -268 -517
rect -228 -557 -172 -517
rect -132 -557 -76 -517
rect -36 -557 -5 -517
rect -586 -613 -5 -557
rect -586 -653 -556 -613
rect -516 -653 -460 -613
rect -420 -653 -364 -613
rect -324 -653 -268 -613
rect -228 -653 -172 -613
rect -132 -653 -76 -613
rect -36 -653 -5 -613
rect -586 -709 -5 -653
rect -586 -749 -556 -709
rect -516 -749 -460 -709
rect -420 -749 -364 -709
rect -324 -749 -268 -709
rect -228 -749 -172 -709
rect -132 -749 -76 -709
rect -36 -749 -5 -709
rect -586 -805 -5 -749
rect -586 -845 -556 -805
rect -516 -845 -460 -805
rect -420 -845 -364 -805
rect -324 -845 -268 -805
rect -228 -845 -172 -805
rect -132 -845 -76 -805
rect -36 -845 -5 -805
rect -586 -901 -5 -845
rect -586 -941 -556 -901
rect -516 -941 -460 -901
rect -420 -941 -364 -901
rect -324 -941 -268 -901
rect -228 -941 -172 -901
rect -132 -941 -76 -901
rect -36 -941 -5 -901
rect -586 -997 -5 -941
rect -586 -1037 -556 -997
rect -516 -1037 -460 -997
rect -420 -1037 -364 -997
rect -324 -1037 -268 -997
rect -228 -1037 -172 -997
rect -132 -1037 -76 -997
rect -36 -1037 -5 -997
rect -586 -1075 -5 -1037
<< via1 >>
rect -556 1363 -516 1403
rect -460 1363 -420 1403
rect -364 1363 -324 1403
rect -268 1363 -228 1403
rect -172 1363 -132 1403
rect -76 1363 -36 1403
rect -556 1267 -516 1307
rect -460 1267 -420 1307
rect -364 1267 -324 1307
rect -268 1267 -228 1307
rect -172 1267 -132 1307
rect -76 1267 -36 1307
rect -556 1171 -516 1211
rect -460 1171 -420 1211
rect -364 1171 -324 1211
rect -268 1171 -228 1211
rect -172 1171 -132 1211
rect -76 1171 -36 1211
rect -556 1075 -516 1115
rect -460 1075 -420 1115
rect -364 1075 -324 1115
rect -268 1075 -228 1115
rect -172 1075 -132 1115
rect -76 1075 -36 1115
rect -556 979 -516 1019
rect -460 979 -420 1019
rect -364 979 -324 1019
rect -268 979 -228 1019
rect -172 979 -132 1019
rect -76 979 -36 1019
rect -556 883 -516 923
rect -460 883 -420 923
rect -364 883 -324 923
rect -268 883 -228 923
rect -172 883 -132 923
rect -76 883 -36 923
rect -556 787 -516 827
rect -460 787 -420 827
rect -364 787 -324 827
rect -268 787 -228 827
rect -172 787 -132 827
rect -76 787 -36 827
rect -556 691 -516 731
rect -460 691 -420 731
rect -364 691 -324 731
rect -268 691 -228 731
rect -172 691 -132 731
rect -76 691 -36 731
rect -556 595 -516 635
rect -460 595 -420 635
rect -364 595 -324 635
rect -268 595 -228 635
rect -172 595 -132 635
rect -76 595 -36 635
rect -556 499 -516 539
rect -460 499 -420 539
rect -364 499 -324 539
rect -268 499 -228 539
rect -172 499 -132 539
rect -76 499 -36 539
rect -556 403 -516 443
rect -460 403 -420 443
rect -364 403 -324 443
rect -268 403 -228 443
rect -172 403 -132 443
rect -76 403 -36 443
rect -556 307 -516 347
rect -460 307 -420 347
rect -364 307 -324 347
rect -268 307 -228 347
rect -172 326 -132 347
rect -76 326 -36 347
rect -172 307 -167 326
rect -167 307 -132 326
rect -76 307 -63 326
rect -63 307 -36 326
rect -556 211 -516 251
rect -460 211 -420 251
rect -364 211 -324 251
rect -268 211 -228 251
rect -172 226 -167 251
rect -167 226 -132 251
rect -76 226 -63 251
rect -63 226 -36 251
rect -172 211 -132 226
rect -76 211 -36 226
rect -556 115 -516 155
rect -460 115 -420 155
rect -364 115 -324 155
rect -268 115 -228 155
rect -172 122 -132 155
rect -76 122 -36 155
rect -172 115 -167 122
rect -167 115 -132 122
rect -76 115 -63 122
rect -63 115 -36 122
rect -556 19 -516 59
rect -460 19 -420 59
rect -364 19 -324 59
rect -268 19 -228 59
rect -172 54 -132 59
rect -76 54 -36 59
rect -172 22 -167 54
rect -167 22 -132 54
rect -76 22 -63 54
rect -63 22 -36 54
rect -172 19 -132 22
rect -76 19 -36 22
rect -556 -77 -516 -37
rect -460 -77 -420 -37
rect -364 -77 -324 -37
rect -268 -77 -228 -37
rect -172 -77 -132 -37
rect -76 -77 -36 -37
rect -556 -173 -516 -133
rect -460 -173 -420 -133
rect -364 -173 -324 -133
rect -268 -173 -228 -133
rect -172 -173 -132 -133
rect -76 -173 -36 -133
rect -556 -269 -516 -229
rect -460 -269 -420 -229
rect -364 -269 -324 -229
rect -268 -269 -228 -229
rect -172 -269 -132 -229
rect -76 -269 -36 -229
rect 371 546 411 586
rect 467 546 507 586
rect 563 546 603 586
rect 371 450 411 490
rect 467 450 507 490
rect 563 450 603 490
rect 371 354 411 394
rect 467 354 507 394
rect 563 354 603 394
rect 371 294 374 298
rect 374 294 410 298
rect 410 294 411 298
rect 467 294 478 298
rect 478 294 507 298
rect 371 258 411 294
rect 467 258 507 294
rect 563 258 603 298
rect 371 190 411 202
rect 467 190 507 202
rect 371 162 374 190
rect 374 162 410 190
rect 410 162 411 190
rect 467 162 478 190
rect 478 162 507 190
rect 563 162 603 202
rect 371 90 374 106
rect 374 90 410 106
rect 410 90 411 106
rect 467 90 478 106
rect 478 90 507 106
rect 371 66 411 90
rect 467 66 507 90
rect 563 66 603 106
rect 371 -30 411 10
rect 467 -30 507 10
rect 563 -30 603 10
rect 371 -126 411 -86
rect 467 -126 507 -86
rect 563 -126 603 -86
rect 371 -222 411 -182
rect 467 -222 507 -182
rect 563 -222 603 -182
rect -556 -365 -516 -325
rect -460 -365 -420 -325
rect -364 -365 -324 -325
rect -268 -365 -228 -325
rect -172 -365 -132 -325
rect -76 -365 -36 -325
rect -556 -461 -516 -421
rect -460 -461 -420 -421
rect -364 -461 -324 -421
rect -268 -461 -228 -421
rect -172 -461 -132 -421
rect -76 -461 -36 -421
rect -556 -557 -516 -517
rect -460 -557 -420 -517
rect -364 -557 -324 -517
rect -268 -557 -228 -517
rect -172 -557 -132 -517
rect -76 -557 -36 -517
rect -556 -653 -516 -613
rect -460 -653 -420 -613
rect -364 -653 -324 -613
rect -268 -653 -228 -613
rect -172 -653 -132 -613
rect -76 -653 -36 -613
rect -556 -749 -516 -709
rect -460 -749 -420 -709
rect -364 -749 -324 -709
rect -268 -749 -228 -709
rect -172 -749 -132 -709
rect -76 -749 -36 -709
rect -556 -845 -516 -805
rect -460 -845 -420 -805
rect -364 -845 -324 -805
rect -268 -845 -228 -805
rect -172 -845 -132 -805
rect -76 -845 -36 -805
rect -556 -941 -516 -901
rect -460 -941 -420 -901
rect -364 -941 -324 -901
rect -268 -941 -228 -901
rect -172 -941 -132 -901
rect -76 -941 -36 -901
rect -556 -1037 -516 -997
rect -460 -1037 -420 -997
rect -364 -1037 -324 -997
rect -268 -1037 -228 -997
rect -172 -1037 -132 -997
rect -76 -1037 -36 -997
<< metal2 >>
rect -586 1403 -5 1441
rect -586 1363 -556 1403
rect -516 1363 -460 1403
rect -420 1363 -364 1403
rect -324 1363 -268 1403
rect -228 1363 -172 1403
rect -132 1363 -76 1403
rect -36 1363 -5 1403
rect -586 1307 -5 1363
rect -586 1267 -556 1307
rect -516 1267 -460 1307
rect -420 1267 -364 1307
rect -324 1267 -268 1307
rect -228 1267 -172 1307
rect -132 1267 -76 1307
rect -36 1267 -5 1307
rect -586 1211 -5 1267
rect -586 1171 -556 1211
rect -516 1171 -460 1211
rect -420 1171 -364 1211
rect -324 1171 -268 1211
rect -228 1171 -172 1211
rect -132 1171 -76 1211
rect -36 1171 -5 1211
rect -586 1115 -5 1171
rect -586 1075 -556 1115
rect -516 1075 -460 1115
rect -420 1075 -364 1115
rect -324 1075 -268 1115
rect -228 1075 -172 1115
rect -132 1075 -76 1115
rect -36 1075 -5 1115
rect -586 1019 -5 1075
rect -586 979 -556 1019
rect -516 979 -460 1019
rect -420 979 -364 1019
rect -324 979 -268 1019
rect -228 979 -172 1019
rect -132 979 -76 1019
rect -36 979 -5 1019
rect -586 923 -5 979
rect -586 883 -556 923
rect -516 883 -460 923
rect -420 883 -364 923
rect -324 883 -268 923
rect -228 883 -172 923
rect -132 883 -76 923
rect -36 883 -5 923
rect -586 827 -5 883
rect -586 787 -556 827
rect -516 787 -460 827
rect -420 787 -364 827
rect -324 787 -268 827
rect -228 787 -172 827
rect -132 787 -76 827
rect -36 787 -5 827
rect -586 731 -5 787
rect -586 691 -556 731
rect -516 691 -460 731
rect -420 691 -364 731
rect -324 691 -268 731
rect -228 691 -172 731
rect -132 691 -76 731
rect -36 691 -5 731
rect -586 635 -5 691
rect -586 595 -556 635
rect -516 595 -460 635
rect -420 595 -364 635
rect -324 595 -268 635
rect -228 595 -172 635
rect -132 595 -76 635
rect -36 595 -5 635
rect -586 539 -5 595
rect -586 499 -556 539
rect -516 499 -460 539
rect -420 499 -364 539
rect -324 499 -268 539
rect -228 499 -172 539
rect -132 499 -76 539
rect -36 499 -5 539
rect -586 443 -5 499
rect -586 403 -556 443
rect -516 403 -460 443
rect -420 403 -364 443
rect -324 403 -268 443
rect -228 403 -172 443
rect -132 403 -76 443
rect -36 403 -5 443
rect -586 347 -5 403
rect -586 307 -556 347
rect -516 307 -460 347
rect -420 307 -364 347
rect -324 307 -268 347
rect -228 307 -172 347
rect -132 307 -76 347
rect -36 307 -5 347
rect -586 251 -5 307
rect -586 211 -556 251
rect -516 211 -460 251
rect -420 211 -364 251
rect -324 211 -268 251
rect -228 211 -172 251
rect -132 211 -76 251
rect -36 211 -5 251
rect -586 155 -5 211
rect -586 115 -556 155
rect -516 115 -460 155
rect -420 115 -364 155
rect -324 115 -268 155
rect -228 115 -172 155
rect -132 115 -76 155
rect -36 115 -5 155
rect -586 59 -5 115
rect -586 19 -556 59
rect -516 19 -460 59
rect -420 19 -364 59
rect -324 19 -268 59
rect -228 19 -172 59
rect -132 19 -76 59
rect -36 19 -5 59
rect -586 -37 -5 19
rect -586 -77 -556 -37
rect -516 -77 -460 -37
rect -420 -77 -364 -37
rect -324 -77 -268 -37
rect -228 -77 -172 -37
rect -132 -77 -76 -37
rect -36 -77 -5 -37
rect -586 -133 -5 -77
rect -586 -173 -556 -133
rect -516 -173 -460 -133
rect -420 -173 -364 -133
rect -324 -173 -268 -133
rect -228 -173 -172 -133
rect -132 -173 -76 -133
rect -36 -173 -5 -133
rect -586 -229 -5 -173
rect -586 -269 -556 -229
rect -516 -269 -460 -229
rect -420 -269 -364 -229
rect -324 -269 -268 -229
rect -228 -269 -172 -229
rect -132 -269 -76 -229
rect -36 -269 -5 -229
rect 317 586 657 622
rect 317 546 371 586
rect 411 546 467 586
rect 507 546 563 586
rect 603 546 657 586
rect 317 490 657 546
rect 317 450 371 490
rect 411 450 467 490
rect 507 450 563 490
rect 603 450 657 490
rect 317 394 657 450
rect 317 354 371 394
rect 411 354 467 394
rect 507 354 563 394
rect 603 354 657 394
rect 317 298 657 354
rect 317 258 371 298
rect 411 258 467 298
rect 507 258 563 298
rect 603 258 657 298
rect 317 202 657 258
rect 317 162 371 202
rect 411 162 467 202
rect 507 162 563 202
rect 603 162 657 202
rect 317 106 657 162
rect 317 66 371 106
rect 411 66 467 106
rect 507 66 563 106
rect 603 66 657 106
rect 317 10 657 66
rect 317 -30 371 10
rect 411 -30 467 10
rect 507 -30 563 10
rect 603 -30 657 10
rect 317 -86 657 -30
rect 317 -126 371 -86
rect 411 -126 467 -86
rect 507 -126 563 -86
rect 603 -126 657 -86
rect 317 -182 657 -126
rect 317 -222 371 -182
rect 411 -222 467 -182
rect 507 -222 563 -182
rect 603 -222 657 -182
rect 317 -258 657 -222
rect -586 -325 -5 -269
rect -586 -365 -556 -325
rect -516 -365 -460 -325
rect -420 -365 -364 -325
rect -324 -365 -268 -325
rect -228 -365 -172 -325
rect -132 -365 -76 -325
rect -36 -365 -5 -325
rect -586 -421 -5 -365
rect -586 -461 -556 -421
rect -516 -461 -460 -421
rect -420 -461 -364 -421
rect -324 -461 -268 -421
rect -228 -461 -172 -421
rect -132 -461 -76 -421
rect -36 -461 -5 -421
rect -586 -517 -5 -461
rect -586 -557 -556 -517
rect -516 -557 -460 -517
rect -420 -557 -364 -517
rect -324 -557 -268 -517
rect -228 -557 -172 -517
rect -132 -557 -76 -517
rect -36 -557 -5 -517
rect -586 -613 -5 -557
rect -586 -653 -556 -613
rect -516 -653 -460 -613
rect -420 -653 -364 -613
rect -324 -653 -268 -613
rect -228 -653 -172 -613
rect -132 -653 -76 -613
rect -36 -653 -5 -613
rect -586 -709 -5 -653
rect -586 -749 -556 -709
rect -516 -749 -460 -709
rect -420 -749 -364 -709
rect -324 -749 -268 -709
rect -228 -749 -172 -709
rect -132 -749 -76 -709
rect -36 -749 -5 -709
rect -586 -805 -5 -749
rect -586 -845 -556 -805
rect -516 -845 -460 -805
rect -420 -845 -364 -805
rect -324 -845 -268 -805
rect -228 -845 -172 -805
rect -132 -845 -76 -805
rect -36 -845 -5 -805
rect -586 -901 -5 -845
rect -586 -941 -556 -901
rect -516 -941 -460 -901
rect -420 -941 -364 -901
rect -324 -941 -268 -901
rect -228 -941 -172 -901
rect -132 -941 -76 -901
rect -36 -941 -5 -901
rect -586 -997 -5 -941
rect -586 -1037 -556 -997
rect -516 -1037 -460 -997
rect -420 -1037 -364 -997
rect -324 -1037 -268 -997
rect -228 -1037 -172 -997
rect -132 -1037 -76 -997
rect -36 -1037 -5 -997
rect -586 -1075 -5 -1037
<< via2 >>
rect -556 1363 -516 1403
rect -460 1363 -420 1403
rect -364 1363 -324 1403
rect -268 1363 -228 1403
rect -172 1363 -132 1403
rect -76 1363 -36 1403
rect -556 1267 -516 1307
rect -460 1267 -420 1307
rect -364 1267 -324 1307
rect -268 1267 -228 1307
rect -172 1267 -132 1307
rect -76 1267 -36 1307
rect -556 1171 -516 1211
rect -460 1171 -420 1211
rect -364 1171 -324 1211
rect -268 1171 -228 1211
rect -172 1171 -132 1211
rect -76 1171 -36 1211
rect -556 1075 -516 1115
rect -460 1075 -420 1115
rect -364 1075 -324 1115
rect -268 1075 -228 1115
rect -172 1075 -132 1115
rect -76 1075 -36 1115
rect -556 979 -516 1019
rect -460 979 -420 1019
rect -364 979 -324 1019
rect -268 979 -228 1019
rect -172 979 -132 1019
rect -76 979 -36 1019
rect -556 883 -516 923
rect -460 883 -420 923
rect -364 883 -324 923
rect -268 883 -228 923
rect -172 883 -132 923
rect -76 883 -36 923
rect -556 787 -516 827
rect -460 787 -420 827
rect -364 787 -324 827
rect -268 787 -228 827
rect -172 787 -132 827
rect -76 787 -36 827
rect -556 691 -516 731
rect -460 691 -420 731
rect -364 691 -324 731
rect -268 691 -228 731
rect -172 691 -132 731
rect -76 691 -36 731
rect -556 595 -516 635
rect -460 595 -420 635
rect -364 595 -324 635
rect -268 595 -228 635
rect -172 595 -132 635
rect -76 595 -36 635
rect -556 499 -516 539
rect -460 499 -420 539
rect -364 499 -324 539
rect -268 499 -228 539
rect -172 499 -132 539
rect -76 499 -36 539
rect -556 403 -516 443
rect -460 403 -420 443
rect -364 403 -324 443
rect -268 403 -228 443
rect -172 403 -132 443
rect -76 403 -36 443
rect -556 307 -516 347
rect -460 307 -420 347
rect -364 307 -324 347
rect -268 307 -228 347
rect -172 307 -132 347
rect -76 307 -36 347
rect -556 211 -516 251
rect -460 211 -420 251
rect -364 211 -324 251
rect -268 211 -228 251
rect -172 211 -132 251
rect -76 211 -36 251
rect -556 115 -516 155
rect -460 115 -420 155
rect -364 115 -324 155
rect -268 115 -228 155
rect -172 115 -132 155
rect -76 115 -36 155
rect -556 19 -516 59
rect -460 19 -420 59
rect -364 19 -324 59
rect -268 19 -228 59
rect -172 19 -132 59
rect -76 19 -36 59
rect -556 -77 -516 -37
rect -460 -77 -420 -37
rect -364 -77 -324 -37
rect -268 -77 -228 -37
rect -172 -77 -132 -37
rect -76 -77 -36 -37
rect -556 -173 -516 -133
rect -460 -173 -420 -133
rect -364 -173 -324 -133
rect -268 -173 -228 -133
rect -172 -173 -132 -133
rect -76 -173 -36 -133
rect -556 -269 -516 -229
rect -460 -269 -420 -229
rect -364 -269 -324 -229
rect -268 -269 -228 -229
rect -172 -269 -132 -229
rect -76 -269 -36 -229
rect 371 546 411 586
rect 467 546 507 586
rect 563 546 603 586
rect 371 450 411 490
rect 467 450 507 490
rect 563 450 603 490
rect 371 354 411 394
rect 467 354 507 394
rect 563 354 603 394
rect 371 258 411 298
rect 467 258 507 298
rect 563 258 603 298
rect 371 162 411 202
rect 467 162 507 202
rect 563 162 603 202
rect 371 66 411 106
rect 467 66 507 106
rect 563 66 603 106
rect 371 -30 411 10
rect 467 -30 507 10
rect 563 -30 603 10
rect 371 -126 411 -86
rect 467 -126 507 -86
rect 563 -126 603 -86
rect 371 -222 411 -182
rect 467 -222 507 -182
rect 563 -222 603 -182
rect -556 -365 -516 -325
rect -460 -365 -420 -325
rect -364 -365 -324 -325
rect -268 -365 -228 -325
rect -172 -365 -132 -325
rect -76 -365 -36 -325
rect -556 -461 -516 -421
rect -460 -461 -420 -421
rect -364 -461 -324 -421
rect -268 -461 -228 -421
rect -172 -461 -132 -421
rect -76 -461 -36 -421
rect -556 -557 -516 -517
rect -460 -557 -420 -517
rect -364 -557 -324 -517
rect -268 -557 -228 -517
rect -172 -557 -132 -517
rect -76 -557 -36 -517
rect -556 -653 -516 -613
rect -460 -653 -420 -613
rect -364 -653 -324 -613
rect -268 -653 -228 -613
rect -172 -653 -132 -613
rect -76 -653 -36 -613
rect -556 -749 -516 -709
rect -460 -749 -420 -709
rect -364 -749 -324 -709
rect -268 -749 -228 -709
rect -172 -749 -132 -709
rect -76 -749 -36 -709
rect -556 -845 -516 -805
rect -460 -845 -420 -805
rect -364 -845 -324 -805
rect -268 -845 -228 -805
rect -172 -845 -132 -805
rect -76 -845 -36 -805
rect -556 -941 -516 -901
rect -460 -941 -420 -901
rect -364 -941 -324 -901
rect -268 -941 -228 -901
rect -172 -941 -132 -901
rect -76 -941 -36 -901
rect -556 -1037 -516 -997
rect -460 -1037 -420 -997
rect -364 -1037 -324 -997
rect -268 -1037 -228 -997
rect -172 -1037 -132 -997
rect -76 -1037 -36 -997
<< metal3 >>
rect -586 1403 -5 1441
rect -586 1363 -556 1403
rect -516 1363 -460 1403
rect -420 1363 -364 1403
rect -324 1363 -268 1403
rect -228 1363 -172 1403
rect -132 1363 -76 1403
rect -36 1363 -5 1403
rect -586 1307 -5 1363
rect -586 1267 -556 1307
rect -516 1267 -460 1307
rect -420 1267 -364 1307
rect -324 1267 -268 1307
rect -228 1267 -172 1307
rect -132 1267 -76 1307
rect -36 1267 -5 1307
rect -586 1211 -5 1267
rect -586 1171 -556 1211
rect -516 1171 -460 1211
rect -420 1171 -364 1211
rect -324 1171 -268 1211
rect -228 1171 -172 1211
rect -132 1171 -76 1211
rect -36 1171 -5 1211
rect -586 1115 -5 1171
rect -586 1075 -556 1115
rect -516 1075 -460 1115
rect -420 1075 -364 1115
rect -324 1075 -268 1115
rect -228 1075 -172 1115
rect -132 1075 -76 1115
rect -36 1075 -5 1115
rect -586 1019 -5 1075
rect -586 979 -556 1019
rect -516 979 -460 1019
rect -420 979 -364 1019
rect -324 979 -268 1019
rect -228 979 -172 1019
rect -132 979 -76 1019
rect -36 979 -5 1019
rect -586 923 -5 979
rect -586 883 -556 923
rect -516 883 -460 923
rect -420 883 -364 923
rect -324 883 -268 923
rect -228 883 -172 923
rect -132 883 -76 923
rect -36 883 -5 923
rect -586 827 -5 883
rect -586 787 -556 827
rect -516 787 -460 827
rect -420 787 -364 827
rect -324 787 -268 827
rect -228 787 -172 827
rect -132 787 -76 827
rect -36 787 -5 827
rect -586 731 -5 787
rect -586 691 -556 731
rect -516 691 -460 731
rect -420 691 -364 731
rect -324 691 -268 731
rect -228 691 -172 731
rect -132 691 -76 731
rect -36 691 -5 731
rect -586 635 -5 691
rect -586 595 -556 635
rect -516 595 -460 635
rect -420 595 -364 635
rect -324 595 -268 635
rect -228 595 -172 635
rect -132 595 -76 635
rect -36 595 -5 635
rect -586 539 -5 595
rect -586 499 -556 539
rect -516 499 -460 539
rect -420 499 -364 539
rect -324 499 -268 539
rect -228 499 -172 539
rect -132 499 -76 539
rect -36 499 -5 539
rect -586 443 -5 499
rect -586 403 -556 443
rect -516 403 -460 443
rect -420 403 -364 443
rect -324 403 -268 443
rect -228 403 -172 443
rect -132 403 -76 443
rect -36 403 -5 443
rect -586 347 -5 403
rect -586 307 -556 347
rect -516 307 -460 347
rect -420 307 -364 347
rect -324 307 -268 347
rect -228 307 -172 347
rect -132 307 -76 347
rect -36 307 -5 347
rect -586 251 -5 307
rect -586 211 -556 251
rect -516 211 -460 251
rect -420 211 -364 251
rect -324 211 -268 251
rect -228 211 -172 251
rect -132 211 -76 251
rect -36 211 -5 251
rect -586 155 -5 211
rect -586 115 -556 155
rect -516 115 -460 155
rect -420 115 -364 155
rect -324 115 -268 155
rect -228 115 -172 155
rect -132 115 -76 155
rect -36 115 -5 155
rect -586 59 -5 115
rect -586 19 -556 59
rect -516 19 -460 59
rect -420 19 -364 59
rect -324 19 -268 59
rect -228 19 -172 59
rect -132 19 -76 59
rect -36 19 -5 59
rect -586 -37 -5 19
rect -586 -77 -556 -37
rect -516 -77 -460 -37
rect -420 -77 -364 -37
rect -324 -77 -268 -37
rect -228 -77 -172 -37
rect -132 -77 -76 -37
rect -36 -77 -5 -37
rect -586 -133 -5 -77
rect -586 -173 -556 -133
rect -516 -173 -460 -133
rect -420 -173 -364 -133
rect -324 -173 -268 -133
rect -228 -173 -172 -133
rect -132 -173 -76 -133
rect -36 -173 -5 -133
rect -586 -229 -5 -173
rect -586 -269 -556 -229
rect -516 -269 -460 -229
rect -420 -269 -364 -229
rect -324 -269 -268 -229
rect -228 -269 -172 -229
rect -132 -269 -76 -229
rect -36 -269 -5 -229
rect 317 586 657 622
rect 317 546 371 586
rect 411 546 467 586
rect 507 546 563 586
rect 603 546 657 586
rect 317 490 657 546
rect 317 450 371 490
rect 411 450 467 490
rect 507 450 563 490
rect 603 450 657 490
rect 317 394 657 450
rect 317 354 371 394
rect 411 354 467 394
rect 507 354 563 394
rect 603 354 657 394
rect 317 298 657 354
rect 317 258 371 298
rect 411 258 467 298
rect 507 258 563 298
rect 603 258 657 298
rect 317 202 657 258
rect 317 162 371 202
rect 411 162 467 202
rect 507 162 563 202
rect 603 162 657 202
rect 317 106 657 162
rect 317 66 371 106
rect 411 66 467 106
rect 507 66 563 106
rect 603 66 657 106
rect 317 10 657 66
rect 317 -30 371 10
rect 411 -30 467 10
rect 507 -30 563 10
rect 603 -30 657 10
rect 317 -86 657 -30
rect 317 -126 371 -86
rect 411 -126 467 -86
rect 507 -126 563 -86
rect 603 -126 657 -86
rect 317 -182 657 -126
rect 317 -222 371 -182
rect 411 -222 467 -182
rect 507 -222 563 -182
rect 603 -222 657 -182
rect 317 -258 657 -222
rect -586 -325 -5 -269
rect -586 -365 -556 -325
rect -516 -365 -460 -325
rect -420 -365 -364 -325
rect -324 -365 -268 -325
rect -228 -365 -172 -325
rect -132 -365 -76 -325
rect -36 -365 -5 -325
rect -586 -421 -5 -365
rect -586 -461 -556 -421
rect -516 -461 -460 -421
rect -420 -461 -364 -421
rect -324 -461 -268 -421
rect -228 -461 -172 -421
rect -132 -461 -76 -421
rect -36 -461 -5 -421
rect -586 -517 -5 -461
rect -586 -557 -556 -517
rect -516 -557 -460 -517
rect -420 -557 -364 -517
rect -324 -557 -268 -517
rect -228 -557 -172 -517
rect -132 -557 -76 -517
rect -36 -557 -5 -517
rect -586 -613 -5 -557
rect -586 -653 -556 -613
rect -516 -653 -460 -613
rect -420 -653 -364 -613
rect -324 -653 -268 -613
rect -228 -653 -172 -613
rect -132 -653 -76 -613
rect -36 -653 -5 -613
rect -586 -709 -5 -653
rect -586 -749 -556 -709
rect -516 -749 -460 -709
rect -420 -749 -364 -709
rect -324 -749 -268 -709
rect -228 -749 -172 -709
rect -132 -749 -76 -709
rect -36 -749 -5 -709
rect -586 -805 -5 -749
rect -586 -845 -556 -805
rect -516 -845 -460 -805
rect -420 -845 -364 -805
rect -324 -845 -268 -805
rect -228 -845 -172 -805
rect -132 -845 -76 -805
rect -36 -845 -5 -805
rect -586 -901 -5 -845
rect -586 -941 -556 -901
rect -516 -941 -460 -901
rect -420 -941 -364 -901
rect -324 -941 -268 -901
rect -228 -941 -172 -901
rect -132 -941 -76 -901
rect -36 -941 -5 -901
rect -586 -997 -5 -941
rect -586 -1037 -556 -997
rect -516 -1037 -460 -997
rect -420 -1037 -364 -997
rect -324 -1037 -268 -997
rect -228 -1037 -172 -997
rect -132 -1037 -76 -997
rect -36 -1037 -5 -997
rect -586 -1075 -5 -1037
<< fillblock >>
rect -284 -194 596 542
<< labels >>
flabel metal3 s -586 -1075 -427 1441 0 FreeSans 1000 0 0 0 T1
port 1 nsew
flabel metal3 s 527 -258 657 622 0 FreeSans 1000 0 0 0 T2
port 2 nsew
<< properties >>
string device primitive
string GDS_END 26478
string GDS_FILE fuse_prim.gds
string GDS_START 110
<< end >>
