magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2005 2604 4524
<< nwell >>
rect -124 1152 604 2524
<< pwell >>
rect -5 107 315 1054
rect -5 -5 485 107
<< nmos >>
rect 89 242 115 1028
rect 191 242 217 1028
<< pmos >>
rect 89 1276 115 2158
rect 191 1276 217 2158
<< ndiff >>
rect 21 288 89 1028
rect 21 256 35 288
rect 67 256 89 288
rect 21 242 89 256
rect 115 999 191 1028
rect 115 967 137 999
rect 169 967 191 999
rect 115 931 191 967
rect 115 899 137 931
rect 169 899 191 931
rect 115 863 191 899
rect 115 831 137 863
rect 169 831 191 863
rect 115 795 191 831
rect 115 763 137 795
rect 169 763 191 795
rect 115 727 191 763
rect 115 695 137 727
rect 169 695 191 727
rect 115 659 191 695
rect 115 627 137 659
rect 169 627 191 659
rect 115 591 191 627
rect 115 559 137 591
rect 169 559 191 591
rect 115 523 191 559
rect 115 491 137 523
rect 169 491 191 523
rect 115 455 191 491
rect 115 423 137 455
rect 169 423 191 455
rect 115 387 191 423
rect 115 355 137 387
rect 169 355 191 387
rect 115 242 191 355
rect 217 288 289 1028
rect 217 256 243 288
rect 275 256 289 288
rect 217 242 289 256
<< pdiff >>
rect 21 2144 89 2158
rect 21 2112 35 2144
rect 67 2112 89 2144
rect 21 1276 89 2112
rect 115 1276 191 2158
rect 217 2031 289 2158
rect 217 1999 243 2031
rect 275 1999 289 2031
rect 217 1963 289 1999
rect 217 1931 243 1963
rect 275 1931 289 1963
rect 217 1895 289 1931
rect 217 1863 243 1895
rect 275 1863 289 1895
rect 217 1827 289 1863
rect 217 1795 243 1827
rect 275 1795 289 1827
rect 217 1759 289 1795
rect 217 1727 243 1759
rect 275 1727 289 1759
rect 217 1691 289 1727
rect 217 1659 243 1691
rect 275 1659 289 1691
rect 217 1623 289 1659
rect 217 1591 243 1623
rect 275 1591 289 1623
rect 217 1555 289 1591
rect 217 1523 243 1555
rect 275 1523 289 1555
rect 217 1487 289 1523
rect 217 1455 243 1487
rect 275 1455 289 1487
rect 217 1419 289 1455
rect 217 1387 243 1419
rect 275 1387 289 1419
rect 217 1351 289 1387
rect 217 1319 243 1351
rect 275 1319 289 1351
rect 217 1276 289 1319
<< ndiffc >>
rect 35 256 67 288
rect 137 967 169 999
rect 137 899 169 931
rect 137 831 169 863
rect 137 763 169 795
rect 137 695 169 727
rect 137 627 169 659
rect 137 559 169 591
rect 137 491 169 523
rect 137 423 169 455
rect 137 355 169 387
rect 243 256 275 288
<< pdiffc >>
rect 35 2112 67 2144
rect 243 1999 275 2031
rect 243 1931 275 1963
rect 243 1863 275 1895
rect 243 1795 275 1827
rect 243 1727 275 1759
rect 243 1659 275 1691
rect 243 1591 275 1623
rect 243 1523 275 1555
rect 243 1455 275 1487
rect 243 1387 275 1419
rect 243 1319 275 1351
<< psubdiff >>
rect 21 67 459 81
rect 21 35 54 67
rect 86 35 122 67
rect 154 35 190 67
rect 222 35 258 67
rect 290 35 326 67
rect 358 35 394 67
rect 426 35 459 67
rect 21 21 459 35
<< nsubdiff >>
rect 21 2365 459 2379
rect 21 2333 54 2365
rect 86 2333 122 2365
rect 154 2333 190 2365
rect 222 2333 258 2365
rect 290 2333 326 2365
rect 358 2333 394 2365
rect 426 2333 459 2365
rect 21 2319 459 2333
<< psubdiffcont >>
rect 54 35 86 67
rect 122 35 154 67
rect 190 35 222 67
rect 258 35 290 67
rect 326 35 358 67
rect 394 35 426 67
<< nsubdiffcont >>
rect 54 2333 86 2365
rect 122 2333 154 2365
rect 190 2333 222 2365
rect 258 2333 290 2365
rect 326 2333 358 2365
rect 394 2333 426 2365
<< poly >>
rect 89 2158 115 2194
rect 191 2158 217 2194
rect 89 1182 115 1276
rect 191 1182 217 1276
rect 21 1168 115 1182
rect 21 1136 35 1168
rect 67 1136 115 1168
rect 21 1122 115 1136
rect 151 1168 217 1182
rect 151 1136 165 1168
rect 197 1136 217 1168
rect 151 1122 217 1136
rect 89 1028 115 1122
rect 191 1028 217 1122
rect 89 206 115 242
rect 191 206 217 242
<< polycont >>
rect 35 1136 67 1168
rect 165 1136 197 1168
<< metal1 >>
rect 0 2365 480 2400
rect 0 2333 54 2365
rect 86 2333 122 2365
rect 154 2333 190 2365
rect 222 2333 258 2365
rect 290 2333 326 2365
rect 358 2333 394 2365
rect 426 2333 480 2365
rect 0 2144 480 2333
rect 0 2112 35 2144
rect 67 2112 480 2144
rect 30 1168 72 2076
rect 30 1136 35 1168
rect 67 1136 72 1168
rect 30 324 72 1136
rect 160 1168 202 2076
rect 160 1136 165 1168
rect 197 1136 202 1168
rect 160 1051 202 1136
rect 238 2031 280 2076
rect 238 1999 243 2031
rect 275 1999 280 2031
rect 238 1963 280 1999
rect 238 1931 243 1963
rect 275 1931 280 1963
rect 238 1895 280 1931
rect 238 1863 243 1895
rect 275 1863 280 1895
rect 238 1827 280 1863
rect 238 1795 243 1827
rect 275 1795 280 1827
rect 238 1759 280 1795
rect 238 1727 243 1759
rect 275 1727 280 1759
rect 238 1691 280 1727
rect 238 1659 243 1691
rect 275 1659 280 1691
rect 238 1623 280 1659
rect 238 1591 243 1623
rect 275 1591 280 1623
rect 238 1555 280 1591
rect 238 1523 243 1555
rect 275 1523 280 1555
rect 238 1487 280 1523
rect 238 1455 243 1487
rect 275 1455 280 1487
rect 238 1419 280 1455
rect 238 1387 243 1419
rect 275 1387 280 1419
rect 238 1351 280 1387
rect 238 1319 243 1351
rect 275 1319 280 1351
rect 238 1015 280 1319
rect 137 999 280 1015
rect 169 967 280 999
rect 137 931 280 967
rect 169 899 280 931
rect 137 863 280 899
rect 169 831 280 863
rect 137 795 280 831
rect 169 763 280 795
rect 137 727 280 763
rect 169 695 280 727
rect 137 659 280 695
rect 169 627 280 659
rect 137 591 280 627
rect 169 559 280 591
rect 137 523 280 559
rect 169 491 280 523
rect 137 455 280 491
rect 169 423 280 455
rect 137 387 280 423
rect 169 355 280 387
rect 137 324 280 355
rect 0 256 35 288
rect 67 256 243 288
rect 275 256 480 288
rect 0 67 480 256
rect 0 35 54 67
rect 86 35 122 67
rect 154 35 190 67
rect 222 35 258 67
rect 290 35 326 67
rect 358 35 394 67
rect 426 35 480 67
rect 0 0 480 35
<< labels >>
flabel metal1 s 160 1051 202 2076 0 FreeSans 800 0 0 0 i1
port 5 nsew
flabel metal1 s 238 324 280 2076 0 FreeSans 800 0 0 0 nq
port 3 nsew
rlabel metal1 s 30 324 72 2076 4 i0
port 4 nsew
rlabel metal1 s 0 2112 480 2400 4 vdd
port 1 nsew
rlabel metal1 s 0 0 480 288 4 vss
port 2 nsew
flabel comment s 74 52 74 52 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 22701262
string GDS_FILE sg13g2_io.gds
string GDS_START 22697160
<< end >>
