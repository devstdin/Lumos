magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 34 56 350 292
rect -26 -56 410 56
<< nmos >>
rect 128 118 154 266
rect 230 118 256 266
<< pmos >>
rect 128 412 154 636
rect 230 412 256 636
<< ndiff >>
rect 60 245 128 266
rect 60 213 74 245
rect 106 213 128 245
rect 60 166 128 213
rect 60 134 74 166
rect 106 134 128 166
rect 60 118 128 134
rect 154 118 230 266
rect 256 245 324 266
rect 256 213 278 245
rect 310 213 324 245
rect 256 166 324 213
rect 256 134 278 166
rect 310 134 324 166
rect 256 118 324 134
<< pdiff >>
rect 60 622 128 636
rect 60 590 74 622
rect 106 590 128 622
rect 60 540 128 590
rect 60 508 74 540
rect 106 508 128 540
rect 60 458 128 508
rect 60 426 74 458
rect 106 426 128 458
rect 60 412 128 426
rect 154 622 230 636
rect 154 590 176 622
rect 208 590 230 622
rect 154 540 230 590
rect 154 508 176 540
rect 208 508 230 540
rect 154 458 230 508
rect 154 426 176 458
rect 208 426 230 458
rect 154 412 230 426
rect 256 622 324 636
rect 256 590 278 622
rect 310 590 324 622
rect 256 540 324 590
rect 256 508 278 540
rect 310 508 324 540
rect 256 458 324 508
rect 256 426 278 458
rect 310 426 324 458
rect 256 412 324 426
<< ndiffc >>
rect 74 213 106 245
rect 74 134 106 166
rect 278 213 310 245
rect 278 134 310 166
<< pdiffc >>
rect 74 590 106 622
rect 74 508 106 540
rect 74 426 106 458
rect 176 590 208 622
rect 176 508 208 540
rect 176 426 208 458
rect 278 590 310 622
rect 278 508 310 540
rect 278 426 310 458
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 128 636 154 672
rect 230 636 256 672
rect 128 351 154 412
rect 66 337 154 351
rect 66 305 80 337
rect 112 305 154 337
rect 66 291 154 305
rect 128 266 154 291
rect 230 351 256 412
rect 230 337 312 351
rect 230 305 266 337
rect 298 305 312 337
rect 230 291 312 305
rect 230 266 256 291
rect 128 82 154 118
rect 230 82 256 118
<< polycont >>
rect 80 305 112 337
rect 266 305 298 337
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 64 622 116 712
rect 64 590 74 622
rect 106 590 116 622
rect 64 540 116 590
rect 64 508 74 540
rect 106 508 116 540
rect 64 458 116 508
rect 64 426 74 458
rect 106 426 116 458
rect 64 416 116 426
rect 166 622 218 632
rect 166 590 176 622
rect 208 590 218 622
rect 166 540 218 590
rect 166 508 176 540
rect 208 508 218 540
rect 166 458 218 508
rect 166 426 176 458
rect 208 426 218 458
rect 66 337 124 380
rect 66 305 80 337
rect 112 305 124 337
rect 66 294 124 305
rect 64 245 116 255
rect 64 213 74 245
rect 106 213 116 245
rect 64 166 116 213
rect 166 249 218 426
rect 268 622 320 712
rect 268 590 278 622
rect 310 590 320 622
rect 268 540 320 590
rect 268 508 278 540
rect 310 508 320 540
rect 268 458 320 508
rect 268 426 278 458
rect 310 426 320 458
rect 268 416 320 426
rect 254 337 320 380
rect 254 305 266 337
rect 298 305 320 337
rect 254 294 320 305
rect 166 245 320 249
rect 166 213 278 245
rect 310 213 320 245
rect 166 212 320 213
rect 64 134 74 166
rect 106 134 116 166
rect 64 44 116 134
rect 268 166 320 212
rect 268 134 278 166
rect 310 134 320 166
rect 268 124 320 134
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 166 273 218 632 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 254 294 320 380 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 66 294 124 380 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 173970
string GDS_FILE 6_final.gds
string GDS_START 170172
<< end >>
