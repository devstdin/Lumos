magic
tech ihp-sg13g2
timestamp 1757240632
<< error_p >>
rect -23 2765 23 2791
rect 77 2765 123 2791
rect -23 -2791 23 -2765
rect 77 -2791 123 -2765
<< psubdiff >>
rect -115 2876 215 2883
rect -115 2860 -78 2876
rect 178 2860 215 2876
rect -115 2853 215 2860
rect -115 2846 -85 2853
rect -115 -2846 -108 2846
rect -92 -2846 -85 2846
rect 185 2846 215 2853
rect -115 -2853 -85 -2846
rect 185 -2846 192 2846
rect 208 -2846 215 2846
rect 185 -2853 215 -2846
rect -115 -2860 215 -2853
rect -115 -2876 -78 -2860
rect 178 -2876 215 -2860
rect -115 -2883 215 -2876
<< psubdiffcont >>
rect -78 2860 178 2876
rect -108 -2846 -92 2846
rect 192 -2846 208 2846
rect -78 -2876 178 -2860
<< poly >>
rect -25 2786 25 2793
rect -25 2770 -18 2786
rect 18 2770 25 2786
rect -25 2750 25 2770
rect -25 -2770 25 -2750
rect -25 -2786 -18 -2770
rect 18 -2786 25 -2770
rect -25 -2793 25 -2786
rect 75 2786 125 2793
rect 75 2770 82 2786
rect 118 2770 125 2786
rect 75 2750 125 2770
rect 75 -2770 125 -2750
rect 75 -2786 82 -2770
rect 118 -2786 125 -2770
rect 75 -2793 125 -2786
<< polycont >>
rect -18 2770 18 2786
rect -18 -2786 18 -2770
rect 82 2770 118 2786
rect 82 -2786 118 -2770
<< xpolyres >>
rect -25 -2750 25 2750
rect 75 -2750 125 2750
<< metal1 >>
rect -113 2876 213 2881
rect -113 2860 -78 2876
rect 178 2860 213 2876
rect -113 2855 213 2860
rect -113 2846 -87 2855
rect -113 -2846 -108 2846
rect -92 -2846 -87 2846
rect 187 2846 213 2855
rect -113 -2855 -87 -2846
rect 187 -2846 192 2846
rect 208 -2846 213 2846
rect 187 -2855 213 -2846
rect -113 -2860 213 -2855
rect -113 -2876 -78 -2860
rect 178 -2876 213 -2860
rect -113 -2881 213 -2876
<< properties >>
string gencell rhigh
string library sg13g2_devstdin
string parameters w 0.5 l 55 nx 2 dx 0.5 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class resistor endcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
