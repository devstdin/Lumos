magic
tech ihp-sg13g2
magscale 1 2
timestamp 1749416725
<< error_p >>
rect -2510 13390 -2501 13399
rect 2501 13390 2510 13399
rect 2930 13390 2939 13399
rect 7941 13390 7950 13399
rect 8370 13390 8379 13399
rect 13381 13390 13390 13399
rect -2519 13381 -2510 13390
rect 2510 13381 2519 13390
rect -2519 8370 -2510 8379
rect 2510 8370 2519 8379
rect 2921 8370 2930 8379
rect 7950 8370 7959 8379
rect 8361 8370 8370 8379
rect 13390 8370 13399 8379
rect -2510 8361 -2501 8370
rect 2501 8361 2510 8370
rect 2930 8361 2939 8370
rect 7941 8361 7950 8370
rect 8370 8361 8379 8370
rect 13381 8361 13390 8370
rect -2510 7950 -2501 7959
rect 2501 7950 2510 7959
rect 2930 7950 2939 7959
rect 7941 7950 7950 7959
rect 8370 7950 8379 7959
rect 13381 7950 13390 7959
rect -2519 7941 -2510 7950
rect 2510 7941 2519 7950
rect -2519 2930 -2510 2939
rect 2510 2930 2519 2939
rect 2921 2930 2930 2939
rect 7950 2930 7959 2939
rect 8361 2930 8370 2939
rect 13390 2930 13399 2939
rect -2510 2921 -2501 2930
rect 2501 2921 2510 2930
rect 2930 2921 2939 2930
rect 7941 2921 7950 2930
rect 8370 2921 8379 2930
rect 13381 2921 13390 2930
rect -2510 2510 -2501 2519
rect 2501 2510 2510 2519
rect 2930 2510 2939 2519
rect 7941 2510 7950 2519
rect 8370 2510 8379 2519
rect 13381 2510 13390 2519
rect -2519 2501 -2510 2510
rect 2510 2501 2519 2510
rect -2519 -2510 -2510 -2501
rect 2510 -2510 2519 -2501
rect 2921 -2510 2930 -2501
rect 7950 -2510 7959 -2501
rect 8361 -2510 8370 -2501
rect 13390 -2510 13399 -2501
rect -2510 -2519 -2501 -2510
rect 2501 -2519 2510 -2510
rect 2930 -2519 2939 -2510
rect 7941 -2519 7950 -2510
rect 8370 -2519 8379 -2510
rect 13381 -2519 13390 -2510
<< via4 >>
rect -2510 8370 2510 13390
rect 2930 8370 7950 13390
rect 8370 8370 13390 13390
rect -2510 2930 2510 7950
rect 2930 2930 7950 7950
rect 8370 2930 13390 7950
rect -2510 -2510 2510 2510
rect 2930 -2510 7950 2510
rect 8370 -2510 13390 2510
<< metal5 >>
rect -2520 13390 2520 13400
rect -2520 8370 -2510 13390
rect 2510 8370 2520 13390
rect -2520 8360 2520 8370
rect 2920 13390 7960 13400
rect 2920 8370 2930 13390
rect 7950 8370 7960 13390
rect 2920 8360 7960 8370
rect 8360 13390 13400 13400
rect 8360 8370 8370 13390
rect 13390 8370 13400 13390
rect 8360 8360 13400 8370
rect -2520 7950 2520 7960
rect -2520 2930 -2510 7950
rect 2510 2930 2520 7950
rect -2520 2920 2520 2930
rect 2920 7950 7960 7960
rect 2920 2930 2930 7950
rect 7950 2930 7960 7950
rect 2920 2920 7960 2930
rect 8360 7950 13400 7960
rect 8360 2930 8370 7950
rect 13390 2930 13400 7950
rect 8360 2920 13400 2930
rect -2520 2510 2520 2520
rect -2520 -2510 -2510 2510
rect 2510 -2510 2520 2510
rect -2520 -2520 2520 -2510
rect 2920 2510 7960 2520
rect 2920 -2510 2930 2510
rect 7950 -2510 7960 2510
rect 2920 -2520 7960 -2510
rect 8360 2510 13400 2520
rect 8360 -2510 8370 2510
rect 13390 -2510 13400 2510
rect 8360 -2520 13400 -2510
<< mimcap >>
rect -2400 13208 2400 13280
rect -2400 8552 -2328 13208
rect 2328 8552 2400 13208
rect -2400 8480 2400 8552
rect 3040 13208 7840 13280
rect 3040 8552 3112 13208
rect 7768 8552 7840 13208
rect 3040 8480 7840 8552
rect 8480 13208 13280 13280
rect 8480 8552 8552 13208
rect 13208 8552 13280 13208
rect 8480 8480 13280 8552
rect -2400 7768 2400 7840
rect -2400 3112 -2328 7768
rect 2328 3112 2400 7768
rect -2400 3040 2400 3112
rect 3040 7768 7840 7840
rect 3040 3112 3112 7768
rect 7768 3112 7840 7768
rect 3040 3040 7840 3112
rect 8480 7768 13280 7840
rect 8480 3112 8552 7768
rect 13208 3112 13280 7768
rect 8480 3040 13280 3112
rect -2400 2328 2400 2400
rect -2400 -2328 -2328 2328
rect 2328 -2328 2400 2328
rect -2400 -2400 2400 -2328
rect 3040 2328 7840 2400
rect 3040 -2328 3112 2328
rect 7768 -2328 7840 2328
rect 3040 -2400 7840 -2328
rect 8480 2328 13280 2400
rect 8480 -2328 8552 2328
rect 13208 -2328 13280 2328
rect 8480 -2400 13280 -2328
<< mimcapcontact >>
rect -2328 8552 2328 13208
rect 3112 8552 7768 13208
rect 8552 8552 13208 13208
rect -2328 3112 2328 7768
rect 3112 3112 7768 7768
rect 8552 3112 13208 7768
rect -2328 -2328 2328 2328
rect 3112 -2328 7768 2328
rect 8552 -2328 13208 2328
<< properties >>
string gencell cmim
string library sg13g2_devstdin
string parameters w 24 l 24 nx 3 dx 2 ny 3 dy 2 wmin 1.14 lmin 1.14 class capacitor topcc 100 botcc 100
<< end >>
