magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2124 18124 4104
<< nwell >>
rect -124 1788 16124 2104
rect -124 192 192 1788
rect 15808 192 16124 1788
rect -124 -124 16124 192
<< pwell >>
rect 334 1526 15666 1646
rect 334 454 454 1526
rect 2960 1237 3168 1526
rect 5679 454 10321 1526
rect 15546 454 15666 1526
rect 334 334 15666 454
<< hvnmos >>
rect 5799 550 5919 1430
rect 6155 550 6275 1430
rect 6403 550 6523 1430
rect 6759 550 6879 1430
rect 7007 550 7127 1430
rect 7363 550 7483 1430
rect 7611 550 7731 1430
rect 7967 550 8087 1430
rect 8215 550 8335 1430
rect 8571 550 8691 1430
rect 8819 550 8939 1430
rect 9175 550 9295 1430
rect 9423 550 9543 1430
rect 9779 550 9899 1430
rect 10027 550 10147 1430
<< hvndiff >>
rect 5705 1414 5799 1430
rect 5705 1382 5719 1414
rect 5751 1382 5799 1414
rect 5705 1346 5799 1382
rect 5705 1314 5719 1346
rect 5751 1314 5799 1346
rect 5705 1278 5799 1314
rect 5705 1246 5719 1278
rect 5751 1246 5799 1278
rect 5705 1210 5799 1246
rect 5705 1178 5719 1210
rect 5751 1178 5799 1210
rect 5705 1142 5799 1178
rect 5705 1110 5719 1142
rect 5751 1110 5799 1142
rect 5705 1074 5799 1110
rect 5705 1042 5719 1074
rect 5751 1042 5799 1074
rect 5705 1006 5799 1042
rect 5705 974 5719 1006
rect 5751 974 5799 1006
rect 5705 938 5799 974
rect 5705 906 5719 938
rect 5751 906 5799 938
rect 5705 870 5799 906
rect 5705 838 5719 870
rect 5751 838 5799 870
rect 5705 802 5799 838
rect 5705 770 5719 802
rect 5751 770 5799 802
rect 5705 734 5799 770
rect 5705 702 5719 734
rect 5751 702 5799 734
rect 5705 666 5799 702
rect 5705 634 5719 666
rect 5751 634 5799 666
rect 5705 598 5799 634
rect 5705 566 5719 598
rect 5751 566 5799 598
rect 5705 550 5799 566
rect 5919 1414 6155 1430
rect 5919 1382 6021 1414
rect 6053 1382 6155 1414
rect 5919 1346 6155 1382
rect 5919 1314 6021 1346
rect 6053 1314 6155 1346
rect 5919 1278 6155 1314
rect 5919 1246 6021 1278
rect 6053 1246 6155 1278
rect 5919 1210 6155 1246
rect 5919 1178 6021 1210
rect 6053 1178 6155 1210
rect 5919 1142 6155 1178
rect 5919 1110 6021 1142
rect 6053 1110 6155 1142
rect 5919 1074 6155 1110
rect 5919 1042 6021 1074
rect 6053 1042 6155 1074
rect 5919 1006 6155 1042
rect 5919 974 6021 1006
rect 6053 974 6155 1006
rect 5919 938 6155 974
rect 5919 906 6021 938
rect 6053 906 6155 938
rect 5919 870 6155 906
rect 5919 838 6021 870
rect 6053 838 6155 870
rect 5919 802 6155 838
rect 5919 770 6021 802
rect 6053 770 6155 802
rect 5919 734 6155 770
rect 5919 702 6021 734
rect 6053 702 6155 734
rect 5919 666 6155 702
rect 5919 634 6021 666
rect 6053 634 6155 666
rect 5919 598 6155 634
rect 5919 566 6021 598
rect 6053 566 6155 598
rect 5919 550 6155 566
rect 6275 1414 6403 1430
rect 6275 1382 6323 1414
rect 6355 1382 6403 1414
rect 6275 1346 6403 1382
rect 6275 1314 6323 1346
rect 6355 1314 6403 1346
rect 6275 1278 6403 1314
rect 6275 1246 6323 1278
rect 6355 1246 6403 1278
rect 6275 1210 6403 1246
rect 6275 1178 6323 1210
rect 6355 1178 6403 1210
rect 6275 1142 6403 1178
rect 6275 1110 6323 1142
rect 6355 1110 6403 1142
rect 6275 1074 6403 1110
rect 6275 1042 6323 1074
rect 6355 1042 6403 1074
rect 6275 1006 6403 1042
rect 6275 974 6323 1006
rect 6355 974 6403 1006
rect 6275 938 6403 974
rect 6275 906 6323 938
rect 6355 906 6403 938
rect 6275 870 6403 906
rect 6275 838 6323 870
rect 6355 838 6403 870
rect 6275 802 6403 838
rect 6275 770 6323 802
rect 6355 770 6403 802
rect 6275 734 6403 770
rect 6275 702 6323 734
rect 6355 702 6403 734
rect 6275 666 6403 702
rect 6275 634 6323 666
rect 6355 634 6403 666
rect 6275 598 6403 634
rect 6275 566 6323 598
rect 6355 566 6403 598
rect 6275 550 6403 566
rect 6523 1414 6759 1430
rect 6523 1382 6625 1414
rect 6657 1382 6759 1414
rect 6523 1346 6759 1382
rect 6523 1314 6625 1346
rect 6657 1314 6759 1346
rect 6523 1278 6759 1314
rect 6523 1246 6625 1278
rect 6657 1246 6759 1278
rect 6523 1210 6759 1246
rect 6523 1178 6625 1210
rect 6657 1178 6759 1210
rect 6523 1142 6759 1178
rect 6523 1110 6625 1142
rect 6657 1110 6759 1142
rect 6523 1074 6759 1110
rect 6523 1042 6625 1074
rect 6657 1042 6759 1074
rect 6523 1006 6759 1042
rect 6523 974 6625 1006
rect 6657 974 6759 1006
rect 6523 938 6759 974
rect 6523 906 6625 938
rect 6657 906 6759 938
rect 6523 870 6759 906
rect 6523 838 6625 870
rect 6657 838 6759 870
rect 6523 802 6759 838
rect 6523 770 6625 802
rect 6657 770 6759 802
rect 6523 734 6759 770
rect 6523 702 6625 734
rect 6657 702 6759 734
rect 6523 666 6759 702
rect 6523 634 6625 666
rect 6657 634 6759 666
rect 6523 598 6759 634
rect 6523 566 6625 598
rect 6657 566 6759 598
rect 6523 550 6759 566
rect 6879 1414 7007 1430
rect 6879 1382 6927 1414
rect 6959 1382 7007 1414
rect 6879 1346 7007 1382
rect 6879 1314 6927 1346
rect 6959 1314 7007 1346
rect 6879 1278 7007 1314
rect 6879 1246 6927 1278
rect 6959 1246 7007 1278
rect 6879 1210 7007 1246
rect 6879 1178 6927 1210
rect 6959 1178 7007 1210
rect 6879 1142 7007 1178
rect 6879 1110 6927 1142
rect 6959 1110 7007 1142
rect 6879 1074 7007 1110
rect 6879 1042 6927 1074
rect 6959 1042 7007 1074
rect 6879 1006 7007 1042
rect 6879 974 6927 1006
rect 6959 974 7007 1006
rect 6879 938 7007 974
rect 6879 906 6927 938
rect 6959 906 7007 938
rect 6879 870 7007 906
rect 6879 838 6927 870
rect 6959 838 7007 870
rect 6879 802 7007 838
rect 6879 770 6927 802
rect 6959 770 7007 802
rect 6879 734 7007 770
rect 6879 702 6927 734
rect 6959 702 7007 734
rect 6879 666 7007 702
rect 6879 634 6927 666
rect 6959 634 7007 666
rect 6879 598 7007 634
rect 6879 566 6927 598
rect 6959 566 7007 598
rect 6879 550 7007 566
rect 7127 1414 7363 1430
rect 7127 1382 7229 1414
rect 7261 1382 7363 1414
rect 7127 1346 7363 1382
rect 7127 1314 7229 1346
rect 7261 1314 7363 1346
rect 7127 1278 7363 1314
rect 7127 1246 7229 1278
rect 7261 1246 7363 1278
rect 7127 1210 7363 1246
rect 7127 1178 7229 1210
rect 7261 1178 7363 1210
rect 7127 1142 7363 1178
rect 7127 1110 7229 1142
rect 7261 1110 7363 1142
rect 7127 1074 7363 1110
rect 7127 1042 7229 1074
rect 7261 1042 7363 1074
rect 7127 1006 7363 1042
rect 7127 974 7229 1006
rect 7261 974 7363 1006
rect 7127 938 7363 974
rect 7127 906 7229 938
rect 7261 906 7363 938
rect 7127 870 7363 906
rect 7127 838 7229 870
rect 7261 838 7363 870
rect 7127 802 7363 838
rect 7127 770 7229 802
rect 7261 770 7363 802
rect 7127 734 7363 770
rect 7127 702 7229 734
rect 7261 702 7363 734
rect 7127 666 7363 702
rect 7127 634 7229 666
rect 7261 634 7363 666
rect 7127 598 7363 634
rect 7127 566 7229 598
rect 7261 566 7363 598
rect 7127 550 7363 566
rect 7483 1414 7611 1430
rect 7483 1382 7531 1414
rect 7563 1382 7611 1414
rect 7483 1346 7611 1382
rect 7483 1314 7531 1346
rect 7563 1314 7611 1346
rect 7483 1278 7611 1314
rect 7483 1246 7531 1278
rect 7563 1246 7611 1278
rect 7483 1210 7611 1246
rect 7483 1178 7531 1210
rect 7563 1178 7611 1210
rect 7483 1142 7611 1178
rect 7483 1110 7531 1142
rect 7563 1110 7611 1142
rect 7483 1074 7611 1110
rect 7483 1042 7531 1074
rect 7563 1042 7611 1074
rect 7483 1006 7611 1042
rect 7483 974 7531 1006
rect 7563 974 7611 1006
rect 7483 938 7611 974
rect 7483 906 7531 938
rect 7563 906 7611 938
rect 7483 870 7611 906
rect 7483 838 7531 870
rect 7563 838 7611 870
rect 7483 802 7611 838
rect 7483 770 7531 802
rect 7563 770 7611 802
rect 7483 734 7611 770
rect 7483 702 7531 734
rect 7563 702 7611 734
rect 7483 666 7611 702
rect 7483 634 7531 666
rect 7563 634 7611 666
rect 7483 598 7611 634
rect 7483 566 7531 598
rect 7563 566 7611 598
rect 7483 550 7611 566
rect 7731 1414 7967 1430
rect 7731 1382 7833 1414
rect 7865 1382 7967 1414
rect 7731 1346 7967 1382
rect 7731 1314 7833 1346
rect 7865 1314 7967 1346
rect 7731 1278 7967 1314
rect 7731 1246 7833 1278
rect 7865 1246 7967 1278
rect 7731 1210 7967 1246
rect 7731 1178 7833 1210
rect 7865 1178 7967 1210
rect 7731 1142 7967 1178
rect 7731 1110 7833 1142
rect 7865 1110 7967 1142
rect 7731 1074 7967 1110
rect 7731 1042 7833 1074
rect 7865 1042 7967 1074
rect 7731 1006 7967 1042
rect 7731 974 7833 1006
rect 7865 974 7967 1006
rect 7731 938 7967 974
rect 7731 906 7833 938
rect 7865 906 7967 938
rect 7731 870 7967 906
rect 7731 838 7833 870
rect 7865 838 7967 870
rect 7731 802 7967 838
rect 7731 770 7833 802
rect 7865 770 7967 802
rect 7731 734 7967 770
rect 7731 702 7833 734
rect 7865 702 7967 734
rect 7731 666 7967 702
rect 7731 634 7833 666
rect 7865 634 7967 666
rect 7731 598 7967 634
rect 7731 566 7833 598
rect 7865 566 7967 598
rect 7731 550 7967 566
rect 8087 1414 8215 1430
rect 8087 1382 8135 1414
rect 8167 1382 8215 1414
rect 8087 1346 8215 1382
rect 8087 1314 8135 1346
rect 8167 1314 8215 1346
rect 8087 1278 8215 1314
rect 8087 1246 8135 1278
rect 8167 1246 8215 1278
rect 8087 1210 8215 1246
rect 8087 1178 8135 1210
rect 8167 1178 8215 1210
rect 8087 1142 8215 1178
rect 8087 1110 8135 1142
rect 8167 1110 8215 1142
rect 8087 1074 8215 1110
rect 8087 1042 8135 1074
rect 8167 1042 8215 1074
rect 8087 1006 8215 1042
rect 8087 974 8135 1006
rect 8167 974 8215 1006
rect 8087 938 8215 974
rect 8087 906 8135 938
rect 8167 906 8215 938
rect 8087 870 8215 906
rect 8087 838 8135 870
rect 8167 838 8215 870
rect 8087 802 8215 838
rect 8087 770 8135 802
rect 8167 770 8215 802
rect 8087 734 8215 770
rect 8087 702 8135 734
rect 8167 702 8215 734
rect 8087 666 8215 702
rect 8087 634 8135 666
rect 8167 634 8215 666
rect 8087 598 8215 634
rect 8087 566 8135 598
rect 8167 566 8215 598
rect 8087 550 8215 566
rect 8335 1414 8571 1430
rect 8335 1382 8437 1414
rect 8469 1382 8571 1414
rect 8335 1346 8571 1382
rect 8335 1314 8437 1346
rect 8469 1314 8571 1346
rect 8335 1278 8571 1314
rect 8335 1246 8437 1278
rect 8469 1246 8571 1278
rect 8335 1210 8571 1246
rect 8335 1178 8437 1210
rect 8469 1178 8571 1210
rect 8335 1142 8571 1178
rect 8335 1110 8437 1142
rect 8469 1110 8571 1142
rect 8335 1074 8571 1110
rect 8335 1042 8437 1074
rect 8469 1042 8571 1074
rect 8335 1006 8571 1042
rect 8335 974 8437 1006
rect 8469 974 8571 1006
rect 8335 938 8571 974
rect 8335 906 8437 938
rect 8469 906 8571 938
rect 8335 870 8571 906
rect 8335 838 8437 870
rect 8469 838 8571 870
rect 8335 802 8571 838
rect 8335 770 8437 802
rect 8469 770 8571 802
rect 8335 734 8571 770
rect 8335 702 8437 734
rect 8469 702 8571 734
rect 8335 666 8571 702
rect 8335 634 8437 666
rect 8469 634 8571 666
rect 8335 598 8571 634
rect 8335 566 8437 598
rect 8469 566 8571 598
rect 8335 550 8571 566
rect 8691 1414 8819 1430
rect 8691 1382 8739 1414
rect 8771 1382 8819 1414
rect 8691 1346 8819 1382
rect 8691 1314 8739 1346
rect 8771 1314 8819 1346
rect 8691 1278 8819 1314
rect 8691 1246 8739 1278
rect 8771 1246 8819 1278
rect 8691 1210 8819 1246
rect 8691 1178 8739 1210
rect 8771 1178 8819 1210
rect 8691 1142 8819 1178
rect 8691 1110 8739 1142
rect 8771 1110 8819 1142
rect 8691 1074 8819 1110
rect 8691 1042 8739 1074
rect 8771 1042 8819 1074
rect 8691 1006 8819 1042
rect 8691 974 8739 1006
rect 8771 974 8819 1006
rect 8691 938 8819 974
rect 8691 906 8739 938
rect 8771 906 8819 938
rect 8691 870 8819 906
rect 8691 838 8739 870
rect 8771 838 8819 870
rect 8691 802 8819 838
rect 8691 770 8739 802
rect 8771 770 8819 802
rect 8691 734 8819 770
rect 8691 702 8739 734
rect 8771 702 8819 734
rect 8691 666 8819 702
rect 8691 634 8739 666
rect 8771 634 8819 666
rect 8691 598 8819 634
rect 8691 566 8739 598
rect 8771 566 8819 598
rect 8691 550 8819 566
rect 8939 1414 9175 1430
rect 8939 1382 9041 1414
rect 9073 1382 9175 1414
rect 8939 1346 9175 1382
rect 8939 1314 9041 1346
rect 9073 1314 9175 1346
rect 8939 1278 9175 1314
rect 8939 1246 9041 1278
rect 9073 1246 9175 1278
rect 8939 1210 9175 1246
rect 8939 1178 9041 1210
rect 9073 1178 9175 1210
rect 8939 1142 9175 1178
rect 8939 1110 9041 1142
rect 9073 1110 9175 1142
rect 8939 1074 9175 1110
rect 8939 1042 9041 1074
rect 9073 1042 9175 1074
rect 8939 1006 9175 1042
rect 8939 974 9041 1006
rect 9073 974 9175 1006
rect 8939 938 9175 974
rect 8939 906 9041 938
rect 9073 906 9175 938
rect 8939 870 9175 906
rect 8939 838 9041 870
rect 9073 838 9175 870
rect 8939 802 9175 838
rect 8939 770 9041 802
rect 9073 770 9175 802
rect 8939 734 9175 770
rect 8939 702 9041 734
rect 9073 702 9175 734
rect 8939 666 9175 702
rect 8939 634 9041 666
rect 9073 634 9175 666
rect 8939 598 9175 634
rect 8939 566 9041 598
rect 9073 566 9175 598
rect 8939 550 9175 566
rect 9295 1414 9423 1430
rect 9295 1382 9343 1414
rect 9375 1382 9423 1414
rect 9295 1346 9423 1382
rect 9295 1314 9343 1346
rect 9375 1314 9423 1346
rect 9295 1278 9423 1314
rect 9295 1246 9343 1278
rect 9375 1246 9423 1278
rect 9295 1210 9423 1246
rect 9295 1178 9343 1210
rect 9375 1178 9423 1210
rect 9295 1142 9423 1178
rect 9295 1110 9343 1142
rect 9375 1110 9423 1142
rect 9295 1074 9423 1110
rect 9295 1042 9343 1074
rect 9375 1042 9423 1074
rect 9295 1006 9423 1042
rect 9295 974 9343 1006
rect 9375 974 9423 1006
rect 9295 938 9423 974
rect 9295 906 9343 938
rect 9375 906 9423 938
rect 9295 870 9423 906
rect 9295 838 9343 870
rect 9375 838 9423 870
rect 9295 802 9423 838
rect 9295 770 9343 802
rect 9375 770 9423 802
rect 9295 734 9423 770
rect 9295 702 9343 734
rect 9375 702 9423 734
rect 9295 666 9423 702
rect 9295 634 9343 666
rect 9375 634 9423 666
rect 9295 598 9423 634
rect 9295 566 9343 598
rect 9375 566 9423 598
rect 9295 550 9423 566
rect 9543 1414 9779 1430
rect 9543 1382 9645 1414
rect 9677 1382 9779 1414
rect 9543 1346 9779 1382
rect 9543 1314 9645 1346
rect 9677 1314 9779 1346
rect 9543 1278 9779 1314
rect 9543 1246 9645 1278
rect 9677 1246 9779 1278
rect 9543 1210 9779 1246
rect 9543 1178 9645 1210
rect 9677 1178 9779 1210
rect 9543 1142 9779 1178
rect 9543 1110 9645 1142
rect 9677 1110 9779 1142
rect 9543 1074 9779 1110
rect 9543 1042 9645 1074
rect 9677 1042 9779 1074
rect 9543 1006 9779 1042
rect 9543 974 9645 1006
rect 9677 974 9779 1006
rect 9543 938 9779 974
rect 9543 906 9645 938
rect 9677 906 9779 938
rect 9543 870 9779 906
rect 9543 838 9645 870
rect 9677 838 9779 870
rect 9543 802 9779 838
rect 9543 770 9645 802
rect 9677 770 9779 802
rect 9543 734 9779 770
rect 9543 702 9645 734
rect 9677 702 9779 734
rect 9543 666 9779 702
rect 9543 634 9645 666
rect 9677 634 9779 666
rect 9543 598 9779 634
rect 9543 566 9645 598
rect 9677 566 9779 598
rect 9543 550 9779 566
rect 9899 1414 10027 1430
rect 9899 1382 9947 1414
rect 9979 1382 10027 1414
rect 9899 1346 10027 1382
rect 9899 1314 9947 1346
rect 9979 1314 10027 1346
rect 9899 1278 10027 1314
rect 9899 1246 9947 1278
rect 9979 1246 10027 1278
rect 9899 1210 10027 1246
rect 9899 1178 9947 1210
rect 9979 1178 10027 1210
rect 9899 1142 10027 1178
rect 9899 1110 9947 1142
rect 9979 1110 10027 1142
rect 9899 1074 10027 1110
rect 9899 1042 9947 1074
rect 9979 1042 10027 1074
rect 9899 1006 10027 1042
rect 9899 974 9947 1006
rect 9979 974 10027 1006
rect 9899 938 10027 974
rect 9899 906 9947 938
rect 9979 906 10027 938
rect 9899 870 10027 906
rect 9899 838 9947 870
rect 9979 838 10027 870
rect 9899 802 10027 838
rect 9899 770 9947 802
rect 9979 770 10027 802
rect 9899 734 10027 770
rect 9899 702 9947 734
rect 9979 702 10027 734
rect 9899 666 10027 702
rect 9899 634 9947 666
rect 9979 634 10027 666
rect 9899 598 10027 634
rect 9899 566 9947 598
rect 9979 566 10027 598
rect 9899 550 10027 566
rect 10147 1414 10295 1430
rect 10147 1382 10249 1414
rect 10281 1382 10295 1414
rect 10147 1346 10295 1382
rect 10147 1314 10249 1346
rect 10281 1314 10295 1346
rect 10147 1278 10295 1314
rect 10147 1246 10249 1278
rect 10281 1246 10295 1278
rect 10147 1210 10295 1246
rect 10147 1178 10249 1210
rect 10281 1178 10295 1210
rect 10147 1142 10295 1178
rect 10147 1110 10249 1142
rect 10281 1110 10295 1142
rect 10147 1074 10295 1110
rect 10147 1042 10249 1074
rect 10281 1042 10295 1074
rect 10147 1006 10295 1042
rect 10147 974 10249 1006
rect 10281 974 10295 1006
rect 10147 938 10295 974
rect 10147 906 10249 938
rect 10281 906 10295 938
rect 10147 870 10295 906
rect 10147 838 10249 870
rect 10281 838 10295 870
rect 10147 802 10295 838
rect 10147 770 10249 802
rect 10281 770 10295 802
rect 10147 734 10295 770
rect 10147 702 10249 734
rect 10281 702 10295 734
rect 10147 666 10295 702
rect 10147 634 10249 666
rect 10281 634 10295 666
rect 10147 598 10295 634
rect 10147 566 10249 598
rect 10281 566 10295 598
rect 10147 550 10295 566
<< hvndiffc >>
rect 5719 1382 5751 1414
rect 5719 1314 5751 1346
rect 5719 1246 5751 1278
rect 5719 1178 5751 1210
rect 5719 1110 5751 1142
rect 5719 1042 5751 1074
rect 5719 974 5751 1006
rect 5719 906 5751 938
rect 5719 838 5751 870
rect 5719 770 5751 802
rect 5719 702 5751 734
rect 5719 634 5751 666
rect 5719 566 5751 598
rect 6021 1382 6053 1414
rect 6021 1314 6053 1346
rect 6021 1246 6053 1278
rect 6021 1178 6053 1210
rect 6021 1110 6053 1142
rect 6021 1042 6053 1074
rect 6021 974 6053 1006
rect 6021 906 6053 938
rect 6021 838 6053 870
rect 6021 770 6053 802
rect 6021 702 6053 734
rect 6021 634 6053 666
rect 6021 566 6053 598
rect 6323 1382 6355 1414
rect 6323 1314 6355 1346
rect 6323 1246 6355 1278
rect 6323 1178 6355 1210
rect 6323 1110 6355 1142
rect 6323 1042 6355 1074
rect 6323 974 6355 1006
rect 6323 906 6355 938
rect 6323 838 6355 870
rect 6323 770 6355 802
rect 6323 702 6355 734
rect 6323 634 6355 666
rect 6323 566 6355 598
rect 6625 1382 6657 1414
rect 6625 1314 6657 1346
rect 6625 1246 6657 1278
rect 6625 1178 6657 1210
rect 6625 1110 6657 1142
rect 6625 1042 6657 1074
rect 6625 974 6657 1006
rect 6625 906 6657 938
rect 6625 838 6657 870
rect 6625 770 6657 802
rect 6625 702 6657 734
rect 6625 634 6657 666
rect 6625 566 6657 598
rect 6927 1382 6959 1414
rect 6927 1314 6959 1346
rect 6927 1246 6959 1278
rect 6927 1178 6959 1210
rect 6927 1110 6959 1142
rect 6927 1042 6959 1074
rect 6927 974 6959 1006
rect 6927 906 6959 938
rect 6927 838 6959 870
rect 6927 770 6959 802
rect 6927 702 6959 734
rect 6927 634 6959 666
rect 6927 566 6959 598
rect 7229 1382 7261 1414
rect 7229 1314 7261 1346
rect 7229 1246 7261 1278
rect 7229 1178 7261 1210
rect 7229 1110 7261 1142
rect 7229 1042 7261 1074
rect 7229 974 7261 1006
rect 7229 906 7261 938
rect 7229 838 7261 870
rect 7229 770 7261 802
rect 7229 702 7261 734
rect 7229 634 7261 666
rect 7229 566 7261 598
rect 7531 1382 7563 1414
rect 7531 1314 7563 1346
rect 7531 1246 7563 1278
rect 7531 1178 7563 1210
rect 7531 1110 7563 1142
rect 7531 1042 7563 1074
rect 7531 974 7563 1006
rect 7531 906 7563 938
rect 7531 838 7563 870
rect 7531 770 7563 802
rect 7531 702 7563 734
rect 7531 634 7563 666
rect 7531 566 7563 598
rect 7833 1382 7865 1414
rect 7833 1314 7865 1346
rect 7833 1246 7865 1278
rect 7833 1178 7865 1210
rect 7833 1110 7865 1142
rect 7833 1042 7865 1074
rect 7833 974 7865 1006
rect 7833 906 7865 938
rect 7833 838 7865 870
rect 7833 770 7865 802
rect 7833 702 7865 734
rect 7833 634 7865 666
rect 7833 566 7865 598
rect 8135 1382 8167 1414
rect 8135 1314 8167 1346
rect 8135 1246 8167 1278
rect 8135 1178 8167 1210
rect 8135 1110 8167 1142
rect 8135 1042 8167 1074
rect 8135 974 8167 1006
rect 8135 906 8167 938
rect 8135 838 8167 870
rect 8135 770 8167 802
rect 8135 702 8167 734
rect 8135 634 8167 666
rect 8135 566 8167 598
rect 8437 1382 8469 1414
rect 8437 1314 8469 1346
rect 8437 1246 8469 1278
rect 8437 1178 8469 1210
rect 8437 1110 8469 1142
rect 8437 1042 8469 1074
rect 8437 974 8469 1006
rect 8437 906 8469 938
rect 8437 838 8469 870
rect 8437 770 8469 802
rect 8437 702 8469 734
rect 8437 634 8469 666
rect 8437 566 8469 598
rect 8739 1382 8771 1414
rect 8739 1314 8771 1346
rect 8739 1246 8771 1278
rect 8739 1178 8771 1210
rect 8739 1110 8771 1142
rect 8739 1042 8771 1074
rect 8739 974 8771 1006
rect 8739 906 8771 938
rect 8739 838 8771 870
rect 8739 770 8771 802
rect 8739 702 8771 734
rect 8739 634 8771 666
rect 8739 566 8771 598
rect 9041 1382 9073 1414
rect 9041 1314 9073 1346
rect 9041 1246 9073 1278
rect 9041 1178 9073 1210
rect 9041 1110 9073 1142
rect 9041 1042 9073 1074
rect 9041 974 9073 1006
rect 9041 906 9073 938
rect 9041 838 9073 870
rect 9041 770 9073 802
rect 9041 702 9073 734
rect 9041 634 9073 666
rect 9041 566 9073 598
rect 9343 1382 9375 1414
rect 9343 1314 9375 1346
rect 9343 1246 9375 1278
rect 9343 1178 9375 1210
rect 9343 1110 9375 1142
rect 9343 1042 9375 1074
rect 9343 974 9375 1006
rect 9343 906 9375 938
rect 9343 838 9375 870
rect 9343 770 9375 802
rect 9343 702 9375 734
rect 9343 634 9375 666
rect 9343 566 9375 598
rect 9645 1382 9677 1414
rect 9645 1314 9677 1346
rect 9645 1246 9677 1278
rect 9645 1178 9677 1210
rect 9645 1110 9677 1142
rect 9645 1042 9677 1074
rect 9645 974 9677 1006
rect 9645 906 9677 938
rect 9645 838 9677 870
rect 9645 770 9677 802
rect 9645 702 9677 734
rect 9645 634 9677 666
rect 9645 566 9677 598
rect 9947 1382 9979 1414
rect 9947 1314 9979 1346
rect 9947 1246 9979 1278
rect 9947 1178 9979 1210
rect 9947 1110 9979 1142
rect 9947 1042 9979 1074
rect 9947 974 9979 1006
rect 9947 906 9979 938
rect 9947 838 9979 870
rect 9947 770 9979 802
rect 9947 702 9979 734
rect 9947 634 9979 666
rect 9947 566 9979 598
rect 10249 1382 10281 1414
rect 10249 1314 10281 1346
rect 10249 1246 10281 1278
rect 10249 1178 10281 1210
rect 10249 1110 10281 1142
rect 10249 1042 10281 1074
rect 10249 974 10281 1006
rect 10249 906 10281 938
rect 10249 838 10281 870
rect 10249 770 10281 802
rect 10249 702 10281 734
rect 10249 634 10281 666
rect 10249 566 10281 598
<< psubdiff >>
rect 360 1602 15640 1620
rect 360 1570 402 1602
rect 434 1570 470 1602
rect 502 1570 538 1602
rect 570 1570 606 1602
rect 638 1570 674 1602
rect 706 1570 742 1602
rect 774 1570 810 1602
rect 842 1570 878 1602
rect 910 1570 946 1602
rect 978 1570 1014 1602
rect 1046 1570 1082 1602
rect 1114 1570 1150 1602
rect 1182 1570 1218 1602
rect 1250 1570 1286 1602
rect 1318 1570 1354 1602
rect 1386 1570 1422 1602
rect 1454 1570 1490 1602
rect 1522 1570 1558 1602
rect 1590 1570 1626 1602
rect 1658 1570 1694 1602
rect 1726 1570 1762 1602
rect 1794 1570 1830 1602
rect 1862 1570 1898 1602
rect 1930 1570 1966 1602
rect 1998 1570 2034 1602
rect 2066 1570 2102 1602
rect 2134 1570 2170 1602
rect 2202 1570 2238 1602
rect 2270 1570 2306 1602
rect 2338 1570 2374 1602
rect 2406 1570 2442 1602
rect 2474 1570 2510 1602
rect 2542 1570 2578 1602
rect 2610 1570 2646 1602
rect 2678 1570 2714 1602
rect 2746 1570 2782 1602
rect 2814 1570 2850 1602
rect 2882 1570 2918 1602
rect 2950 1570 2986 1602
rect 3018 1570 3054 1602
rect 3086 1570 3122 1602
rect 3154 1570 3190 1602
rect 3222 1570 3258 1602
rect 3290 1570 3326 1602
rect 3358 1570 3394 1602
rect 3426 1570 3462 1602
rect 3494 1570 3530 1602
rect 3562 1570 3598 1602
rect 3630 1570 3666 1602
rect 3698 1570 3734 1602
rect 3766 1570 3802 1602
rect 3834 1570 3870 1602
rect 3902 1570 3938 1602
rect 3970 1570 4006 1602
rect 4038 1570 4074 1602
rect 4106 1570 4142 1602
rect 4174 1570 4210 1602
rect 4242 1570 4278 1602
rect 4310 1570 4346 1602
rect 4378 1570 4414 1602
rect 4446 1570 4482 1602
rect 4514 1570 4550 1602
rect 4582 1570 4618 1602
rect 4650 1570 4686 1602
rect 4718 1570 4754 1602
rect 4786 1570 4822 1602
rect 4854 1570 4890 1602
rect 4922 1570 4958 1602
rect 4990 1570 5026 1602
rect 5058 1570 5094 1602
rect 5126 1570 5162 1602
rect 5194 1570 5230 1602
rect 5262 1570 5298 1602
rect 5330 1570 5366 1602
rect 5398 1570 5434 1602
rect 5466 1570 5502 1602
rect 5534 1570 5570 1602
rect 5602 1570 5638 1602
rect 5670 1570 5706 1602
rect 5738 1570 5774 1602
rect 5806 1570 5842 1602
rect 5874 1570 5910 1602
rect 5942 1570 5978 1602
rect 6010 1570 6046 1602
rect 6078 1570 6114 1602
rect 6146 1570 6182 1602
rect 6214 1570 6250 1602
rect 6282 1570 6318 1602
rect 6350 1570 6386 1602
rect 6418 1570 6454 1602
rect 6486 1570 6522 1602
rect 6554 1570 6590 1602
rect 6622 1570 6658 1602
rect 6690 1570 6726 1602
rect 6758 1570 6794 1602
rect 6826 1570 6862 1602
rect 6894 1570 6930 1602
rect 6962 1570 6998 1602
rect 7030 1570 7066 1602
rect 7098 1570 7134 1602
rect 7166 1570 7202 1602
rect 7234 1570 7270 1602
rect 7302 1570 7338 1602
rect 7370 1570 7406 1602
rect 7438 1570 7474 1602
rect 7506 1570 7542 1602
rect 7574 1570 7610 1602
rect 7642 1570 7678 1602
rect 7710 1570 7746 1602
rect 7778 1570 7814 1602
rect 7846 1570 7882 1602
rect 7914 1570 7950 1602
rect 7982 1570 8018 1602
rect 8050 1570 8086 1602
rect 8118 1570 8154 1602
rect 8186 1570 8222 1602
rect 8254 1570 8290 1602
rect 8322 1570 8358 1602
rect 8390 1570 8426 1602
rect 8458 1570 8494 1602
rect 8526 1570 8562 1602
rect 8594 1570 8630 1602
rect 8662 1570 8698 1602
rect 8730 1570 8766 1602
rect 8798 1570 8834 1602
rect 8866 1570 8902 1602
rect 8934 1570 8970 1602
rect 9002 1570 9038 1602
rect 9070 1570 9106 1602
rect 9138 1570 9174 1602
rect 9206 1570 9242 1602
rect 9274 1570 9310 1602
rect 9342 1570 9378 1602
rect 9410 1570 9446 1602
rect 9478 1570 9514 1602
rect 9546 1570 9582 1602
rect 9614 1570 9650 1602
rect 9682 1570 9718 1602
rect 9750 1570 9786 1602
rect 9818 1570 9854 1602
rect 9886 1570 9922 1602
rect 9954 1570 9990 1602
rect 10022 1570 10058 1602
rect 10090 1570 10126 1602
rect 10158 1570 10194 1602
rect 10226 1570 10262 1602
rect 10294 1570 10330 1602
rect 10362 1570 10398 1602
rect 10430 1570 10466 1602
rect 10498 1570 10534 1602
rect 10566 1570 10602 1602
rect 10634 1570 10670 1602
rect 10702 1570 10738 1602
rect 10770 1570 10806 1602
rect 10838 1570 10874 1602
rect 10906 1570 10942 1602
rect 10974 1570 11010 1602
rect 11042 1570 11078 1602
rect 11110 1570 11146 1602
rect 11178 1570 11214 1602
rect 11246 1570 11282 1602
rect 11314 1570 11350 1602
rect 11382 1570 11418 1602
rect 11450 1570 11486 1602
rect 11518 1570 11554 1602
rect 11586 1570 11622 1602
rect 11654 1570 11690 1602
rect 11722 1570 11758 1602
rect 11790 1570 11826 1602
rect 11858 1570 11894 1602
rect 11926 1570 11962 1602
rect 11994 1570 12030 1602
rect 12062 1570 12098 1602
rect 12130 1570 12166 1602
rect 12198 1570 12234 1602
rect 12266 1570 12302 1602
rect 12334 1570 12370 1602
rect 12402 1570 12438 1602
rect 12470 1570 12506 1602
rect 12538 1570 12574 1602
rect 12606 1570 12642 1602
rect 12674 1570 12710 1602
rect 12742 1570 12778 1602
rect 12810 1570 12846 1602
rect 12878 1570 12914 1602
rect 12946 1570 12982 1602
rect 13014 1570 13050 1602
rect 13082 1570 13118 1602
rect 13150 1570 13186 1602
rect 13218 1570 13254 1602
rect 13286 1570 13322 1602
rect 13354 1570 13390 1602
rect 13422 1570 13458 1602
rect 13490 1570 13526 1602
rect 13558 1570 13594 1602
rect 13626 1570 13662 1602
rect 13694 1570 13730 1602
rect 13762 1570 13798 1602
rect 13830 1570 13866 1602
rect 13898 1570 13934 1602
rect 13966 1570 14002 1602
rect 14034 1570 14070 1602
rect 14102 1570 14138 1602
rect 14170 1570 14206 1602
rect 14238 1570 14274 1602
rect 14306 1570 14342 1602
rect 14374 1570 14410 1602
rect 14442 1570 14478 1602
rect 14510 1570 14546 1602
rect 14578 1570 14614 1602
rect 14646 1570 14682 1602
rect 14714 1570 14750 1602
rect 14782 1570 14818 1602
rect 14850 1570 14886 1602
rect 14918 1570 14954 1602
rect 14986 1570 15022 1602
rect 15054 1570 15090 1602
rect 15122 1570 15158 1602
rect 15190 1570 15226 1602
rect 15258 1570 15294 1602
rect 15326 1570 15362 1602
rect 15394 1570 15430 1602
rect 15462 1570 15498 1602
rect 15530 1570 15566 1602
rect 15598 1570 15640 1602
rect 360 1552 15640 1570
rect 360 1516 428 1552
rect 360 1484 378 1516
rect 410 1484 428 1516
rect 15572 1516 15640 1552
rect 360 1448 428 1484
rect 360 1416 378 1448
rect 410 1416 428 1448
rect 15572 1484 15590 1516
rect 15622 1484 15640 1516
rect 15572 1448 15640 1484
rect 360 1380 428 1416
rect 360 1348 378 1380
rect 410 1348 428 1380
rect 360 1312 428 1348
rect 360 1280 378 1312
rect 410 1280 428 1312
rect 360 1244 428 1280
rect 360 1212 378 1244
rect 410 1212 428 1244
rect 360 1176 428 1212
rect 360 1144 378 1176
rect 410 1144 428 1176
rect 360 1108 428 1144
rect 360 1076 378 1108
rect 410 1076 428 1108
rect 360 1040 428 1076
rect 360 1008 378 1040
rect 410 1008 428 1040
rect 360 972 428 1008
rect 360 940 378 972
rect 410 940 428 972
rect 360 904 428 940
rect 360 872 378 904
rect 410 872 428 904
rect 360 836 428 872
rect 360 804 378 836
rect 410 804 428 836
rect 360 768 428 804
rect 360 736 378 768
rect 410 736 428 768
rect 360 700 428 736
rect 360 668 378 700
rect 410 668 428 700
rect 360 632 428 668
rect 360 600 378 632
rect 410 600 428 632
rect 360 564 428 600
rect 360 532 378 564
rect 410 532 428 564
rect 15572 1416 15590 1448
rect 15622 1416 15640 1448
rect 15572 1380 15640 1416
rect 15572 1348 15590 1380
rect 15622 1348 15640 1380
rect 15572 1312 15640 1348
rect 15572 1280 15590 1312
rect 15622 1280 15640 1312
rect 15572 1244 15640 1280
rect 15572 1212 15590 1244
rect 15622 1212 15640 1244
rect 15572 1176 15640 1212
rect 15572 1144 15590 1176
rect 15622 1144 15640 1176
rect 15572 1108 15640 1144
rect 15572 1076 15590 1108
rect 15622 1076 15640 1108
rect 15572 1040 15640 1076
rect 15572 1008 15590 1040
rect 15622 1008 15640 1040
rect 15572 972 15640 1008
rect 15572 940 15590 972
rect 15622 940 15640 972
rect 15572 904 15640 940
rect 15572 872 15590 904
rect 15622 872 15640 904
rect 15572 836 15640 872
rect 15572 804 15590 836
rect 15622 804 15640 836
rect 15572 768 15640 804
rect 15572 736 15590 768
rect 15622 736 15640 768
rect 15572 700 15640 736
rect 15572 668 15590 700
rect 15622 668 15640 700
rect 15572 632 15640 668
rect 15572 600 15590 632
rect 15622 600 15640 632
rect 15572 564 15640 600
rect 360 496 428 532
rect 360 464 378 496
rect 410 464 428 496
rect 15572 532 15590 564
rect 15622 532 15640 564
rect 15572 496 15640 532
rect 360 428 428 464
rect 15572 464 15590 496
rect 15622 464 15640 496
rect 15572 428 15640 464
rect 360 410 15640 428
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 360 15640 378
<< nsubdiff >>
rect 0 1962 16000 1980
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 15932 360 16000 396
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< psubdiffcont >>
rect 402 1570 434 1602
rect 470 1570 502 1602
rect 538 1570 570 1602
rect 606 1570 638 1602
rect 674 1570 706 1602
rect 742 1570 774 1602
rect 810 1570 842 1602
rect 878 1570 910 1602
rect 946 1570 978 1602
rect 1014 1570 1046 1602
rect 1082 1570 1114 1602
rect 1150 1570 1182 1602
rect 1218 1570 1250 1602
rect 1286 1570 1318 1602
rect 1354 1570 1386 1602
rect 1422 1570 1454 1602
rect 1490 1570 1522 1602
rect 1558 1570 1590 1602
rect 1626 1570 1658 1602
rect 1694 1570 1726 1602
rect 1762 1570 1794 1602
rect 1830 1570 1862 1602
rect 1898 1570 1930 1602
rect 1966 1570 1998 1602
rect 2034 1570 2066 1602
rect 2102 1570 2134 1602
rect 2170 1570 2202 1602
rect 2238 1570 2270 1602
rect 2306 1570 2338 1602
rect 2374 1570 2406 1602
rect 2442 1570 2474 1602
rect 2510 1570 2542 1602
rect 2578 1570 2610 1602
rect 2646 1570 2678 1602
rect 2714 1570 2746 1602
rect 2782 1570 2814 1602
rect 2850 1570 2882 1602
rect 2918 1570 2950 1602
rect 2986 1570 3018 1602
rect 3054 1570 3086 1602
rect 3122 1570 3154 1602
rect 3190 1570 3222 1602
rect 3258 1570 3290 1602
rect 3326 1570 3358 1602
rect 3394 1570 3426 1602
rect 3462 1570 3494 1602
rect 3530 1570 3562 1602
rect 3598 1570 3630 1602
rect 3666 1570 3698 1602
rect 3734 1570 3766 1602
rect 3802 1570 3834 1602
rect 3870 1570 3902 1602
rect 3938 1570 3970 1602
rect 4006 1570 4038 1602
rect 4074 1570 4106 1602
rect 4142 1570 4174 1602
rect 4210 1570 4242 1602
rect 4278 1570 4310 1602
rect 4346 1570 4378 1602
rect 4414 1570 4446 1602
rect 4482 1570 4514 1602
rect 4550 1570 4582 1602
rect 4618 1570 4650 1602
rect 4686 1570 4718 1602
rect 4754 1570 4786 1602
rect 4822 1570 4854 1602
rect 4890 1570 4922 1602
rect 4958 1570 4990 1602
rect 5026 1570 5058 1602
rect 5094 1570 5126 1602
rect 5162 1570 5194 1602
rect 5230 1570 5262 1602
rect 5298 1570 5330 1602
rect 5366 1570 5398 1602
rect 5434 1570 5466 1602
rect 5502 1570 5534 1602
rect 5570 1570 5602 1602
rect 5638 1570 5670 1602
rect 5706 1570 5738 1602
rect 5774 1570 5806 1602
rect 5842 1570 5874 1602
rect 5910 1570 5942 1602
rect 5978 1570 6010 1602
rect 6046 1570 6078 1602
rect 6114 1570 6146 1602
rect 6182 1570 6214 1602
rect 6250 1570 6282 1602
rect 6318 1570 6350 1602
rect 6386 1570 6418 1602
rect 6454 1570 6486 1602
rect 6522 1570 6554 1602
rect 6590 1570 6622 1602
rect 6658 1570 6690 1602
rect 6726 1570 6758 1602
rect 6794 1570 6826 1602
rect 6862 1570 6894 1602
rect 6930 1570 6962 1602
rect 6998 1570 7030 1602
rect 7066 1570 7098 1602
rect 7134 1570 7166 1602
rect 7202 1570 7234 1602
rect 7270 1570 7302 1602
rect 7338 1570 7370 1602
rect 7406 1570 7438 1602
rect 7474 1570 7506 1602
rect 7542 1570 7574 1602
rect 7610 1570 7642 1602
rect 7678 1570 7710 1602
rect 7746 1570 7778 1602
rect 7814 1570 7846 1602
rect 7882 1570 7914 1602
rect 7950 1570 7982 1602
rect 8018 1570 8050 1602
rect 8086 1570 8118 1602
rect 8154 1570 8186 1602
rect 8222 1570 8254 1602
rect 8290 1570 8322 1602
rect 8358 1570 8390 1602
rect 8426 1570 8458 1602
rect 8494 1570 8526 1602
rect 8562 1570 8594 1602
rect 8630 1570 8662 1602
rect 8698 1570 8730 1602
rect 8766 1570 8798 1602
rect 8834 1570 8866 1602
rect 8902 1570 8934 1602
rect 8970 1570 9002 1602
rect 9038 1570 9070 1602
rect 9106 1570 9138 1602
rect 9174 1570 9206 1602
rect 9242 1570 9274 1602
rect 9310 1570 9342 1602
rect 9378 1570 9410 1602
rect 9446 1570 9478 1602
rect 9514 1570 9546 1602
rect 9582 1570 9614 1602
rect 9650 1570 9682 1602
rect 9718 1570 9750 1602
rect 9786 1570 9818 1602
rect 9854 1570 9886 1602
rect 9922 1570 9954 1602
rect 9990 1570 10022 1602
rect 10058 1570 10090 1602
rect 10126 1570 10158 1602
rect 10194 1570 10226 1602
rect 10262 1570 10294 1602
rect 10330 1570 10362 1602
rect 10398 1570 10430 1602
rect 10466 1570 10498 1602
rect 10534 1570 10566 1602
rect 10602 1570 10634 1602
rect 10670 1570 10702 1602
rect 10738 1570 10770 1602
rect 10806 1570 10838 1602
rect 10874 1570 10906 1602
rect 10942 1570 10974 1602
rect 11010 1570 11042 1602
rect 11078 1570 11110 1602
rect 11146 1570 11178 1602
rect 11214 1570 11246 1602
rect 11282 1570 11314 1602
rect 11350 1570 11382 1602
rect 11418 1570 11450 1602
rect 11486 1570 11518 1602
rect 11554 1570 11586 1602
rect 11622 1570 11654 1602
rect 11690 1570 11722 1602
rect 11758 1570 11790 1602
rect 11826 1570 11858 1602
rect 11894 1570 11926 1602
rect 11962 1570 11994 1602
rect 12030 1570 12062 1602
rect 12098 1570 12130 1602
rect 12166 1570 12198 1602
rect 12234 1570 12266 1602
rect 12302 1570 12334 1602
rect 12370 1570 12402 1602
rect 12438 1570 12470 1602
rect 12506 1570 12538 1602
rect 12574 1570 12606 1602
rect 12642 1570 12674 1602
rect 12710 1570 12742 1602
rect 12778 1570 12810 1602
rect 12846 1570 12878 1602
rect 12914 1570 12946 1602
rect 12982 1570 13014 1602
rect 13050 1570 13082 1602
rect 13118 1570 13150 1602
rect 13186 1570 13218 1602
rect 13254 1570 13286 1602
rect 13322 1570 13354 1602
rect 13390 1570 13422 1602
rect 13458 1570 13490 1602
rect 13526 1570 13558 1602
rect 13594 1570 13626 1602
rect 13662 1570 13694 1602
rect 13730 1570 13762 1602
rect 13798 1570 13830 1602
rect 13866 1570 13898 1602
rect 13934 1570 13966 1602
rect 14002 1570 14034 1602
rect 14070 1570 14102 1602
rect 14138 1570 14170 1602
rect 14206 1570 14238 1602
rect 14274 1570 14306 1602
rect 14342 1570 14374 1602
rect 14410 1570 14442 1602
rect 14478 1570 14510 1602
rect 14546 1570 14578 1602
rect 14614 1570 14646 1602
rect 14682 1570 14714 1602
rect 14750 1570 14782 1602
rect 14818 1570 14850 1602
rect 14886 1570 14918 1602
rect 14954 1570 14986 1602
rect 15022 1570 15054 1602
rect 15090 1570 15122 1602
rect 15158 1570 15190 1602
rect 15226 1570 15258 1602
rect 15294 1570 15326 1602
rect 15362 1570 15394 1602
rect 15430 1570 15462 1602
rect 15498 1570 15530 1602
rect 15566 1570 15598 1602
rect 378 1484 410 1516
rect 378 1416 410 1448
rect 15590 1484 15622 1516
rect 378 1348 410 1380
rect 378 1280 410 1312
rect 378 1212 410 1244
rect 378 1144 410 1176
rect 378 1076 410 1108
rect 378 1008 410 1040
rect 378 940 410 972
rect 378 872 410 904
rect 378 804 410 836
rect 378 736 410 768
rect 378 668 410 700
rect 378 600 410 632
rect 378 532 410 564
rect 15590 1416 15622 1448
rect 15590 1348 15622 1380
rect 15590 1280 15622 1312
rect 15590 1212 15622 1244
rect 15590 1144 15622 1176
rect 15590 1076 15622 1108
rect 15590 1008 15622 1040
rect 15590 940 15622 972
rect 15590 872 15622 904
rect 15590 804 15622 836
rect 15590 736 15622 768
rect 15590 668 15622 700
rect 15590 600 15622 632
rect 378 464 410 496
rect 15590 532 15622 564
rect 15590 464 15622 496
rect 402 378 434 410
rect 470 378 502 410
rect 538 378 570 410
rect 606 378 638 410
rect 674 378 706 410
rect 742 378 774 410
rect 810 378 842 410
rect 878 378 910 410
rect 946 378 978 410
rect 1014 378 1046 410
rect 1082 378 1114 410
rect 1150 378 1182 410
rect 1218 378 1250 410
rect 1286 378 1318 410
rect 1354 378 1386 410
rect 1422 378 1454 410
rect 1490 378 1522 410
rect 1558 378 1590 410
rect 1626 378 1658 410
rect 1694 378 1726 410
rect 1762 378 1794 410
rect 1830 378 1862 410
rect 1898 378 1930 410
rect 1966 378 1998 410
rect 2034 378 2066 410
rect 2102 378 2134 410
rect 2170 378 2202 410
rect 2238 378 2270 410
rect 2306 378 2338 410
rect 2374 378 2406 410
rect 2442 378 2474 410
rect 2510 378 2542 410
rect 2578 378 2610 410
rect 2646 378 2678 410
rect 2714 378 2746 410
rect 2782 378 2814 410
rect 2850 378 2882 410
rect 2918 378 2950 410
rect 2986 378 3018 410
rect 3054 378 3086 410
rect 3122 378 3154 410
rect 3190 378 3222 410
rect 3258 378 3290 410
rect 3326 378 3358 410
rect 3394 378 3426 410
rect 3462 378 3494 410
rect 3530 378 3562 410
rect 3598 378 3630 410
rect 3666 378 3698 410
rect 3734 378 3766 410
rect 3802 378 3834 410
rect 3870 378 3902 410
rect 3938 378 3970 410
rect 4006 378 4038 410
rect 4074 378 4106 410
rect 4142 378 4174 410
rect 4210 378 4242 410
rect 4278 378 4310 410
rect 4346 378 4378 410
rect 4414 378 4446 410
rect 4482 378 4514 410
rect 4550 378 4582 410
rect 4618 378 4650 410
rect 4686 378 4718 410
rect 4754 378 4786 410
rect 4822 378 4854 410
rect 4890 378 4922 410
rect 4958 378 4990 410
rect 5026 378 5058 410
rect 5094 378 5126 410
rect 5162 378 5194 410
rect 5230 378 5262 410
rect 5298 378 5330 410
rect 5366 378 5398 410
rect 5434 378 5466 410
rect 5502 378 5534 410
rect 5570 378 5602 410
rect 5638 378 5670 410
rect 5706 378 5738 410
rect 5774 378 5806 410
rect 5842 378 5874 410
rect 5910 378 5942 410
rect 5978 378 6010 410
rect 6046 378 6078 410
rect 6114 378 6146 410
rect 6182 378 6214 410
rect 6250 378 6282 410
rect 6318 378 6350 410
rect 6386 378 6418 410
rect 6454 378 6486 410
rect 6522 378 6554 410
rect 6590 378 6622 410
rect 6658 378 6690 410
rect 6726 378 6758 410
rect 6794 378 6826 410
rect 6862 378 6894 410
rect 6930 378 6962 410
rect 6998 378 7030 410
rect 7066 378 7098 410
rect 7134 378 7166 410
rect 7202 378 7234 410
rect 7270 378 7302 410
rect 7338 378 7370 410
rect 7406 378 7438 410
rect 7474 378 7506 410
rect 7542 378 7574 410
rect 7610 378 7642 410
rect 7678 378 7710 410
rect 7746 378 7778 410
rect 7814 378 7846 410
rect 7882 378 7914 410
rect 7950 378 7982 410
rect 8018 378 8050 410
rect 8086 378 8118 410
rect 8154 378 8186 410
rect 8222 378 8254 410
rect 8290 378 8322 410
rect 8358 378 8390 410
rect 8426 378 8458 410
rect 8494 378 8526 410
rect 8562 378 8594 410
rect 8630 378 8662 410
rect 8698 378 8730 410
rect 8766 378 8798 410
rect 8834 378 8866 410
rect 8902 378 8934 410
rect 8970 378 9002 410
rect 9038 378 9070 410
rect 9106 378 9138 410
rect 9174 378 9206 410
rect 9242 378 9274 410
rect 9310 378 9342 410
rect 9378 378 9410 410
rect 9446 378 9478 410
rect 9514 378 9546 410
rect 9582 378 9614 410
rect 9650 378 9682 410
rect 9718 378 9750 410
rect 9786 378 9818 410
rect 9854 378 9886 410
rect 9922 378 9954 410
rect 9990 378 10022 410
rect 10058 378 10090 410
rect 10126 378 10158 410
rect 10194 378 10226 410
rect 10262 378 10294 410
rect 10330 378 10362 410
rect 10398 378 10430 410
rect 10466 378 10498 410
rect 10534 378 10566 410
rect 10602 378 10634 410
rect 10670 378 10702 410
rect 10738 378 10770 410
rect 10806 378 10838 410
rect 10874 378 10906 410
rect 10942 378 10974 410
rect 11010 378 11042 410
rect 11078 378 11110 410
rect 11146 378 11178 410
rect 11214 378 11246 410
rect 11282 378 11314 410
rect 11350 378 11382 410
rect 11418 378 11450 410
rect 11486 378 11518 410
rect 11554 378 11586 410
rect 11622 378 11654 410
rect 11690 378 11722 410
rect 11758 378 11790 410
rect 11826 378 11858 410
rect 11894 378 11926 410
rect 11962 378 11994 410
rect 12030 378 12062 410
rect 12098 378 12130 410
rect 12166 378 12198 410
rect 12234 378 12266 410
rect 12302 378 12334 410
rect 12370 378 12402 410
rect 12438 378 12470 410
rect 12506 378 12538 410
rect 12574 378 12606 410
rect 12642 378 12674 410
rect 12710 378 12742 410
rect 12778 378 12810 410
rect 12846 378 12878 410
rect 12914 378 12946 410
rect 12982 378 13014 410
rect 13050 378 13082 410
rect 13118 378 13150 410
rect 13186 378 13218 410
rect 13254 378 13286 410
rect 13322 378 13354 410
rect 13390 378 13422 410
rect 13458 378 13490 410
rect 13526 378 13558 410
rect 13594 378 13626 410
rect 13662 378 13694 410
rect 13730 378 13762 410
rect 13798 378 13830 410
rect 13866 378 13898 410
rect 13934 378 13966 410
rect 14002 378 14034 410
rect 14070 378 14102 410
rect 14138 378 14170 410
rect 14206 378 14238 410
rect 14274 378 14306 410
rect 14342 378 14374 410
rect 14410 378 14442 410
rect 14478 378 14510 410
rect 14546 378 14578 410
rect 14614 378 14646 410
rect 14682 378 14714 410
rect 14750 378 14782 410
rect 14818 378 14850 410
rect 14886 378 14918 410
rect 14954 378 14986 410
rect 15022 378 15054 410
rect 15090 378 15122 410
rect 15158 378 15190 410
rect 15226 378 15258 410
rect 15294 378 15326 410
rect 15362 378 15394 410
rect 15430 378 15462 410
rect 15498 378 15530 410
rect 15566 378 15598 410
<< nsubdiffcont >>
rect 28 1930 60 1962
rect 96 1930 128 1962
rect 164 1930 196 1962
rect 232 1930 264 1962
rect 300 1930 332 1962
rect 368 1930 400 1962
rect 436 1930 468 1962
rect 504 1930 536 1962
rect 572 1930 604 1962
rect 640 1930 672 1962
rect 708 1930 740 1962
rect 776 1930 808 1962
rect 844 1930 876 1962
rect 912 1930 944 1962
rect 980 1930 1012 1962
rect 1048 1930 1080 1962
rect 1116 1930 1148 1962
rect 1184 1930 1216 1962
rect 1252 1930 1284 1962
rect 1320 1930 1352 1962
rect 1388 1930 1420 1962
rect 1456 1930 1488 1962
rect 1524 1930 1556 1962
rect 1592 1930 1624 1962
rect 1660 1930 1692 1962
rect 1728 1930 1760 1962
rect 1796 1930 1828 1962
rect 1864 1930 1896 1962
rect 1932 1930 1964 1962
rect 2000 1930 2032 1962
rect 2068 1930 2100 1962
rect 2136 1930 2168 1962
rect 2204 1930 2236 1962
rect 2272 1930 2304 1962
rect 2340 1930 2372 1962
rect 2408 1930 2440 1962
rect 2476 1930 2508 1962
rect 2544 1930 2576 1962
rect 2612 1930 2644 1962
rect 2680 1930 2712 1962
rect 2748 1930 2780 1962
rect 2816 1930 2848 1962
rect 2884 1930 2916 1962
rect 2952 1930 2984 1962
rect 3020 1930 3052 1962
rect 3088 1930 3120 1962
rect 3156 1930 3188 1962
rect 3224 1930 3256 1962
rect 3292 1930 3324 1962
rect 3360 1930 3392 1962
rect 3428 1930 3460 1962
rect 3496 1930 3528 1962
rect 3564 1930 3596 1962
rect 3632 1930 3664 1962
rect 3700 1930 3732 1962
rect 3768 1930 3800 1962
rect 3836 1930 3868 1962
rect 3904 1930 3936 1962
rect 3972 1930 4004 1962
rect 4040 1930 4072 1962
rect 4108 1930 4140 1962
rect 4176 1930 4208 1962
rect 4244 1930 4276 1962
rect 4312 1930 4344 1962
rect 4380 1930 4412 1962
rect 4448 1930 4480 1962
rect 4516 1930 4548 1962
rect 4584 1930 4616 1962
rect 4652 1930 4684 1962
rect 4720 1930 4752 1962
rect 4788 1930 4820 1962
rect 4856 1930 4888 1962
rect 4924 1930 4956 1962
rect 4992 1930 5024 1962
rect 5060 1930 5092 1962
rect 5128 1930 5160 1962
rect 5196 1930 5228 1962
rect 5264 1930 5296 1962
rect 5332 1930 5364 1962
rect 5400 1930 5432 1962
rect 5468 1930 5500 1962
rect 5536 1930 5568 1962
rect 5604 1930 5636 1962
rect 5672 1930 5704 1962
rect 5740 1930 5772 1962
rect 5808 1930 5840 1962
rect 5876 1930 5908 1962
rect 5944 1930 5976 1962
rect 6012 1930 6044 1962
rect 6080 1930 6112 1962
rect 6148 1930 6180 1962
rect 6216 1930 6248 1962
rect 6284 1930 6316 1962
rect 6352 1930 6384 1962
rect 6420 1930 6452 1962
rect 6488 1930 6520 1962
rect 6556 1930 6588 1962
rect 6624 1930 6656 1962
rect 6692 1930 6724 1962
rect 6760 1930 6792 1962
rect 6828 1930 6860 1962
rect 6896 1930 6928 1962
rect 6964 1930 6996 1962
rect 7032 1930 7064 1962
rect 7100 1930 7132 1962
rect 7168 1930 7200 1962
rect 7236 1930 7268 1962
rect 7304 1930 7336 1962
rect 7372 1930 7404 1962
rect 7440 1930 7472 1962
rect 7508 1930 7540 1962
rect 7576 1930 7608 1962
rect 7644 1930 7676 1962
rect 7712 1930 7744 1962
rect 7780 1930 7812 1962
rect 7848 1930 7880 1962
rect 7916 1930 7948 1962
rect 7984 1930 8016 1962
rect 8052 1930 8084 1962
rect 8120 1930 8152 1962
rect 8188 1930 8220 1962
rect 8256 1930 8288 1962
rect 8324 1930 8356 1962
rect 8392 1930 8424 1962
rect 8460 1930 8492 1962
rect 8528 1930 8560 1962
rect 8596 1930 8628 1962
rect 8664 1930 8696 1962
rect 8732 1930 8764 1962
rect 8800 1930 8832 1962
rect 8868 1930 8900 1962
rect 8936 1930 8968 1962
rect 9004 1930 9036 1962
rect 9072 1930 9104 1962
rect 9140 1930 9172 1962
rect 9208 1930 9240 1962
rect 9276 1930 9308 1962
rect 9344 1930 9376 1962
rect 9412 1930 9444 1962
rect 9480 1930 9512 1962
rect 9548 1930 9580 1962
rect 9616 1930 9648 1962
rect 9684 1930 9716 1962
rect 9752 1930 9784 1962
rect 9820 1930 9852 1962
rect 9888 1930 9920 1962
rect 9956 1930 9988 1962
rect 10024 1930 10056 1962
rect 10092 1930 10124 1962
rect 10160 1930 10192 1962
rect 10228 1930 10260 1962
rect 10296 1930 10328 1962
rect 10364 1930 10396 1962
rect 10432 1930 10464 1962
rect 10500 1930 10532 1962
rect 10568 1930 10600 1962
rect 10636 1930 10668 1962
rect 10704 1930 10736 1962
rect 10772 1930 10804 1962
rect 10840 1930 10872 1962
rect 10908 1930 10940 1962
rect 10976 1930 11008 1962
rect 11044 1930 11076 1962
rect 11112 1930 11144 1962
rect 11180 1930 11212 1962
rect 11248 1930 11280 1962
rect 11316 1930 11348 1962
rect 11384 1930 11416 1962
rect 11452 1930 11484 1962
rect 11520 1930 11552 1962
rect 11588 1930 11620 1962
rect 11656 1930 11688 1962
rect 11724 1930 11756 1962
rect 11792 1930 11824 1962
rect 11860 1930 11892 1962
rect 11928 1930 11960 1962
rect 11996 1930 12028 1962
rect 12064 1930 12096 1962
rect 12132 1930 12164 1962
rect 12200 1930 12232 1962
rect 12268 1930 12300 1962
rect 12336 1930 12368 1962
rect 12404 1930 12436 1962
rect 12472 1930 12504 1962
rect 12540 1930 12572 1962
rect 12608 1930 12640 1962
rect 12676 1930 12708 1962
rect 12744 1930 12776 1962
rect 12812 1930 12844 1962
rect 12880 1930 12912 1962
rect 12948 1930 12980 1962
rect 13016 1930 13048 1962
rect 13084 1930 13116 1962
rect 13152 1930 13184 1962
rect 13220 1930 13252 1962
rect 13288 1930 13320 1962
rect 13356 1930 13388 1962
rect 13424 1930 13456 1962
rect 13492 1930 13524 1962
rect 13560 1930 13592 1962
rect 13628 1930 13660 1962
rect 13696 1930 13728 1962
rect 13764 1930 13796 1962
rect 13832 1930 13864 1962
rect 13900 1930 13932 1962
rect 13968 1930 14000 1962
rect 14036 1930 14068 1962
rect 14104 1930 14136 1962
rect 14172 1930 14204 1962
rect 14240 1930 14272 1962
rect 14308 1930 14340 1962
rect 14376 1930 14408 1962
rect 14444 1930 14476 1962
rect 14512 1930 14544 1962
rect 14580 1930 14612 1962
rect 14648 1930 14680 1962
rect 14716 1930 14748 1962
rect 14784 1930 14816 1962
rect 14852 1930 14884 1962
rect 14920 1930 14952 1962
rect 14988 1930 15020 1962
rect 15056 1930 15088 1962
rect 15124 1930 15156 1962
rect 15192 1930 15224 1962
rect 15260 1930 15292 1962
rect 15328 1930 15360 1962
rect 15396 1930 15428 1962
rect 15464 1930 15496 1962
rect 15532 1930 15564 1962
rect 15600 1930 15632 1962
rect 15668 1930 15700 1962
rect 15736 1930 15768 1962
rect 15804 1930 15836 1962
rect 15872 1930 15904 1962
rect 15940 1930 15972 1962
rect 18 1824 50 1856
rect 18 1756 50 1788
rect 18 1688 50 1720
rect 18 1620 50 1652
rect 15950 1824 15982 1856
rect 15950 1756 15982 1788
rect 15950 1688 15982 1720
rect 15950 1620 15982 1652
rect 18 1552 50 1584
rect 18 1484 50 1516
rect 18 1416 50 1448
rect 18 1348 50 1380
rect 18 1280 50 1312
rect 18 1212 50 1244
rect 18 1144 50 1176
rect 18 1076 50 1108
rect 18 1008 50 1040
rect 18 940 50 972
rect 18 872 50 904
rect 18 804 50 836
rect 18 736 50 768
rect 18 668 50 700
rect 18 600 50 632
rect 18 532 50 564
rect 18 464 50 496
rect 18 396 50 428
rect 15950 1552 15982 1584
rect 15950 1484 15982 1516
rect 15950 1416 15982 1448
rect 15950 1348 15982 1380
rect 15950 1280 15982 1312
rect 15950 1212 15982 1244
rect 15950 1144 15982 1176
rect 15950 1076 15982 1108
rect 15950 1008 15982 1040
rect 15950 940 15982 972
rect 15950 872 15982 904
rect 15950 804 15982 836
rect 15950 736 15982 768
rect 15950 668 15982 700
rect 15950 600 15982 632
rect 15950 532 15982 564
rect 15950 464 15982 496
rect 15950 396 15982 428
rect 18 328 50 360
rect 18 260 50 292
rect 18 192 50 224
rect 18 124 50 156
rect 15950 328 15982 360
rect 15950 260 15982 292
rect 15950 192 15982 224
rect 15950 124 15982 156
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< poly >>
rect 5799 1490 5919 1504
rect 5799 1458 5843 1490
rect 5875 1458 5919 1490
rect 5799 1430 5919 1458
rect 6155 1490 6275 1504
rect 6155 1458 6199 1490
rect 6231 1458 6275 1490
rect 6155 1430 6275 1458
rect 6403 1490 6523 1504
rect 6403 1458 6447 1490
rect 6479 1458 6523 1490
rect 6403 1430 6523 1458
rect 6759 1490 6879 1504
rect 6759 1458 6803 1490
rect 6835 1458 6879 1490
rect 6759 1430 6879 1458
rect 7007 1490 7127 1504
rect 7007 1458 7051 1490
rect 7083 1458 7127 1490
rect 7007 1430 7127 1458
rect 7363 1490 7483 1504
rect 7363 1458 7407 1490
rect 7439 1458 7483 1490
rect 7363 1430 7483 1458
rect 7611 1490 7731 1504
rect 7611 1458 7655 1490
rect 7687 1458 7731 1490
rect 7611 1430 7731 1458
rect 7967 1490 8087 1504
rect 7967 1458 8011 1490
rect 8043 1458 8087 1490
rect 7967 1430 8087 1458
rect 8215 1490 8335 1504
rect 8215 1458 8259 1490
rect 8291 1458 8335 1490
rect 8215 1430 8335 1458
rect 8571 1490 8691 1504
rect 8571 1458 8615 1490
rect 8647 1458 8691 1490
rect 8571 1430 8691 1458
rect 8819 1490 8939 1504
rect 8819 1458 8863 1490
rect 8895 1458 8939 1490
rect 8819 1430 8939 1458
rect 9175 1490 9295 1504
rect 9175 1458 9219 1490
rect 9251 1458 9295 1490
rect 9175 1430 9295 1458
rect 9423 1490 9543 1504
rect 9423 1458 9467 1490
rect 9499 1458 9543 1490
rect 9423 1430 9543 1458
rect 9779 1490 9899 1504
rect 9779 1458 9823 1490
rect 9855 1458 9899 1490
rect 9779 1430 9899 1458
rect 10027 1490 10147 1504
rect 10027 1458 10071 1490
rect 10103 1458 10147 1490
rect 10027 1430 10147 1458
rect 5799 522 5919 550
rect 5799 490 5843 522
rect 5875 490 5919 522
rect 5799 476 5919 490
rect 6155 522 6275 550
rect 6155 490 6199 522
rect 6231 490 6275 522
rect 6155 476 6275 490
rect 6403 522 6523 550
rect 6403 490 6447 522
rect 6479 490 6523 522
rect 6403 476 6523 490
rect 6759 522 6879 550
rect 6759 490 6803 522
rect 6835 490 6879 522
rect 6759 476 6879 490
rect 7007 522 7127 550
rect 7007 490 7051 522
rect 7083 490 7127 522
rect 7007 476 7127 490
rect 7363 522 7483 550
rect 7363 490 7407 522
rect 7439 490 7483 522
rect 7363 476 7483 490
rect 7611 522 7731 550
rect 7611 490 7655 522
rect 7687 490 7731 522
rect 7611 476 7731 490
rect 7967 522 8087 550
rect 7967 490 8011 522
rect 8043 490 8087 522
rect 7967 476 8087 490
rect 8215 522 8335 550
rect 8215 490 8259 522
rect 8291 490 8335 522
rect 8215 476 8335 490
rect 8571 522 8691 550
rect 8571 490 8615 522
rect 8647 490 8691 522
rect 8571 476 8691 490
rect 8819 522 8939 550
rect 8819 490 8863 522
rect 8895 490 8939 522
rect 8819 476 8939 490
rect 9175 522 9295 550
rect 9175 490 9219 522
rect 9251 490 9295 522
rect 9175 476 9295 490
rect 9423 522 9543 550
rect 9423 490 9467 522
rect 9499 490 9543 522
rect 9423 476 9543 490
rect 9779 522 9899 550
rect 9779 490 9823 522
rect 9855 490 9899 522
rect 9779 476 9899 490
rect 10027 522 10147 550
rect 10027 490 10071 522
rect 10103 490 10147 522
rect 10027 476 10147 490
<< polycont >>
rect 5843 1458 5875 1490
rect 6199 1458 6231 1490
rect 6447 1458 6479 1490
rect 6803 1458 6835 1490
rect 7051 1458 7083 1490
rect 7407 1458 7439 1490
rect 7655 1458 7687 1490
rect 8011 1458 8043 1490
rect 8259 1458 8291 1490
rect 8615 1458 8647 1490
rect 8863 1458 8895 1490
rect 9219 1458 9251 1490
rect 9467 1458 9499 1490
rect 9823 1458 9855 1490
rect 10071 1458 10103 1490
rect 5843 490 5875 522
rect 6199 490 6231 522
rect 6447 490 6479 522
rect 6803 490 6835 522
rect 7051 490 7083 522
rect 7407 490 7439 522
rect 7655 490 7687 522
rect 8011 490 8043 522
rect 8259 490 8291 522
rect 8615 490 8647 522
rect 8863 490 8895 522
rect 9219 490 9251 522
rect 9467 490 9499 522
rect 9823 490 9855 522
rect 10071 490 10103 522
<< ndiode >>
rect 2986 1391 3142 1419
rect 2986 1359 3014 1391
rect 3046 1359 3082 1391
rect 3114 1359 3142 1391
rect 2986 1323 3142 1359
rect 2986 1291 3014 1323
rect 3046 1291 3082 1323
rect 3114 1291 3142 1323
rect 2986 1263 3142 1291
<< ndiodecont >>
rect 3014 1359 3046 1391
rect 3082 1359 3114 1391
rect 3014 1291 3046 1323
rect 3082 1291 3114 1323
<< metal1 >>
rect 0 1962 16000 1980
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 360 1606 15640 1620
rect 360 1602 5715 1606
rect 5755 1602 6319 1606
rect 6359 1602 6923 1606
rect 6963 1602 7527 1606
rect 7567 1602 8131 1606
rect 8171 1602 8735 1606
rect 8775 1602 9339 1606
rect 9379 1602 9943 1606
rect 9983 1602 15640 1606
rect 360 1570 402 1602
rect 434 1570 470 1602
rect 502 1570 538 1602
rect 570 1570 606 1602
rect 638 1570 674 1602
rect 706 1570 742 1602
rect 774 1570 810 1602
rect 842 1570 878 1602
rect 910 1570 946 1602
rect 978 1570 1014 1602
rect 1046 1570 1082 1602
rect 1114 1570 1150 1602
rect 1182 1570 1218 1602
rect 1250 1570 1286 1602
rect 1318 1570 1354 1602
rect 1386 1570 1422 1602
rect 1454 1570 1490 1602
rect 1522 1570 1558 1602
rect 1590 1570 1626 1602
rect 1658 1570 1694 1602
rect 1726 1570 1762 1602
rect 1794 1570 1830 1602
rect 1862 1570 1898 1602
rect 1930 1570 1966 1602
rect 1998 1570 2034 1602
rect 2066 1570 2102 1602
rect 2134 1570 2170 1602
rect 2202 1570 2238 1602
rect 2270 1570 2306 1602
rect 2338 1570 2374 1602
rect 2406 1570 2442 1602
rect 2474 1570 2510 1602
rect 2542 1570 2578 1602
rect 2610 1570 2646 1602
rect 2678 1570 2714 1602
rect 2746 1570 2782 1602
rect 2814 1570 2850 1602
rect 2882 1570 2918 1602
rect 2950 1570 2986 1602
rect 3018 1570 3054 1602
rect 3086 1570 3122 1602
rect 3154 1570 3190 1602
rect 3222 1570 3258 1602
rect 3290 1570 3326 1602
rect 3358 1570 3394 1602
rect 3426 1570 3462 1602
rect 3494 1570 3530 1602
rect 3562 1570 3598 1602
rect 3630 1570 3666 1602
rect 3698 1570 3734 1602
rect 3766 1570 3802 1602
rect 3834 1570 3870 1602
rect 3902 1570 3938 1602
rect 3970 1570 4006 1602
rect 4038 1570 4074 1602
rect 4106 1570 4142 1602
rect 4174 1570 4210 1602
rect 4242 1570 4278 1602
rect 4310 1570 4346 1602
rect 4378 1570 4414 1602
rect 4446 1570 4482 1602
rect 4514 1570 4550 1602
rect 4582 1570 4618 1602
rect 4650 1570 4686 1602
rect 4718 1570 4754 1602
rect 4786 1570 4822 1602
rect 4854 1570 4890 1602
rect 4922 1570 4958 1602
rect 4990 1570 5026 1602
rect 5058 1570 5094 1602
rect 5126 1570 5162 1602
rect 5194 1570 5230 1602
rect 5262 1570 5298 1602
rect 5330 1570 5366 1602
rect 5398 1570 5434 1602
rect 5466 1570 5502 1602
rect 5534 1570 5570 1602
rect 5602 1570 5638 1602
rect 5670 1570 5706 1602
rect 5755 1570 5774 1602
rect 5806 1570 5842 1602
rect 5874 1570 5910 1602
rect 5942 1570 5978 1602
rect 6010 1570 6046 1602
rect 6078 1570 6114 1602
rect 6146 1570 6182 1602
rect 6214 1570 6250 1602
rect 6282 1570 6318 1602
rect 6359 1570 6386 1602
rect 6418 1570 6454 1602
rect 6486 1570 6522 1602
rect 6554 1570 6590 1602
rect 6622 1570 6658 1602
rect 6690 1570 6726 1602
rect 6758 1570 6794 1602
rect 6826 1570 6862 1602
rect 6894 1570 6923 1602
rect 6963 1570 6998 1602
rect 7030 1570 7066 1602
rect 7098 1570 7134 1602
rect 7166 1570 7202 1602
rect 7234 1570 7270 1602
rect 7302 1570 7338 1602
rect 7370 1570 7406 1602
rect 7438 1570 7474 1602
rect 7506 1570 7527 1602
rect 7574 1570 7610 1602
rect 7642 1570 7678 1602
rect 7710 1570 7746 1602
rect 7778 1570 7814 1602
rect 7846 1570 7882 1602
rect 7914 1570 7950 1602
rect 7982 1570 8018 1602
rect 8050 1570 8086 1602
rect 8118 1570 8131 1602
rect 8186 1570 8222 1602
rect 8254 1570 8290 1602
rect 8322 1570 8358 1602
rect 8390 1570 8426 1602
rect 8458 1570 8494 1602
rect 8526 1570 8562 1602
rect 8594 1570 8630 1602
rect 8662 1570 8698 1602
rect 8730 1570 8735 1602
rect 8798 1570 8834 1602
rect 8866 1570 8902 1602
rect 8934 1570 8970 1602
rect 9002 1570 9038 1602
rect 9070 1570 9106 1602
rect 9138 1570 9174 1602
rect 9206 1570 9242 1602
rect 9274 1570 9310 1602
rect 9410 1570 9446 1602
rect 9478 1570 9514 1602
rect 9546 1570 9582 1602
rect 9614 1570 9650 1602
rect 9682 1570 9718 1602
rect 9750 1570 9786 1602
rect 9818 1570 9854 1602
rect 9886 1570 9922 1602
rect 9983 1570 9990 1602
rect 10022 1570 10058 1602
rect 10090 1570 10126 1602
rect 10158 1570 10194 1602
rect 10226 1570 10262 1602
rect 10294 1570 10330 1602
rect 10362 1570 10398 1602
rect 10430 1570 10466 1602
rect 10498 1570 10534 1602
rect 10566 1570 10602 1602
rect 10634 1570 10670 1602
rect 10702 1570 10738 1602
rect 10770 1570 10806 1602
rect 10838 1570 10874 1602
rect 10906 1570 10942 1602
rect 10974 1570 11010 1602
rect 11042 1570 11078 1602
rect 11110 1570 11146 1602
rect 11178 1570 11214 1602
rect 11246 1570 11282 1602
rect 11314 1570 11350 1602
rect 11382 1570 11418 1602
rect 11450 1570 11486 1602
rect 11518 1570 11554 1602
rect 11586 1570 11622 1602
rect 11654 1570 11690 1602
rect 11722 1570 11758 1602
rect 11790 1570 11826 1602
rect 11858 1570 11894 1602
rect 11926 1570 11962 1602
rect 11994 1570 12030 1602
rect 12062 1570 12098 1602
rect 12130 1570 12166 1602
rect 12198 1570 12234 1602
rect 12266 1570 12302 1602
rect 12334 1570 12370 1602
rect 12402 1570 12438 1602
rect 12470 1570 12506 1602
rect 12538 1570 12574 1602
rect 12606 1570 12642 1602
rect 12674 1570 12710 1602
rect 12742 1570 12778 1602
rect 12810 1570 12846 1602
rect 12878 1570 12914 1602
rect 12946 1570 12982 1602
rect 13014 1570 13050 1602
rect 13082 1570 13118 1602
rect 13150 1570 13186 1602
rect 13218 1570 13254 1602
rect 13286 1570 13322 1602
rect 13354 1570 13390 1602
rect 13422 1570 13458 1602
rect 13490 1570 13526 1602
rect 13558 1570 13594 1602
rect 13626 1570 13662 1602
rect 13694 1570 13730 1602
rect 13762 1570 13798 1602
rect 13830 1570 13866 1602
rect 13898 1570 13934 1602
rect 13966 1570 14002 1602
rect 14034 1570 14070 1602
rect 14102 1570 14138 1602
rect 14170 1570 14206 1602
rect 14238 1570 14274 1602
rect 14306 1570 14342 1602
rect 14374 1570 14410 1602
rect 14442 1570 14478 1602
rect 14510 1570 14546 1602
rect 14578 1570 14614 1602
rect 14646 1570 14682 1602
rect 14714 1570 14750 1602
rect 14782 1570 14818 1602
rect 14850 1570 14886 1602
rect 14918 1570 14954 1602
rect 14986 1570 15022 1602
rect 15054 1570 15090 1602
rect 15122 1570 15158 1602
rect 15190 1570 15226 1602
rect 15258 1570 15294 1602
rect 15326 1570 15362 1602
rect 15394 1570 15430 1602
rect 15462 1570 15498 1602
rect 15530 1570 15566 1602
rect 15598 1570 15640 1602
rect 360 1566 5715 1570
rect 5755 1566 6319 1570
rect 6359 1566 6923 1570
rect 6963 1566 7527 1570
rect 7567 1566 8131 1570
rect 8171 1566 8735 1570
rect 8775 1566 9339 1570
rect 9379 1566 9943 1570
rect 9983 1566 15640 1570
rect 360 1552 15640 1566
rect 360 1516 428 1552
rect 360 1484 378 1516
rect 410 1484 428 1516
rect 15572 1516 15640 1552
rect 360 1448 428 1484
rect 360 1416 378 1448
rect 410 1416 428 1448
rect 360 1380 428 1416
rect 3045 1490 10103 1506
rect 3045 1474 5843 1490
rect 3045 1464 3087 1474
rect 3045 1391 3046 1464
rect 360 1348 378 1380
rect 410 1348 428 1380
rect 360 1312 428 1348
rect 360 1280 378 1312
rect 410 1280 428 1312
rect 3004 1342 3046 1391
rect 3086 1391 3087 1464
rect 5875 1474 6199 1490
rect 5714 1420 5756 1430
rect 3086 1342 3124 1391
rect 3004 1291 3124 1342
rect 360 1244 428 1280
rect 360 1212 378 1244
rect 410 1212 428 1244
rect 360 1176 428 1212
rect 360 1144 378 1176
rect 410 1144 428 1176
rect 360 1108 428 1144
rect 360 1076 378 1108
rect 410 1076 428 1108
rect 360 1040 428 1076
rect 360 1008 378 1040
rect 410 1008 428 1040
rect 360 972 428 1008
rect 360 940 378 972
rect 410 940 428 972
rect 360 904 428 940
rect 360 872 378 904
rect 410 872 428 904
rect 360 836 428 872
rect 360 804 378 836
rect 410 804 428 836
rect 360 768 428 804
rect 360 736 378 768
rect 410 736 428 768
rect 360 700 428 736
rect 360 668 378 700
rect 410 668 428 700
rect 360 632 428 668
rect 360 600 378 632
rect 410 600 428 632
rect 360 564 428 600
rect 360 532 378 564
rect 410 532 428 564
rect 5714 560 5715 1420
rect 5755 560 5756 1420
rect 5714 550 5756 560
rect 360 496 428 532
rect 360 464 378 496
rect 410 464 428 496
rect 5843 522 5875 1458
rect 6231 1474 6447 1490
rect 5975 1420 6099 1430
rect 5975 560 5976 1420
rect 6098 560 6099 1420
rect 5975 550 6099 560
rect 5843 474 5875 490
rect 6199 522 6231 1458
rect 6479 1474 6803 1490
rect 6318 1420 6360 1430
rect 6318 560 6319 1420
rect 6359 560 6360 1420
rect 6318 550 6360 560
rect 6199 474 6231 490
rect 6447 522 6479 1458
rect 6835 1474 7051 1490
rect 6579 1420 6703 1430
rect 6579 560 6580 1420
rect 6702 560 6703 1420
rect 6579 550 6703 560
rect 6447 474 6479 490
rect 6803 522 6835 1458
rect 7083 1474 7407 1490
rect 6922 1420 6964 1430
rect 6922 560 6923 1420
rect 6963 560 6964 1420
rect 6922 550 6964 560
rect 6803 474 6835 490
rect 7051 522 7083 1458
rect 7439 1474 7655 1490
rect 7183 1420 7307 1430
rect 7183 560 7184 1420
rect 7306 560 7307 1420
rect 7183 550 7307 560
rect 7051 474 7083 490
rect 7407 522 7439 1458
rect 7687 1474 8011 1490
rect 7526 1420 7568 1430
rect 7526 560 7527 1420
rect 7567 560 7568 1420
rect 7526 550 7568 560
rect 7407 474 7439 490
rect 7655 522 7687 1458
rect 8043 1474 8259 1490
rect 7787 1420 7911 1430
rect 7787 560 7788 1420
rect 7910 560 7911 1420
rect 7787 550 7911 560
rect 7655 474 7687 490
rect 8011 522 8043 1458
rect 8291 1474 8615 1490
rect 8130 1420 8172 1430
rect 8130 560 8131 1420
rect 8171 560 8172 1420
rect 8130 550 8172 560
rect 8011 474 8043 490
rect 8259 522 8291 1458
rect 8647 1474 8863 1490
rect 8391 1420 8515 1430
rect 8391 560 8392 1420
rect 8514 560 8515 1420
rect 8391 550 8515 560
rect 8259 474 8291 490
rect 8615 522 8647 1458
rect 8895 1474 9219 1490
rect 8734 1420 8776 1430
rect 8734 560 8735 1420
rect 8775 560 8776 1420
rect 8734 550 8776 560
rect 8615 474 8647 490
rect 8863 522 8895 1458
rect 9251 1474 9467 1490
rect 8995 1420 9119 1430
rect 8995 560 8996 1420
rect 9118 560 9119 1420
rect 8995 550 9119 560
rect 8863 474 8895 490
rect 9219 522 9251 1458
rect 9499 1474 9823 1490
rect 9338 1420 9380 1430
rect 9338 560 9339 1420
rect 9379 560 9380 1420
rect 9338 550 9380 560
rect 9219 474 9251 490
rect 9467 522 9499 1458
rect 9855 1474 10071 1490
rect 9599 1420 9723 1430
rect 9599 560 9600 1420
rect 9722 560 9723 1420
rect 9599 550 9723 560
rect 9467 474 9499 490
rect 9823 522 9855 1458
rect 9942 1420 9984 1430
rect 9942 560 9943 1420
rect 9983 560 9984 1420
rect 9942 550 9984 560
rect 9823 474 9855 490
rect 10071 522 10103 1458
rect 15572 1484 15590 1516
rect 15622 1484 15640 1516
rect 15572 1448 15640 1484
rect 10203 1420 10327 1430
rect 10203 560 10204 1420
rect 10326 560 10327 1420
rect 10203 550 10327 560
rect 15572 1416 15590 1448
rect 15622 1416 15640 1448
rect 15572 1380 15640 1416
rect 15572 1348 15590 1380
rect 15622 1348 15640 1380
rect 15572 1312 15640 1348
rect 15572 1280 15590 1312
rect 15622 1280 15640 1312
rect 15572 1244 15640 1280
rect 15572 1212 15590 1244
rect 15622 1212 15640 1244
rect 15572 1176 15640 1212
rect 15572 1144 15590 1176
rect 15622 1144 15640 1176
rect 15572 1108 15640 1144
rect 15572 1076 15590 1108
rect 15622 1076 15640 1108
rect 15572 1040 15640 1076
rect 15572 1008 15590 1040
rect 15622 1008 15640 1040
rect 15572 972 15640 1008
rect 15572 940 15590 972
rect 15622 940 15640 972
rect 15572 904 15640 940
rect 15572 872 15590 904
rect 15622 872 15640 904
rect 15572 836 15640 872
rect 15572 804 15590 836
rect 15622 804 15640 836
rect 15572 768 15640 804
rect 15572 736 15590 768
rect 15622 736 15640 768
rect 15572 700 15640 736
rect 15572 668 15590 700
rect 15622 668 15640 700
rect 15572 632 15640 668
rect 15572 600 15590 632
rect 15622 600 15640 632
rect 15572 564 15640 600
rect 10071 474 10103 490
rect 15572 532 15590 564
rect 15622 532 15640 564
rect 15572 496 15640 532
rect 360 428 428 464
rect 15572 464 15590 496
rect 15622 464 15640 496
rect 15572 428 15640 464
rect 360 414 15640 428
rect 360 410 5715 414
rect 5755 410 6319 414
rect 6359 410 6923 414
rect 6963 410 7527 414
rect 7567 410 8131 414
rect 8171 410 8735 414
rect 8775 410 9339 414
rect 9379 410 9943 414
rect 9983 410 15640 414
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5755 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6359 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6923 410
rect 6963 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7527 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8131 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8735 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9983 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 374 5715 378
rect 5755 374 6319 378
rect 6359 374 6923 378
rect 6963 374 7527 378
rect 7567 374 8131 378
rect 8171 374 8735 378
rect 8775 374 9339 378
rect 9379 374 9943 378
rect 9983 374 15640 378
rect 360 360 15640 374
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 15932 360 16000 396
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 5715 1602 5755 1606
rect 6319 1602 6359 1606
rect 6923 1602 6963 1606
rect 7527 1602 7567 1606
rect 8131 1602 8171 1606
rect 8735 1602 8775 1606
rect 9339 1602 9379 1606
rect 9943 1602 9983 1606
rect 5715 1570 5738 1602
rect 5738 1570 5755 1602
rect 6319 1570 6350 1602
rect 6350 1570 6359 1602
rect 6923 1570 6930 1602
rect 6930 1570 6962 1602
rect 6962 1570 6963 1602
rect 7527 1570 7542 1602
rect 7542 1570 7567 1602
rect 8131 1570 8154 1602
rect 8154 1570 8171 1602
rect 8735 1570 8766 1602
rect 8766 1570 8775 1602
rect 9339 1570 9342 1602
rect 9342 1570 9378 1602
rect 9378 1570 9379 1602
rect 9943 1570 9954 1602
rect 9954 1570 9983 1602
rect 5715 1566 5755 1570
rect 6319 1566 6359 1570
rect 6923 1566 6963 1570
rect 7527 1566 7567 1570
rect 8131 1566 8171 1570
rect 8735 1566 8775 1570
rect 9339 1566 9379 1570
rect 9943 1566 9983 1570
rect 3046 1342 3086 1464
rect 5715 1414 5755 1420
rect 5715 1382 5719 1414
rect 5719 1382 5751 1414
rect 5751 1382 5755 1414
rect 5715 1346 5755 1382
rect 5715 1314 5719 1346
rect 5719 1314 5751 1346
rect 5751 1314 5755 1346
rect 5715 1278 5755 1314
rect 5715 1246 5719 1278
rect 5719 1246 5751 1278
rect 5751 1246 5755 1278
rect 5715 1210 5755 1246
rect 5715 1178 5719 1210
rect 5719 1178 5751 1210
rect 5751 1178 5755 1210
rect 5715 1142 5755 1178
rect 5715 1110 5719 1142
rect 5719 1110 5751 1142
rect 5751 1110 5755 1142
rect 5715 1074 5755 1110
rect 5715 1042 5719 1074
rect 5719 1042 5751 1074
rect 5751 1042 5755 1074
rect 5715 1006 5755 1042
rect 5715 974 5719 1006
rect 5719 974 5751 1006
rect 5751 974 5755 1006
rect 5715 938 5755 974
rect 5715 906 5719 938
rect 5719 906 5751 938
rect 5751 906 5755 938
rect 5715 870 5755 906
rect 5715 838 5719 870
rect 5719 838 5751 870
rect 5751 838 5755 870
rect 5715 802 5755 838
rect 5715 770 5719 802
rect 5719 770 5751 802
rect 5751 770 5755 802
rect 5715 734 5755 770
rect 5715 702 5719 734
rect 5719 702 5751 734
rect 5751 702 5755 734
rect 5715 666 5755 702
rect 5715 634 5719 666
rect 5719 634 5751 666
rect 5751 634 5755 666
rect 5715 598 5755 634
rect 5715 566 5719 598
rect 5719 566 5751 598
rect 5751 566 5755 598
rect 5715 560 5755 566
rect 5976 1414 6098 1420
rect 5976 1382 6021 1414
rect 6021 1382 6053 1414
rect 6053 1382 6098 1414
rect 5976 1346 6098 1382
rect 5976 1314 6021 1346
rect 6021 1314 6053 1346
rect 6053 1314 6098 1346
rect 5976 1278 6098 1314
rect 5976 1246 6021 1278
rect 6021 1246 6053 1278
rect 6053 1246 6098 1278
rect 5976 1210 6098 1246
rect 5976 1178 6021 1210
rect 6021 1178 6053 1210
rect 6053 1178 6098 1210
rect 5976 1142 6098 1178
rect 5976 1110 6021 1142
rect 6021 1110 6053 1142
rect 6053 1110 6098 1142
rect 5976 1074 6098 1110
rect 5976 1042 6021 1074
rect 6021 1042 6053 1074
rect 6053 1042 6098 1074
rect 5976 1006 6098 1042
rect 5976 974 6021 1006
rect 6021 974 6053 1006
rect 6053 974 6098 1006
rect 5976 938 6098 974
rect 5976 906 6021 938
rect 6021 906 6053 938
rect 6053 906 6098 938
rect 5976 870 6098 906
rect 5976 838 6021 870
rect 6021 838 6053 870
rect 6053 838 6098 870
rect 5976 802 6098 838
rect 5976 770 6021 802
rect 6021 770 6053 802
rect 6053 770 6098 802
rect 5976 734 6098 770
rect 5976 702 6021 734
rect 6021 702 6053 734
rect 6053 702 6098 734
rect 5976 666 6098 702
rect 5976 634 6021 666
rect 6021 634 6053 666
rect 6053 634 6098 666
rect 5976 598 6098 634
rect 5976 566 6021 598
rect 6021 566 6053 598
rect 6053 566 6098 598
rect 5976 560 6098 566
rect 6319 1414 6359 1420
rect 6319 1382 6323 1414
rect 6323 1382 6355 1414
rect 6355 1382 6359 1414
rect 6319 1346 6359 1382
rect 6319 1314 6323 1346
rect 6323 1314 6355 1346
rect 6355 1314 6359 1346
rect 6319 1278 6359 1314
rect 6319 1246 6323 1278
rect 6323 1246 6355 1278
rect 6355 1246 6359 1278
rect 6319 1210 6359 1246
rect 6319 1178 6323 1210
rect 6323 1178 6355 1210
rect 6355 1178 6359 1210
rect 6319 1142 6359 1178
rect 6319 1110 6323 1142
rect 6323 1110 6355 1142
rect 6355 1110 6359 1142
rect 6319 1074 6359 1110
rect 6319 1042 6323 1074
rect 6323 1042 6355 1074
rect 6355 1042 6359 1074
rect 6319 1006 6359 1042
rect 6319 974 6323 1006
rect 6323 974 6355 1006
rect 6355 974 6359 1006
rect 6319 938 6359 974
rect 6319 906 6323 938
rect 6323 906 6355 938
rect 6355 906 6359 938
rect 6319 870 6359 906
rect 6319 838 6323 870
rect 6323 838 6355 870
rect 6355 838 6359 870
rect 6319 802 6359 838
rect 6319 770 6323 802
rect 6323 770 6355 802
rect 6355 770 6359 802
rect 6319 734 6359 770
rect 6319 702 6323 734
rect 6323 702 6355 734
rect 6355 702 6359 734
rect 6319 666 6359 702
rect 6319 634 6323 666
rect 6323 634 6355 666
rect 6355 634 6359 666
rect 6319 598 6359 634
rect 6319 566 6323 598
rect 6323 566 6355 598
rect 6355 566 6359 598
rect 6319 560 6359 566
rect 6580 1414 6702 1420
rect 6580 1382 6625 1414
rect 6625 1382 6657 1414
rect 6657 1382 6702 1414
rect 6580 1346 6702 1382
rect 6580 1314 6625 1346
rect 6625 1314 6657 1346
rect 6657 1314 6702 1346
rect 6580 1278 6702 1314
rect 6580 1246 6625 1278
rect 6625 1246 6657 1278
rect 6657 1246 6702 1278
rect 6580 1210 6702 1246
rect 6580 1178 6625 1210
rect 6625 1178 6657 1210
rect 6657 1178 6702 1210
rect 6580 1142 6702 1178
rect 6580 1110 6625 1142
rect 6625 1110 6657 1142
rect 6657 1110 6702 1142
rect 6580 1074 6702 1110
rect 6580 1042 6625 1074
rect 6625 1042 6657 1074
rect 6657 1042 6702 1074
rect 6580 1006 6702 1042
rect 6580 974 6625 1006
rect 6625 974 6657 1006
rect 6657 974 6702 1006
rect 6580 938 6702 974
rect 6580 906 6625 938
rect 6625 906 6657 938
rect 6657 906 6702 938
rect 6580 870 6702 906
rect 6580 838 6625 870
rect 6625 838 6657 870
rect 6657 838 6702 870
rect 6580 802 6702 838
rect 6580 770 6625 802
rect 6625 770 6657 802
rect 6657 770 6702 802
rect 6580 734 6702 770
rect 6580 702 6625 734
rect 6625 702 6657 734
rect 6657 702 6702 734
rect 6580 666 6702 702
rect 6580 634 6625 666
rect 6625 634 6657 666
rect 6657 634 6702 666
rect 6580 598 6702 634
rect 6580 566 6625 598
rect 6625 566 6657 598
rect 6657 566 6702 598
rect 6580 560 6702 566
rect 6923 1414 6963 1420
rect 6923 1382 6927 1414
rect 6927 1382 6959 1414
rect 6959 1382 6963 1414
rect 6923 1346 6963 1382
rect 6923 1314 6927 1346
rect 6927 1314 6959 1346
rect 6959 1314 6963 1346
rect 6923 1278 6963 1314
rect 6923 1246 6927 1278
rect 6927 1246 6959 1278
rect 6959 1246 6963 1278
rect 6923 1210 6963 1246
rect 6923 1178 6927 1210
rect 6927 1178 6959 1210
rect 6959 1178 6963 1210
rect 6923 1142 6963 1178
rect 6923 1110 6927 1142
rect 6927 1110 6959 1142
rect 6959 1110 6963 1142
rect 6923 1074 6963 1110
rect 6923 1042 6927 1074
rect 6927 1042 6959 1074
rect 6959 1042 6963 1074
rect 6923 1006 6963 1042
rect 6923 974 6927 1006
rect 6927 974 6959 1006
rect 6959 974 6963 1006
rect 6923 938 6963 974
rect 6923 906 6927 938
rect 6927 906 6959 938
rect 6959 906 6963 938
rect 6923 870 6963 906
rect 6923 838 6927 870
rect 6927 838 6959 870
rect 6959 838 6963 870
rect 6923 802 6963 838
rect 6923 770 6927 802
rect 6927 770 6959 802
rect 6959 770 6963 802
rect 6923 734 6963 770
rect 6923 702 6927 734
rect 6927 702 6959 734
rect 6959 702 6963 734
rect 6923 666 6963 702
rect 6923 634 6927 666
rect 6927 634 6959 666
rect 6959 634 6963 666
rect 6923 598 6963 634
rect 6923 566 6927 598
rect 6927 566 6959 598
rect 6959 566 6963 598
rect 6923 560 6963 566
rect 7184 1414 7306 1420
rect 7184 1382 7229 1414
rect 7229 1382 7261 1414
rect 7261 1382 7306 1414
rect 7184 1346 7306 1382
rect 7184 1314 7229 1346
rect 7229 1314 7261 1346
rect 7261 1314 7306 1346
rect 7184 1278 7306 1314
rect 7184 1246 7229 1278
rect 7229 1246 7261 1278
rect 7261 1246 7306 1278
rect 7184 1210 7306 1246
rect 7184 1178 7229 1210
rect 7229 1178 7261 1210
rect 7261 1178 7306 1210
rect 7184 1142 7306 1178
rect 7184 1110 7229 1142
rect 7229 1110 7261 1142
rect 7261 1110 7306 1142
rect 7184 1074 7306 1110
rect 7184 1042 7229 1074
rect 7229 1042 7261 1074
rect 7261 1042 7306 1074
rect 7184 1006 7306 1042
rect 7184 974 7229 1006
rect 7229 974 7261 1006
rect 7261 974 7306 1006
rect 7184 938 7306 974
rect 7184 906 7229 938
rect 7229 906 7261 938
rect 7261 906 7306 938
rect 7184 870 7306 906
rect 7184 838 7229 870
rect 7229 838 7261 870
rect 7261 838 7306 870
rect 7184 802 7306 838
rect 7184 770 7229 802
rect 7229 770 7261 802
rect 7261 770 7306 802
rect 7184 734 7306 770
rect 7184 702 7229 734
rect 7229 702 7261 734
rect 7261 702 7306 734
rect 7184 666 7306 702
rect 7184 634 7229 666
rect 7229 634 7261 666
rect 7261 634 7306 666
rect 7184 598 7306 634
rect 7184 566 7229 598
rect 7229 566 7261 598
rect 7261 566 7306 598
rect 7184 560 7306 566
rect 7527 1414 7567 1420
rect 7527 1382 7531 1414
rect 7531 1382 7563 1414
rect 7563 1382 7567 1414
rect 7527 1346 7567 1382
rect 7527 1314 7531 1346
rect 7531 1314 7563 1346
rect 7563 1314 7567 1346
rect 7527 1278 7567 1314
rect 7527 1246 7531 1278
rect 7531 1246 7563 1278
rect 7563 1246 7567 1278
rect 7527 1210 7567 1246
rect 7527 1178 7531 1210
rect 7531 1178 7563 1210
rect 7563 1178 7567 1210
rect 7527 1142 7567 1178
rect 7527 1110 7531 1142
rect 7531 1110 7563 1142
rect 7563 1110 7567 1142
rect 7527 1074 7567 1110
rect 7527 1042 7531 1074
rect 7531 1042 7563 1074
rect 7563 1042 7567 1074
rect 7527 1006 7567 1042
rect 7527 974 7531 1006
rect 7531 974 7563 1006
rect 7563 974 7567 1006
rect 7527 938 7567 974
rect 7527 906 7531 938
rect 7531 906 7563 938
rect 7563 906 7567 938
rect 7527 870 7567 906
rect 7527 838 7531 870
rect 7531 838 7563 870
rect 7563 838 7567 870
rect 7527 802 7567 838
rect 7527 770 7531 802
rect 7531 770 7563 802
rect 7563 770 7567 802
rect 7527 734 7567 770
rect 7527 702 7531 734
rect 7531 702 7563 734
rect 7563 702 7567 734
rect 7527 666 7567 702
rect 7527 634 7531 666
rect 7531 634 7563 666
rect 7563 634 7567 666
rect 7527 598 7567 634
rect 7527 566 7531 598
rect 7531 566 7563 598
rect 7563 566 7567 598
rect 7527 560 7567 566
rect 7788 1414 7910 1420
rect 7788 1382 7833 1414
rect 7833 1382 7865 1414
rect 7865 1382 7910 1414
rect 7788 1346 7910 1382
rect 7788 1314 7833 1346
rect 7833 1314 7865 1346
rect 7865 1314 7910 1346
rect 7788 1278 7910 1314
rect 7788 1246 7833 1278
rect 7833 1246 7865 1278
rect 7865 1246 7910 1278
rect 7788 1210 7910 1246
rect 7788 1178 7833 1210
rect 7833 1178 7865 1210
rect 7865 1178 7910 1210
rect 7788 1142 7910 1178
rect 7788 1110 7833 1142
rect 7833 1110 7865 1142
rect 7865 1110 7910 1142
rect 7788 1074 7910 1110
rect 7788 1042 7833 1074
rect 7833 1042 7865 1074
rect 7865 1042 7910 1074
rect 7788 1006 7910 1042
rect 7788 974 7833 1006
rect 7833 974 7865 1006
rect 7865 974 7910 1006
rect 7788 938 7910 974
rect 7788 906 7833 938
rect 7833 906 7865 938
rect 7865 906 7910 938
rect 7788 870 7910 906
rect 7788 838 7833 870
rect 7833 838 7865 870
rect 7865 838 7910 870
rect 7788 802 7910 838
rect 7788 770 7833 802
rect 7833 770 7865 802
rect 7865 770 7910 802
rect 7788 734 7910 770
rect 7788 702 7833 734
rect 7833 702 7865 734
rect 7865 702 7910 734
rect 7788 666 7910 702
rect 7788 634 7833 666
rect 7833 634 7865 666
rect 7865 634 7910 666
rect 7788 598 7910 634
rect 7788 566 7833 598
rect 7833 566 7865 598
rect 7865 566 7910 598
rect 7788 560 7910 566
rect 8131 1414 8171 1420
rect 8131 1382 8135 1414
rect 8135 1382 8167 1414
rect 8167 1382 8171 1414
rect 8131 1346 8171 1382
rect 8131 1314 8135 1346
rect 8135 1314 8167 1346
rect 8167 1314 8171 1346
rect 8131 1278 8171 1314
rect 8131 1246 8135 1278
rect 8135 1246 8167 1278
rect 8167 1246 8171 1278
rect 8131 1210 8171 1246
rect 8131 1178 8135 1210
rect 8135 1178 8167 1210
rect 8167 1178 8171 1210
rect 8131 1142 8171 1178
rect 8131 1110 8135 1142
rect 8135 1110 8167 1142
rect 8167 1110 8171 1142
rect 8131 1074 8171 1110
rect 8131 1042 8135 1074
rect 8135 1042 8167 1074
rect 8167 1042 8171 1074
rect 8131 1006 8171 1042
rect 8131 974 8135 1006
rect 8135 974 8167 1006
rect 8167 974 8171 1006
rect 8131 938 8171 974
rect 8131 906 8135 938
rect 8135 906 8167 938
rect 8167 906 8171 938
rect 8131 870 8171 906
rect 8131 838 8135 870
rect 8135 838 8167 870
rect 8167 838 8171 870
rect 8131 802 8171 838
rect 8131 770 8135 802
rect 8135 770 8167 802
rect 8167 770 8171 802
rect 8131 734 8171 770
rect 8131 702 8135 734
rect 8135 702 8167 734
rect 8167 702 8171 734
rect 8131 666 8171 702
rect 8131 634 8135 666
rect 8135 634 8167 666
rect 8167 634 8171 666
rect 8131 598 8171 634
rect 8131 566 8135 598
rect 8135 566 8167 598
rect 8167 566 8171 598
rect 8131 560 8171 566
rect 8392 1414 8514 1420
rect 8392 1382 8437 1414
rect 8437 1382 8469 1414
rect 8469 1382 8514 1414
rect 8392 1346 8514 1382
rect 8392 1314 8437 1346
rect 8437 1314 8469 1346
rect 8469 1314 8514 1346
rect 8392 1278 8514 1314
rect 8392 1246 8437 1278
rect 8437 1246 8469 1278
rect 8469 1246 8514 1278
rect 8392 1210 8514 1246
rect 8392 1178 8437 1210
rect 8437 1178 8469 1210
rect 8469 1178 8514 1210
rect 8392 1142 8514 1178
rect 8392 1110 8437 1142
rect 8437 1110 8469 1142
rect 8469 1110 8514 1142
rect 8392 1074 8514 1110
rect 8392 1042 8437 1074
rect 8437 1042 8469 1074
rect 8469 1042 8514 1074
rect 8392 1006 8514 1042
rect 8392 974 8437 1006
rect 8437 974 8469 1006
rect 8469 974 8514 1006
rect 8392 938 8514 974
rect 8392 906 8437 938
rect 8437 906 8469 938
rect 8469 906 8514 938
rect 8392 870 8514 906
rect 8392 838 8437 870
rect 8437 838 8469 870
rect 8469 838 8514 870
rect 8392 802 8514 838
rect 8392 770 8437 802
rect 8437 770 8469 802
rect 8469 770 8514 802
rect 8392 734 8514 770
rect 8392 702 8437 734
rect 8437 702 8469 734
rect 8469 702 8514 734
rect 8392 666 8514 702
rect 8392 634 8437 666
rect 8437 634 8469 666
rect 8469 634 8514 666
rect 8392 598 8514 634
rect 8392 566 8437 598
rect 8437 566 8469 598
rect 8469 566 8514 598
rect 8392 560 8514 566
rect 8735 1414 8775 1420
rect 8735 1382 8739 1414
rect 8739 1382 8771 1414
rect 8771 1382 8775 1414
rect 8735 1346 8775 1382
rect 8735 1314 8739 1346
rect 8739 1314 8771 1346
rect 8771 1314 8775 1346
rect 8735 1278 8775 1314
rect 8735 1246 8739 1278
rect 8739 1246 8771 1278
rect 8771 1246 8775 1278
rect 8735 1210 8775 1246
rect 8735 1178 8739 1210
rect 8739 1178 8771 1210
rect 8771 1178 8775 1210
rect 8735 1142 8775 1178
rect 8735 1110 8739 1142
rect 8739 1110 8771 1142
rect 8771 1110 8775 1142
rect 8735 1074 8775 1110
rect 8735 1042 8739 1074
rect 8739 1042 8771 1074
rect 8771 1042 8775 1074
rect 8735 1006 8775 1042
rect 8735 974 8739 1006
rect 8739 974 8771 1006
rect 8771 974 8775 1006
rect 8735 938 8775 974
rect 8735 906 8739 938
rect 8739 906 8771 938
rect 8771 906 8775 938
rect 8735 870 8775 906
rect 8735 838 8739 870
rect 8739 838 8771 870
rect 8771 838 8775 870
rect 8735 802 8775 838
rect 8735 770 8739 802
rect 8739 770 8771 802
rect 8771 770 8775 802
rect 8735 734 8775 770
rect 8735 702 8739 734
rect 8739 702 8771 734
rect 8771 702 8775 734
rect 8735 666 8775 702
rect 8735 634 8739 666
rect 8739 634 8771 666
rect 8771 634 8775 666
rect 8735 598 8775 634
rect 8735 566 8739 598
rect 8739 566 8771 598
rect 8771 566 8775 598
rect 8735 560 8775 566
rect 8996 1414 9118 1420
rect 8996 1382 9041 1414
rect 9041 1382 9073 1414
rect 9073 1382 9118 1414
rect 8996 1346 9118 1382
rect 8996 1314 9041 1346
rect 9041 1314 9073 1346
rect 9073 1314 9118 1346
rect 8996 1278 9118 1314
rect 8996 1246 9041 1278
rect 9041 1246 9073 1278
rect 9073 1246 9118 1278
rect 8996 1210 9118 1246
rect 8996 1178 9041 1210
rect 9041 1178 9073 1210
rect 9073 1178 9118 1210
rect 8996 1142 9118 1178
rect 8996 1110 9041 1142
rect 9041 1110 9073 1142
rect 9073 1110 9118 1142
rect 8996 1074 9118 1110
rect 8996 1042 9041 1074
rect 9041 1042 9073 1074
rect 9073 1042 9118 1074
rect 8996 1006 9118 1042
rect 8996 974 9041 1006
rect 9041 974 9073 1006
rect 9073 974 9118 1006
rect 8996 938 9118 974
rect 8996 906 9041 938
rect 9041 906 9073 938
rect 9073 906 9118 938
rect 8996 870 9118 906
rect 8996 838 9041 870
rect 9041 838 9073 870
rect 9073 838 9118 870
rect 8996 802 9118 838
rect 8996 770 9041 802
rect 9041 770 9073 802
rect 9073 770 9118 802
rect 8996 734 9118 770
rect 8996 702 9041 734
rect 9041 702 9073 734
rect 9073 702 9118 734
rect 8996 666 9118 702
rect 8996 634 9041 666
rect 9041 634 9073 666
rect 9073 634 9118 666
rect 8996 598 9118 634
rect 8996 566 9041 598
rect 9041 566 9073 598
rect 9073 566 9118 598
rect 8996 560 9118 566
rect 9339 1414 9379 1420
rect 9339 1382 9343 1414
rect 9343 1382 9375 1414
rect 9375 1382 9379 1414
rect 9339 1346 9379 1382
rect 9339 1314 9343 1346
rect 9343 1314 9375 1346
rect 9375 1314 9379 1346
rect 9339 1278 9379 1314
rect 9339 1246 9343 1278
rect 9343 1246 9375 1278
rect 9375 1246 9379 1278
rect 9339 1210 9379 1246
rect 9339 1178 9343 1210
rect 9343 1178 9375 1210
rect 9375 1178 9379 1210
rect 9339 1142 9379 1178
rect 9339 1110 9343 1142
rect 9343 1110 9375 1142
rect 9375 1110 9379 1142
rect 9339 1074 9379 1110
rect 9339 1042 9343 1074
rect 9343 1042 9375 1074
rect 9375 1042 9379 1074
rect 9339 1006 9379 1042
rect 9339 974 9343 1006
rect 9343 974 9375 1006
rect 9375 974 9379 1006
rect 9339 938 9379 974
rect 9339 906 9343 938
rect 9343 906 9375 938
rect 9375 906 9379 938
rect 9339 870 9379 906
rect 9339 838 9343 870
rect 9343 838 9375 870
rect 9375 838 9379 870
rect 9339 802 9379 838
rect 9339 770 9343 802
rect 9343 770 9375 802
rect 9375 770 9379 802
rect 9339 734 9379 770
rect 9339 702 9343 734
rect 9343 702 9375 734
rect 9375 702 9379 734
rect 9339 666 9379 702
rect 9339 634 9343 666
rect 9343 634 9375 666
rect 9375 634 9379 666
rect 9339 598 9379 634
rect 9339 566 9343 598
rect 9343 566 9375 598
rect 9375 566 9379 598
rect 9339 560 9379 566
rect 9600 1414 9722 1420
rect 9600 1382 9645 1414
rect 9645 1382 9677 1414
rect 9677 1382 9722 1414
rect 9600 1346 9722 1382
rect 9600 1314 9645 1346
rect 9645 1314 9677 1346
rect 9677 1314 9722 1346
rect 9600 1278 9722 1314
rect 9600 1246 9645 1278
rect 9645 1246 9677 1278
rect 9677 1246 9722 1278
rect 9600 1210 9722 1246
rect 9600 1178 9645 1210
rect 9645 1178 9677 1210
rect 9677 1178 9722 1210
rect 9600 1142 9722 1178
rect 9600 1110 9645 1142
rect 9645 1110 9677 1142
rect 9677 1110 9722 1142
rect 9600 1074 9722 1110
rect 9600 1042 9645 1074
rect 9645 1042 9677 1074
rect 9677 1042 9722 1074
rect 9600 1006 9722 1042
rect 9600 974 9645 1006
rect 9645 974 9677 1006
rect 9677 974 9722 1006
rect 9600 938 9722 974
rect 9600 906 9645 938
rect 9645 906 9677 938
rect 9677 906 9722 938
rect 9600 870 9722 906
rect 9600 838 9645 870
rect 9645 838 9677 870
rect 9677 838 9722 870
rect 9600 802 9722 838
rect 9600 770 9645 802
rect 9645 770 9677 802
rect 9677 770 9722 802
rect 9600 734 9722 770
rect 9600 702 9645 734
rect 9645 702 9677 734
rect 9677 702 9722 734
rect 9600 666 9722 702
rect 9600 634 9645 666
rect 9645 634 9677 666
rect 9677 634 9722 666
rect 9600 598 9722 634
rect 9600 566 9645 598
rect 9645 566 9677 598
rect 9677 566 9722 598
rect 9600 560 9722 566
rect 9943 1414 9983 1420
rect 9943 1382 9947 1414
rect 9947 1382 9979 1414
rect 9979 1382 9983 1414
rect 9943 1346 9983 1382
rect 9943 1314 9947 1346
rect 9947 1314 9979 1346
rect 9979 1314 9983 1346
rect 9943 1278 9983 1314
rect 9943 1246 9947 1278
rect 9947 1246 9979 1278
rect 9979 1246 9983 1278
rect 9943 1210 9983 1246
rect 9943 1178 9947 1210
rect 9947 1178 9979 1210
rect 9979 1178 9983 1210
rect 9943 1142 9983 1178
rect 9943 1110 9947 1142
rect 9947 1110 9979 1142
rect 9979 1110 9983 1142
rect 9943 1074 9983 1110
rect 9943 1042 9947 1074
rect 9947 1042 9979 1074
rect 9979 1042 9983 1074
rect 9943 1006 9983 1042
rect 9943 974 9947 1006
rect 9947 974 9979 1006
rect 9979 974 9983 1006
rect 9943 938 9983 974
rect 9943 906 9947 938
rect 9947 906 9979 938
rect 9979 906 9983 938
rect 9943 870 9983 906
rect 9943 838 9947 870
rect 9947 838 9979 870
rect 9979 838 9983 870
rect 9943 802 9983 838
rect 9943 770 9947 802
rect 9947 770 9979 802
rect 9979 770 9983 802
rect 9943 734 9983 770
rect 9943 702 9947 734
rect 9947 702 9979 734
rect 9979 702 9983 734
rect 9943 666 9983 702
rect 9943 634 9947 666
rect 9947 634 9979 666
rect 9979 634 9983 666
rect 9943 598 9983 634
rect 9943 566 9947 598
rect 9947 566 9979 598
rect 9979 566 9983 598
rect 9943 560 9983 566
rect 10204 1414 10326 1420
rect 10204 1382 10249 1414
rect 10249 1382 10281 1414
rect 10281 1382 10326 1414
rect 10204 1346 10326 1382
rect 10204 1314 10249 1346
rect 10249 1314 10281 1346
rect 10281 1314 10326 1346
rect 10204 1278 10326 1314
rect 10204 1246 10249 1278
rect 10249 1246 10281 1278
rect 10281 1246 10326 1278
rect 10204 1210 10326 1246
rect 10204 1178 10249 1210
rect 10249 1178 10281 1210
rect 10281 1178 10326 1210
rect 10204 1142 10326 1178
rect 10204 1110 10249 1142
rect 10249 1110 10281 1142
rect 10281 1110 10326 1142
rect 10204 1074 10326 1110
rect 10204 1042 10249 1074
rect 10249 1042 10281 1074
rect 10281 1042 10326 1074
rect 10204 1006 10326 1042
rect 10204 974 10249 1006
rect 10249 974 10281 1006
rect 10281 974 10326 1006
rect 10204 938 10326 974
rect 10204 906 10249 938
rect 10249 906 10281 938
rect 10281 906 10326 938
rect 10204 870 10326 906
rect 10204 838 10249 870
rect 10249 838 10281 870
rect 10281 838 10326 870
rect 10204 802 10326 838
rect 10204 770 10249 802
rect 10249 770 10281 802
rect 10281 770 10326 802
rect 10204 734 10326 770
rect 10204 702 10249 734
rect 10249 702 10281 734
rect 10281 702 10326 734
rect 10204 666 10326 702
rect 10204 634 10249 666
rect 10249 634 10281 666
rect 10281 634 10326 666
rect 10204 598 10326 634
rect 10204 566 10249 598
rect 10249 566 10281 598
rect 10281 566 10326 598
rect 10204 560 10326 566
rect 5715 410 5755 414
rect 6319 410 6359 414
rect 6923 410 6963 414
rect 7527 410 7567 414
rect 8131 410 8171 414
rect 8735 410 8775 414
rect 9339 410 9379 414
rect 9943 410 9983 414
rect 5715 378 5738 410
rect 5738 378 5755 410
rect 6319 378 6350 410
rect 6350 378 6359 410
rect 6923 378 6930 410
rect 6930 378 6962 410
rect 6962 378 6963 410
rect 7527 378 7542 410
rect 7542 378 7567 410
rect 8131 378 8154 410
rect 8154 378 8171 410
rect 8735 378 8766 410
rect 8766 378 8775 410
rect 9339 378 9342 410
rect 9342 378 9378 410
rect 9378 378 9379 410
rect 9943 378 9954 410
rect 9954 378 9983 410
rect 5715 374 5755 378
rect 6319 374 6359 378
rect 6923 374 6963 378
rect 7527 374 7567 378
rect 8131 374 8171 378
rect 8735 374 8775 378
rect 9339 374 9379 378
rect 9943 374 9983 378
<< metal2 >>
rect 3046 1464 3086 1980
rect 3046 1333 3086 1342
rect 5715 1953 5755 1980
rect 5976 1420 6098 1980
rect 5976 551 6098 560
rect 6319 1953 6359 1980
rect 5715 0 5755 27
rect 6580 1420 6702 1980
rect 6580 551 6702 560
rect 6923 1953 6963 1980
rect 6319 0 6359 27
rect 7184 1420 7306 1980
rect 7184 551 7306 560
rect 7527 1953 7567 1980
rect 6923 0 6963 27
rect 7788 1420 7910 1980
rect 7788 551 7910 560
rect 8131 1953 8171 1980
rect 7527 0 7567 27
rect 8392 1420 8514 1980
rect 8392 551 8514 560
rect 8735 1953 8775 1980
rect 8131 0 8171 27
rect 8996 1420 9118 1980
rect 8996 551 9118 560
rect 9339 1953 9379 1980
rect 8735 0 8775 27
rect 9600 1420 9722 1980
rect 9600 551 9722 560
rect 9943 1953 9983 1980
rect 9339 0 9379 27
rect 10204 1420 10326 1980
rect 10204 551 10326 560
rect 9943 0 9983 27
<< via2 >>
rect 5715 1606 5755 1953
rect 5715 1566 5755 1606
rect 5715 1420 5755 1566
rect 5715 560 5755 1420
rect 5715 414 5755 560
rect 6319 1606 6359 1953
rect 6319 1566 6359 1606
rect 6319 1420 6359 1566
rect 6319 560 6359 1420
rect 5715 374 5755 414
rect 5715 27 5755 374
rect 6319 414 6359 560
rect 6923 1606 6963 1953
rect 6923 1566 6963 1606
rect 6923 1420 6963 1566
rect 6923 560 6963 1420
rect 6319 374 6359 414
rect 6319 27 6359 374
rect 6923 414 6963 560
rect 7527 1606 7567 1953
rect 7527 1566 7567 1606
rect 7527 1420 7567 1566
rect 7527 560 7567 1420
rect 6923 374 6963 414
rect 6923 27 6963 374
rect 7527 414 7567 560
rect 8131 1606 8171 1953
rect 8131 1566 8171 1606
rect 8131 1420 8171 1566
rect 8131 560 8171 1420
rect 7527 374 7567 414
rect 7527 27 7567 374
rect 8131 414 8171 560
rect 8735 1606 8775 1953
rect 8735 1566 8775 1606
rect 8735 1420 8775 1566
rect 8735 560 8775 1420
rect 8131 374 8171 414
rect 8131 27 8171 374
rect 8735 414 8775 560
rect 9339 1606 9379 1953
rect 9339 1566 9379 1606
rect 9339 1420 9379 1566
rect 9339 560 9379 1420
rect 8735 374 8775 414
rect 8735 27 8775 374
rect 9339 414 9379 560
rect 9943 1606 9983 1953
rect 9943 1566 9983 1606
rect 9943 1420 9983 1566
rect 9943 560 9983 1420
rect 9339 374 9379 414
rect 9339 27 9379 374
rect 9943 414 9983 560
rect 9943 374 9983 414
rect 9943 27 9983 374
<< metal3 >>
rect 5715 1953 5755 1962
rect 5715 18 5755 27
rect 6319 1953 6359 1962
rect 6319 18 6359 27
rect 6923 1953 6963 1962
rect 6923 18 6963 27
rect 7527 1953 7567 1962
rect 7527 18 7567 27
rect 8131 1953 8171 1962
rect 8131 18 8171 27
rect 8735 1953 8775 1962
rect 8735 18 8775 27
rect 9339 1953 9379 1962
rect 9339 18 9379 27
rect 9943 1953 9983 1962
rect 9943 18 9983 27
<< labels >>
flabel metal2 s 10204 551 10326 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 9600 551 9722 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 8996 551 9118 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 8392 551 8514 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 7788 551 7910 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 6580 551 6702 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 7184 551 7306 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
rlabel metal2 s 3046 1333 3086 1980 4 gate
port 3 nsew
rlabel metal2 s 5976 551 6098 1980 4 pad
port 2 nsew
rlabel comment s 394 394 394 394 4 sub!
flabel comment s 3064 1341 3064 1341 0 FreeSans 400 0 0 0 dant
flabel metal1 s 485 1556 801 1613 0 FreeSans 51 0 0 0 iovss
port 1 nsew
<< properties >>
string device primitive
string GDS_END 26431256
string GDS_FILE sg13g2_io.gds
string GDS_START 26313724
<< end >>
