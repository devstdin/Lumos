magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756676971
<< error_p >>
rect -67745 131856 135535 132116
rect -67745 131276 -67485 131856
rect -68585 131016 -67485 131276
rect -67453 131564 135243 131824
rect -68585 130436 -68325 131016
rect -67453 130984 -67193 131564
rect -69425 130176 -68325 130436
rect -68293 130724 -67193 130984
rect 134983 130984 135243 131564
rect 135275 131276 135535 131856
rect 135275 131016 136375 131276
rect 134983 130724 136083 130984
rect -69425 129596 -69165 130176
rect -68293 130144 -68033 130724
rect -70265 129336 -69165 129596
rect -69133 129884 -68033 130144
rect 135823 130144 136083 130724
rect 136115 130436 136375 131016
rect 136115 130176 137215 130436
rect 135823 129884 136923 130144
rect -70265 128756 -70005 129336
rect -69133 129304 -68873 129884
rect -71105 128496 -70005 128756
rect -69973 129044 -68873 129304
rect 136663 129304 136923 129884
rect 136955 129596 137215 130176
rect 136955 129336 138055 129596
rect 136663 129044 137763 129304
rect -71105 -58264 -70845 128496
rect -69973 128464 -69713 129044
rect -70813 128204 -69713 128464
rect 137503 128464 137763 129044
rect 137795 128756 138055 129336
rect 137795 128496 138895 128756
rect 137503 128204 138603 128464
rect -70813 -57972 -70553 128204
rect 138343 -57972 138603 128204
rect -70813 -58232 -69713 -57972
rect -71105 -58524 -70005 -58264
rect -70265 -59104 -70005 -58524
rect -69973 -58812 -69713 -58232
rect 137503 -58232 138603 -57972
rect 137503 -58812 137763 -58232
rect 138635 -58264 138895 128496
rect -69973 -59072 -68873 -58812
rect -70265 -59364 -69165 -59104
rect -69425 -59944 -69165 -59364
rect -69133 -59652 -68873 -59072
rect 136663 -59072 137763 -58812
rect 137795 -58524 138895 -58264
rect 136663 -59652 136923 -59072
rect 137795 -59104 138055 -58524
rect -69133 -59912 -68033 -59652
rect -69425 -60204 -68325 -59944
rect -68585 -60784 -68325 -60204
rect -68293 -60492 -68033 -59912
rect 135823 -59912 136923 -59652
rect 136955 -59364 138055 -59104
rect 135823 -60492 136083 -59912
rect 136955 -59944 137215 -59364
rect -68293 -60752 -67193 -60492
rect -68585 -61044 -67485 -60784
rect -67745 -61624 -67485 -61044
rect -67453 -61332 -67193 -60752
rect 134983 -60752 136083 -60492
rect 136115 -60204 137215 -59944
rect 134983 -61332 135243 -60752
rect 136115 -60784 136375 -60204
rect -67453 -61592 135243 -61332
rect 135275 -61044 136375 -60784
rect 135275 -61624 135535 -61044
rect -67745 -61884 135535 -61624
<< sealcont >>
rect -67485 131824 135275 131856
rect -67485 131016 -67453 131824
rect -68325 130984 -67453 131016
rect 135243 131016 135275 131824
rect 135243 130984 136115 131016
rect -68325 130176 -68293 130984
rect -69165 130144 -68293 130176
rect 136083 130176 136115 130984
rect 136083 130144 136955 130176
rect -69165 129336 -69133 130144
rect -70005 129304 -69133 129336
rect 136923 129336 136955 130144
rect 136923 129304 137795 129336
rect -70005 128496 -69973 129304
rect -70845 128464 -69973 128496
rect 137763 128496 137795 129304
rect 137763 128464 138635 128496
rect -70845 -58232 -70813 128464
rect 138603 -58232 138635 128464
rect -70845 -58264 -69973 -58232
rect -70005 -59072 -69973 -58264
rect 137763 -58264 138635 -58232
rect 137763 -59072 137795 -58264
rect -70005 -59104 -69133 -59072
rect -69165 -59912 -69133 -59104
rect 136923 -59104 137795 -59072
rect 136923 -59912 136955 -59104
rect -69165 -59944 -68293 -59912
rect -68325 -60752 -68293 -59944
rect 136083 -59944 136955 -59912
rect 136083 -60752 136115 -59944
rect -68325 -60784 -67453 -60752
rect -67485 -61592 -67453 -60784
rect 135243 -60784 136115 -60752
rect 135243 -61592 135275 -60784
rect -67485 -61624 135275 -61592
<< metal1 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67447 131416 135237 131818
rect -68725 130576 -68325 131016
rect -67447 130978 -67045 131416
rect -69565 130176 -68325 130576
rect -68287 130576 -67045 130978
rect 134835 130978 135237 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 136077 130978
rect -69565 129736 -69165 130176
rect -68287 130138 -67885 130576
rect -70405 129336 -69165 129736
rect -69127 129736 -67885 130138
rect 135675 130138 136077 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136917 130138
rect -70405 128896 -70005 129336
rect -69127 129298 -68725 129736
rect -71245 128496 -70005 128896
rect -69967 128896 -68725 129298
rect 136515 129298 136917 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137757 129298
rect -71245 -58264 -70845 128496
rect -69967 128458 -69565 128896
rect -70807 128056 -69565 128458
rect 137355 128458 137757 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138597 128458
rect -70807 -57824 -70405 128056
rect 138195 -57824 138597 128056
rect -70807 -58226 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69967 -58664 -69565 -58226
rect 137355 -58226 138597 -57824
rect 137355 -58664 137757 -58226
rect 138635 -58264 139035 128496
rect -69967 -59066 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -69127 -59504 -68725 -59066
rect 136515 -59066 137757 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136917 -59066
rect 137795 -59104 138195 -58664
rect -69127 -59906 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68287 -60344 -67885 -59906
rect 135675 -59906 136917 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 136077 -59906
rect 136955 -59944 137355 -59504
rect -68287 -60746 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67447 -61184 -67045 -60746
rect 134835 -60746 136077 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135237 -60746
rect 136115 -60784 136515 -60344
rect -67447 -61586 135237 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia1 >>
rect -67485 131818 135275 131856
rect -67485 131016 -67447 131818
rect -68325 130978 -67447 131016
rect -68325 130176 -68287 130978
rect 135237 131016 135275 131818
rect 135237 130978 136115 131016
rect -69165 130138 -68287 130176
rect -69165 129336 -69127 130138
rect 136077 130176 136115 130978
rect 136077 130138 136955 130176
rect -70005 129298 -69127 129336
rect -70005 128496 -69967 129298
rect 136917 129336 136955 130138
rect 136917 129298 137795 129336
rect -70845 128458 -69967 128496
rect -70845 -58226 -70807 128458
rect 137757 128496 137795 129298
rect 137757 128458 138635 128496
rect -70845 -58264 -69967 -58226
rect -70005 -59066 -69967 -58264
rect 138597 -58226 138635 128458
rect 137757 -58264 138635 -58226
rect -70005 -59104 -69127 -59066
rect -69165 -59906 -69127 -59104
rect 137757 -59066 137795 -58264
rect 136917 -59104 137795 -59066
rect -69165 -59944 -68287 -59906
rect -68325 -60746 -68287 -59944
rect 136917 -59906 136955 -59104
rect 136077 -59944 136955 -59906
rect -68325 -60784 -67447 -60746
rect -67485 -61586 -67447 -60784
rect 136077 -60746 136115 -59944
rect 135237 -60784 136115 -60746
rect 135237 -61586 135275 -60784
rect -67485 -61624 135275 -61586
<< metal2 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67447 131416 135237 131818
rect -68725 130576 -68325 131016
rect -67447 130978 -67045 131416
rect -69565 130176 -68325 130576
rect -68287 130576 -67045 130978
rect 134835 130978 135237 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 136077 130978
rect -69565 129736 -69165 130176
rect -68287 130138 -67885 130576
rect -70405 129336 -69165 129736
rect -69127 129736 -67885 130138
rect 135675 130138 136077 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136917 130138
rect -70405 128896 -70005 129336
rect -69127 129298 -68725 129736
rect -71245 128496 -70005 128896
rect -69967 128896 -68725 129298
rect 136515 129298 136917 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137757 129298
rect -71245 -58264 -70845 128496
rect -69967 128458 -69565 128896
rect -70807 128056 -69565 128458
rect 137355 128458 137757 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138597 128458
rect -70807 -57824 -70405 128056
rect 138195 -57824 138597 128056
rect -70807 -58226 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69967 -58664 -69565 -58226
rect 137355 -58226 138597 -57824
rect 137355 -58664 137757 -58226
rect 138635 -58264 139035 128496
rect -69967 -59066 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -69127 -59504 -68725 -59066
rect 136515 -59066 137757 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136917 -59066
rect 137795 -59104 138195 -58664
rect -69127 -59906 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68287 -60344 -67885 -59906
rect 135675 -59906 136917 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 136077 -59906
rect 136955 -59944 137355 -59504
rect -68287 -60746 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67447 -61184 -67045 -60746
rect 134835 -60746 136077 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135237 -60746
rect 136115 -60784 136515 -60344
rect -67447 -61586 135237 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia2 >>
rect -67485 131818 135275 131856
rect -67485 131016 -67447 131818
rect -68325 130978 -67447 131016
rect -68325 130176 -68287 130978
rect 135237 131016 135275 131818
rect 135237 130978 136115 131016
rect -69165 130138 -68287 130176
rect -69165 129336 -69127 130138
rect 136077 130176 136115 130978
rect 136077 130138 136955 130176
rect -70005 129298 -69127 129336
rect -70005 128496 -69967 129298
rect 136917 129336 136955 130138
rect 136917 129298 137795 129336
rect -70845 128458 -69967 128496
rect -70845 -58226 -70807 128458
rect 137757 128496 137795 129298
rect 137757 128458 138635 128496
rect -70845 -58264 -69967 -58226
rect -70005 -59066 -69967 -58264
rect 138597 -58226 138635 128458
rect 137757 -58264 138635 -58226
rect -70005 -59104 -69127 -59066
rect -69165 -59906 -69127 -59104
rect 137757 -59066 137795 -58264
rect 136917 -59104 137795 -59066
rect -69165 -59944 -68287 -59906
rect -68325 -60746 -68287 -59944
rect 136917 -59906 136955 -59104
rect 136077 -59944 136955 -59906
rect -68325 -60784 -67447 -60746
rect -67485 -61586 -67447 -60784
rect 136077 -60746 136115 -59944
rect 135237 -60784 136115 -60746
rect 135237 -61586 135275 -60784
rect -67485 -61624 135275 -61586
<< metal3 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67447 131416 135237 131818
rect -68725 130576 -68325 131016
rect -67447 130978 -67045 131416
rect -69565 130176 -68325 130576
rect -68287 130576 -67045 130978
rect 134835 130978 135237 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 136077 130978
rect -69565 129736 -69165 130176
rect -68287 130138 -67885 130576
rect -70405 129336 -69165 129736
rect -69127 129736 -67885 130138
rect 135675 130138 136077 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136917 130138
rect -70405 128896 -70005 129336
rect -69127 129298 -68725 129736
rect -71245 128496 -70005 128896
rect -69967 128896 -68725 129298
rect 136515 129298 136917 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137757 129298
rect -71245 -58264 -70845 128496
rect -69967 128458 -69565 128896
rect -70807 128056 -69565 128458
rect 137355 128458 137757 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138597 128458
rect -70807 -57824 -70405 128056
rect 138195 -57824 138597 128056
rect -70807 -58226 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69967 -58664 -69565 -58226
rect 137355 -58226 138597 -57824
rect 137355 -58664 137757 -58226
rect 138635 -58264 139035 128496
rect -69967 -59066 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -69127 -59504 -68725 -59066
rect 136515 -59066 137757 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136917 -59066
rect 137795 -59104 138195 -58664
rect -69127 -59906 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68287 -60344 -67885 -59906
rect 135675 -59906 136917 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 136077 -59906
rect 136955 -59944 137355 -59504
rect -68287 -60746 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67447 -61184 -67045 -60746
rect 134835 -60746 136077 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135237 -60746
rect 136115 -60784 136515 -60344
rect -67447 -61586 135237 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia3 >>
rect -67485 131818 135275 131856
rect -67485 131016 -67447 131818
rect -68325 130978 -67447 131016
rect -68325 130176 -68287 130978
rect 135237 131016 135275 131818
rect 135237 130978 136115 131016
rect -69165 130138 -68287 130176
rect -69165 129336 -69127 130138
rect 136077 130176 136115 130978
rect 136077 130138 136955 130176
rect -70005 129298 -69127 129336
rect -70005 128496 -69967 129298
rect 136917 129336 136955 130138
rect 136917 129298 137795 129336
rect -70845 128458 -69967 128496
rect -70845 -58226 -70807 128458
rect 137757 128496 137795 129298
rect 137757 128458 138635 128496
rect -70845 -58264 -69967 -58226
rect -70005 -59066 -69967 -58264
rect 138597 -58226 138635 128458
rect 137757 -58264 138635 -58226
rect -70005 -59104 -69127 -59066
rect -69165 -59906 -69127 -59104
rect 137757 -59066 137795 -58264
rect 136917 -59104 137795 -59066
rect -69165 -59944 -68287 -59906
rect -68325 -60746 -68287 -59944
rect 136917 -59906 136955 -59104
rect 136077 -59944 136955 -59906
rect -68325 -60784 -67447 -60746
rect -67485 -61586 -67447 -60784
rect 136077 -60746 136115 -59944
rect 135237 -60784 136115 -60746
rect 135237 -61586 135275 -60784
rect -67485 -61624 135275 -61586
<< metal4 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67447 131416 135237 131818
rect -68725 130576 -68325 131016
rect -67447 130978 -67045 131416
rect -69565 130176 -68325 130576
rect -68287 130576 -67045 130978
rect 134835 130978 135237 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 136077 130978
rect -69565 129736 -69165 130176
rect -68287 130138 -67885 130576
rect -70405 129336 -69165 129736
rect -69127 129736 -67885 130138
rect 135675 130138 136077 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136917 130138
rect -70405 128896 -70005 129336
rect -69127 129298 -68725 129736
rect -71245 128496 -70005 128896
rect -69967 128896 -68725 129298
rect 136515 129298 136917 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137757 129298
rect -71245 -58264 -70845 128496
rect -69967 128458 -69565 128896
rect -70807 128056 -69565 128458
rect 137355 128458 137757 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138597 128458
rect -70807 -57824 -70405 128056
rect 138195 -57824 138597 128056
rect -70807 -58226 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69967 -58664 -69565 -58226
rect 137355 -58226 138597 -57824
rect 137355 -58664 137757 -58226
rect 138635 -58264 139035 128496
rect -69967 -59066 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -69127 -59504 -68725 -59066
rect 136515 -59066 137757 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136917 -59066
rect 137795 -59104 138195 -58664
rect -69127 -59906 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68287 -60344 -67885 -59906
rect 135675 -59906 136917 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 136077 -59906
rect 136955 -59944 137355 -59504
rect -68287 -60746 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67447 -61184 -67045 -60746
rect 134835 -60746 136077 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135237 -60746
rect 136115 -60784 136515 -60344
rect -67447 -61586 135237 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia4 >>
rect -67485 131818 135275 131856
rect -67485 131016 -67447 131818
rect -68325 130978 -67447 131016
rect -68325 130176 -68287 130978
rect 135237 131016 135275 131818
rect 135237 130978 136115 131016
rect -69165 130138 -68287 130176
rect -69165 129336 -69127 130138
rect 136077 130176 136115 130978
rect 136077 130138 136955 130176
rect -70005 129298 -69127 129336
rect -70005 128496 -69967 129298
rect 136917 129336 136955 130138
rect 136917 129298 137795 129336
rect -70845 128458 -69967 128496
rect -70845 -58226 -70807 128458
rect 137757 128496 137795 129298
rect 137757 128458 138635 128496
rect -70845 -58264 -69967 -58226
rect -70005 -59066 -69967 -58264
rect 138597 -58226 138635 128458
rect 137757 -58264 138635 -58226
rect -70005 -59104 -69127 -59066
rect -69165 -59906 -69127 -59104
rect 137757 -59066 137795 -58264
rect 136917 -59104 137795 -59066
rect -69165 -59944 -68287 -59906
rect -68325 -60746 -68287 -59944
rect 136917 -59906 136955 -59104
rect 136077 -59944 136955 -59906
rect -68325 -60784 -67447 -60746
rect -67485 -61586 -67447 -60784
rect 136077 -60746 136115 -59944
rect 135237 -60784 136115 -60746
rect 135237 -61586 135275 -60784
rect -67485 -61624 135275 -61586
<< metal5 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67401 131416 135191 131772
rect -68725 130576 -68325 131016
rect -67401 130932 -67045 131416
rect -69565 130176 -68325 130576
rect -68241 130576 -67045 130932
rect 134835 130932 135191 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 136031 130932
rect -69565 129736 -69165 130176
rect -68241 130092 -67885 130576
rect -70405 129336 -69165 129736
rect -69081 129736 -67885 130092
rect 135675 130092 136031 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136871 130092
rect -70405 128896 -70005 129336
rect -69081 129252 -68725 129736
rect -71245 128496 -70005 128896
rect -69921 128896 -68725 129252
rect 136515 129252 136871 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137711 129252
rect -71245 -58264 -70845 128496
rect -69921 128412 -69565 128896
rect -70761 128056 -69565 128412
rect 137355 128412 137711 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138551 128412
rect -70761 -57824 -70405 128056
rect 138195 -57824 138551 128056
rect -70761 -58180 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69921 -58664 -69565 -58180
rect 137355 -58180 138551 -57824
rect 137355 -58664 137711 -58180
rect 138635 -58264 139035 128496
rect -69921 -59020 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -69081 -59504 -68725 -59020
rect 136515 -59020 137711 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136871 -59020
rect 137795 -59104 138195 -58664
rect -69081 -59860 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68241 -60344 -67885 -59860
rect 135675 -59860 136871 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 136031 -59860
rect 136955 -59944 137355 -59504
rect -68241 -60700 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67401 -61184 -67045 -60700
rect 134835 -60700 136031 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135191 -60700
rect 136115 -60784 136515 -60344
rect -67401 -61540 135191 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia5 >>
rect -67485 131772 135275 131856
rect -67485 131016 -67401 131772
rect -68325 130932 -67401 131016
rect -68325 130176 -68241 130932
rect 135191 131016 135275 131772
rect 135191 130932 136115 131016
rect -69165 130092 -68241 130176
rect -69165 129336 -69081 130092
rect 136031 130176 136115 130932
rect 136031 130092 136955 130176
rect -70005 129252 -69081 129336
rect -70005 128496 -69921 129252
rect 136871 129336 136955 130092
rect 136871 129252 137795 129336
rect -70845 128412 -69921 128496
rect -70845 -58180 -70761 128412
rect 137711 128496 137795 129252
rect 137711 128412 138635 128496
rect -70845 -58264 -69921 -58180
rect -70005 -59020 -69921 -58264
rect 138551 -58180 138635 128412
rect 137711 -58264 138635 -58180
rect -70005 -59104 -69081 -59020
rect -69165 -59860 -69081 -59104
rect 137711 -59020 137795 -58264
rect 136871 -59104 137795 -59020
rect -69165 -59944 -68241 -59860
rect -68325 -60700 -68241 -59944
rect 136871 -59860 136955 -59104
rect 136031 -59944 136955 -59860
rect -68325 -60784 -67401 -60700
rect -67485 -61540 -67401 -60784
rect 136031 -60700 136115 -59944
rect 135191 -60784 136115 -60700
rect 135191 -61540 135275 -60784
rect -67485 -61624 135275 -61540
<< metal6 >>
rect -67885 131856 135675 132256
rect -67885 131416 -67485 131856
rect -68725 131016 -67485 131416
rect -67305 131416 135095 131676
rect -68725 130576 -68325 131016
rect -67305 130836 -67045 131416
rect -69565 130176 -68325 130576
rect -68145 130576 -67045 130836
rect 134835 130836 135095 131416
rect 135275 131416 135675 131856
rect 135275 131016 136515 131416
rect 134835 130576 135935 130836
rect -69565 129736 -69165 130176
rect -68145 129996 -67885 130576
rect -70405 129336 -69165 129736
rect -68985 129736 -67885 129996
rect 135675 129996 135935 130576
rect 136115 130576 136515 131016
rect 136115 130176 137355 130576
rect 135675 129736 136775 129996
rect -70405 128896 -70005 129336
rect -68985 129156 -68725 129736
rect -71245 128496 -70005 128896
rect -69825 128896 -68725 129156
rect 136515 129156 136775 129736
rect 136955 129736 137355 130176
rect 136955 129336 138195 129736
rect 136515 128896 137615 129156
rect -71245 -58264 -70845 128496
rect -69825 128316 -69565 128896
rect -70665 128056 -69565 128316
rect 137355 128316 137615 128896
rect 137795 128896 138195 129336
rect 137795 128496 139035 128896
rect 137355 128056 138455 128316
rect -70665 -57824 -70405 128056
rect 138195 -57824 138455 128056
rect -70665 -58084 -69565 -57824
rect -71245 -58664 -70005 -58264
rect -70405 -59104 -70005 -58664
rect -69825 -58664 -69565 -58084
rect 137355 -58084 138455 -57824
rect 137355 -58664 137615 -58084
rect 138635 -58264 139035 128496
rect -69825 -58924 -68725 -58664
rect -70405 -59504 -69165 -59104
rect -69565 -59944 -69165 -59504
rect -68985 -59504 -68725 -58924
rect 136515 -58924 137615 -58664
rect 137795 -58664 139035 -58264
rect 136515 -59504 136775 -58924
rect 137795 -59104 138195 -58664
rect -68985 -59764 -67885 -59504
rect -69565 -60344 -68325 -59944
rect -68725 -60784 -68325 -60344
rect -68145 -60344 -67885 -59764
rect 135675 -59764 136775 -59504
rect 136955 -59504 138195 -59104
rect 135675 -60344 135935 -59764
rect 136955 -59944 137355 -59504
rect -68145 -60604 -67045 -60344
rect -68725 -61184 -67485 -60784
rect -67885 -61624 -67485 -61184
rect -67305 -61184 -67045 -60604
rect 134835 -60604 135935 -60344
rect 136115 -60344 137355 -59944
rect 134835 -61184 135095 -60604
rect 136115 -60784 136515 -60344
rect -67305 -61444 135095 -61184
rect 135275 -61184 136515 -60784
rect 135275 -61624 135675 -61184
rect -67885 -62024 135675 -61624
<< sealvia6 >>
rect -67485 131676 135275 131856
rect -67485 131016 -67305 131676
rect -68325 130836 -67305 131016
rect -68325 130176 -68145 130836
rect 135095 131016 135275 131676
rect 135095 130836 136115 131016
rect -69165 129996 -68145 130176
rect -69165 129336 -68985 129996
rect 135935 130176 136115 130836
rect 135935 129996 136955 130176
rect -70005 129156 -68985 129336
rect -70005 128496 -69825 129156
rect 136775 129336 136955 129996
rect 136775 129156 137795 129336
rect -70845 128316 -69825 128496
rect -70845 -58084 -70665 128316
rect 137615 128496 137795 129156
rect 137615 128316 138635 128496
rect -70845 -58264 -69825 -58084
rect -70005 -58924 -69825 -58264
rect 138455 -58084 138635 128316
rect 137615 -58264 138635 -58084
rect -70005 -59104 -68985 -58924
rect -69165 -59764 -68985 -59104
rect 137615 -58924 137795 -58264
rect 136775 -59104 137795 -58924
rect -69165 -59944 -68145 -59764
rect -68325 -60604 -68145 -59944
rect 136775 -59764 136955 -59104
rect 135935 -59944 136955 -59764
rect -68325 -60784 -67305 -60604
rect -67485 -61444 -67305 -60784
rect 135935 -60604 136115 -59944
rect 135095 -60784 136115 -60604
rect 135095 -61444 135275 -60784
rect -67485 -61624 135275 -61444
<< metal7 >>
rect -67885 131416 135675 132256
rect -68725 130576 -67045 131416
rect 134835 130576 136515 131416
rect -69565 129736 -67885 130576
rect 135675 129736 137355 130576
rect -70405 128896 -68725 129736
rect 136515 128896 138195 129736
rect -71245 128056 -69565 128896
rect 137355 128056 139035 128896
rect -71245 -57824 -70405 128056
rect 138195 -57824 139035 128056
rect -71245 -58664 -69565 -57824
rect 137355 -58664 139035 -57824
rect -70405 -59504 -68725 -58664
rect 136515 -59504 138195 -58664
rect -69565 -60344 -67885 -59504
rect 135675 -60344 137355 -59504
rect -68725 -61184 -67045 -60344
rect 134835 -61184 136515 -60344
rect -67885 -62024 135675 -61184
<< seal >>
rect -69325 132856 137115 133696
rect -70165 132016 -68485 132856
rect -71005 131176 -69325 132016
rect 136275 132016 137955 132856
rect -71845 130336 -70165 131176
rect 137115 131176 138795 132016
rect -72685 129496 -71005 130336
rect 137955 130336 139635 131176
rect -72685 -59264 -71845 129496
rect 138795 129496 140475 130336
rect -72685 -60104 -71005 -59264
rect 139635 -59264 140475 129496
rect -71845 -60944 -70165 -60104
rect 138795 -60104 140475 -59264
rect -71005 -61784 -69325 -60944
rect 137955 -60944 139635 -60104
rect -70165 -62624 -68485 -61784
rect 137115 -61784 138795 -60944
rect 136275 -62624 137955 -61784
rect -69325 -63464 137115 -62624
<< end >>
