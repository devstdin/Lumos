magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 45 56 475 300
rect -26 -56 506 56
<< nmos >>
rect 139 120 165 274
rect 253 120 279 274
rect 355 120 381 274
<< pmos >>
rect 139 412 165 636
rect 253 412 279 636
rect 355 412 381 636
<< ndiff >>
rect 71 234 139 274
rect 71 202 85 234
rect 117 202 139 234
rect 71 166 139 202
rect 71 134 85 166
rect 117 134 139 166
rect 71 120 139 134
rect 165 234 253 274
rect 165 202 199 234
rect 231 202 253 234
rect 165 166 253 202
rect 165 134 199 166
rect 231 134 253 166
rect 165 120 253 134
rect 279 166 355 274
rect 279 134 301 166
rect 333 134 355 166
rect 279 120 355 134
rect 381 234 449 274
rect 381 202 403 234
rect 435 202 449 234
rect 381 166 449 202
rect 381 134 403 166
rect 435 134 449 166
rect 381 120 449 134
<< pdiff >>
rect 71 622 139 636
rect 71 590 85 622
rect 117 590 139 622
rect 71 554 139 590
rect 71 522 85 554
rect 117 522 139 554
rect 71 486 139 522
rect 71 454 85 486
rect 117 454 139 486
rect 71 412 139 454
rect 165 412 253 636
rect 279 412 355 636
rect 381 622 449 636
rect 381 590 403 622
rect 435 590 449 622
rect 381 554 449 590
rect 381 522 403 554
rect 435 522 449 554
rect 381 486 449 522
rect 381 454 403 486
rect 435 454 449 486
rect 381 412 449 454
<< ndiffc >>
rect 85 202 117 234
rect 85 134 117 166
rect 199 202 231 234
rect 199 134 231 166
rect 301 134 333 166
rect 403 202 435 234
rect 403 134 435 166
<< pdiffc >>
rect 85 590 117 622
rect 85 522 117 554
rect 85 454 117 486
rect 403 590 435 622
rect 403 522 435 554
rect 403 454 435 486
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 139 636 165 672
rect 253 636 279 672
rect 355 636 381 672
rect 139 370 165 412
rect 71 356 165 370
rect 71 324 85 356
rect 117 324 165 356
rect 71 310 165 324
rect 139 274 165 310
rect 253 370 279 412
rect 355 370 381 412
rect 253 356 313 370
rect 253 324 267 356
rect 299 324 313 356
rect 253 310 313 324
rect 355 356 415 370
rect 355 324 369 356
rect 401 324 415 356
rect 355 310 415 324
rect 253 274 279 310
rect 355 274 381 310
rect 139 60 165 120
rect 253 60 279 120
rect 355 60 381 120
<< polycont >>
rect 85 324 117 356
rect 267 324 299 356
rect 369 324 401 356
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 75 622 127 712
rect 75 590 85 622
rect 117 590 127 622
rect 75 554 127 590
rect 75 522 85 554
rect 117 522 127 554
rect 393 622 445 626
rect 393 590 403 622
rect 435 590 445 622
rect 393 554 445 590
rect 393 533 403 554
rect 75 486 127 522
rect 75 454 85 486
rect 117 454 127 486
rect 75 441 127 454
rect 189 522 403 533
rect 435 522 445 554
rect 189 486 445 522
rect 189 476 403 486
rect 68 356 124 370
rect 68 324 85 356
rect 117 324 124 356
rect 68 303 124 324
rect 189 244 224 476
rect 393 454 403 476
rect 435 454 445 486
rect 393 444 445 454
rect 260 356 316 370
rect 260 324 267 356
rect 299 324 316 356
rect 260 303 316 324
rect 356 356 412 370
rect 356 324 369 356
rect 401 324 412 356
rect 356 303 412 324
rect 75 234 127 244
rect 75 202 85 234
rect 117 202 127 234
rect 75 166 127 202
rect 75 134 85 166
rect 117 134 127 166
rect 75 44 127 134
rect 189 234 445 244
rect 189 202 199 234
rect 231 212 403 234
rect 231 202 241 212
rect 189 166 241 202
rect 393 202 403 212
rect 435 202 445 234
rect 189 134 199 166
rect 231 134 241 166
rect 189 124 241 134
rect 291 166 343 176
rect 291 134 301 166
rect 333 134 343 166
rect 291 44 343 134
rect 393 166 445 202
rect 393 134 403 166
rect 435 134 445 166
rect 393 124 445 134
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 68 303 124 370 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 192 476 445 533 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 260 303 316 370 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 356 303 412 370 0 FreeSans 400 0 0 0 C
port 5 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 149040
string GDS_FILE 6_final.gds
string GDS_START 144572
<< end >>
