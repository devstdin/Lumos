magic
tech ihp-sg13g2
timestamp 1748595295
<< error_p >>
rect -18 280 -13 285
rect 13 280 18 285
rect 160 280 165 285
rect 191 280 196 285
rect 338 280 343 285
rect 369 280 374 285
rect 516 280 521 285
rect 547 280 552 285
rect 694 280 699 285
rect 725 280 730 285
rect 872 280 877 285
rect 903 280 908 285
rect 1050 280 1055 285
rect 1081 280 1086 285
rect -23 275 23 280
rect 155 275 201 280
rect 333 275 379 280
rect 511 275 557 280
rect 689 275 735 280
rect 867 275 913 280
rect 1045 275 1091 280
rect -18 269 18 275
rect 160 269 196 275
rect 338 269 374 275
rect 516 269 552 275
rect 694 269 730 275
rect 872 269 908 275
rect 1050 269 1086 275
rect -23 264 23 269
rect 155 264 201 269
rect 333 264 379 269
rect 511 264 557 269
rect 689 264 735 269
rect 867 264 913 269
rect 1045 264 1091 269
rect -18 259 -13 264
rect 13 259 18 264
rect 160 259 165 264
rect 191 259 196 264
rect 338 259 343 264
rect 369 259 374 264
rect 516 259 521 264
rect 547 259 552 264
rect 694 259 699 264
rect 725 259 730 264
rect 872 259 877 264
rect 903 259 908 264
rect 1050 259 1055 264
rect 1081 259 1086 264
rect -52 243 -47 248
rect -41 243 -36 248
rect 36 243 41 248
rect 47 243 52 248
rect 126 243 131 248
rect 137 243 142 248
rect 214 243 219 248
rect 225 243 230 248
rect 304 243 309 248
rect 315 243 320 248
rect 392 243 397 248
rect 403 243 408 248
rect 482 243 487 248
rect 493 243 498 248
rect 570 243 575 248
rect 581 243 586 248
rect 660 243 665 248
rect 671 243 676 248
rect 748 243 753 248
rect 759 243 764 248
rect 838 243 843 248
rect 849 243 854 248
rect 926 243 931 248
rect 937 243 942 248
rect 1016 243 1021 248
rect 1027 243 1032 248
rect 1104 243 1109 248
rect 1115 243 1120 248
rect -57 238 -52 243
rect -36 238 -31 243
rect 31 238 36 243
rect 52 238 57 243
rect 121 238 126 243
rect 142 238 147 243
rect 209 238 214 243
rect 230 238 235 243
rect 299 238 304 243
rect 320 238 325 243
rect 387 238 392 243
rect 408 238 413 243
rect 477 238 482 243
rect 498 238 503 243
rect 565 238 570 243
rect 586 238 591 243
rect 655 238 660 243
rect 676 238 681 243
rect 743 238 748 243
rect 764 238 769 243
rect 833 238 838 243
rect 854 238 859 243
rect 921 238 926 243
rect 942 238 947 243
rect 1011 238 1016 243
rect 1032 238 1037 243
rect 1099 238 1104 243
rect 1120 238 1125 243
rect -57 -243 -52 -238
rect -36 -243 -31 -238
rect 31 -243 36 -238
rect 52 -243 57 -238
rect 121 -243 126 -238
rect 142 -243 147 -238
rect 209 -243 214 -238
rect 230 -243 235 -238
rect 299 -243 304 -238
rect 320 -243 325 -238
rect 387 -243 392 -238
rect 408 -243 413 -238
rect 477 -243 482 -238
rect 498 -243 503 -238
rect 565 -243 570 -238
rect 586 -243 591 -238
rect 655 -243 660 -238
rect 676 -243 681 -238
rect 743 -243 748 -238
rect 764 -243 769 -238
rect 833 -243 838 -238
rect 854 -243 859 -238
rect 921 -243 926 -238
rect 942 -243 947 -238
rect 1011 -243 1016 -238
rect 1032 -243 1037 -238
rect 1099 -243 1104 -238
rect 1120 -243 1125 -238
rect -52 -248 -47 -243
rect -41 -248 -36 -243
rect 36 -248 41 -243
rect 47 -248 52 -243
rect 126 -248 131 -243
rect 137 -248 142 -243
rect 214 -248 219 -243
rect 225 -248 230 -243
rect 304 -248 309 -243
rect 315 -248 320 -243
rect 392 -248 397 -243
rect 403 -248 408 -243
rect 482 -248 487 -243
rect 493 -248 498 -243
rect 570 -248 575 -243
rect 581 -248 586 -243
rect 660 -248 665 -243
rect 671 -248 676 -243
rect 748 -248 753 -243
rect 759 -248 764 -243
rect 838 -248 843 -243
rect 849 -248 854 -243
rect 926 -248 931 -243
rect 937 -248 942 -243
rect 1016 -248 1021 -243
rect 1027 -248 1032 -243
rect 1104 -248 1109 -243
rect 1115 -248 1120 -243
rect -18 -264 -13 -259
rect 13 -264 18 -259
rect 160 -264 165 -259
rect 191 -264 196 -259
rect 338 -264 343 -259
rect 369 -264 374 -259
rect 516 -264 521 -259
rect 547 -264 552 -259
rect 694 -264 699 -259
rect 725 -264 730 -259
rect 872 -264 877 -259
rect 903 -264 908 -259
rect 1050 -264 1055 -259
rect 1081 -264 1086 -259
rect -23 -269 23 -264
rect 155 -269 201 -264
rect 333 -269 379 -264
rect 511 -269 557 -264
rect 689 -269 735 -264
rect 867 -269 913 -264
rect 1045 -269 1091 -264
rect -18 -275 18 -269
rect 160 -275 196 -269
rect 338 -275 374 -269
rect 516 -275 552 -269
rect 694 -275 730 -269
rect 872 -275 908 -269
rect 1050 -275 1086 -269
rect -23 -280 23 -275
rect 155 -280 201 -275
rect 333 -280 379 -275
rect 511 -280 557 -275
rect 689 -280 735 -275
rect 867 -280 913 -275
rect 1045 -280 1091 -275
rect -18 -285 -13 -280
rect 13 -285 18 -280
rect 160 -285 165 -280
rect 191 -285 196 -280
rect 338 -285 343 -280
rect 369 -285 374 -280
rect 516 -285 521 -280
rect 547 -285 552 -280
rect 694 -285 699 -280
rect 725 -285 730 -280
rect 872 -285 877 -280
rect 903 -285 908 -280
rect 1050 -285 1055 -280
rect 1081 -285 1086 -280
<< nwell >>
rect -232 -412 1300 412
<< hvpmos >>
rect -25 -250 25 250
rect 153 -250 203 250
rect 331 -250 381 250
rect 509 -250 559 250
rect 687 -250 737 250
rect 865 -250 915 250
rect 1043 -250 1093 250
<< hvpdiff >>
rect -59 243 -25 250
rect -59 -243 -52 243
rect -36 -243 -25 243
rect -59 -250 -25 -243
rect 25 243 59 250
rect 25 -243 36 243
rect 52 -243 59 243
rect 25 -250 59 -243
rect 119 243 153 250
rect 119 -243 126 243
rect 142 -243 153 243
rect 119 -250 153 -243
rect 203 243 237 250
rect 203 -243 214 243
rect 230 -243 237 243
rect 203 -250 237 -243
rect 297 243 331 250
rect 297 -243 304 243
rect 320 -243 331 243
rect 297 -250 331 -243
rect 381 243 415 250
rect 381 -243 392 243
rect 408 -243 415 243
rect 381 -250 415 -243
rect 475 243 509 250
rect 475 -243 482 243
rect 498 -243 509 243
rect 475 -250 509 -243
rect 559 243 593 250
rect 559 -243 570 243
rect 586 -243 593 243
rect 559 -250 593 -243
rect 653 243 687 250
rect 653 -243 660 243
rect 676 -243 687 243
rect 653 -250 687 -243
rect 737 243 771 250
rect 737 -243 748 243
rect 764 -243 771 243
rect 737 -250 771 -243
rect 831 243 865 250
rect 831 -243 838 243
rect 854 -243 865 243
rect 831 -250 865 -243
rect 915 243 949 250
rect 915 -243 926 243
rect 942 -243 949 243
rect 915 -250 949 -243
rect 1009 243 1043 250
rect 1009 -243 1016 243
rect 1032 -243 1043 243
rect 1009 -250 1043 -243
rect 1093 243 1127 250
rect 1093 -243 1104 243
rect 1120 -243 1127 243
rect 1093 -250 1127 -243
<< hvpdiffc >>
rect -52 -243 -36 243
rect 36 -243 52 243
rect 126 -243 142 243
rect 214 -243 230 243
rect 304 -243 320 243
rect 392 -243 408 243
rect 482 -243 498 243
rect 570 -243 586 243
rect 660 -243 676 243
rect 748 -243 764 243
rect 838 -243 854 243
rect 926 -243 942 243
rect 1016 -243 1032 243
rect 1104 -243 1120 243
<< nsubdiff >>
rect -170 343 1238 350
rect -170 327 -133 343
rect 1201 327 1238 343
rect -170 320 1238 327
rect -170 313 -140 320
rect -170 -313 -163 313
rect -147 -313 -140 313
rect 1208 313 1238 320
rect -170 -320 -140 -313
rect 1208 -313 1215 313
rect 1231 -313 1238 313
rect 1208 -320 1238 -313
rect -170 -327 1238 -320
rect -170 -343 -133 -327
rect 1201 -343 1238 -327
rect -170 -350 1238 -343
<< nsubdiffcont >>
rect -133 327 1201 343
rect -163 -313 -147 313
rect 1215 -313 1231 313
rect -133 -343 1201 -327
<< poly >>
rect -25 280 25 287
rect -25 264 -18 280
rect 18 264 25 280
rect -25 250 25 264
rect 153 280 203 287
rect 153 264 160 280
rect 196 264 203 280
rect 153 250 203 264
rect 331 280 381 287
rect 331 264 338 280
rect 374 264 381 280
rect 331 250 381 264
rect 509 280 559 287
rect 509 264 516 280
rect 552 264 559 280
rect 509 250 559 264
rect 687 280 737 287
rect 687 264 694 280
rect 730 264 737 280
rect 687 250 737 264
rect 865 280 915 287
rect 865 264 872 280
rect 908 264 915 280
rect 865 250 915 264
rect 1043 280 1093 287
rect 1043 264 1050 280
rect 1086 264 1093 280
rect 1043 250 1093 264
rect -25 -264 25 -250
rect -25 -280 -18 -264
rect 18 -280 25 -264
rect -25 -287 25 -280
rect 153 -264 203 -250
rect 153 -280 160 -264
rect 196 -280 203 -264
rect 153 -287 203 -280
rect 331 -264 381 -250
rect 331 -280 338 -264
rect 374 -280 381 -264
rect 331 -287 381 -280
rect 509 -264 559 -250
rect 509 -280 516 -264
rect 552 -280 559 -264
rect 509 -287 559 -280
rect 687 -264 737 -250
rect 687 -280 694 -264
rect 730 -280 737 -264
rect 687 -287 737 -280
rect 865 -264 915 -250
rect 865 -280 872 -264
rect 908 -280 915 -264
rect 865 -287 915 -280
rect 1043 -264 1093 -250
rect 1043 -280 1050 -264
rect 1086 -280 1093 -264
rect 1043 -287 1093 -280
<< polycont >>
rect -18 264 18 280
rect 160 264 196 280
rect 338 264 374 280
rect 516 264 552 280
rect 694 264 730 280
rect 872 264 908 280
rect 1050 264 1086 280
rect -18 -280 18 -264
rect 160 -280 196 -264
rect 338 -280 374 -264
rect 516 -280 552 -264
rect 694 -280 730 -264
rect 872 -280 908 -264
rect 1050 -280 1086 -264
<< metal1 >>
rect -168 343 1236 348
rect -168 327 -133 343
rect 1201 327 1236 343
rect -168 322 1236 327
rect -168 313 -142 322
rect -168 -313 -163 313
rect -147 -313 -142 313
rect 1210 313 1236 322
rect -168 -322 -142 -313
rect 1210 -313 1215 313
rect 1231 -313 1236 313
rect 1210 -322 1236 -313
rect -168 -327 1236 -322
rect -168 -343 -133 -327
rect 1201 -343 1236 -327
rect -168 -348 1236 -343
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 5 l 0.5 nf 1 nx 7 dx 0.6 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 1
<< end >>
