magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< nwell >>
rect 8084 51 8269 648
rect 0 -101 8269 51
rect 8084 -697 8269 -101
rect 8265 -4031 9253 -3934
<< metal1 >>
rect -1927 -859 -1022 801
rect -260 481 9253 801
rect -260 -569 180 481
rect 350 128 392 481
rect 428 342 560 394
rect 458 106 530 342
rect 428 54 560 106
rect 596 54 638 320
rect 688 128 730 481
rect 766 342 898 394
rect 796 106 868 342
rect 766 54 898 106
rect 934 54 976 320
rect 1026 128 1068 481
rect 1104 342 1236 394
rect 1134 106 1206 342
rect 1104 54 1236 106
rect 1272 54 1314 320
rect 1364 128 1406 481
rect 1442 342 1574 394
rect 1472 106 1544 342
rect 1442 54 1574 106
rect 1610 54 1652 320
rect 1702 128 1744 481
rect 1780 342 1912 394
rect 1810 106 1882 342
rect 1780 54 1912 106
rect 1948 54 1990 320
rect 2040 128 2082 481
rect 2118 342 2250 394
rect 2148 106 2220 342
rect 2118 54 2250 106
rect 2286 54 2328 320
rect 2378 128 2420 481
rect 2456 342 2588 394
rect 2486 106 2558 342
rect 2456 54 2588 106
rect 2624 54 2666 320
rect 2716 128 2758 481
rect 2794 342 2926 394
rect 2824 106 2896 342
rect 2794 54 2926 106
rect 2962 54 3004 320
rect 3054 128 3096 481
rect 3132 342 3264 394
rect 3162 106 3234 342
rect 3132 54 3264 106
rect 3300 54 3342 320
rect 3392 128 3434 481
rect 3470 342 3602 394
rect 3500 106 3572 342
rect 3470 54 3602 106
rect 3638 54 3680 320
rect 3730 128 3772 481
rect 3808 342 3940 394
rect 3838 106 3910 342
rect 3808 54 3940 106
rect 350 -15 3940 54
rect 350 -369 392 -15
rect 428 -113 2926 -64
rect 428 -155 560 -113
rect 2794 -155 2926 -113
rect 458 -391 530 -155
rect 596 -187 701 -177
rect 596 -391 648 -187
rect 428 -433 648 -391
rect 691 -433 701 -187
rect 2646 -187 2758 -177
rect 2646 -359 2656 -187
rect 2702 -359 2758 -187
rect 2646 -369 2758 -359
rect 2824 -391 2896 -155
rect 3976 -171 4018 320
rect 4068 128 4110 476
rect 4146 342 4278 394
rect 4176 106 4248 342
rect 4146 54 4278 106
rect 4314 54 4356 320
rect 4406 128 4448 476
rect 4484 342 4616 394
rect 4514 106 4586 342
rect 4484 54 4616 106
rect 4652 54 4694 320
rect 4744 128 4786 476
rect 4822 342 4954 394
rect 4852 106 4924 342
rect 4822 54 4954 106
rect 4990 54 5032 320
rect 5082 128 5124 476
rect 5160 342 5292 394
rect 5190 106 5262 342
rect 5160 54 5292 106
rect 5328 54 5370 320
rect 5420 128 5462 476
rect 5498 342 5630 394
rect 5528 106 5600 342
rect 5498 54 5630 106
rect 5666 54 5708 320
rect 5758 128 5800 476
rect 5836 342 5968 394
rect 5866 106 5938 342
rect 5836 54 5968 106
rect 6004 54 6046 320
rect 6096 128 6138 476
rect 6174 342 6306 394
rect 6204 106 6276 342
rect 6174 54 6306 106
rect 6342 54 6384 320
rect 6434 128 6476 476
rect 6512 342 6644 394
rect 6542 106 6614 342
rect 6512 54 6644 106
rect 6680 54 6722 320
rect 6772 128 6814 476
rect 6850 342 6982 394
rect 6880 106 6952 342
rect 6850 54 6982 106
rect 7018 54 7060 320
rect 7110 128 7152 476
rect 7188 342 7320 394
rect 7218 106 7290 342
rect 7188 54 7320 106
rect 7356 54 7398 320
rect 7448 128 7490 476
rect 7526 342 7658 394
rect 7556 106 7628 342
rect 7526 54 7658 106
rect 2962 -240 4018 -171
rect 4068 -15 7658 54
rect 4068 -171 4110 -15
rect 5160 -113 7658 -63
rect 5160 -155 5292 -113
rect 7526 -155 7658 -113
rect 4068 -240 5124 -171
rect 2962 -369 3004 -240
rect 5082 -369 5124 -240
rect 5190 -391 5262 -155
rect 5328 -187 5433 -177
rect 5328 -391 5380 -187
rect 428 -443 701 -433
rect 2794 -443 2926 -391
rect 5160 -433 5380 -391
rect 5423 -433 5433 -187
rect 7378 -187 7490 -177
rect 7378 -359 7388 -187
rect 7434 -359 7490 -187
rect 7378 -369 7490 -359
rect 7556 -391 7628 -155
rect 7694 -369 7736 320
rect 5160 -443 5433 -433
rect 7526 -443 7658 -391
rect 7912 -568 8445 481
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect 242 -869 3940 -859
rect 242 -937 252 -869
rect 301 -902 3940 -869
rect 301 -937 311 -902
rect 242 -947 311 -937
rect 428 -944 560 -902
rect -1927 -1310 -1022 -1228
rect 350 -1310 392 -966
rect 458 -1180 530 -944
rect 596 -1158 638 -902
rect 766 -944 898 -902
rect 428 -1232 560 -1180
rect 688 -1310 730 -966
rect 796 -1180 868 -944
rect 934 -1158 976 -902
rect 1104 -944 1236 -902
rect 766 -1232 898 -1180
rect 1026 -1310 1068 -966
rect 1134 -1180 1206 -944
rect 1272 -1158 1314 -902
rect 1442 -944 1574 -902
rect 1104 -1232 1236 -1180
rect 1364 -1310 1406 -966
rect 1472 -1180 1544 -944
rect 1610 -1158 1652 -902
rect 1780 -944 1912 -902
rect 1442 -1232 1574 -1180
rect 1702 -1310 1744 -966
rect 1810 -1180 1882 -944
rect 1948 -1158 1990 -902
rect 2118 -944 2250 -902
rect 1780 -1232 1912 -1180
rect 2040 -1310 2082 -966
rect 2148 -1180 2220 -944
rect 2286 -1158 2328 -902
rect 2456 -944 2588 -902
rect 2118 -1232 2250 -1180
rect 2378 -1310 2420 -966
rect 2486 -1180 2558 -944
rect 2624 -1158 2666 -902
rect 2794 -944 2926 -902
rect 2456 -1232 2588 -1180
rect 2716 -1310 2758 -966
rect 2824 -1180 2896 -944
rect 2962 -1158 3004 -902
rect 3132 -944 3264 -902
rect 2794 -1232 2926 -1180
rect 3054 -1310 3096 -966
rect 3162 -1180 3234 -944
rect 3300 -1158 3342 -902
rect 3470 -944 3602 -902
rect 3132 -1232 3264 -1180
rect 3392 -1310 3434 -966
rect 3500 -1180 3572 -944
rect 3638 -1158 3680 -902
rect 3808 -944 3940 -902
rect 4146 -902 7658 -859
rect 4146 -944 4278 -902
rect 3470 -1232 3602 -1180
rect 3730 -1310 3772 -966
rect 3838 -1180 3910 -944
rect 3976 -1003 4022 -966
rect 3954 -1013 4022 -1003
rect 3954 -1111 3964 -1013
rect 4012 -1111 4022 -1013
rect 3954 -1121 4022 -1111
rect 3976 -1158 4022 -1121
rect 3808 -1232 3940 -1180
rect 4068 -1310 4110 -966
rect 4176 -1180 4248 -944
rect 4314 -1003 4360 -902
rect 4484 -944 4616 -902
rect 4292 -1013 4360 -1003
rect 4292 -1111 4302 -1013
rect 4350 -1111 4360 -1013
rect 4292 -1121 4360 -1111
rect 4314 -1158 4360 -1121
rect 4146 -1232 4278 -1180
rect 4406 -1310 4448 -966
rect 4514 -1180 4586 -944
rect 4652 -1158 4694 -902
rect 4822 -944 4954 -902
rect 4484 -1232 4616 -1180
rect 4744 -1310 4786 -966
rect 4852 -1180 4924 -944
rect 4990 -1158 5032 -902
rect 5160 -944 5292 -902
rect 4822 -1232 4954 -1180
rect 5082 -1310 5124 -966
rect 5190 -1180 5262 -944
rect 5328 -1158 5370 -902
rect 5498 -944 5630 -902
rect 5160 -1232 5292 -1180
rect 5420 -1310 5462 -966
rect 5528 -1180 5600 -944
rect 5666 -1158 5708 -902
rect 5836 -944 5968 -902
rect 5498 -1232 5630 -1180
rect 5758 -1310 5800 -966
rect 5866 -1180 5938 -944
rect 6004 -1158 6046 -902
rect 6174 -944 6306 -902
rect 5836 -1232 5968 -1180
rect 6096 -1310 6138 -966
rect 6204 -1180 6276 -944
rect 6342 -1158 6384 -902
rect 6512 -944 6644 -902
rect 6174 -1232 6306 -1180
rect 6434 -1310 6476 -966
rect 6542 -1180 6614 -944
rect 6680 -1158 6722 -902
rect 6850 -944 6982 -902
rect 6512 -1232 6644 -1180
rect 6772 -1310 6814 -966
rect 6880 -1180 6952 -944
rect 7018 -1158 7060 -902
rect 7188 -944 7320 -902
rect 6850 -1232 6982 -1180
rect 7110 -1310 7152 -966
rect 7218 -1180 7290 -944
rect 7356 -1158 7398 -902
rect 7526 -944 7658 -902
rect 7188 -1232 7320 -1180
rect 7448 -1310 7490 -966
rect 7556 -1180 7628 -944
rect 7694 -972 7786 -962
rect 7694 -1152 7704 -972
rect 7776 -1152 7786 -972
rect 7694 -1162 7786 -1152
rect 7526 -1232 7658 -1180
rect -1927 -1654 8169 -1310
rect 7825 -4821 8169 -1654
rect 8286 -4349 8445 -568
rect 8565 320 8611 480
rect 8693 342 8825 394
rect 8565 -1672 8657 320
rect 8719 -1694 8799 342
rect 8693 -1736 8825 -1694
rect 8527 -1746 8825 -1736
rect 8527 -1790 8537 -1746
rect 8615 -1790 8825 -1746
rect 8527 -1800 8825 -1790
rect 8693 -1842 8825 -1800
rect 8565 -3856 8657 -1864
rect 8565 -4003 8625 -3856
rect 8719 -3878 8799 -1842
rect 8861 -3856 8953 320
rect 8693 -3930 8825 -3878
rect 8565 -4045 8825 -4003
rect 8693 -4087 8825 -4045
rect 8519 -4115 8657 -4105
rect 8519 -4195 8529 -4115
rect 8601 -4195 8657 -4115
rect 8519 -4205 8657 -4195
rect 8719 -4223 8799 -4087
rect 8907 -4105 8953 -3856
rect 8861 -4205 8953 -4105
rect 8693 -4233 8825 -4223
rect 8693 -4303 8703 -4233
rect 8815 -4303 8825 -4233
rect 8693 -4313 8825 -4303
rect 9078 -4349 9253 481
rect 8286 -4359 9253 -4349
rect 8286 -4444 8574 -4359
rect 8661 -4444 9253 -4359
rect 8286 -4454 9253 -4444
rect 7825 -4831 9253 -4821
rect 7825 -4916 8422 -4831
rect 8509 -4916 9253 -4831
rect 7825 -4926 9253 -4916
rect 7825 -5124 8442 -4926
rect 8692 -4972 8824 -4962
rect 8692 -5042 8702 -4972
rect 8814 -5042 8824 -4972
rect 8692 -5052 8824 -5042
rect 8286 -9742 8442 -5124
rect 8518 -5080 8656 -5070
rect 8518 -5160 8528 -5080
rect 8600 -5160 8656 -5080
rect 8518 -5170 8656 -5160
rect 8718 -5188 8798 -5052
rect 8860 -5170 8952 -5070
rect 8692 -5230 8824 -5188
rect 8564 -5272 8824 -5230
rect 8564 -5416 8624 -5272
rect 8692 -5394 8824 -5342
rect 8564 -7408 8656 -5416
rect 8718 -7430 8798 -5394
rect 8906 -5416 8952 -5170
rect 8692 -7472 8824 -7430
rect 8526 -7482 8824 -7472
rect 8526 -7526 8536 -7482
rect 8614 -7526 8824 -7482
rect 8526 -7536 8824 -7526
rect 8692 -7578 8824 -7536
rect 8564 -9592 8656 -7600
rect 8564 -9742 8610 -9592
rect 8718 -9614 8798 -7578
rect 8860 -9592 8952 -5416
rect 8692 -9666 8824 -9614
rect 9072 -9742 9253 -4926
rect 8286 -9940 9253 -9742
<< via1 >>
rect 648 -433 691 -187
rect 2656 -359 2702 -187
rect 5380 -433 5423 -187
rect 7388 -359 7434 -187
rect -1845 -1228 -1104 -859
rect 252 -937 301 -869
rect 3964 -1111 4012 -1013
rect 4302 -1111 4350 -1013
rect 7704 -1152 7776 -972
rect 8537 -1790 8615 -1746
rect 8529 -4195 8601 -4115
rect 8703 -4303 8815 -4233
rect 8574 -4444 8661 -4359
rect 8422 -4916 8509 -4831
rect 8702 -5042 8814 -4972
rect 8528 -5160 8600 -5080
rect 8536 -7526 8614 -7482
<< metal2 >>
rect -1927 -859 -1022 -777
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect -734 -859 -541 801
rect 638 -187 701 -177
rect 638 -433 648 -187
rect 691 -433 701 -187
rect 638 -622 701 -433
rect 2646 -187 2712 -177
rect 2646 -359 2656 -187
rect 2702 -359 2712 -187
rect 2646 -481 2712 -359
rect 5370 -187 5433 -177
rect 5370 -433 5380 -187
rect 5423 -433 5433 -187
rect 2646 -547 4360 -481
rect 638 -685 4022 -622
rect -734 -869 311 -859
rect -734 -937 252 -869
rect 301 -937 311 -869
rect -734 -1052 311 -937
rect 3976 -1003 4022 -685
rect 4314 -1003 4360 -547
rect 5370 -622 5433 -433
rect 7378 -187 7444 -177
rect 7378 -359 7388 -187
rect 7434 -359 7444 -187
rect 7378 -481 7444 -359
rect 7378 -547 8001 -481
rect 5370 -685 7786 -622
rect 7740 -962 7786 -685
rect 3954 -1013 4022 -1003
rect 3954 -1111 3964 -1013
rect 4012 -1111 4022 -1013
rect 3954 -1121 4022 -1111
rect 4292 -1013 4360 -1003
rect 4292 -1111 4302 -1013
rect 4350 -1111 4360 -1013
rect 4292 -1121 4360 -1111
rect 7694 -972 7786 -962
rect 7694 -1152 7704 -972
rect 7776 -1152 7786 -972
rect 7694 -1162 7786 -1152
rect -1927 -1310 -1022 -1228
rect 7871 -1736 8001 -547
rect 7871 -1746 8625 -1736
rect 7871 -1790 8537 -1746
rect 8615 -1790 8625 -1746
rect 7871 -1800 8625 -1790
rect 8121 -5937 8265 -1800
rect 8473 -4115 8611 -4105
rect 8473 -4195 8529 -4115
rect 8601 -4195 8611 -4115
rect 8473 -4205 8611 -4195
rect 8473 -4821 8519 -4205
rect 8693 -4233 8825 -4223
rect 8693 -4303 8703 -4233
rect 8815 -4303 8825 -4233
rect 8693 -4313 8825 -4303
rect 8412 -4831 8519 -4821
rect 8412 -4916 8422 -4831
rect 8509 -4916 8519 -4831
rect 8412 -4926 8519 -4916
rect 8564 -4359 8671 -4349
rect 8564 -4444 8574 -4359
rect 8661 -4444 8671 -4359
rect 8564 -4454 8671 -4444
rect 8564 -5070 8610 -4454
rect 8718 -4532 8799 -4313
rect 8718 -4752 9253 -4532
rect 8718 -4962 8799 -4752
rect 8692 -4972 8824 -4962
rect 8692 -5042 8702 -4972
rect 8814 -5042 8824 -4972
rect 8692 -5052 8824 -5042
rect 8518 -5080 8610 -5070
rect 8518 -5160 8528 -5080
rect 8600 -5160 8610 -5080
rect 8518 -5170 8610 -5160
rect 8121 -7526 8131 -5937
rect 8255 -7472 8265 -5937
rect 8255 -7482 8624 -7472
rect 8255 -7526 8536 -7482
rect 8614 -7526 8624 -7482
rect 8121 -7536 8624 -7526
<< via2 >>
rect -1845 -1228 -1104 -859
rect 8131 -7526 8255 -5937
<< metal3 >>
rect -1927 -859 -1022 -777
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect -1927 -1310 -1022 -1228
rect 7599 -5937 8265 -5927
rect 7599 -5947 8131 -5937
rect 7599 -7516 7619 -5947
rect 7599 -7526 8131 -7516
rect 8255 -7526 8265 -5937
rect 7599 -7536 8265 -7526
<< via3 >>
rect -1845 -1228 -1104 -859
rect 7619 -7516 8131 -5947
rect 8131 -7516 8245 -5947
<< metal4 >>
rect -1927 -859 -1022 -777
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect -1927 -1310 -1022 -1228
rect -9582 -3087 -5342 -1487
rect -5142 -3087 -902 -1487
rect -702 -3087 3538 -1487
rect 3738 -3087 7978 -1487
rect -9582 -4127 7978 -3087
rect -9582 -5727 -5342 -4127
rect -5142 -5727 -902 -4127
rect -702 -5727 3538 -4127
rect 3738 -5727 7978 -4127
rect -7982 -5927 -6942 -5727
rect 5338 -5927 6378 -5727
rect -9582 -7527 -5342 -5927
rect -5142 -7527 -902 -5927
rect -702 -7527 3538 -5927
rect 3738 -5947 8265 -5927
rect 3738 -7516 7619 -5947
rect 8245 -7516 8265 -5947
rect 3738 -7527 8265 -7516
rect -9582 -7536 8265 -7527
rect -9582 -8567 7978 -7536
rect -9582 -10167 -5342 -8567
rect -5142 -10167 -902 -8567
rect -702 -10167 3538 -8567
rect 3738 -10167 7978 -8567
<< via4 >>
rect -1845 -1228 -1104 -859
<< metal5 >>
rect -1927 -859 -1022 -777
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect -1927 -1310 -1022 -1228
<< via5 >>
rect -1845 -1228 -1104 -859
<< metal6 >>
rect -1927 -859 -1022 -777
rect -1927 -1228 -1845 -859
rect -1104 -1228 -1022 -859
rect -1927 -1607 -1022 -1228
rect -9462 -3087 -5462 -1607
rect -5022 -3087 -1022 -1607
rect -582 -3087 3418 -1607
rect 3858 -3087 7858 -1607
rect -9462 -4127 7858 -3087
rect -9462 -5607 -5462 -4127
rect -5022 -5607 -1022 -4127
rect -582 -5607 3418 -4127
rect 3858 -5607 7858 -4127
rect -7982 -6047 -6942 -5607
rect 5338 -6047 6378 -5607
rect -9462 -7527 -5462 -6047
rect -5022 -7527 -1022 -6047
rect -582 -7527 3418 -6047
rect 3858 -7527 7858 -6047
rect -9462 -8567 7858 -7527
rect -9462 -10047 -5462 -8567
rect -5022 -10047 -1022 -8567
rect -582 -10047 3418 -8567
rect 3858 -10047 7858 -8567
use cmim_XD4LYE  cmim_XD4LYE_0
timestamp 1757240632
transform 0 1 -7462 -1 0 -3607
box -2120 -2120 6560 15440
use hvnmos_4SCLER  hvnmos_4SCLER_0
timestamp 1757240632
transform 1 0 8758 0 1 -5120
box -370 -124 370 250
use hvnmos_NH3G3K  hvnmos_NH3G3K_0
timestamp 1757240632
transform 1 0 8758 0 1 -8596
box -370 -1200 370 3258
use hvnmos_WF38FF  hvnmos_WF38FF_0
timestamp 1757240632
transform 1 0 494 0 1 -1062
box -370 -300 7468 300
use hvpmos_7J3G3K  hvpmos_7J3G3K_0
timestamp 1757240632
transform 1 0 8759 0 1 -2860
box -494 -1124 494 3508
use hvpmos_MRCLER  hvpmos_MRCLER_0
timestamp 1757240632
transform 1 0 8759 0 1 -4155
box -494 -374 494 174
use hvpmos_UG3GPR  hvpmos_UG3GPR_0
timestamp 1757240632
transform 1 0 494 0 1 -273
box -494 -424 7592 224
use hvpmos_XF38FF  hvpmos_XF38FF_0
timestamp 1757240632
transform 1 0 494 0 1 224
box -494 -224 7592 424
<< labels >>
flabel metal1 -260 568 253 801 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal1 -1927 568 -1022 801 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal2 -734 568 -541 801 0 FreeSans 800 0 0 0 IBIAS
port 2 nsew
flabel metal2 8799 -4752 9253 -4532 0 FreeSans 800 0 0 0 RESET
port 3 nsew
<< end >>
