magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 1200 834
<< pwell >>
rect 19 56 1152 314
rect -26 -56 1178 56
<< nmos >>
rect 114 140 140 288
rect 216 140 242 288
rect 420 140 446 288
rect 522 140 548 288
rect 624 140 650 288
rect 726 140 752 288
rect 930 140 956 288
rect 1032 140 1058 288
<< pmos >>
rect 114 412 140 636
rect 216 412 242 636
rect 420 412 446 636
rect 522 412 548 636
rect 624 412 650 636
rect 726 412 752 636
rect 930 412 956 636
rect 1032 412 1058 636
<< ndiff >>
rect 45 254 114 288
rect 45 222 60 254
rect 92 222 114 254
rect 45 186 114 222
rect 45 154 60 186
rect 92 154 114 186
rect 45 140 114 154
rect 140 254 216 288
rect 140 222 162 254
rect 194 222 216 254
rect 140 186 216 222
rect 140 154 162 186
rect 194 154 216 186
rect 140 140 216 154
rect 242 186 420 288
rect 242 154 264 186
rect 296 154 366 186
rect 398 154 420 186
rect 242 140 420 154
rect 446 254 522 288
rect 446 222 468 254
rect 500 222 522 254
rect 446 186 522 222
rect 446 154 468 186
rect 500 154 522 186
rect 446 140 522 154
rect 548 186 624 288
rect 548 154 570 186
rect 602 154 624 186
rect 548 140 624 154
rect 650 254 726 288
rect 650 222 672 254
rect 704 222 726 254
rect 650 186 726 222
rect 650 154 672 186
rect 704 154 726 186
rect 650 140 726 154
rect 752 186 930 288
rect 752 154 774 186
rect 806 154 876 186
rect 908 154 930 186
rect 752 140 930 154
rect 956 254 1032 288
rect 956 222 978 254
rect 1010 222 1032 254
rect 956 186 1032 222
rect 956 154 978 186
rect 1010 154 1032 186
rect 956 140 1032 154
rect 1058 254 1126 288
rect 1058 222 1080 254
rect 1112 222 1126 254
rect 1058 186 1126 222
rect 1058 154 1080 186
rect 1112 154 1126 186
rect 1058 140 1126 154
<< pdiff >>
rect 45 622 114 636
rect 45 590 60 622
rect 92 590 114 622
rect 45 554 114 590
rect 45 522 60 554
rect 92 522 114 554
rect 45 486 114 522
rect 45 454 60 486
rect 92 454 114 486
rect 45 412 114 454
rect 140 622 216 636
rect 140 590 162 622
rect 194 590 216 622
rect 140 554 216 590
rect 140 522 162 554
rect 194 522 216 554
rect 140 486 216 522
rect 140 454 162 486
rect 194 454 216 486
rect 140 412 216 454
rect 242 622 310 636
rect 242 590 264 622
rect 296 590 310 622
rect 242 554 310 590
rect 242 522 264 554
rect 296 522 310 554
rect 242 412 310 522
rect 352 622 420 636
rect 352 590 366 622
rect 398 590 420 622
rect 352 554 420 590
rect 352 522 366 554
rect 398 522 420 554
rect 352 412 420 522
rect 446 554 522 636
rect 446 522 468 554
rect 500 522 522 554
rect 446 486 522 522
rect 446 454 468 486
rect 500 454 522 486
rect 446 412 522 454
rect 548 622 624 636
rect 548 590 570 622
rect 602 590 624 622
rect 548 554 624 590
rect 548 522 570 554
rect 602 522 624 554
rect 548 486 624 522
rect 548 454 570 486
rect 602 454 624 486
rect 548 412 624 454
rect 650 554 726 636
rect 650 522 672 554
rect 704 522 726 554
rect 650 486 726 522
rect 650 454 672 486
rect 704 454 726 486
rect 650 412 726 454
rect 752 622 820 636
rect 752 590 774 622
rect 806 590 820 622
rect 752 554 820 590
rect 752 522 774 554
rect 806 522 820 554
rect 752 412 820 522
rect 862 622 930 636
rect 862 590 876 622
rect 908 590 930 622
rect 862 554 930 590
rect 862 522 876 554
rect 908 522 930 554
rect 862 486 930 522
rect 862 454 876 486
rect 908 454 930 486
rect 862 412 930 454
rect 956 554 1032 636
rect 956 522 978 554
rect 1010 522 1032 554
rect 956 486 1032 522
rect 956 454 978 486
rect 1010 454 1032 486
rect 956 412 1032 454
rect 1058 622 1126 636
rect 1058 590 1080 622
rect 1112 590 1126 622
rect 1058 554 1126 590
rect 1058 522 1080 554
rect 1112 522 1126 554
rect 1058 486 1126 522
rect 1058 454 1080 486
rect 1112 454 1126 486
rect 1058 412 1126 454
<< ndiffc >>
rect 60 222 92 254
rect 60 154 92 186
rect 162 222 194 254
rect 162 154 194 186
rect 264 154 296 186
rect 366 154 398 186
rect 468 222 500 254
rect 468 154 500 186
rect 570 154 602 186
rect 672 222 704 254
rect 672 154 704 186
rect 774 154 806 186
rect 876 154 908 186
rect 978 222 1010 254
rect 978 154 1010 186
rect 1080 222 1112 254
rect 1080 154 1112 186
<< pdiffc >>
rect 60 590 92 622
rect 60 522 92 554
rect 60 454 92 486
rect 162 590 194 622
rect 162 522 194 554
rect 162 454 194 486
rect 264 590 296 622
rect 264 522 296 554
rect 366 590 398 622
rect 366 522 398 554
rect 468 522 500 554
rect 468 454 500 486
rect 570 590 602 622
rect 570 522 602 554
rect 570 454 602 486
rect 672 522 704 554
rect 672 454 704 486
rect 774 590 806 622
rect 774 522 806 554
rect 876 590 908 622
rect 876 522 908 554
rect 876 454 908 486
rect 978 522 1010 554
rect 978 454 1010 486
rect 1080 590 1112 622
rect 1080 522 1112 554
rect 1080 454 1112 486
<< psubdiff >>
rect 0 16 1152 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1152 16
rect 0 -30 1152 -16
<< nsubdiff >>
rect 0 772 1152 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1152 772
rect 0 726 1152 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
<< poly >>
rect 114 636 140 672
rect 216 636 242 672
rect 420 636 446 672
rect 522 636 548 672
rect 624 636 650 672
rect 726 636 752 672
rect 930 636 956 672
rect 1032 636 1058 672
rect 114 380 140 412
rect 216 380 242 412
rect 114 366 242 380
rect 114 334 128 366
rect 160 334 196 366
rect 228 334 242 366
rect 114 320 242 334
rect 114 288 140 320
rect 216 288 242 320
rect 420 380 446 412
rect 522 380 548 412
rect 420 366 548 380
rect 420 334 434 366
rect 466 334 502 366
rect 534 334 548 366
rect 420 320 548 334
rect 420 288 446 320
rect 522 288 548 320
rect 624 380 650 412
rect 726 380 752 412
rect 930 380 956 412
rect 1032 380 1058 412
rect 624 366 752 380
rect 624 334 638 366
rect 670 334 706 366
rect 738 334 752 366
rect 624 320 752 334
rect 872 366 1058 380
rect 872 334 886 366
rect 918 334 1058 366
rect 872 320 1058 334
rect 624 288 650 320
rect 726 288 752 320
rect 930 288 956 320
rect 1032 288 1058 320
rect 114 104 140 140
rect 216 104 242 140
rect 420 104 446 140
rect 522 104 548 140
rect 624 104 650 140
rect 726 104 752 140
rect 930 104 956 140
rect 1032 104 1058 140
<< polycont >>
rect 128 334 160 366
rect 196 334 228 366
rect 434 334 466 366
rect 502 334 534 366
rect 638 334 670 366
rect 706 334 738 366
rect 886 334 918 366
<< metal1 >>
rect 0 772 1152 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1152 772
rect 0 712 1152 740
rect 50 622 102 712
rect 50 590 60 622
rect 92 590 102 622
rect 50 554 102 590
rect 50 522 60 554
rect 92 522 102 554
rect 50 486 102 522
rect 50 454 60 486
rect 92 454 102 486
rect 50 444 102 454
rect 152 622 204 632
rect 152 590 162 622
rect 194 590 204 622
rect 152 554 204 590
rect 152 522 162 554
rect 194 522 204 554
rect 152 486 204 522
rect 254 622 306 712
rect 254 590 264 622
rect 296 590 306 622
rect 254 554 306 590
rect 254 522 264 554
rect 296 522 306 554
rect 254 512 306 522
rect 356 622 816 636
rect 356 590 366 622
rect 398 600 570 622
rect 398 590 408 600
rect 356 554 408 590
rect 560 590 570 600
rect 602 600 774 622
rect 602 590 612 600
rect 356 522 366 554
rect 398 522 408 554
rect 356 512 408 522
rect 458 554 510 564
rect 458 522 468 554
rect 500 522 510 554
rect 152 454 162 486
rect 194 476 204 486
rect 458 486 510 522
rect 458 476 468 486
rect 194 454 468 476
rect 500 454 510 486
rect 152 436 510 454
rect 560 554 612 590
rect 764 590 774 600
rect 806 590 816 622
rect 560 522 570 554
rect 602 522 612 554
rect 560 486 612 522
rect 560 454 570 486
rect 602 454 612 486
rect 560 444 612 454
rect 662 554 714 564
rect 662 522 672 554
rect 704 522 714 554
rect 662 486 714 522
rect 764 554 816 590
rect 764 522 774 554
rect 806 522 816 554
rect 764 512 816 522
rect 866 622 1122 632
rect 866 590 876 622
rect 908 600 1080 622
rect 908 590 918 600
rect 866 554 918 590
rect 1070 590 1080 600
rect 1112 590 1122 622
rect 866 522 876 554
rect 908 522 918 554
rect 662 454 672 486
rect 704 476 714 486
rect 866 486 918 522
rect 866 476 876 486
rect 704 454 876 476
rect 908 454 918 486
rect 662 436 918 454
rect 968 554 1020 564
rect 968 522 978 554
rect 1010 522 1020 554
rect 968 486 1020 522
rect 968 454 978 486
rect 1010 454 1020 486
rect 118 366 238 376
rect 118 334 128 366
rect 160 334 196 366
rect 228 334 238 366
rect 118 312 238 334
rect 424 366 544 376
rect 424 334 434 366
rect 466 334 502 366
rect 534 334 544 366
rect 424 312 544 334
rect 628 366 748 376
rect 628 334 638 366
rect 670 334 706 366
rect 738 334 748 366
rect 628 312 748 334
rect 805 366 928 376
rect 805 334 886 366
rect 918 334 928 366
rect 805 312 928 334
rect 968 368 1020 454
rect 1070 554 1122 590
rect 1070 522 1080 554
rect 1112 522 1122 554
rect 1070 486 1122 522
rect 1070 454 1080 486
rect 1112 454 1122 486
rect 1070 416 1122 454
rect 968 304 1097 368
rect 968 270 1020 304
rect 50 254 102 264
rect 50 222 60 254
rect 92 222 102 254
rect 50 186 102 222
rect 50 154 60 186
rect 92 154 102 186
rect 50 44 102 154
rect 152 254 1020 270
rect 152 222 162 254
rect 194 232 468 254
rect 194 222 204 232
rect 152 186 204 222
rect 458 222 468 232
rect 500 232 672 254
rect 500 222 510 232
rect 152 154 162 186
rect 194 154 204 186
rect 152 144 204 154
rect 254 186 408 196
rect 254 154 264 186
rect 296 154 366 186
rect 398 154 408 186
rect 254 44 408 154
rect 458 186 510 222
rect 662 222 672 232
rect 704 232 978 254
rect 704 222 714 232
rect 458 154 468 186
rect 500 154 510 186
rect 458 144 510 154
rect 560 186 612 196
rect 560 154 570 186
rect 602 154 612 186
rect 560 44 612 154
rect 662 186 714 222
rect 968 222 978 232
rect 1010 222 1020 254
rect 662 154 672 186
rect 704 154 714 186
rect 662 144 714 154
rect 764 186 918 196
rect 764 154 774 186
rect 806 154 876 186
rect 908 154 918 186
rect 764 44 918 154
rect 968 186 1020 222
rect 968 154 978 186
rect 1010 154 1020 186
rect 968 144 1020 154
rect 1070 254 1122 264
rect 1070 222 1080 254
rect 1112 222 1122 254
rect 1070 186 1122 222
rect 1070 154 1080 186
rect 1112 154 1122 186
rect 1070 44 1122 154
rect 0 16 1152 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1152 16
rect 0 -44 1152 -16
<< labels >>
flabel metal1 s 1020 304 1097 368 0 FreeSans 500 0 0 0 Y
port 2 nsew
flabel metal1 s 0 -44 1152 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 805 312 928 376 0 FreeSans 500 0 0 0 D
port 4 nsew
flabel metal1 s 0 712 1152 800 0 FreeSans 500 0 0 0 VDD
port 5 nsew
flabel metal1 s 424 312 544 376 0 FreeSans 500 0 0 0 B
port 6 nsew
flabel metal1 s 118 312 238 376 0 FreeSans 500 0 0 0 A
port 7 nsew
flabel metal1 s 255 756 255 756 0 FreeSans 400 0 0 0 VDD
flabel metal1 s 417 1 417 1 0 FreeSans 500 0 0 0 VSS
flabel metal1 s 628 312 748 376 0 FreeSans 500 0 0 0 C
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 756
string GDS_END 182242
string GDS_FILE 6_final.gds
string GDS_START 174016
<< end >>
