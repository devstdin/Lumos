magic
tech ihp-sg13g2
timestamp 1749416725
<< error_p >>
rect -18 1622 -13 1627
rect 13 1622 18 1627
rect 140 1622 145 1627
rect 171 1622 176 1627
rect 298 1622 303 1627
rect 329 1622 334 1627
rect 456 1622 461 1627
rect 487 1622 492 1627
rect 614 1622 619 1627
rect 645 1622 650 1627
rect 772 1622 777 1627
rect 803 1622 808 1627
rect 930 1622 935 1627
rect 961 1622 966 1627
rect 1088 1622 1093 1627
rect 1119 1622 1124 1627
rect 1246 1622 1251 1627
rect 1277 1622 1282 1627
rect 1404 1622 1409 1627
rect 1435 1622 1440 1627
rect 1562 1622 1567 1627
rect 1593 1622 1598 1627
rect 1720 1622 1725 1627
rect 1751 1622 1756 1627
rect 1878 1622 1883 1627
rect 1909 1622 1914 1627
rect 2036 1622 2041 1627
rect 2067 1622 2072 1627
rect 2194 1622 2199 1627
rect 2225 1622 2230 1627
rect 2352 1622 2357 1627
rect 2383 1622 2388 1627
rect 2510 1622 2515 1627
rect 2541 1622 2546 1627
rect 2668 1622 2673 1627
rect 2699 1622 2704 1627
rect 2826 1622 2831 1627
rect 2857 1622 2862 1627
rect 2984 1622 2989 1627
rect 3015 1622 3020 1627
rect -23 1617 23 1622
rect 135 1617 181 1622
rect 293 1617 339 1622
rect 451 1617 497 1622
rect 609 1617 655 1622
rect 767 1617 813 1622
rect 925 1617 971 1622
rect 1083 1617 1129 1622
rect 1241 1617 1287 1622
rect 1399 1617 1445 1622
rect 1557 1617 1603 1622
rect 1715 1617 1761 1622
rect 1873 1617 1919 1622
rect 2031 1617 2077 1622
rect 2189 1617 2235 1622
rect 2347 1617 2393 1622
rect 2505 1617 2551 1622
rect 2663 1617 2709 1622
rect 2821 1617 2867 1622
rect 2979 1617 3025 1622
rect -18 1611 18 1617
rect 140 1611 176 1617
rect 298 1611 334 1617
rect 456 1611 492 1617
rect 614 1611 650 1617
rect 772 1611 808 1617
rect 930 1611 966 1617
rect 1088 1611 1124 1617
rect 1246 1611 1282 1617
rect 1404 1611 1440 1617
rect 1562 1611 1598 1617
rect 1720 1611 1756 1617
rect 1878 1611 1914 1617
rect 2036 1611 2072 1617
rect 2194 1611 2230 1617
rect 2352 1611 2388 1617
rect 2510 1611 2546 1617
rect 2668 1611 2704 1617
rect 2826 1611 2862 1617
rect 2984 1611 3020 1617
rect -23 1606 23 1611
rect 135 1606 181 1611
rect 293 1606 339 1611
rect 451 1606 497 1611
rect 609 1606 655 1611
rect 767 1606 813 1611
rect 925 1606 971 1611
rect 1083 1606 1129 1611
rect 1241 1606 1287 1611
rect 1399 1606 1445 1611
rect 1557 1606 1603 1611
rect 1715 1606 1761 1611
rect 1873 1606 1919 1611
rect 2031 1606 2077 1611
rect 2189 1606 2235 1611
rect 2347 1606 2393 1611
rect 2505 1606 2551 1611
rect 2663 1606 2709 1611
rect 2821 1606 2867 1611
rect 2979 1606 3025 1611
rect -18 1601 -13 1606
rect 13 1601 18 1606
rect 140 1601 145 1606
rect 171 1601 176 1606
rect 298 1601 303 1606
rect 329 1601 334 1606
rect 456 1601 461 1606
rect 487 1601 492 1606
rect 614 1601 619 1606
rect 645 1601 650 1606
rect 772 1601 777 1606
rect 803 1601 808 1606
rect 930 1601 935 1606
rect 961 1601 966 1606
rect 1088 1601 1093 1606
rect 1119 1601 1124 1606
rect 1246 1601 1251 1606
rect 1277 1601 1282 1606
rect 1404 1601 1409 1606
rect 1435 1601 1440 1606
rect 1562 1601 1567 1606
rect 1593 1601 1598 1606
rect 1720 1601 1725 1606
rect 1751 1601 1756 1606
rect 1878 1601 1883 1606
rect 1909 1601 1914 1606
rect 2036 1601 2041 1606
rect 2067 1601 2072 1606
rect 2194 1601 2199 1606
rect 2225 1601 2230 1606
rect 2352 1601 2357 1606
rect 2383 1601 2388 1606
rect 2510 1601 2515 1606
rect 2541 1601 2546 1606
rect 2668 1601 2673 1606
rect 2699 1601 2704 1606
rect 2826 1601 2831 1606
rect 2857 1601 2862 1606
rect 2984 1601 2989 1606
rect 3015 1601 3020 1606
rect -52 1585 -47 1590
rect -41 1585 -36 1590
rect 36 1585 41 1590
rect 47 1585 52 1590
rect 106 1585 111 1590
rect 117 1585 122 1590
rect 194 1585 199 1590
rect 205 1585 210 1590
rect 264 1585 269 1590
rect 275 1585 280 1590
rect 352 1585 357 1590
rect 363 1585 368 1590
rect 422 1585 427 1590
rect 433 1585 438 1590
rect 510 1585 515 1590
rect 521 1585 526 1590
rect 580 1585 585 1590
rect 591 1585 596 1590
rect 668 1585 673 1590
rect 679 1585 684 1590
rect 738 1585 743 1590
rect 749 1585 754 1590
rect 826 1585 831 1590
rect 837 1585 842 1590
rect 896 1585 901 1590
rect 907 1585 912 1590
rect 984 1585 989 1590
rect 995 1585 1000 1590
rect 1054 1585 1059 1590
rect 1065 1585 1070 1590
rect 1142 1585 1147 1590
rect 1153 1585 1158 1590
rect 1212 1585 1217 1590
rect 1223 1585 1228 1590
rect 1300 1585 1305 1590
rect 1311 1585 1316 1590
rect 1370 1585 1375 1590
rect 1381 1585 1386 1590
rect 1458 1585 1463 1590
rect 1469 1585 1474 1590
rect 1528 1585 1533 1590
rect 1539 1585 1544 1590
rect 1616 1585 1621 1590
rect 1627 1585 1632 1590
rect 1686 1585 1691 1590
rect 1697 1585 1702 1590
rect 1774 1585 1779 1590
rect 1785 1585 1790 1590
rect 1844 1585 1849 1590
rect 1855 1585 1860 1590
rect 1932 1585 1937 1590
rect 1943 1585 1948 1590
rect 2002 1585 2007 1590
rect 2013 1585 2018 1590
rect 2090 1585 2095 1590
rect 2101 1585 2106 1590
rect 2160 1585 2165 1590
rect 2171 1585 2176 1590
rect 2248 1585 2253 1590
rect 2259 1585 2264 1590
rect 2318 1585 2323 1590
rect 2329 1585 2334 1590
rect 2406 1585 2411 1590
rect 2417 1585 2422 1590
rect 2476 1585 2481 1590
rect 2487 1585 2492 1590
rect 2564 1585 2569 1590
rect 2575 1585 2580 1590
rect 2634 1585 2639 1590
rect 2645 1585 2650 1590
rect 2722 1585 2727 1590
rect 2733 1585 2738 1590
rect 2792 1585 2797 1590
rect 2803 1585 2808 1590
rect 2880 1585 2885 1590
rect 2891 1585 2896 1590
rect 2950 1585 2955 1590
rect 2961 1585 2966 1590
rect 3038 1585 3043 1590
rect 3049 1585 3054 1590
rect -57 1580 -52 1585
rect -36 1580 -31 1585
rect 31 1580 36 1585
rect 52 1580 57 1585
rect 101 1580 106 1585
rect 122 1580 127 1585
rect 189 1580 194 1585
rect 210 1580 215 1585
rect 259 1580 264 1585
rect 280 1580 285 1585
rect 347 1580 352 1585
rect 368 1580 373 1585
rect 417 1580 422 1585
rect 438 1580 443 1585
rect 505 1580 510 1585
rect 526 1580 531 1585
rect 575 1580 580 1585
rect 596 1580 601 1585
rect 663 1580 668 1585
rect 684 1580 689 1585
rect 733 1580 738 1585
rect 754 1580 759 1585
rect 821 1580 826 1585
rect 842 1580 847 1585
rect 891 1580 896 1585
rect 912 1580 917 1585
rect 979 1580 984 1585
rect 1000 1580 1005 1585
rect 1049 1580 1054 1585
rect 1070 1580 1075 1585
rect 1137 1580 1142 1585
rect 1158 1580 1163 1585
rect 1207 1580 1212 1585
rect 1228 1580 1233 1585
rect 1295 1580 1300 1585
rect 1316 1580 1321 1585
rect 1365 1580 1370 1585
rect 1386 1580 1391 1585
rect 1453 1580 1458 1585
rect 1474 1580 1479 1585
rect 1523 1580 1528 1585
rect 1544 1580 1549 1585
rect 1611 1580 1616 1585
rect 1632 1580 1637 1585
rect 1681 1580 1686 1585
rect 1702 1580 1707 1585
rect 1769 1580 1774 1585
rect 1790 1580 1795 1585
rect 1839 1580 1844 1585
rect 1860 1580 1865 1585
rect 1927 1580 1932 1585
rect 1948 1580 1953 1585
rect 1997 1580 2002 1585
rect 2018 1580 2023 1585
rect 2085 1580 2090 1585
rect 2106 1580 2111 1585
rect 2155 1580 2160 1585
rect 2176 1580 2181 1585
rect 2243 1580 2248 1585
rect 2264 1580 2269 1585
rect 2313 1580 2318 1585
rect 2334 1580 2339 1585
rect 2401 1580 2406 1585
rect 2422 1580 2427 1585
rect 2471 1580 2476 1585
rect 2492 1580 2497 1585
rect 2559 1580 2564 1585
rect 2580 1580 2585 1585
rect 2629 1580 2634 1585
rect 2650 1580 2655 1585
rect 2717 1580 2722 1585
rect 2738 1580 2743 1585
rect 2787 1580 2792 1585
rect 2808 1580 2813 1585
rect 2875 1580 2880 1585
rect 2896 1580 2901 1585
rect 2945 1580 2950 1585
rect 2966 1580 2971 1585
rect 3033 1580 3038 1585
rect 3054 1580 3059 1585
rect -57 599 -52 604
rect -36 599 -31 604
rect 31 599 36 604
rect 52 599 57 604
rect 101 599 106 604
rect 122 599 127 604
rect 189 599 194 604
rect 210 599 215 604
rect 259 599 264 604
rect 280 599 285 604
rect 347 599 352 604
rect 368 599 373 604
rect 417 599 422 604
rect 438 599 443 604
rect 505 599 510 604
rect 526 599 531 604
rect 575 599 580 604
rect 596 599 601 604
rect 663 599 668 604
rect 684 599 689 604
rect 733 599 738 604
rect 754 599 759 604
rect 821 599 826 604
rect 842 599 847 604
rect 891 599 896 604
rect 912 599 917 604
rect 979 599 984 604
rect 1000 599 1005 604
rect 1049 599 1054 604
rect 1070 599 1075 604
rect 1137 599 1142 604
rect 1158 599 1163 604
rect 1207 599 1212 604
rect 1228 599 1233 604
rect 1295 599 1300 604
rect 1316 599 1321 604
rect 1365 599 1370 604
rect 1386 599 1391 604
rect 1453 599 1458 604
rect 1474 599 1479 604
rect 1523 599 1528 604
rect 1544 599 1549 604
rect 1611 599 1616 604
rect 1632 599 1637 604
rect 1681 599 1686 604
rect 1702 599 1707 604
rect 1769 599 1774 604
rect 1790 599 1795 604
rect 1839 599 1844 604
rect 1860 599 1865 604
rect 1927 599 1932 604
rect 1948 599 1953 604
rect 1997 599 2002 604
rect 2018 599 2023 604
rect 2085 599 2090 604
rect 2106 599 2111 604
rect 2155 599 2160 604
rect 2176 599 2181 604
rect 2243 599 2248 604
rect 2264 599 2269 604
rect 2313 599 2318 604
rect 2334 599 2339 604
rect 2401 599 2406 604
rect 2422 599 2427 604
rect 2471 599 2476 604
rect 2492 599 2497 604
rect 2559 599 2564 604
rect 2580 599 2585 604
rect 2629 599 2634 604
rect 2650 599 2655 604
rect 2717 599 2722 604
rect 2738 599 2743 604
rect 2787 599 2792 604
rect 2808 599 2813 604
rect 2875 599 2880 604
rect 2896 599 2901 604
rect 2945 599 2950 604
rect 2966 599 2971 604
rect 3033 599 3038 604
rect 3054 599 3059 604
rect -52 594 -47 599
rect -41 594 -36 599
rect 36 594 41 599
rect 47 594 52 599
rect 106 594 111 599
rect 117 594 122 599
rect 194 594 199 599
rect 205 594 210 599
rect 264 594 269 599
rect 275 594 280 599
rect 352 594 357 599
rect 363 594 368 599
rect 422 594 427 599
rect 433 594 438 599
rect 510 594 515 599
rect 521 594 526 599
rect 580 594 585 599
rect 591 594 596 599
rect 668 594 673 599
rect 679 594 684 599
rect 738 594 743 599
rect 749 594 754 599
rect 826 594 831 599
rect 837 594 842 599
rect 896 594 901 599
rect 907 594 912 599
rect 984 594 989 599
rect 995 594 1000 599
rect 1054 594 1059 599
rect 1065 594 1070 599
rect 1142 594 1147 599
rect 1153 594 1158 599
rect 1212 594 1217 599
rect 1223 594 1228 599
rect 1300 594 1305 599
rect 1311 594 1316 599
rect 1370 594 1375 599
rect 1381 594 1386 599
rect 1458 594 1463 599
rect 1469 594 1474 599
rect 1528 594 1533 599
rect 1539 594 1544 599
rect 1616 594 1621 599
rect 1627 594 1632 599
rect 1686 594 1691 599
rect 1697 594 1702 599
rect 1774 594 1779 599
rect 1785 594 1790 599
rect 1844 594 1849 599
rect 1855 594 1860 599
rect 1932 594 1937 599
rect 1943 594 1948 599
rect 2002 594 2007 599
rect 2013 594 2018 599
rect 2090 594 2095 599
rect 2101 594 2106 599
rect 2160 594 2165 599
rect 2171 594 2176 599
rect 2248 594 2253 599
rect 2259 594 2264 599
rect 2318 594 2323 599
rect 2329 594 2334 599
rect 2406 594 2411 599
rect 2417 594 2422 599
rect 2476 594 2481 599
rect 2487 594 2492 599
rect 2564 594 2569 599
rect 2575 594 2580 599
rect 2634 594 2639 599
rect 2645 594 2650 599
rect 2722 594 2727 599
rect 2733 594 2738 599
rect 2792 594 2797 599
rect 2803 594 2808 599
rect 2880 594 2885 599
rect 2891 594 2896 599
rect 2950 594 2955 599
rect 2961 594 2966 599
rect 3038 594 3043 599
rect 3049 594 3054 599
rect -18 578 -13 583
rect 13 578 18 583
rect 140 578 145 583
rect 171 578 176 583
rect 298 578 303 583
rect 329 578 334 583
rect 456 578 461 583
rect 487 578 492 583
rect 614 578 619 583
rect 645 578 650 583
rect 772 578 777 583
rect 803 578 808 583
rect 930 578 935 583
rect 961 578 966 583
rect 1088 578 1093 583
rect 1119 578 1124 583
rect 1246 578 1251 583
rect 1277 578 1282 583
rect 1404 578 1409 583
rect 1435 578 1440 583
rect 1562 578 1567 583
rect 1593 578 1598 583
rect 1720 578 1725 583
rect 1751 578 1756 583
rect 1878 578 1883 583
rect 1909 578 1914 583
rect 2036 578 2041 583
rect 2067 578 2072 583
rect 2194 578 2199 583
rect 2225 578 2230 583
rect 2352 578 2357 583
rect 2383 578 2388 583
rect 2510 578 2515 583
rect 2541 578 2546 583
rect 2668 578 2673 583
rect 2699 578 2704 583
rect 2826 578 2831 583
rect 2857 578 2862 583
rect 2984 578 2989 583
rect 3015 578 3020 583
rect -23 573 23 578
rect 135 573 181 578
rect 293 573 339 578
rect 451 573 497 578
rect 609 573 655 578
rect 767 573 813 578
rect 925 573 971 578
rect 1083 573 1129 578
rect 1241 573 1287 578
rect 1399 573 1445 578
rect 1557 573 1603 578
rect 1715 573 1761 578
rect 1873 573 1919 578
rect 2031 573 2077 578
rect 2189 573 2235 578
rect 2347 573 2393 578
rect 2505 573 2551 578
rect 2663 573 2709 578
rect 2821 573 2867 578
rect 2979 573 3025 578
rect -18 567 18 573
rect 140 567 176 573
rect 298 567 334 573
rect 456 567 492 573
rect 614 567 650 573
rect 772 567 808 573
rect 930 567 966 573
rect 1088 567 1124 573
rect 1246 567 1282 573
rect 1404 567 1440 573
rect 1562 567 1598 573
rect 1720 567 1756 573
rect 1878 567 1914 573
rect 2036 567 2072 573
rect 2194 567 2230 573
rect 2352 567 2388 573
rect 2510 567 2546 573
rect 2668 567 2704 573
rect 2826 567 2862 573
rect 2984 567 3020 573
rect -23 562 23 567
rect 135 562 181 567
rect 293 562 339 567
rect 451 562 497 567
rect 609 562 655 567
rect 767 562 813 567
rect 925 562 971 567
rect 1083 562 1129 567
rect 1241 562 1287 567
rect 1399 562 1445 567
rect 1557 562 1603 567
rect 1715 562 1761 567
rect 1873 562 1919 567
rect 2031 562 2077 567
rect 2189 562 2235 567
rect 2347 562 2393 567
rect 2505 562 2551 567
rect 2663 562 2709 567
rect 2821 562 2867 567
rect 2979 562 3025 567
rect -18 557 -13 562
rect 13 557 18 562
rect 140 557 145 562
rect 171 557 176 562
rect 298 557 303 562
rect 329 557 334 562
rect 456 557 461 562
rect 487 557 492 562
rect 614 557 619 562
rect 645 557 650 562
rect 772 557 777 562
rect 803 557 808 562
rect 930 557 935 562
rect 961 557 966 562
rect 1088 557 1093 562
rect 1119 557 1124 562
rect 1246 557 1251 562
rect 1277 557 1282 562
rect 1404 557 1409 562
rect 1435 557 1440 562
rect 1562 557 1567 562
rect 1593 557 1598 562
rect 1720 557 1725 562
rect 1751 557 1756 562
rect 1878 557 1883 562
rect 1909 557 1914 562
rect 2036 557 2041 562
rect 2067 557 2072 562
rect 2194 557 2199 562
rect 2225 557 2230 562
rect 2352 557 2357 562
rect 2383 557 2388 562
rect 2510 557 2515 562
rect 2541 557 2546 562
rect 2668 557 2673 562
rect 2699 557 2704 562
rect 2826 557 2831 562
rect 2857 557 2862 562
rect 2984 557 2989 562
rect 3015 557 3020 562
rect -18 530 -13 535
rect 13 530 18 535
rect 140 530 145 535
rect 171 530 176 535
rect 298 530 303 535
rect 329 530 334 535
rect 456 530 461 535
rect 487 530 492 535
rect 614 530 619 535
rect 645 530 650 535
rect 772 530 777 535
rect 803 530 808 535
rect 930 530 935 535
rect 961 530 966 535
rect 1088 530 1093 535
rect 1119 530 1124 535
rect 1246 530 1251 535
rect 1277 530 1282 535
rect 1404 530 1409 535
rect 1435 530 1440 535
rect 1562 530 1567 535
rect 1593 530 1598 535
rect 1720 530 1725 535
rect 1751 530 1756 535
rect 1878 530 1883 535
rect 1909 530 1914 535
rect 2036 530 2041 535
rect 2067 530 2072 535
rect 2194 530 2199 535
rect 2225 530 2230 535
rect 2352 530 2357 535
rect 2383 530 2388 535
rect 2510 530 2515 535
rect 2541 530 2546 535
rect 2668 530 2673 535
rect 2699 530 2704 535
rect 2826 530 2831 535
rect 2857 530 2862 535
rect 2984 530 2989 535
rect 3015 530 3020 535
rect -23 525 23 530
rect 135 525 181 530
rect 293 525 339 530
rect 451 525 497 530
rect 609 525 655 530
rect 767 525 813 530
rect 925 525 971 530
rect 1083 525 1129 530
rect 1241 525 1287 530
rect 1399 525 1445 530
rect 1557 525 1603 530
rect 1715 525 1761 530
rect 1873 525 1919 530
rect 2031 525 2077 530
rect 2189 525 2235 530
rect 2347 525 2393 530
rect 2505 525 2551 530
rect 2663 525 2709 530
rect 2821 525 2867 530
rect 2979 525 3025 530
rect -18 519 18 525
rect 140 519 176 525
rect 298 519 334 525
rect 456 519 492 525
rect 614 519 650 525
rect 772 519 808 525
rect 930 519 966 525
rect 1088 519 1124 525
rect 1246 519 1282 525
rect 1404 519 1440 525
rect 1562 519 1598 525
rect 1720 519 1756 525
rect 1878 519 1914 525
rect 2036 519 2072 525
rect 2194 519 2230 525
rect 2352 519 2388 525
rect 2510 519 2546 525
rect 2668 519 2704 525
rect 2826 519 2862 525
rect 2984 519 3020 525
rect -23 514 23 519
rect 135 514 181 519
rect 293 514 339 519
rect 451 514 497 519
rect 609 514 655 519
rect 767 514 813 519
rect 925 514 971 519
rect 1083 514 1129 519
rect 1241 514 1287 519
rect 1399 514 1445 519
rect 1557 514 1603 519
rect 1715 514 1761 519
rect 1873 514 1919 519
rect 2031 514 2077 519
rect 2189 514 2235 519
rect 2347 514 2393 519
rect 2505 514 2551 519
rect 2663 514 2709 519
rect 2821 514 2867 519
rect 2979 514 3025 519
rect -18 509 -13 514
rect 13 509 18 514
rect 140 509 145 514
rect 171 509 176 514
rect 298 509 303 514
rect 329 509 334 514
rect 456 509 461 514
rect 487 509 492 514
rect 614 509 619 514
rect 645 509 650 514
rect 772 509 777 514
rect 803 509 808 514
rect 930 509 935 514
rect 961 509 966 514
rect 1088 509 1093 514
rect 1119 509 1124 514
rect 1246 509 1251 514
rect 1277 509 1282 514
rect 1404 509 1409 514
rect 1435 509 1440 514
rect 1562 509 1567 514
rect 1593 509 1598 514
rect 1720 509 1725 514
rect 1751 509 1756 514
rect 1878 509 1883 514
rect 1909 509 1914 514
rect 2036 509 2041 514
rect 2067 509 2072 514
rect 2194 509 2199 514
rect 2225 509 2230 514
rect 2352 509 2357 514
rect 2383 509 2388 514
rect 2510 509 2515 514
rect 2541 509 2546 514
rect 2668 509 2673 514
rect 2699 509 2704 514
rect 2826 509 2831 514
rect 2857 509 2862 514
rect 2984 509 2989 514
rect 3015 509 3020 514
rect -52 493 -47 498
rect -41 493 -36 498
rect 36 493 41 498
rect 47 493 52 498
rect 106 493 111 498
rect 117 493 122 498
rect 194 493 199 498
rect 205 493 210 498
rect 264 493 269 498
rect 275 493 280 498
rect 352 493 357 498
rect 363 493 368 498
rect 422 493 427 498
rect 433 493 438 498
rect 510 493 515 498
rect 521 493 526 498
rect 580 493 585 498
rect 591 493 596 498
rect 668 493 673 498
rect 679 493 684 498
rect 738 493 743 498
rect 749 493 754 498
rect 826 493 831 498
rect 837 493 842 498
rect 896 493 901 498
rect 907 493 912 498
rect 984 493 989 498
rect 995 493 1000 498
rect 1054 493 1059 498
rect 1065 493 1070 498
rect 1142 493 1147 498
rect 1153 493 1158 498
rect 1212 493 1217 498
rect 1223 493 1228 498
rect 1300 493 1305 498
rect 1311 493 1316 498
rect 1370 493 1375 498
rect 1381 493 1386 498
rect 1458 493 1463 498
rect 1469 493 1474 498
rect 1528 493 1533 498
rect 1539 493 1544 498
rect 1616 493 1621 498
rect 1627 493 1632 498
rect 1686 493 1691 498
rect 1697 493 1702 498
rect 1774 493 1779 498
rect 1785 493 1790 498
rect 1844 493 1849 498
rect 1855 493 1860 498
rect 1932 493 1937 498
rect 1943 493 1948 498
rect 2002 493 2007 498
rect 2013 493 2018 498
rect 2090 493 2095 498
rect 2101 493 2106 498
rect 2160 493 2165 498
rect 2171 493 2176 498
rect 2248 493 2253 498
rect 2259 493 2264 498
rect 2318 493 2323 498
rect 2329 493 2334 498
rect 2406 493 2411 498
rect 2417 493 2422 498
rect 2476 493 2481 498
rect 2487 493 2492 498
rect 2564 493 2569 498
rect 2575 493 2580 498
rect 2634 493 2639 498
rect 2645 493 2650 498
rect 2722 493 2727 498
rect 2733 493 2738 498
rect 2792 493 2797 498
rect 2803 493 2808 498
rect 2880 493 2885 498
rect 2891 493 2896 498
rect 2950 493 2955 498
rect 2961 493 2966 498
rect 3038 493 3043 498
rect 3049 493 3054 498
rect -57 488 -52 493
rect -36 488 -31 493
rect 31 488 36 493
rect 52 488 57 493
rect 101 488 106 493
rect 122 488 127 493
rect 189 488 194 493
rect 210 488 215 493
rect 259 488 264 493
rect 280 488 285 493
rect 347 488 352 493
rect 368 488 373 493
rect 417 488 422 493
rect 438 488 443 493
rect 505 488 510 493
rect 526 488 531 493
rect 575 488 580 493
rect 596 488 601 493
rect 663 488 668 493
rect 684 488 689 493
rect 733 488 738 493
rect 754 488 759 493
rect 821 488 826 493
rect 842 488 847 493
rect 891 488 896 493
rect 912 488 917 493
rect 979 488 984 493
rect 1000 488 1005 493
rect 1049 488 1054 493
rect 1070 488 1075 493
rect 1137 488 1142 493
rect 1158 488 1163 493
rect 1207 488 1212 493
rect 1228 488 1233 493
rect 1295 488 1300 493
rect 1316 488 1321 493
rect 1365 488 1370 493
rect 1386 488 1391 493
rect 1453 488 1458 493
rect 1474 488 1479 493
rect 1523 488 1528 493
rect 1544 488 1549 493
rect 1611 488 1616 493
rect 1632 488 1637 493
rect 1681 488 1686 493
rect 1702 488 1707 493
rect 1769 488 1774 493
rect 1790 488 1795 493
rect 1839 488 1844 493
rect 1860 488 1865 493
rect 1927 488 1932 493
rect 1948 488 1953 493
rect 1997 488 2002 493
rect 2018 488 2023 493
rect 2085 488 2090 493
rect 2106 488 2111 493
rect 2155 488 2160 493
rect 2176 488 2181 493
rect 2243 488 2248 493
rect 2264 488 2269 493
rect 2313 488 2318 493
rect 2334 488 2339 493
rect 2401 488 2406 493
rect 2422 488 2427 493
rect 2471 488 2476 493
rect 2492 488 2497 493
rect 2559 488 2564 493
rect 2580 488 2585 493
rect 2629 488 2634 493
rect 2650 488 2655 493
rect 2717 488 2722 493
rect 2738 488 2743 493
rect 2787 488 2792 493
rect 2808 488 2813 493
rect 2875 488 2880 493
rect 2896 488 2901 493
rect 2945 488 2950 493
rect 2966 488 2971 493
rect 3033 488 3038 493
rect 3054 488 3059 493
rect -57 -493 -52 -488
rect -36 -493 -31 -488
rect 31 -493 36 -488
rect 52 -493 57 -488
rect 101 -493 106 -488
rect 122 -493 127 -488
rect 189 -493 194 -488
rect 210 -493 215 -488
rect 259 -493 264 -488
rect 280 -493 285 -488
rect 347 -493 352 -488
rect 368 -493 373 -488
rect 417 -493 422 -488
rect 438 -493 443 -488
rect 505 -493 510 -488
rect 526 -493 531 -488
rect 575 -493 580 -488
rect 596 -493 601 -488
rect 663 -493 668 -488
rect 684 -493 689 -488
rect 733 -493 738 -488
rect 754 -493 759 -488
rect 821 -493 826 -488
rect 842 -493 847 -488
rect 891 -493 896 -488
rect 912 -493 917 -488
rect 979 -493 984 -488
rect 1000 -493 1005 -488
rect 1049 -493 1054 -488
rect 1070 -493 1075 -488
rect 1137 -493 1142 -488
rect 1158 -493 1163 -488
rect 1207 -493 1212 -488
rect 1228 -493 1233 -488
rect 1295 -493 1300 -488
rect 1316 -493 1321 -488
rect 1365 -493 1370 -488
rect 1386 -493 1391 -488
rect 1453 -493 1458 -488
rect 1474 -493 1479 -488
rect 1523 -493 1528 -488
rect 1544 -493 1549 -488
rect 1611 -493 1616 -488
rect 1632 -493 1637 -488
rect 1681 -493 1686 -488
rect 1702 -493 1707 -488
rect 1769 -493 1774 -488
rect 1790 -493 1795 -488
rect 1839 -493 1844 -488
rect 1860 -493 1865 -488
rect 1927 -493 1932 -488
rect 1948 -493 1953 -488
rect 1997 -493 2002 -488
rect 2018 -493 2023 -488
rect 2085 -493 2090 -488
rect 2106 -493 2111 -488
rect 2155 -493 2160 -488
rect 2176 -493 2181 -488
rect 2243 -493 2248 -488
rect 2264 -493 2269 -488
rect 2313 -493 2318 -488
rect 2334 -493 2339 -488
rect 2401 -493 2406 -488
rect 2422 -493 2427 -488
rect 2471 -493 2476 -488
rect 2492 -493 2497 -488
rect 2559 -493 2564 -488
rect 2580 -493 2585 -488
rect 2629 -493 2634 -488
rect 2650 -493 2655 -488
rect 2717 -493 2722 -488
rect 2738 -493 2743 -488
rect 2787 -493 2792 -488
rect 2808 -493 2813 -488
rect 2875 -493 2880 -488
rect 2896 -493 2901 -488
rect 2945 -493 2950 -488
rect 2966 -493 2971 -488
rect 3033 -493 3038 -488
rect 3054 -493 3059 -488
rect -52 -498 -47 -493
rect -41 -498 -36 -493
rect 36 -498 41 -493
rect 47 -498 52 -493
rect 106 -498 111 -493
rect 117 -498 122 -493
rect 194 -498 199 -493
rect 205 -498 210 -493
rect 264 -498 269 -493
rect 275 -498 280 -493
rect 352 -498 357 -493
rect 363 -498 368 -493
rect 422 -498 427 -493
rect 433 -498 438 -493
rect 510 -498 515 -493
rect 521 -498 526 -493
rect 580 -498 585 -493
rect 591 -498 596 -493
rect 668 -498 673 -493
rect 679 -498 684 -493
rect 738 -498 743 -493
rect 749 -498 754 -493
rect 826 -498 831 -493
rect 837 -498 842 -493
rect 896 -498 901 -493
rect 907 -498 912 -493
rect 984 -498 989 -493
rect 995 -498 1000 -493
rect 1054 -498 1059 -493
rect 1065 -498 1070 -493
rect 1142 -498 1147 -493
rect 1153 -498 1158 -493
rect 1212 -498 1217 -493
rect 1223 -498 1228 -493
rect 1300 -498 1305 -493
rect 1311 -498 1316 -493
rect 1370 -498 1375 -493
rect 1381 -498 1386 -493
rect 1458 -498 1463 -493
rect 1469 -498 1474 -493
rect 1528 -498 1533 -493
rect 1539 -498 1544 -493
rect 1616 -498 1621 -493
rect 1627 -498 1632 -493
rect 1686 -498 1691 -493
rect 1697 -498 1702 -493
rect 1774 -498 1779 -493
rect 1785 -498 1790 -493
rect 1844 -498 1849 -493
rect 1855 -498 1860 -493
rect 1932 -498 1937 -493
rect 1943 -498 1948 -493
rect 2002 -498 2007 -493
rect 2013 -498 2018 -493
rect 2090 -498 2095 -493
rect 2101 -498 2106 -493
rect 2160 -498 2165 -493
rect 2171 -498 2176 -493
rect 2248 -498 2253 -493
rect 2259 -498 2264 -493
rect 2318 -498 2323 -493
rect 2329 -498 2334 -493
rect 2406 -498 2411 -493
rect 2417 -498 2422 -493
rect 2476 -498 2481 -493
rect 2487 -498 2492 -493
rect 2564 -498 2569 -493
rect 2575 -498 2580 -493
rect 2634 -498 2639 -493
rect 2645 -498 2650 -493
rect 2722 -498 2727 -493
rect 2733 -498 2738 -493
rect 2792 -498 2797 -493
rect 2803 -498 2808 -493
rect 2880 -498 2885 -493
rect 2891 -498 2896 -493
rect 2950 -498 2955 -493
rect 2961 -498 2966 -493
rect 3038 -498 3043 -493
rect 3049 -498 3054 -493
rect -18 -514 -13 -509
rect 13 -514 18 -509
rect 140 -514 145 -509
rect 171 -514 176 -509
rect 298 -514 303 -509
rect 329 -514 334 -509
rect 456 -514 461 -509
rect 487 -514 492 -509
rect 614 -514 619 -509
rect 645 -514 650 -509
rect 772 -514 777 -509
rect 803 -514 808 -509
rect 930 -514 935 -509
rect 961 -514 966 -509
rect 1088 -514 1093 -509
rect 1119 -514 1124 -509
rect 1246 -514 1251 -509
rect 1277 -514 1282 -509
rect 1404 -514 1409 -509
rect 1435 -514 1440 -509
rect 1562 -514 1567 -509
rect 1593 -514 1598 -509
rect 1720 -514 1725 -509
rect 1751 -514 1756 -509
rect 1878 -514 1883 -509
rect 1909 -514 1914 -509
rect 2036 -514 2041 -509
rect 2067 -514 2072 -509
rect 2194 -514 2199 -509
rect 2225 -514 2230 -509
rect 2352 -514 2357 -509
rect 2383 -514 2388 -509
rect 2510 -514 2515 -509
rect 2541 -514 2546 -509
rect 2668 -514 2673 -509
rect 2699 -514 2704 -509
rect 2826 -514 2831 -509
rect 2857 -514 2862 -509
rect 2984 -514 2989 -509
rect 3015 -514 3020 -509
rect -23 -519 23 -514
rect 135 -519 181 -514
rect 293 -519 339 -514
rect 451 -519 497 -514
rect 609 -519 655 -514
rect 767 -519 813 -514
rect 925 -519 971 -514
rect 1083 -519 1129 -514
rect 1241 -519 1287 -514
rect 1399 -519 1445 -514
rect 1557 -519 1603 -514
rect 1715 -519 1761 -514
rect 1873 -519 1919 -514
rect 2031 -519 2077 -514
rect 2189 -519 2235 -514
rect 2347 -519 2393 -514
rect 2505 -519 2551 -514
rect 2663 -519 2709 -514
rect 2821 -519 2867 -514
rect 2979 -519 3025 -514
rect -18 -525 18 -519
rect 140 -525 176 -519
rect 298 -525 334 -519
rect 456 -525 492 -519
rect 614 -525 650 -519
rect 772 -525 808 -519
rect 930 -525 966 -519
rect 1088 -525 1124 -519
rect 1246 -525 1282 -519
rect 1404 -525 1440 -519
rect 1562 -525 1598 -519
rect 1720 -525 1756 -519
rect 1878 -525 1914 -519
rect 2036 -525 2072 -519
rect 2194 -525 2230 -519
rect 2352 -525 2388 -519
rect 2510 -525 2546 -519
rect 2668 -525 2704 -519
rect 2826 -525 2862 -519
rect 2984 -525 3020 -519
rect -23 -530 23 -525
rect 135 -530 181 -525
rect 293 -530 339 -525
rect 451 -530 497 -525
rect 609 -530 655 -525
rect 767 -530 813 -525
rect 925 -530 971 -525
rect 1083 -530 1129 -525
rect 1241 -530 1287 -525
rect 1399 -530 1445 -525
rect 1557 -530 1603 -525
rect 1715 -530 1761 -525
rect 1873 -530 1919 -525
rect 2031 -530 2077 -525
rect 2189 -530 2235 -525
rect 2347 -530 2393 -525
rect 2505 -530 2551 -525
rect 2663 -530 2709 -525
rect 2821 -530 2867 -525
rect 2979 -530 3025 -525
rect -18 -535 -13 -530
rect 13 -535 18 -530
rect 140 -535 145 -530
rect 171 -535 176 -530
rect 298 -535 303 -530
rect 329 -535 334 -530
rect 456 -535 461 -530
rect 487 -535 492 -530
rect 614 -535 619 -530
rect 645 -535 650 -530
rect 772 -535 777 -530
rect 803 -535 808 -530
rect 930 -535 935 -530
rect 961 -535 966 -530
rect 1088 -535 1093 -530
rect 1119 -535 1124 -530
rect 1246 -535 1251 -530
rect 1277 -535 1282 -530
rect 1404 -535 1409 -530
rect 1435 -535 1440 -530
rect 1562 -535 1567 -530
rect 1593 -535 1598 -530
rect 1720 -535 1725 -530
rect 1751 -535 1756 -530
rect 1878 -535 1883 -530
rect 1909 -535 1914 -530
rect 2036 -535 2041 -530
rect 2067 -535 2072 -530
rect 2194 -535 2199 -530
rect 2225 -535 2230 -530
rect 2352 -535 2357 -530
rect 2383 -535 2388 -530
rect 2510 -535 2515 -530
rect 2541 -535 2546 -530
rect 2668 -535 2673 -530
rect 2699 -535 2704 -530
rect 2826 -535 2831 -530
rect 2857 -535 2862 -530
rect 2984 -535 2989 -530
rect 3015 -535 3020 -530
<< nwell >>
rect -205 -651 3207 1743
<< hvpmos >>
rect -25 592 25 1592
rect 133 592 183 1592
rect 291 592 341 1592
rect 449 592 499 1592
rect 607 592 657 1592
rect 765 592 815 1592
rect 923 592 973 1592
rect 1081 592 1131 1592
rect 1239 592 1289 1592
rect 1397 592 1447 1592
rect 1555 592 1605 1592
rect 1713 592 1763 1592
rect 1871 592 1921 1592
rect 2029 592 2079 1592
rect 2187 592 2237 1592
rect 2345 592 2395 1592
rect 2503 592 2553 1592
rect 2661 592 2711 1592
rect 2819 592 2869 1592
rect 2977 592 3027 1592
rect -25 -500 25 500
rect 133 -500 183 500
rect 291 -500 341 500
rect 449 -500 499 500
rect 607 -500 657 500
rect 765 -500 815 500
rect 923 -500 973 500
rect 1081 -500 1131 500
rect 1239 -500 1289 500
rect 1397 -500 1447 500
rect 1555 -500 1605 500
rect 1713 -500 1763 500
rect 1871 -500 1921 500
rect 2029 -500 2079 500
rect 2187 -500 2237 500
rect 2345 -500 2395 500
rect 2503 -500 2553 500
rect 2661 -500 2711 500
rect 2819 -500 2869 500
rect 2977 -500 3027 500
<< hvpdiff >>
rect -59 1585 -25 1592
rect -59 599 -52 1585
rect -36 599 -25 1585
rect -59 592 -25 599
rect 25 1585 59 1592
rect 25 599 36 1585
rect 52 599 59 1585
rect 25 592 59 599
rect 99 1585 133 1592
rect 99 599 106 1585
rect 122 599 133 1585
rect 99 592 133 599
rect 183 1585 217 1592
rect 183 599 194 1585
rect 210 599 217 1585
rect 183 592 217 599
rect 257 1585 291 1592
rect 257 599 264 1585
rect 280 599 291 1585
rect 257 592 291 599
rect 341 1585 375 1592
rect 341 599 352 1585
rect 368 599 375 1585
rect 341 592 375 599
rect 415 1585 449 1592
rect 415 599 422 1585
rect 438 599 449 1585
rect 415 592 449 599
rect 499 1585 533 1592
rect 499 599 510 1585
rect 526 599 533 1585
rect 499 592 533 599
rect 573 1585 607 1592
rect 573 599 580 1585
rect 596 599 607 1585
rect 573 592 607 599
rect 657 1585 691 1592
rect 657 599 668 1585
rect 684 599 691 1585
rect 657 592 691 599
rect 731 1585 765 1592
rect 731 599 738 1585
rect 754 599 765 1585
rect 731 592 765 599
rect 815 1585 849 1592
rect 815 599 826 1585
rect 842 599 849 1585
rect 815 592 849 599
rect 889 1585 923 1592
rect 889 599 896 1585
rect 912 599 923 1585
rect 889 592 923 599
rect 973 1585 1007 1592
rect 973 599 984 1585
rect 1000 599 1007 1585
rect 973 592 1007 599
rect 1047 1585 1081 1592
rect 1047 599 1054 1585
rect 1070 599 1081 1585
rect 1047 592 1081 599
rect 1131 1585 1165 1592
rect 1131 599 1142 1585
rect 1158 599 1165 1585
rect 1131 592 1165 599
rect 1205 1585 1239 1592
rect 1205 599 1212 1585
rect 1228 599 1239 1585
rect 1205 592 1239 599
rect 1289 1585 1323 1592
rect 1289 599 1300 1585
rect 1316 599 1323 1585
rect 1289 592 1323 599
rect 1363 1585 1397 1592
rect 1363 599 1370 1585
rect 1386 599 1397 1585
rect 1363 592 1397 599
rect 1447 1585 1481 1592
rect 1447 599 1458 1585
rect 1474 599 1481 1585
rect 1447 592 1481 599
rect 1521 1585 1555 1592
rect 1521 599 1528 1585
rect 1544 599 1555 1585
rect 1521 592 1555 599
rect 1605 1585 1639 1592
rect 1605 599 1616 1585
rect 1632 599 1639 1585
rect 1605 592 1639 599
rect 1679 1585 1713 1592
rect 1679 599 1686 1585
rect 1702 599 1713 1585
rect 1679 592 1713 599
rect 1763 1585 1797 1592
rect 1763 599 1774 1585
rect 1790 599 1797 1585
rect 1763 592 1797 599
rect 1837 1585 1871 1592
rect 1837 599 1844 1585
rect 1860 599 1871 1585
rect 1837 592 1871 599
rect 1921 1585 1955 1592
rect 1921 599 1932 1585
rect 1948 599 1955 1585
rect 1921 592 1955 599
rect 1995 1585 2029 1592
rect 1995 599 2002 1585
rect 2018 599 2029 1585
rect 1995 592 2029 599
rect 2079 1585 2113 1592
rect 2079 599 2090 1585
rect 2106 599 2113 1585
rect 2079 592 2113 599
rect 2153 1585 2187 1592
rect 2153 599 2160 1585
rect 2176 599 2187 1585
rect 2153 592 2187 599
rect 2237 1585 2271 1592
rect 2237 599 2248 1585
rect 2264 599 2271 1585
rect 2237 592 2271 599
rect 2311 1585 2345 1592
rect 2311 599 2318 1585
rect 2334 599 2345 1585
rect 2311 592 2345 599
rect 2395 1585 2429 1592
rect 2395 599 2406 1585
rect 2422 599 2429 1585
rect 2395 592 2429 599
rect 2469 1585 2503 1592
rect 2469 599 2476 1585
rect 2492 599 2503 1585
rect 2469 592 2503 599
rect 2553 1585 2587 1592
rect 2553 599 2564 1585
rect 2580 599 2587 1585
rect 2553 592 2587 599
rect 2627 1585 2661 1592
rect 2627 599 2634 1585
rect 2650 599 2661 1585
rect 2627 592 2661 599
rect 2711 1585 2745 1592
rect 2711 599 2722 1585
rect 2738 599 2745 1585
rect 2711 592 2745 599
rect 2785 1585 2819 1592
rect 2785 599 2792 1585
rect 2808 599 2819 1585
rect 2785 592 2819 599
rect 2869 1585 2903 1592
rect 2869 599 2880 1585
rect 2896 599 2903 1585
rect 2869 592 2903 599
rect 2943 1585 2977 1592
rect 2943 599 2950 1585
rect 2966 599 2977 1585
rect 2943 592 2977 599
rect 3027 1585 3061 1592
rect 3027 599 3038 1585
rect 3054 599 3061 1585
rect 3027 592 3061 599
rect -59 493 -25 500
rect -59 -493 -52 493
rect -36 -493 -25 493
rect -59 -500 -25 -493
rect 25 493 59 500
rect 25 -493 36 493
rect 52 -493 59 493
rect 25 -500 59 -493
rect 99 493 133 500
rect 99 -493 106 493
rect 122 -493 133 493
rect 99 -500 133 -493
rect 183 493 217 500
rect 183 -493 194 493
rect 210 -493 217 493
rect 183 -500 217 -493
rect 257 493 291 500
rect 257 -493 264 493
rect 280 -493 291 493
rect 257 -500 291 -493
rect 341 493 375 500
rect 341 -493 352 493
rect 368 -493 375 493
rect 341 -500 375 -493
rect 415 493 449 500
rect 415 -493 422 493
rect 438 -493 449 493
rect 415 -500 449 -493
rect 499 493 533 500
rect 499 -493 510 493
rect 526 -493 533 493
rect 499 -500 533 -493
rect 573 493 607 500
rect 573 -493 580 493
rect 596 -493 607 493
rect 573 -500 607 -493
rect 657 493 691 500
rect 657 -493 668 493
rect 684 -493 691 493
rect 657 -500 691 -493
rect 731 493 765 500
rect 731 -493 738 493
rect 754 -493 765 493
rect 731 -500 765 -493
rect 815 493 849 500
rect 815 -493 826 493
rect 842 -493 849 493
rect 815 -500 849 -493
rect 889 493 923 500
rect 889 -493 896 493
rect 912 -493 923 493
rect 889 -500 923 -493
rect 973 493 1007 500
rect 973 -493 984 493
rect 1000 -493 1007 493
rect 973 -500 1007 -493
rect 1047 493 1081 500
rect 1047 -493 1054 493
rect 1070 -493 1081 493
rect 1047 -500 1081 -493
rect 1131 493 1165 500
rect 1131 -493 1142 493
rect 1158 -493 1165 493
rect 1131 -500 1165 -493
rect 1205 493 1239 500
rect 1205 -493 1212 493
rect 1228 -493 1239 493
rect 1205 -500 1239 -493
rect 1289 493 1323 500
rect 1289 -493 1300 493
rect 1316 -493 1323 493
rect 1289 -500 1323 -493
rect 1363 493 1397 500
rect 1363 -493 1370 493
rect 1386 -493 1397 493
rect 1363 -500 1397 -493
rect 1447 493 1481 500
rect 1447 -493 1458 493
rect 1474 -493 1481 493
rect 1447 -500 1481 -493
rect 1521 493 1555 500
rect 1521 -493 1528 493
rect 1544 -493 1555 493
rect 1521 -500 1555 -493
rect 1605 493 1639 500
rect 1605 -493 1616 493
rect 1632 -493 1639 493
rect 1605 -500 1639 -493
rect 1679 493 1713 500
rect 1679 -493 1686 493
rect 1702 -493 1713 493
rect 1679 -500 1713 -493
rect 1763 493 1797 500
rect 1763 -493 1774 493
rect 1790 -493 1797 493
rect 1763 -500 1797 -493
rect 1837 493 1871 500
rect 1837 -493 1844 493
rect 1860 -493 1871 493
rect 1837 -500 1871 -493
rect 1921 493 1955 500
rect 1921 -493 1932 493
rect 1948 -493 1955 493
rect 1921 -500 1955 -493
rect 1995 493 2029 500
rect 1995 -493 2002 493
rect 2018 -493 2029 493
rect 1995 -500 2029 -493
rect 2079 493 2113 500
rect 2079 -493 2090 493
rect 2106 -493 2113 493
rect 2079 -500 2113 -493
rect 2153 493 2187 500
rect 2153 -493 2160 493
rect 2176 -493 2187 493
rect 2153 -500 2187 -493
rect 2237 493 2271 500
rect 2237 -493 2248 493
rect 2264 -493 2271 493
rect 2237 -500 2271 -493
rect 2311 493 2345 500
rect 2311 -493 2318 493
rect 2334 -493 2345 493
rect 2311 -500 2345 -493
rect 2395 493 2429 500
rect 2395 -493 2406 493
rect 2422 -493 2429 493
rect 2395 -500 2429 -493
rect 2469 493 2503 500
rect 2469 -493 2476 493
rect 2492 -493 2503 493
rect 2469 -500 2503 -493
rect 2553 493 2587 500
rect 2553 -493 2564 493
rect 2580 -493 2587 493
rect 2553 -500 2587 -493
rect 2627 493 2661 500
rect 2627 -493 2634 493
rect 2650 -493 2661 493
rect 2627 -500 2661 -493
rect 2711 493 2745 500
rect 2711 -493 2722 493
rect 2738 -493 2745 493
rect 2711 -500 2745 -493
rect 2785 493 2819 500
rect 2785 -493 2792 493
rect 2808 -493 2819 493
rect 2785 -500 2819 -493
rect 2869 493 2903 500
rect 2869 -493 2880 493
rect 2896 -493 2903 493
rect 2869 -500 2903 -493
rect 2943 493 2977 500
rect 2943 -493 2950 493
rect 2966 -493 2977 493
rect 2943 -500 2977 -493
rect 3027 493 3061 500
rect 3027 -493 3038 493
rect 3054 -493 3061 493
rect 3027 -500 3061 -493
<< hvpdiffc >>
rect -52 599 -36 1585
rect 36 599 52 1585
rect 106 599 122 1585
rect 194 599 210 1585
rect 264 599 280 1585
rect 352 599 368 1585
rect 422 599 438 1585
rect 510 599 526 1585
rect 580 599 596 1585
rect 668 599 684 1585
rect 738 599 754 1585
rect 826 599 842 1585
rect 896 599 912 1585
rect 984 599 1000 1585
rect 1054 599 1070 1585
rect 1142 599 1158 1585
rect 1212 599 1228 1585
rect 1300 599 1316 1585
rect 1370 599 1386 1585
rect 1458 599 1474 1585
rect 1528 599 1544 1585
rect 1616 599 1632 1585
rect 1686 599 1702 1585
rect 1774 599 1790 1585
rect 1844 599 1860 1585
rect 1932 599 1948 1585
rect 2002 599 2018 1585
rect 2090 599 2106 1585
rect 2160 599 2176 1585
rect 2248 599 2264 1585
rect 2318 599 2334 1585
rect 2406 599 2422 1585
rect 2476 599 2492 1585
rect 2564 599 2580 1585
rect 2634 599 2650 1585
rect 2722 599 2738 1585
rect 2792 599 2808 1585
rect 2880 599 2896 1585
rect 2950 599 2966 1585
rect 3038 599 3054 1585
rect -52 -493 -36 493
rect 36 -493 52 493
rect 106 -493 122 493
rect 194 -493 210 493
rect 264 -493 280 493
rect 352 -493 368 493
rect 422 -493 438 493
rect 510 -493 526 493
rect 580 -493 596 493
rect 668 -493 684 493
rect 738 -493 754 493
rect 826 -493 842 493
rect 896 -493 912 493
rect 984 -493 1000 493
rect 1054 -493 1070 493
rect 1142 -493 1158 493
rect 1212 -493 1228 493
rect 1300 -493 1316 493
rect 1370 -493 1386 493
rect 1458 -493 1474 493
rect 1528 -493 1544 493
rect 1616 -493 1632 493
rect 1686 -493 1702 493
rect 1774 -493 1790 493
rect 1844 -493 1860 493
rect 1932 -493 1948 493
rect 2002 -493 2018 493
rect 2090 -493 2106 493
rect 2160 -493 2176 493
rect 2248 -493 2264 493
rect 2318 -493 2334 493
rect 2406 -493 2422 493
rect 2476 -493 2492 493
rect 2564 -493 2580 493
rect 2634 -493 2650 493
rect 2722 -493 2738 493
rect 2792 -493 2808 493
rect 2880 -493 2896 493
rect 2950 -493 2966 493
rect 3038 -493 3054 493
<< nsubdiff >>
rect -143 1674 3145 1681
rect -143 1658 -106 1674
rect 3108 1658 3145 1674
rect -143 1651 3145 1658
rect -143 1644 -113 1651
rect -143 -552 -136 1644
rect -120 -552 -113 1644
rect 3115 1644 3145 1651
rect -143 -559 -113 -552
rect 3115 -552 3122 1644
rect 3138 -552 3145 1644
rect 3115 -559 3145 -552
rect -143 -566 3145 -559
rect -143 -582 -106 -566
rect 3108 -582 3145 -566
rect -143 -589 3145 -582
<< nsubdiffcont >>
rect -106 1658 3108 1674
rect -136 -552 -120 1644
rect 3122 -552 3138 1644
rect -106 -582 3108 -566
<< poly >>
rect -25 1622 25 1629
rect -25 1606 -18 1622
rect 18 1606 25 1622
rect -25 1592 25 1606
rect 133 1622 183 1629
rect 133 1606 140 1622
rect 176 1606 183 1622
rect 133 1592 183 1606
rect 291 1622 341 1629
rect 291 1606 298 1622
rect 334 1606 341 1622
rect 291 1592 341 1606
rect 449 1622 499 1629
rect 449 1606 456 1622
rect 492 1606 499 1622
rect 449 1592 499 1606
rect 607 1622 657 1629
rect 607 1606 614 1622
rect 650 1606 657 1622
rect 607 1592 657 1606
rect 765 1622 815 1629
rect 765 1606 772 1622
rect 808 1606 815 1622
rect 765 1592 815 1606
rect 923 1622 973 1629
rect 923 1606 930 1622
rect 966 1606 973 1622
rect 923 1592 973 1606
rect 1081 1622 1131 1629
rect 1081 1606 1088 1622
rect 1124 1606 1131 1622
rect 1081 1592 1131 1606
rect 1239 1622 1289 1629
rect 1239 1606 1246 1622
rect 1282 1606 1289 1622
rect 1239 1592 1289 1606
rect 1397 1622 1447 1629
rect 1397 1606 1404 1622
rect 1440 1606 1447 1622
rect 1397 1592 1447 1606
rect 1555 1622 1605 1629
rect 1555 1606 1562 1622
rect 1598 1606 1605 1622
rect 1555 1592 1605 1606
rect 1713 1622 1763 1629
rect 1713 1606 1720 1622
rect 1756 1606 1763 1622
rect 1713 1592 1763 1606
rect 1871 1622 1921 1629
rect 1871 1606 1878 1622
rect 1914 1606 1921 1622
rect 1871 1592 1921 1606
rect 2029 1622 2079 1629
rect 2029 1606 2036 1622
rect 2072 1606 2079 1622
rect 2029 1592 2079 1606
rect 2187 1622 2237 1629
rect 2187 1606 2194 1622
rect 2230 1606 2237 1622
rect 2187 1592 2237 1606
rect 2345 1622 2395 1629
rect 2345 1606 2352 1622
rect 2388 1606 2395 1622
rect 2345 1592 2395 1606
rect 2503 1622 2553 1629
rect 2503 1606 2510 1622
rect 2546 1606 2553 1622
rect 2503 1592 2553 1606
rect 2661 1622 2711 1629
rect 2661 1606 2668 1622
rect 2704 1606 2711 1622
rect 2661 1592 2711 1606
rect 2819 1622 2869 1629
rect 2819 1606 2826 1622
rect 2862 1606 2869 1622
rect 2819 1592 2869 1606
rect 2977 1622 3027 1629
rect 2977 1606 2984 1622
rect 3020 1606 3027 1622
rect 2977 1592 3027 1606
rect -25 578 25 592
rect -25 562 -18 578
rect 18 562 25 578
rect -25 555 25 562
rect 133 578 183 592
rect 133 562 140 578
rect 176 562 183 578
rect 133 555 183 562
rect 291 578 341 592
rect 291 562 298 578
rect 334 562 341 578
rect 291 555 341 562
rect 449 578 499 592
rect 449 562 456 578
rect 492 562 499 578
rect 449 555 499 562
rect 607 578 657 592
rect 607 562 614 578
rect 650 562 657 578
rect 607 555 657 562
rect 765 578 815 592
rect 765 562 772 578
rect 808 562 815 578
rect 765 555 815 562
rect 923 578 973 592
rect 923 562 930 578
rect 966 562 973 578
rect 923 555 973 562
rect 1081 578 1131 592
rect 1081 562 1088 578
rect 1124 562 1131 578
rect 1081 555 1131 562
rect 1239 578 1289 592
rect 1239 562 1246 578
rect 1282 562 1289 578
rect 1239 555 1289 562
rect 1397 578 1447 592
rect 1397 562 1404 578
rect 1440 562 1447 578
rect 1397 555 1447 562
rect 1555 578 1605 592
rect 1555 562 1562 578
rect 1598 562 1605 578
rect 1555 555 1605 562
rect 1713 578 1763 592
rect 1713 562 1720 578
rect 1756 562 1763 578
rect 1713 555 1763 562
rect 1871 578 1921 592
rect 1871 562 1878 578
rect 1914 562 1921 578
rect 1871 555 1921 562
rect 2029 578 2079 592
rect 2029 562 2036 578
rect 2072 562 2079 578
rect 2029 555 2079 562
rect 2187 578 2237 592
rect 2187 562 2194 578
rect 2230 562 2237 578
rect 2187 555 2237 562
rect 2345 578 2395 592
rect 2345 562 2352 578
rect 2388 562 2395 578
rect 2345 555 2395 562
rect 2503 578 2553 592
rect 2503 562 2510 578
rect 2546 562 2553 578
rect 2503 555 2553 562
rect 2661 578 2711 592
rect 2661 562 2668 578
rect 2704 562 2711 578
rect 2661 555 2711 562
rect 2819 578 2869 592
rect 2819 562 2826 578
rect 2862 562 2869 578
rect 2819 555 2869 562
rect 2977 578 3027 592
rect 2977 562 2984 578
rect 3020 562 3027 578
rect 2977 555 3027 562
rect -25 530 25 537
rect -25 514 -18 530
rect 18 514 25 530
rect -25 500 25 514
rect 133 530 183 537
rect 133 514 140 530
rect 176 514 183 530
rect 133 500 183 514
rect 291 530 341 537
rect 291 514 298 530
rect 334 514 341 530
rect 291 500 341 514
rect 449 530 499 537
rect 449 514 456 530
rect 492 514 499 530
rect 449 500 499 514
rect 607 530 657 537
rect 607 514 614 530
rect 650 514 657 530
rect 607 500 657 514
rect 765 530 815 537
rect 765 514 772 530
rect 808 514 815 530
rect 765 500 815 514
rect 923 530 973 537
rect 923 514 930 530
rect 966 514 973 530
rect 923 500 973 514
rect 1081 530 1131 537
rect 1081 514 1088 530
rect 1124 514 1131 530
rect 1081 500 1131 514
rect 1239 530 1289 537
rect 1239 514 1246 530
rect 1282 514 1289 530
rect 1239 500 1289 514
rect 1397 530 1447 537
rect 1397 514 1404 530
rect 1440 514 1447 530
rect 1397 500 1447 514
rect 1555 530 1605 537
rect 1555 514 1562 530
rect 1598 514 1605 530
rect 1555 500 1605 514
rect 1713 530 1763 537
rect 1713 514 1720 530
rect 1756 514 1763 530
rect 1713 500 1763 514
rect 1871 530 1921 537
rect 1871 514 1878 530
rect 1914 514 1921 530
rect 1871 500 1921 514
rect 2029 530 2079 537
rect 2029 514 2036 530
rect 2072 514 2079 530
rect 2029 500 2079 514
rect 2187 530 2237 537
rect 2187 514 2194 530
rect 2230 514 2237 530
rect 2187 500 2237 514
rect 2345 530 2395 537
rect 2345 514 2352 530
rect 2388 514 2395 530
rect 2345 500 2395 514
rect 2503 530 2553 537
rect 2503 514 2510 530
rect 2546 514 2553 530
rect 2503 500 2553 514
rect 2661 530 2711 537
rect 2661 514 2668 530
rect 2704 514 2711 530
rect 2661 500 2711 514
rect 2819 530 2869 537
rect 2819 514 2826 530
rect 2862 514 2869 530
rect 2819 500 2869 514
rect 2977 530 3027 537
rect 2977 514 2984 530
rect 3020 514 3027 530
rect 2977 500 3027 514
rect -25 -514 25 -500
rect -25 -530 -18 -514
rect 18 -530 25 -514
rect -25 -537 25 -530
rect 133 -514 183 -500
rect 133 -530 140 -514
rect 176 -530 183 -514
rect 133 -537 183 -530
rect 291 -514 341 -500
rect 291 -530 298 -514
rect 334 -530 341 -514
rect 291 -537 341 -530
rect 449 -514 499 -500
rect 449 -530 456 -514
rect 492 -530 499 -514
rect 449 -537 499 -530
rect 607 -514 657 -500
rect 607 -530 614 -514
rect 650 -530 657 -514
rect 607 -537 657 -530
rect 765 -514 815 -500
rect 765 -530 772 -514
rect 808 -530 815 -514
rect 765 -537 815 -530
rect 923 -514 973 -500
rect 923 -530 930 -514
rect 966 -530 973 -514
rect 923 -537 973 -530
rect 1081 -514 1131 -500
rect 1081 -530 1088 -514
rect 1124 -530 1131 -514
rect 1081 -537 1131 -530
rect 1239 -514 1289 -500
rect 1239 -530 1246 -514
rect 1282 -530 1289 -514
rect 1239 -537 1289 -530
rect 1397 -514 1447 -500
rect 1397 -530 1404 -514
rect 1440 -530 1447 -514
rect 1397 -537 1447 -530
rect 1555 -514 1605 -500
rect 1555 -530 1562 -514
rect 1598 -530 1605 -514
rect 1555 -537 1605 -530
rect 1713 -514 1763 -500
rect 1713 -530 1720 -514
rect 1756 -530 1763 -514
rect 1713 -537 1763 -530
rect 1871 -514 1921 -500
rect 1871 -530 1878 -514
rect 1914 -530 1921 -514
rect 1871 -537 1921 -530
rect 2029 -514 2079 -500
rect 2029 -530 2036 -514
rect 2072 -530 2079 -514
rect 2029 -537 2079 -530
rect 2187 -514 2237 -500
rect 2187 -530 2194 -514
rect 2230 -530 2237 -514
rect 2187 -537 2237 -530
rect 2345 -514 2395 -500
rect 2345 -530 2352 -514
rect 2388 -530 2395 -514
rect 2345 -537 2395 -530
rect 2503 -514 2553 -500
rect 2503 -530 2510 -514
rect 2546 -530 2553 -514
rect 2503 -537 2553 -530
rect 2661 -514 2711 -500
rect 2661 -530 2668 -514
rect 2704 -530 2711 -514
rect 2661 -537 2711 -530
rect 2819 -514 2869 -500
rect 2819 -530 2826 -514
rect 2862 -530 2869 -514
rect 2819 -537 2869 -530
rect 2977 -514 3027 -500
rect 2977 -530 2984 -514
rect 3020 -530 3027 -514
rect 2977 -537 3027 -530
<< polycont >>
rect -18 1606 18 1622
rect 140 1606 176 1622
rect 298 1606 334 1622
rect 456 1606 492 1622
rect 614 1606 650 1622
rect 772 1606 808 1622
rect 930 1606 966 1622
rect 1088 1606 1124 1622
rect 1246 1606 1282 1622
rect 1404 1606 1440 1622
rect 1562 1606 1598 1622
rect 1720 1606 1756 1622
rect 1878 1606 1914 1622
rect 2036 1606 2072 1622
rect 2194 1606 2230 1622
rect 2352 1606 2388 1622
rect 2510 1606 2546 1622
rect 2668 1606 2704 1622
rect 2826 1606 2862 1622
rect 2984 1606 3020 1622
rect -18 562 18 578
rect 140 562 176 578
rect 298 562 334 578
rect 456 562 492 578
rect 614 562 650 578
rect 772 562 808 578
rect 930 562 966 578
rect 1088 562 1124 578
rect 1246 562 1282 578
rect 1404 562 1440 578
rect 1562 562 1598 578
rect 1720 562 1756 578
rect 1878 562 1914 578
rect 2036 562 2072 578
rect 2194 562 2230 578
rect 2352 562 2388 578
rect 2510 562 2546 578
rect 2668 562 2704 578
rect 2826 562 2862 578
rect 2984 562 3020 578
rect -18 514 18 530
rect 140 514 176 530
rect 298 514 334 530
rect 456 514 492 530
rect 614 514 650 530
rect 772 514 808 530
rect 930 514 966 530
rect 1088 514 1124 530
rect 1246 514 1282 530
rect 1404 514 1440 530
rect 1562 514 1598 530
rect 1720 514 1756 530
rect 1878 514 1914 530
rect 2036 514 2072 530
rect 2194 514 2230 530
rect 2352 514 2388 530
rect 2510 514 2546 530
rect 2668 514 2704 530
rect 2826 514 2862 530
rect 2984 514 3020 530
rect -18 -530 18 -514
rect 140 -530 176 -514
rect 298 -530 334 -514
rect 456 -530 492 -514
rect 614 -530 650 -514
rect 772 -530 808 -514
rect 930 -530 966 -514
rect 1088 -530 1124 -514
rect 1246 -530 1282 -514
rect 1404 -530 1440 -514
rect 1562 -530 1598 -514
rect 1720 -530 1756 -514
rect 1878 -530 1914 -514
rect 2036 -530 2072 -514
rect 2194 -530 2230 -514
rect 2352 -530 2388 -514
rect 2510 -530 2546 -514
rect 2668 -530 2704 -514
rect 2826 -530 2862 -514
rect 2984 -530 3020 -514
<< metal1 >>
rect -141 1674 3143 1679
rect -141 1658 -106 1674
rect 3108 1658 3143 1674
rect -141 1653 3143 1658
rect -141 1644 -115 1653
rect -141 -552 -136 1644
rect -120 -552 -115 1644
rect 3117 1644 3143 1653
rect -141 -561 -115 -552
rect 3117 -552 3122 1644
rect 3138 -552 3143 1644
rect 3117 -561 3143 -552
rect -141 -566 3143 -561
rect -141 -582 -106 -566
rect 3108 -582 3143 -566
rect -141 -587 3143 -582
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 10 l 0.5 nf 1 nx 20 dx 0.4 ny 2 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
