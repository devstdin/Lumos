magic
tech ihp-sg13g2
timestamp 1748519341
<< error_p >>
rect -93 530 -88 535
rect 88 530 93 535
rect 255 530 260 535
rect 436 530 441 535
rect 603 530 608 535
rect 784 530 789 535
rect 951 530 956 535
rect 1132 530 1137 535
rect -98 525 -93 530
rect 93 525 98 530
rect 250 525 255 530
rect 441 525 446 530
rect 598 525 603 530
rect 789 525 794 530
rect 946 525 951 530
rect 1137 525 1142 530
rect -98 514 -93 519
rect 93 514 98 519
rect 250 514 255 519
rect 441 514 446 519
rect 598 514 603 519
rect 789 514 794 519
rect 946 514 951 519
rect 1137 514 1142 519
rect -93 509 -88 514
rect 88 509 93 514
rect 255 509 260 514
rect 436 509 441 514
rect 603 509 608 514
rect 784 509 789 514
rect 951 509 956 514
rect 1132 509 1137 514
rect -127 493 -122 498
rect -116 493 -111 498
rect 111 493 116 498
rect 122 493 127 498
rect 221 493 226 498
rect 232 493 237 498
rect 459 493 464 498
rect 470 493 475 498
rect 569 493 574 498
rect 580 493 585 498
rect 807 493 812 498
rect 818 493 823 498
rect 917 493 922 498
rect 928 493 933 498
rect 1155 493 1160 498
rect 1166 493 1171 498
rect -132 488 -127 493
rect -111 488 -106 493
rect 106 488 111 493
rect 127 488 132 493
rect 216 488 221 493
rect 237 488 242 493
rect 454 488 459 493
rect 475 488 480 493
rect 564 488 569 493
rect 585 488 590 493
rect 802 488 807 493
rect 823 488 828 493
rect 912 488 917 493
rect 933 488 938 493
rect 1150 488 1155 493
rect 1171 488 1176 493
rect -132 -493 -127 -488
rect -111 -493 -106 -488
rect 106 -493 111 -488
rect 127 -493 132 -488
rect 216 -493 221 -488
rect 237 -493 242 -488
rect 454 -493 459 -488
rect 475 -493 480 -488
rect 564 -493 569 -488
rect 585 -493 590 -488
rect 802 -493 807 -488
rect 823 -493 828 -488
rect 912 -493 917 -488
rect 933 -493 938 -488
rect 1150 -493 1155 -488
rect 1171 -493 1176 -488
rect -127 -498 -122 -493
rect -116 -498 -111 -493
rect 111 -498 116 -493
rect 122 -498 127 -493
rect 221 -498 226 -493
rect 232 -498 237 -493
rect 459 -498 464 -493
rect 470 -498 475 -493
rect 569 -498 574 -493
rect 580 -498 585 -493
rect 807 -498 812 -493
rect 818 -498 823 -493
rect 917 -498 922 -493
rect 928 -498 933 -493
rect 1155 -498 1160 -493
rect 1166 -498 1171 -493
rect -93 -514 -88 -509
rect 88 -514 93 -509
rect 255 -514 260 -509
rect 436 -514 441 -509
rect 603 -514 608 -509
rect 784 -514 789 -509
rect 951 -514 956 -509
rect 1132 -514 1137 -509
rect -98 -519 -93 -514
rect 93 -519 98 -514
rect 250 -519 255 -514
rect 441 -519 446 -514
rect 598 -519 603 -514
rect 789 -519 794 -514
rect 946 -519 951 -514
rect 1137 -519 1142 -514
rect -98 -530 -93 -525
rect 93 -530 98 -525
rect 250 -530 255 -525
rect 441 -530 446 -525
rect 598 -530 603 -525
rect 789 -530 794 -525
rect 946 -530 951 -525
rect 1137 -530 1142 -525
rect -93 -535 -88 -530
rect 88 -535 93 -530
rect 255 -535 260 -530
rect 436 -535 441 -530
rect 603 -535 608 -530
rect 784 -535 789 -530
rect 951 -535 956 -530
rect 1132 -535 1137 -530
<< hvnmos >>
rect -100 -500 100 500
rect 248 -500 448 500
rect 596 -500 796 500
rect 944 -500 1144 500
<< hvndiff >>
rect -134 493 -100 500
rect -134 -493 -127 493
rect -111 -493 -100 493
rect -134 -500 -100 -493
rect 100 493 134 500
rect 100 -493 111 493
rect 127 -493 134 493
rect 100 -500 134 -493
rect 214 493 248 500
rect 214 -493 221 493
rect 237 -493 248 493
rect 214 -500 248 -493
rect 448 493 482 500
rect 448 -493 459 493
rect 475 -493 482 493
rect 448 -500 482 -493
rect 562 493 596 500
rect 562 -493 569 493
rect 585 -493 596 493
rect 562 -500 596 -493
rect 796 493 830 500
rect 796 -493 807 493
rect 823 -493 830 493
rect 796 -500 830 -493
rect 910 493 944 500
rect 910 -493 917 493
rect 933 -493 944 493
rect 910 -500 944 -493
rect 1144 493 1178 500
rect 1144 -493 1155 493
rect 1171 -493 1178 493
rect 1144 -500 1178 -493
<< hvndiffc >>
rect -127 -493 -111 493
rect 111 -493 127 493
rect 221 -493 237 493
rect 459 -493 475 493
rect 569 -493 585 493
rect 807 -493 823 493
rect 917 -493 933 493
rect 1155 -493 1171 493
<< psubdiff >>
rect -326 626 1178 633
rect -326 610 -289 626
rect 1171 610 1178 626
rect -326 603 1178 610
rect -326 596 -296 603
rect -326 -596 -319 596
rect -303 -596 -296 596
rect -326 -603 -296 -596
rect -326 -610 1178 -603
rect -326 -626 -289 -610
rect 1171 -626 1178 -610
rect -326 -633 1178 -626
<< psubdiffcont >>
rect -289 610 1171 626
rect -319 -596 -303 596
rect -289 -626 1171 -610
<< poly >>
rect -100 530 100 537
rect -100 514 -93 530
rect 93 514 100 530
rect -100 500 100 514
rect 248 530 448 537
rect 248 514 255 530
rect 441 514 448 530
rect 248 500 448 514
rect 596 530 796 537
rect 596 514 603 530
rect 789 514 796 530
rect 596 500 796 514
rect 944 530 1144 537
rect 944 514 951 530
rect 1137 514 1144 530
rect 944 500 1144 514
rect -100 -514 100 -500
rect -100 -530 -93 -514
rect 93 -530 100 -514
rect -100 -537 100 -530
rect 248 -514 448 -500
rect 248 -530 255 -514
rect 441 -530 448 -514
rect 248 -537 448 -530
rect 596 -514 796 -500
rect 596 -530 603 -514
rect 789 -530 796 -514
rect 596 -537 796 -530
rect 944 -514 1144 -500
rect 944 -530 951 -514
rect 1137 -530 1144 -514
rect 944 -537 1144 -530
<< polycont >>
rect -93 514 93 530
rect 255 514 441 530
rect 603 514 789 530
rect 951 514 1137 530
rect -93 -530 93 -514
rect 255 -530 441 -514
rect 603 -530 789 -514
rect 951 -530 1137 -514
<< metal1 >>
rect -324 626 1176 631
rect -324 610 -289 626
rect 1171 610 1176 626
rect -324 605 1176 610
rect -324 596 -298 605
rect -324 -596 -319 596
rect -303 -596 -298 596
rect -324 -605 -298 -596
rect -324 -610 1176 -605
rect -324 -626 -289 -610
rect 1171 -626 1176 -610
rect -324 -631 1176 -626
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 10 l 2 nf 1 nx 4 dx 0.8 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 3 glc 1 grc 0 gtc 1 gbc 1
<< end >>
