magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2026 -2026 18026 5878
<< nwell >>
rect 236 236 15764 3616
<< pwell >>
rect -26 3758 16026 3878
rect -26 94 94 3758
rect 15906 94 16026 3758
rect -26 -26 16026 94
<< hvpmos >>
rect 6856 1970 6976 3302
rect 7212 1970 7332 3302
rect 7460 1970 7580 3302
rect 7816 1970 7936 3302
rect 8064 1970 8184 3302
rect 8420 1970 8540 3302
rect 8668 1970 8788 3302
rect 9024 1970 9144 3302
rect 6856 550 6976 1882
rect 7212 550 7332 1882
rect 7460 550 7580 1882
rect 7816 550 7936 1882
rect 8064 550 8184 1882
rect 8420 550 8540 1882
rect 8668 550 8788 1882
rect 9024 550 9144 1882
<< hvpdiff >>
rect 6762 3264 6856 3302
rect 6762 3232 6776 3264
rect 6808 3232 6856 3264
rect 6762 3196 6856 3232
rect 6762 3164 6776 3196
rect 6808 3164 6856 3196
rect 6762 3128 6856 3164
rect 6762 3096 6776 3128
rect 6808 3096 6856 3128
rect 6762 3060 6856 3096
rect 6762 3028 6776 3060
rect 6808 3028 6856 3060
rect 6762 2992 6856 3028
rect 6762 2960 6776 2992
rect 6808 2960 6856 2992
rect 6762 2924 6856 2960
rect 6762 2892 6776 2924
rect 6808 2892 6856 2924
rect 6762 2856 6856 2892
rect 6762 2824 6776 2856
rect 6808 2824 6856 2856
rect 6762 2788 6856 2824
rect 6762 2756 6776 2788
rect 6808 2756 6856 2788
rect 6762 2720 6856 2756
rect 6762 2688 6776 2720
rect 6808 2688 6856 2720
rect 6762 2652 6856 2688
rect 6762 2620 6776 2652
rect 6808 2620 6856 2652
rect 6762 2584 6856 2620
rect 6762 2552 6776 2584
rect 6808 2552 6856 2584
rect 6762 2516 6856 2552
rect 6762 2484 6776 2516
rect 6808 2484 6856 2516
rect 6762 2448 6856 2484
rect 6762 2416 6776 2448
rect 6808 2416 6856 2448
rect 6762 2380 6856 2416
rect 6762 2348 6776 2380
rect 6808 2348 6856 2380
rect 6762 2312 6856 2348
rect 6762 2280 6776 2312
rect 6808 2280 6856 2312
rect 6762 2244 6856 2280
rect 6762 2212 6776 2244
rect 6808 2212 6856 2244
rect 6762 2176 6856 2212
rect 6762 2144 6776 2176
rect 6808 2144 6856 2176
rect 6762 2108 6856 2144
rect 6762 2076 6776 2108
rect 6808 2076 6856 2108
rect 6762 2040 6856 2076
rect 6762 2008 6776 2040
rect 6808 2008 6856 2040
rect 6762 1970 6856 2008
rect 6976 3264 7212 3302
rect 6976 3232 7078 3264
rect 7110 3232 7212 3264
rect 6976 3196 7212 3232
rect 6976 3164 7078 3196
rect 7110 3164 7212 3196
rect 6976 3128 7212 3164
rect 6976 3096 7078 3128
rect 7110 3096 7212 3128
rect 6976 3060 7212 3096
rect 6976 3028 7078 3060
rect 7110 3028 7212 3060
rect 6976 2992 7212 3028
rect 6976 2960 7078 2992
rect 7110 2960 7212 2992
rect 6976 2924 7212 2960
rect 6976 2892 7078 2924
rect 7110 2892 7212 2924
rect 6976 2856 7212 2892
rect 6976 2824 7078 2856
rect 7110 2824 7212 2856
rect 6976 2788 7212 2824
rect 6976 2756 7078 2788
rect 7110 2756 7212 2788
rect 6976 2720 7212 2756
rect 6976 2688 7078 2720
rect 7110 2688 7212 2720
rect 6976 2652 7212 2688
rect 6976 2620 7078 2652
rect 7110 2620 7212 2652
rect 6976 2584 7212 2620
rect 6976 2552 7078 2584
rect 7110 2552 7212 2584
rect 6976 2516 7212 2552
rect 6976 2484 7078 2516
rect 7110 2484 7212 2516
rect 6976 2448 7212 2484
rect 6976 2416 7078 2448
rect 7110 2416 7212 2448
rect 6976 2380 7212 2416
rect 6976 2348 7078 2380
rect 7110 2348 7212 2380
rect 6976 2312 7212 2348
rect 6976 2280 7078 2312
rect 7110 2280 7212 2312
rect 6976 2244 7212 2280
rect 6976 2212 7078 2244
rect 7110 2212 7212 2244
rect 6976 2176 7212 2212
rect 6976 2144 7078 2176
rect 7110 2144 7212 2176
rect 6976 2108 7212 2144
rect 6976 2076 7078 2108
rect 7110 2076 7212 2108
rect 6976 2040 7212 2076
rect 6976 2008 7078 2040
rect 7110 2008 7212 2040
rect 6976 1970 7212 2008
rect 7332 3264 7460 3302
rect 7332 3232 7380 3264
rect 7412 3232 7460 3264
rect 7332 3196 7460 3232
rect 7332 3164 7380 3196
rect 7412 3164 7460 3196
rect 7332 3128 7460 3164
rect 7332 3096 7380 3128
rect 7412 3096 7460 3128
rect 7332 3060 7460 3096
rect 7332 3028 7380 3060
rect 7412 3028 7460 3060
rect 7332 2992 7460 3028
rect 7332 2960 7380 2992
rect 7412 2960 7460 2992
rect 7332 2924 7460 2960
rect 7332 2892 7380 2924
rect 7412 2892 7460 2924
rect 7332 2856 7460 2892
rect 7332 2824 7380 2856
rect 7412 2824 7460 2856
rect 7332 2788 7460 2824
rect 7332 2756 7380 2788
rect 7412 2756 7460 2788
rect 7332 2720 7460 2756
rect 7332 2688 7380 2720
rect 7412 2688 7460 2720
rect 7332 2652 7460 2688
rect 7332 2620 7380 2652
rect 7412 2620 7460 2652
rect 7332 2584 7460 2620
rect 7332 2552 7380 2584
rect 7412 2552 7460 2584
rect 7332 2516 7460 2552
rect 7332 2484 7380 2516
rect 7412 2484 7460 2516
rect 7332 2448 7460 2484
rect 7332 2416 7380 2448
rect 7412 2416 7460 2448
rect 7332 2380 7460 2416
rect 7332 2348 7380 2380
rect 7412 2348 7460 2380
rect 7332 2312 7460 2348
rect 7332 2280 7380 2312
rect 7412 2280 7460 2312
rect 7332 2244 7460 2280
rect 7332 2212 7380 2244
rect 7412 2212 7460 2244
rect 7332 2176 7460 2212
rect 7332 2144 7380 2176
rect 7412 2144 7460 2176
rect 7332 2108 7460 2144
rect 7332 2076 7380 2108
rect 7412 2076 7460 2108
rect 7332 2040 7460 2076
rect 7332 2008 7380 2040
rect 7412 2008 7460 2040
rect 7332 1970 7460 2008
rect 7580 3264 7816 3302
rect 7580 3232 7682 3264
rect 7714 3232 7816 3264
rect 7580 3196 7816 3232
rect 7580 3164 7682 3196
rect 7714 3164 7816 3196
rect 7580 3128 7816 3164
rect 7580 3096 7682 3128
rect 7714 3096 7816 3128
rect 7580 3060 7816 3096
rect 7580 3028 7682 3060
rect 7714 3028 7816 3060
rect 7580 2992 7816 3028
rect 7580 2960 7682 2992
rect 7714 2960 7816 2992
rect 7580 2924 7816 2960
rect 7580 2892 7682 2924
rect 7714 2892 7816 2924
rect 7580 2856 7816 2892
rect 7580 2824 7682 2856
rect 7714 2824 7816 2856
rect 7580 2788 7816 2824
rect 7580 2756 7682 2788
rect 7714 2756 7816 2788
rect 7580 2720 7816 2756
rect 7580 2688 7682 2720
rect 7714 2688 7816 2720
rect 7580 2652 7816 2688
rect 7580 2620 7682 2652
rect 7714 2620 7816 2652
rect 7580 2584 7816 2620
rect 7580 2552 7682 2584
rect 7714 2552 7816 2584
rect 7580 2516 7816 2552
rect 7580 2484 7682 2516
rect 7714 2484 7816 2516
rect 7580 2448 7816 2484
rect 7580 2416 7682 2448
rect 7714 2416 7816 2448
rect 7580 2380 7816 2416
rect 7580 2348 7682 2380
rect 7714 2348 7816 2380
rect 7580 2312 7816 2348
rect 7580 2280 7682 2312
rect 7714 2280 7816 2312
rect 7580 2244 7816 2280
rect 7580 2212 7682 2244
rect 7714 2212 7816 2244
rect 7580 2176 7816 2212
rect 7580 2144 7682 2176
rect 7714 2144 7816 2176
rect 7580 2108 7816 2144
rect 7580 2076 7682 2108
rect 7714 2076 7816 2108
rect 7580 2040 7816 2076
rect 7580 2008 7682 2040
rect 7714 2008 7816 2040
rect 7580 1970 7816 2008
rect 7936 3264 8064 3302
rect 7936 3232 7984 3264
rect 8016 3232 8064 3264
rect 7936 3196 8064 3232
rect 7936 3164 7984 3196
rect 8016 3164 8064 3196
rect 7936 3128 8064 3164
rect 7936 3096 7984 3128
rect 8016 3096 8064 3128
rect 7936 3060 8064 3096
rect 7936 3028 7984 3060
rect 8016 3028 8064 3060
rect 7936 2992 8064 3028
rect 7936 2960 7984 2992
rect 8016 2960 8064 2992
rect 7936 2924 8064 2960
rect 7936 2892 7984 2924
rect 8016 2892 8064 2924
rect 7936 2856 8064 2892
rect 7936 2824 7984 2856
rect 8016 2824 8064 2856
rect 7936 2788 8064 2824
rect 7936 2756 7984 2788
rect 8016 2756 8064 2788
rect 7936 2720 8064 2756
rect 7936 2688 7984 2720
rect 8016 2688 8064 2720
rect 7936 2652 8064 2688
rect 7936 2620 7984 2652
rect 8016 2620 8064 2652
rect 7936 2584 8064 2620
rect 7936 2552 7984 2584
rect 8016 2552 8064 2584
rect 7936 2516 8064 2552
rect 7936 2484 7984 2516
rect 8016 2484 8064 2516
rect 7936 2448 8064 2484
rect 7936 2416 7984 2448
rect 8016 2416 8064 2448
rect 7936 2380 8064 2416
rect 7936 2348 7984 2380
rect 8016 2348 8064 2380
rect 7936 2312 8064 2348
rect 7936 2280 7984 2312
rect 8016 2280 8064 2312
rect 7936 2244 8064 2280
rect 7936 2212 7984 2244
rect 8016 2212 8064 2244
rect 7936 2176 8064 2212
rect 7936 2144 7984 2176
rect 8016 2144 8064 2176
rect 7936 2108 8064 2144
rect 7936 2076 7984 2108
rect 8016 2076 8064 2108
rect 7936 2040 8064 2076
rect 7936 2008 7984 2040
rect 8016 2008 8064 2040
rect 7936 1970 8064 2008
rect 8184 3264 8420 3302
rect 8184 3232 8286 3264
rect 8318 3232 8420 3264
rect 8184 3196 8420 3232
rect 8184 3164 8286 3196
rect 8318 3164 8420 3196
rect 8184 3128 8420 3164
rect 8184 3096 8286 3128
rect 8318 3096 8420 3128
rect 8184 3060 8420 3096
rect 8184 3028 8286 3060
rect 8318 3028 8420 3060
rect 8184 2992 8420 3028
rect 8184 2960 8286 2992
rect 8318 2960 8420 2992
rect 8184 2924 8420 2960
rect 8184 2892 8286 2924
rect 8318 2892 8420 2924
rect 8184 2856 8420 2892
rect 8184 2824 8286 2856
rect 8318 2824 8420 2856
rect 8184 2788 8420 2824
rect 8184 2756 8286 2788
rect 8318 2756 8420 2788
rect 8184 2720 8420 2756
rect 8184 2688 8286 2720
rect 8318 2688 8420 2720
rect 8184 2652 8420 2688
rect 8184 2620 8286 2652
rect 8318 2620 8420 2652
rect 8184 2584 8420 2620
rect 8184 2552 8286 2584
rect 8318 2552 8420 2584
rect 8184 2516 8420 2552
rect 8184 2484 8286 2516
rect 8318 2484 8420 2516
rect 8184 2448 8420 2484
rect 8184 2416 8286 2448
rect 8318 2416 8420 2448
rect 8184 2380 8420 2416
rect 8184 2348 8286 2380
rect 8318 2348 8420 2380
rect 8184 2312 8420 2348
rect 8184 2280 8286 2312
rect 8318 2280 8420 2312
rect 8184 2244 8420 2280
rect 8184 2212 8286 2244
rect 8318 2212 8420 2244
rect 8184 2176 8420 2212
rect 8184 2144 8286 2176
rect 8318 2144 8420 2176
rect 8184 2108 8420 2144
rect 8184 2076 8286 2108
rect 8318 2076 8420 2108
rect 8184 2040 8420 2076
rect 8184 2008 8286 2040
rect 8318 2008 8420 2040
rect 8184 1970 8420 2008
rect 8540 3264 8668 3302
rect 8540 3232 8588 3264
rect 8620 3232 8668 3264
rect 8540 3196 8668 3232
rect 8540 3164 8588 3196
rect 8620 3164 8668 3196
rect 8540 3128 8668 3164
rect 8540 3096 8588 3128
rect 8620 3096 8668 3128
rect 8540 3060 8668 3096
rect 8540 3028 8588 3060
rect 8620 3028 8668 3060
rect 8540 2992 8668 3028
rect 8540 2960 8588 2992
rect 8620 2960 8668 2992
rect 8540 2924 8668 2960
rect 8540 2892 8588 2924
rect 8620 2892 8668 2924
rect 8540 2856 8668 2892
rect 8540 2824 8588 2856
rect 8620 2824 8668 2856
rect 8540 2788 8668 2824
rect 8540 2756 8588 2788
rect 8620 2756 8668 2788
rect 8540 2720 8668 2756
rect 8540 2688 8588 2720
rect 8620 2688 8668 2720
rect 8540 2652 8668 2688
rect 8540 2620 8588 2652
rect 8620 2620 8668 2652
rect 8540 2584 8668 2620
rect 8540 2552 8588 2584
rect 8620 2552 8668 2584
rect 8540 2516 8668 2552
rect 8540 2484 8588 2516
rect 8620 2484 8668 2516
rect 8540 2448 8668 2484
rect 8540 2416 8588 2448
rect 8620 2416 8668 2448
rect 8540 2380 8668 2416
rect 8540 2348 8588 2380
rect 8620 2348 8668 2380
rect 8540 2312 8668 2348
rect 8540 2280 8588 2312
rect 8620 2280 8668 2312
rect 8540 2244 8668 2280
rect 8540 2212 8588 2244
rect 8620 2212 8668 2244
rect 8540 2176 8668 2212
rect 8540 2144 8588 2176
rect 8620 2144 8668 2176
rect 8540 2108 8668 2144
rect 8540 2076 8588 2108
rect 8620 2076 8668 2108
rect 8540 2040 8668 2076
rect 8540 2008 8588 2040
rect 8620 2008 8668 2040
rect 8540 1970 8668 2008
rect 8788 3264 9024 3302
rect 8788 3232 8890 3264
rect 8922 3232 9024 3264
rect 8788 3196 9024 3232
rect 8788 3164 8890 3196
rect 8922 3164 9024 3196
rect 8788 3128 9024 3164
rect 8788 3096 8890 3128
rect 8922 3096 9024 3128
rect 8788 3060 9024 3096
rect 8788 3028 8890 3060
rect 8922 3028 9024 3060
rect 8788 2992 9024 3028
rect 8788 2960 8890 2992
rect 8922 2960 9024 2992
rect 8788 2924 9024 2960
rect 8788 2892 8890 2924
rect 8922 2892 9024 2924
rect 8788 2856 9024 2892
rect 8788 2824 8890 2856
rect 8922 2824 9024 2856
rect 8788 2788 9024 2824
rect 8788 2756 8890 2788
rect 8922 2756 9024 2788
rect 8788 2720 9024 2756
rect 8788 2688 8890 2720
rect 8922 2688 9024 2720
rect 8788 2652 9024 2688
rect 8788 2620 8890 2652
rect 8922 2620 9024 2652
rect 8788 2584 9024 2620
rect 8788 2552 8890 2584
rect 8922 2552 9024 2584
rect 8788 2516 9024 2552
rect 8788 2484 8890 2516
rect 8922 2484 9024 2516
rect 8788 2448 9024 2484
rect 8788 2416 8890 2448
rect 8922 2416 9024 2448
rect 8788 2380 9024 2416
rect 8788 2348 8890 2380
rect 8922 2348 9024 2380
rect 8788 2312 9024 2348
rect 8788 2280 8890 2312
rect 8922 2280 9024 2312
rect 8788 2244 9024 2280
rect 8788 2212 8890 2244
rect 8922 2212 9024 2244
rect 8788 2176 9024 2212
rect 8788 2144 8890 2176
rect 8922 2144 9024 2176
rect 8788 2108 9024 2144
rect 8788 2076 8890 2108
rect 8922 2076 9024 2108
rect 8788 2040 9024 2076
rect 8788 2008 8890 2040
rect 8922 2008 9024 2040
rect 8788 1970 9024 2008
rect 9144 3264 9238 3302
rect 9144 3232 9192 3264
rect 9224 3232 9238 3264
rect 9144 3196 9238 3232
rect 9144 3164 9192 3196
rect 9224 3164 9238 3196
rect 9144 3128 9238 3164
rect 9144 3096 9192 3128
rect 9224 3096 9238 3128
rect 9144 3060 9238 3096
rect 9144 3028 9192 3060
rect 9224 3028 9238 3060
rect 9144 2992 9238 3028
rect 9144 2960 9192 2992
rect 9224 2960 9238 2992
rect 9144 2924 9238 2960
rect 9144 2892 9192 2924
rect 9224 2892 9238 2924
rect 9144 2856 9238 2892
rect 9144 2824 9192 2856
rect 9224 2824 9238 2856
rect 9144 2788 9238 2824
rect 9144 2756 9192 2788
rect 9224 2756 9238 2788
rect 9144 2720 9238 2756
rect 9144 2688 9192 2720
rect 9224 2688 9238 2720
rect 9144 2652 9238 2688
rect 9144 2620 9192 2652
rect 9224 2620 9238 2652
rect 9144 2584 9238 2620
rect 9144 2552 9192 2584
rect 9224 2552 9238 2584
rect 9144 2516 9238 2552
rect 9144 2484 9192 2516
rect 9224 2484 9238 2516
rect 9144 2448 9238 2484
rect 9144 2416 9192 2448
rect 9224 2416 9238 2448
rect 9144 2380 9238 2416
rect 9144 2348 9192 2380
rect 9224 2348 9238 2380
rect 9144 2312 9238 2348
rect 9144 2280 9192 2312
rect 9224 2280 9238 2312
rect 9144 2244 9238 2280
rect 9144 2212 9192 2244
rect 9224 2212 9238 2244
rect 9144 2176 9238 2212
rect 9144 2144 9192 2176
rect 9224 2144 9238 2176
rect 9144 2108 9238 2144
rect 9144 2076 9192 2108
rect 9224 2076 9238 2108
rect 9144 2040 9238 2076
rect 9144 2008 9192 2040
rect 9224 2008 9238 2040
rect 9144 1970 9238 2008
rect 6762 1844 6856 1882
rect 6762 1812 6776 1844
rect 6808 1812 6856 1844
rect 6762 1776 6856 1812
rect 6762 1744 6776 1776
rect 6808 1744 6856 1776
rect 6762 1708 6856 1744
rect 6762 1676 6776 1708
rect 6808 1676 6856 1708
rect 6762 1640 6856 1676
rect 6762 1608 6776 1640
rect 6808 1608 6856 1640
rect 6762 1572 6856 1608
rect 6762 1540 6776 1572
rect 6808 1540 6856 1572
rect 6762 1504 6856 1540
rect 6762 1472 6776 1504
rect 6808 1472 6856 1504
rect 6762 1436 6856 1472
rect 6762 1404 6776 1436
rect 6808 1404 6856 1436
rect 6762 1368 6856 1404
rect 6762 1336 6776 1368
rect 6808 1336 6856 1368
rect 6762 1300 6856 1336
rect 6762 1268 6776 1300
rect 6808 1268 6856 1300
rect 6762 1232 6856 1268
rect 6762 1200 6776 1232
rect 6808 1200 6856 1232
rect 6762 1164 6856 1200
rect 6762 1132 6776 1164
rect 6808 1132 6856 1164
rect 6762 1096 6856 1132
rect 6762 1064 6776 1096
rect 6808 1064 6856 1096
rect 6762 1028 6856 1064
rect 6762 996 6776 1028
rect 6808 996 6856 1028
rect 6762 960 6856 996
rect 6762 928 6776 960
rect 6808 928 6856 960
rect 6762 892 6856 928
rect 6762 860 6776 892
rect 6808 860 6856 892
rect 6762 824 6856 860
rect 6762 792 6776 824
rect 6808 792 6856 824
rect 6762 756 6856 792
rect 6762 724 6776 756
rect 6808 724 6856 756
rect 6762 688 6856 724
rect 6762 656 6776 688
rect 6808 656 6856 688
rect 6762 620 6856 656
rect 6762 588 6776 620
rect 6808 588 6856 620
rect 6762 550 6856 588
rect 6976 1844 7212 1882
rect 6976 1812 7078 1844
rect 7110 1812 7212 1844
rect 6976 1776 7212 1812
rect 6976 1744 7078 1776
rect 7110 1744 7212 1776
rect 6976 1708 7212 1744
rect 6976 1676 7078 1708
rect 7110 1676 7212 1708
rect 6976 1640 7212 1676
rect 6976 1608 7078 1640
rect 7110 1608 7212 1640
rect 6976 1572 7212 1608
rect 6976 1540 7078 1572
rect 7110 1540 7212 1572
rect 6976 1504 7212 1540
rect 6976 1472 7078 1504
rect 7110 1472 7212 1504
rect 6976 1436 7212 1472
rect 6976 1404 7078 1436
rect 7110 1404 7212 1436
rect 6976 1368 7212 1404
rect 6976 1336 7078 1368
rect 7110 1336 7212 1368
rect 6976 1300 7212 1336
rect 6976 1268 7078 1300
rect 7110 1268 7212 1300
rect 6976 1232 7212 1268
rect 6976 1200 7078 1232
rect 7110 1200 7212 1232
rect 6976 1164 7212 1200
rect 6976 1132 7078 1164
rect 7110 1132 7212 1164
rect 6976 1096 7212 1132
rect 6976 1064 7078 1096
rect 7110 1064 7212 1096
rect 6976 1028 7212 1064
rect 6976 996 7078 1028
rect 7110 996 7212 1028
rect 6976 960 7212 996
rect 6976 928 7078 960
rect 7110 928 7212 960
rect 6976 892 7212 928
rect 6976 860 7078 892
rect 7110 860 7212 892
rect 6976 824 7212 860
rect 6976 792 7078 824
rect 7110 792 7212 824
rect 6976 756 7212 792
rect 6976 724 7078 756
rect 7110 724 7212 756
rect 6976 688 7212 724
rect 6976 656 7078 688
rect 7110 656 7212 688
rect 6976 620 7212 656
rect 6976 588 7078 620
rect 7110 588 7212 620
rect 6976 550 7212 588
rect 7332 1844 7460 1882
rect 7332 1812 7380 1844
rect 7412 1812 7460 1844
rect 7332 1776 7460 1812
rect 7332 1744 7380 1776
rect 7412 1744 7460 1776
rect 7332 1708 7460 1744
rect 7332 1676 7380 1708
rect 7412 1676 7460 1708
rect 7332 1640 7460 1676
rect 7332 1608 7380 1640
rect 7412 1608 7460 1640
rect 7332 1572 7460 1608
rect 7332 1540 7380 1572
rect 7412 1540 7460 1572
rect 7332 1504 7460 1540
rect 7332 1472 7380 1504
rect 7412 1472 7460 1504
rect 7332 1436 7460 1472
rect 7332 1404 7380 1436
rect 7412 1404 7460 1436
rect 7332 1368 7460 1404
rect 7332 1336 7380 1368
rect 7412 1336 7460 1368
rect 7332 1300 7460 1336
rect 7332 1268 7380 1300
rect 7412 1268 7460 1300
rect 7332 1232 7460 1268
rect 7332 1200 7380 1232
rect 7412 1200 7460 1232
rect 7332 1164 7460 1200
rect 7332 1132 7380 1164
rect 7412 1132 7460 1164
rect 7332 1096 7460 1132
rect 7332 1064 7380 1096
rect 7412 1064 7460 1096
rect 7332 1028 7460 1064
rect 7332 996 7380 1028
rect 7412 996 7460 1028
rect 7332 960 7460 996
rect 7332 928 7380 960
rect 7412 928 7460 960
rect 7332 892 7460 928
rect 7332 860 7380 892
rect 7412 860 7460 892
rect 7332 824 7460 860
rect 7332 792 7380 824
rect 7412 792 7460 824
rect 7332 756 7460 792
rect 7332 724 7380 756
rect 7412 724 7460 756
rect 7332 688 7460 724
rect 7332 656 7380 688
rect 7412 656 7460 688
rect 7332 620 7460 656
rect 7332 588 7380 620
rect 7412 588 7460 620
rect 7332 550 7460 588
rect 7580 1844 7816 1882
rect 7580 1812 7682 1844
rect 7714 1812 7816 1844
rect 7580 1776 7816 1812
rect 7580 1744 7682 1776
rect 7714 1744 7816 1776
rect 7580 1708 7816 1744
rect 7580 1676 7682 1708
rect 7714 1676 7816 1708
rect 7580 1640 7816 1676
rect 7580 1608 7682 1640
rect 7714 1608 7816 1640
rect 7580 1572 7816 1608
rect 7580 1540 7682 1572
rect 7714 1540 7816 1572
rect 7580 1504 7816 1540
rect 7580 1472 7682 1504
rect 7714 1472 7816 1504
rect 7580 1436 7816 1472
rect 7580 1404 7682 1436
rect 7714 1404 7816 1436
rect 7580 1368 7816 1404
rect 7580 1336 7682 1368
rect 7714 1336 7816 1368
rect 7580 1300 7816 1336
rect 7580 1268 7682 1300
rect 7714 1268 7816 1300
rect 7580 1232 7816 1268
rect 7580 1200 7682 1232
rect 7714 1200 7816 1232
rect 7580 1164 7816 1200
rect 7580 1132 7682 1164
rect 7714 1132 7816 1164
rect 7580 1096 7816 1132
rect 7580 1064 7682 1096
rect 7714 1064 7816 1096
rect 7580 1028 7816 1064
rect 7580 996 7682 1028
rect 7714 996 7816 1028
rect 7580 960 7816 996
rect 7580 928 7682 960
rect 7714 928 7816 960
rect 7580 892 7816 928
rect 7580 860 7682 892
rect 7714 860 7816 892
rect 7580 824 7816 860
rect 7580 792 7682 824
rect 7714 792 7816 824
rect 7580 756 7816 792
rect 7580 724 7682 756
rect 7714 724 7816 756
rect 7580 688 7816 724
rect 7580 656 7682 688
rect 7714 656 7816 688
rect 7580 620 7816 656
rect 7580 588 7682 620
rect 7714 588 7816 620
rect 7580 550 7816 588
rect 7936 1844 8064 1882
rect 7936 1812 7984 1844
rect 8016 1812 8064 1844
rect 7936 1776 8064 1812
rect 7936 1744 7984 1776
rect 8016 1744 8064 1776
rect 7936 1708 8064 1744
rect 7936 1676 7984 1708
rect 8016 1676 8064 1708
rect 7936 1640 8064 1676
rect 7936 1608 7984 1640
rect 8016 1608 8064 1640
rect 7936 1572 8064 1608
rect 7936 1540 7984 1572
rect 8016 1540 8064 1572
rect 7936 1504 8064 1540
rect 7936 1472 7984 1504
rect 8016 1472 8064 1504
rect 7936 1436 8064 1472
rect 7936 1404 7984 1436
rect 8016 1404 8064 1436
rect 7936 1368 8064 1404
rect 7936 1336 7984 1368
rect 8016 1336 8064 1368
rect 7936 1300 8064 1336
rect 7936 1268 7984 1300
rect 8016 1268 8064 1300
rect 7936 1232 8064 1268
rect 7936 1200 7984 1232
rect 8016 1200 8064 1232
rect 7936 1164 8064 1200
rect 7936 1132 7984 1164
rect 8016 1132 8064 1164
rect 7936 1096 8064 1132
rect 7936 1064 7984 1096
rect 8016 1064 8064 1096
rect 7936 1028 8064 1064
rect 7936 996 7984 1028
rect 8016 996 8064 1028
rect 7936 960 8064 996
rect 7936 928 7984 960
rect 8016 928 8064 960
rect 7936 892 8064 928
rect 7936 860 7984 892
rect 8016 860 8064 892
rect 7936 824 8064 860
rect 7936 792 7984 824
rect 8016 792 8064 824
rect 7936 756 8064 792
rect 7936 724 7984 756
rect 8016 724 8064 756
rect 7936 688 8064 724
rect 7936 656 7984 688
rect 8016 656 8064 688
rect 7936 620 8064 656
rect 7936 588 7984 620
rect 8016 588 8064 620
rect 7936 550 8064 588
rect 8184 1844 8420 1882
rect 8184 1812 8286 1844
rect 8318 1812 8420 1844
rect 8184 1776 8420 1812
rect 8184 1744 8286 1776
rect 8318 1744 8420 1776
rect 8184 1708 8420 1744
rect 8184 1676 8286 1708
rect 8318 1676 8420 1708
rect 8184 1640 8420 1676
rect 8184 1608 8286 1640
rect 8318 1608 8420 1640
rect 8184 1572 8420 1608
rect 8184 1540 8286 1572
rect 8318 1540 8420 1572
rect 8184 1504 8420 1540
rect 8184 1472 8286 1504
rect 8318 1472 8420 1504
rect 8184 1436 8420 1472
rect 8184 1404 8286 1436
rect 8318 1404 8420 1436
rect 8184 1368 8420 1404
rect 8184 1336 8286 1368
rect 8318 1336 8420 1368
rect 8184 1300 8420 1336
rect 8184 1268 8286 1300
rect 8318 1268 8420 1300
rect 8184 1232 8420 1268
rect 8184 1200 8286 1232
rect 8318 1200 8420 1232
rect 8184 1164 8420 1200
rect 8184 1132 8286 1164
rect 8318 1132 8420 1164
rect 8184 1096 8420 1132
rect 8184 1064 8286 1096
rect 8318 1064 8420 1096
rect 8184 1028 8420 1064
rect 8184 996 8286 1028
rect 8318 996 8420 1028
rect 8184 960 8420 996
rect 8184 928 8286 960
rect 8318 928 8420 960
rect 8184 892 8420 928
rect 8184 860 8286 892
rect 8318 860 8420 892
rect 8184 824 8420 860
rect 8184 792 8286 824
rect 8318 792 8420 824
rect 8184 756 8420 792
rect 8184 724 8286 756
rect 8318 724 8420 756
rect 8184 688 8420 724
rect 8184 656 8286 688
rect 8318 656 8420 688
rect 8184 620 8420 656
rect 8184 588 8286 620
rect 8318 588 8420 620
rect 8184 550 8420 588
rect 8540 1844 8668 1882
rect 8540 1812 8588 1844
rect 8620 1812 8668 1844
rect 8540 1776 8668 1812
rect 8540 1744 8588 1776
rect 8620 1744 8668 1776
rect 8540 1708 8668 1744
rect 8540 1676 8588 1708
rect 8620 1676 8668 1708
rect 8540 1640 8668 1676
rect 8540 1608 8588 1640
rect 8620 1608 8668 1640
rect 8540 1572 8668 1608
rect 8540 1540 8588 1572
rect 8620 1540 8668 1572
rect 8540 1504 8668 1540
rect 8540 1472 8588 1504
rect 8620 1472 8668 1504
rect 8540 1436 8668 1472
rect 8540 1404 8588 1436
rect 8620 1404 8668 1436
rect 8540 1368 8668 1404
rect 8540 1336 8588 1368
rect 8620 1336 8668 1368
rect 8540 1300 8668 1336
rect 8540 1268 8588 1300
rect 8620 1268 8668 1300
rect 8540 1232 8668 1268
rect 8540 1200 8588 1232
rect 8620 1200 8668 1232
rect 8540 1164 8668 1200
rect 8540 1132 8588 1164
rect 8620 1132 8668 1164
rect 8540 1096 8668 1132
rect 8540 1064 8588 1096
rect 8620 1064 8668 1096
rect 8540 1028 8668 1064
rect 8540 996 8588 1028
rect 8620 996 8668 1028
rect 8540 960 8668 996
rect 8540 928 8588 960
rect 8620 928 8668 960
rect 8540 892 8668 928
rect 8540 860 8588 892
rect 8620 860 8668 892
rect 8540 824 8668 860
rect 8540 792 8588 824
rect 8620 792 8668 824
rect 8540 756 8668 792
rect 8540 724 8588 756
rect 8620 724 8668 756
rect 8540 688 8668 724
rect 8540 656 8588 688
rect 8620 656 8668 688
rect 8540 620 8668 656
rect 8540 588 8588 620
rect 8620 588 8668 620
rect 8540 550 8668 588
rect 8788 1844 9024 1882
rect 8788 1812 8890 1844
rect 8922 1812 9024 1844
rect 8788 1776 9024 1812
rect 8788 1744 8890 1776
rect 8922 1744 9024 1776
rect 8788 1708 9024 1744
rect 8788 1676 8890 1708
rect 8922 1676 9024 1708
rect 8788 1640 9024 1676
rect 8788 1608 8890 1640
rect 8922 1608 9024 1640
rect 8788 1572 9024 1608
rect 8788 1540 8890 1572
rect 8922 1540 9024 1572
rect 8788 1504 9024 1540
rect 8788 1472 8890 1504
rect 8922 1472 9024 1504
rect 8788 1436 9024 1472
rect 8788 1404 8890 1436
rect 8922 1404 9024 1436
rect 8788 1368 9024 1404
rect 8788 1336 8890 1368
rect 8922 1336 9024 1368
rect 8788 1300 9024 1336
rect 8788 1268 8890 1300
rect 8922 1268 9024 1300
rect 8788 1232 9024 1268
rect 8788 1200 8890 1232
rect 8922 1200 9024 1232
rect 8788 1164 9024 1200
rect 8788 1132 8890 1164
rect 8922 1132 9024 1164
rect 8788 1096 9024 1132
rect 8788 1064 8890 1096
rect 8922 1064 9024 1096
rect 8788 1028 9024 1064
rect 8788 996 8890 1028
rect 8922 996 9024 1028
rect 8788 960 9024 996
rect 8788 928 8890 960
rect 8922 928 9024 960
rect 8788 892 9024 928
rect 8788 860 8890 892
rect 8922 860 9024 892
rect 8788 824 9024 860
rect 8788 792 8890 824
rect 8922 792 9024 824
rect 8788 756 9024 792
rect 8788 724 8890 756
rect 8922 724 9024 756
rect 8788 688 9024 724
rect 8788 656 8890 688
rect 8922 656 9024 688
rect 8788 620 9024 656
rect 8788 588 8890 620
rect 8922 588 9024 620
rect 8788 550 9024 588
rect 9144 1844 9238 1882
rect 9144 1812 9192 1844
rect 9224 1812 9238 1844
rect 9144 1776 9238 1812
rect 9144 1744 9192 1776
rect 9224 1744 9238 1776
rect 9144 1708 9238 1744
rect 9144 1676 9192 1708
rect 9224 1676 9238 1708
rect 9144 1640 9238 1676
rect 9144 1608 9192 1640
rect 9224 1608 9238 1640
rect 9144 1572 9238 1608
rect 9144 1540 9192 1572
rect 9224 1540 9238 1572
rect 9144 1504 9238 1540
rect 9144 1472 9192 1504
rect 9224 1472 9238 1504
rect 9144 1436 9238 1472
rect 9144 1404 9192 1436
rect 9224 1404 9238 1436
rect 9144 1368 9238 1404
rect 9144 1336 9192 1368
rect 9224 1336 9238 1368
rect 9144 1300 9238 1336
rect 9144 1268 9192 1300
rect 9224 1268 9238 1300
rect 9144 1232 9238 1268
rect 9144 1200 9192 1232
rect 9224 1200 9238 1232
rect 9144 1164 9238 1200
rect 9144 1132 9192 1164
rect 9224 1132 9238 1164
rect 9144 1096 9238 1132
rect 9144 1064 9192 1096
rect 9224 1064 9238 1096
rect 9144 1028 9238 1064
rect 9144 996 9192 1028
rect 9224 996 9238 1028
rect 9144 960 9238 996
rect 9144 928 9192 960
rect 9224 928 9238 960
rect 9144 892 9238 928
rect 9144 860 9192 892
rect 9224 860 9238 892
rect 9144 824 9238 860
rect 9144 792 9192 824
rect 9224 792 9238 824
rect 9144 756 9238 792
rect 9144 724 9192 756
rect 9224 724 9238 756
rect 9144 688 9238 724
rect 9144 656 9192 688
rect 9224 656 9238 688
rect 9144 620 9238 656
rect 9144 588 9192 620
rect 9224 588 9238 620
rect 9144 550 9238 588
<< hvpdiffc >>
rect 6776 3232 6808 3264
rect 6776 3164 6808 3196
rect 6776 3096 6808 3128
rect 6776 3028 6808 3060
rect 6776 2960 6808 2992
rect 6776 2892 6808 2924
rect 6776 2824 6808 2856
rect 6776 2756 6808 2788
rect 6776 2688 6808 2720
rect 6776 2620 6808 2652
rect 6776 2552 6808 2584
rect 6776 2484 6808 2516
rect 6776 2416 6808 2448
rect 6776 2348 6808 2380
rect 6776 2280 6808 2312
rect 6776 2212 6808 2244
rect 6776 2144 6808 2176
rect 6776 2076 6808 2108
rect 6776 2008 6808 2040
rect 7078 3232 7110 3264
rect 7078 3164 7110 3196
rect 7078 3096 7110 3128
rect 7078 3028 7110 3060
rect 7078 2960 7110 2992
rect 7078 2892 7110 2924
rect 7078 2824 7110 2856
rect 7078 2756 7110 2788
rect 7078 2688 7110 2720
rect 7078 2620 7110 2652
rect 7078 2552 7110 2584
rect 7078 2484 7110 2516
rect 7078 2416 7110 2448
rect 7078 2348 7110 2380
rect 7078 2280 7110 2312
rect 7078 2212 7110 2244
rect 7078 2144 7110 2176
rect 7078 2076 7110 2108
rect 7078 2008 7110 2040
rect 7380 3232 7412 3264
rect 7380 3164 7412 3196
rect 7380 3096 7412 3128
rect 7380 3028 7412 3060
rect 7380 2960 7412 2992
rect 7380 2892 7412 2924
rect 7380 2824 7412 2856
rect 7380 2756 7412 2788
rect 7380 2688 7412 2720
rect 7380 2620 7412 2652
rect 7380 2552 7412 2584
rect 7380 2484 7412 2516
rect 7380 2416 7412 2448
rect 7380 2348 7412 2380
rect 7380 2280 7412 2312
rect 7380 2212 7412 2244
rect 7380 2144 7412 2176
rect 7380 2076 7412 2108
rect 7380 2008 7412 2040
rect 7682 3232 7714 3264
rect 7682 3164 7714 3196
rect 7682 3096 7714 3128
rect 7682 3028 7714 3060
rect 7682 2960 7714 2992
rect 7682 2892 7714 2924
rect 7682 2824 7714 2856
rect 7682 2756 7714 2788
rect 7682 2688 7714 2720
rect 7682 2620 7714 2652
rect 7682 2552 7714 2584
rect 7682 2484 7714 2516
rect 7682 2416 7714 2448
rect 7682 2348 7714 2380
rect 7682 2280 7714 2312
rect 7682 2212 7714 2244
rect 7682 2144 7714 2176
rect 7682 2076 7714 2108
rect 7682 2008 7714 2040
rect 7984 3232 8016 3264
rect 7984 3164 8016 3196
rect 7984 3096 8016 3128
rect 7984 3028 8016 3060
rect 7984 2960 8016 2992
rect 7984 2892 8016 2924
rect 7984 2824 8016 2856
rect 7984 2756 8016 2788
rect 7984 2688 8016 2720
rect 7984 2620 8016 2652
rect 7984 2552 8016 2584
rect 7984 2484 8016 2516
rect 7984 2416 8016 2448
rect 7984 2348 8016 2380
rect 7984 2280 8016 2312
rect 7984 2212 8016 2244
rect 7984 2144 8016 2176
rect 7984 2076 8016 2108
rect 7984 2008 8016 2040
rect 8286 3232 8318 3264
rect 8286 3164 8318 3196
rect 8286 3096 8318 3128
rect 8286 3028 8318 3060
rect 8286 2960 8318 2992
rect 8286 2892 8318 2924
rect 8286 2824 8318 2856
rect 8286 2756 8318 2788
rect 8286 2688 8318 2720
rect 8286 2620 8318 2652
rect 8286 2552 8318 2584
rect 8286 2484 8318 2516
rect 8286 2416 8318 2448
rect 8286 2348 8318 2380
rect 8286 2280 8318 2312
rect 8286 2212 8318 2244
rect 8286 2144 8318 2176
rect 8286 2076 8318 2108
rect 8286 2008 8318 2040
rect 8588 3232 8620 3264
rect 8588 3164 8620 3196
rect 8588 3096 8620 3128
rect 8588 3028 8620 3060
rect 8588 2960 8620 2992
rect 8588 2892 8620 2924
rect 8588 2824 8620 2856
rect 8588 2756 8620 2788
rect 8588 2688 8620 2720
rect 8588 2620 8620 2652
rect 8588 2552 8620 2584
rect 8588 2484 8620 2516
rect 8588 2416 8620 2448
rect 8588 2348 8620 2380
rect 8588 2280 8620 2312
rect 8588 2212 8620 2244
rect 8588 2144 8620 2176
rect 8588 2076 8620 2108
rect 8588 2008 8620 2040
rect 8890 3232 8922 3264
rect 8890 3164 8922 3196
rect 8890 3096 8922 3128
rect 8890 3028 8922 3060
rect 8890 2960 8922 2992
rect 8890 2892 8922 2924
rect 8890 2824 8922 2856
rect 8890 2756 8922 2788
rect 8890 2688 8922 2720
rect 8890 2620 8922 2652
rect 8890 2552 8922 2584
rect 8890 2484 8922 2516
rect 8890 2416 8922 2448
rect 8890 2348 8922 2380
rect 8890 2280 8922 2312
rect 8890 2212 8922 2244
rect 8890 2144 8922 2176
rect 8890 2076 8922 2108
rect 8890 2008 8922 2040
rect 9192 3232 9224 3264
rect 9192 3164 9224 3196
rect 9192 3096 9224 3128
rect 9192 3028 9224 3060
rect 9192 2960 9224 2992
rect 9192 2892 9224 2924
rect 9192 2824 9224 2856
rect 9192 2756 9224 2788
rect 9192 2688 9224 2720
rect 9192 2620 9224 2652
rect 9192 2552 9224 2584
rect 9192 2484 9224 2516
rect 9192 2416 9224 2448
rect 9192 2348 9224 2380
rect 9192 2280 9224 2312
rect 9192 2212 9224 2244
rect 9192 2144 9224 2176
rect 9192 2076 9224 2108
rect 9192 2008 9224 2040
rect 6776 1812 6808 1844
rect 6776 1744 6808 1776
rect 6776 1676 6808 1708
rect 6776 1608 6808 1640
rect 6776 1540 6808 1572
rect 6776 1472 6808 1504
rect 6776 1404 6808 1436
rect 6776 1336 6808 1368
rect 6776 1268 6808 1300
rect 6776 1200 6808 1232
rect 6776 1132 6808 1164
rect 6776 1064 6808 1096
rect 6776 996 6808 1028
rect 6776 928 6808 960
rect 6776 860 6808 892
rect 6776 792 6808 824
rect 6776 724 6808 756
rect 6776 656 6808 688
rect 6776 588 6808 620
rect 7078 1812 7110 1844
rect 7078 1744 7110 1776
rect 7078 1676 7110 1708
rect 7078 1608 7110 1640
rect 7078 1540 7110 1572
rect 7078 1472 7110 1504
rect 7078 1404 7110 1436
rect 7078 1336 7110 1368
rect 7078 1268 7110 1300
rect 7078 1200 7110 1232
rect 7078 1132 7110 1164
rect 7078 1064 7110 1096
rect 7078 996 7110 1028
rect 7078 928 7110 960
rect 7078 860 7110 892
rect 7078 792 7110 824
rect 7078 724 7110 756
rect 7078 656 7110 688
rect 7078 588 7110 620
rect 7380 1812 7412 1844
rect 7380 1744 7412 1776
rect 7380 1676 7412 1708
rect 7380 1608 7412 1640
rect 7380 1540 7412 1572
rect 7380 1472 7412 1504
rect 7380 1404 7412 1436
rect 7380 1336 7412 1368
rect 7380 1268 7412 1300
rect 7380 1200 7412 1232
rect 7380 1132 7412 1164
rect 7380 1064 7412 1096
rect 7380 996 7412 1028
rect 7380 928 7412 960
rect 7380 860 7412 892
rect 7380 792 7412 824
rect 7380 724 7412 756
rect 7380 656 7412 688
rect 7380 588 7412 620
rect 7682 1812 7714 1844
rect 7682 1744 7714 1776
rect 7682 1676 7714 1708
rect 7682 1608 7714 1640
rect 7682 1540 7714 1572
rect 7682 1472 7714 1504
rect 7682 1404 7714 1436
rect 7682 1336 7714 1368
rect 7682 1268 7714 1300
rect 7682 1200 7714 1232
rect 7682 1132 7714 1164
rect 7682 1064 7714 1096
rect 7682 996 7714 1028
rect 7682 928 7714 960
rect 7682 860 7714 892
rect 7682 792 7714 824
rect 7682 724 7714 756
rect 7682 656 7714 688
rect 7682 588 7714 620
rect 7984 1812 8016 1844
rect 7984 1744 8016 1776
rect 7984 1676 8016 1708
rect 7984 1608 8016 1640
rect 7984 1540 8016 1572
rect 7984 1472 8016 1504
rect 7984 1404 8016 1436
rect 7984 1336 8016 1368
rect 7984 1268 8016 1300
rect 7984 1200 8016 1232
rect 7984 1132 8016 1164
rect 7984 1064 8016 1096
rect 7984 996 8016 1028
rect 7984 928 8016 960
rect 7984 860 8016 892
rect 7984 792 8016 824
rect 7984 724 8016 756
rect 7984 656 8016 688
rect 7984 588 8016 620
rect 8286 1812 8318 1844
rect 8286 1744 8318 1776
rect 8286 1676 8318 1708
rect 8286 1608 8318 1640
rect 8286 1540 8318 1572
rect 8286 1472 8318 1504
rect 8286 1404 8318 1436
rect 8286 1336 8318 1368
rect 8286 1268 8318 1300
rect 8286 1200 8318 1232
rect 8286 1132 8318 1164
rect 8286 1064 8318 1096
rect 8286 996 8318 1028
rect 8286 928 8318 960
rect 8286 860 8318 892
rect 8286 792 8318 824
rect 8286 724 8318 756
rect 8286 656 8318 688
rect 8286 588 8318 620
rect 8588 1812 8620 1844
rect 8588 1744 8620 1776
rect 8588 1676 8620 1708
rect 8588 1608 8620 1640
rect 8588 1540 8620 1572
rect 8588 1472 8620 1504
rect 8588 1404 8620 1436
rect 8588 1336 8620 1368
rect 8588 1268 8620 1300
rect 8588 1200 8620 1232
rect 8588 1132 8620 1164
rect 8588 1064 8620 1096
rect 8588 996 8620 1028
rect 8588 928 8620 960
rect 8588 860 8620 892
rect 8588 792 8620 824
rect 8588 724 8620 756
rect 8588 656 8620 688
rect 8588 588 8620 620
rect 8890 1812 8922 1844
rect 8890 1744 8922 1776
rect 8890 1676 8922 1708
rect 8890 1608 8922 1640
rect 8890 1540 8922 1572
rect 8890 1472 8922 1504
rect 8890 1404 8922 1436
rect 8890 1336 8922 1368
rect 8890 1268 8922 1300
rect 8890 1200 8922 1232
rect 8890 1132 8922 1164
rect 8890 1064 8922 1096
rect 8890 996 8922 1028
rect 8890 928 8922 960
rect 8890 860 8922 892
rect 8890 792 8922 824
rect 8890 724 8922 756
rect 8890 656 8922 688
rect 8890 588 8922 620
rect 9192 1812 9224 1844
rect 9192 1744 9224 1776
rect 9192 1676 9224 1708
rect 9192 1608 9224 1640
rect 9192 1540 9224 1572
rect 9192 1472 9224 1504
rect 9192 1404 9224 1436
rect 9192 1336 9224 1368
rect 9192 1268 9224 1300
rect 9192 1200 9224 1232
rect 9192 1132 9224 1164
rect 9192 1064 9224 1096
rect 9192 996 9224 1028
rect 9192 928 9224 960
rect 9192 860 9224 892
rect 9192 792 9224 824
rect 9192 724 9224 756
rect 9192 656 9224 688
rect 9192 588 9224 620
<< psubdiff >>
rect 0 3834 16000 3852
rect 0 3802 28 3834
rect 60 3802 96 3834
rect 128 3802 164 3834
rect 196 3802 232 3834
rect 264 3802 300 3834
rect 332 3802 368 3834
rect 400 3802 436 3834
rect 468 3802 504 3834
rect 536 3802 572 3834
rect 604 3802 640 3834
rect 672 3802 708 3834
rect 740 3802 776 3834
rect 808 3802 844 3834
rect 876 3802 912 3834
rect 944 3802 980 3834
rect 1012 3802 1048 3834
rect 1080 3802 1116 3834
rect 1148 3802 1184 3834
rect 1216 3802 1252 3834
rect 1284 3802 1320 3834
rect 1352 3802 1388 3834
rect 1420 3802 1456 3834
rect 1488 3802 1524 3834
rect 1556 3802 1592 3834
rect 1624 3802 1660 3834
rect 1692 3802 1728 3834
rect 1760 3802 1796 3834
rect 1828 3802 1864 3834
rect 1896 3802 1932 3834
rect 1964 3802 2000 3834
rect 2032 3802 2068 3834
rect 2100 3802 2136 3834
rect 2168 3802 2204 3834
rect 2236 3802 2272 3834
rect 2304 3802 2340 3834
rect 2372 3802 2408 3834
rect 2440 3802 2476 3834
rect 2508 3802 2544 3834
rect 2576 3802 2612 3834
rect 2644 3802 2680 3834
rect 2712 3802 2748 3834
rect 2780 3802 2816 3834
rect 2848 3802 2884 3834
rect 2916 3802 2952 3834
rect 2984 3802 3020 3834
rect 3052 3802 3088 3834
rect 3120 3802 3156 3834
rect 3188 3802 3224 3834
rect 3256 3802 3292 3834
rect 3324 3802 3360 3834
rect 3392 3802 3428 3834
rect 3460 3802 3496 3834
rect 3528 3802 3564 3834
rect 3596 3802 3632 3834
rect 3664 3802 3700 3834
rect 3732 3802 3768 3834
rect 3800 3802 3836 3834
rect 3868 3802 3904 3834
rect 3936 3802 3972 3834
rect 4004 3802 4040 3834
rect 4072 3802 4108 3834
rect 4140 3802 4176 3834
rect 4208 3802 4244 3834
rect 4276 3802 4312 3834
rect 4344 3802 4380 3834
rect 4412 3802 4448 3834
rect 4480 3802 4516 3834
rect 4548 3802 4584 3834
rect 4616 3802 4652 3834
rect 4684 3802 4720 3834
rect 4752 3802 4788 3834
rect 4820 3802 4856 3834
rect 4888 3802 4924 3834
rect 4956 3802 4992 3834
rect 5024 3802 5060 3834
rect 5092 3802 5128 3834
rect 5160 3802 5196 3834
rect 5228 3802 5264 3834
rect 5296 3802 5332 3834
rect 5364 3802 5400 3834
rect 5432 3802 5468 3834
rect 5500 3802 5536 3834
rect 5568 3802 5604 3834
rect 5636 3802 5672 3834
rect 5704 3802 5740 3834
rect 5772 3802 5808 3834
rect 5840 3802 5876 3834
rect 5908 3802 5944 3834
rect 5976 3802 6012 3834
rect 6044 3802 6080 3834
rect 6112 3802 6148 3834
rect 6180 3802 6216 3834
rect 6248 3802 6284 3834
rect 6316 3802 6352 3834
rect 6384 3802 6420 3834
rect 6452 3802 6488 3834
rect 6520 3802 6556 3834
rect 6588 3802 6624 3834
rect 6656 3802 6692 3834
rect 6724 3802 6760 3834
rect 6792 3802 6828 3834
rect 6860 3802 6896 3834
rect 6928 3802 6964 3834
rect 6996 3802 7032 3834
rect 7064 3802 7100 3834
rect 7132 3802 7168 3834
rect 7200 3802 7236 3834
rect 7268 3802 7304 3834
rect 7336 3802 7372 3834
rect 7404 3802 7440 3834
rect 7472 3802 7508 3834
rect 7540 3802 7576 3834
rect 7608 3802 7644 3834
rect 7676 3802 7712 3834
rect 7744 3802 7780 3834
rect 7812 3802 7848 3834
rect 7880 3802 7916 3834
rect 7948 3802 7984 3834
rect 8016 3802 8052 3834
rect 8084 3802 8120 3834
rect 8152 3802 8188 3834
rect 8220 3802 8256 3834
rect 8288 3802 8324 3834
rect 8356 3802 8392 3834
rect 8424 3802 8460 3834
rect 8492 3802 8528 3834
rect 8560 3802 8596 3834
rect 8628 3802 8664 3834
rect 8696 3802 8732 3834
rect 8764 3802 8800 3834
rect 8832 3802 8868 3834
rect 8900 3802 8936 3834
rect 8968 3802 9004 3834
rect 9036 3802 9072 3834
rect 9104 3802 9140 3834
rect 9172 3802 9208 3834
rect 9240 3802 9276 3834
rect 9308 3802 9344 3834
rect 9376 3802 9412 3834
rect 9444 3802 9480 3834
rect 9512 3802 9548 3834
rect 9580 3802 9616 3834
rect 9648 3802 9684 3834
rect 9716 3802 9752 3834
rect 9784 3802 9820 3834
rect 9852 3802 9888 3834
rect 9920 3802 9956 3834
rect 9988 3802 10024 3834
rect 10056 3802 10092 3834
rect 10124 3802 10160 3834
rect 10192 3802 10228 3834
rect 10260 3802 10296 3834
rect 10328 3802 10364 3834
rect 10396 3802 10432 3834
rect 10464 3802 10500 3834
rect 10532 3802 10568 3834
rect 10600 3802 10636 3834
rect 10668 3802 10704 3834
rect 10736 3802 10772 3834
rect 10804 3802 10840 3834
rect 10872 3802 10908 3834
rect 10940 3802 10976 3834
rect 11008 3802 11044 3834
rect 11076 3802 11112 3834
rect 11144 3802 11180 3834
rect 11212 3802 11248 3834
rect 11280 3802 11316 3834
rect 11348 3802 11384 3834
rect 11416 3802 11452 3834
rect 11484 3802 11520 3834
rect 11552 3802 11588 3834
rect 11620 3802 11656 3834
rect 11688 3802 11724 3834
rect 11756 3802 11792 3834
rect 11824 3802 11860 3834
rect 11892 3802 11928 3834
rect 11960 3802 11996 3834
rect 12028 3802 12064 3834
rect 12096 3802 12132 3834
rect 12164 3802 12200 3834
rect 12232 3802 12268 3834
rect 12300 3802 12336 3834
rect 12368 3802 12404 3834
rect 12436 3802 12472 3834
rect 12504 3802 12540 3834
rect 12572 3802 12608 3834
rect 12640 3802 12676 3834
rect 12708 3802 12744 3834
rect 12776 3802 12812 3834
rect 12844 3802 12880 3834
rect 12912 3802 12948 3834
rect 12980 3802 13016 3834
rect 13048 3802 13084 3834
rect 13116 3802 13152 3834
rect 13184 3802 13220 3834
rect 13252 3802 13288 3834
rect 13320 3802 13356 3834
rect 13388 3802 13424 3834
rect 13456 3802 13492 3834
rect 13524 3802 13560 3834
rect 13592 3802 13628 3834
rect 13660 3802 13696 3834
rect 13728 3802 13764 3834
rect 13796 3802 13832 3834
rect 13864 3802 13900 3834
rect 13932 3802 13968 3834
rect 14000 3802 14036 3834
rect 14068 3802 14104 3834
rect 14136 3802 14172 3834
rect 14204 3802 14240 3834
rect 14272 3802 14308 3834
rect 14340 3802 14376 3834
rect 14408 3802 14444 3834
rect 14476 3802 14512 3834
rect 14544 3802 14580 3834
rect 14612 3802 14648 3834
rect 14680 3802 14716 3834
rect 14748 3802 14784 3834
rect 14816 3802 14852 3834
rect 14884 3802 14920 3834
rect 14952 3802 14988 3834
rect 15020 3802 15056 3834
rect 15088 3802 15124 3834
rect 15156 3802 15192 3834
rect 15224 3802 15260 3834
rect 15292 3802 15328 3834
rect 15360 3802 15396 3834
rect 15428 3802 15464 3834
rect 15496 3802 15532 3834
rect 15564 3802 15600 3834
rect 15632 3802 15668 3834
rect 15700 3802 15736 3834
rect 15768 3802 15804 3834
rect 15836 3802 15872 3834
rect 15904 3802 15940 3834
rect 15972 3802 16000 3834
rect 0 3784 16000 3802
rect 0 3744 68 3784
rect 0 3712 18 3744
rect 50 3712 68 3744
rect 0 3676 68 3712
rect 0 3644 18 3676
rect 50 3644 68 3676
rect 0 3608 68 3644
rect 0 3576 18 3608
rect 50 3576 68 3608
rect 0 3540 68 3576
rect 0 3508 18 3540
rect 50 3508 68 3540
rect 0 3472 68 3508
rect 15932 3744 16000 3784
rect 15932 3712 15950 3744
rect 15982 3712 16000 3744
rect 15932 3676 16000 3712
rect 15932 3644 15950 3676
rect 15982 3644 16000 3676
rect 15932 3608 16000 3644
rect 15932 3576 15950 3608
rect 15982 3576 16000 3608
rect 15932 3540 16000 3576
rect 15932 3508 15950 3540
rect 15982 3508 16000 3540
rect 0 3440 18 3472
rect 50 3440 68 3472
rect 0 3404 68 3440
rect 0 3372 18 3404
rect 50 3372 68 3404
rect 0 3336 68 3372
rect 0 3304 18 3336
rect 50 3304 68 3336
rect 0 3268 68 3304
rect 0 3236 18 3268
rect 50 3236 68 3268
rect 0 3200 68 3236
rect 0 3168 18 3200
rect 50 3168 68 3200
rect 0 3132 68 3168
rect 0 3100 18 3132
rect 50 3100 68 3132
rect 0 3064 68 3100
rect 0 3032 18 3064
rect 50 3032 68 3064
rect 0 2996 68 3032
rect 0 2964 18 2996
rect 50 2964 68 2996
rect 0 2928 68 2964
rect 0 2896 18 2928
rect 50 2896 68 2928
rect 0 2860 68 2896
rect 0 2828 18 2860
rect 50 2828 68 2860
rect 0 2792 68 2828
rect 0 2760 18 2792
rect 50 2760 68 2792
rect 0 2724 68 2760
rect 0 2692 18 2724
rect 50 2692 68 2724
rect 0 2656 68 2692
rect 0 2624 18 2656
rect 50 2624 68 2656
rect 0 2588 68 2624
rect 0 2556 18 2588
rect 50 2556 68 2588
rect 0 2520 68 2556
rect 0 2488 18 2520
rect 50 2488 68 2520
rect 0 2452 68 2488
rect 0 2420 18 2452
rect 50 2420 68 2452
rect 0 2384 68 2420
rect 0 2352 18 2384
rect 50 2352 68 2384
rect 0 2316 68 2352
rect 0 2284 18 2316
rect 50 2284 68 2316
rect 0 2248 68 2284
rect 0 2216 18 2248
rect 50 2216 68 2248
rect 0 2180 68 2216
rect 0 2148 18 2180
rect 50 2148 68 2180
rect 0 2112 68 2148
rect 0 2080 18 2112
rect 50 2080 68 2112
rect 0 2044 68 2080
rect 0 2012 18 2044
rect 50 2012 68 2044
rect 0 1976 68 2012
rect 0 1944 18 1976
rect 50 1944 68 1976
rect 0 1908 68 1944
rect 0 1876 18 1908
rect 50 1876 68 1908
rect 0 1840 68 1876
rect 0 1808 18 1840
rect 50 1808 68 1840
rect 0 1772 68 1808
rect 0 1740 18 1772
rect 50 1740 68 1772
rect 0 1704 68 1740
rect 0 1672 18 1704
rect 50 1672 68 1704
rect 0 1636 68 1672
rect 0 1604 18 1636
rect 50 1604 68 1636
rect 0 1568 68 1604
rect 0 1536 18 1568
rect 50 1536 68 1568
rect 0 1500 68 1536
rect 0 1468 18 1500
rect 50 1468 68 1500
rect 0 1432 68 1468
rect 0 1400 18 1432
rect 50 1400 68 1432
rect 0 1364 68 1400
rect 0 1332 18 1364
rect 50 1332 68 1364
rect 0 1296 68 1332
rect 0 1264 18 1296
rect 50 1264 68 1296
rect 0 1228 68 1264
rect 0 1196 18 1228
rect 50 1196 68 1228
rect 0 1160 68 1196
rect 0 1128 18 1160
rect 50 1128 68 1160
rect 0 1092 68 1128
rect 0 1060 18 1092
rect 50 1060 68 1092
rect 0 1024 68 1060
rect 0 992 18 1024
rect 50 992 68 1024
rect 0 956 68 992
rect 0 924 18 956
rect 50 924 68 956
rect 0 888 68 924
rect 0 856 18 888
rect 50 856 68 888
rect 0 820 68 856
rect 0 788 18 820
rect 50 788 68 820
rect 0 752 68 788
rect 0 720 18 752
rect 50 720 68 752
rect 0 684 68 720
rect 0 652 18 684
rect 50 652 68 684
rect 0 616 68 652
rect 0 584 18 616
rect 50 584 68 616
rect 0 548 68 584
rect 0 516 18 548
rect 50 516 68 548
rect 0 480 68 516
rect 0 448 18 480
rect 50 448 68 480
rect 0 412 68 448
rect 0 380 18 412
rect 50 380 68 412
rect 0 344 68 380
rect 15932 3472 16000 3508
rect 15932 3440 15950 3472
rect 15982 3440 16000 3472
rect 15932 3404 16000 3440
rect 15932 3372 15950 3404
rect 15982 3372 16000 3404
rect 15932 3336 16000 3372
rect 15932 3304 15950 3336
rect 15982 3304 16000 3336
rect 15932 3268 16000 3304
rect 15932 3236 15950 3268
rect 15982 3236 16000 3268
rect 15932 3200 16000 3236
rect 15932 3168 15950 3200
rect 15982 3168 16000 3200
rect 15932 3132 16000 3168
rect 15932 3100 15950 3132
rect 15982 3100 16000 3132
rect 15932 3064 16000 3100
rect 15932 3032 15950 3064
rect 15982 3032 16000 3064
rect 15932 2996 16000 3032
rect 15932 2964 15950 2996
rect 15982 2964 16000 2996
rect 15932 2928 16000 2964
rect 15932 2896 15950 2928
rect 15982 2896 16000 2928
rect 15932 2860 16000 2896
rect 15932 2828 15950 2860
rect 15982 2828 16000 2860
rect 15932 2792 16000 2828
rect 15932 2760 15950 2792
rect 15982 2760 16000 2792
rect 15932 2724 16000 2760
rect 15932 2692 15950 2724
rect 15982 2692 16000 2724
rect 15932 2656 16000 2692
rect 15932 2624 15950 2656
rect 15982 2624 16000 2656
rect 15932 2588 16000 2624
rect 15932 2556 15950 2588
rect 15982 2556 16000 2588
rect 15932 2520 16000 2556
rect 15932 2488 15950 2520
rect 15982 2488 16000 2520
rect 15932 2452 16000 2488
rect 15932 2420 15950 2452
rect 15982 2420 16000 2452
rect 15932 2384 16000 2420
rect 15932 2352 15950 2384
rect 15982 2352 16000 2384
rect 15932 2316 16000 2352
rect 15932 2284 15950 2316
rect 15982 2284 16000 2316
rect 15932 2248 16000 2284
rect 15932 2216 15950 2248
rect 15982 2216 16000 2248
rect 15932 2180 16000 2216
rect 15932 2148 15950 2180
rect 15982 2148 16000 2180
rect 15932 2112 16000 2148
rect 15932 2080 15950 2112
rect 15982 2080 16000 2112
rect 15932 2044 16000 2080
rect 15932 2012 15950 2044
rect 15982 2012 16000 2044
rect 15932 1976 16000 2012
rect 15932 1944 15950 1976
rect 15982 1944 16000 1976
rect 15932 1908 16000 1944
rect 15932 1876 15950 1908
rect 15982 1876 16000 1908
rect 15932 1840 16000 1876
rect 15932 1808 15950 1840
rect 15982 1808 16000 1840
rect 15932 1772 16000 1808
rect 15932 1740 15950 1772
rect 15982 1740 16000 1772
rect 15932 1704 16000 1740
rect 15932 1672 15950 1704
rect 15982 1672 16000 1704
rect 15932 1636 16000 1672
rect 15932 1604 15950 1636
rect 15982 1604 16000 1636
rect 15932 1568 16000 1604
rect 15932 1536 15950 1568
rect 15982 1536 16000 1568
rect 15932 1500 16000 1536
rect 15932 1468 15950 1500
rect 15982 1468 16000 1500
rect 15932 1432 16000 1468
rect 15932 1400 15950 1432
rect 15982 1400 16000 1432
rect 15932 1364 16000 1400
rect 15932 1332 15950 1364
rect 15982 1332 16000 1364
rect 15932 1296 16000 1332
rect 15932 1264 15950 1296
rect 15982 1264 16000 1296
rect 15932 1228 16000 1264
rect 15932 1196 15950 1228
rect 15982 1196 16000 1228
rect 15932 1160 16000 1196
rect 15932 1128 15950 1160
rect 15982 1128 16000 1160
rect 15932 1092 16000 1128
rect 15932 1060 15950 1092
rect 15982 1060 16000 1092
rect 15932 1024 16000 1060
rect 15932 992 15950 1024
rect 15982 992 16000 1024
rect 15932 956 16000 992
rect 15932 924 15950 956
rect 15982 924 16000 956
rect 15932 888 16000 924
rect 15932 856 15950 888
rect 15982 856 16000 888
rect 15932 820 16000 856
rect 15932 788 15950 820
rect 15982 788 16000 820
rect 15932 752 16000 788
rect 15932 720 15950 752
rect 15982 720 16000 752
rect 15932 684 16000 720
rect 15932 652 15950 684
rect 15982 652 16000 684
rect 15932 616 16000 652
rect 15932 584 15950 616
rect 15982 584 16000 616
rect 15932 548 16000 584
rect 15932 516 15950 548
rect 15982 516 16000 548
rect 15932 480 16000 516
rect 15932 448 15950 480
rect 15982 448 16000 480
rect 15932 412 16000 448
rect 15932 380 15950 412
rect 15982 380 16000 412
rect 0 312 18 344
rect 50 312 68 344
rect 0 276 68 312
rect 0 244 18 276
rect 50 244 68 276
rect 0 208 68 244
rect 0 176 18 208
rect 50 176 68 208
rect 0 140 68 176
rect 0 108 18 140
rect 50 108 68 140
rect 0 68 68 108
rect 15932 344 16000 380
rect 15932 312 15950 344
rect 15982 312 16000 344
rect 15932 276 16000 312
rect 15932 244 15950 276
rect 15982 244 16000 276
rect 15932 208 16000 244
rect 15932 176 15950 208
rect 15982 176 16000 208
rect 15932 140 16000 176
rect 15932 108 15950 140
rect 15982 108 16000 140
rect 15932 68 16000 108
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< nsubdiff >>
rect 360 3474 15640 3492
rect 360 3442 402 3474
rect 434 3442 470 3474
rect 502 3442 538 3474
rect 570 3442 606 3474
rect 638 3442 674 3474
rect 706 3442 742 3474
rect 774 3442 810 3474
rect 842 3442 878 3474
rect 910 3442 946 3474
rect 978 3442 1014 3474
rect 1046 3442 1082 3474
rect 1114 3442 1150 3474
rect 1182 3442 1218 3474
rect 1250 3442 1286 3474
rect 1318 3442 1354 3474
rect 1386 3442 1422 3474
rect 1454 3442 1490 3474
rect 1522 3442 1558 3474
rect 1590 3442 1626 3474
rect 1658 3442 1694 3474
rect 1726 3442 1762 3474
rect 1794 3442 1830 3474
rect 1862 3442 1898 3474
rect 1930 3442 1966 3474
rect 1998 3442 2034 3474
rect 2066 3442 2102 3474
rect 2134 3442 2170 3474
rect 2202 3442 2238 3474
rect 2270 3442 2306 3474
rect 2338 3442 2374 3474
rect 2406 3442 2442 3474
rect 2474 3442 2510 3474
rect 2542 3442 2578 3474
rect 2610 3442 2646 3474
rect 2678 3442 2714 3474
rect 2746 3442 2782 3474
rect 2814 3442 2850 3474
rect 2882 3442 2918 3474
rect 2950 3442 2986 3474
rect 3018 3442 3054 3474
rect 3086 3442 3122 3474
rect 3154 3442 3190 3474
rect 3222 3442 3258 3474
rect 3290 3442 3326 3474
rect 3358 3442 3394 3474
rect 3426 3442 3462 3474
rect 3494 3442 3530 3474
rect 3562 3442 3598 3474
rect 3630 3442 3666 3474
rect 3698 3442 3734 3474
rect 3766 3442 3802 3474
rect 3834 3442 3870 3474
rect 3902 3442 3938 3474
rect 3970 3442 4006 3474
rect 4038 3442 4074 3474
rect 4106 3442 4142 3474
rect 4174 3442 4210 3474
rect 4242 3442 4278 3474
rect 4310 3442 4346 3474
rect 4378 3442 4414 3474
rect 4446 3442 4482 3474
rect 4514 3442 4550 3474
rect 4582 3442 4618 3474
rect 4650 3442 4686 3474
rect 4718 3442 4754 3474
rect 4786 3442 4822 3474
rect 4854 3442 4890 3474
rect 4922 3442 4958 3474
rect 4990 3442 5026 3474
rect 5058 3442 5094 3474
rect 5126 3442 5162 3474
rect 5194 3442 5230 3474
rect 5262 3442 5298 3474
rect 5330 3442 5366 3474
rect 5398 3442 5434 3474
rect 5466 3442 5502 3474
rect 5534 3442 5570 3474
rect 5602 3442 5638 3474
rect 5670 3442 5706 3474
rect 5738 3442 5774 3474
rect 5806 3442 5842 3474
rect 5874 3442 5910 3474
rect 5942 3442 5978 3474
rect 6010 3442 6046 3474
rect 6078 3442 6114 3474
rect 6146 3442 6182 3474
rect 6214 3442 6250 3474
rect 6282 3442 6318 3474
rect 6350 3442 6386 3474
rect 6418 3442 6454 3474
rect 6486 3442 6522 3474
rect 6554 3442 6590 3474
rect 6622 3442 6658 3474
rect 6690 3442 6726 3474
rect 6758 3442 6794 3474
rect 6826 3442 6862 3474
rect 6894 3442 6930 3474
rect 6962 3442 6998 3474
rect 7030 3442 7066 3474
rect 7098 3442 7134 3474
rect 7166 3442 7202 3474
rect 7234 3442 7270 3474
rect 7302 3442 7338 3474
rect 7370 3442 7406 3474
rect 7438 3442 7474 3474
rect 7506 3442 7542 3474
rect 7574 3442 7610 3474
rect 7642 3442 7678 3474
rect 7710 3442 7746 3474
rect 7778 3442 7814 3474
rect 7846 3442 7882 3474
rect 7914 3442 7950 3474
rect 7982 3442 8018 3474
rect 8050 3442 8086 3474
rect 8118 3442 8154 3474
rect 8186 3442 8222 3474
rect 8254 3442 8290 3474
rect 8322 3442 8358 3474
rect 8390 3442 8426 3474
rect 8458 3442 8494 3474
rect 8526 3442 8562 3474
rect 8594 3442 8630 3474
rect 8662 3442 8698 3474
rect 8730 3442 8766 3474
rect 8798 3442 8834 3474
rect 8866 3442 8902 3474
rect 8934 3442 8970 3474
rect 9002 3442 9038 3474
rect 9070 3442 9106 3474
rect 9138 3442 9174 3474
rect 9206 3442 9242 3474
rect 9274 3442 9310 3474
rect 9342 3442 9378 3474
rect 9410 3442 9446 3474
rect 9478 3442 9514 3474
rect 9546 3442 9582 3474
rect 9614 3442 9650 3474
rect 9682 3442 9718 3474
rect 9750 3442 9786 3474
rect 9818 3442 9854 3474
rect 9886 3442 9922 3474
rect 9954 3442 9990 3474
rect 10022 3442 10058 3474
rect 10090 3442 10126 3474
rect 10158 3442 10194 3474
rect 10226 3442 10262 3474
rect 10294 3442 10330 3474
rect 10362 3442 10398 3474
rect 10430 3442 10466 3474
rect 10498 3442 10534 3474
rect 10566 3442 10602 3474
rect 10634 3442 10670 3474
rect 10702 3442 10738 3474
rect 10770 3442 10806 3474
rect 10838 3442 10874 3474
rect 10906 3442 10942 3474
rect 10974 3442 11010 3474
rect 11042 3442 11078 3474
rect 11110 3442 11146 3474
rect 11178 3442 11214 3474
rect 11246 3442 11282 3474
rect 11314 3442 11350 3474
rect 11382 3442 11418 3474
rect 11450 3442 11486 3474
rect 11518 3442 11554 3474
rect 11586 3442 11622 3474
rect 11654 3442 11690 3474
rect 11722 3442 11758 3474
rect 11790 3442 11826 3474
rect 11858 3442 11894 3474
rect 11926 3442 11962 3474
rect 11994 3442 12030 3474
rect 12062 3442 12098 3474
rect 12130 3442 12166 3474
rect 12198 3442 12234 3474
rect 12266 3442 12302 3474
rect 12334 3442 12370 3474
rect 12402 3442 12438 3474
rect 12470 3442 12506 3474
rect 12538 3442 12574 3474
rect 12606 3442 12642 3474
rect 12674 3442 12710 3474
rect 12742 3442 12778 3474
rect 12810 3442 12846 3474
rect 12878 3442 12914 3474
rect 12946 3442 12982 3474
rect 13014 3442 13050 3474
rect 13082 3442 13118 3474
rect 13150 3442 13186 3474
rect 13218 3442 13254 3474
rect 13286 3442 13322 3474
rect 13354 3442 13390 3474
rect 13422 3442 13458 3474
rect 13490 3442 13526 3474
rect 13558 3442 13594 3474
rect 13626 3442 13662 3474
rect 13694 3442 13730 3474
rect 13762 3442 13798 3474
rect 13830 3442 13866 3474
rect 13898 3442 13934 3474
rect 13966 3442 14002 3474
rect 14034 3442 14070 3474
rect 14102 3442 14138 3474
rect 14170 3442 14206 3474
rect 14238 3442 14274 3474
rect 14306 3442 14342 3474
rect 14374 3442 14410 3474
rect 14442 3442 14478 3474
rect 14510 3442 14546 3474
rect 14578 3442 14614 3474
rect 14646 3442 14682 3474
rect 14714 3442 14750 3474
rect 14782 3442 14818 3474
rect 14850 3442 14886 3474
rect 14918 3442 14954 3474
rect 14986 3442 15022 3474
rect 15054 3442 15090 3474
rect 15122 3442 15158 3474
rect 15190 3442 15226 3474
rect 15258 3442 15294 3474
rect 15326 3442 15362 3474
rect 15394 3442 15430 3474
rect 15462 3442 15498 3474
rect 15530 3442 15566 3474
rect 15598 3442 15640 3474
rect 360 3424 15640 3442
rect 360 3370 428 3424
rect 360 3338 378 3370
rect 410 3338 428 3370
rect 360 3302 428 3338
rect 15572 3370 15640 3424
rect 15572 3338 15590 3370
rect 15622 3338 15640 3370
rect 15572 3302 15640 3338
rect 360 3270 378 3302
rect 410 3270 428 3302
rect 360 3234 428 3270
rect 360 3202 378 3234
rect 410 3202 428 3234
rect 360 3166 428 3202
rect 360 3134 378 3166
rect 410 3134 428 3166
rect 360 3098 428 3134
rect 360 3066 378 3098
rect 410 3066 428 3098
rect 360 3030 428 3066
rect 360 2998 378 3030
rect 410 2998 428 3030
rect 360 2962 428 2998
rect 360 2930 378 2962
rect 410 2930 428 2962
rect 360 2894 428 2930
rect 360 2862 378 2894
rect 410 2862 428 2894
rect 360 2826 428 2862
rect 360 2794 378 2826
rect 410 2794 428 2826
rect 360 2758 428 2794
rect 360 2726 378 2758
rect 410 2726 428 2758
rect 360 2690 428 2726
rect 360 2658 378 2690
rect 410 2658 428 2690
rect 360 2622 428 2658
rect 360 2590 378 2622
rect 410 2590 428 2622
rect 360 2554 428 2590
rect 360 2522 378 2554
rect 410 2522 428 2554
rect 360 2486 428 2522
rect 360 2454 378 2486
rect 410 2454 428 2486
rect 360 2418 428 2454
rect 360 2386 378 2418
rect 410 2386 428 2418
rect 360 2350 428 2386
rect 360 2318 378 2350
rect 410 2318 428 2350
rect 360 2282 428 2318
rect 360 2250 378 2282
rect 410 2250 428 2282
rect 360 2214 428 2250
rect 360 2182 378 2214
rect 410 2182 428 2214
rect 360 2146 428 2182
rect 360 2114 378 2146
rect 410 2114 428 2146
rect 360 2078 428 2114
rect 360 2046 378 2078
rect 410 2046 428 2078
rect 360 2010 428 2046
rect 360 1978 378 2010
rect 410 1978 428 2010
rect 360 1942 428 1978
rect 15572 3270 15590 3302
rect 15622 3270 15640 3302
rect 15572 3234 15640 3270
rect 15572 3202 15590 3234
rect 15622 3202 15640 3234
rect 15572 3166 15640 3202
rect 15572 3134 15590 3166
rect 15622 3134 15640 3166
rect 15572 3098 15640 3134
rect 15572 3066 15590 3098
rect 15622 3066 15640 3098
rect 15572 3030 15640 3066
rect 15572 2998 15590 3030
rect 15622 2998 15640 3030
rect 15572 2962 15640 2998
rect 15572 2930 15590 2962
rect 15622 2930 15640 2962
rect 15572 2894 15640 2930
rect 15572 2862 15590 2894
rect 15622 2862 15640 2894
rect 15572 2826 15640 2862
rect 15572 2794 15590 2826
rect 15622 2794 15640 2826
rect 15572 2758 15640 2794
rect 15572 2726 15590 2758
rect 15622 2726 15640 2758
rect 15572 2690 15640 2726
rect 15572 2658 15590 2690
rect 15622 2658 15640 2690
rect 15572 2622 15640 2658
rect 15572 2590 15590 2622
rect 15622 2590 15640 2622
rect 15572 2554 15640 2590
rect 15572 2522 15590 2554
rect 15622 2522 15640 2554
rect 15572 2486 15640 2522
rect 15572 2454 15590 2486
rect 15622 2454 15640 2486
rect 15572 2418 15640 2454
rect 15572 2386 15590 2418
rect 15622 2386 15640 2418
rect 15572 2350 15640 2386
rect 15572 2318 15590 2350
rect 15622 2318 15640 2350
rect 15572 2282 15640 2318
rect 15572 2250 15590 2282
rect 15622 2250 15640 2282
rect 15572 2214 15640 2250
rect 15572 2182 15590 2214
rect 15622 2182 15640 2214
rect 15572 2146 15640 2182
rect 15572 2114 15590 2146
rect 15622 2114 15640 2146
rect 15572 2078 15640 2114
rect 15572 2046 15590 2078
rect 15622 2046 15640 2078
rect 15572 2010 15640 2046
rect 15572 1978 15590 2010
rect 15622 1978 15640 2010
rect 360 1910 378 1942
rect 410 1910 428 1942
rect 360 1874 428 1910
rect 15572 1942 15640 1978
rect 15572 1910 15590 1942
rect 15622 1910 15640 1942
rect 360 1842 378 1874
rect 410 1842 428 1874
rect 360 1806 428 1842
rect 360 1774 378 1806
rect 410 1774 428 1806
rect 360 1738 428 1774
rect 360 1706 378 1738
rect 410 1706 428 1738
rect 360 1670 428 1706
rect 360 1638 378 1670
rect 410 1638 428 1670
rect 360 1602 428 1638
rect 360 1570 378 1602
rect 410 1570 428 1602
rect 360 1534 428 1570
rect 360 1502 378 1534
rect 410 1502 428 1534
rect 360 1466 428 1502
rect 360 1434 378 1466
rect 410 1434 428 1466
rect 360 1398 428 1434
rect 360 1366 378 1398
rect 410 1366 428 1398
rect 360 1330 428 1366
rect 360 1298 378 1330
rect 410 1298 428 1330
rect 360 1262 428 1298
rect 360 1230 378 1262
rect 410 1230 428 1262
rect 360 1194 428 1230
rect 360 1162 378 1194
rect 410 1162 428 1194
rect 360 1126 428 1162
rect 360 1094 378 1126
rect 410 1094 428 1126
rect 360 1058 428 1094
rect 360 1026 378 1058
rect 410 1026 428 1058
rect 360 990 428 1026
rect 360 958 378 990
rect 410 958 428 990
rect 360 922 428 958
rect 360 890 378 922
rect 410 890 428 922
rect 360 854 428 890
rect 360 822 378 854
rect 410 822 428 854
rect 360 786 428 822
rect 360 754 378 786
rect 410 754 428 786
rect 360 718 428 754
rect 360 686 378 718
rect 410 686 428 718
rect 360 650 428 686
rect 360 618 378 650
rect 410 618 428 650
rect 360 582 428 618
rect 360 550 378 582
rect 410 550 428 582
rect 15572 1874 15640 1910
rect 15572 1842 15590 1874
rect 15622 1842 15640 1874
rect 15572 1806 15640 1842
rect 15572 1774 15590 1806
rect 15622 1774 15640 1806
rect 15572 1738 15640 1774
rect 15572 1706 15590 1738
rect 15622 1706 15640 1738
rect 15572 1670 15640 1706
rect 15572 1638 15590 1670
rect 15622 1638 15640 1670
rect 15572 1602 15640 1638
rect 15572 1570 15590 1602
rect 15622 1570 15640 1602
rect 15572 1534 15640 1570
rect 15572 1502 15590 1534
rect 15622 1502 15640 1534
rect 15572 1466 15640 1502
rect 15572 1434 15590 1466
rect 15622 1434 15640 1466
rect 15572 1398 15640 1434
rect 15572 1366 15590 1398
rect 15622 1366 15640 1398
rect 15572 1330 15640 1366
rect 15572 1298 15590 1330
rect 15622 1298 15640 1330
rect 15572 1262 15640 1298
rect 15572 1230 15590 1262
rect 15622 1230 15640 1262
rect 15572 1194 15640 1230
rect 15572 1162 15590 1194
rect 15622 1162 15640 1194
rect 15572 1126 15640 1162
rect 15572 1094 15590 1126
rect 15622 1094 15640 1126
rect 15572 1058 15640 1094
rect 15572 1026 15590 1058
rect 15622 1026 15640 1058
rect 15572 990 15640 1026
rect 15572 958 15590 990
rect 15622 958 15640 990
rect 15572 922 15640 958
rect 15572 890 15590 922
rect 15622 890 15640 922
rect 15572 854 15640 890
rect 15572 822 15590 854
rect 15622 822 15640 854
rect 15572 786 15640 822
rect 15572 754 15590 786
rect 15622 754 15640 786
rect 15572 718 15640 754
rect 15572 686 15590 718
rect 15622 686 15640 718
rect 15572 650 15640 686
rect 15572 618 15590 650
rect 15622 618 15640 650
rect 15572 582 15640 618
rect 15572 550 15590 582
rect 15622 550 15640 582
rect 360 514 428 550
rect 360 482 378 514
rect 410 482 428 514
rect 360 428 428 482
rect 15572 514 15640 550
rect 15572 482 15590 514
rect 15622 482 15640 514
rect 15572 428 15640 482
rect 360 410 15640 428
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6794 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7406 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 7982 378 8018 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8594 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9206 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 360 15640 378
<< psubdiffcont >>
rect 28 3802 60 3834
rect 96 3802 128 3834
rect 164 3802 196 3834
rect 232 3802 264 3834
rect 300 3802 332 3834
rect 368 3802 400 3834
rect 436 3802 468 3834
rect 504 3802 536 3834
rect 572 3802 604 3834
rect 640 3802 672 3834
rect 708 3802 740 3834
rect 776 3802 808 3834
rect 844 3802 876 3834
rect 912 3802 944 3834
rect 980 3802 1012 3834
rect 1048 3802 1080 3834
rect 1116 3802 1148 3834
rect 1184 3802 1216 3834
rect 1252 3802 1284 3834
rect 1320 3802 1352 3834
rect 1388 3802 1420 3834
rect 1456 3802 1488 3834
rect 1524 3802 1556 3834
rect 1592 3802 1624 3834
rect 1660 3802 1692 3834
rect 1728 3802 1760 3834
rect 1796 3802 1828 3834
rect 1864 3802 1896 3834
rect 1932 3802 1964 3834
rect 2000 3802 2032 3834
rect 2068 3802 2100 3834
rect 2136 3802 2168 3834
rect 2204 3802 2236 3834
rect 2272 3802 2304 3834
rect 2340 3802 2372 3834
rect 2408 3802 2440 3834
rect 2476 3802 2508 3834
rect 2544 3802 2576 3834
rect 2612 3802 2644 3834
rect 2680 3802 2712 3834
rect 2748 3802 2780 3834
rect 2816 3802 2848 3834
rect 2884 3802 2916 3834
rect 2952 3802 2984 3834
rect 3020 3802 3052 3834
rect 3088 3802 3120 3834
rect 3156 3802 3188 3834
rect 3224 3802 3256 3834
rect 3292 3802 3324 3834
rect 3360 3802 3392 3834
rect 3428 3802 3460 3834
rect 3496 3802 3528 3834
rect 3564 3802 3596 3834
rect 3632 3802 3664 3834
rect 3700 3802 3732 3834
rect 3768 3802 3800 3834
rect 3836 3802 3868 3834
rect 3904 3802 3936 3834
rect 3972 3802 4004 3834
rect 4040 3802 4072 3834
rect 4108 3802 4140 3834
rect 4176 3802 4208 3834
rect 4244 3802 4276 3834
rect 4312 3802 4344 3834
rect 4380 3802 4412 3834
rect 4448 3802 4480 3834
rect 4516 3802 4548 3834
rect 4584 3802 4616 3834
rect 4652 3802 4684 3834
rect 4720 3802 4752 3834
rect 4788 3802 4820 3834
rect 4856 3802 4888 3834
rect 4924 3802 4956 3834
rect 4992 3802 5024 3834
rect 5060 3802 5092 3834
rect 5128 3802 5160 3834
rect 5196 3802 5228 3834
rect 5264 3802 5296 3834
rect 5332 3802 5364 3834
rect 5400 3802 5432 3834
rect 5468 3802 5500 3834
rect 5536 3802 5568 3834
rect 5604 3802 5636 3834
rect 5672 3802 5704 3834
rect 5740 3802 5772 3834
rect 5808 3802 5840 3834
rect 5876 3802 5908 3834
rect 5944 3802 5976 3834
rect 6012 3802 6044 3834
rect 6080 3802 6112 3834
rect 6148 3802 6180 3834
rect 6216 3802 6248 3834
rect 6284 3802 6316 3834
rect 6352 3802 6384 3834
rect 6420 3802 6452 3834
rect 6488 3802 6520 3834
rect 6556 3802 6588 3834
rect 6624 3802 6656 3834
rect 6692 3802 6724 3834
rect 6760 3802 6792 3834
rect 6828 3802 6860 3834
rect 6896 3802 6928 3834
rect 6964 3802 6996 3834
rect 7032 3802 7064 3834
rect 7100 3802 7132 3834
rect 7168 3802 7200 3834
rect 7236 3802 7268 3834
rect 7304 3802 7336 3834
rect 7372 3802 7404 3834
rect 7440 3802 7472 3834
rect 7508 3802 7540 3834
rect 7576 3802 7608 3834
rect 7644 3802 7676 3834
rect 7712 3802 7744 3834
rect 7780 3802 7812 3834
rect 7848 3802 7880 3834
rect 7916 3802 7948 3834
rect 7984 3802 8016 3834
rect 8052 3802 8084 3834
rect 8120 3802 8152 3834
rect 8188 3802 8220 3834
rect 8256 3802 8288 3834
rect 8324 3802 8356 3834
rect 8392 3802 8424 3834
rect 8460 3802 8492 3834
rect 8528 3802 8560 3834
rect 8596 3802 8628 3834
rect 8664 3802 8696 3834
rect 8732 3802 8764 3834
rect 8800 3802 8832 3834
rect 8868 3802 8900 3834
rect 8936 3802 8968 3834
rect 9004 3802 9036 3834
rect 9072 3802 9104 3834
rect 9140 3802 9172 3834
rect 9208 3802 9240 3834
rect 9276 3802 9308 3834
rect 9344 3802 9376 3834
rect 9412 3802 9444 3834
rect 9480 3802 9512 3834
rect 9548 3802 9580 3834
rect 9616 3802 9648 3834
rect 9684 3802 9716 3834
rect 9752 3802 9784 3834
rect 9820 3802 9852 3834
rect 9888 3802 9920 3834
rect 9956 3802 9988 3834
rect 10024 3802 10056 3834
rect 10092 3802 10124 3834
rect 10160 3802 10192 3834
rect 10228 3802 10260 3834
rect 10296 3802 10328 3834
rect 10364 3802 10396 3834
rect 10432 3802 10464 3834
rect 10500 3802 10532 3834
rect 10568 3802 10600 3834
rect 10636 3802 10668 3834
rect 10704 3802 10736 3834
rect 10772 3802 10804 3834
rect 10840 3802 10872 3834
rect 10908 3802 10940 3834
rect 10976 3802 11008 3834
rect 11044 3802 11076 3834
rect 11112 3802 11144 3834
rect 11180 3802 11212 3834
rect 11248 3802 11280 3834
rect 11316 3802 11348 3834
rect 11384 3802 11416 3834
rect 11452 3802 11484 3834
rect 11520 3802 11552 3834
rect 11588 3802 11620 3834
rect 11656 3802 11688 3834
rect 11724 3802 11756 3834
rect 11792 3802 11824 3834
rect 11860 3802 11892 3834
rect 11928 3802 11960 3834
rect 11996 3802 12028 3834
rect 12064 3802 12096 3834
rect 12132 3802 12164 3834
rect 12200 3802 12232 3834
rect 12268 3802 12300 3834
rect 12336 3802 12368 3834
rect 12404 3802 12436 3834
rect 12472 3802 12504 3834
rect 12540 3802 12572 3834
rect 12608 3802 12640 3834
rect 12676 3802 12708 3834
rect 12744 3802 12776 3834
rect 12812 3802 12844 3834
rect 12880 3802 12912 3834
rect 12948 3802 12980 3834
rect 13016 3802 13048 3834
rect 13084 3802 13116 3834
rect 13152 3802 13184 3834
rect 13220 3802 13252 3834
rect 13288 3802 13320 3834
rect 13356 3802 13388 3834
rect 13424 3802 13456 3834
rect 13492 3802 13524 3834
rect 13560 3802 13592 3834
rect 13628 3802 13660 3834
rect 13696 3802 13728 3834
rect 13764 3802 13796 3834
rect 13832 3802 13864 3834
rect 13900 3802 13932 3834
rect 13968 3802 14000 3834
rect 14036 3802 14068 3834
rect 14104 3802 14136 3834
rect 14172 3802 14204 3834
rect 14240 3802 14272 3834
rect 14308 3802 14340 3834
rect 14376 3802 14408 3834
rect 14444 3802 14476 3834
rect 14512 3802 14544 3834
rect 14580 3802 14612 3834
rect 14648 3802 14680 3834
rect 14716 3802 14748 3834
rect 14784 3802 14816 3834
rect 14852 3802 14884 3834
rect 14920 3802 14952 3834
rect 14988 3802 15020 3834
rect 15056 3802 15088 3834
rect 15124 3802 15156 3834
rect 15192 3802 15224 3834
rect 15260 3802 15292 3834
rect 15328 3802 15360 3834
rect 15396 3802 15428 3834
rect 15464 3802 15496 3834
rect 15532 3802 15564 3834
rect 15600 3802 15632 3834
rect 15668 3802 15700 3834
rect 15736 3802 15768 3834
rect 15804 3802 15836 3834
rect 15872 3802 15904 3834
rect 15940 3802 15972 3834
rect 18 3712 50 3744
rect 18 3644 50 3676
rect 18 3576 50 3608
rect 18 3508 50 3540
rect 15950 3712 15982 3744
rect 15950 3644 15982 3676
rect 15950 3576 15982 3608
rect 15950 3508 15982 3540
rect 18 3440 50 3472
rect 18 3372 50 3404
rect 18 3304 50 3336
rect 18 3236 50 3268
rect 18 3168 50 3200
rect 18 3100 50 3132
rect 18 3032 50 3064
rect 18 2964 50 2996
rect 18 2896 50 2928
rect 18 2828 50 2860
rect 18 2760 50 2792
rect 18 2692 50 2724
rect 18 2624 50 2656
rect 18 2556 50 2588
rect 18 2488 50 2520
rect 18 2420 50 2452
rect 18 2352 50 2384
rect 18 2284 50 2316
rect 18 2216 50 2248
rect 18 2148 50 2180
rect 18 2080 50 2112
rect 18 2012 50 2044
rect 18 1944 50 1976
rect 18 1876 50 1908
rect 18 1808 50 1840
rect 18 1740 50 1772
rect 18 1672 50 1704
rect 18 1604 50 1636
rect 18 1536 50 1568
rect 18 1468 50 1500
rect 18 1400 50 1432
rect 18 1332 50 1364
rect 18 1264 50 1296
rect 18 1196 50 1228
rect 18 1128 50 1160
rect 18 1060 50 1092
rect 18 992 50 1024
rect 18 924 50 956
rect 18 856 50 888
rect 18 788 50 820
rect 18 720 50 752
rect 18 652 50 684
rect 18 584 50 616
rect 18 516 50 548
rect 18 448 50 480
rect 18 380 50 412
rect 15950 3440 15982 3472
rect 15950 3372 15982 3404
rect 15950 3304 15982 3336
rect 15950 3236 15982 3268
rect 15950 3168 15982 3200
rect 15950 3100 15982 3132
rect 15950 3032 15982 3064
rect 15950 2964 15982 2996
rect 15950 2896 15982 2928
rect 15950 2828 15982 2860
rect 15950 2760 15982 2792
rect 15950 2692 15982 2724
rect 15950 2624 15982 2656
rect 15950 2556 15982 2588
rect 15950 2488 15982 2520
rect 15950 2420 15982 2452
rect 15950 2352 15982 2384
rect 15950 2284 15982 2316
rect 15950 2216 15982 2248
rect 15950 2148 15982 2180
rect 15950 2080 15982 2112
rect 15950 2012 15982 2044
rect 15950 1944 15982 1976
rect 15950 1876 15982 1908
rect 15950 1808 15982 1840
rect 15950 1740 15982 1772
rect 15950 1672 15982 1704
rect 15950 1604 15982 1636
rect 15950 1536 15982 1568
rect 15950 1468 15982 1500
rect 15950 1400 15982 1432
rect 15950 1332 15982 1364
rect 15950 1264 15982 1296
rect 15950 1196 15982 1228
rect 15950 1128 15982 1160
rect 15950 1060 15982 1092
rect 15950 992 15982 1024
rect 15950 924 15982 956
rect 15950 856 15982 888
rect 15950 788 15982 820
rect 15950 720 15982 752
rect 15950 652 15982 684
rect 15950 584 15982 616
rect 15950 516 15982 548
rect 15950 448 15982 480
rect 15950 380 15982 412
rect 18 312 50 344
rect 18 244 50 276
rect 18 176 50 208
rect 18 108 50 140
rect 15950 312 15982 344
rect 15950 244 15982 276
rect 15950 176 15982 208
rect 15950 108 15982 140
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< nsubdiffcont >>
rect 402 3442 434 3474
rect 470 3442 502 3474
rect 538 3442 570 3474
rect 606 3442 638 3474
rect 674 3442 706 3474
rect 742 3442 774 3474
rect 810 3442 842 3474
rect 878 3442 910 3474
rect 946 3442 978 3474
rect 1014 3442 1046 3474
rect 1082 3442 1114 3474
rect 1150 3442 1182 3474
rect 1218 3442 1250 3474
rect 1286 3442 1318 3474
rect 1354 3442 1386 3474
rect 1422 3442 1454 3474
rect 1490 3442 1522 3474
rect 1558 3442 1590 3474
rect 1626 3442 1658 3474
rect 1694 3442 1726 3474
rect 1762 3442 1794 3474
rect 1830 3442 1862 3474
rect 1898 3442 1930 3474
rect 1966 3442 1998 3474
rect 2034 3442 2066 3474
rect 2102 3442 2134 3474
rect 2170 3442 2202 3474
rect 2238 3442 2270 3474
rect 2306 3442 2338 3474
rect 2374 3442 2406 3474
rect 2442 3442 2474 3474
rect 2510 3442 2542 3474
rect 2578 3442 2610 3474
rect 2646 3442 2678 3474
rect 2714 3442 2746 3474
rect 2782 3442 2814 3474
rect 2850 3442 2882 3474
rect 2918 3442 2950 3474
rect 2986 3442 3018 3474
rect 3054 3442 3086 3474
rect 3122 3442 3154 3474
rect 3190 3442 3222 3474
rect 3258 3442 3290 3474
rect 3326 3442 3358 3474
rect 3394 3442 3426 3474
rect 3462 3442 3494 3474
rect 3530 3442 3562 3474
rect 3598 3442 3630 3474
rect 3666 3442 3698 3474
rect 3734 3442 3766 3474
rect 3802 3442 3834 3474
rect 3870 3442 3902 3474
rect 3938 3442 3970 3474
rect 4006 3442 4038 3474
rect 4074 3442 4106 3474
rect 4142 3442 4174 3474
rect 4210 3442 4242 3474
rect 4278 3442 4310 3474
rect 4346 3442 4378 3474
rect 4414 3442 4446 3474
rect 4482 3442 4514 3474
rect 4550 3442 4582 3474
rect 4618 3442 4650 3474
rect 4686 3442 4718 3474
rect 4754 3442 4786 3474
rect 4822 3442 4854 3474
rect 4890 3442 4922 3474
rect 4958 3442 4990 3474
rect 5026 3442 5058 3474
rect 5094 3442 5126 3474
rect 5162 3442 5194 3474
rect 5230 3442 5262 3474
rect 5298 3442 5330 3474
rect 5366 3442 5398 3474
rect 5434 3442 5466 3474
rect 5502 3442 5534 3474
rect 5570 3442 5602 3474
rect 5638 3442 5670 3474
rect 5706 3442 5738 3474
rect 5774 3442 5806 3474
rect 5842 3442 5874 3474
rect 5910 3442 5942 3474
rect 5978 3442 6010 3474
rect 6046 3442 6078 3474
rect 6114 3442 6146 3474
rect 6182 3442 6214 3474
rect 6250 3442 6282 3474
rect 6318 3442 6350 3474
rect 6386 3442 6418 3474
rect 6454 3442 6486 3474
rect 6522 3442 6554 3474
rect 6590 3442 6622 3474
rect 6658 3442 6690 3474
rect 6726 3442 6758 3474
rect 6794 3442 6826 3474
rect 6862 3442 6894 3474
rect 6930 3442 6962 3474
rect 6998 3442 7030 3474
rect 7066 3442 7098 3474
rect 7134 3442 7166 3474
rect 7202 3442 7234 3474
rect 7270 3442 7302 3474
rect 7338 3442 7370 3474
rect 7406 3442 7438 3474
rect 7474 3442 7506 3474
rect 7542 3442 7574 3474
rect 7610 3442 7642 3474
rect 7678 3442 7710 3474
rect 7746 3442 7778 3474
rect 7814 3442 7846 3474
rect 7882 3442 7914 3474
rect 7950 3442 7982 3474
rect 8018 3442 8050 3474
rect 8086 3442 8118 3474
rect 8154 3442 8186 3474
rect 8222 3442 8254 3474
rect 8290 3442 8322 3474
rect 8358 3442 8390 3474
rect 8426 3442 8458 3474
rect 8494 3442 8526 3474
rect 8562 3442 8594 3474
rect 8630 3442 8662 3474
rect 8698 3442 8730 3474
rect 8766 3442 8798 3474
rect 8834 3442 8866 3474
rect 8902 3442 8934 3474
rect 8970 3442 9002 3474
rect 9038 3442 9070 3474
rect 9106 3442 9138 3474
rect 9174 3442 9206 3474
rect 9242 3442 9274 3474
rect 9310 3442 9342 3474
rect 9378 3442 9410 3474
rect 9446 3442 9478 3474
rect 9514 3442 9546 3474
rect 9582 3442 9614 3474
rect 9650 3442 9682 3474
rect 9718 3442 9750 3474
rect 9786 3442 9818 3474
rect 9854 3442 9886 3474
rect 9922 3442 9954 3474
rect 9990 3442 10022 3474
rect 10058 3442 10090 3474
rect 10126 3442 10158 3474
rect 10194 3442 10226 3474
rect 10262 3442 10294 3474
rect 10330 3442 10362 3474
rect 10398 3442 10430 3474
rect 10466 3442 10498 3474
rect 10534 3442 10566 3474
rect 10602 3442 10634 3474
rect 10670 3442 10702 3474
rect 10738 3442 10770 3474
rect 10806 3442 10838 3474
rect 10874 3442 10906 3474
rect 10942 3442 10974 3474
rect 11010 3442 11042 3474
rect 11078 3442 11110 3474
rect 11146 3442 11178 3474
rect 11214 3442 11246 3474
rect 11282 3442 11314 3474
rect 11350 3442 11382 3474
rect 11418 3442 11450 3474
rect 11486 3442 11518 3474
rect 11554 3442 11586 3474
rect 11622 3442 11654 3474
rect 11690 3442 11722 3474
rect 11758 3442 11790 3474
rect 11826 3442 11858 3474
rect 11894 3442 11926 3474
rect 11962 3442 11994 3474
rect 12030 3442 12062 3474
rect 12098 3442 12130 3474
rect 12166 3442 12198 3474
rect 12234 3442 12266 3474
rect 12302 3442 12334 3474
rect 12370 3442 12402 3474
rect 12438 3442 12470 3474
rect 12506 3442 12538 3474
rect 12574 3442 12606 3474
rect 12642 3442 12674 3474
rect 12710 3442 12742 3474
rect 12778 3442 12810 3474
rect 12846 3442 12878 3474
rect 12914 3442 12946 3474
rect 12982 3442 13014 3474
rect 13050 3442 13082 3474
rect 13118 3442 13150 3474
rect 13186 3442 13218 3474
rect 13254 3442 13286 3474
rect 13322 3442 13354 3474
rect 13390 3442 13422 3474
rect 13458 3442 13490 3474
rect 13526 3442 13558 3474
rect 13594 3442 13626 3474
rect 13662 3442 13694 3474
rect 13730 3442 13762 3474
rect 13798 3442 13830 3474
rect 13866 3442 13898 3474
rect 13934 3442 13966 3474
rect 14002 3442 14034 3474
rect 14070 3442 14102 3474
rect 14138 3442 14170 3474
rect 14206 3442 14238 3474
rect 14274 3442 14306 3474
rect 14342 3442 14374 3474
rect 14410 3442 14442 3474
rect 14478 3442 14510 3474
rect 14546 3442 14578 3474
rect 14614 3442 14646 3474
rect 14682 3442 14714 3474
rect 14750 3442 14782 3474
rect 14818 3442 14850 3474
rect 14886 3442 14918 3474
rect 14954 3442 14986 3474
rect 15022 3442 15054 3474
rect 15090 3442 15122 3474
rect 15158 3442 15190 3474
rect 15226 3442 15258 3474
rect 15294 3442 15326 3474
rect 15362 3442 15394 3474
rect 15430 3442 15462 3474
rect 15498 3442 15530 3474
rect 15566 3442 15598 3474
rect 378 3338 410 3370
rect 15590 3338 15622 3370
rect 378 3270 410 3302
rect 378 3202 410 3234
rect 378 3134 410 3166
rect 378 3066 410 3098
rect 378 2998 410 3030
rect 378 2930 410 2962
rect 378 2862 410 2894
rect 378 2794 410 2826
rect 378 2726 410 2758
rect 378 2658 410 2690
rect 378 2590 410 2622
rect 378 2522 410 2554
rect 378 2454 410 2486
rect 378 2386 410 2418
rect 378 2318 410 2350
rect 378 2250 410 2282
rect 378 2182 410 2214
rect 378 2114 410 2146
rect 378 2046 410 2078
rect 378 1978 410 2010
rect 15590 3270 15622 3302
rect 15590 3202 15622 3234
rect 15590 3134 15622 3166
rect 15590 3066 15622 3098
rect 15590 2998 15622 3030
rect 15590 2930 15622 2962
rect 15590 2862 15622 2894
rect 15590 2794 15622 2826
rect 15590 2726 15622 2758
rect 15590 2658 15622 2690
rect 15590 2590 15622 2622
rect 15590 2522 15622 2554
rect 15590 2454 15622 2486
rect 15590 2386 15622 2418
rect 15590 2318 15622 2350
rect 15590 2250 15622 2282
rect 15590 2182 15622 2214
rect 15590 2114 15622 2146
rect 15590 2046 15622 2078
rect 15590 1978 15622 2010
rect 378 1910 410 1942
rect 15590 1910 15622 1942
rect 378 1842 410 1874
rect 378 1774 410 1806
rect 378 1706 410 1738
rect 378 1638 410 1670
rect 378 1570 410 1602
rect 378 1502 410 1534
rect 378 1434 410 1466
rect 378 1366 410 1398
rect 378 1298 410 1330
rect 378 1230 410 1262
rect 378 1162 410 1194
rect 378 1094 410 1126
rect 378 1026 410 1058
rect 378 958 410 990
rect 378 890 410 922
rect 378 822 410 854
rect 378 754 410 786
rect 378 686 410 718
rect 378 618 410 650
rect 378 550 410 582
rect 15590 1842 15622 1874
rect 15590 1774 15622 1806
rect 15590 1706 15622 1738
rect 15590 1638 15622 1670
rect 15590 1570 15622 1602
rect 15590 1502 15622 1534
rect 15590 1434 15622 1466
rect 15590 1366 15622 1398
rect 15590 1298 15622 1330
rect 15590 1230 15622 1262
rect 15590 1162 15622 1194
rect 15590 1094 15622 1126
rect 15590 1026 15622 1058
rect 15590 958 15622 990
rect 15590 890 15622 922
rect 15590 822 15622 854
rect 15590 754 15622 786
rect 15590 686 15622 718
rect 15590 618 15622 650
rect 15590 550 15622 582
rect 378 482 410 514
rect 15590 482 15622 514
rect 402 378 434 410
rect 470 378 502 410
rect 538 378 570 410
rect 606 378 638 410
rect 674 378 706 410
rect 742 378 774 410
rect 810 378 842 410
rect 878 378 910 410
rect 946 378 978 410
rect 1014 378 1046 410
rect 1082 378 1114 410
rect 1150 378 1182 410
rect 1218 378 1250 410
rect 1286 378 1318 410
rect 1354 378 1386 410
rect 1422 378 1454 410
rect 1490 378 1522 410
rect 1558 378 1590 410
rect 1626 378 1658 410
rect 1694 378 1726 410
rect 1762 378 1794 410
rect 1830 378 1862 410
rect 1898 378 1930 410
rect 1966 378 1998 410
rect 2034 378 2066 410
rect 2102 378 2134 410
rect 2170 378 2202 410
rect 2238 378 2270 410
rect 2306 378 2338 410
rect 2374 378 2406 410
rect 2442 378 2474 410
rect 2510 378 2542 410
rect 2578 378 2610 410
rect 2646 378 2678 410
rect 2714 378 2746 410
rect 2782 378 2814 410
rect 2850 378 2882 410
rect 2918 378 2950 410
rect 2986 378 3018 410
rect 3054 378 3086 410
rect 3122 378 3154 410
rect 3190 378 3222 410
rect 3258 378 3290 410
rect 3326 378 3358 410
rect 3394 378 3426 410
rect 3462 378 3494 410
rect 3530 378 3562 410
rect 3598 378 3630 410
rect 3666 378 3698 410
rect 3734 378 3766 410
rect 3802 378 3834 410
rect 3870 378 3902 410
rect 3938 378 3970 410
rect 4006 378 4038 410
rect 4074 378 4106 410
rect 4142 378 4174 410
rect 4210 378 4242 410
rect 4278 378 4310 410
rect 4346 378 4378 410
rect 4414 378 4446 410
rect 4482 378 4514 410
rect 4550 378 4582 410
rect 4618 378 4650 410
rect 4686 378 4718 410
rect 4754 378 4786 410
rect 4822 378 4854 410
rect 4890 378 4922 410
rect 4958 378 4990 410
rect 5026 378 5058 410
rect 5094 378 5126 410
rect 5162 378 5194 410
rect 5230 378 5262 410
rect 5298 378 5330 410
rect 5366 378 5398 410
rect 5434 378 5466 410
rect 5502 378 5534 410
rect 5570 378 5602 410
rect 5638 378 5670 410
rect 5706 378 5738 410
rect 5774 378 5806 410
rect 5842 378 5874 410
rect 5910 378 5942 410
rect 5978 378 6010 410
rect 6046 378 6078 410
rect 6114 378 6146 410
rect 6182 378 6214 410
rect 6250 378 6282 410
rect 6318 378 6350 410
rect 6386 378 6418 410
rect 6454 378 6486 410
rect 6522 378 6554 410
rect 6590 378 6622 410
rect 6658 378 6690 410
rect 6726 378 6758 410
rect 6794 378 6826 410
rect 6862 378 6894 410
rect 6930 378 6962 410
rect 6998 378 7030 410
rect 7066 378 7098 410
rect 7134 378 7166 410
rect 7202 378 7234 410
rect 7270 378 7302 410
rect 7338 378 7370 410
rect 7406 378 7438 410
rect 7474 378 7506 410
rect 7542 378 7574 410
rect 7610 378 7642 410
rect 7678 378 7710 410
rect 7746 378 7778 410
rect 7814 378 7846 410
rect 7882 378 7914 410
rect 7950 378 7982 410
rect 8018 378 8050 410
rect 8086 378 8118 410
rect 8154 378 8186 410
rect 8222 378 8254 410
rect 8290 378 8322 410
rect 8358 378 8390 410
rect 8426 378 8458 410
rect 8494 378 8526 410
rect 8562 378 8594 410
rect 8630 378 8662 410
rect 8698 378 8730 410
rect 8766 378 8798 410
rect 8834 378 8866 410
rect 8902 378 8934 410
rect 8970 378 9002 410
rect 9038 378 9070 410
rect 9106 378 9138 410
rect 9174 378 9206 410
rect 9242 378 9274 410
rect 9310 378 9342 410
rect 9378 378 9410 410
rect 9446 378 9478 410
rect 9514 378 9546 410
rect 9582 378 9614 410
rect 9650 378 9682 410
rect 9718 378 9750 410
rect 9786 378 9818 410
rect 9854 378 9886 410
rect 9922 378 9954 410
rect 9990 378 10022 410
rect 10058 378 10090 410
rect 10126 378 10158 410
rect 10194 378 10226 410
rect 10262 378 10294 410
rect 10330 378 10362 410
rect 10398 378 10430 410
rect 10466 378 10498 410
rect 10534 378 10566 410
rect 10602 378 10634 410
rect 10670 378 10702 410
rect 10738 378 10770 410
rect 10806 378 10838 410
rect 10874 378 10906 410
rect 10942 378 10974 410
rect 11010 378 11042 410
rect 11078 378 11110 410
rect 11146 378 11178 410
rect 11214 378 11246 410
rect 11282 378 11314 410
rect 11350 378 11382 410
rect 11418 378 11450 410
rect 11486 378 11518 410
rect 11554 378 11586 410
rect 11622 378 11654 410
rect 11690 378 11722 410
rect 11758 378 11790 410
rect 11826 378 11858 410
rect 11894 378 11926 410
rect 11962 378 11994 410
rect 12030 378 12062 410
rect 12098 378 12130 410
rect 12166 378 12198 410
rect 12234 378 12266 410
rect 12302 378 12334 410
rect 12370 378 12402 410
rect 12438 378 12470 410
rect 12506 378 12538 410
rect 12574 378 12606 410
rect 12642 378 12674 410
rect 12710 378 12742 410
rect 12778 378 12810 410
rect 12846 378 12878 410
rect 12914 378 12946 410
rect 12982 378 13014 410
rect 13050 378 13082 410
rect 13118 378 13150 410
rect 13186 378 13218 410
rect 13254 378 13286 410
rect 13322 378 13354 410
rect 13390 378 13422 410
rect 13458 378 13490 410
rect 13526 378 13558 410
rect 13594 378 13626 410
rect 13662 378 13694 410
rect 13730 378 13762 410
rect 13798 378 13830 410
rect 13866 378 13898 410
rect 13934 378 13966 410
rect 14002 378 14034 410
rect 14070 378 14102 410
rect 14138 378 14170 410
rect 14206 378 14238 410
rect 14274 378 14306 410
rect 14342 378 14374 410
rect 14410 378 14442 410
rect 14478 378 14510 410
rect 14546 378 14578 410
rect 14614 378 14646 410
rect 14682 378 14714 410
rect 14750 378 14782 410
rect 14818 378 14850 410
rect 14886 378 14918 410
rect 14954 378 14986 410
rect 15022 378 15054 410
rect 15090 378 15122 410
rect 15158 378 15190 410
rect 15226 378 15258 410
rect 15294 378 15326 410
rect 15362 378 15394 410
rect 15430 378 15462 410
rect 15498 378 15530 410
rect 15566 378 15598 410
<< poly >>
rect 6856 3362 6976 3376
rect 6856 3330 6900 3362
rect 6932 3330 6976 3362
rect 6856 3302 6976 3330
rect 7212 3362 7332 3376
rect 7212 3330 7256 3362
rect 7288 3330 7332 3362
rect 7212 3302 7332 3330
rect 7460 3362 7580 3376
rect 7460 3330 7504 3362
rect 7536 3330 7580 3362
rect 7460 3302 7580 3330
rect 7816 3362 7936 3376
rect 7816 3330 7860 3362
rect 7892 3330 7936 3362
rect 7816 3302 7936 3330
rect 8064 3362 8184 3376
rect 8064 3330 8108 3362
rect 8140 3330 8184 3362
rect 8064 3302 8184 3330
rect 8420 3362 8540 3376
rect 8420 3330 8464 3362
rect 8496 3330 8540 3362
rect 8420 3302 8540 3330
rect 8668 3362 8788 3376
rect 8668 3330 8712 3362
rect 8744 3330 8788 3362
rect 8668 3302 8788 3330
rect 9024 3362 9144 3376
rect 9024 3330 9068 3362
rect 9100 3330 9144 3362
rect 9024 3302 9144 3330
rect 6856 1942 6976 1970
rect 6856 1910 6900 1942
rect 6932 1910 6976 1942
rect 6856 1882 6976 1910
rect 7212 1942 7332 1970
rect 7212 1910 7256 1942
rect 7288 1910 7332 1942
rect 7212 1882 7332 1910
rect 7460 1942 7580 1970
rect 7460 1910 7504 1942
rect 7536 1910 7580 1942
rect 7460 1882 7580 1910
rect 7816 1942 7936 1970
rect 7816 1910 7860 1942
rect 7892 1910 7936 1942
rect 7816 1882 7936 1910
rect 8064 1942 8184 1970
rect 8064 1910 8108 1942
rect 8140 1910 8184 1942
rect 8064 1882 8184 1910
rect 8420 1942 8540 1970
rect 8420 1910 8464 1942
rect 8496 1910 8540 1942
rect 8420 1882 8540 1910
rect 8668 1942 8788 1970
rect 8668 1910 8712 1942
rect 8744 1910 8788 1942
rect 8668 1882 8788 1910
rect 9024 1942 9144 1970
rect 9024 1910 9068 1942
rect 9100 1910 9144 1942
rect 9024 1882 9144 1910
rect 6856 522 6976 550
rect 6856 490 6900 522
rect 6932 490 6976 522
rect 6856 476 6976 490
rect 7212 522 7332 550
rect 7212 490 7256 522
rect 7288 490 7332 522
rect 7212 476 7332 490
rect 7460 522 7580 550
rect 7460 490 7504 522
rect 7536 490 7580 522
rect 7460 476 7580 490
rect 7816 522 7936 550
rect 7816 490 7860 522
rect 7892 490 7936 522
rect 7816 476 7936 490
rect 8064 522 8184 550
rect 8064 490 8108 522
rect 8140 490 8184 522
rect 8064 476 8184 490
rect 8420 522 8540 550
rect 8420 490 8464 522
rect 8496 490 8540 522
rect 8420 476 8540 490
rect 8668 522 8788 550
rect 8668 490 8712 522
rect 8744 490 8788 522
rect 8668 476 8788 490
rect 9024 522 9144 550
rect 9024 490 9068 522
rect 9100 490 9144 522
rect 9024 476 9144 490
<< polycont >>
rect 6900 3330 6932 3362
rect 7256 3330 7288 3362
rect 7504 3330 7536 3362
rect 7860 3330 7892 3362
rect 8108 3330 8140 3362
rect 8464 3330 8496 3362
rect 8712 3330 8744 3362
rect 9068 3330 9100 3362
rect 6900 1910 6932 1942
rect 7256 1910 7288 1942
rect 7504 1910 7536 1942
rect 7860 1910 7892 1942
rect 8108 1910 8140 1942
rect 8464 1910 8496 1942
rect 8712 1910 8744 1942
rect 9068 1910 9100 1942
rect 6900 490 6932 522
rect 7256 490 7288 522
rect 7504 490 7536 522
rect 7860 490 7892 522
rect 8108 490 8140 522
rect 8464 490 8496 522
rect 8712 490 8744 522
rect 9068 490 9100 522
<< pdiode >>
rect 3548 3236 3644 3268
rect 3548 3204 3580 3236
rect 3612 3204 3644 3236
rect 3548 3172 3644 3204
<< pdiodecont >>
rect 3580 3204 3612 3236
<< metal1 >>
rect 0 3834 16000 3852
rect 0 3802 28 3834
rect 60 3802 96 3834
rect 128 3802 164 3834
rect 196 3802 232 3834
rect 264 3802 300 3834
rect 332 3802 368 3834
rect 400 3802 436 3834
rect 468 3802 504 3834
rect 536 3802 572 3834
rect 604 3802 640 3834
rect 672 3802 708 3834
rect 740 3802 776 3834
rect 808 3802 844 3834
rect 876 3802 912 3834
rect 944 3802 980 3834
rect 1012 3802 1048 3834
rect 1080 3802 1116 3834
rect 1148 3802 1184 3834
rect 1216 3802 1252 3834
rect 1284 3802 1320 3834
rect 1352 3802 1388 3834
rect 1420 3802 1456 3834
rect 1488 3802 1524 3834
rect 1556 3802 1592 3834
rect 1624 3802 1660 3834
rect 1692 3802 1728 3834
rect 1760 3802 1796 3834
rect 1828 3802 1864 3834
rect 1896 3802 1932 3834
rect 1964 3802 2000 3834
rect 2032 3802 2068 3834
rect 2100 3802 2136 3834
rect 2168 3802 2204 3834
rect 2236 3802 2272 3834
rect 2304 3802 2340 3834
rect 2372 3802 2408 3834
rect 2440 3802 2476 3834
rect 2508 3802 2544 3834
rect 2576 3802 2612 3834
rect 2644 3802 2680 3834
rect 2712 3802 2748 3834
rect 2780 3802 2816 3834
rect 2848 3802 2884 3834
rect 2916 3802 2952 3834
rect 2984 3802 3020 3834
rect 3052 3802 3088 3834
rect 3120 3802 3156 3834
rect 3188 3802 3224 3834
rect 3256 3802 3292 3834
rect 3324 3802 3360 3834
rect 3392 3802 3428 3834
rect 3460 3802 3496 3834
rect 3528 3802 3564 3834
rect 3596 3802 3632 3834
rect 3664 3802 3700 3834
rect 3732 3802 3768 3834
rect 3800 3802 3836 3834
rect 3868 3802 3904 3834
rect 3936 3802 3972 3834
rect 4004 3802 4040 3834
rect 4072 3802 4108 3834
rect 4140 3802 4176 3834
rect 4208 3802 4244 3834
rect 4276 3802 4312 3834
rect 4344 3802 4380 3834
rect 4412 3802 4448 3834
rect 4480 3802 4516 3834
rect 4548 3802 4584 3834
rect 4616 3802 4652 3834
rect 4684 3802 4720 3834
rect 4752 3802 4788 3834
rect 4820 3802 4856 3834
rect 4888 3802 4924 3834
rect 4956 3802 4992 3834
rect 5024 3802 5060 3834
rect 5092 3802 5128 3834
rect 5160 3802 5196 3834
rect 5228 3802 5264 3834
rect 5296 3802 5332 3834
rect 5364 3802 5400 3834
rect 5432 3802 5468 3834
rect 5500 3802 5536 3834
rect 5568 3802 5604 3834
rect 5636 3802 5672 3834
rect 5704 3802 5740 3834
rect 5772 3802 5808 3834
rect 5840 3802 5876 3834
rect 5908 3802 5944 3834
rect 5976 3802 6012 3834
rect 6044 3802 6080 3834
rect 6112 3802 6148 3834
rect 6180 3802 6216 3834
rect 6248 3802 6284 3834
rect 6316 3802 6352 3834
rect 6384 3802 6420 3834
rect 6452 3802 6488 3834
rect 6520 3802 6556 3834
rect 6588 3802 6624 3834
rect 6656 3802 6692 3834
rect 6724 3802 6760 3834
rect 6792 3802 6828 3834
rect 6860 3802 6896 3834
rect 6928 3802 6964 3834
rect 6996 3802 7032 3834
rect 7064 3802 7100 3834
rect 7132 3802 7168 3834
rect 7200 3802 7236 3834
rect 7268 3802 7304 3834
rect 7336 3802 7372 3834
rect 7404 3802 7440 3834
rect 7472 3802 7508 3834
rect 7540 3802 7576 3834
rect 7608 3802 7644 3834
rect 7676 3802 7712 3834
rect 7744 3802 7780 3834
rect 7812 3802 7848 3834
rect 7880 3802 7916 3834
rect 7948 3802 7984 3834
rect 8016 3802 8052 3834
rect 8084 3802 8120 3834
rect 8152 3802 8188 3834
rect 8220 3802 8256 3834
rect 8288 3802 8324 3834
rect 8356 3802 8392 3834
rect 8424 3802 8460 3834
rect 8492 3802 8528 3834
rect 8560 3802 8596 3834
rect 8628 3802 8664 3834
rect 8696 3802 8732 3834
rect 8764 3802 8800 3834
rect 8832 3802 8868 3834
rect 8900 3802 8936 3834
rect 8968 3802 9004 3834
rect 9036 3802 9072 3834
rect 9104 3802 9140 3834
rect 9172 3802 9208 3834
rect 9240 3802 9276 3834
rect 9308 3802 9344 3834
rect 9376 3802 9412 3834
rect 9444 3802 9480 3834
rect 9512 3802 9548 3834
rect 9580 3802 9616 3834
rect 9648 3802 9684 3834
rect 9716 3802 9752 3834
rect 9784 3802 9820 3834
rect 9852 3802 9888 3834
rect 9920 3802 9956 3834
rect 9988 3802 10024 3834
rect 10056 3802 10092 3834
rect 10124 3802 10160 3834
rect 10192 3802 10228 3834
rect 10260 3802 10296 3834
rect 10328 3802 10364 3834
rect 10396 3802 10432 3834
rect 10464 3802 10500 3834
rect 10532 3802 10568 3834
rect 10600 3802 10636 3834
rect 10668 3802 10704 3834
rect 10736 3802 10772 3834
rect 10804 3802 10840 3834
rect 10872 3802 10908 3834
rect 10940 3802 10976 3834
rect 11008 3802 11044 3834
rect 11076 3802 11112 3834
rect 11144 3802 11180 3834
rect 11212 3802 11248 3834
rect 11280 3802 11316 3834
rect 11348 3802 11384 3834
rect 11416 3802 11452 3834
rect 11484 3802 11520 3834
rect 11552 3802 11588 3834
rect 11620 3802 11656 3834
rect 11688 3802 11724 3834
rect 11756 3802 11792 3834
rect 11824 3802 11860 3834
rect 11892 3802 11928 3834
rect 11960 3802 11996 3834
rect 12028 3802 12064 3834
rect 12096 3802 12132 3834
rect 12164 3802 12200 3834
rect 12232 3802 12268 3834
rect 12300 3802 12336 3834
rect 12368 3802 12404 3834
rect 12436 3802 12472 3834
rect 12504 3802 12540 3834
rect 12572 3802 12608 3834
rect 12640 3802 12676 3834
rect 12708 3802 12744 3834
rect 12776 3802 12812 3834
rect 12844 3802 12880 3834
rect 12912 3802 12948 3834
rect 12980 3802 13016 3834
rect 13048 3802 13084 3834
rect 13116 3802 13152 3834
rect 13184 3802 13220 3834
rect 13252 3802 13288 3834
rect 13320 3802 13356 3834
rect 13388 3802 13424 3834
rect 13456 3802 13492 3834
rect 13524 3802 13560 3834
rect 13592 3802 13628 3834
rect 13660 3802 13696 3834
rect 13728 3802 13764 3834
rect 13796 3802 13832 3834
rect 13864 3802 13900 3834
rect 13932 3802 13968 3834
rect 14000 3802 14036 3834
rect 14068 3802 14104 3834
rect 14136 3802 14172 3834
rect 14204 3802 14240 3834
rect 14272 3802 14308 3834
rect 14340 3802 14376 3834
rect 14408 3802 14444 3834
rect 14476 3802 14512 3834
rect 14544 3802 14580 3834
rect 14612 3802 14648 3834
rect 14680 3802 14716 3834
rect 14748 3802 14784 3834
rect 14816 3802 14852 3834
rect 14884 3802 14920 3834
rect 14952 3802 14988 3834
rect 15020 3802 15056 3834
rect 15088 3802 15124 3834
rect 15156 3802 15192 3834
rect 15224 3802 15260 3834
rect 15292 3802 15328 3834
rect 15360 3802 15396 3834
rect 15428 3802 15464 3834
rect 15496 3802 15532 3834
rect 15564 3802 15600 3834
rect 15632 3802 15668 3834
rect 15700 3802 15736 3834
rect 15768 3802 15804 3834
rect 15836 3802 15872 3834
rect 15904 3802 15940 3834
rect 15972 3802 16000 3834
rect 0 3784 16000 3802
rect 0 3744 68 3784
rect 0 3712 18 3744
rect 50 3712 68 3744
rect 0 3676 68 3712
rect 0 3644 18 3676
rect 50 3644 68 3676
rect 0 3608 68 3644
rect 0 3576 18 3608
rect 50 3576 68 3608
rect 0 3540 68 3576
rect 0 3508 18 3540
rect 50 3508 68 3540
rect 0 3472 68 3508
rect 15932 3744 16000 3784
rect 15932 3712 15950 3744
rect 15982 3712 16000 3744
rect 15932 3676 16000 3712
rect 15932 3644 15950 3676
rect 15982 3644 16000 3676
rect 15932 3608 16000 3644
rect 15932 3576 15950 3608
rect 15982 3576 16000 3608
rect 15932 3540 16000 3576
rect 15932 3508 15950 3540
rect 15982 3508 16000 3540
rect 0 3440 18 3472
rect 50 3440 68 3472
rect 0 3404 68 3440
rect 0 3372 18 3404
rect 50 3372 68 3404
rect 0 3336 68 3372
rect 0 3304 18 3336
rect 50 3304 68 3336
rect 0 3268 68 3304
rect 0 3236 18 3268
rect 50 3236 68 3268
rect 0 3200 68 3236
rect 0 3168 18 3200
rect 50 3168 68 3200
rect 0 3132 68 3168
rect 0 3100 18 3132
rect 50 3100 68 3132
rect 0 3064 68 3100
rect 0 3032 18 3064
rect 50 3032 68 3064
rect 0 2996 68 3032
rect 0 2964 18 2996
rect 50 2964 68 2996
rect 0 2928 68 2964
rect 0 2896 18 2928
rect 50 2896 68 2928
rect 0 2860 68 2896
rect 0 2828 18 2860
rect 50 2828 68 2860
rect 0 2792 68 2828
rect 0 2760 18 2792
rect 50 2760 68 2792
rect 0 2724 68 2760
rect 0 2692 18 2724
rect 50 2692 68 2724
rect 0 2656 68 2692
rect 0 2624 18 2656
rect 50 2624 68 2656
rect 0 2588 68 2624
rect 0 2556 18 2588
rect 50 2556 68 2588
rect 0 2520 68 2556
rect 0 2488 18 2520
rect 50 2488 68 2520
rect 0 2452 68 2488
rect 0 2420 18 2452
rect 50 2420 68 2452
rect 0 2384 68 2420
rect 0 2352 18 2384
rect 50 2352 68 2384
rect 0 2316 68 2352
rect 0 2284 18 2316
rect 50 2284 68 2316
rect 0 2248 68 2284
rect 0 2216 18 2248
rect 50 2216 68 2248
rect 0 2180 68 2216
rect 0 2148 18 2180
rect 50 2148 68 2180
rect 0 2112 68 2148
rect 0 2080 18 2112
rect 50 2080 68 2112
rect 0 2044 68 2080
rect 0 2012 18 2044
rect 50 2012 68 2044
rect 0 1976 68 2012
rect 0 1944 18 1976
rect 50 1944 68 1976
rect 0 1908 68 1944
rect 0 1876 18 1908
rect 50 1876 68 1908
rect 0 1840 68 1876
rect 0 1808 18 1840
rect 50 1808 68 1840
rect 0 1772 68 1808
rect 0 1740 18 1772
rect 50 1740 68 1772
rect 0 1704 68 1740
rect 0 1672 18 1704
rect 50 1672 68 1704
rect 0 1636 68 1672
rect 0 1604 18 1636
rect 50 1604 68 1636
rect 0 1568 68 1604
rect 0 1536 18 1568
rect 50 1536 68 1568
rect 0 1500 68 1536
rect 0 1468 18 1500
rect 50 1468 68 1500
rect 0 1432 68 1468
rect 0 1400 18 1432
rect 50 1400 68 1432
rect 0 1364 68 1400
rect 0 1332 18 1364
rect 50 1332 68 1364
rect 0 1296 68 1332
rect 0 1264 18 1296
rect 50 1264 68 1296
rect 0 1228 68 1264
rect 0 1196 18 1228
rect 50 1196 68 1228
rect 0 1160 68 1196
rect 0 1128 18 1160
rect 50 1128 68 1160
rect 0 1092 68 1128
rect 0 1060 18 1092
rect 50 1060 68 1092
rect 0 1024 68 1060
rect 0 992 18 1024
rect 50 992 68 1024
rect 0 956 68 992
rect 0 924 18 956
rect 50 924 68 956
rect 0 888 68 924
rect 0 856 18 888
rect 50 856 68 888
rect 0 820 68 856
rect 0 788 18 820
rect 50 788 68 820
rect 0 752 68 788
rect 0 720 18 752
rect 50 720 68 752
rect 0 684 68 720
rect 0 652 18 684
rect 50 652 68 684
rect 0 616 68 652
rect 0 584 18 616
rect 50 584 68 616
rect 0 548 68 584
rect 0 516 18 548
rect 50 516 68 548
rect 0 480 68 516
rect 0 448 18 480
rect 50 448 68 480
rect 0 412 68 448
rect 0 380 18 412
rect 50 380 68 412
rect 0 344 68 380
rect 360 3478 15640 3492
rect 360 3474 6772 3478
rect 6812 3474 7376 3478
rect 7416 3474 7980 3478
rect 8020 3474 8584 3478
rect 8624 3474 9188 3478
rect 9228 3474 15640 3478
rect 360 3442 402 3474
rect 434 3442 470 3474
rect 502 3442 538 3474
rect 570 3442 606 3474
rect 638 3442 674 3474
rect 706 3442 742 3474
rect 774 3442 810 3474
rect 842 3442 878 3474
rect 910 3442 946 3474
rect 978 3442 1014 3474
rect 1046 3442 1082 3474
rect 1114 3442 1150 3474
rect 1182 3442 1218 3474
rect 1250 3442 1286 3474
rect 1318 3442 1354 3474
rect 1386 3442 1422 3474
rect 1454 3442 1490 3474
rect 1522 3442 1558 3474
rect 1590 3442 1626 3474
rect 1658 3442 1694 3474
rect 1726 3442 1762 3474
rect 1794 3442 1830 3474
rect 1862 3442 1898 3474
rect 1930 3442 1966 3474
rect 1998 3442 2034 3474
rect 2066 3442 2102 3474
rect 2134 3442 2170 3474
rect 2202 3442 2238 3474
rect 2270 3442 2306 3474
rect 2338 3442 2374 3474
rect 2406 3442 2442 3474
rect 2474 3442 2510 3474
rect 2542 3442 2578 3474
rect 2610 3442 2646 3474
rect 2678 3442 2714 3474
rect 2746 3442 2782 3474
rect 2814 3442 2850 3474
rect 2882 3442 2918 3474
rect 2950 3442 2986 3474
rect 3018 3442 3054 3474
rect 3086 3442 3122 3474
rect 3154 3442 3190 3474
rect 3222 3442 3258 3474
rect 3290 3442 3326 3474
rect 3358 3442 3394 3474
rect 3426 3442 3462 3474
rect 3494 3442 3530 3474
rect 3562 3442 3598 3474
rect 3630 3442 3666 3474
rect 3698 3442 3734 3474
rect 3766 3442 3802 3474
rect 3834 3442 3870 3474
rect 3902 3442 3938 3474
rect 3970 3442 4006 3474
rect 4038 3442 4074 3474
rect 4106 3442 4142 3474
rect 4174 3442 4210 3474
rect 4242 3442 4278 3474
rect 4310 3442 4346 3474
rect 4378 3442 4414 3474
rect 4446 3442 4482 3474
rect 4514 3442 4550 3474
rect 4582 3442 4618 3474
rect 4650 3442 4686 3474
rect 4718 3442 4754 3474
rect 4786 3442 4822 3474
rect 4854 3442 4890 3474
rect 4922 3442 4958 3474
rect 4990 3442 5026 3474
rect 5058 3442 5094 3474
rect 5126 3442 5162 3474
rect 5194 3442 5230 3474
rect 5262 3442 5298 3474
rect 5330 3442 5366 3474
rect 5398 3442 5434 3474
rect 5466 3442 5502 3474
rect 5534 3442 5570 3474
rect 5602 3442 5638 3474
rect 5670 3442 5706 3474
rect 5738 3442 5774 3474
rect 5806 3442 5842 3474
rect 5874 3442 5910 3474
rect 5942 3442 5978 3474
rect 6010 3442 6046 3474
rect 6078 3442 6114 3474
rect 6146 3442 6182 3474
rect 6214 3442 6250 3474
rect 6282 3442 6318 3474
rect 6350 3442 6386 3474
rect 6418 3442 6454 3474
rect 6486 3442 6522 3474
rect 6554 3442 6590 3474
rect 6622 3442 6658 3474
rect 6690 3442 6726 3474
rect 6758 3442 6772 3474
rect 6826 3442 6862 3474
rect 6894 3442 6930 3474
rect 6962 3442 6998 3474
rect 7030 3442 7066 3474
rect 7098 3442 7134 3474
rect 7166 3442 7202 3474
rect 7234 3442 7270 3474
rect 7302 3442 7338 3474
rect 7370 3442 7376 3474
rect 7438 3442 7474 3474
rect 7506 3442 7542 3474
rect 7574 3442 7610 3474
rect 7642 3442 7678 3474
rect 7710 3442 7746 3474
rect 7778 3442 7814 3474
rect 7846 3442 7882 3474
rect 7914 3442 7950 3474
rect 8050 3442 8086 3474
rect 8118 3442 8154 3474
rect 8186 3442 8222 3474
rect 8254 3442 8290 3474
rect 8322 3442 8358 3474
rect 8390 3442 8426 3474
rect 8458 3442 8494 3474
rect 8526 3442 8562 3474
rect 8624 3442 8630 3474
rect 8662 3442 8698 3474
rect 8730 3442 8766 3474
rect 8798 3442 8834 3474
rect 8866 3442 8902 3474
rect 8934 3442 8970 3474
rect 9002 3442 9038 3474
rect 9070 3442 9106 3474
rect 9138 3442 9174 3474
rect 9228 3442 9242 3474
rect 9274 3442 9310 3474
rect 9342 3442 9378 3474
rect 9410 3442 9446 3474
rect 9478 3442 9514 3474
rect 9546 3442 9582 3474
rect 9614 3442 9650 3474
rect 9682 3442 9718 3474
rect 9750 3442 9786 3474
rect 9818 3442 9854 3474
rect 9886 3442 9922 3474
rect 9954 3442 9990 3474
rect 10022 3442 10058 3474
rect 10090 3442 10126 3474
rect 10158 3442 10194 3474
rect 10226 3442 10262 3474
rect 10294 3442 10330 3474
rect 10362 3442 10398 3474
rect 10430 3442 10466 3474
rect 10498 3442 10534 3474
rect 10566 3442 10602 3474
rect 10634 3442 10670 3474
rect 10702 3442 10738 3474
rect 10770 3442 10806 3474
rect 10838 3442 10874 3474
rect 10906 3442 10942 3474
rect 10974 3442 11010 3474
rect 11042 3442 11078 3474
rect 11110 3442 11146 3474
rect 11178 3442 11214 3474
rect 11246 3442 11282 3474
rect 11314 3442 11350 3474
rect 11382 3442 11418 3474
rect 11450 3442 11486 3474
rect 11518 3442 11554 3474
rect 11586 3442 11622 3474
rect 11654 3442 11690 3474
rect 11722 3442 11758 3474
rect 11790 3442 11826 3474
rect 11858 3442 11894 3474
rect 11926 3442 11962 3474
rect 11994 3442 12030 3474
rect 12062 3442 12098 3474
rect 12130 3442 12166 3474
rect 12198 3442 12234 3474
rect 12266 3442 12302 3474
rect 12334 3442 12370 3474
rect 12402 3442 12438 3474
rect 12470 3442 12506 3474
rect 12538 3442 12574 3474
rect 12606 3442 12642 3474
rect 12674 3442 12710 3474
rect 12742 3442 12778 3474
rect 12810 3442 12846 3474
rect 12878 3442 12914 3474
rect 12946 3442 12982 3474
rect 13014 3442 13050 3474
rect 13082 3442 13118 3474
rect 13150 3442 13186 3474
rect 13218 3442 13254 3474
rect 13286 3442 13322 3474
rect 13354 3442 13390 3474
rect 13422 3442 13458 3474
rect 13490 3442 13526 3474
rect 13558 3442 13594 3474
rect 13626 3442 13662 3474
rect 13694 3442 13730 3474
rect 13762 3442 13798 3474
rect 13830 3442 13866 3474
rect 13898 3442 13934 3474
rect 13966 3442 14002 3474
rect 14034 3442 14070 3474
rect 14102 3442 14138 3474
rect 14170 3442 14206 3474
rect 14238 3442 14274 3474
rect 14306 3442 14342 3474
rect 14374 3442 14410 3474
rect 14442 3442 14478 3474
rect 14510 3442 14546 3474
rect 14578 3442 14614 3474
rect 14646 3442 14682 3474
rect 14714 3442 14750 3474
rect 14782 3442 14818 3474
rect 14850 3442 14886 3474
rect 14918 3442 14954 3474
rect 14986 3442 15022 3474
rect 15054 3442 15090 3474
rect 15122 3442 15158 3474
rect 15190 3442 15226 3474
rect 15258 3442 15294 3474
rect 15326 3442 15362 3474
rect 15394 3442 15430 3474
rect 15462 3442 15498 3474
rect 15530 3442 15566 3474
rect 15598 3442 15640 3474
rect 360 3438 6772 3442
rect 6812 3438 7376 3442
rect 7416 3438 7980 3442
rect 8020 3438 8584 3442
rect 8624 3438 9188 3442
rect 9228 3438 15640 3442
rect 360 3424 15640 3438
rect 360 3370 428 3424
rect 360 3338 378 3370
rect 410 3338 428 3370
rect 360 3302 428 3338
rect 360 3270 378 3302
rect 410 3270 428 3302
rect 360 3234 428 3270
rect 3574 3362 9100 3378
rect 3574 3346 6900 3362
rect 3574 3336 3616 3346
rect 3574 3236 3575 3336
rect 360 3202 378 3234
rect 410 3202 428 3234
rect 3570 3214 3575 3236
rect 3615 3236 3616 3336
rect 6932 3346 7256 3362
rect 6771 3264 6813 3280
rect 3615 3214 3622 3236
rect 3570 3204 3622 3214
rect 6771 3232 6776 3264
rect 6808 3232 6813 3264
rect 6771 3230 6813 3232
rect 360 3166 428 3202
rect 3574 3172 3616 3204
rect 360 3134 378 3166
rect 410 3134 428 3166
rect 360 3098 428 3134
rect 360 3066 378 3098
rect 410 3066 428 3098
rect 360 3030 428 3066
rect 360 2998 378 3030
rect 410 2998 428 3030
rect 360 2962 428 2998
rect 360 2930 378 2962
rect 410 2930 428 2962
rect 360 2894 428 2930
rect 360 2862 378 2894
rect 410 2862 428 2894
rect 360 2826 428 2862
rect 360 2794 378 2826
rect 410 2794 428 2826
rect 360 2758 428 2794
rect 360 2726 378 2758
rect 410 2726 428 2758
rect 360 2690 428 2726
rect 360 2658 378 2690
rect 410 2658 428 2690
rect 360 2622 428 2658
rect 360 2590 378 2622
rect 410 2590 428 2622
rect 360 2554 428 2590
rect 360 2522 378 2554
rect 410 2522 428 2554
rect 360 2486 428 2522
rect 360 2454 378 2486
rect 410 2454 428 2486
rect 360 2418 428 2454
rect 360 2386 378 2418
rect 410 2386 428 2418
rect 360 2350 428 2386
rect 360 2318 378 2350
rect 410 2318 428 2350
rect 360 2282 428 2318
rect 360 2250 378 2282
rect 410 2250 428 2282
rect 360 2214 428 2250
rect 360 2182 378 2214
rect 410 2182 428 2214
rect 360 2146 428 2182
rect 360 2114 378 2146
rect 410 2114 428 2146
rect 360 2078 428 2114
rect 360 2046 378 2078
rect 410 2046 428 2078
rect 360 2010 428 2046
rect 360 1978 378 2010
rect 410 1978 428 2010
rect 6771 2042 6772 3230
rect 6812 2042 6813 3230
rect 6771 2040 6813 2042
rect 6771 2008 6776 2040
rect 6808 2008 6813 2040
rect 6771 1992 6813 2008
rect 360 1942 428 1978
rect 360 1910 378 1942
rect 410 1910 428 1942
rect 360 1874 428 1910
rect 360 1842 378 1874
rect 410 1842 428 1874
rect 6900 1942 6932 3330
rect 7288 3346 7504 3362
rect 7032 3264 7156 3280
rect 7032 3232 7078 3264
rect 7110 3232 7156 3264
rect 7032 3230 7156 3232
rect 7032 2042 7033 3230
rect 7155 2042 7156 3230
rect 7032 2040 7156 2042
rect 7032 2008 7078 2040
rect 7110 2008 7156 2040
rect 7032 1992 7156 2008
rect 360 1806 428 1842
rect 360 1774 378 1806
rect 410 1774 428 1806
rect 360 1738 428 1774
rect 360 1706 378 1738
rect 410 1706 428 1738
rect 360 1670 428 1706
rect 360 1638 378 1670
rect 410 1638 428 1670
rect 360 1602 428 1638
rect 360 1570 378 1602
rect 410 1570 428 1602
rect 360 1534 428 1570
rect 360 1502 378 1534
rect 410 1502 428 1534
rect 360 1466 428 1502
rect 360 1434 378 1466
rect 410 1434 428 1466
rect 360 1398 428 1434
rect 360 1366 378 1398
rect 410 1366 428 1398
rect 360 1330 428 1366
rect 360 1298 378 1330
rect 410 1298 428 1330
rect 360 1262 428 1298
rect 360 1230 378 1262
rect 410 1230 428 1262
rect 360 1194 428 1230
rect 360 1162 378 1194
rect 410 1162 428 1194
rect 360 1126 428 1162
rect 360 1094 378 1126
rect 410 1094 428 1126
rect 360 1058 428 1094
rect 360 1026 378 1058
rect 410 1026 428 1058
rect 360 990 428 1026
rect 360 958 378 990
rect 410 958 428 990
rect 360 922 428 958
rect 360 890 378 922
rect 410 890 428 922
rect 360 854 428 890
rect 360 822 378 854
rect 410 822 428 854
rect 360 786 428 822
rect 360 754 378 786
rect 410 754 428 786
rect 360 718 428 754
rect 360 686 378 718
rect 410 686 428 718
rect 360 650 428 686
rect 360 618 378 650
rect 410 618 428 650
rect 360 582 428 618
rect 360 550 378 582
rect 410 550 428 582
rect 6771 1844 6813 1860
rect 6771 1812 6776 1844
rect 6808 1812 6813 1844
rect 6771 1810 6813 1812
rect 6771 622 6772 1810
rect 6812 622 6813 1810
rect 6771 620 6813 622
rect 6771 588 6776 620
rect 6808 588 6813 620
rect 6771 572 6813 588
rect 360 514 428 550
rect 360 482 378 514
rect 410 482 428 514
rect 360 428 428 482
rect 6900 522 6932 1910
rect 7256 1942 7288 3330
rect 7536 3346 7860 3362
rect 7375 3264 7417 3280
rect 7375 3232 7380 3264
rect 7412 3232 7417 3264
rect 7375 3230 7417 3232
rect 7375 2042 7376 3230
rect 7416 2042 7417 3230
rect 7375 2040 7417 2042
rect 7375 2008 7380 2040
rect 7412 2008 7417 2040
rect 7375 1992 7417 2008
rect 7032 1844 7156 1860
rect 7032 1812 7078 1844
rect 7110 1812 7156 1844
rect 7032 1810 7156 1812
rect 7032 622 7033 1810
rect 7155 622 7156 1810
rect 7032 620 7156 622
rect 7032 588 7078 620
rect 7110 588 7156 620
rect 7032 572 7156 588
rect 6900 474 6932 490
rect 7256 522 7288 1910
rect 7504 1942 7536 3330
rect 7892 3346 8108 3362
rect 7636 3264 7760 3280
rect 7636 3232 7682 3264
rect 7714 3232 7760 3264
rect 7636 3230 7760 3232
rect 7636 2042 7637 3230
rect 7759 2042 7760 3230
rect 7636 2040 7760 2042
rect 7636 2008 7682 2040
rect 7714 2008 7760 2040
rect 7636 1992 7760 2008
rect 7375 1844 7417 1860
rect 7375 1812 7380 1844
rect 7412 1812 7417 1844
rect 7375 1810 7417 1812
rect 7375 622 7376 1810
rect 7416 622 7417 1810
rect 7375 620 7417 622
rect 7375 588 7380 620
rect 7412 588 7417 620
rect 7375 572 7417 588
rect 7256 474 7288 490
rect 7504 522 7536 1910
rect 7860 1942 7892 3330
rect 8140 3346 8464 3362
rect 7979 3264 8021 3280
rect 7979 3232 7984 3264
rect 8016 3232 8021 3264
rect 7979 3230 8021 3232
rect 7979 2042 7980 3230
rect 8020 2042 8021 3230
rect 7979 2040 8021 2042
rect 7979 2008 7984 2040
rect 8016 2008 8021 2040
rect 7979 1992 8021 2008
rect 7636 1844 7760 1860
rect 7636 1812 7682 1844
rect 7714 1812 7760 1844
rect 7636 1810 7760 1812
rect 7636 622 7637 1810
rect 7759 622 7760 1810
rect 7636 620 7760 622
rect 7636 588 7682 620
rect 7714 588 7760 620
rect 7636 572 7760 588
rect 7504 474 7536 490
rect 7860 522 7892 1910
rect 8108 1942 8140 3330
rect 8496 3346 8712 3362
rect 8240 3264 8364 3280
rect 8240 3232 8286 3264
rect 8318 3232 8364 3264
rect 8240 3230 8364 3232
rect 8240 2042 8241 3230
rect 8363 2042 8364 3230
rect 8240 2040 8364 2042
rect 8240 2008 8286 2040
rect 8318 2008 8364 2040
rect 8240 1992 8364 2008
rect 7979 1844 8021 1860
rect 7979 1812 7984 1844
rect 8016 1812 8021 1844
rect 7979 1810 8021 1812
rect 7979 622 7980 1810
rect 8020 622 8021 1810
rect 7979 620 8021 622
rect 7979 588 7984 620
rect 8016 588 8021 620
rect 7979 572 8021 588
rect 7860 474 7892 490
rect 8108 522 8140 1910
rect 8464 1942 8496 3330
rect 8744 3346 9068 3362
rect 8583 3264 8625 3280
rect 8583 3232 8588 3264
rect 8620 3232 8625 3264
rect 8583 3230 8625 3232
rect 8583 2042 8584 3230
rect 8624 2042 8625 3230
rect 8583 2040 8625 2042
rect 8583 2008 8588 2040
rect 8620 2008 8625 2040
rect 8583 1992 8625 2008
rect 8240 1844 8364 1860
rect 8240 1812 8286 1844
rect 8318 1812 8364 1844
rect 8240 1810 8364 1812
rect 8240 622 8241 1810
rect 8363 622 8364 1810
rect 8240 620 8364 622
rect 8240 588 8286 620
rect 8318 588 8364 620
rect 8240 572 8364 588
rect 8108 474 8140 490
rect 8464 522 8496 1910
rect 8712 1942 8744 3330
rect 8844 3264 8968 3280
rect 8844 3232 8890 3264
rect 8922 3232 8968 3264
rect 8844 3230 8968 3232
rect 8844 2042 8845 3230
rect 8967 2042 8968 3230
rect 8844 2040 8968 2042
rect 8844 2008 8890 2040
rect 8922 2008 8968 2040
rect 8844 1992 8968 2008
rect 8583 1844 8625 1860
rect 8583 1812 8588 1844
rect 8620 1812 8625 1844
rect 8583 1810 8625 1812
rect 8583 622 8584 1810
rect 8624 622 8625 1810
rect 8583 620 8625 622
rect 8583 588 8588 620
rect 8620 588 8625 620
rect 8583 572 8625 588
rect 8464 474 8496 490
rect 8712 522 8744 1910
rect 9068 1942 9100 3330
rect 15572 3370 15640 3424
rect 15572 3338 15590 3370
rect 15622 3338 15640 3370
rect 15572 3302 15640 3338
rect 9187 3264 9229 3280
rect 9187 3232 9192 3264
rect 9224 3232 9229 3264
rect 9187 3230 9229 3232
rect 9187 2042 9188 3230
rect 9228 2042 9229 3230
rect 9187 2040 9229 2042
rect 9187 2008 9192 2040
rect 9224 2008 9229 2040
rect 9187 1992 9229 2008
rect 15572 3270 15590 3302
rect 15622 3270 15640 3302
rect 15572 3234 15640 3270
rect 15572 3202 15590 3234
rect 15622 3202 15640 3234
rect 15572 3166 15640 3202
rect 15572 3134 15590 3166
rect 15622 3134 15640 3166
rect 15572 3098 15640 3134
rect 15572 3066 15590 3098
rect 15622 3066 15640 3098
rect 15572 3030 15640 3066
rect 15572 2998 15590 3030
rect 15622 2998 15640 3030
rect 15572 2962 15640 2998
rect 15572 2930 15590 2962
rect 15622 2930 15640 2962
rect 15572 2894 15640 2930
rect 15572 2862 15590 2894
rect 15622 2862 15640 2894
rect 15572 2826 15640 2862
rect 15572 2794 15590 2826
rect 15622 2794 15640 2826
rect 15572 2758 15640 2794
rect 15572 2726 15590 2758
rect 15622 2726 15640 2758
rect 15572 2690 15640 2726
rect 15572 2658 15590 2690
rect 15622 2658 15640 2690
rect 15572 2622 15640 2658
rect 15572 2590 15590 2622
rect 15622 2590 15640 2622
rect 15572 2554 15640 2590
rect 15572 2522 15590 2554
rect 15622 2522 15640 2554
rect 15572 2486 15640 2522
rect 15572 2454 15590 2486
rect 15622 2454 15640 2486
rect 15572 2418 15640 2454
rect 15572 2386 15590 2418
rect 15622 2386 15640 2418
rect 15572 2350 15640 2386
rect 15572 2318 15590 2350
rect 15622 2318 15640 2350
rect 15572 2282 15640 2318
rect 15572 2250 15590 2282
rect 15622 2250 15640 2282
rect 15572 2214 15640 2250
rect 15572 2182 15590 2214
rect 15622 2182 15640 2214
rect 15572 2146 15640 2182
rect 15572 2114 15590 2146
rect 15622 2114 15640 2146
rect 15572 2078 15640 2114
rect 15572 2046 15590 2078
rect 15622 2046 15640 2078
rect 15572 2010 15640 2046
rect 8844 1844 8968 1860
rect 8844 1812 8890 1844
rect 8922 1812 8968 1844
rect 8844 1810 8968 1812
rect 8844 622 8845 1810
rect 8967 622 8968 1810
rect 8844 620 8968 622
rect 8844 588 8890 620
rect 8922 588 8968 620
rect 8844 572 8968 588
rect 8712 474 8744 490
rect 9068 522 9100 1910
rect 15572 1978 15590 2010
rect 15622 1978 15640 2010
rect 15572 1942 15640 1978
rect 15572 1910 15590 1942
rect 15622 1910 15640 1942
rect 15572 1874 15640 1910
rect 9187 1844 9229 1860
rect 9187 1812 9192 1844
rect 9224 1812 9229 1844
rect 9187 1810 9229 1812
rect 9187 622 9188 1810
rect 9228 622 9229 1810
rect 9187 620 9229 622
rect 9187 588 9192 620
rect 9224 588 9229 620
rect 9187 572 9229 588
rect 15572 1842 15590 1874
rect 15622 1842 15640 1874
rect 15572 1806 15640 1842
rect 15572 1774 15590 1806
rect 15622 1774 15640 1806
rect 15572 1738 15640 1774
rect 15572 1706 15590 1738
rect 15622 1706 15640 1738
rect 15572 1670 15640 1706
rect 15572 1638 15590 1670
rect 15622 1638 15640 1670
rect 15572 1602 15640 1638
rect 15572 1570 15590 1602
rect 15622 1570 15640 1602
rect 15572 1534 15640 1570
rect 15572 1502 15590 1534
rect 15622 1502 15640 1534
rect 15572 1466 15640 1502
rect 15572 1434 15590 1466
rect 15622 1434 15640 1466
rect 15572 1398 15640 1434
rect 15572 1366 15590 1398
rect 15622 1366 15640 1398
rect 15572 1330 15640 1366
rect 15572 1298 15590 1330
rect 15622 1298 15640 1330
rect 15572 1262 15640 1298
rect 15572 1230 15590 1262
rect 15622 1230 15640 1262
rect 15572 1194 15640 1230
rect 15572 1162 15590 1194
rect 15622 1162 15640 1194
rect 15572 1126 15640 1162
rect 15572 1094 15590 1126
rect 15622 1094 15640 1126
rect 15572 1058 15640 1094
rect 15572 1026 15590 1058
rect 15622 1026 15640 1058
rect 15572 990 15640 1026
rect 15572 958 15590 990
rect 15622 958 15640 990
rect 15572 922 15640 958
rect 15572 890 15590 922
rect 15622 890 15640 922
rect 15572 854 15640 890
rect 15572 822 15590 854
rect 15622 822 15640 854
rect 15572 786 15640 822
rect 15572 754 15590 786
rect 15622 754 15640 786
rect 15572 718 15640 754
rect 15572 686 15590 718
rect 15622 686 15640 718
rect 15572 650 15640 686
rect 15572 618 15590 650
rect 15622 618 15640 650
rect 15572 582 15640 618
rect 9068 474 9100 490
rect 15572 550 15590 582
rect 15622 550 15640 582
rect 15572 514 15640 550
rect 15572 482 15590 514
rect 15622 482 15640 514
rect 15572 428 15640 482
rect 360 414 15640 428
rect 360 410 6772 414
rect 6812 410 7376 414
rect 7416 410 7980 414
rect 8020 410 8584 414
rect 8624 410 9188 414
rect 9228 410 15640 414
rect 360 378 402 410
rect 434 378 470 410
rect 502 378 538 410
rect 570 378 606 410
rect 638 378 674 410
rect 706 378 742 410
rect 774 378 810 410
rect 842 378 878 410
rect 910 378 946 410
rect 978 378 1014 410
rect 1046 378 1082 410
rect 1114 378 1150 410
rect 1182 378 1218 410
rect 1250 378 1286 410
rect 1318 378 1354 410
rect 1386 378 1422 410
rect 1454 378 1490 410
rect 1522 378 1558 410
rect 1590 378 1626 410
rect 1658 378 1694 410
rect 1726 378 1762 410
rect 1794 378 1830 410
rect 1862 378 1898 410
rect 1930 378 1966 410
rect 1998 378 2034 410
rect 2066 378 2102 410
rect 2134 378 2170 410
rect 2202 378 2238 410
rect 2270 378 2306 410
rect 2338 378 2374 410
rect 2406 378 2442 410
rect 2474 378 2510 410
rect 2542 378 2578 410
rect 2610 378 2646 410
rect 2678 378 2714 410
rect 2746 378 2782 410
rect 2814 378 2850 410
rect 2882 378 2918 410
rect 2950 378 2986 410
rect 3018 378 3054 410
rect 3086 378 3122 410
rect 3154 378 3190 410
rect 3222 378 3258 410
rect 3290 378 3326 410
rect 3358 378 3394 410
rect 3426 378 3462 410
rect 3494 378 3530 410
rect 3562 378 3598 410
rect 3630 378 3666 410
rect 3698 378 3734 410
rect 3766 378 3802 410
rect 3834 378 3870 410
rect 3902 378 3938 410
rect 3970 378 4006 410
rect 4038 378 4074 410
rect 4106 378 4142 410
rect 4174 378 4210 410
rect 4242 378 4278 410
rect 4310 378 4346 410
rect 4378 378 4414 410
rect 4446 378 4482 410
rect 4514 378 4550 410
rect 4582 378 4618 410
rect 4650 378 4686 410
rect 4718 378 4754 410
rect 4786 378 4822 410
rect 4854 378 4890 410
rect 4922 378 4958 410
rect 4990 378 5026 410
rect 5058 378 5094 410
rect 5126 378 5162 410
rect 5194 378 5230 410
rect 5262 378 5298 410
rect 5330 378 5366 410
rect 5398 378 5434 410
rect 5466 378 5502 410
rect 5534 378 5570 410
rect 5602 378 5638 410
rect 5670 378 5706 410
rect 5738 378 5774 410
rect 5806 378 5842 410
rect 5874 378 5910 410
rect 5942 378 5978 410
rect 6010 378 6046 410
rect 6078 378 6114 410
rect 6146 378 6182 410
rect 6214 378 6250 410
rect 6282 378 6318 410
rect 6350 378 6386 410
rect 6418 378 6454 410
rect 6486 378 6522 410
rect 6554 378 6590 410
rect 6622 378 6658 410
rect 6690 378 6726 410
rect 6758 378 6772 410
rect 6826 378 6862 410
rect 6894 378 6930 410
rect 6962 378 6998 410
rect 7030 378 7066 410
rect 7098 378 7134 410
rect 7166 378 7202 410
rect 7234 378 7270 410
rect 7302 378 7338 410
rect 7370 378 7376 410
rect 7438 378 7474 410
rect 7506 378 7542 410
rect 7574 378 7610 410
rect 7642 378 7678 410
rect 7710 378 7746 410
rect 7778 378 7814 410
rect 7846 378 7882 410
rect 7914 378 7950 410
rect 8050 378 8086 410
rect 8118 378 8154 410
rect 8186 378 8222 410
rect 8254 378 8290 410
rect 8322 378 8358 410
rect 8390 378 8426 410
rect 8458 378 8494 410
rect 8526 378 8562 410
rect 8624 378 8630 410
rect 8662 378 8698 410
rect 8730 378 8766 410
rect 8798 378 8834 410
rect 8866 378 8902 410
rect 8934 378 8970 410
rect 9002 378 9038 410
rect 9070 378 9106 410
rect 9138 378 9174 410
rect 9228 378 9242 410
rect 9274 378 9310 410
rect 9342 378 9378 410
rect 9410 378 9446 410
rect 9478 378 9514 410
rect 9546 378 9582 410
rect 9614 378 9650 410
rect 9682 378 9718 410
rect 9750 378 9786 410
rect 9818 378 9854 410
rect 9886 378 9922 410
rect 9954 378 9990 410
rect 10022 378 10058 410
rect 10090 378 10126 410
rect 10158 378 10194 410
rect 10226 378 10262 410
rect 10294 378 10330 410
rect 10362 378 10398 410
rect 10430 378 10466 410
rect 10498 378 10534 410
rect 10566 378 10602 410
rect 10634 378 10670 410
rect 10702 378 10738 410
rect 10770 378 10806 410
rect 10838 378 10874 410
rect 10906 378 10942 410
rect 10974 378 11010 410
rect 11042 378 11078 410
rect 11110 378 11146 410
rect 11178 378 11214 410
rect 11246 378 11282 410
rect 11314 378 11350 410
rect 11382 378 11418 410
rect 11450 378 11486 410
rect 11518 378 11554 410
rect 11586 378 11622 410
rect 11654 378 11690 410
rect 11722 378 11758 410
rect 11790 378 11826 410
rect 11858 378 11894 410
rect 11926 378 11962 410
rect 11994 378 12030 410
rect 12062 378 12098 410
rect 12130 378 12166 410
rect 12198 378 12234 410
rect 12266 378 12302 410
rect 12334 378 12370 410
rect 12402 378 12438 410
rect 12470 378 12506 410
rect 12538 378 12574 410
rect 12606 378 12642 410
rect 12674 378 12710 410
rect 12742 378 12778 410
rect 12810 378 12846 410
rect 12878 378 12914 410
rect 12946 378 12982 410
rect 13014 378 13050 410
rect 13082 378 13118 410
rect 13150 378 13186 410
rect 13218 378 13254 410
rect 13286 378 13322 410
rect 13354 378 13390 410
rect 13422 378 13458 410
rect 13490 378 13526 410
rect 13558 378 13594 410
rect 13626 378 13662 410
rect 13694 378 13730 410
rect 13762 378 13798 410
rect 13830 378 13866 410
rect 13898 378 13934 410
rect 13966 378 14002 410
rect 14034 378 14070 410
rect 14102 378 14138 410
rect 14170 378 14206 410
rect 14238 378 14274 410
rect 14306 378 14342 410
rect 14374 378 14410 410
rect 14442 378 14478 410
rect 14510 378 14546 410
rect 14578 378 14614 410
rect 14646 378 14682 410
rect 14714 378 14750 410
rect 14782 378 14818 410
rect 14850 378 14886 410
rect 14918 378 14954 410
rect 14986 378 15022 410
rect 15054 378 15090 410
rect 15122 378 15158 410
rect 15190 378 15226 410
rect 15258 378 15294 410
rect 15326 378 15362 410
rect 15394 378 15430 410
rect 15462 378 15498 410
rect 15530 378 15566 410
rect 15598 378 15640 410
rect 360 374 6772 378
rect 6812 374 7376 378
rect 7416 374 7980 378
rect 8020 374 8584 378
rect 8624 374 9188 378
rect 9228 374 15640 378
rect 360 360 15640 374
rect 15932 3472 16000 3508
rect 15932 3440 15950 3472
rect 15982 3440 16000 3472
rect 15932 3404 16000 3440
rect 15932 3372 15950 3404
rect 15982 3372 16000 3404
rect 15932 3336 16000 3372
rect 15932 3304 15950 3336
rect 15982 3304 16000 3336
rect 15932 3268 16000 3304
rect 15932 3236 15950 3268
rect 15982 3236 16000 3268
rect 15932 3200 16000 3236
rect 15932 3168 15950 3200
rect 15982 3168 16000 3200
rect 15932 3132 16000 3168
rect 15932 3100 15950 3132
rect 15982 3100 16000 3132
rect 15932 3064 16000 3100
rect 15932 3032 15950 3064
rect 15982 3032 16000 3064
rect 15932 2996 16000 3032
rect 15932 2964 15950 2996
rect 15982 2964 16000 2996
rect 15932 2928 16000 2964
rect 15932 2896 15950 2928
rect 15982 2896 16000 2928
rect 15932 2860 16000 2896
rect 15932 2828 15950 2860
rect 15982 2828 16000 2860
rect 15932 2792 16000 2828
rect 15932 2760 15950 2792
rect 15982 2760 16000 2792
rect 15932 2724 16000 2760
rect 15932 2692 15950 2724
rect 15982 2692 16000 2724
rect 15932 2656 16000 2692
rect 15932 2624 15950 2656
rect 15982 2624 16000 2656
rect 15932 2588 16000 2624
rect 15932 2556 15950 2588
rect 15982 2556 16000 2588
rect 15932 2520 16000 2556
rect 15932 2488 15950 2520
rect 15982 2488 16000 2520
rect 15932 2452 16000 2488
rect 15932 2420 15950 2452
rect 15982 2420 16000 2452
rect 15932 2384 16000 2420
rect 15932 2352 15950 2384
rect 15982 2352 16000 2384
rect 15932 2316 16000 2352
rect 15932 2284 15950 2316
rect 15982 2284 16000 2316
rect 15932 2248 16000 2284
rect 15932 2216 15950 2248
rect 15982 2216 16000 2248
rect 15932 2180 16000 2216
rect 15932 2148 15950 2180
rect 15982 2148 16000 2180
rect 15932 2112 16000 2148
rect 15932 2080 15950 2112
rect 15982 2080 16000 2112
rect 15932 2044 16000 2080
rect 15932 2012 15950 2044
rect 15982 2012 16000 2044
rect 15932 1976 16000 2012
rect 15932 1944 15950 1976
rect 15982 1944 16000 1976
rect 15932 1908 16000 1944
rect 15932 1876 15950 1908
rect 15982 1876 16000 1908
rect 15932 1840 16000 1876
rect 15932 1808 15950 1840
rect 15982 1808 16000 1840
rect 15932 1772 16000 1808
rect 15932 1740 15950 1772
rect 15982 1740 16000 1772
rect 15932 1704 16000 1740
rect 15932 1672 15950 1704
rect 15982 1672 16000 1704
rect 15932 1636 16000 1672
rect 15932 1604 15950 1636
rect 15982 1604 16000 1636
rect 15932 1568 16000 1604
rect 15932 1536 15950 1568
rect 15982 1536 16000 1568
rect 15932 1500 16000 1536
rect 15932 1468 15950 1500
rect 15982 1468 16000 1500
rect 15932 1432 16000 1468
rect 15932 1400 15950 1432
rect 15982 1400 16000 1432
rect 15932 1364 16000 1400
rect 15932 1332 15950 1364
rect 15982 1332 16000 1364
rect 15932 1296 16000 1332
rect 15932 1264 15950 1296
rect 15982 1264 16000 1296
rect 15932 1228 16000 1264
rect 15932 1196 15950 1228
rect 15982 1196 16000 1228
rect 15932 1160 16000 1196
rect 15932 1128 15950 1160
rect 15982 1128 16000 1160
rect 15932 1092 16000 1128
rect 15932 1060 15950 1092
rect 15982 1060 16000 1092
rect 15932 1024 16000 1060
rect 15932 992 15950 1024
rect 15982 992 16000 1024
rect 15932 956 16000 992
rect 15932 924 15950 956
rect 15982 924 16000 956
rect 15932 888 16000 924
rect 15932 856 15950 888
rect 15982 856 16000 888
rect 15932 820 16000 856
rect 15932 788 15950 820
rect 15982 788 16000 820
rect 15932 752 16000 788
rect 15932 720 15950 752
rect 15982 720 16000 752
rect 15932 684 16000 720
rect 15932 652 15950 684
rect 15982 652 16000 684
rect 15932 616 16000 652
rect 15932 584 15950 616
rect 15982 584 16000 616
rect 15932 548 16000 584
rect 15932 516 15950 548
rect 15982 516 16000 548
rect 15932 480 16000 516
rect 15932 448 15950 480
rect 15982 448 16000 480
rect 15932 412 16000 448
rect 15932 380 15950 412
rect 15982 380 16000 412
rect 0 312 18 344
rect 50 312 68 344
rect 0 276 68 312
rect 0 244 18 276
rect 50 244 68 276
rect 0 208 68 244
rect 0 176 18 208
rect 50 176 68 208
rect 0 140 68 176
rect 0 108 18 140
rect 50 108 68 140
rect 0 68 68 108
rect 15932 344 16000 380
rect 15932 312 15950 344
rect 15982 312 16000 344
rect 15932 276 16000 312
rect 15932 244 15950 276
rect 15982 244 16000 276
rect 15932 208 16000 244
rect 15932 176 15950 208
rect 15982 176 16000 208
rect 15932 140 16000 176
rect 15932 108 15950 140
rect 15982 108 16000 140
rect 15932 68 16000 108
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 0 16000 18
<< via1 >>
rect 6772 3474 6812 3478
rect 7376 3474 7416 3478
rect 7980 3474 8020 3478
rect 8584 3474 8624 3478
rect 9188 3474 9228 3478
rect 6772 3442 6794 3474
rect 6794 3442 6812 3474
rect 7376 3442 7406 3474
rect 7406 3442 7416 3474
rect 7980 3442 7982 3474
rect 7982 3442 8018 3474
rect 8018 3442 8020 3474
rect 8584 3442 8594 3474
rect 8594 3442 8624 3474
rect 9188 3442 9206 3474
rect 9206 3442 9228 3474
rect 6772 3438 6812 3442
rect 7376 3438 7416 3442
rect 7980 3438 8020 3442
rect 8584 3438 8624 3442
rect 9188 3438 9228 3442
rect 3575 3214 3615 3336
rect 6772 3196 6812 3230
rect 6772 3164 6776 3196
rect 6776 3164 6808 3196
rect 6808 3164 6812 3196
rect 6772 3128 6812 3164
rect 6772 3096 6776 3128
rect 6776 3096 6808 3128
rect 6808 3096 6812 3128
rect 6772 3060 6812 3096
rect 6772 3028 6776 3060
rect 6776 3028 6808 3060
rect 6808 3028 6812 3060
rect 6772 2992 6812 3028
rect 6772 2960 6776 2992
rect 6776 2960 6808 2992
rect 6808 2960 6812 2992
rect 6772 2924 6812 2960
rect 6772 2892 6776 2924
rect 6776 2892 6808 2924
rect 6808 2892 6812 2924
rect 6772 2856 6812 2892
rect 6772 2824 6776 2856
rect 6776 2824 6808 2856
rect 6808 2824 6812 2856
rect 6772 2788 6812 2824
rect 6772 2756 6776 2788
rect 6776 2756 6808 2788
rect 6808 2756 6812 2788
rect 6772 2720 6812 2756
rect 6772 2688 6776 2720
rect 6776 2688 6808 2720
rect 6808 2688 6812 2720
rect 6772 2652 6812 2688
rect 6772 2620 6776 2652
rect 6776 2620 6808 2652
rect 6808 2620 6812 2652
rect 6772 2584 6812 2620
rect 6772 2552 6776 2584
rect 6776 2552 6808 2584
rect 6808 2552 6812 2584
rect 6772 2516 6812 2552
rect 6772 2484 6776 2516
rect 6776 2484 6808 2516
rect 6808 2484 6812 2516
rect 6772 2448 6812 2484
rect 6772 2416 6776 2448
rect 6776 2416 6808 2448
rect 6808 2416 6812 2448
rect 6772 2380 6812 2416
rect 6772 2348 6776 2380
rect 6776 2348 6808 2380
rect 6808 2348 6812 2380
rect 6772 2312 6812 2348
rect 6772 2280 6776 2312
rect 6776 2280 6808 2312
rect 6808 2280 6812 2312
rect 6772 2244 6812 2280
rect 6772 2212 6776 2244
rect 6776 2212 6808 2244
rect 6808 2212 6812 2244
rect 6772 2176 6812 2212
rect 6772 2144 6776 2176
rect 6776 2144 6808 2176
rect 6808 2144 6812 2176
rect 6772 2108 6812 2144
rect 6772 2076 6776 2108
rect 6776 2076 6808 2108
rect 6808 2076 6812 2108
rect 6772 2042 6812 2076
rect 7033 3196 7155 3230
rect 7033 3164 7078 3196
rect 7078 3164 7110 3196
rect 7110 3164 7155 3196
rect 7033 3128 7155 3164
rect 7033 3096 7078 3128
rect 7078 3096 7110 3128
rect 7110 3096 7155 3128
rect 7033 3060 7155 3096
rect 7033 3028 7078 3060
rect 7078 3028 7110 3060
rect 7110 3028 7155 3060
rect 7033 2992 7155 3028
rect 7033 2960 7078 2992
rect 7078 2960 7110 2992
rect 7110 2960 7155 2992
rect 7033 2924 7155 2960
rect 7033 2892 7078 2924
rect 7078 2892 7110 2924
rect 7110 2892 7155 2924
rect 7033 2856 7155 2892
rect 7033 2824 7078 2856
rect 7078 2824 7110 2856
rect 7110 2824 7155 2856
rect 7033 2788 7155 2824
rect 7033 2756 7078 2788
rect 7078 2756 7110 2788
rect 7110 2756 7155 2788
rect 7033 2720 7155 2756
rect 7033 2688 7078 2720
rect 7078 2688 7110 2720
rect 7110 2688 7155 2720
rect 7033 2652 7155 2688
rect 7033 2620 7078 2652
rect 7078 2620 7110 2652
rect 7110 2620 7155 2652
rect 7033 2584 7155 2620
rect 7033 2552 7078 2584
rect 7078 2552 7110 2584
rect 7110 2552 7155 2584
rect 7033 2516 7155 2552
rect 7033 2484 7078 2516
rect 7078 2484 7110 2516
rect 7110 2484 7155 2516
rect 7033 2448 7155 2484
rect 7033 2416 7078 2448
rect 7078 2416 7110 2448
rect 7110 2416 7155 2448
rect 7033 2380 7155 2416
rect 7033 2348 7078 2380
rect 7078 2348 7110 2380
rect 7110 2348 7155 2380
rect 7033 2312 7155 2348
rect 7033 2280 7078 2312
rect 7078 2280 7110 2312
rect 7110 2280 7155 2312
rect 7033 2244 7155 2280
rect 7033 2212 7078 2244
rect 7078 2212 7110 2244
rect 7110 2212 7155 2244
rect 7033 2176 7155 2212
rect 7033 2144 7078 2176
rect 7078 2144 7110 2176
rect 7110 2144 7155 2176
rect 7033 2108 7155 2144
rect 7033 2076 7078 2108
rect 7078 2076 7110 2108
rect 7110 2076 7155 2108
rect 7033 2042 7155 2076
rect 6772 1776 6812 1810
rect 6772 1744 6776 1776
rect 6776 1744 6808 1776
rect 6808 1744 6812 1776
rect 6772 1708 6812 1744
rect 6772 1676 6776 1708
rect 6776 1676 6808 1708
rect 6808 1676 6812 1708
rect 6772 1640 6812 1676
rect 6772 1608 6776 1640
rect 6776 1608 6808 1640
rect 6808 1608 6812 1640
rect 6772 1572 6812 1608
rect 6772 1540 6776 1572
rect 6776 1540 6808 1572
rect 6808 1540 6812 1572
rect 6772 1504 6812 1540
rect 6772 1472 6776 1504
rect 6776 1472 6808 1504
rect 6808 1472 6812 1504
rect 6772 1436 6812 1472
rect 6772 1404 6776 1436
rect 6776 1404 6808 1436
rect 6808 1404 6812 1436
rect 6772 1368 6812 1404
rect 6772 1336 6776 1368
rect 6776 1336 6808 1368
rect 6808 1336 6812 1368
rect 6772 1300 6812 1336
rect 6772 1268 6776 1300
rect 6776 1268 6808 1300
rect 6808 1268 6812 1300
rect 6772 1232 6812 1268
rect 6772 1200 6776 1232
rect 6776 1200 6808 1232
rect 6808 1200 6812 1232
rect 6772 1164 6812 1200
rect 6772 1132 6776 1164
rect 6776 1132 6808 1164
rect 6808 1132 6812 1164
rect 6772 1096 6812 1132
rect 6772 1064 6776 1096
rect 6776 1064 6808 1096
rect 6808 1064 6812 1096
rect 6772 1028 6812 1064
rect 6772 996 6776 1028
rect 6776 996 6808 1028
rect 6808 996 6812 1028
rect 6772 960 6812 996
rect 6772 928 6776 960
rect 6776 928 6808 960
rect 6808 928 6812 960
rect 6772 892 6812 928
rect 6772 860 6776 892
rect 6776 860 6808 892
rect 6808 860 6812 892
rect 6772 824 6812 860
rect 6772 792 6776 824
rect 6776 792 6808 824
rect 6808 792 6812 824
rect 6772 756 6812 792
rect 6772 724 6776 756
rect 6776 724 6808 756
rect 6808 724 6812 756
rect 6772 688 6812 724
rect 6772 656 6776 688
rect 6776 656 6808 688
rect 6808 656 6812 688
rect 6772 622 6812 656
rect 7376 3196 7416 3230
rect 7376 3164 7380 3196
rect 7380 3164 7412 3196
rect 7412 3164 7416 3196
rect 7376 3128 7416 3164
rect 7376 3096 7380 3128
rect 7380 3096 7412 3128
rect 7412 3096 7416 3128
rect 7376 3060 7416 3096
rect 7376 3028 7380 3060
rect 7380 3028 7412 3060
rect 7412 3028 7416 3060
rect 7376 2992 7416 3028
rect 7376 2960 7380 2992
rect 7380 2960 7412 2992
rect 7412 2960 7416 2992
rect 7376 2924 7416 2960
rect 7376 2892 7380 2924
rect 7380 2892 7412 2924
rect 7412 2892 7416 2924
rect 7376 2856 7416 2892
rect 7376 2824 7380 2856
rect 7380 2824 7412 2856
rect 7412 2824 7416 2856
rect 7376 2788 7416 2824
rect 7376 2756 7380 2788
rect 7380 2756 7412 2788
rect 7412 2756 7416 2788
rect 7376 2720 7416 2756
rect 7376 2688 7380 2720
rect 7380 2688 7412 2720
rect 7412 2688 7416 2720
rect 7376 2652 7416 2688
rect 7376 2620 7380 2652
rect 7380 2620 7412 2652
rect 7412 2620 7416 2652
rect 7376 2584 7416 2620
rect 7376 2552 7380 2584
rect 7380 2552 7412 2584
rect 7412 2552 7416 2584
rect 7376 2516 7416 2552
rect 7376 2484 7380 2516
rect 7380 2484 7412 2516
rect 7412 2484 7416 2516
rect 7376 2448 7416 2484
rect 7376 2416 7380 2448
rect 7380 2416 7412 2448
rect 7412 2416 7416 2448
rect 7376 2380 7416 2416
rect 7376 2348 7380 2380
rect 7380 2348 7412 2380
rect 7412 2348 7416 2380
rect 7376 2312 7416 2348
rect 7376 2280 7380 2312
rect 7380 2280 7412 2312
rect 7412 2280 7416 2312
rect 7376 2244 7416 2280
rect 7376 2212 7380 2244
rect 7380 2212 7412 2244
rect 7412 2212 7416 2244
rect 7376 2176 7416 2212
rect 7376 2144 7380 2176
rect 7380 2144 7412 2176
rect 7412 2144 7416 2176
rect 7376 2108 7416 2144
rect 7376 2076 7380 2108
rect 7380 2076 7412 2108
rect 7412 2076 7416 2108
rect 7376 2042 7416 2076
rect 7033 1776 7155 1810
rect 7033 1744 7078 1776
rect 7078 1744 7110 1776
rect 7110 1744 7155 1776
rect 7033 1708 7155 1744
rect 7033 1676 7078 1708
rect 7078 1676 7110 1708
rect 7110 1676 7155 1708
rect 7033 1640 7155 1676
rect 7033 1608 7078 1640
rect 7078 1608 7110 1640
rect 7110 1608 7155 1640
rect 7033 1572 7155 1608
rect 7033 1540 7078 1572
rect 7078 1540 7110 1572
rect 7110 1540 7155 1572
rect 7033 1504 7155 1540
rect 7033 1472 7078 1504
rect 7078 1472 7110 1504
rect 7110 1472 7155 1504
rect 7033 1436 7155 1472
rect 7033 1404 7078 1436
rect 7078 1404 7110 1436
rect 7110 1404 7155 1436
rect 7033 1368 7155 1404
rect 7033 1336 7078 1368
rect 7078 1336 7110 1368
rect 7110 1336 7155 1368
rect 7033 1300 7155 1336
rect 7033 1268 7078 1300
rect 7078 1268 7110 1300
rect 7110 1268 7155 1300
rect 7033 1232 7155 1268
rect 7033 1200 7078 1232
rect 7078 1200 7110 1232
rect 7110 1200 7155 1232
rect 7033 1164 7155 1200
rect 7033 1132 7078 1164
rect 7078 1132 7110 1164
rect 7110 1132 7155 1164
rect 7033 1096 7155 1132
rect 7033 1064 7078 1096
rect 7078 1064 7110 1096
rect 7110 1064 7155 1096
rect 7033 1028 7155 1064
rect 7033 996 7078 1028
rect 7078 996 7110 1028
rect 7110 996 7155 1028
rect 7033 960 7155 996
rect 7033 928 7078 960
rect 7078 928 7110 960
rect 7110 928 7155 960
rect 7033 892 7155 928
rect 7033 860 7078 892
rect 7078 860 7110 892
rect 7110 860 7155 892
rect 7033 824 7155 860
rect 7033 792 7078 824
rect 7078 792 7110 824
rect 7110 792 7155 824
rect 7033 756 7155 792
rect 7033 724 7078 756
rect 7078 724 7110 756
rect 7110 724 7155 756
rect 7033 688 7155 724
rect 7033 656 7078 688
rect 7078 656 7110 688
rect 7110 656 7155 688
rect 7033 622 7155 656
rect 7637 3196 7759 3230
rect 7637 3164 7682 3196
rect 7682 3164 7714 3196
rect 7714 3164 7759 3196
rect 7637 3128 7759 3164
rect 7637 3096 7682 3128
rect 7682 3096 7714 3128
rect 7714 3096 7759 3128
rect 7637 3060 7759 3096
rect 7637 3028 7682 3060
rect 7682 3028 7714 3060
rect 7714 3028 7759 3060
rect 7637 2992 7759 3028
rect 7637 2960 7682 2992
rect 7682 2960 7714 2992
rect 7714 2960 7759 2992
rect 7637 2924 7759 2960
rect 7637 2892 7682 2924
rect 7682 2892 7714 2924
rect 7714 2892 7759 2924
rect 7637 2856 7759 2892
rect 7637 2824 7682 2856
rect 7682 2824 7714 2856
rect 7714 2824 7759 2856
rect 7637 2788 7759 2824
rect 7637 2756 7682 2788
rect 7682 2756 7714 2788
rect 7714 2756 7759 2788
rect 7637 2720 7759 2756
rect 7637 2688 7682 2720
rect 7682 2688 7714 2720
rect 7714 2688 7759 2720
rect 7637 2652 7759 2688
rect 7637 2620 7682 2652
rect 7682 2620 7714 2652
rect 7714 2620 7759 2652
rect 7637 2584 7759 2620
rect 7637 2552 7682 2584
rect 7682 2552 7714 2584
rect 7714 2552 7759 2584
rect 7637 2516 7759 2552
rect 7637 2484 7682 2516
rect 7682 2484 7714 2516
rect 7714 2484 7759 2516
rect 7637 2448 7759 2484
rect 7637 2416 7682 2448
rect 7682 2416 7714 2448
rect 7714 2416 7759 2448
rect 7637 2380 7759 2416
rect 7637 2348 7682 2380
rect 7682 2348 7714 2380
rect 7714 2348 7759 2380
rect 7637 2312 7759 2348
rect 7637 2280 7682 2312
rect 7682 2280 7714 2312
rect 7714 2280 7759 2312
rect 7637 2244 7759 2280
rect 7637 2212 7682 2244
rect 7682 2212 7714 2244
rect 7714 2212 7759 2244
rect 7637 2176 7759 2212
rect 7637 2144 7682 2176
rect 7682 2144 7714 2176
rect 7714 2144 7759 2176
rect 7637 2108 7759 2144
rect 7637 2076 7682 2108
rect 7682 2076 7714 2108
rect 7714 2076 7759 2108
rect 7637 2042 7759 2076
rect 7376 1776 7416 1810
rect 7376 1744 7380 1776
rect 7380 1744 7412 1776
rect 7412 1744 7416 1776
rect 7376 1708 7416 1744
rect 7376 1676 7380 1708
rect 7380 1676 7412 1708
rect 7412 1676 7416 1708
rect 7376 1640 7416 1676
rect 7376 1608 7380 1640
rect 7380 1608 7412 1640
rect 7412 1608 7416 1640
rect 7376 1572 7416 1608
rect 7376 1540 7380 1572
rect 7380 1540 7412 1572
rect 7412 1540 7416 1572
rect 7376 1504 7416 1540
rect 7376 1472 7380 1504
rect 7380 1472 7412 1504
rect 7412 1472 7416 1504
rect 7376 1436 7416 1472
rect 7376 1404 7380 1436
rect 7380 1404 7412 1436
rect 7412 1404 7416 1436
rect 7376 1368 7416 1404
rect 7376 1336 7380 1368
rect 7380 1336 7412 1368
rect 7412 1336 7416 1368
rect 7376 1300 7416 1336
rect 7376 1268 7380 1300
rect 7380 1268 7412 1300
rect 7412 1268 7416 1300
rect 7376 1232 7416 1268
rect 7376 1200 7380 1232
rect 7380 1200 7412 1232
rect 7412 1200 7416 1232
rect 7376 1164 7416 1200
rect 7376 1132 7380 1164
rect 7380 1132 7412 1164
rect 7412 1132 7416 1164
rect 7376 1096 7416 1132
rect 7376 1064 7380 1096
rect 7380 1064 7412 1096
rect 7412 1064 7416 1096
rect 7376 1028 7416 1064
rect 7376 996 7380 1028
rect 7380 996 7412 1028
rect 7412 996 7416 1028
rect 7376 960 7416 996
rect 7376 928 7380 960
rect 7380 928 7412 960
rect 7412 928 7416 960
rect 7376 892 7416 928
rect 7376 860 7380 892
rect 7380 860 7412 892
rect 7412 860 7416 892
rect 7376 824 7416 860
rect 7376 792 7380 824
rect 7380 792 7412 824
rect 7412 792 7416 824
rect 7376 756 7416 792
rect 7376 724 7380 756
rect 7380 724 7412 756
rect 7412 724 7416 756
rect 7376 688 7416 724
rect 7376 656 7380 688
rect 7380 656 7412 688
rect 7412 656 7416 688
rect 7376 622 7416 656
rect 7980 3196 8020 3230
rect 7980 3164 7984 3196
rect 7984 3164 8016 3196
rect 8016 3164 8020 3196
rect 7980 3128 8020 3164
rect 7980 3096 7984 3128
rect 7984 3096 8016 3128
rect 8016 3096 8020 3128
rect 7980 3060 8020 3096
rect 7980 3028 7984 3060
rect 7984 3028 8016 3060
rect 8016 3028 8020 3060
rect 7980 2992 8020 3028
rect 7980 2960 7984 2992
rect 7984 2960 8016 2992
rect 8016 2960 8020 2992
rect 7980 2924 8020 2960
rect 7980 2892 7984 2924
rect 7984 2892 8016 2924
rect 8016 2892 8020 2924
rect 7980 2856 8020 2892
rect 7980 2824 7984 2856
rect 7984 2824 8016 2856
rect 8016 2824 8020 2856
rect 7980 2788 8020 2824
rect 7980 2756 7984 2788
rect 7984 2756 8016 2788
rect 8016 2756 8020 2788
rect 7980 2720 8020 2756
rect 7980 2688 7984 2720
rect 7984 2688 8016 2720
rect 8016 2688 8020 2720
rect 7980 2652 8020 2688
rect 7980 2620 7984 2652
rect 7984 2620 8016 2652
rect 8016 2620 8020 2652
rect 7980 2584 8020 2620
rect 7980 2552 7984 2584
rect 7984 2552 8016 2584
rect 8016 2552 8020 2584
rect 7980 2516 8020 2552
rect 7980 2484 7984 2516
rect 7984 2484 8016 2516
rect 8016 2484 8020 2516
rect 7980 2448 8020 2484
rect 7980 2416 7984 2448
rect 7984 2416 8016 2448
rect 8016 2416 8020 2448
rect 7980 2380 8020 2416
rect 7980 2348 7984 2380
rect 7984 2348 8016 2380
rect 8016 2348 8020 2380
rect 7980 2312 8020 2348
rect 7980 2280 7984 2312
rect 7984 2280 8016 2312
rect 8016 2280 8020 2312
rect 7980 2244 8020 2280
rect 7980 2212 7984 2244
rect 7984 2212 8016 2244
rect 8016 2212 8020 2244
rect 7980 2176 8020 2212
rect 7980 2144 7984 2176
rect 7984 2144 8016 2176
rect 8016 2144 8020 2176
rect 7980 2108 8020 2144
rect 7980 2076 7984 2108
rect 7984 2076 8016 2108
rect 8016 2076 8020 2108
rect 7980 2042 8020 2076
rect 7637 1776 7759 1810
rect 7637 1744 7682 1776
rect 7682 1744 7714 1776
rect 7714 1744 7759 1776
rect 7637 1708 7759 1744
rect 7637 1676 7682 1708
rect 7682 1676 7714 1708
rect 7714 1676 7759 1708
rect 7637 1640 7759 1676
rect 7637 1608 7682 1640
rect 7682 1608 7714 1640
rect 7714 1608 7759 1640
rect 7637 1572 7759 1608
rect 7637 1540 7682 1572
rect 7682 1540 7714 1572
rect 7714 1540 7759 1572
rect 7637 1504 7759 1540
rect 7637 1472 7682 1504
rect 7682 1472 7714 1504
rect 7714 1472 7759 1504
rect 7637 1436 7759 1472
rect 7637 1404 7682 1436
rect 7682 1404 7714 1436
rect 7714 1404 7759 1436
rect 7637 1368 7759 1404
rect 7637 1336 7682 1368
rect 7682 1336 7714 1368
rect 7714 1336 7759 1368
rect 7637 1300 7759 1336
rect 7637 1268 7682 1300
rect 7682 1268 7714 1300
rect 7714 1268 7759 1300
rect 7637 1232 7759 1268
rect 7637 1200 7682 1232
rect 7682 1200 7714 1232
rect 7714 1200 7759 1232
rect 7637 1164 7759 1200
rect 7637 1132 7682 1164
rect 7682 1132 7714 1164
rect 7714 1132 7759 1164
rect 7637 1096 7759 1132
rect 7637 1064 7682 1096
rect 7682 1064 7714 1096
rect 7714 1064 7759 1096
rect 7637 1028 7759 1064
rect 7637 996 7682 1028
rect 7682 996 7714 1028
rect 7714 996 7759 1028
rect 7637 960 7759 996
rect 7637 928 7682 960
rect 7682 928 7714 960
rect 7714 928 7759 960
rect 7637 892 7759 928
rect 7637 860 7682 892
rect 7682 860 7714 892
rect 7714 860 7759 892
rect 7637 824 7759 860
rect 7637 792 7682 824
rect 7682 792 7714 824
rect 7714 792 7759 824
rect 7637 756 7759 792
rect 7637 724 7682 756
rect 7682 724 7714 756
rect 7714 724 7759 756
rect 7637 688 7759 724
rect 7637 656 7682 688
rect 7682 656 7714 688
rect 7714 656 7759 688
rect 7637 622 7759 656
rect 8241 3196 8363 3230
rect 8241 3164 8286 3196
rect 8286 3164 8318 3196
rect 8318 3164 8363 3196
rect 8241 3128 8363 3164
rect 8241 3096 8286 3128
rect 8286 3096 8318 3128
rect 8318 3096 8363 3128
rect 8241 3060 8363 3096
rect 8241 3028 8286 3060
rect 8286 3028 8318 3060
rect 8318 3028 8363 3060
rect 8241 2992 8363 3028
rect 8241 2960 8286 2992
rect 8286 2960 8318 2992
rect 8318 2960 8363 2992
rect 8241 2924 8363 2960
rect 8241 2892 8286 2924
rect 8286 2892 8318 2924
rect 8318 2892 8363 2924
rect 8241 2856 8363 2892
rect 8241 2824 8286 2856
rect 8286 2824 8318 2856
rect 8318 2824 8363 2856
rect 8241 2788 8363 2824
rect 8241 2756 8286 2788
rect 8286 2756 8318 2788
rect 8318 2756 8363 2788
rect 8241 2720 8363 2756
rect 8241 2688 8286 2720
rect 8286 2688 8318 2720
rect 8318 2688 8363 2720
rect 8241 2652 8363 2688
rect 8241 2620 8286 2652
rect 8286 2620 8318 2652
rect 8318 2620 8363 2652
rect 8241 2584 8363 2620
rect 8241 2552 8286 2584
rect 8286 2552 8318 2584
rect 8318 2552 8363 2584
rect 8241 2516 8363 2552
rect 8241 2484 8286 2516
rect 8286 2484 8318 2516
rect 8318 2484 8363 2516
rect 8241 2448 8363 2484
rect 8241 2416 8286 2448
rect 8286 2416 8318 2448
rect 8318 2416 8363 2448
rect 8241 2380 8363 2416
rect 8241 2348 8286 2380
rect 8286 2348 8318 2380
rect 8318 2348 8363 2380
rect 8241 2312 8363 2348
rect 8241 2280 8286 2312
rect 8286 2280 8318 2312
rect 8318 2280 8363 2312
rect 8241 2244 8363 2280
rect 8241 2212 8286 2244
rect 8286 2212 8318 2244
rect 8318 2212 8363 2244
rect 8241 2176 8363 2212
rect 8241 2144 8286 2176
rect 8286 2144 8318 2176
rect 8318 2144 8363 2176
rect 8241 2108 8363 2144
rect 8241 2076 8286 2108
rect 8286 2076 8318 2108
rect 8318 2076 8363 2108
rect 8241 2042 8363 2076
rect 7980 1776 8020 1810
rect 7980 1744 7984 1776
rect 7984 1744 8016 1776
rect 8016 1744 8020 1776
rect 7980 1708 8020 1744
rect 7980 1676 7984 1708
rect 7984 1676 8016 1708
rect 8016 1676 8020 1708
rect 7980 1640 8020 1676
rect 7980 1608 7984 1640
rect 7984 1608 8016 1640
rect 8016 1608 8020 1640
rect 7980 1572 8020 1608
rect 7980 1540 7984 1572
rect 7984 1540 8016 1572
rect 8016 1540 8020 1572
rect 7980 1504 8020 1540
rect 7980 1472 7984 1504
rect 7984 1472 8016 1504
rect 8016 1472 8020 1504
rect 7980 1436 8020 1472
rect 7980 1404 7984 1436
rect 7984 1404 8016 1436
rect 8016 1404 8020 1436
rect 7980 1368 8020 1404
rect 7980 1336 7984 1368
rect 7984 1336 8016 1368
rect 8016 1336 8020 1368
rect 7980 1300 8020 1336
rect 7980 1268 7984 1300
rect 7984 1268 8016 1300
rect 8016 1268 8020 1300
rect 7980 1232 8020 1268
rect 7980 1200 7984 1232
rect 7984 1200 8016 1232
rect 8016 1200 8020 1232
rect 7980 1164 8020 1200
rect 7980 1132 7984 1164
rect 7984 1132 8016 1164
rect 8016 1132 8020 1164
rect 7980 1096 8020 1132
rect 7980 1064 7984 1096
rect 7984 1064 8016 1096
rect 8016 1064 8020 1096
rect 7980 1028 8020 1064
rect 7980 996 7984 1028
rect 7984 996 8016 1028
rect 8016 996 8020 1028
rect 7980 960 8020 996
rect 7980 928 7984 960
rect 7984 928 8016 960
rect 8016 928 8020 960
rect 7980 892 8020 928
rect 7980 860 7984 892
rect 7984 860 8016 892
rect 8016 860 8020 892
rect 7980 824 8020 860
rect 7980 792 7984 824
rect 7984 792 8016 824
rect 8016 792 8020 824
rect 7980 756 8020 792
rect 7980 724 7984 756
rect 7984 724 8016 756
rect 8016 724 8020 756
rect 7980 688 8020 724
rect 7980 656 7984 688
rect 7984 656 8016 688
rect 8016 656 8020 688
rect 7980 622 8020 656
rect 8584 3196 8624 3230
rect 8584 3164 8588 3196
rect 8588 3164 8620 3196
rect 8620 3164 8624 3196
rect 8584 3128 8624 3164
rect 8584 3096 8588 3128
rect 8588 3096 8620 3128
rect 8620 3096 8624 3128
rect 8584 3060 8624 3096
rect 8584 3028 8588 3060
rect 8588 3028 8620 3060
rect 8620 3028 8624 3060
rect 8584 2992 8624 3028
rect 8584 2960 8588 2992
rect 8588 2960 8620 2992
rect 8620 2960 8624 2992
rect 8584 2924 8624 2960
rect 8584 2892 8588 2924
rect 8588 2892 8620 2924
rect 8620 2892 8624 2924
rect 8584 2856 8624 2892
rect 8584 2824 8588 2856
rect 8588 2824 8620 2856
rect 8620 2824 8624 2856
rect 8584 2788 8624 2824
rect 8584 2756 8588 2788
rect 8588 2756 8620 2788
rect 8620 2756 8624 2788
rect 8584 2720 8624 2756
rect 8584 2688 8588 2720
rect 8588 2688 8620 2720
rect 8620 2688 8624 2720
rect 8584 2652 8624 2688
rect 8584 2620 8588 2652
rect 8588 2620 8620 2652
rect 8620 2620 8624 2652
rect 8584 2584 8624 2620
rect 8584 2552 8588 2584
rect 8588 2552 8620 2584
rect 8620 2552 8624 2584
rect 8584 2516 8624 2552
rect 8584 2484 8588 2516
rect 8588 2484 8620 2516
rect 8620 2484 8624 2516
rect 8584 2448 8624 2484
rect 8584 2416 8588 2448
rect 8588 2416 8620 2448
rect 8620 2416 8624 2448
rect 8584 2380 8624 2416
rect 8584 2348 8588 2380
rect 8588 2348 8620 2380
rect 8620 2348 8624 2380
rect 8584 2312 8624 2348
rect 8584 2280 8588 2312
rect 8588 2280 8620 2312
rect 8620 2280 8624 2312
rect 8584 2244 8624 2280
rect 8584 2212 8588 2244
rect 8588 2212 8620 2244
rect 8620 2212 8624 2244
rect 8584 2176 8624 2212
rect 8584 2144 8588 2176
rect 8588 2144 8620 2176
rect 8620 2144 8624 2176
rect 8584 2108 8624 2144
rect 8584 2076 8588 2108
rect 8588 2076 8620 2108
rect 8620 2076 8624 2108
rect 8584 2042 8624 2076
rect 8241 1776 8363 1810
rect 8241 1744 8286 1776
rect 8286 1744 8318 1776
rect 8318 1744 8363 1776
rect 8241 1708 8363 1744
rect 8241 1676 8286 1708
rect 8286 1676 8318 1708
rect 8318 1676 8363 1708
rect 8241 1640 8363 1676
rect 8241 1608 8286 1640
rect 8286 1608 8318 1640
rect 8318 1608 8363 1640
rect 8241 1572 8363 1608
rect 8241 1540 8286 1572
rect 8286 1540 8318 1572
rect 8318 1540 8363 1572
rect 8241 1504 8363 1540
rect 8241 1472 8286 1504
rect 8286 1472 8318 1504
rect 8318 1472 8363 1504
rect 8241 1436 8363 1472
rect 8241 1404 8286 1436
rect 8286 1404 8318 1436
rect 8318 1404 8363 1436
rect 8241 1368 8363 1404
rect 8241 1336 8286 1368
rect 8286 1336 8318 1368
rect 8318 1336 8363 1368
rect 8241 1300 8363 1336
rect 8241 1268 8286 1300
rect 8286 1268 8318 1300
rect 8318 1268 8363 1300
rect 8241 1232 8363 1268
rect 8241 1200 8286 1232
rect 8286 1200 8318 1232
rect 8318 1200 8363 1232
rect 8241 1164 8363 1200
rect 8241 1132 8286 1164
rect 8286 1132 8318 1164
rect 8318 1132 8363 1164
rect 8241 1096 8363 1132
rect 8241 1064 8286 1096
rect 8286 1064 8318 1096
rect 8318 1064 8363 1096
rect 8241 1028 8363 1064
rect 8241 996 8286 1028
rect 8286 996 8318 1028
rect 8318 996 8363 1028
rect 8241 960 8363 996
rect 8241 928 8286 960
rect 8286 928 8318 960
rect 8318 928 8363 960
rect 8241 892 8363 928
rect 8241 860 8286 892
rect 8286 860 8318 892
rect 8318 860 8363 892
rect 8241 824 8363 860
rect 8241 792 8286 824
rect 8286 792 8318 824
rect 8318 792 8363 824
rect 8241 756 8363 792
rect 8241 724 8286 756
rect 8286 724 8318 756
rect 8318 724 8363 756
rect 8241 688 8363 724
rect 8241 656 8286 688
rect 8286 656 8318 688
rect 8318 656 8363 688
rect 8241 622 8363 656
rect 8845 3196 8967 3230
rect 8845 3164 8890 3196
rect 8890 3164 8922 3196
rect 8922 3164 8967 3196
rect 8845 3128 8967 3164
rect 8845 3096 8890 3128
rect 8890 3096 8922 3128
rect 8922 3096 8967 3128
rect 8845 3060 8967 3096
rect 8845 3028 8890 3060
rect 8890 3028 8922 3060
rect 8922 3028 8967 3060
rect 8845 2992 8967 3028
rect 8845 2960 8890 2992
rect 8890 2960 8922 2992
rect 8922 2960 8967 2992
rect 8845 2924 8967 2960
rect 8845 2892 8890 2924
rect 8890 2892 8922 2924
rect 8922 2892 8967 2924
rect 8845 2856 8967 2892
rect 8845 2824 8890 2856
rect 8890 2824 8922 2856
rect 8922 2824 8967 2856
rect 8845 2788 8967 2824
rect 8845 2756 8890 2788
rect 8890 2756 8922 2788
rect 8922 2756 8967 2788
rect 8845 2720 8967 2756
rect 8845 2688 8890 2720
rect 8890 2688 8922 2720
rect 8922 2688 8967 2720
rect 8845 2652 8967 2688
rect 8845 2620 8890 2652
rect 8890 2620 8922 2652
rect 8922 2620 8967 2652
rect 8845 2584 8967 2620
rect 8845 2552 8890 2584
rect 8890 2552 8922 2584
rect 8922 2552 8967 2584
rect 8845 2516 8967 2552
rect 8845 2484 8890 2516
rect 8890 2484 8922 2516
rect 8922 2484 8967 2516
rect 8845 2448 8967 2484
rect 8845 2416 8890 2448
rect 8890 2416 8922 2448
rect 8922 2416 8967 2448
rect 8845 2380 8967 2416
rect 8845 2348 8890 2380
rect 8890 2348 8922 2380
rect 8922 2348 8967 2380
rect 8845 2312 8967 2348
rect 8845 2280 8890 2312
rect 8890 2280 8922 2312
rect 8922 2280 8967 2312
rect 8845 2244 8967 2280
rect 8845 2212 8890 2244
rect 8890 2212 8922 2244
rect 8922 2212 8967 2244
rect 8845 2176 8967 2212
rect 8845 2144 8890 2176
rect 8890 2144 8922 2176
rect 8922 2144 8967 2176
rect 8845 2108 8967 2144
rect 8845 2076 8890 2108
rect 8890 2076 8922 2108
rect 8922 2076 8967 2108
rect 8845 2042 8967 2076
rect 8584 1776 8624 1810
rect 8584 1744 8588 1776
rect 8588 1744 8620 1776
rect 8620 1744 8624 1776
rect 8584 1708 8624 1744
rect 8584 1676 8588 1708
rect 8588 1676 8620 1708
rect 8620 1676 8624 1708
rect 8584 1640 8624 1676
rect 8584 1608 8588 1640
rect 8588 1608 8620 1640
rect 8620 1608 8624 1640
rect 8584 1572 8624 1608
rect 8584 1540 8588 1572
rect 8588 1540 8620 1572
rect 8620 1540 8624 1572
rect 8584 1504 8624 1540
rect 8584 1472 8588 1504
rect 8588 1472 8620 1504
rect 8620 1472 8624 1504
rect 8584 1436 8624 1472
rect 8584 1404 8588 1436
rect 8588 1404 8620 1436
rect 8620 1404 8624 1436
rect 8584 1368 8624 1404
rect 8584 1336 8588 1368
rect 8588 1336 8620 1368
rect 8620 1336 8624 1368
rect 8584 1300 8624 1336
rect 8584 1268 8588 1300
rect 8588 1268 8620 1300
rect 8620 1268 8624 1300
rect 8584 1232 8624 1268
rect 8584 1200 8588 1232
rect 8588 1200 8620 1232
rect 8620 1200 8624 1232
rect 8584 1164 8624 1200
rect 8584 1132 8588 1164
rect 8588 1132 8620 1164
rect 8620 1132 8624 1164
rect 8584 1096 8624 1132
rect 8584 1064 8588 1096
rect 8588 1064 8620 1096
rect 8620 1064 8624 1096
rect 8584 1028 8624 1064
rect 8584 996 8588 1028
rect 8588 996 8620 1028
rect 8620 996 8624 1028
rect 8584 960 8624 996
rect 8584 928 8588 960
rect 8588 928 8620 960
rect 8620 928 8624 960
rect 8584 892 8624 928
rect 8584 860 8588 892
rect 8588 860 8620 892
rect 8620 860 8624 892
rect 8584 824 8624 860
rect 8584 792 8588 824
rect 8588 792 8620 824
rect 8620 792 8624 824
rect 8584 756 8624 792
rect 8584 724 8588 756
rect 8588 724 8620 756
rect 8620 724 8624 756
rect 8584 688 8624 724
rect 8584 656 8588 688
rect 8588 656 8620 688
rect 8620 656 8624 688
rect 8584 622 8624 656
rect 9188 3196 9228 3230
rect 9188 3164 9192 3196
rect 9192 3164 9224 3196
rect 9224 3164 9228 3196
rect 9188 3128 9228 3164
rect 9188 3096 9192 3128
rect 9192 3096 9224 3128
rect 9224 3096 9228 3128
rect 9188 3060 9228 3096
rect 9188 3028 9192 3060
rect 9192 3028 9224 3060
rect 9224 3028 9228 3060
rect 9188 2992 9228 3028
rect 9188 2960 9192 2992
rect 9192 2960 9224 2992
rect 9224 2960 9228 2992
rect 9188 2924 9228 2960
rect 9188 2892 9192 2924
rect 9192 2892 9224 2924
rect 9224 2892 9228 2924
rect 9188 2856 9228 2892
rect 9188 2824 9192 2856
rect 9192 2824 9224 2856
rect 9224 2824 9228 2856
rect 9188 2788 9228 2824
rect 9188 2756 9192 2788
rect 9192 2756 9224 2788
rect 9224 2756 9228 2788
rect 9188 2720 9228 2756
rect 9188 2688 9192 2720
rect 9192 2688 9224 2720
rect 9224 2688 9228 2720
rect 9188 2652 9228 2688
rect 9188 2620 9192 2652
rect 9192 2620 9224 2652
rect 9224 2620 9228 2652
rect 9188 2584 9228 2620
rect 9188 2552 9192 2584
rect 9192 2552 9224 2584
rect 9224 2552 9228 2584
rect 9188 2516 9228 2552
rect 9188 2484 9192 2516
rect 9192 2484 9224 2516
rect 9224 2484 9228 2516
rect 9188 2448 9228 2484
rect 9188 2416 9192 2448
rect 9192 2416 9224 2448
rect 9224 2416 9228 2448
rect 9188 2380 9228 2416
rect 9188 2348 9192 2380
rect 9192 2348 9224 2380
rect 9224 2348 9228 2380
rect 9188 2312 9228 2348
rect 9188 2280 9192 2312
rect 9192 2280 9224 2312
rect 9224 2280 9228 2312
rect 9188 2244 9228 2280
rect 9188 2212 9192 2244
rect 9192 2212 9224 2244
rect 9224 2212 9228 2244
rect 9188 2176 9228 2212
rect 9188 2144 9192 2176
rect 9192 2144 9224 2176
rect 9224 2144 9228 2176
rect 9188 2108 9228 2144
rect 9188 2076 9192 2108
rect 9192 2076 9224 2108
rect 9224 2076 9228 2108
rect 9188 2042 9228 2076
rect 8845 1776 8967 1810
rect 8845 1744 8890 1776
rect 8890 1744 8922 1776
rect 8922 1744 8967 1776
rect 8845 1708 8967 1744
rect 8845 1676 8890 1708
rect 8890 1676 8922 1708
rect 8922 1676 8967 1708
rect 8845 1640 8967 1676
rect 8845 1608 8890 1640
rect 8890 1608 8922 1640
rect 8922 1608 8967 1640
rect 8845 1572 8967 1608
rect 8845 1540 8890 1572
rect 8890 1540 8922 1572
rect 8922 1540 8967 1572
rect 8845 1504 8967 1540
rect 8845 1472 8890 1504
rect 8890 1472 8922 1504
rect 8922 1472 8967 1504
rect 8845 1436 8967 1472
rect 8845 1404 8890 1436
rect 8890 1404 8922 1436
rect 8922 1404 8967 1436
rect 8845 1368 8967 1404
rect 8845 1336 8890 1368
rect 8890 1336 8922 1368
rect 8922 1336 8967 1368
rect 8845 1300 8967 1336
rect 8845 1268 8890 1300
rect 8890 1268 8922 1300
rect 8922 1268 8967 1300
rect 8845 1232 8967 1268
rect 8845 1200 8890 1232
rect 8890 1200 8922 1232
rect 8922 1200 8967 1232
rect 8845 1164 8967 1200
rect 8845 1132 8890 1164
rect 8890 1132 8922 1164
rect 8922 1132 8967 1164
rect 8845 1096 8967 1132
rect 8845 1064 8890 1096
rect 8890 1064 8922 1096
rect 8922 1064 8967 1096
rect 8845 1028 8967 1064
rect 8845 996 8890 1028
rect 8890 996 8922 1028
rect 8922 996 8967 1028
rect 8845 960 8967 996
rect 8845 928 8890 960
rect 8890 928 8922 960
rect 8922 928 8967 960
rect 8845 892 8967 928
rect 8845 860 8890 892
rect 8890 860 8922 892
rect 8922 860 8967 892
rect 8845 824 8967 860
rect 8845 792 8890 824
rect 8890 792 8922 824
rect 8922 792 8967 824
rect 8845 756 8967 792
rect 8845 724 8890 756
rect 8890 724 8922 756
rect 8922 724 8967 756
rect 8845 688 8967 724
rect 8845 656 8890 688
rect 8890 656 8922 688
rect 8922 656 8967 688
rect 8845 622 8967 656
rect 9188 1776 9228 1810
rect 9188 1744 9192 1776
rect 9192 1744 9224 1776
rect 9224 1744 9228 1776
rect 9188 1708 9228 1744
rect 9188 1676 9192 1708
rect 9192 1676 9224 1708
rect 9224 1676 9228 1708
rect 9188 1640 9228 1676
rect 9188 1608 9192 1640
rect 9192 1608 9224 1640
rect 9224 1608 9228 1640
rect 9188 1572 9228 1608
rect 9188 1540 9192 1572
rect 9192 1540 9224 1572
rect 9224 1540 9228 1572
rect 9188 1504 9228 1540
rect 9188 1472 9192 1504
rect 9192 1472 9224 1504
rect 9224 1472 9228 1504
rect 9188 1436 9228 1472
rect 9188 1404 9192 1436
rect 9192 1404 9224 1436
rect 9224 1404 9228 1436
rect 9188 1368 9228 1404
rect 9188 1336 9192 1368
rect 9192 1336 9224 1368
rect 9224 1336 9228 1368
rect 9188 1300 9228 1336
rect 9188 1268 9192 1300
rect 9192 1268 9224 1300
rect 9224 1268 9228 1300
rect 9188 1232 9228 1268
rect 9188 1200 9192 1232
rect 9192 1200 9224 1232
rect 9224 1200 9228 1232
rect 9188 1164 9228 1200
rect 9188 1132 9192 1164
rect 9192 1132 9224 1164
rect 9224 1132 9228 1164
rect 9188 1096 9228 1132
rect 9188 1064 9192 1096
rect 9192 1064 9224 1096
rect 9224 1064 9228 1096
rect 9188 1028 9228 1064
rect 9188 996 9192 1028
rect 9192 996 9224 1028
rect 9224 996 9228 1028
rect 9188 960 9228 996
rect 9188 928 9192 960
rect 9192 928 9224 960
rect 9224 928 9228 960
rect 9188 892 9228 928
rect 9188 860 9192 892
rect 9192 860 9224 892
rect 9224 860 9228 892
rect 9188 824 9228 860
rect 9188 792 9192 824
rect 9192 792 9224 824
rect 9224 792 9228 824
rect 9188 756 9228 792
rect 9188 724 9192 756
rect 9192 724 9224 756
rect 9224 724 9228 756
rect 9188 688 9228 724
rect 9188 656 9192 688
rect 9192 656 9224 688
rect 9224 656 9228 688
rect 9188 622 9228 656
rect 6772 410 6812 414
rect 7376 410 7416 414
rect 7980 410 8020 414
rect 8584 410 8624 414
rect 9188 410 9228 414
rect 6772 378 6794 410
rect 6794 378 6812 410
rect 7376 378 7406 410
rect 7406 378 7416 410
rect 7980 378 7982 410
rect 7982 378 8018 410
rect 8018 378 8020 410
rect 8584 378 8594 410
rect 8594 378 8624 410
rect 9188 378 9206 410
rect 9206 378 9228 410
rect 6772 374 6812 378
rect 7376 374 7416 378
rect 7980 374 8020 378
rect 8584 374 8624 378
rect 9188 374 9228 378
<< metal2 >>
rect 3575 3336 3615 3852
rect 3575 3205 3615 3214
rect 6772 3832 6812 3852
rect 7033 3230 7155 3852
rect 7033 1810 7155 2042
rect 7033 613 7155 622
rect 7376 3832 7416 3852
rect 6772 0 6812 20
rect 7637 3230 7759 3852
rect 7637 1810 7759 2042
rect 7637 613 7759 622
rect 7980 3832 8020 3852
rect 7376 0 7416 20
rect 8241 3230 8363 3852
rect 8241 1810 8363 2042
rect 8241 613 8363 622
rect 8584 3832 8624 3852
rect 7980 0 8020 20
rect 8845 3230 8967 3852
rect 8845 1810 8967 2042
rect 8845 613 8967 622
rect 9188 3832 9228 3852
rect 8584 0 8624 20
rect 9188 0 9228 20
<< via2 >>
rect 6772 3478 6812 3832
rect 6772 3438 6812 3478
rect 6772 3230 6812 3438
rect 6772 2042 6812 3230
rect 6772 1810 6812 2042
rect 6772 622 6812 1810
rect 6772 414 6812 622
rect 7376 3478 7416 3832
rect 7376 3438 7416 3478
rect 7376 3230 7416 3438
rect 7376 2042 7416 3230
rect 7376 1810 7416 2042
rect 7376 622 7416 1810
rect 6772 374 6812 414
rect 6772 20 6812 374
rect 7376 414 7416 622
rect 7980 3478 8020 3832
rect 7980 3438 8020 3478
rect 7980 3230 8020 3438
rect 7980 2042 8020 3230
rect 7980 1810 8020 2042
rect 7980 622 8020 1810
rect 7376 374 7416 414
rect 7376 20 7416 374
rect 7980 414 8020 622
rect 8584 3478 8624 3832
rect 8584 3438 8624 3478
rect 8584 3230 8624 3438
rect 8584 2042 8624 3230
rect 8584 1810 8624 2042
rect 8584 622 8624 1810
rect 7980 374 8020 414
rect 7980 20 8020 374
rect 8584 414 8624 622
rect 9188 3478 9228 3832
rect 9188 3438 9228 3478
rect 9188 3230 9228 3438
rect 9188 2042 9228 3230
rect 9188 1810 9228 2042
rect 9188 622 9228 1810
rect 8584 374 8624 414
rect 8584 20 8624 374
rect 9188 414 9228 622
rect 9188 374 9228 414
rect 9188 20 9228 374
<< metal3 >>
rect 6772 3832 6812 3841
rect 6772 11 6812 20
rect 7376 3832 7416 3841
rect 7376 11 7416 20
rect 7980 3832 8020 3841
rect 7980 11 8020 20
rect 8584 3832 8624 3841
rect 8584 11 8624 20
rect 9188 3832 9228 3841
rect 9188 11 9228 20
<< labels >>
flabel metal2 s 8845 613 8967 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
flabel metal2 s 8241 613 8363 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
rlabel metal2 s 3575 3205 3615 3852 4 gate
port 4 nsew
rlabel metal2 s 7033 613 7155 3852 4 pad
port 3 nsew
flabel metal2 s 7637 613 7759 3852 0 FreeSans 800 0 0 0 pad
port 3 nsew
rlabel comment s 34 34 34 34 4 sub!
flabel comment s 3596 3220 3596 3220 0 FreeSans 400 0 0 0 dpant
flabel metal1 s 1081 3424 1535 3492 0 FreeSans 800 0 0 0 iovdd
port 2 nsew
flabel metal1 s 1052 3784 1505 3852 0 FreeSans 800 0 0 0 iovss
port 1 nsew
<< properties >>
string device primitive
string GDS_END 36349708
string GDS_FILE sg13g2_io.gds
string GDS_START 36208426
<< end >>
