magic
tech ihp-sg13g2
timestamp 1752440150
<< error_p >>
rect -18 130 -13 135
rect 13 130 18 135
rect -23 125 23 130
rect -18 119 18 125
rect -23 114 23 119
rect -18 109 -13 114
rect 13 109 18 114
rect -52 93 -47 98
rect -41 93 -36 98
rect 36 93 41 98
rect 47 93 52 98
rect -57 88 -52 93
rect -36 88 -31 93
rect 31 88 36 93
rect 52 88 57 93
rect -57 -93 -52 -88
rect -36 -93 -31 -88
rect 31 -93 36 -88
rect 52 -93 57 -88
rect -52 -98 -47 -93
rect -41 -98 -36 -93
rect 36 -98 41 -93
rect 47 -98 52 -93
rect -18 -114 -13 -109
rect 13 -114 18 -109
rect -23 -119 23 -114
rect -18 -125 18 -119
rect -23 -130 23 -125
rect -18 -135 -13 -130
rect 13 -135 18 -130
<< hvnmos >>
rect -25 -100 25 100
<< hvndiff >>
rect -59 93 -25 100
rect -59 -93 -52 93
rect -36 -93 -25 93
rect -59 -100 -25 -93
rect 25 93 59 100
rect 25 -93 36 93
rect 52 -93 59 93
rect 25 -100 59 -93
<< hvndiffc >>
rect -52 -93 -36 93
rect 36 -93 52 93
<< psubdiff >>
rect -59 182 59 189
rect -59 166 -52 182
rect 52 166 59 182
rect -59 159 59 166
rect -59 -166 59 -159
rect -59 -182 -52 -166
rect 52 -182 59 -166
rect -59 -189 59 -182
<< psubdiffcont >>
rect -52 166 52 182
rect -52 -182 52 -166
<< poly >>
rect -25 130 25 137
rect -25 114 -18 130
rect 18 114 25 130
rect -25 100 25 114
rect -25 -114 25 -100
rect -25 -130 -18 -114
rect 18 -130 25 -114
rect -25 -137 25 -130
<< polycont >>
rect -18 114 18 130
rect -18 -130 18 -114
<< metal1 >>
rect -57 182 57 187
rect -57 166 -52 182
rect 52 166 57 182
rect -57 161 57 166
rect -57 -166 57 -161
rect -57 -182 -52 -166
rect 52 -182 57 -166
rect -57 -187 57 -182
<< properties >>
string gencell hvnmos
string library sg13g2_devstdin
string parameters w 2 l 0.5 nf 1 nx 1 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 0 grc 0 gtc 1 gbc 1
<< end >>
