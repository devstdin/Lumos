magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757240632
<< error_p >>
rect -1486 11980 -1476 11990
rect 1476 11980 1486 11990
rect -1496 11970 -1486 11980
rect 1486 11970 1496 11980
rect -1496 11948 -1486 11958
rect 1486 11948 1496 11958
rect -1486 11938 -1476 11948
rect 1476 11938 1486 11948
rect -1554 11906 -1544 11916
rect -1532 11906 -1522 11916
rect 1522 11906 1532 11916
rect 1544 11906 1554 11916
rect -1564 11896 -1554 11906
rect -1522 11896 -1512 11906
rect 1512 11896 1522 11906
rect 1554 11896 1564 11906
rect -1564 9934 -1554 9944
rect -1522 9934 -1512 9944
rect 1512 9934 1522 9944
rect 1554 9934 1564 9944
rect -1554 9924 -1544 9934
rect -1532 9924 -1522 9934
rect 1522 9924 1532 9934
rect 1544 9924 1554 9934
rect -1486 9892 -1476 9902
rect 1476 9892 1486 9902
rect -1496 9882 -1486 9892
rect 1486 9882 1496 9892
rect -1496 9860 -1486 9870
rect 1486 9860 1496 9870
rect -1486 9850 -1476 9860
rect 1476 9850 1486 9860
rect -1486 9796 -1476 9806
rect 1476 9796 1486 9806
rect -1496 9786 -1486 9796
rect 1486 9786 1496 9796
rect -1496 9764 -1486 9774
rect 1486 9764 1496 9774
rect -1486 9754 -1476 9764
rect 1476 9754 1486 9764
rect -1554 9722 -1544 9732
rect -1532 9722 -1522 9732
rect 1522 9722 1532 9732
rect 1544 9722 1554 9732
rect -1564 9712 -1554 9722
rect -1522 9712 -1512 9722
rect 1512 9712 1522 9722
rect 1554 9712 1564 9722
rect -1564 7750 -1554 7760
rect -1522 7750 -1512 7760
rect 1512 7750 1522 7760
rect 1554 7750 1564 7760
rect -1554 7740 -1544 7750
rect -1532 7740 -1522 7750
rect 1522 7740 1532 7750
rect 1544 7740 1554 7750
rect -1486 7708 -1476 7718
rect 1476 7708 1486 7718
rect -1496 7698 -1486 7708
rect 1486 7698 1496 7708
rect -1496 7676 -1486 7686
rect 1486 7676 1496 7686
rect -1486 7666 -1476 7676
rect 1476 7666 1486 7676
rect -1486 7612 -1476 7622
rect 1476 7612 1486 7622
rect -1496 7602 -1486 7612
rect 1486 7602 1496 7612
rect -1496 7580 -1486 7590
rect 1486 7580 1496 7590
rect -1486 7570 -1476 7580
rect 1476 7570 1486 7580
rect -1554 7538 -1544 7548
rect -1532 7538 -1522 7548
rect 1522 7538 1532 7548
rect 1544 7538 1554 7548
rect -1564 7528 -1554 7538
rect -1522 7528 -1512 7538
rect 1512 7528 1522 7538
rect 1554 7528 1564 7538
rect -1564 5566 -1554 5576
rect -1522 5566 -1512 5576
rect 1512 5566 1522 5576
rect 1554 5566 1564 5576
rect -1554 5556 -1544 5566
rect -1532 5556 -1522 5566
rect 1522 5556 1532 5566
rect 1544 5556 1554 5566
rect -1486 5524 -1476 5534
rect 1476 5524 1486 5534
rect -1496 5514 -1486 5524
rect 1486 5514 1496 5524
rect -1496 5492 -1486 5502
rect 1486 5492 1496 5502
rect -1486 5482 -1476 5492
rect 1476 5482 1486 5492
rect -1486 5428 -1476 5438
rect 1476 5428 1486 5438
rect -1496 5418 -1486 5428
rect 1486 5418 1496 5428
rect -1496 5396 -1486 5406
rect 1486 5396 1496 5406
rect -1486 5386 -1476 5396
rect 1476 5386 1486 5396
rect -1554 5354 -1544 5364
rect -1532 5354 -1522 5364
rect 1522 5354 1532 5364
rect 1544 5354 1554 5364
rect -1564 5344 -1554 5354
rect -1522 5344 -1512 5354
rect 1512 5344 1522 5354
rect 1554 5344 1564 5354
rect -1564 3382 -1554 3392
rect -1522 3382 -1512 3392
rect 1512 3382 1522 3392
rect 1554 3382 1564 3392
rect -1554 3372 -1544 3382
rect -1532 3372 -1522 3382
rect 1522 3372 1532 3382
rect 1544 3372 1554 3382
rect -1486 3340 -1476 3350
rect 1476 3340 1486 3350
rect -1496 3330 -1486 3340
rect 1486 3330 1496 3340
rect -1496 3308 -1486 3318
rect 1486 3308 1496 3318
rect -1486 3298 -1476 3308
rect 1476 3298 1486 3308
rect -1486 3244 -1476 3254
rect 1476 3244 1486 3254
rect -1496 3234 -1486 3244
rect 1486 3234 1496 3244
rect -1496 3212 -1486 3222
rect 1486 3212 1496 3222
rect -1486 3202 -1476 3212
rect 1476 3202 1486 3212
rect -1554 3170 -1544 3180
rect -1532 3170 -1522 3180
rect 1522 3170 1532 3180
rect 1544 3170 1554 3180
rect -1564 3160 -1554 3170
rect -1522 3160 -1512 3170
rect 1512 3160 1522 3170
rect 1554 3160 1564 3170
rect -1564 1198 -1554 1208
rect -1522 1198 -1512 1208
rect 1512 1198 1522 1208
rect 1554 1198 1564 1208
rect -1554 1188 -1544 1198
rect -1532 1188 -1522 1198
rect 1522 1188 1532 1198
rect 1544 1188 1554 1198
rect -1486 1156 -1476 1166
rect 1476 1156 1486 1166
rect -1496 1146 -1486 1156
rect 1486 1146 1496 1156
rect -1496 1124 -1486 1134
rect 1486 1124 1496 1134
rect -1486 1114 -1476 1124
rect 1476 1114 1486 1124
rect -1486 1060 -1476 1070
rect 1476 1060 1486 1070
rect -1496 1050 -1486 1060
rect 1486 1050 1496 1060
rect -1496 1028 -1486 1038
rect 1486 1028 1496 1038
rect -1486 1018 -1476 1028
rect 1476 1018 1486 1028
rect -1554 986 -1544 996
rect -1532 986 -1522 996
rect 1522 986 1532 996
rect 1544 986 1554 996
rect -1564 976 -1554 986
rect -1522 976 -1512 986
rect 1512 976 1522 986
rect 1554 976 1564 986
rect -1564 -986 -1554 -976
rect -1522 -986 -1512 -976
rect 1512 -986 1522 -976
rect 1554 -986 1564 -976
rect -1554 -996 -1544 -986
rect -1532 -996 -1522 -986
rect 1522 -996 1532 -986
rect 1544 -996 1554 -986
rect -1486 -1028 -1476 -1018
rect 1476 -1028 1486 -1018
rect -1496 -1038 -1486 -1028
rect 1486 -1038 1496 -1028
rect -1496 -1060 -1486 -1050
rect 1486 -1060 1496 -1050
rect -1486 -1070 -1476 -1060
rect 1476 -1070 1486 -1060
<< nwell >>
rect -1878 -1074 1878 12229
rect -1692 -1124 1692 -1074
<< hvpmos >>
rect -1500 9920 1500 11920
rect -1500 7736 1500 9736
rect -1500 5552 1500 7552
rect -1500 3368 1500 5368
rect -1500 1184 1500 3184
rect -1500 -1000 1500 1000
<< hvpdiff >>
rect -1568 11906 -1500 11920
rect -1568 9934 -1554 11906
rect -1522 9934 -1500 11906
rect -1568 9920 -1500 9934
rect 1500 11906 1568 11920
rect 1500 9934 1522 11906
rect 1554 9934 1568 11906
rect 1500 9920 1568 9934
rect -1568 9722 -1500 9736
rect -1568 7750 -1554 9722
rect -1522 7750 -1500 9722
rect -1568 7736 -1500 7750
rect 1500 9722 1568 9736
rect 1500 7750 1522 9722
rect 1554 7750 1568 9722
rect 1500 7736 1568 7750
rect -1568 7538 -1500 7552
rect -1568 5566 -1554 7538
rect -1522 5566 -1500 7538
rect -1568 5552 -1500 5566
rect 1500 7538 1568 7552
rect 1500 5566 1522 7538
rect 1554 5566 1568 7538
rect 1500 5552 1568 5566
rect -1568 5354 -1500 5368
rect -1568 3382 -1554 5354
rect -1522 3382 -1500 5354
rect -1568 3368 -1500 3382
rect 1500 5354 1568 5368
rect 1500 3382 1522 5354
rect 1554 3382 1568 5354
rect 1500 3368 1568 3382
rect -1568 3170 -1500 3184
rect -1568 1198 -1554 3170
rect -1522 1198 -1500 3170
rect -1568 1184 -1500 1198
rect 1500 3170 1568 3184
rect 1500 1198 1522 3170
rect 1554 1198 1568 3170
rect 1500 1184 1568 1198
rect -1568 986 -1500 1000
rect -1568 -986 -1554 986
rect -1522 -986 -1500 986
rect -1568 -1000 -1500 -986
rect 1500 986 1568 1000
rect 1500 -986 1522 986
rect 1554 -986 1568 986
rect 1500 -1000 1568 -986
<< hvpdiffc >>
rect -1554 9934 -1522 11906
rect 1522 9934 1554 11906
rect -1554 7750 -1522 9722
rect 1522 7750 1554 9722
rect -1554 5566 -1522 7538
rect 1522 5566 1554 7538
rect -1554 3382 -1522 5354
rect 1522 3382 1554 5354
rect -1554 1198 -1522 3170
rect 1522 1198 1554 3170
rect -1554 -986 -1522 986
rect 1522 -986 1554 986
<< nsubdiff >>
rect -1754 12091 1754 12105
rect -1754 12059 -1680 12091
rect 1680 12059 1754 12091
rect -1754 12045 1754 12059
rect -1754 12031 -1694 12045
rect -1754 -936 -1740 12031
rect -1708 -936 -1694 12031
rect 1694 12031 1754 12045
rect -1754 -950 -1694 -936
rect 1694 -936 1708 12031
rect 1740 -936 1754 12031
rect 1694 -950 1754 -936
<< nsubdiffcont >>
rect -1680 12059 1680 12091
rect -1740 -936 -1708 12031
rect 1708 -936 1740 12031
<< poly >>
rect -1500 11980 1500 11994
rect -1500 11948 -1486 11980
rect 1486 11948 1500 11980
rect -1500 11920 1500 11948
rect -1500 9892 1500 9920
rect -1500 9860 -1486 9892
rect 1486 9860 1500 9892
rect -1500 9846 1500 9860
rect -1500 9796 1500 9810
rect -1500 9764 -1486 9796
rect 1486 9764 1500 9796
rect -1500 9736 1500 9764
rect -1500 7708 1500 7736
rect -1500 7676 -1486 7708
rect 1486 7676 1500 7708
rect -1500 7662 1500 7676
rect -1500 7612 1500 7626
rect -1500 7580 -1486 7612
rect 1486 7580 1500 7612
rect -1500 7552 1500 7580
rect -1500 5524 1500 5552
rect -1500 5492 -1486 5524
rect 1486 5492 1500 5524
rect -1500 5478 1500 5492
rect -1500 5428 1500 5442
rect -1500 5396 -1486 5428
rect 1486 5396 1500 5428
rect -1500 5368 1500 5396
rect -1500 3340 1500 3368
rect -1500 3308 -1486 3340
rect 1486 3308 1500 3340
rect -1500 3294 1500 3308
rect -1500 3244 1500 3258
rect -1500 3212 -1486 3244
rect 1486 3212 1500 3244
rect -1500 3184 1500 3212
rect -1500 1156 1500 1184
rect -1500 1124 -1486 1156
rect 1486 1124 1500 1156
rect -1500 1110 1500 1124
rect -1500 1060 1500 1074
rect -1500 1028 -1486 1060
rect 1486 1028 1500 1060
rect -1500 1000 1500 1028
rect -1500 -1028 1500 -1000
rect -1500 -1060 -1486 -1028
rect 1486 -1060 1500 -1028
rect -1500 -1074 1500 -1060
<< polycont >>
rect -1486 11948 1486 11980
rect -1486 9860 1486 9892
rect -1486 9764 1486 9796
rect -1486 7676 1486 7708
rect -1486 7580 1486 7612
rect -1486 5492 1486 5524
rect -1486 5396 1486 5428
rect -1486 3308 1486 3340
rect -1486 3212 1486 3244
rect -1486 1124 1486 1156
rect -1486 1028 1486 1060
rect -1486 -1060 1486 -1028
<< metal1 >>
rect -1750 12091 1750 12101
rect -1750 12059 -1680 12091
rect 1680 12059 1750 12091
rect -1750 12049 1750 12059
rect -1750 12031 -1698 12049
rect -1750 -936 -1740 12031
rect -1708 -936 -1698 12031
rect 1698 12031 1750 12049
rect -1750 -946 -1698 -936
rect 1698 -936 1708 12031
rect 1740 -936 1750 12031
rect 1698 -946 1750 -936
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 10 l 15 nf 1 nx 1 dx 0.21 ny 6 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.1666 glc 1 grc 1 gtc 1 gbc 0
<< end >>
