magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -2005 2604 4524
<< nwell >>
rect -124 1152 604 2524
<< pwell >>
rect -5 107 315 1054
rect -5 -5 485 107
<< nmos >>
rect 89 242 115 1028
rect 191 242 217 1028
<< pmos >>
rect 89 1276 115 2158
rect 191 1276 217 2158
<< ndiff >>
rect 21 288 89 1028
rect 21 256 35 288
rect 67 256 89 288
rect 21 242 89 256
rect 115 242 191 1028
rect 217 999 289 1028
rect 217 967 243 999
rect 275 967 289 999
rect 217 931 289 967
rect 217 899 243 931
rect 275 899 289 931
rect 217 863 289 899
rect 217 831 243 863
rect 275 831 289 863
rect 217 795 289 831
rect 217 763 243 795
rect 275 763 289 795
rect 217 727 289 763
rect 217 695 243 727
rect 275 695 289 727
rect 217 659 289 695
rect 217 627 243 659
rect 275 627 289 659
rect 217 591 289 627
rect 217 559 243 591
rect 275 559 289 591
rect 217 523 289 559
rect 217 491 243 523
rect 275 491 289 523
rect 217 455 289 491
rect 217 423 243 455
rect 275 423 289 455
rect 217 387 289 423
rect 217 355 243 387
rect 275 355 289 387
rect 217 242 289 355
<< pdiff >>
rect 21 2144 89 2158
rect 21 2112 35 2144
rect 67 2112 89 2144
rect 21 1276 89 2112
rect 115 2031 191 2158
rect 115 1999 137 2031
rect 169 1999 191 2031
rect 115 1963 191 1999
rect 115 1931 137 1963
rect 169 1931 191 1963
rect 115 1895 191 1931
rect 115 1863 137 1895
rect 169 1863 191 1895
rect 115 1827 191 1863
rect 115 1795 137 1827
rect 169 1795 191 1827
rect 115 1759 191 1795
rect 115 1727 137 1759
rect 169 1727 191 1759
rect 115 1691 191 1727
rect 115 1659 137 1691
rect 169 1659 191 1691
rect 115 1623 191 1659
rect 115 1591 137 1623
rect 169 1591 191 1623
rect 115 1555 191 1591
rect 115 1523 137 1555
rect 169 1523 191 1555
rect 115 1487 191 1523
rect 115 1455 137 1487
rect 169 1455 191 1487
rect 115 1419 191 1455
rect 115 1387 137 1419
rect 169 1387 191 1419
rect 115 1351 191 1387
rect 115 1319 137 1351
rect 169 1319 191 1351
rect 115 1276 191 1319
rect 217 2144 289 2158
rect 217 2112 243 2144
rect 275 2112 289 2144
rect 217 1276 289 2112
<< ndiffc >>
rect 35 256 67 288
rect 243 967 275 999
rect 243 899 275 931
rect 243 831 275 863
rect 243 763 275 795
rect 243 695 275 727
rect 243 627 275 659
rect 243 559 275 591
rect 243 491 275 523
rect 243 423 275 455
rect 243 355 275 387
<< pdiffc >>
rect 35 2112 67 2144
rect 137 1999 169 2031
rect 137 1931 169 1963
rect 137 1863 169 1895
rect 137 1795 169 1827
rect 137 1727 169 1759
rect 137 1659 169 1691
rect 137 1591 169 1623
rect 137 1523 169 1555
rect 137 1455 169 1487
rect 137 1387 169 1419
rect 137 1319 169 1351
rect 243 2112 275 2144
<< psubdiff >>
rect 21 67 459 81
rect 21 35 54 67
rect 86 35 122 67
rect 154 35 190 67
rect 222 35 258 67
rect 290 35 326 67
rect 358 35 394 67
rect 426 35 459 67
rect 21 21 459 35
<< nsubdiff >>
rect 21 2365 459 2379
rect 21 2333 54 2365
rect 86 2333 122 2365
rect 154 2333 190 2365
rect 222 2333 258 2365
rect 290 2333 326 2365
rect 358 2333 394 2365
rect 426 2333 459 2365
rect 21 2319 459 2333
<< psubdiffcont >>
rect 54 35 86 67
rect 122 35 154 67
rect 190 35 222 67
rect 258 35 290 67
rect 326 35 358 67
rect 394 35 426 67
<< nsubdiffcont >>
rect 54 2333 86 2365
rect 122 2333 154 2365
rect 190 2333 222 2365
rect 258 2333 290 2365
rect 326 2333 358 2365
rect 394 2333 426 2365
<< poly >>
rect 89 2158 115 2194
rect 191 2158 217 2194
rect 89 1182 115 1276
rect 191 1182 217 1276
rect 21 1168 115 1182
rect 21 1136 35 1168
rect 67 1136 115 1168
rect 21 1122 115 1136
rect 151 1168 217 1182
rect 151 1136 165 1168
rect 197 1136 217 1168
rect 151 1122 217 1136
rect 89 1028 115 1122
rect 191 1028 217 1122
rect 89 206 115 242
rect 191 206 217 242
<< polycont >>
rect 35 1136 67 1168
rect 165 1136 197 1168
<< metal1 >>
rect 0 2365 480 2400
rect 0 2333 54 2365
rect 86 2333 122 2365
rect 154 2333 190 2365
rect 222 2333 258 2365
rect 290 2333 326 2365
rect 358 2333 394 2365
rect 426 2333 480 2365
rect 0 2144 480 2333
rect 0 2112 35 2144
rect 67 2112 243 2144
rect 275 2112 480 2144
rect 30 1168 72 2076
rect 137 2031 280 2076
rect 169 1999 280 2031
rect 137 1963 280 1999
rect 169 1931 280 1963
rect 137 1895 280 1931
rect 169 1863 280 1895
rect 137 1827 280 1863
rect 169 1795 280 1827
rect 137 1759 280 1795
rect 169 1727 280 1759
rect 137 1691 280 1727
rect 169 1659 280 1691
rect 137 1623 280 1659
rect 169 1591 280 1623
rect 137 1555 280 1591
rect 169 1523 280 1555
rect 137 1487 280 1523
rect 169 1455 280 1487
rect 137 1419 280 1455
rect 169 1387 280 1419
rect 137 1351 280 1387
rect 169 1319 280 1351
rect 137 1303 280 1319
rect 30 1136 35 1168
rect 67 1136 72 1168
rect 30 324 72 1136
rect 160 1168 202 1267
rect 160 1136 165 1168
rect 197 1136 202 1168
rect 160 324 202 1136
rect 238 999 280 1303
rect 238 967 243 999
rect 275 967 280 999
rect 238 931 280 967
rect 238 899 243 931
rect 275 899 280 931
rect 238 863 280 899
rect 238 831 243 863
rect 275 831 280 863
rect 238 795 280 831
rect 238 763 243 795
rect 275 763 280 795
rect 238 727 280 763
rect 238 695 243 727
rect 275 695 280 727
rect 238 659 280 695
rect 238 627 243 659
rect 275 627 280 659
rect 238 591 280 627
rect 238 559 243 591
rect 275 559 280 591
rect 238 523 280 559
rect 238 491 243 523
rect 275 491 280 523
rect 238 455 280 491
rect 238 423 243 455
rect 275 423 280 455
rect 238 387 280 423
rect 238 355 243 387
rect 275 355 280 387
rect 238 324 280 355
rect 0 256 35 288
rect 67 256 480 288
rect 0 67 480 256
rect 0 35 54 67
rect 86 35 122 67
rect 154 35 190 67
rect 222 35 258 67
rect 290 35 326 67
rect 358 35 394 67
rect 426 35 480 67
rect 0 0 480 35
<< labels >>
flabel metal1 s 238 324 280 2076 0 FreeSans 800 0 0 0 nq
port 3 nsew
flabel metal1 s 160 324 202 1267 0 FreeSans 800 0 0 0 i1
port 5 nsew
rlabel metal1 s 30 324 72 2076 4 i0
port 4 nsew
rlabel metal1 s 0 2112 480 2400 4 vdd
port 1 nsew
rlabel metal1 s 0 0 480 288 4 vss
port 2 nsew
flabel comment s 72 58 72 58 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 22706678
string GDS_FILE sg13g2_io.gds
string GDS_START 22702576
<< end >>
