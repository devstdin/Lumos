magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 6 56 570 270
rect -26 -56 602 56
<< nmos >>
rect 101 96 127 244
rect 202 96 228 244
rect 372 96 398 244
rect 450 96 476 244
<< pmos >>
rect 101 436 127 660
rect 224 436 250 660
rect 326 436 352 660
rect 450 436 476 660
<< ndiff >>
rect 32 210 101 244
rect 32 178 46 210
rect 78 178 101 210
rect 32 142 101 178
rect 32 110 46 142
rect 78 110 101 142
rect 32 96 101 110
rect 127 96 202 244
rect 228 210 372 244
rect 228 178 250 210
rect 282 178 318 210
rect 350 178 372 210
rect 228 96 372 178
rect 398 96 450 244
rect 476 210 544 244
rect 476 178 498 210
rect 530 178 544 210
rect 476 142 544 178
rect 476 110 498 142
rect 530 110 544 142
rect 476 96 544 110
<< pdiff >>
rect 33 646 101 660
rect 33 614 47 646
rect 79 614 101 646
rect 33 578 101 614
rect 33 546 47 578
rect 79 546 101 578
rect 33 502 101 546
rect 33 470 47 502
rect 79 470 101 502
rect 33 436 101 470
rect 127 646 224 660
rect 127 614 170 646
rect 202 614 224 646
rect 127 578 224 614
rect 127 546 170 578
rect 202 546 224 578
rect 127 436 224 546
rect 250 570 326 660
rect 250 538 272 570
rect 304 538 326 570
rect 250 502 326 538
rect 250 470 272 502
rect 304 470 326 502
rect 250 436 326 470
rect 352 646 450 660
rect 352 614 374 646
rect 406 614 450 646
rect 352 578 450 614
rect 352 546 374 578
rect 406 546 450 578
rect 352 436 450 546
rect 476 646 544 660
rect 476 614 498 646
rect 530 614 544 646
rect 476 578 544 614
rect 476 546 498 578
rect 530 546 544 578
rect 476 502 544 546
rect 476 470 498 502
rect 530 470 544 502
rect 476 436 544 470
<< ndiffc >>
rect 46 178 78 210
rect 46 110 78 142
rect 250 178 282 210
rect 318 178 350 210
rect 498 178 530 210
rect 498 110 530 142
<< pdiffc >>
rect 47 614 79 646
rect 47 546 79 578
rect 47 470 79 502
rect 170 614 202 646
rect 170 546 202 578
rect 272 538 304 570
rect 272 470 304 502
rect 374 614 406 646
rect 374 546 406 578
rect 498 614 530 646
rect 498 546 530 578
rect 498 470 530 502
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 101 660 127 696
rect 224 660 250 696
rect 326 660 352 696
rect 450 660 476 696
rect 101 422 127 436
rect 34 408 127 422
rect 224 418 250 436
rect 34 376 48 408
rect 80 396 127 408
rect 190 404 250 418
rect 80 376 95 396
rect 34 362 95 376
rect 190 372 204 404
rect 236 372 250 404
rect 326 414 352 436
rect 450 414 476 436
rect 326 400 414 414
rect 326 380 368 400
rect 190 350 250 372
rect 140 326 250 350
rect 101 322 250 326
rect 286 368 368 380
rect 400 368 414 400
rect 286 354 414 368
rect 450 400 544 414
rect 450 368 498 400
rect 530 368 544 400
rect 450 354 544 368
rect 101 298 166 322
rect 101 244 127 298
rect 286 286 312 354
rect 202 258 312 286
rect 354 304 414 318
rect 354 272 368 304
rect 400 272 414 304
rect 354 258 414 272
rect 202 244 228 258
rect 372 244 398 258
rect 450 244 476 354
rect 101 60 127 96
rect 202 60 228 96
rect 372 60 398 96
rect 450 60 476 96
<< polycont >>
rect 48 376 80 408
rect 204 372 236 404
rect 368 368 400 400
rect 498 368 530 400
rect 368 272 400 304
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 36 646 90 712
rect 36 614 47 646
rect 79 614 90 646
rect 36 578 90 614
rect 36 546 47 578
rect 79 546 90 578
rect 36 502 90 546
rect 160 646 416 656
rect 160 614 170 646
rect 202 617 374 646
rect 202 614 212 617
rect 160 578 212 614
rect 364 614 374 617
rect 406 614 416 646
rect 160 546 170 578
rect 202 546 212 578
rect 160 536 212 546
rect 262 570 320 580
rect 262 538 272 570
rect 304 538 320 570
rect 36 470 47 502
rect 79 470 90 502
rect 36 460 90 470
rect 262 502 320 538
rect 364 578 416 614
rect 364 546 374 578
rect 406 546 416 578
rect 364 536 416 546
rect 488 646 540 712
rect 488 614 498 646
rect 530 614 540 646
rect 488 578 540 614
rect 488 546 498 578
rect 530 546 540 578
rect 262 470 272 502
rect 304 470 320 502
rect 488 502 540 546
rect 262 460 320 470
rect 164 414 223 451
rect 34 408 128 414
rect 34 376 48 408
rect 80 376 128 408
rect 34 312 128 376
rect 164 404 248 414
rect 164 372 204 404
rect 236 372 248 404
rect 164 357 248 372
rect 84 298 128 312
rect 84 266 156 298
rect 36 210 88 220
rect 36 178 46 210
rect 78 178 88 210
rect 36 142 88 178
rect 36 110 46 142
rect 78 110 88 142
rect 36 44 88 110
rect 124 128 156 266
rect 284 220 320 460
rect 356 400 416 488
rect 488 470 498 502
rect 530 470 540 502
rect 488 460 540 470
rect 356 368 368 400
rect 400 368 416 400
rect 356 354 416 368
rect 454 400 544 414
rect 454 368 498 400
rect 530 368 544 400
rect 358 304 418 312
rect 358 272 368 304
rect 400 272 418 304
rect 358 266 418 272
rect 454 266 544 368
rect 250 210 350 220
rect 282 178 318 210
rect 250 168 350 178
rect 386 128 418 266
rect 124 96 418 128
rect 488 210 540 220
rect 488 178 498 210
rect 530 178 540 210
rect 488 142 540 178
rect 488 110 498 142
rect 530 110 540 142
rect 488 44 540 110
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 262 460 320 580 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 454 266 544 414 0 FreeSans 400 0 0 0 A2
port 3 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 164 357 223 451 0 FreeSans 400 0 0 0 B1
port 5 nsew
flabel metal1 s 34 312 128 414 0 FreeSans 400 0 0 0 A1
port 6 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 7 nsew
flabel metal1 s 356 354 416 488 0 FreeSans 400 0 0 0 B2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 212220
string GDS_FILE 6_final.gds
string GDS_START 207146
<< end >>
