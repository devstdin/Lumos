magic
tech ihp-sg13g2
timestamp 1749470838
<< error_p >>
rect -18 536 -13 541
rect 13 536 18 541
rect 50 536 55 541
rect 81 536 86 541
rect 118 536 123 541
rect 149 536 154 541
rect 186 536 191 541
rect 217 536 222 541
rect 254 536 259 541
rect 285 536 290 541
rect -23 531 23 536
rect 45 531 91 536
rect 113 531 159 536
rect 181 531 227 536
rect 249 531 295 536
rect -18 525 18 531
rect 50 525 86 531
rect 118 525 154 531
rect 186 525 222 531
rect 254 525 290 531
rect -23 520 23 525
rect 45 520 91 525
rect 113 520 159 525
rect 181 520 227 525
rect 249 520 295 525
rect -18 515 -13 520
rect 13 515 18 520
rect 50 515 55 520
rect 81 515 86 520
rect 118 515 123 520
rect 149 515 154 520
rect 186 515 191 520
rect 217 515 222 520
rect 254 515 259 520
rect 285 515 290 520
rect -18 -520 -13 -515
rect 13 -520 18 -515
rect 50 -520 55 -515
rect 81 -520 86 -515
rect 118 -520 123 -515
rect 149 -520 154 -515
rect 186 -520 191 -515
rect 217 -520 222 -515
rect 254 -520 259 -515
rect 285 -520 290 -515
rect -23 -525 23 -520
rect 45 -525 91 -520
rect 113 -525 159 -520
rect 181 -525 227 -520
rect 249 -525 295 -520
rect -18 -531 18 -525
rect 50 -531 86 -525
rect 118 -531 154 -525
rect 186 -531 222 -525
rect 254 -531 290 -525
rect -23 -536 23 -531
rect 45 -536 91 -531
rect 113 -536 159 -531
rect 181 -536 227 -531
rect 249 -536 295 -531
rect -18 -541 -13 -536
rect 13 -541 18 -536
rect 50 -541 55 -536
rect 81 -541 86 -536
rect 118 -541 123 -536
rect 149 -541 154 -536
rect 186 -541 191 -536
rect 217 -541 222 -536
rect 254 -541 259 -536
rect 285 -541 290 -536
<< psubdiff >>
rect -115 626 387 633
rect -115 610 -78 626
rect 350 610 387 626
rect -115 603 387 610
rect -115 596 -85 603
rect -115 -596 -108 596
rect -92 -596 -85 596
rect 357 596 387 603
rect -115 -603 -85 -596
rect 357 -596 364 596
rect 380 -596 387 596
rect 357 -603 387 -596
rect -115 -610 387 -603
rect -115 -626 -78 -610
rect 350 -626 387 -610
rect -115 -633 387 -626
<< psubdiffcont >>
rect -78 610 350 626
rect -108 -596 -92 596
rect 364 -596 380 596
rect -78 -626 350 -610
<< poly >>
rect -25 536 25 543
rect -25 520 -18 536
rect 18 520 25 536
rect -25 500 25 520
rect -25 -520 25 -500
rect -25 -536 -18 -520
rect 18 -536 25 -520
rect -25 -543 25 -536
rect 43 536 93 543
rect 43 520 50 536
rect 86 520 93 536
rect 43 500 93 520
rect 43 -520 93 -500
rect 43 -536 50 -520
rect 86 -536 93 -520
rect 43 -543 93 -536
rect 111 536 161 543
rect 111 520 118 536
rect 154 520 161 536
rect 111 500 161 520
rect 111 -520 161 -500
rect 111 -536 118 -520
rect 154 -536 161 -520
rect 111 -543 161 -536
rect 179 536 229 543
rect 179 520 186 536
rect 222 520 229 536
rect 179 500 229 520
rect 179 -520 229 -500
rect 179 -536 186 -520
rect 222 -536 229 -520
rect 179 -543 229 -536
rect 247 536 297 543
rect 247 520 254 536
rect 290 520 297 536
rect 247 500 297 520
rect 247 -520 297 -500
rect 247 -536 254 -520
rect 290 -536 297 -520
rect 247 -543 297 -536
<< polycont >>
rect -18 520 18 536
rect -18 -536 18 -520
rect 50 520 86 536
rect 50 -536 86 -520
rect 118 520 154 536
rect 118 -536 154 -520
rect 186 520 222 536
rect 186 -536 222 -520
rect 254 520 290 536
rect 254 -536 290 -520
<< xpolyres >>
rect -25 -500 25 500
rect 43 -500 93 500
rect 111 -500 161 500
rect 179 -500 229 500
rect 247 -500 297 500
<< metal1 >>
rect -113 626 385 631
rect -113 610 -78 626
rect 350 610 385 626
rect -113 605 385 610
rect -113 596 -87 605
rect -113 -596 -108 596
rect -92 -596 -87 596
rect 359 596 385 605
rect -113 -605 -87 -596
rect 359 -596 364 596
rect 380 -596 385 596
rect 359 -605 385 -596
rect -113 -610 385 -605
rect -113 -626 -78 -610
rect 350 -626 385 -610
rect -113 -631 385 -626
<< properties >>
string gencell rhigh
string library sg13g2_devstdin
string parameters w 0.5 l 10 nx 5 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class resistor endcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
