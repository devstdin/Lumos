magic
tech ihp-sg13g2
timestamp 1757240632
<< error_p >>
rect -33 80 -28 85
rect 28 80 33 85
rect 1150 80 1155 85
rect 1211 80 1216 85
rect 2333 80 2338 85
rect 2394 80 2399 85
rect 3516 80 3521 85
rect 3577 80 3582 85
rect -38 75 -33 80
rect 33 75 38 80
rect 1145 75 1150 80
rect 1216 75 1221 80
rect 2328 75 2333 80
rect 2399 75 2404 80
rect 3511 75 3516 80
rect 3582 75 3587 80
rect -38 64 -33 69
rect 33 64 38 69
rect 1145 64 1150 69
rect 1216 64 1221 69
rect 2328 64 2333 69
rect 2399 64 2404 69
rect 3511 64 3516 69
rect 3582 64 3587 69
rect -33 59 -28 64
rect 28 59 33 64
rect 1150 59 1155 64
rect 1211 59 1216 64
rect 2333 59 2338 64
rect 2394 59 2399 64
rect 3516 59 3521 64
rect 3577 59 3582 64
rect -67 43 -62 48
rect -56 43 -51 48
rect 51 43 56 48
rect 62 43 67 48
rect 1116 43 1121 48
rect 1127 43 1132 48
rect 1234 43 1239 48
rect 1245 43 1250 48
rect 2299 43 2304 48
rect 2310 43 2315 48
rect 2417 43 2422 48
rect 2428 43 2433 48
rect 3482 43 3487 48
rect 3493 43 3498 48
rect 3600 43 3605 48
rect 3611 43 3616 48
rect -72 38 -67 43
rect -51 38 -46 43
rect 46 38 51 43
rect 67 38 72 43
rect 1111 38 1116 43
rect 1132 38 1137 43
rect 1229 38 1234 43
rect 1250 38 1255 43
rect 2294 38 2299 43
rect 2315 38 2320 43
rect 2412 38 2417 43
rect 2433 38 2438 43
rect 3477 38 3482 43
rect 3498 38 3503 43
rect 3595 38 3600 43
rect 3616 38 3621 43
rect -72 -43 -67 -38
rect -51 -43 -46 -38
rect 46 -43 51 -38
rect 67 -43 72 -38
rect 1111 -43 1116 -38
rect 1132 -43 1137 -38
rect 1229 -43 1234 -38
rect 1250 -43 1255 -38
rect 2294 -43 2299 -38
rect 2315 -43 2320 -38
rect 2412 -43 2417 -38
rect 2433 -43 2438 -38
rect 3477 -43 3482 -38
rect 3498 -43 3503 -38
rect 3595 -43 3600 -38
rect 3616 -43 3621 -38
rect -67 -48 -62 -43
rect -56 -48 -51 -43
rect 51 -48 56 -43
rect 62 -48 67 -43
rect 1116 -48 1121 -43
rect 1127 -48 1132 -43
rect 1234 -48 1239 -43
rect 1245 -48 1250 -43
rect 2299 -48 2304 -43
rect 2310 -48 2315 -43
rect 2417 -48 2422 -43
rect 2428 -48 2433 -43
rect 3482 -48 3487 -43
rect 3493 -48 3498 -43
rect 3600 -48 3605 -43
rect 3611 -48 3616 -43
rect -33 -64 -28 -59
rect 28 -64 33 -59
rect 1150 -64 1155 -59
rect 1211 -64 1216 -59
rect 2333 -64 2338 -59
rect 2394 -64 2399 -59
rect 3516 -64 3521 -59
rect 3577 -64 3582 -59
rect -38 -69 -33 -64
rect 33 -69 38 -64
rect 1145 -69 1150 -64
rect 1216 -69 1221 -64
rect 2328 -69 2333 -64
rect 2399 -69 2404 -64
rect 3511 -69 3516 -64
rect 3582 -69 3587 -64
rect -38 -80 -33 -75
rect 33 -80 38 -75
rect 1145 -80 1150 -75
rect 1216 -80 1221 -75
rect 2328 -80 2333 -75
rect 2399 -80 2404 -75
rect 3511 -80 3516 -75
rect 3582 -80 3587 -75
rect -33 -85 -28 -80
rect 28 -85 33 -80
rect 1150 -85 1155 -80
rect 1211 -85 1216 -80
rect 2333 -85 2338 -80
rect 2394 -85 2399 -80
rect 3516 -85 3521 -80
rect 3577 -85 3582 -80
<< nwell >>
rect -136 87 136 112
rect 1047 87 1319 112
rect 2230 87 2502 112
rect 3413 87 3685 112
rect -247 -212 3796 87
<< hvpmos >>
rect -40 -50 40 50
rect 1143 -50 1223 50
rect 2326 -50 2406 50
rect 3509 -50 3589 50
<< hvpdiff >>
rect -74 43 -40 50
rect -74 -43 -67 43
rect -51 -43 -40 43
rect -74 -50 -40 -43
rect 40 43 74 50
rect 40 -43 51 43
rect 67 -43 74 43
rect 40 -50 74 -43
rect 1109 43 1143 50
rect 1109 -43 1116 43
rect 1132 -43 1143 43
rect 1109 -50 1143 -43
rect 1223 43 1257 50
rect 1223 -43 1234 43
rect 1250 -43 1257 43
rect 1223 -50 1257 -43
rect 2292 43 2326 50
rect 2292 -43 2299 43
rect 2315 -43 2326 43
rect 2292 -50 2326 -43
rect 2406 43 2440 50
rect 2406 -43 2417 43
rect 2433 -43 2440 43
rect 2406 -50 2440 -43
rect 3475 43 3509 50
rect 3475 -43 3482 43
rect 3498 -43 3509 43
rect 3475 -50 3509 -43
rect 3589 43 3623 50
rect 3589 -43 3600 43
rect 3616 -43 3623 43
rect 3589 -50 3623 -43
<< hvpdiffc >>
rect -67 -43 -51 43
rect 51 -43 67 43
rect 1116 -43 1132 43
rect 1234 -43 1250 43
rect 2299 -43 2315 43
rect 2417 -43 2433 43
rect 3482 -43 3498 43
rect 3600 -43 3616 43
<< nsubdiff >>
rect -185 18 -155 25
rect -185 -113 -178 18
rect -162 -113 -155 18
rect 3704 18 3734 25
rect -185 -120 -155 -113
rect 3704 -113 3711 18
rect 3727 -113 3734 18
rect 3704 -120 3734 -113
rect -185 -127 3734 -120
rect -185 -143 -148 -127
rect 3697 -143 3734 -127
rect -185 -150 3734 -143
<< nsubdiffcont >>
rect -178 -113 -162 18
rect 3711 -113 3727 18
rect -148 -143 3697 -127
<< poly >>
rect -40 80 40 87
rect -40 64 -33 80
rect 33 64 40 80
rect -40 50 40 64
rect 1143 80 1223 87
rect 1143 64 1150 80
rect 1216 64 1223 80
rect 1143 50 1223 64
rect 2326 80 2406 87
rect 2326 64 2333 80
rect 2399 64 2406 80
rect 2326 50 2406 64
rect 3509 80 3589 87
rect 3509 64 3516 80
rect 3582 64 3589 80
rect 3509 50 3589 64
rect -40 -64 40 -50
rect -40 -80 -33 -64
rect 33 -80 40 -64
rect -40 -87 40 -80
rect 1143 -64 1223 -50
rect 1143 -80 1150 -64
rect 1216 -80 1223 -64
rect 1143 -87 1223 -80
rect 2326 -64 2406 -50
rect 2326 -80 2333 -64
rect 2399 -80 2406 -64
rect 2326 -87 2406 -80
rect 3509 -64 3589 -50
rect 3509 -80 3516 -64
rect 3582 -80 3589 -64
rect 3509 -87 3589 -80
<< polycont >>
rect -33 64 33 80
rect 1150 64 1216 80
rect 2333 64 2399 80
rect 3516 64 3582 80
rect -33 -80 33 -64
rect 1150 -80 1216 -64
rect 2333 -80 2399 -64
rect 3516 -80 3582 -64
<< metal1 >>
rect -183 18 -157 23
rect -183 -113 -178 18
rect -162 -113 -157 18
rect 3706 18 3732 23
rect -183 -122 -157 -113
rect 3706 -113 3711 18
rect 3727 -113 3732 18
rect 3706 -122 3732 -113
rect -183 -127 3732 -122
rect -183 -143 -148 -127
rect 3697 -143 3732 -127
rect -183 -148 3732 -143
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 1 l 0.8 nf 1 nx 4 dx 10.35 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 0 gbc 1
<< end >>
