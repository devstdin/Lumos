magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 32 292 324 314
rect 32 56 745 292
rect -26 -56 794 56
<< nmos >>
rect 129 160 155 288
rect 204 160 230 288
rect 409 118 435 266
rect 523 118 549 266
rect 625 118 651 266
<< pmos >>
rect 166 429 192 597
rect 268 429 294 597
rect 409 412 435 636
rect 486 412 512 636
rect 598 412 624 636
<< ndiff >>
rect 58 274 129 288
rect 58 242 75 274
rect 107 242 129 274
rect 58 206 129 242
rect 58 174 75 206
rect 107 174 129 206
rect 58 160 129 174
rect 155 160 204 288
rect 230 206 298 288
rect 230 174 252 206
rect 284 174 298 206
rect 230 160 298 174
rect 341 195 409 266
rect 341 163 355 195
rect 387 163 409 195
rect 341 118 409 163
rect 435 128 523 266
rect 435 118 463 128
rect 449 96 463 118
rect 495 118 523 128
rect 549 195 625 266
rect 549 163 571 195
rect 603 163 625 195
rect 549 118 625 163
rect 651 232 719 266
rect 651 200 673 232
rect 705 200 719 232
rect 651 164 719 200
rect 651 132 673 164
rect 705 132 719 164
rect 651 118 719 132
rect 495 96 509 118
rect 449 82 509 96
<< pdiff >>
rect 341 622 409 636
rect 341 597 355 622
rect 58 583 166 597
rect 58 551 74 583
rect 106 551 166 583
rect 58 515 166 551
rect 58 483 74 515
rect 106 483 166 515
rect 58 429 166 483
rect 192 583 268 597
rect 192 551 214 583
rect 246 551 268 583
rect 192 515 268 551
rect 192 483 214 515
rect 246 483 268 515
rect 192 429 268 483
rect 294 590 355 597
rect 387 590 409 622
rect 294 554 409 590
rect 294 522 355 554
rect 387 522 409 554
rect 294 429 409 522
rect 341 412 409 429
rect 435 412 486 636
rect 512 622 598 636
rect 512 590 544 622
rect 576 590 598 622
rect 512 554 598 590
rect 512 522 544 554
rect 576 522 598 554
rect 512 486 598 522
rect 512 454 544 486
rect 576 454 598 486
rect 512 412 598 454
rect 624 622 692 636
rect 624 590 646 622
rect 678 590 692 622
rect 624 554 692 590
rect 624 522 646 554
rect 678 522 692 554
rect 624 412 692 522
<< ndiffc >>
rect 75 242 107 274
rect 75 174 107 206
rect 252 174 284 206
rect 355 163 387 195
rect 463 96 495 128
rect 571 163 603 195
rect 673 200 705 232
rect 673 132 705 164
<< pdiffc >>
rect 74 551 106 583
rect 74 483 106 515
rect 214 551 246 583
rect 214 483 246 515
rect 355 590 387 622
rect 355 522 387 554
rect 544 590 576 622
rect 544 522 576 554
rect 544 454 576 486
rect 646 590 678 622
rect 646 522 678 554
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 409 636 435 672
rect 486 636 512 672
rect 598 636 624 672
rect 166 597 192 633
rect 268 597 294 633
rect 166 414 192 429
rect 129 382 192 414
rect 129 288 155 382
rect 268 377 294 429
rect 409 377 435 412
rect 486 377 512 412
rect 248 363 314 377
rect 248 343 265 363
rect 204 331 265 343
rect 297 331 314 363
rect 204 317 314 331
rect 362 363 435 377
rect 362 331 379 363
rect 411 331 435 363
rect 362 317 435 331
rect 471 363 531 377
rect 598 370 624 412
rect 471 331 485 363
rect 517 352 531 363
rect 594 353 660 370
rect 517 331 549 352
rect 471 317 549 331
rect 204 288 230 317
rect 409 266 435 317
rect 523 266 549 317
rect 594 321 611 353
rect 643 321 660 353
rect 594 304 660 321
rect 625 266 651 304
rect 129 88 155 160
rect 204 124 230 160
rect 409 88 435 118
rect 129 62 435 88
rect 523 82 549 118
rect 625 82 651 118
<< polycont >>
rect 265 331 297 363
rect 379 331 411 363
rect 485 331 517 363
rect 611 321 643 353
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 64 583 116 712
rect 345 622 397 712
rect 64 551 74 583
rect 106 551 116 583
rect 64 515 116 551
rect 64 483 74 515
rect 106 483 116 515
rect 204 583 256 593
rect 204 551 214 583
rect 246 551 256 583
rect 204 515 256 551
rect 204 513 214 515
rect 64 473 116 483
rect 160 483 214 513
rect 246 483 256 515
rect 345 590 355 622
rect 387 590 397 622
rect 345 554 397 590
rect 345 522 355 554
rect 387 522 397 554
rect 345 512 397 522
rect 534 622 600 632
rect 534 590 544 622
rect 576 590 600 622
rect 534 554 600 590
rect 534 522 544 554
rect 576 522 600 554
rect 160 473 256 483
rect 534 486 600 522
rect 636 622 688 712
rect 636 590 646 622
rect 678 590 688 622
rect 636 554 688 590
rect 636 522 646 554
rect 678 522 688 554
rect 636 512 688 522
rect 64 274 117 284
rect 64 242 75 274
rect 107 242 117 274
rect 64 206 117 242
rect 64 174 75 206
rect 107 174 117 206
rect 64 44 117 174
rect 160 199 192 473
rect 534 454 544 486
rect 576 454 600 486
rect 534 448 600 454
rect 284 416 496 448
rect 534 416 714 448
rect 284 380 316 416
rect 248 363 316 380
rect 248 331 265 363
rect 297 331 316 363
rect 248 305 316 331
rect 352 363 415 380
rect 352 331 379 363
rect 411 331 415 363
rect 352 305 415 331
rect 464 373 496 416
rect 464 363 527 373
rect 464 331 485 363
rect 517 331 527 363
rect 464 321 527 331
rect 586 353 646 363
rect 586 321 611 353
rect 643 321 646 353
rect 586 311 646 321
rect 586 268 620 311
rect 242 236 620 268
rect 682 242 714 416
rect 242 206 294 236
rect 242 199 252 206
rect 160 174 252 199
rect 284 174 294 206
rect 663 232 714 242
rect 663 200 673 232
rect 705 200 714 232
rect 160 167 294 174
rect 345 195 613 200
rect 345 163 355 195
rect 387 166 571 195
rect 387 163 405 166
rect 345 160 405 163
rect 554 163 571 166
rect 603 163 613 195
rect 554 158 613 163
rect 663 164 714 200
rect 663 132 673 164
rect 705 132 714 164
rect 453 128 505 130
rect 453 96 463 128
rect 495 96 505 128
rect 663 122 714 132
rect 453 44 505 96
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 534 416 600 632 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 248 305 316 380 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 352 305 415 380 0 FreeSans 400 0 0 0 A
port 5 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 155316
string GDS_FILE 6_final.gds
string GDS_START 149086
<< end >>
