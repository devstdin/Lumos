magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 63 56 481 292
rect -26 -56 506 56
<< nmos >>
rect 157 118 183 266
rect 259 118 285 266
rect 361 138 387 266
<< pmos >>
rect 157 412 183 636
rect 259 412 285 636
rect 361 427 387 627
<< ndiff >>
rect 89 252 157 266
rect 89 220 103 252
rect 135 220 157 252
rect 89 164 157 220
rect 89 132 103 164
rect 135 132 157 164
rect 89 118 157 132
rect 183 252 259 266
rect 183 220 205 252
rect 237 220 259 252
rect 183 164 259 220
rect 183 132 205 164
rect 237 132 259 164
rect 183 118 259 132
rect 285 183 361 266
rect 285 151 307 183
rect 339 151 361 183
rect 285 138 361 151
rect 387 252 455 266
rect 387 220 409 252
rect 441 220 455 252
rect 387 184 455 220
rect 387 152 409 184
rect 441 152 455 184
rect 387 138 455 152
rect 285 118 347 138
<< pdiff >>
rect 26 622 157 636
rect 26 590 40 622
rect 72 590 157 622
rect 26 554 157 590
rect 26 522 40 554
rect 72 522 157 554
rect 26 412 157 522
rect 183 458 259 636
rect 183 426 205 458
rect 237 426 259 458
rect 183 412 259 426
rect 285 627 347 636
rect 285 613 361 627
rect 285 581 307 613
rect 339 581 361 613
rect 285 427 361 581
rect 387 609 455 627
rect 387 577 409 609
rect 441 577 455 609
rect 387 541 455 577
rect 387 509 409 541
rect 441 509 455 541
rect 387 473 455 509
rect 387 441 409 473
rect 441 441 455 473
rect 387 427 455 441
rect 285 412 347 427
<< ndiffc >>
rect 103 220 135 252
rect 103 132 135 164
rect 205 220 237 252
rect 205 132 237 164
rect 307 151 339 183
rect 409 220 441 252
rect 409 152 441 184
<< pdiffc >>
rect 40 590 72 622
rect 40 522 72 554
rect 205 426 237 458
rect 307 581 339 613
rect 409 577 441 609
rect 409 509 441 541
rect 409 441 441 473
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 157 636 183 672
rect 259 636 285 672
rect 361 627 387 663
rect 157 370 183 412
rect 259 370 285 412
rect 41 353 285 370
rect 41 321 55 353
rect 87 321 285 353
rect 41 304 285 321
rect 157 266 183 304
rect 259 266 285 304
rect 361 377 387 427
rect 361 363 428 377
rect 361 331 382 363
rect 414 331 428 363
rect 361 317 428 331
rect 361 266 387 317
rect 157 82 183 118
rect 259 82 285 118
rect 361 102 387 138
<< polycont >>
rect 55 321 87 353
rect 382 331 414 363
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 30 622 82 712
rect 30 590 40 622
rect 72 590 82 622
rect 30 554 82 590
rect 297 613 349 712
rect 297 581 307 613
rect 339 581 349 613
rect 297 579 349 581
rect 394 609 452 620
rect 30 522 40 554
rect 72 522 82 554
rect 394 577 409 609
rect 441 577 452 609
rect 394 542 452 577
rect 30 512 82 522
rect 121 541 452 542
rect 121 510 409 541
rect 121 475 153 510
rect 45 443 153 475
rect 195 458 247 468
rect 45 353 97 443
rect 195 426 205 458
rect 237 426 247 458
rect 195 370 247 426
rect 45 321 55 353
rect 87 321 97 353
rect 45 311 97 321
rect 134 304 247 370
rect 93 252 145 262
rect 93 220 103 252
rect 135 220 145 252
rect 93 164 145 220
rect 93 132 103 164
rect 135 132 145 164
rect 93 44 145 132
rect 195 252 247 304
rect 195 220 205 252
rect 237 220 247 252
rect 283 262 315 510
rect 394 509 409 510
rect 441 509 452 541
rect 394 473 452 509
rect 394 441 409 473
rect 441 441 452 473
rect 394 436 452 441
rect 351 363 428 374
rect 351 331 382 363
rect 414 331 428 363
rect 351 298 428 331
rect 283 252 451 262
rect 283 229 409 252
rect 195 164 247 220
rect 399 220 409 229
rect 441 220 451 252
rect 195 132 205 164
rect 237 132 247 164
rect 195 122 247 132
rect 297 183 349 193
rect 297 151 307 183
rect 339 151 349 183
rect 297 44 349 151
rect 399 184 451 220
rect 399 152 409 184
rect 441 152 451 184
rect 399 144 451 152
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 134 304 247 370 0 FreeSans 400 0 0 0 X
port 4 nsew
flabel metal1 s 351 298 428 374 0 FreeSans 400 0 0 0 A
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 79354
string GDS_FILE 6_final.gds
string GDS_START 75138
<< end >>
