magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753301161
<< nwell >>
rect 9537 380 10387 1568
<< metal1 >>
rect 482 12448 4647 12458
rect 482 12400 4470 12448
rect 4637 12400 4647 12448
rect 482 12390 4647 12400
rect 4896 12448 9066 12458
rect 4896 12400 4906 12448
rect 5078 12400 9066 12448
rect 4896 12390 9066 12400
rect 482 12364 554 12390
rect 760 12364 832 12390
rect 1038 12364 1110 12390
rect 1316 12364 1388 12390
rect 1594 12364 1666 12390
rect 1872 12364 1944 12390
rect 2150 12364 2222 12390
rect 2428 12364 2500 12390
rect 2706 12364 2778 12390
rect 2984 12364 3056 12390
rect 3262 12364 3334 12390
rect 3540 12364 3612 12390
rect 3818 12364 3890 12390
rect 4096 12364 4168 12390
rect 4374 12364 4446 12390
rect 5102 12364 5174 12390
rect 5380 12364 5452 12390
rect 5658 12364 5730 12390
rect 5936 12364 6008 12390
rect 6214 12364 6286 12390
rect 6492 12364 6564 12390
rect 6770 12364 6842 12390
rect 7048 12364 7120 12390
rect 7326 12364 7398 12390
rect 7604 12364 7676 12390
rect 7882 12364 7954 12390
rect 8160 12364 8232 12390
rect 8438 12364 8510 12390
rect 8716 12364 8788 12390
rect 8994 12364 9066 12390
rect 302 11076 456 12332
rect 302 10016 322 11076
rect 436 10016 456 11076
rect 302 8676 456 10016
rect 302 7616 322 8676
rect 436 7616 456 8676
rect 302 6276 456 7616
rect 302 5216 322 6276
rect 436 5216 456 6276
rect 302 3876 456 5216
rect 302 2816 322 3876
rect 436 2816 456 3876
rect 302 1476 456 2816
rect 302 416 322 1476
rect 436 416 456 1476
rect 302 360 456 416
rect 502 328 534 12364
rect 580 12276 734 12332
rect 580 11216 600 12276
rect 714 11216 734 12276
rect 580 9876 734 11216
rect 580 8816 600 9876
rect 714 8816 734 9876
rect 580 7476 734 8816
rect 580 6416 600 7476
rect 714 6416 734 7476
rect 580 5076 734 6416
rect 580 4016 600 5076
rect 714 4016 734 5076
rect 580 2676 734 4016
rect 580 1616 600 2676
rect 714 1616 734 2676
rect 580 360 734 1616
rect 780 328 812 12364
rect 858 11076 1012 12332
rect 858 10016 878 11076
rect 992 10016 1012 11076
rect 858 8676 1012 10016
rect 858 7616 878 8676
rect 992 7616 1012 8676
rect 858 6276 1012 7616
rect 858 5216 878 6276
rect 992 5216 1012 6276
rect 858 3876 1012 5216
rect 858 2816 878 3876
rect 992 2816 1012 3876
rect 858 1476 1012 2816
rect 858 416 878 1476
rect 992 416 1012 1476
rect 858 360 1012 416
rect 1058 328 1090 12364
rect 1136 12276 1290 12332
rect 1136 11216 1156 12276
rect 1270 11216 1290 12276
rect 1136 9876 1290 11216
rect 1136 8816 1156 9876
rect 1270 8816 1290 9876
rect 1136 7476 1290 8816
rect 1136 6416 1156 7476
rect 1270 6416 1290 7476
rect 1136 5076 1290 6416
rect 1136 4016 1156 5076
rect 1270 4016 1290 5076
rect 1136 2676 1290 4016
rect 1136 1616 1156 2676
rect 1270 1616 1290 2676
rect 1136 360 1290 1616
rect 1336 328 1368 12364
rect 1414 11076 1568 12332
rect 1414 10016 1434 11076
rect 1548 10016 1568 11076
rect 1414 8676 1568 10016
rect 1414 7616 1434 8676
rect 1548 7616 1568 8676
rect 1414 6276 1568 7616
rect 1414 5216 1434 6276
rect 1548 5216 1568 6276
rect 1414 3876 1568 5216
rect 1414 2816 1434 3876
rect 1548 2816 1568 3876
rect 1414 1476 1568 2816
rect 1414 416 1434 1476
rect 1548 416 1568 1476
rect 1414 360 1568 416
rect 1614 328 1646 12364
rect 1692 12276 1846 12332
rect 1692 11216 1712 12276
rect 1826 11216 1846 12276
rect 1692 9876 1846 11216
rect 1692 8816 1712 9876
rect 1826 8816 1846 9876
rect 1692 7476 1846 8816
rect 1692 6416 1712 7476
rect 1826 6416 1846 7476
rect 1692 5076 1846 6416
rect 1692 4016 1712 5076
rect 1826 4016 1846 5076
rect 1692 2676 1846 4016
rect 1692 1616 1712 2676
rect 1826 1616 1846 2676
rect 1692 360 1846 1616
rect 1892 328 1924 12364
rect 1970 11076 2124 12332
rect 1970 10016 1990 11076
rect 2104 10016 2124 11076
rect 1970 8676 2124 10016
rect 1970 7616 1990 8676
rect 2104 7616 2124 8676
rect 1970 6276 2124 7616
rect 1970 5216 1990 6276
rect 2104 5216 2124 6276
rect 1970 3876 2124 5216
rect 1970 2816 1990 3876
rect 2104 2816 2124 3876
rect 1970 1476 2124 2816
rect 1970 416 1990 1476
rect 2104 416 2124 1476
rect 1970 360 2124 416
rect 2170 328 2202 12364
rect 2248 12276 2402 12332
rect 2248 11216 2268 12276
rect 2382 11216 2402 12276
rect 2248 9876 2402 11216
rect 2248 8816 2268 9876
rect 2382 8816 2402 9876
rect 2248 7476 2402 8816
rect 2248 6416 2268 7476
rect 2382 6416 2402 7476
rect 2248 5076 2402 6416
rect 2248 4016 2268 5076
rect 2382 4016 2402 5076
rect 2248 2676 2402 4016
rect 2248 1616 2268 2676
rect 2382 1616 2402 2676
rect 2248 360 2402 1616
rect 2448 328 2480 12364
rect 2526 11076 2680 12332
rect 2526 10016 2546 11076
rect 2660 10016 2680 11076
rect 2526 8676 2680 10016
rect 2526 7616 2546 8676
rect 2660 7616 2680 8676
rect 2526 6276 2680 7616
rect 2526 5216 2546 6276
rect 2660 5216 2680 6276
rect 2526 3876 2680 5216
rect 2526 2816 2546 3876
rect 2660 2816 2680 3876
rect 2526 1476 2680 2816
rect 2526 416 2546 1476
rect 2660 416 2680 1476
rect 2526 360 2680 416
rect 2726 328 2758 12364
rect 2804 12276 2958 12332
rect 2804 11216 2824 12276
rect 2938 11216 2958 12276
rect 2804 9876 2958 11216
rect 2804 8816 2824 9876
rect 2938 8816 2958 9876
rect 2804 7476 2958 8816
rect 2804 6416 2824 7476
rect 2938 6416 2958 7476
rect 2804 5076 2958 6416
rect 2804 4016 2824 5076
rect 2938 4016 2958 5076
rect 2804 2676 2958 4016
rect 2804 1616 2824 2676
rect 2938 1616 2958 2676
rect 2804 360 2958 1616
rect 3004 328 3036 12364
rect 3082 11076 3236 12332
rect 3082 10016 3102 11076
rect 3216 10016 3236 11076
rect 3082 8676 3236 10016
rect 3082 7616 3102 8676
rect 3216 7616 3236 8676
rect 3082 6276 3236 7616
rect 3082 5216 3102 6276
rect 3216 5216 3236 6276
rect 3082 3876 3236 5216
rect 3082 2816 3102 3876
rect 3216 2816 3236 3876
rect 3082 1476 3236 2816
rect 3082 416 3102 1476
rect 3216 416 3236 1476
rect 3082 360 3236 416
rect 3282 328 3314 12364
rect 3360 12276 3514 12332
rect 3360 11216 3380 12276
rect 3494 11216 3514 12276
rect 3360 9876 3514 11216
rect 3360 8816 3380 9876
rect 3494 8816 3514 9876
rect 3360 7476 3514 8816
rect 3360 6416 3380 7476
rect 3494 6416 3514 7476
rect 3360 5076 3514 6416
rect 3360 4016 3380 5076
rect 3494 4016 3514 5076
rect 3360 2676 3514 4016
rect 3360 1616 3380 2676
rect 3494 1616 3514 2676
rect 3360 360 3514 1616
rect 3560 328 3592 12364
rect 3638 11076 3792 12332
rect 3638 10016 3658 11076
rect 3772 10016 3792 11076
rect 3638 8676 3792 10016
rect 3638 7616 3658 8676
rect 3772 7616 3792 8676
rect 3638 6276 3792 7616
rect 3638 5216 3658 6276
rect 3772 5216 3792 6276
rect 3638 3876 3792 5216
rect 3638 2816 3658 3876
rect 3772 2816 3792 3876
rect 3638 1476 3792 2816
rect 3638 416 3658 1476
rect 3772 416 3792 1476
rect 3638 360 3792 416
rect 3838 328 3870 12364
rect 3916 12276 4070 12332
rect 3916 11216 3936 12276
rect 4050 11216 4070 12276
rect 3916 9876 4070 11216
rect 3916 8816 3936 9876
rect 4050 8816 4070 9876
rect 3916 7476 4070 8816
rect 3916 6416 3936 7476
rect 4050 6416 4070 7476
rect 3916 5076 4070 6416
rect 3916 4016 3936 5076
rect 4050 4016 4070 5076
rect 3916 2676 4070 4016
rect 3916 1616 3936 2676
rect 4050 1616 4070 2676
rect 3916 360 4070 1616
rect 4116 328 4148 12364
rect 4194 11076 4348 12332
rect 4194 10016 4214 11076
rect 4328 10016 4348 11076
rect 4194 8676 4348 10016
rect 4194 7616 4214 8676
rect 4328 7616 4348 8676
rect 4194 6276 4348 7616
rect 4194 5216 4214 6276
rect 4328 5216 4348 6276
rect 4194 3876 4348 5216
rect 4194 2816 4214 3876
rect 4328 2816 4348 3876
rect 4194 1476 4348 2816
rect 4194 416 4214 1476
rect 4328 416 4348 1476
rect 4194 360 4348 416
rect 4394 328 4426 12364
rect 4472 12276 4626 12332
rect 4472 11216 4492 12276
rect 4606 11216 4626 12276
rect 4472 9876 4626 11216
rect 4472 8816 4492 9876
rect 4606 8816 4626 9876
rect 4472 7476 4626 8816
rect 4472 6416 4492 7476
rect 4606 6416 4626 7476
rect 4472 5076 4626 6416
rect 4472 4016 4492 5076
rect 4606 4016 4626 5076
rect 4472 2676 4626 4016
rect 4472 1616 4492 2676
rect 4606 1616 4626 2676
rect 4472 360 4626 1616
rect 4922 12276 5076 12332
rect 4922 11216 4942 12276
rect 5056 11216 5076 12276
rect 4922 9876 5076 11216
rect 4922 8816 4942 9876
rect 5056 8816 5076 9876
rect 4922 7476 5076 8816
rect 4922 6416 4942 7476
rect 5056 6416 5076 7476
rect 4922 5076 5076 6416
rect 4922 4016 4942 5076
rect 5056 4016 5076 5076
rect 4922 2676 5076 4016
rect 4922 1616 4942 2676
rect 5056 1616 5076 2676
rect 4922 360 5076 1616
rect 5122 328 5154 12364
rect 5200 11076 5354 12332
rect 5200 10016 5220 11076
rect 5334 10016 5354 11076
rect 5200 8676 5354 10016
rect 5200 7616 5220 8676
rect 5334 7616 5354 8676
rect 5200 6276 5354 7616
rect 5200 5216 5220 6276
rect 5334 5216 5354 6276
rect 5200 3876 5354 5216
rect 5200 2816 5220 3876
rect 5334 2816 5354 3876
rect 5200 1476 5354 2816
rect 5200 416 5220 1476
rect 5334 416 5354 1476
rect 5200 360 5354 416
rect 5400 328 5432 12364
rect 5478 12276 5632 12332
rect 5478 11216 5498 12276
rect 5612 11216 5632 12276
rect 5478 9876 5632 11216
rect 5478 8816 5498 9876
rect 5612 8816 5632 9876
rect 5478 7476 5632 8816
rect 5478 6416 5498 7476
rect 5612 6416 5632 7476
rect 5478 5076 5632 6416
rect 5478 4016 5498 5076
rect 5612 4016 5632 5076
rect 5478 2676 5632 4016
rect 5478 1616 5498 2676
rect 5612 1616 5632 2676
rect 5478 360 5632 1616
rect 5678 328 5710 12364
rect 5756 11076 5910 12332
rect 5756 10016 5776 11076
rect 5890 10016 5910 11076
rect 5756 8676 5910 10016
rect 5756 7616 5776 8676
rect 5890 7616 5910 8676
rect 5756 6276 5910 7616
rect 5756 5216 5776 6276
rect 5890 5216 5910 6276
rect 5756 3876 5910 5216
rect 5756 2816 5776 3876
rect 5890 2816 5910 3876
rect 5756 1476 5910 2816
rect 5756 416 5776 1476
rect 5890 416 5910 1476
rect 5756 360 5910 416
rect 5956 328 5988 12364
rect 6034 12276 6188 12332
rect 6034 11216 6054 12276
rect 6168 11216 6188 12276
rect 6034 9876 6188 11216
rect 6034 8816 6054 9876
rect 6168 8816 6188 9876
rect 6034 7476 6188 8816
rect 6034 6416 6054 7476
rect 6168 6416 6188 7476
rect 6034 5076 6188 6416
rect 6034 4016 6054 5076
rect 6168 4016 6188 5076
rect 6034 2676 6188 4016
rect 6034 1616 6054 2676
rect 6168 1616 6188 2676
rect 6034 360 6188 1616
rect 6234 328 6266 12364
rect 6312 11076 6466 12332
rect 6312 10016 6332 11076
rect 6446 10016 6466 11076
rect 6312 8676 6466 10016
rect 6312 7616 6332 8676
rect 6446 7616 6466 8676
rect 6312 6276 6466 7616
rect 6312 5216 6332 6276
rect 6446 5216 6466 6276
rect 6312 3876 6466 5216
rect 6312 2816 6332 3876
rect 6446 2816 6466 3876
rect 6312 1476 6466 2816
rect 6312 416 6332 1476
rect 6446 416 6466 1476
rect 6312 360 6466 416
rect 6512 328 6544 12364
rect 6590 12276 6744 12332
rect 6590 11216 6610 12276
rect 6724 11216 6744 12276
rect 6590 9876 6744 11216
rect 6590 8816 6610 9876
rect 6724 8816 6744 9876
rect 6590 7476 6744 8816
rect 6590 6416 6610 7476
rect 6724 6416 6744 7476
rect 6590 5076 6744 6416
rect 6590 4016 6610 5076
rect 6724 4016 6744 5076
rect 6590 2676 6744 4016
rect 6590 1616 6610 2676
rect 6724 1616 6744 2676
rect 6590 360 6744 1616
rect 6790 328 6822 12364
rect 6868 11076 7022 12332
rect 6868 10016 6888 11076
rect 7002 10016 7022 11076
rect 6868 8676 7022 10016
rect 6868 7616 6888 8676
rect 7002 7616 7022 8676
rect 6868 6276 7022 7616
rect 6868 5216 6888 6276
rect 7002 5216 7022 6276
rect 6868 3876 7022 5216
rect 6868 2816 6888 3876
rect 7002 2816 7022 3876
rect 6868 1476 7022 2816
rect 6868 416 6888 1476
rect 7002 416 7022 1476
rect 6868 360 7022 416
rect 7068 328 7100 12364
rect 7146 12276 7300 12332
rect 7146 11216 7166 12276
rect 7280 11216 7300 12276
rect 7146 9876 7300 11216
rect 7146 8816 7166 9876
rect 7280 8816 7300 9876
rect 7146 7476 7300 8816
rect 7146 6416 7166 7476
rect 7280 6416 7300 7476
rect 7146 5076 7300 6416
rect 7146 4016 7166 5076
rect 7280 4016 7300 5076
rect 7146 2676 7300 4016
rect 7146 1616 7166 2676
rect 7280 1616 7300 2676
rect 7146 360 7300 1616
rect 7346 328 7378 12364
rect 7424 11076 7578 12332
rect 7424 10016 7444 11076
rect 7558 10016 7578 11076
rect 7424 8676 7578 10016
rect 7424 7616 7444 8676
rect 7558 7616 7578 8676
rect 7424 6276 7578 7616
rect 7424 5216 7444 6276
rect 7558 5216 7578 6276
rect 7424 3876 7578 5216
rect 7424 2816 7444 3876
rect 7558 2816 7578 3876
rect 7424 1476 7578 2816
rect 7424 416 7444 1476
rect 7558 416 7578 1476
rect 7424 360 7578 416
rect 7624 328 7656 12364
rect 7702 12276 7856 12332
rect 7702 11216 7722 12276
rect 7836 11216 7856 12276
rect 7702 9876 7856 11216
rect 7702 8816 7722 9876
rect 7836 8816 7856 9876
rect 7702 7476 7856 8816
rect 7702 6416 7722 7476
rect 7836 6416 7856 7476
rect 7702 5076 7856 6416
rect 7702 4016 7722 5076
rect 7836 4016 7856 5076
rect 7702 2676 7856 4016
rect 7702 1616 7722 2676
rect 7836 1616 7856 2676
rect 7702 360 7856 1616
rect 7902 328 7934 12364
rect 7980 11076 8134 12332
rect 7980 10016 8000 11076
rect 8114 10016 8134 11076
rect 7980 8676 8134 10016
rect 7980 7616 8000 8676
rect 8114 7616 8134 8676
rect 7980 6276 8134 7616
rect 7980 5216 8000 6276
rect 8114 5216 8134 6276
rect 7980 3876 8134 5216
rect 7980 2816 8000 3876
rect 8114 2816 8134 3876
rect 7980 1476 8134 2816
rect 7980 416 8000 1476
rect 8114 416 8134 1476
rect 7980 360 8134 416
rect 8180 328 8212 12364
rect 8258 12276 8412 12332
rect 8258 11216 8278 12276
rect 8392 11216 8412 12276
rect 8258 9876 8412 11216
rect 8258 8816 8278 9876
rect 8392 8816 8412 9876
rect 8258 7476 8412 8816
rect 8258 6416 8278 7476
rect 8392 6416 8412 7476
rect 8258 5076 8412 6416
rect 8258 4016 8278 5076
rect 8392 4016 8412 5076
rect 8258 2676 8412 4016
rect 8258 1616 8278 2676
rect 8392 1616 8412 2676
rect 8258 360 8412 1616
rect 8458 328 8490 12364
rect 8536 11076 8690 12332
rect 8536 10016 8556 11076
rect 8670 10016 8690 11076
rect 8536 8676 8690 10016
rect 8536 7616 8556 8676
rect 8670 7616 8690 8676
rect 8536 6276 8690 7616
rect 8536 5216 8556 6276
rect 8670 5216 8690 6276
rect 8536 3876 8690 5216
rect 8536 2816 8556 3876
rect 8670 2816 8690 3876
rect 8536 1476 8690 2816
rect 8536 416 8556 1476
rect 8670 416 8690 1476
rect 8536 360 8690 416
rect 8736 328 8768 12364
rect 8814 12276 8968 12332
rect 8814 11216 8834 12276
rect 8948 11216 8968 12276
rect 8814 9876 8968 11216
rect 8814 8816 8834 9876
rect 8948 8816 8968 9876
rect 8814 7476 8968 8816
rect 8814 6416 8834 7476
rect 8948 6416 8968 7476
rect 8814 5076 8968 6416
rect 8814 4016 8834 5076
rect 8948 4016 8968 5076
rect 8814 2676 8968 4016
rect 8814 1616 8834 2676
rect 8948 1616 8968 2676
rect 8814 360 8968 1616
rect 9014 328 9046 12364
rect 9092 11076 9246 12332
rect 9092 10016 9112 11076
rect 9226 10016 9246 11076
rect 9092 8676 9246 10016
rect 9092 7616 9112 8676
rect 9226 7616 9246 8676
rect 9092 6276 9246 7616
rect 9092 5216 9112 6276
rect 9226 5216 9246 6276
rect 9092 3876 9246 5216
rect 9092 2816 9112 3876
rect 9226 2816 9246 3876
rect 9092 1476 9246 2816
rect 9092 416 9112 1476
rect 9226 416 9246 1476
rect 9092 360 9246 416
rect 9372 12276 9509 12564
rect 9372 11216 9388 12276
rect 9489 11216 9509 12276
rect 9372 9876 9509 11216
rect 9372 8816 9388 9876
rect 9489 8816 9509 9876
rect 9372 7476 9509 8816
rect 9372 6416 9388 7476
rect 9489 6416 9509 7476
rect 9372 5076 9509 6416
rect 9372 4016 9388 5076
rect 9489 4016 9509 5076
rect 9372 2676 9509 4016
rect 9372 1616 9388 2676
rect 9489 1616 9509 2676
rect 9372 1471 9509 1616
rect 9372 1428 10257 1471
rect 9372 1314 9817 1428
rect 9975 1386 10047 1428
rect 482 302 554 328
rect 760 302 832 328
rect 1038 302 1110 328
rect 1316 302 1388 328
rect 1594 302 1666 328
rect 1872 302 1944 328
rect 2150 302 2222 328
rect 2428 302 2500 328
rect 2706 302 2778 328
rect 2984 302 3056 328
rect 3262 302 3334 328
rect 3540 302 3612 328
rect 3818 302 3890 328
rect 4096 302 4168 328
rect 4374 302 4446 328
rect 5102 302 5174 328
rect 5380 302 5452 328
rect 5658 302 5730 328
rect 5936 302 6008 328
rect 6214 302 6286 328
rect 6492 302 6564 328
rect 6770 302 6842 328
rect 7048 302 7120 328
rect 7326 302 7398 328
rect 7604 302 7676 328
rect 7882 302 7954 328
rect 8160 302 8232 328
rect 8438 302 8510 328
rect 8716 302 8788 328
rect 8994 302 9066 328
rect 482 292 4647 302
rect 482 244 4470 292
rect 4637 244 4647 292
rect 482 234 4647 244
rect 4896 292 9309 302
rect 4896 244 4906 292
rect 5078 244 9129 292
rect 9299 244 9309 292
rect 4896 234 9309 244
rect 9372 129 9509 1314
rect 9765 634 9817 1314
rect 9891 1012 9943 1360
rect 10079 1012 10154 1360
rect 9891 949 10154 1012
rect 9891 588 9943 949
rect 10079 588 10154 949
rect 10205 634 10257 1428
rect 9975 469 10047 562
rect 9600 339 10047 469
rect 9600 292 9672 339
rect 9600 134 9610 292
rect 9662 134 9672 292
rect 9600 124 9672 134
rect -3 -709 324 -57
rect 460 -529 512 -237
rect 8572 -247 8705 -237
rect 8572 -319 8582 -247
rect 8695 -319 8705 -247
rect 8572 -329 8705 -319
rect 9743 -288 9795 240
rect 9975 188 10047 339
rect 10106 536 10154 588
rect 10106 335 10518 536
rect 10106 162 10154 335
rect 9891 20 9943 162
rect 10079 20 10154 162
rect 9845 10 10154 20
rect 9845 -62 9855 10
rect 9933 -62 10154 10
rect 9845 -72 10154 -62
rect 9891 -210 9943 -72
rect 10079 -210 10154 -72
rect 9975 -288 10047 -236
rect 10227 -288 10279 240
rect 9743 -437 10279 -288
rect 8572 -529 10279 -437
rect 8752 -709 10279 -529
<< via1 >>
rect 4470 12400 4637 12448
rect 4906 12400 5078 12448
rect 322 10016 436 11076
rect 322 7616 436 8676
rect 322 5216 436 6276
rect 322 2816 436 3876
rect 322 416 436 1476
rect 600 11216 714 12276
rect 600 8816 714 9876
rect 600 6416 714 7476
rect 600 4016 714 5076
rect 600 1616 714 2676
rect 878 10016 992 11076
rect 878 7616 992 8676
rect 878 5216 992 6276
rect 878 2816 992 3876
rect 878 416 992 1476
rect 1156 11216 1270 12276
rect 1156 8816 1270 9876
rect 1156 6416 1270 7476
rect 1156 4016 1270 5076
rect 1156 1616 1270 2676
rect 1434 10016 1548 11076
rect 1434 7616 1548 8676
rect 1434 5216 1548 6276
rect 1434 2816 1548 3876
rect 1434 416 1548 1476
rect 1712 11216 1826 12276
rect 1712 8816 1826 9876
rect 1712 6416 1826 7476
rect 1712 4016 1826 5076
rect 1712 1616 1826 2676
rect 1990 10016 2104 11076
rect 1990 7616 2104 8676
rect 1990 5216 2104 6276
rect 1990 2816 2104 3876
rect 1990 416 2104 1476
rect 2268 11216 2382 12276
rect 2268 8816 2382 9876
rect 2268 6416 2382 7476
rect 2268 4016 2382 5076
rect 2268 1616 2382 2676
rect 2546 10016 2660 11076
rect 2546 7616 2660 8676
rect 2546 5216 2660 6276
rect 2546 2816 2660 3876
rect 2546 416 2660 1476
rect 2824 11216 2938 12276
rect 2824 8816 2938 9876
rect 2824 6416 2938 7476
rect 2824 4016 2938 5076
rect 2824 1616 2938 2676
rect 3102 10016 3216 11076
rect 3102 7616 3216 8676
rect 3102 5216 3216 6276
rect 3102 2816 3216 3876
rect 3102 416 3216 1476
rect 3380 11216 3494 12276
rect 3380 8816 3494 9876
rect 3380 6416 3494 7476
rect 3380 4016 3494 5076
rect 3380 1616 3494 2676
rect 3658 10016 3772 11076
rect 3658 7616 3772 8676
rect 3658 5216 3772 6276
rect 3658 2816 3772 3876
rect 3658 416 3772 1476
rect 3936 11216 4050 12276
rect 3936 8816 4050 9876
rect 3936 6416 4050 7476
rect 3936 4016 4050 5076
rect 3936 1616 4050 2676
rect 4214 10016 4328 11076
rect 4214 7616 4328 8676
rect 4214 5216 4328 6276
rect 4214 2816 4328 3876
rect 4214 416 4328 1476
rect 4492 11216 4606 12276
rect 4492 8816 4606 9876
rect 4492 6416 4606 7476
rect 4492 4016 4606 5076
rect 4492 1616 4606 2676
rect 4942 11216 5056 12276
rect 4942 8816 5056 9876
rect 4942 6416 5056 7476
rect 4942 4016 5056 5076
rect 4942 1616 5056 2676
rect 5220 10016 5334 11076
rect 5220 7616 5334 8676
rect 5220 5216 5334 6276
rect 5220 2816 5334 3876
rect 5220 416 5334 1476
rect 5498 11216 5612 12276
rect 5498 8816 5612 9876
rect 5498 6416 5612 7476
rect 5498 4016 5612 5076
rect 5498 1616 5612 2676
rect 5776 10016 5890 11076
rect 5776 7616 5890 8676
rect 5776 5216 5890 6276
rect 5776 2816 5890 3876
rect 5776 416 5890 1476
rect 6054 11216 6168 12276
rect 6054 8816 6168 9876
rect 6054 6416 6168 7476
rect 6054 4016 6168 5076
rect 6054 1616 6168 2676
rect 6332 10016 6446 11076
rect 6332 7616 6446 8676
rect 6332 5216 6446 6276
rect 6332 2816 6446 3876
rect 6332 416 6446 1476
rect 6610 11216 6724 12276
rect 6610 8816 6724 9876
rect 6610 6416 6724 7476
rect 6610 4016 6724 5076
rect 6610 1616 6724 2676
rect 6888 10016 7002 11076
rect 6888 7616 7002 8676
rect 6888 5216 7002 6276
rect 6888 2816 7002 3876
rect 6888 416 7002 1476
rect 7166 11216 7280 12276
rect 7166 8816 7280 9876
rect 7166 6416 7280 7476
rect 7166 4016 7280 5076
rect 7166 1616 7280 2676
rect 7444 10016 7558 11076
rect 7444 7616 7558 8676
rect 7444 5216 7558 6276
rect 7444 2816 7558 3876
rect 7444 416 7558 1476
rect 7722 11216 7836 12276
rect 7722 8816 7836 9876
rect 7722 6416 7836 7476
rect 7722 4016 7836 5076
rect 7722 1616 7836 2676
rect 8000 10016 8114 11076
rect 8000 7616 8114 8676
rect 8000 5216 8114 6276
rect 8000 2816 8114 3876
rect 8000 416 8114 1476
rect 8278 11216 8392 12276
rect 8278 8816 8392 9876
rect 8278 6416 8392 7476
rect 8278 4016 8392 5076
rect 8278 1616 8392 2676
rect 8556 10016 8670 11076
rect 8556 7616 8670 8676
rect 8556 5216 8670 6276
rect 8556 2816 8670 3876
rect 8556 416 8670 1476
rect 8834 11216 8948 12276
rect 8834 8816 8948 9876
rect 8834 6416 8948 7476
rect 8834 4016 8948 5076
rect 8834 1616 8948 2676
rect 9112 10016 9226 11076
rect 9112 7616 9226 8676
rect 9112 5216 9226 6276
rect 9112 2816 9226 3876
rect 9112 416 9226 1476
rect 9388 11216 9489 12276
rect 9388 8816 9489 9876
rect 9388 6416 9489 7476
rect 9388 4016 9489 5076
rect 9388 1616 9489 2676
rect 4470 244 4637 292
rect 4906 244 5078 292
rect 9129 244 9299 292
rect 9610 134 9662 292
rect 8582 -319 8695 -247
rect 9855 -62 9933 10
<< metal2 >>
rect 4460 12448 5088 12458
rect 4460 12400 4470 12448
rect 4637 12400 4906 12448
rect 5078 12400 5088 12448
rect 4460 12390 5088 12400
rect 302 12276 10525 12296
rect 302 11216 600 12276
rect 714 11216 1156 12276
rect 1270 11216 1712 12276
rect 1826 11216 2268 12276
rect 2382 11216 2824 12276
rect 2938 11216 3380 12276
rect 3494 11216 3936 12276
rect 4050 11216 4492 12276
rect 4606 11216 4942 12276
rect 5056 11216 5498 12276
rect 5612 11216 6054 12276
rect 6168 11216 6610 12276
rect 6724 11216 7166 12276
rect 7280 11216 7722 12276
rect 7836 11216 8278 12276
rect 8392 11216 8834 12276
rect 8948 11216 9388 12276
rect 9489 12203 10525 12276
rect 9489 11216 9585 12203
rect 302 11196 9585 11216
rect -977 11076 9246 11096
rect -977 10997 322 11076
rect -977 496 -877 10997
rect -37 10016 322 10997
rect 436 10016 878 11076
rect 992 10016 1434 11076
rect 1548 10016 1990 11076
rect 2104 10016 2546 11076
rect 2660 10016 3102 11076
rect 3216 10016 3658 11076
rect 3772 10016 4214 11076
rect 4328 10016 5220 11076
rect 5334 10016 5776 11076
rect 5890 10016 6332 11076
rect 6446 10016 6888 11076
rect 7002 10016 7444 11076
rect 7558 10016 8000 11076
rect 8114 10016 8556 11076
rect 8670 10016 9112 11076
rect 9226 10016 9246 11076
rect -37 9996 9246 10016
rect -37 8696 63 9996
rect 9485 9896 9585 11196
rect 302 9876 9585 9896
rect 302 8816 600 9876
rect 714 8816 1156 9876
rect 1270 8816 1712 9876
rect 1826 8816 2268 9876
rect 2382 8816 2824 9876
rect 2938 8816 3380 9876
rect 3494 8816 3936 9876
rect 4050 8816 4492 9876
rect 4606 8816 4942 9876
rect 5056 8816 5498 9876
rect 5612 8816 6054 9876
rect 6168 8816 6610 9876
rect 6724 8816 7166 9876
rect 7280 8816 7722 9876
rect 7836 8816 8278 9876
rect 8392 8816 8834 9876
rect 8948 8816 9388 9876
rect 9489 8816 9585 9876
rect 302 8796 9585 8816
rect -37 8676 9246 8696
rect -37 7616 322 8676
rect 436 7616 878 8676
rect 992 7616 1434 8676
rect 1548 7616 1990 8676
rect 2104 7616 2546 8676
rect 2660 7616 3102 8676
rect 3216 7616 3658 8676
rect 3772 7616 4214 8676
rect 4328 7616 5220 8676
rect 5334 7616 5776 8676
rect 5890 7616 6332 8676
rect 6446 7616 6888 8676
rect 7002 7616 7444 8676
rect 7558 7616 8000 8676
rect 8114 7616 8556 8676
rect 8670 7616 9112 8676
rect 9226 7616 9246 8676
rect -37 7596 9246 7616
rect -37 6296 63 7596
rect 9485 7496 9585 8796
rect 302 7476 9585 7496
rect 302 6416 600 7476
rect 714 6416 1156 7476
rect 1270 6416 1712 7476
rect 1826 6416 2268 7476
rect 2382 6416 2824 7476
rect 2938 6416 3380 7476
rect 3494 6416 3936 7476
rect 4050 6416 4492 7476
rect 4606 6416 4942 7476
rect 5056 6416 5498 7476
rect 5612 6416 6054 7476
rect 6168 6416 6610 7476
rect 6724 6416 7166 7476
rect 7280 6416 7722 7476
rect 7836 6416 8278 7476
rect 8392 6416 8834 7476
rect 8948 6416 9388 7476
rect 9489 6416 9585 7476
rect 302 6396 9585 6416
rect -37 6276 9246 6296
rect -37 5216 322 6276
rect 436 5216 878 6276
rect 992 5216 1434 6276
rect 1548 5216 1990 6276
rect 2104 5216 2546 6276
rect 2660 5216 3102 6276
rect 3216 5216 3658 6276
rect 3772 5216 4214 6276
rect 4328 5216 5220 6276
rect 5334 5216 5776 6276
rect 5890 5216 6332 6276
rect 6446 5216 6888 6276
rect 7002 5216 7444 6276
rect 7558 5216 8000 6276
rect 8114 5216 8556 6276
rect 8670 5216 9112 6276
rect 9226 5216 9246 6276
rect -37 5196 9246 5216
rect -37 3896 63 5196
rect 9485 5096 9585 6396
rect 302 5076 9585 5096
rect 302 4016 600 5076
rect 714 4016 1156 5076
rect 1270 4016 1712 5076
rect 1826 4016 2268 5076
rect 2382 4016 2824 5076
rect 2938 4016 3380 5076
rect 3494 4016 3936 5076
rect 4050 4016 4492 5076
rect 4606 4016 4942 5076
rect 5056 4016 5498 5076
rect 5612 4016 6054 5076
rect 6168 4016 6610 5076
rect 6724 4016 7166 5076
rect 7280 4016 7722 5076
rect 7836 4016 8278 5076
rect 8392 4016 8834 5076
rect 8948 4016 9388 5076
rect 9489 4016 9585 5076
rect 302 3996 9585 4016
rect -37 3876 9246 3896
rect -37 2816 322 3876
rect 436 2816 878 3876
rect 992 2816 1434 3876
rect 1548 2816 1990 3876
rect 2104 2816 2546 3876
rect 2660 2816 3102 3876
rect 3216 2816 3658 3876
rect 3772 2816 4214 3876
rect 4328 2816 5220 3876
rect 5334 2816 5776 3876
rect 5890 2816 6332 3876
rect 6446 2816 6888 3876
rect 7002 2816 7444 3876
rect 7558 2816 8000 3876
rect 8114 2816 8556 3876
rect 8670 2816 9112 3876
rect 9226 2816 9246 3876
rect -37 2796 9246 2816
rect -37 1496 63 2796
rect 9485 2696 9585 3996
rect 302 2676 9585 2696
rect 302 1616 600 2676
rect 714 1616 1156 2676
rect 1270 1616 1712 2676
rect 1826 1616 2268 2676
rect 2382 1616 2824 2676
rect 2938 1616 3380 2676
rect 3494 1616 3936 2676
rect 4050 1616 4492 2676
rect 4606 1616 4942 2676
rect 5056 1616 5498 2676
rect 5612 1616 6054 2676
rect 6168 1616 6610 2676
rect 6724 1616 7166 2676
rect 7280 1616 7722 2676
rect 7836 1616 8278 2676
rect 8392 1616 8834 2676
rect 8948 1616 9388 2676
rect 9489 1696 9585 2676
rect 10425 1696 10525 12203
rect 9489 1616 10525 1696
rect 302 1596 10525 1616
rect -37 1476 9246 1496
rect -37 496 322 1476
rect -977 416 322 496
rect 436 416 878 1476
rect 992 416 1434 1476
rect 1548 416 1990 1476
rect 2104 416 2546 1476
rect 2660 416 3102 1476
rect 3216 416 3658 1476
rect 3772 416 4214 1476
rect 4328 416 5220 1476
rect 5334 416 5776 1476
rect 5890 416 6332 1476
rect 6446 416 6888 1476
rect 7002 416 7444 1476
rect 7558 416 8000 1476
rect 8114 416 8556 1476
rect 8670 416 9112 1476
rect 9226 416 9246 1476
rect -977 396 9246 416
rect 4460 292 5088 302
rect 4460 244 4470 292
rect 4637 244 4906 292
rect 5078 244 5088 292
rect 4460 234 5088 244
rect 9119 292 9672 302
rect 9119 244 9129 292
rect 9299 244 9610 292
rect 9119 134 9610 244
rect 9662 134 9672 292
rect 9119 124 9672 134
rect 9569 10 9943 20
rect 9569 -62 9855 10
rect 9933 -62 9943 10
rect 9569 -72 9943 -62
rect 9569 -237 9661 -72
rect 8572 -247 9661 -237
rect 8572 -319 8582 -247
rect 8695 -319 9661 -247
rect 8572 -329 9661 -319
<< via2 >>
rect 600 11216 714 12276
rect 1156 11216 1270 12276
rect 1712 11216 1826 12276
rect 2268 11216 2382 12276
rect 2824 11216 2938 12276
rect 3380 11216 3494 12276
rect 3936 11216 4050 12276
rect 4492 11216 4606 12276
rect 4942 11216 5056 12276
rect 5498 11216 5612 12276
rect 6054 11216 6168 12276
rect 6610 11216 6724 12276
rect 7166 11216 7280 12276
rect 7722 11216 7836 12276
rect 8278 11216 8392 12276
rect 8834 11216 8948 12276
rect -877 496 -37 10997
rect 322 10016 436 11076
rect 878 10016 992 11076
rect 1434 10016 1548 11076
rect 1990 10016 2104 11076
rect 2546 10016 2660 11076
rect 3102 10016 3216 11076
rect 3658 10016 3772 11076
rect 4214 10016 4328 11076
rect 5220 10016 5334 11076
rect 5776 10016 5890 11076
rect 6332 10016 6446 11076
rect 6888 10016 7002 11076
rect 7444 10016 7558 11076
rect 8000 10016 8114 11076
rect 8556 10016 8670 11076
rect 9112 10016 9226 11076
rect 600 8816 714 9876
rect 1156 8816 1270 9876
rect 1712 8816 1826 9876
rect 2268 8816 2382 9876
rect 2824 8816 2938 9876
rect 3380 8816 3494 9876
rect 3936 8816 4050 9876
rect 4492 8816 4606 9876
rect 4942 8816 5056 9876
rect 5498 8816 5612 9876
rect 6054 8816 6168 9876
rect 6610 8816 6724 9876
rect 7166 8816 7280 9876
rect 7722 8816 7836 9876
rect 8278 8816 8392 9876
rect 8834 8816 8948 9876
rect 322 7616 436 8676
rect 878 7616 992 8676
rect 1434 7616 1548 8676
rect 1990 7616 2104 8676
rect 2546 7616 2660 8676
rect 3102 7616 3216 8676
rect 3658 7616 3772 8676
rect 4214 7616 4328 8676
rect 5220 7616 5334 8676
rect 5776 7616 5890 8676
rect 6332 7616 6446 8676
rect 6888 7616 7002 8676
rect 7444 7616 7558 8676
rect 8000 7616 8114 8676
rect 8556 7616 8670 8676
rect 9112 7616 9226 8676
rect 600 6416 714 7476
rect 1156 6416 1270 7476
rect 1712 6416 1826 7476
rect 2268 6416 2382 7476
rect 2824 6416 2938 7476
rect 3380 6416 3494 7476
rect 3936 6416 4050 7476
rect 4492 6416 4606 7476
rect 4942 6416 5056 7476
rect 5498 6416 5612 7476
rect 6054 6416 6168 7476
rect 6610 6416 6724 7476
rect 7166 6416 7280 7476
rect 7722 6416 7836 7476
rect 8278 6416 8392 7476
rect 8834 6416 8948 7476
rect 322 5216 436 6276
rect 878 5216 992 6276
rect 1434 5216 1548 6276
rect 1990 5216 2104 6276
rect 2546 5216 2660 6276
rect 3102 5216 3216 6276
rect 3658 5216 3772 6276
rect 4214 5216 4328 6276
rect 5220 5216 5334 6276
rect 5776 5216 5890 6276
rect 6332 5216 6446 6276
rect 6888 5216 7002 6276
rect 7444 5216 7558 6276
rect 8000 5216 8114 6276
rect 8556 5216 8670 6276
rect 9112 5216 9226 6276
rect 600 4016 714 5076
rect 1156 4016 1270 5076
rect 1712 4016 1826 5076
rect 2268 4016 2382 5076
rect 2824 4016 2938 5076
rect 3380 4016 3494 5076
rect 3936 4016 4050 5076
rect 4492 4016 4606 5076
rect 4942 4016 5056 5076
rect 5498 4016 5612 5076
rect 6054 4016 6168 5076
rect 6610 4016 6724 5076
rect 7166 4016 7280 5076
rect 7722 4016 7836 5076
rect 8278 4016 8392 5076
rect 8834 4016 8948 5076
rect 322 2816 436 3876
rect 878 2816 992 3876
rect 1434 2816 1548 3876
rect 1990 2816 2104 3876
rect 2546 2816 2660 3876
rect 3102 2816 3216 3876
rect 3658 2816 3772 3876
rect 4214 2816 4328 3876
rect 5220 2816 5334 3876
rect 5776 2816 5890 3876
rect 6332 2816 6446 3876
rect 6888 2816 7002 3876
rect 7444 2816 7558 3876
rect 8000 2816 8114 3876
rect 8556 2816 8670 3876
rect 9112 2816 9226 3876
rect 600 1616 714 2676
rect 1156 1616 1270 2676
rect 1712 1616 1826 2676
rect 2268 1616 2382 2676
rect 2824 1616 2938 2676
rect 3380 1616 3494 2676
rect 3936 1616 4050 2676
rect 4492 1616 4606 2676
rect 4942 1616 5056 2676
rect 5498 1616 5612 2676
rect 6054 1616 6168 2676
rect 6610 1616 6724 2676
rect 7166 1616 7280 2676
rect 7722 1616 7836 2676
rect 8278 1616 8392 2676
rect 8834 1616 8948 2676
rect 9585 1696 10425 12203
rect 322 416 436 1476
rect 878 416 992 1476
rect 1434 416 1548 1476
rect 1990 416 2104 1476
rect 2546 416 2660 1476
rect 3102 416 3216 1476
rect 3658 416 3772 1476
rect 4214 416 4328 1476
rect 5220 416 5334 1476
rect 5776 416 5890 1476
rect 6332 416 6446 1476
rect 6888 416 7002 1476
rect 7444 416 7558 1476
rect 8000 416 8114 1476
rect 8556 416 8670 1476
rect 9112 416 9226 1476
<< metal3 >>
rect 302 12276 10525 12296
rect 302 11216 600 12276
rect 714 11216 1156 12276
rect 1270 11216 1712 12276
rect 1826 11216 2268 12276
rect 2382 11216 2824 12276
rect 2938 11216 3380 12276
rect 3494 11216 3936 12276
rect 4050 11216 4492 12276
rect 4606 11216 4942 12276
rect 5056 11216 5498 12276
rect 5612 11216 6054 12276
rect 6168 11216 6610 12276
rect 6724 11216 7166 12276
rect 7280 11216 7722 12276
rect 7836 11216 8278 12276
rect 8392 11216 8834 12276
rect 8948 12203 10525 12276
rect 8948 11216 9585 12203
rect 302 11196 9585 11216
rect -977 11076 9246 11096
rect -977 10997 322 11076
rect -977 496 -877 10997
rect -37 10016 322 10997
rect 436 10016 878 11076
rect 992 10016 1434 11076
rect 1548 10016 1990 11076
rect 2104 10016 2546 11076
rect 2660 10016 3102 11076
rect 3216 10016 3658 11076
rect 3772 10016 4214 11076
rect 4328 10016 5220 11076
rect 5334 10016 5776 11076
rect 5890 10016 6332 11076
rect 6446 10016 6888 11076
rect 7002 10016 7444 11076
rect 7558 10016 8000 11076
rect 8114 10016 8556 11076
rect 8670 10016 9112 11076
rect 9226 10016 9246 11076
rect -37 9996 9246 10016
rect -37 8696 63 9996
rect 9485 9896 9585 11196
rect 302 9876 9585 9896
rect 302 8816 600 9876
rect 714 8816 1156 9876
rect 1270 8816 1712 9876
rect 1826 8816 2268 9876
rect 2382 8816 2824 9876
rect 2938 8816 3380 9876
rect 3494 8816 3936 9876
rect 4050 8816 4492 9876
rect 4606 8816 4942 9876
rect 5056 8816 5498 9876
rect 5612 8816 6054 9876
rect 6168 8816 6610 9876
rect 6724 8816 7166 9876
rect 7280 8816 7722 9876
rect 7836 8816 8278 9876
rect 8392 8816 8834 9876
rect 8948 8816 9585 9876
rect 302 8796 9585 8816
rect -37 8676 9246 8696
rect -37 7616 322 8676
rect 436 7616 878 8676
rect 992 7616 1434 8676
rect 1548 7616 1990 8676
rect 2104 7616 2546 8676
rect 2660 7616 3102 8676
rect 3216 7616 3658 8676
rect 3772 7616 4214 8676
rect 4328 7616 5220 8676
rect 5334 7616 5776 8676
rect 5890 7616 6332 8676
rect 6446 7616 6888 8676
rect 7002 7616 7444 8676
rect 7558 7616 8000 8676
rect 8114 7616 8556 8676
rect 8670 7616 9112 8676
rect 9226 7616 9246 8676
rect -37 7596 9246 7616
rect -37 6296 63 7596
rect 9485 7496 9585 8796
rect 302 7476 9585 7496
rect 302 6416 600 7476
rect 714 6416 1156 7476
rect 1270 6416 1712 7476
rect 1826 6416 2268 7476
rect 2382 6416 2824 7476
rect 2938 6416 3380 7476
rect 3494 6416 3936 7476
rect 4050 6416 4492 7476
rect 4606 6416 4942 7476
rect 5056 6416 5498 7476
rect 5612 6416 6054 7476
rect 6168 6416 6610 7476
rect 6724 6416 7166 7476
rect 7280 6416 7722 7476
rect 7836 6416 8278 7476
rect 8392 6416 8834 7476
rect 8948 6416 9585 7476
rect 302 6396 9585 6416
rect -37 6276 9246 6296
rect -37 5216 322 6276
rect 436 5216 878 6276
rect 992 5216 1434 6276
rect 1548 5216 1990 6276
rect 2104 5216 2546 6276
rect 2660 5216 3102 6276
rect 3216 5216 3658 6276
rect 3772 5216 4214 6276
rect 4328 5216 5220 6276
rect 5334 5216 5776 6276
rect 5890 5216 6332 6276
rect 6446 5216 6888 6276
rect 7002 5216 7444 6276
rect 7558 5216 8000 6276
rect 8114 5216 8556 6276
rect 8670 5216 9112 6276
rect 9226 5216 9246 6276
rect -37 5196 9246 5216
rect -37 3896 63 5196
rect 9485 5096 9585 6396
rect 302 5076 9585 5096
rect 302 4016 600 5076
rect 714 4016 1156 5076
rect 1270 4016 1712 5076
rect 1826 4016 2268 5076
rect 2382 4016 2824 5076
rect 2938 4016 3380 5076
rect 3494 4016 3936 5076
rect 4050 4016 4492 5076
rect 4606 4016 4942 5076
rect 5056 4016 5498 5076
rect 5612 4016 6054 5076
rect 6168 4016 6610 5076
rect 6724 4016 7166 5076
rect 7280 4016 7722 5076
rect 7836 4016 8278 5076
rect 8392 4016 8834 5076
rect 8948 4016 9585 5076
rect 302 3996 9585 4016
rect -37 3876 9246 3896
rect -37 2816 322 3876
rect 436 2816 878 3876
rect 992 2816 1434 3876
rect 1548 2816 1990 3876
rect 2104 2816 2546 3876
rect 2660 2816 3102 3876
rect 3216 2816 3658 3876
rect 3772 2816 4214 3876
rect 4328 2816 5220 3876
rect 5334 2816 5776 3876
rect 5890 2816 6332 3876
rect 6446 2816 6888 3876
rect 7002 2816 7444 3876
rect 7558 2816 8000 3876
rect 8114 2816 8556 3876
rect 8670 2816 9112 3876
rect 9226 2816 9246 3876
rect -37 2796 9246 2816
rect -37 1496 63 2796
rect 9485 2696 9585 3996
rect 302 2676 9585 2696
rect 302 1616 600 2676
rect 714 1616 1156 2676
rect 1270 1616 1712 2676
rect 1826 1616 2268 2676
rect 2382 1616 2824 2676
rect 2938 1616 3380 2676
rect 3494 1616 3936 2676
rect 4050 1616 4492 2676
rect 4606 1616 4942 2676
rect 5056 1616 5498 2676
rect 5612 1616 6054 2676
rect 6168 1616 6610 2676
rect 6724 1616 7166 2676
rect 7280 1616 7722 2676
rect 7836 1616 8278 2676
rect 8392 1616 8834 2676
rect 8948 1696 9585 2676
rect 10425 1696 10525 12203
rect 8948 1616 10525 1696
rect 302 1596 10525 1616
rect -37 1476 9246 1496
rect -37 496 322 1476
rect -977 416 322 496
rect 436 416 878 1476
rect 992 416 1434 1476
rect 1548 416 1990 1476
rect 2104 416 2546 1476
rect 2660 416 3102 1476
rect 3216 416 3658 1476
rect 3772 416 4214 1476
rect 4328 416 5220 1476
rect 5334 416 5776 1476
rect 5890 416 6332 1476
rect 6446 416 6888 1476
rect 7002 416 7444 1476
rect 7558 416 8000 1476
rect 8114 416 8556 1476
rect 8670 416 9112 1476
rect 9226 416 9246 1476
rect -977 396 9246 416
use hvnmos_LAXGBM  hvnmos_LAXGBM_0
timestamp 1753298217
transform 0 1 10011 -1 0 -24
box -268 -272 268 272
use hvpmos_3RBJXJ  hvpmos_3RBJXJ_0
timestamp 1753298217
transform 0 1 10011 -1 0 974
box -592 -374 592 374
use hvpmos_LSUQBM  hvpmos_LSUQBM_0
timestamp 1753041618
transform 1 0 518 0 1 6346
box -518 -6346 4410 6346
use hvpmos_LSUQBM  hvpmos_LSUQBM_1
timestamp 1753041618
transform 1 0 5138 0 1 6346
box -518 -6346 4410 6346
use rhigh_GGS7YG  rhigh_GGS7YG_0
timestamp 1752520737
transform 0 1 4542 -1 0 -283
box -230 -4266 430 4266
<< labels >>
flabel metal3 -977 396 -439 11095 0 FreeSans 800 0 0 0 VDDSW
port 5 nsew
flabel metal3 9987 1597 10525 12296 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 -3 -709 91 -57 0 FreeSans 800 0 0 0 VSS
port 0 nsew
flabel metal1 10154 335 10518 536 0 FreeSans 320 0 0 0 POWERON
port 6 nsew
<< end >>
