magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 1008 834
<< pwell >>
rect 33 56 945 292
rect -26 -56 986 56
<< nmos >>
rect 127 156 153 266
rect 259 118 285 266
rect 356 118 382 266
rect 470 118 496 266
rect 678 118 704 266
rect 784 118 810 266
<< pmos >>
rect 127 412 153 580
rect 259 412 285 612
rect 418 412 444 612
rect 533 412 559 612
rect 678 412 704 612
rect 784 412 810 636
<< ndiff >>
rect 59 202 127 266
rect 59 170 73 202
rect 105 170 127 202
rect 59 156 127 170
rect 153 232 259 266
rect 153 200 181 232
rect 213 200 259 232
rect 153 164 259 200
rect 153 156 181 164
rect 167 132 181 156
rect 213 132 259 164
rect 167 118 259 132
rect 285 118 356 266
rect 382 164 470 266
rect 382 132 412 164
rect 444 132 470 164
rect 382 118 470 132
rect 496 118 678 266
rect 704 164 784 266
rect 704 132 730 164
rect 762 132 784 164
rect 704 118 784 132
rect 810 232 919 266
rect 810 200 866 232
rect 898 200 919 232
rect 810 164 919 200
rect 810 132 866 164
rect 898 132 919 164
rect 810 118 919 132
<< pdiff >>
rect 718 612 784 636
rect 183 598 259 612
rect 183 580 205 598
rect 59 566 127 580
rect 59 534 73 566
rect 105 534 127 566
rect 59 498 127 534
rect 59 466 73 498
rect 105 466 127 498
rect 59 412 127 466
rect 153 566 205 580
rect 237 566 259 598
rect 153 412 259 566
rect 285 412 418 612
rect 444 579 533 612
rect 444 547 470 579
rect 502 547 533 579
rect 444 511 533 547
rect 444 479 470 511
rect 502 479 533 511
rect 444 412 533 479
rect 559 412 678 612
rect 704 596 784 612
rect 704 564 730 596
rect 762 564 784 596
rect 704 526 784 564
rect 704 494 730 526
rect 762 494 784 526
rect 704 458 784 494
rect 704 426 730 458
rect 762 426 784 458
rect 704 412 784 426
rect 810 596 918 636
rect 810 564 866 596
rect 898 564 918 596
rect 810 526 918 564
rect 810 494 866 526
rect 898 494 918 526
rect 810 458 918 494
rect 810 426 866 458
rect 898 426 918 458
rect 810 412 918 426
<< ndiffc >>
rect 73 170 105 202
rect 181 200 213 232
rect 181 132 213 164
rect 412 132 444 164
rect 730 132 762 164
rect 866 200 898 232
rect 866 132 898 164
<< pdiffc >>
rect 73 534 105 566
rect 73 466 105 498
rect 205 566 237 598
rect 470 547 502 579
rect 470 479 502 511
rect 730 564 762 596
rect 730 494 762 526
rect 730 426 762 458
rect 866 564 898 596
rect 866 494 898 526
rect 866 426 898 458
<< psubdiff >>
rect 0 16 960 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 960 16
rect 0 -30 960 -16
<< nsubdiff >>
rect 0 772 960 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 960 772
rect 0 726 960 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
<< poly >>
rect 127 580 153 616
rect 259 612 285 648
rect 418 612 444 648
rect 533 612 559 648
rect 678 612 704 648
rect 784 636 810 672
rect 127 380 153 412
rect 259 380 285 412
rect 127 362 285 380
rect 127 330 141 362
rect 173 330 285 362
rect 418 354 444 412
rect 533 354 559 412
rect 678 374 704 412
rect 678 356 744 374
rect 127 314 285 330
rect 127 266 153 314
rect 259 266 285 314
rect 322 336 382 350
rect 322 304 336 336
rect 368 304 382 336
rect 322 290 382 304
rect 356 266 382 290
rect 418 336 496 354
rect 418 304 434 336
rect 466 304 496 336
rect 418 288 496 304
rect 533 336 599 354
rect 533 304 553 336
rect 585 304 599 336
rect 533 288 599 304
rect 678 324 694 356
rect 726 324 744 356
rect 678 308 744 324
rect 784 370 810 412
rect 784 352 850 370
rect 784 320 802 352
rect 834 320 850 352
rect 470 266 496 288
rect 678 266 704 308
rect 784 304 850 320
rect 784 266 810 304
rect 127 120 153 156
rect 259 82 285 118
rect 356 82 382 118
rect 470 82 496 118
rect 678 82 704 118
rect 784 82 810 118
<< polycont >>
rect 141 330 173 362
rect 336 304 368 336
rect 434 304 466 336
rect 553 304 585 336
rect 694 324 726 356
rect 802 320 834 352
<< metal1 >>
rect 0 772 960 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 960 772
rect 0 712 960 740
rect 195 598 247 712
rect 59 566 115 576
rect 59 534 73 566
rect 105 534 115 566
rect 195 566 205 598
rect 237 566 247 598
rect 195 556 247 566
rect 296 625 685 659
rect 59 520 115 534
rect 296 520 328 625
rect 59 498 328 520
rect 460 579 512 589
rect 460 547 470 579
rect 502 547 512 579
rect 460 511 512 547
rect 460 501 470 511
rect 59 466 73 498
rect 105 488 328 498
rect 105 466 115 488
rect 59 456 115 466
rect 371 479 470 501
rect 502 479 512 511
rect 371 469 512 479
rect 59 212 91 456
rect 371 452 403 469
rect 257 416 403 452
rect 127 362 221 374
rect 127 330 141 362
rect 173 330 221 362
rect 127 300 221 330
rect 171 232 218 242
rect 59 202 115 212
rect 59 170 73 202
rect 105 170 115 202
rect 59 160 115 170
rect 171 200 181 232
rect 213 200 218 232
rect 171 164 218 200
rect 171 132 181 164
rect 213 132 218 164
rect 171 44 218 132
rect 257 166 290 416
rect 326 336 378 346
rect 326 304 336 336
rect 368 304 378 336
rect 326 294 378 304
rect 342 240 378 294
rect 424 336 507 384
rect 424 304 434 336
rect 466 304 507 336
rect 424 280 507 304
rect 543 336 603 384
rect 543 304 553 336
rect 585 304 603 336
rect 650 374 685 625
rect 726 596 766 712
rect 726 564 730 596
rect 762 564 766 596
rect 726 526 766 564
rect 726 494 730 526
rect 762 494 766 526
rect 726 458 766 494
rect 726 426 730 458
rect 762 426 766 458
rect 726 416 766 426
rect 827 596 918 640
rect 827 564 866 596
rect 898 564 918 596
rect 827 526 918 564
rect 827 494 866 526
rect 898 494 918 526
rect 827 458 918 494
rect 827 426 866 458
rect 898 426 918 458
rect 827 408 918 426
rect 650 356 744 374
rect 650 324 694 356
rect 726 324 744 356
rect 650 308 744 324
rect 789 352 844 370
rect 789 320 802 352
rect 834 320 844 352
rect 543 240 603 304
rect 789 304 844 320
rect 789 240 827 304
rect 880 242 918 408
rect 342 206 603 240
rect 639 206 827 240
rect 863 232 918 242
rect 639 166 673 206
rect 863 200 866 232
rect 898 200 918 232
rect 257 164 673 166
rect 257 132 412 164
rect 444 132 673 164
rect 257 122 673 132
rect 720 164 772 169
rect 720 132 730 164
rect 762 132 772 164
rect 720 44 772 132
rect 863 164 918 200
rect 863 132 866 164
rect 898 132 918 164
rect 863 114 918 132
rect 0 16 960 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 960 16
rect 0 -44 960 -16
<< labels >>
flabel metal1 s 543 206 603 384 0 FreeSans 400 0 0 0 A1
port 2 nsew
flabel metal1 s 827 408 918 640 0 FreeSans 400 0 0 0 X
port 3 nsew
flabel metal1 s 127 300 221 374 0 FreeSans 400 0 0 0 S
port 4 nsew
flabel metal1 s 0 712 960 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -44 960 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 424 280 507 384 0 FreeSans 400 0 0 0 A0
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 960 756
string GDS_END 207100
string GDS_FILE 6_final.gds
string GDS_START 200088
<< end >>
