magic
tech ihp-sg13g2
timestamp 1748543940
<< error_p >>
rect -23 265 23 291
rect 45 265 91 291
rect 113 265 159 291
rect 181 265 227 291
rect 249 265 295 291
rect 317 265 363 291
rect 385 265 431 291
rect 453 265 499 291
rect 521 265 567 291
rect 589 265 635 291
rect -23 -291 23 -265
rect 45 -291 91 -265
rect 113 -291 159 -265
rect 181 -291 227 -265
rect 249 -291 295 -265
rect 317 -291 363 -265
rect 385 -291 431 -265
rect 453 -291 499 -265
rect 521 -291 567 -265
rect 589 -291 635 -265
<< psubdiff >>
rect -115 376 727 383
rect -115 360 -78 376
rect 690 360 727 376
rect -115 353 727 360
rect -115 346 -85 353
rect -115 -346 -108 346
rect -92 -346 -85 346
rect 697 346 727 353
rect -115 -353 -85 -346
rect 697 -346 704 346
rect 720 -346 727 346
rect 697 -353 727 -346
rect -115 -360 727 -353
rect -115 -376 -78 -360
rect 690 -376 727 -360
rect -115 -383 727 -376
<< psubdiffcont >>
rect -78 360 690 376
rect -108 -346 -92 346
rect 704 -346 720 346
rect -78 -376 690 -360
<< poly >>
rect -25 286 25 293
rect -25 270 -18 286
rect 18 270 25 286
rect -25 250 25 270
rect -25 -270 25 -250
rect -25 -286 -18 -270
rect 18 -286 25 -270
rect -25 -293 25 -286
rect 43 286 93 293
rect 43 270 50 286
rect 86 270 93 286
rect 43 250 93 270
rect 43 -270 93 -250
rect 43 -286 50 -270
rect 86 -286 93 -270
rect 43 -293 93 -286
rect 111 286 161 293
rect 111 270 118 286
rect 154 270 161 286
rect 111 250 161 270
rect 111 -270 161 -250
rect 111 -286 118 -270
rect 154 -286 161 -270
rect 111 -293 161 -286
rect 179 286 229 293
rect 179 270 186 286
rect 222 270 229 286
rect 179 250 229 270
rect 179 -270 229 -250
rect 179 -286 186 -270
rect 222 -286 229 -270
rect 179 -293 229 -286
rect 247 286 297 293
rect 247 270 254 286
rect 290 270 297 286
rect 247 250 297 270
rect 247 -270 297 -250
rect 247 -286 254 -270
rect 290 -286 297 -270
rect 247 -293 297 -286
rect 315 286 365 293
rect 315 270 322 286
rect 358 270 365 286
rect 315 250 365 270
rect 315 -270 365 -250
rect 315 -286 322 -270
rect 358 -286 365 -270
rect 315 -293 365 -286
rect 383 286 433 293
rect 383 270 390 286
rect 426 270 433 286
rect 383 250 433 270
rect 383 -270 433 -250
rect 383 -286 390 -270
rect 426 -286 433 -270
rect 383 -293 433 -286
rect 451 286 501 293
rect 451 270 458 286
rect 494 270 501 286
rect 451 250 501 270
rect 451 -270 501 -250
rect 451 -286 458 -270
rect 494 -286 501 -270
rect 451 -293 501 -286
rect 519 286 569 293
rect 519 270 526 286
rect 562 270 569 286
rect 519 250 569 270
rect 519 -270 569 -250
rect 519 -286 526 -270
rect 562 -286 569 -270
rect 519 -293 569 -286
rect 587 286 637 293
rect 587 270 594 286
rect 630 270 637 286
rect 587 250 637 270
rect 587 -270 637 -250
rect 587 -286 594 -270
rect 630 -286 637 -270
rect 587 -293 637 -286
<< polycont >>
rect -18 270 18 286
rect -18 -286 18 -270
rect 50 270 86 286
rect 50 -286 86 -270
rect 118 270 154 286
rect 118 -286 154 -270
rect 186 270 222 286
rect 186 -286 222 -270
rect 254 270 290 286
rect 254 -286 290 -270
rect 322 270 358 286
rect 322 -286 358 -270
rect 390 270 426 286
rect 390 -286 426 -270
rect 458 270 494 286
rect 458 -286 494 -270
rect 526 270 562 286
rect 526 -286 562 -270
rect 594 270 630 286
rect 594 -286 630 -270
<< xpolyres >>
rect -25 -250 25 250
rect 43 -250 93 250
rect 111 -250 161 250
rect 179 -250 229 250
rect 247 -250 297 250
rect 315 -250 365 250
rect 383 -250 433 250
rect 451 -250 501 250
rect 519 -250 569 250
rect 587 -250 637 250
<< metal1 >>
rect -113 376 725 381
rect -113 360 -78 376
rect 690 360 725 376
rect -113 355 725 360
rect -113 346 -87 355
rect -113 -346 -108 346
rect -92 -346 -87 346
rect 699 346 725 355
rect -113 -355 -87 -346
rect 699 -346 704 346
rect 720 -346 725 346
rect 699 -355 725 -346
rect -113 -360 725 -355
rect -113 -376 -78 -360
rect 690 -376 725 -360
rect -113 -381 725 -376
<< properties >>
string gencell rhigh
string library sg13g2_devstdin
string parameters w 0.5 l 5 nx 10 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class resistor endcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
