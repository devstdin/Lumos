magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752439852
<< error_p >>
rect -16 357 -6 367
rect 6 357 16 367
rect -26 347 26 357
rect -16 335 16 347
rect -26 325 26 335
rect -16 315 -6 325
rect 6 315 16 325
rect -67 261 -57 271
rect -45 261 -35 271
rect 35 261 45 271
rect 57 261 67 271
rect -77 251 -67 261
rect -35 251 -25 261
rect 25 251 35 261
rect 67 251 77 261
rect -77 -261 -67 -251
rect -35 -261 -25 -251
rect 25 -261 35 -251
rect 67 -261 77 -251
rect -67 -271 -57 -261
rect -45 -271 -35 -261
rect 35 -271 45 -261
rect 57 -271 67 -261
rect -16 -325 -6 -315
rect 6 -325 16 -315
rect -26 -335 26 -325
rect -16 -347 16 -335
rect -26 -357 26 -347
rect -16 -367 -6 -357
rect 6 -367 16 -357
<< nmos >>
rect -13 -275 13 275
<< ndiff >>
rect -81 261 -13 275
rect -81 -261 -67 261
rect -35 -261 -13 261
rect -81 -275 -13 -261
rect 13 261 81 275
rect 13 -261 35 261
rect 67 -261 81 261
rect 13 -275 81 -261
<< ndiffc >>
rect -67 -261 -35 261
rect 35 -261 67 261
<< psubdiff >>
rect -183 445 183 459
rect -183 413 -109 445
rect 109 413 183 445
rect -183 399 183 413
rect -183 385 -123 399
rect -183 -385 -169 385
rect -137 -385 -123 385
rect 123 385 183 399
rect -183 -399 -123 -385
rect 123 -385 137 385
rect 169 -385 183 385
rect 123 -399 183 -385
rect -183 -413 183 -399
rect -183 -445 -109 -413
rect 109 -445 183 -413
rect -183 -459 183 -445
<< psubdiffcont >>
rect -109 413 109 445
rect -169 -385 -137 385
rect 137 -385 169 385
rect -109 -445 109 -413
<< poly >>
rect -30 357 30 371
rect -30 325 -16 357
rect 16 325 30 357
rect -30 311 30 325
rect -13 275 13 311
rect -13 -311 13 -275
rect -30 -325 30 -311
rect -30 -357 -16 -325
rect 16 -357 30 -325
rect -30 -371 30 -357
<< polycont >>
rect -16 325 16 357
rect -16 -357 16 -325
<< metal1 >>
rect -179 445 179 455
rect -179 413 -109 445
rect 109 413 179 445
rect -179 403 179 413
rect -179 385 -127 403
rect -179 -385 -169 385
rect -137 -385 -127 385
rect 127 385 179 403
rect -179 -403 -127 -385
rect 127 -385 137 385
rect 169 -385 179 385
rect 127 -403 179 -385
rect -179 -413 179 -403
rect -179 -445 -109 -413
rect 109 -445 179 -413
rect -179 -455 179 -445
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 2.75 l 0.13 nf 1 nx 1 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
