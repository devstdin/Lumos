magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752864670
<< error_p >>
rect -36 160 -26 170
rect 26 160 36 170
rect 242 160 252 170
rect 304 160 314 170
rect -46 150 46 160
rect 232 150 324 160
rect -36 138 36 150
rect 242 138 314 150
rect -46 128 46 138
rect 232 128 324 138
rect -36 118 -26 128
rect 26 118 36 128
rect 242 118 252 128
rect 304 118 314 128
rect -104 86 -94 96
rect -82 86 -72 96
rect 72 86 82 96
rect 94 86 104 96
rect 174 86 184 96
rect 196 86 206 96
rect 350 86 360 96
rect 372 86 382 96
rect -114 76 -104 86
rect -72 76 -62 86
rect 62 76 72 86
rect 104 76 114 86
rect 164 76 174 86
rect 206 76 216 86
rect 340 76 350 86
rect 382 76 392 86
rect -114 -86 -104 -76
rect -72 -86 -62 -76
rect 62 -86 72 -76
rect 104 -86 114 -76
rect 164 -86 174 -76
rect 206 -86 216 -76
rect 340 -86 350 -76
rect 382 -86 392 -76
rect -104 -96 -94 -86
rect -82 -96 -72 -86
rect 72 -96 82 -86
rect 94 -96 104 -86
rect 174 -96 184 -86
rect 196 -96 206 -86
rect 350 -96 360 -86
rect 372 -96 382 -86
rect -36 -128 -26 -118
rect 26 -128 36 -118
rect 242 -128 252 -118
rect 304 -128 314 -118
rect -46 -138 46 -128
rect 232 -138 324 -128
rect -36 -150 36 -138
rect 242 -150 314 -138
rect -46 -160 46 -150
rect 232 -160 324 -150
rect -36 -170 -26 -160
rect 26 -170 36 -160
rect 242 -170 252 -160
rect 304 -170 314 -160
<< nmos >>
rect -50 -100 50 100
rect 228 -100 328 100
<< ndiff >>
rect -118 86 -50 100
rect -118 -86 -104 86
rect -72 -86 -50 86
rect -118 -100 -50 -86
rect 50 86 118 100
rect 50 -86 72 86
rect 104 -86 118 86
rect 50 -100 118 -86
rect 160 86 228 100
rect 160 -86 174 86
rect 206 -86 228 86
rect 160 -100 228 -86
rect 328 86 396 100
rect 328 -86 350 86
rect 382 -86 396 86
rect 328 -100 396 -86
<< ndiffc >>
rect -104 -86 -72 86
rect 72 -86 104 86
rect 174 -86 206 86
rect 350 -86 382 86
<< psubdiff >>
rect -241 262 519 276
rect -241 230 -167 262
rect 445 230 519 262
rect -241 216 519 230
rect -241 202 -181 216
rect -241 -202 -227 202
rect -195 -202 -181 202
rect 459 202 519 216
rect -241 -216 -181 -202
rect 459 -202 473 202
rect 505 -202 519 202
rect 459 -216 519 -202
rect -241 -230 519 -216
rect -241 -262 -167 -230
rect 445 -262 519 -230
rect -241 -276 519 -262
<< psubdiffcont >>
rect -167 230 445 262
rect -227 -202 -195 202
rect 473 -202 505 202
rect -167 -262 445 -230
<< poly >>
rect -50 160 50 174
rect -50 128 -36 160
rect 36 128 50 160
rect -50 100 50 128
rect 228 160 328 174
rect 228 128 242 160
rect 314 128 328 160
rect 228 100 328 128
rect -50 -128 50 -100
rect -50 -160 -36 -128
rect 36 -160 50 -128
rect -50 -174 50 -160
rect 228 -128 328 -100
rect 228 -160 242 -128
rect 314 -160 328 -128
rect 228 -174 328 -160
<< polycont >>
rect -36 128 36 160
rect 242 128 314 160
rect -36 -160 36 -128
rect 242 -160 314 -128
<< metal1 >>
rect -237 262 515 272
rect -237 230 -167 262
rect 445 230 515 262
rect -237 220 515 230
rect -237 202 -185 220
rect -237 -202 -227 202
rect -195 -202 -185 202
rect 463 202 515 220
rect -237 -220 -185 -202
rect 463 -202 473 202
rect 505 -202 515 202
rect 463 -220 515 -202
rect -237 -230 515 -220
rect -237 -262 -167 -230
rect 445 -262 515 -230
rect -237 -272 515 -262
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 1 l 0.5 nf 1 nx 2 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 1
<< end >>
