magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2100 -924 2300 37600
<< nwell >>
rect -48 33246 248 33554
rect -100 29546 300 29854
rect -48 1076 248 12324
<< pwell >>
rect 44 31456 156 31524
rect 18 31344 182 31456
rect 44 31072 156 31344
rect 18 12974 182 28060
<< psubdiff >>
rect 84 31384 116 31416
rect 84 31316 116 31348
rect 84 31248 116 31280
rect 84 31180 116 31212
rect 84 31112 116 31144
rect 84 27899 116 27931
rect 84 27831 116 27863
rect 84 27763 116 27795
rect 84 27695 116 27727
rect 84 27627 116 27659
rect 84 27559 116 27591
rect 84 27491 116 27523
rect 84 27423 116 27455
rect 84 27355 116 27387
rect 84 27287 116 27319
rect 84 27219 116 27251
rect 84 27151 116 27183
rect 84 27083 116 27115
rect 84 27015 116 27047
rect 84 26947 116 26979
rect 84 26879 116 26911
rect 84 26811 116 26843
rect 84 26743 116 26775
rect 84 26675 116 26707
rect 84 26607 116 26639
rect 84 26539 116 26571
rect 84 26471 116 26503
rect 84 26403 116 26435
rect 84 26335 116 26367
rect 84 26267 116 26299
rect 84 26199 116 26231
rect 84 26131 116 26163
rect 84 26063 116 26095
rect 84 25995 116 26027
rect 84 25927 116 25959
rect 84 25859 116 25891
rect 84 25791 116 25823
rect 84 25723 116 25755
rect 84 25655 116 25687
rect 84 25587 116 25619
rect 84 25519 116 25551
rect 84 25451 116 25483
rect 84 25383 116 25415
rect 84 25315 116 25347
rect 84 25247 116 25279
rect 84 25179 116 25211
rect 84 25111 116 25143
rect 84 25043 116 25075
rect 84 24975 116 25007
rect 84 24907 116 24939
rect 84 24839 116 24871
rect 84 24771 116 24803
rect 84 24703 116 24735
rect 84 24635 116 24667
rect 84 24567 116 24599
rect 84 24499 116 24531
rect 84 24431 116 24463
rect 84 24363 116 24395
rect 84 24295 116 24327
rect 84 24227 116 24259
rect 84 24159 116 24191
rect 84 24091 116 24123
rect 84 24023 116 24055
rect 84 23955 116 23987
rect 84 23887 116 23919
rect 84 23819 116 23851
rect 84 23751 116 23783
rect 84 23683 116 23715
rect 84 23615 116 23647
rect 84 23547 116 23579
rect 84 23479 116 23511
rect 84 23411 116 23443
rect 84 23343 116 23375
rect 84 23275 116 23307
rect 84 23207 116 23239
rect 84 22788 116 22820
rect 84 22720 116 22752
rect 84 22652 116 22684
rect 84 22584 116 22616
rect 84 22516 116 22548
rect 84 22448 116 22480
rect 84 22380 116 22412
rect 84 22312 116 22344
rect 84 22244 116 22276
rect 84 22176 116 22208
rect 84 22108 116 22140
rect 84 22040 116 22072
rect 84 21972 116 22004
rect 84 21904 116 21936
rect 84 21836 116 21868
rect 84 21768 116 21800
rect 84 21700 116 21732
rect 84 21632 116 21664
rect 84 21564 116 21596
rect 84 21496 116 21528
rect 84 21428 116 21460
rect 84 21360 116 21392
rect 84 21292 116 21324
rect 84 21224 116 21256
rect 84 21156 116 21188
rect 84 21088 116 21120
rect 84 21020 116 21052
rect 84 20952 116 20984
rect 84 20884 116 20916
rect 84 20816 116 20848
rect 84 20748 116 20780
rect 84 20680 116 20712
rect 84 20612 116 20644
rect 84 20544 116 20576
rect 84 20476 116 20508
rect 84 20408 116 20440
rect 84 20340 116 20372
rect 84 20272 116 20304
rect 84 20204 116 20236
rect 84 20136 116 20168
rect 84 20068 116 20100
rect 84 20000 116 20032
rect 84 19932 116 19964
rect 84 19864 116 19896
rect 84 19796 116 19828
rect 84 19728 116 19760
rect 84 19660 116 19692
rect 84 19592 116 19624
rect 84 19524 116 19556
rect 84 19456 116 19488
rect 84 19388 116 19420
rect 84 19320 116 19352
rect 84 19252 116 19284
rect 84 19184 116 19216
rect 84 19116 116 19148
rect 84 19048 116 19080
rect 84 18980 116 19012
rect 84 18912 116 18944
rect 84 18844 116 18876
rect 84 18776 116 18808
rect 84 18708 116 18740
rect 84 18640 116 18672
rect 84 18572 116 18604
rect 84 18504 116 18536
rect 84 18436 116 18468
rect 84 18368 116 18400
rect 84 18300 116 18332
rect 84 18232 116 18264
rect 84 18164 116 18196
rect 84 17770 116 17802
rect 84 17702 116 17734
rect 84 17634 116 17666
rect 84 17566 116 17598
rect 84 17498 116 17530
rect 84 17430 116 17462
rect 84 17362 116 17394
rect 84 17294 116 17326
rect 84 17226 116 17258
rect 84 17158 116 17190
rect 84 17090 116 17122
rect 84 17022 116 17054
rect 84 16954 116 16986
rect 84 16886 116 16918
rect 84 16818 116 16850
rect 84 16750 116 16782
rect 84 16682 116 16714
rect 84 16614 116 16646
rect 84 16546 116 16578
rect 84 16478 116 16510
rect 84 16410 116 16442
rect 84 16342 116 16374
rect 84 16274 116 16306
rect 84 16206 116 16238
rect 84 16138 116 16170
rect 84 16070 116 16102
rect 84 16002 116 16034
rect 84 15934 116 15966
rect 84 15866 116 15898
rect 84 15798 116 15830
rect 84 15730 116 15762
rect 84 15662 116 15694
rect 84 15594 116 15626
rect 84 15526 116 15558
rect 84 15458 116 15490
rect 84 15390 116 15422
rect 84 15322 116 15354
rect 84 15254 116 15286
rect 84 15186 116 15218
rect 84 15118 116 15150
rect 84 15050 116 15082
rect 84 14982 116 15014
rect 84 14914 116 14946
rect 84 14846 116 14878
rect 84 14778 116 14810
rect 84 14710 116 14742
rect 84 14642 116 14674
rect 84 14574 116 14606
rect 84 14506 116 14538
rect 84 14438 116 14470
rect 84 14370 116 14402
rect 84 14302 116 14334
rect 84 14234 116 14266
rect 84 14166 116 14198
rect 84 14098 116 14130
rect 84 14030 116 14062
rect 84 13962 116 13994
rect 84 13894 116 13926
rect 84 13826 116 13858
rect 84 13758 116 13790
rect 84 13690 116 13722
rect 84 13622 116 13654
rect 84 13554 116 13586
rect 84 13486 116 13518
rect 84 13418 116 13450
rect 84 13350 116 13382
rect 84 13282 116 13314
rect 84 13214 116 13246
rect 84 13146 116 13178
rect 84 13078 116 13110
rect 70 31484 130 31498
rect 70 31452 84 31484
rect 116 31452 130 31484
rect 70 31430 130 31452
rect 44 31416 156 31430
rect 44 31384 84 31416
rect 116 31384 156 31416
rect 44 31370 156 31384
rect 70 31348 130 31370
rect 70 31316 84 31348
rect 116 31316 130 31348
rect 70 31280 130 31316
rect 70 31248 84 31280
rect 116 31248 130 31280
rect 70 31212 130 31248
rect 70 31180 84 31212
rect 116 31180 130 31212
rect 70 31144 130 31180
rect 70 31112 84 31144
rect 116 31112 130 31144
rect 70 31098 130 31112
rect 44 27999 156 28034
rect 44 27967 84 27999
rect 116 27967 156 27999
rect 44 27931 156 27967
rect 44 27899 84 27931
rect 116 27899 156 27931
rect 44 27863 156 27899
rect 44 27831 84 27863
rect 116 27831 156 27863
rect 44 27795 156 27831
rect 44 27763 84 27795
rect 116 27763 156 27795
rect 44 27727 156 27763
rect 44 27695 84 27727
rect 116 27695 156 27727
rect 44 27659 156 27695
rect 44 27627 84 27659
rect 116 27627 156 27659
rect 44 27591 156 27627
rect 44 27559 84 27591
rect 116 27559 156 27591
rect 44 27523 156 27559
rect 44 27491 84 27523
rect 116 27491 156 27523
rect 44 27455 156 27491
rect 44 27423 84 27455
rect 116 27423 156 27455
rect 44 27387 156 27423
rect 44 27355 84 27387
rect 116 27355 156 27387
rect 44 27319 156 27355
rect 44 27287 84 27319
rect 116 27287 156 27319
rect 44 27251 156 27287
rect 44 27219 84 27251
rect 116 27219 156 27251
rect 44 27183 156 27219
rect 44 27151 84 27183
rect 116 27151 156 27183
rect 44 27115 156 27151
rect 44 27083 84 27115
rect 116 27083 156 27115
rect 44 27047 156 27083
rect 44 27015 84 27047
rect 116 27015 156 27047
rect 44 26979 156 27015
rect 44 26947 84 26979
rect 116 26947 156 26979
rect 44 26911 156 26947
rect 44 26879 84 26911
rect 116 26879 156 26911
rect 44 26843 156 26879
rect 44 26811 84 26843
rect 116 26811 156 26843
rect 44 26775 156 26811
rect 44 26743 84 26775
rect 116 26743 156 26775
rect 44 26707 156 26743
rect 44 26675 84 26707
rect 116 26675 156 26707
rect 44 26639 156 26675
rect 44 26607 84 26639
rect 116 26607 156 26639
rect 44 26571 156 26607
rect 44 26539 84 26571
rect 116 26539 156 26571
rect 44 26503 156 26539
rect 44 26471 84 26503
rect 116 26471 156 26503
rect 44 26435 156 26471
rect 44 26403 84 26435
rect 116 26403 156 26435
rect 44 26367 156 26403
rect 44 26335 84 26367
rect 116 26335 156 26367
rect 44 26299 156 26335
rect 44 26267 84 26299
rect 116 26267 156 26299
rect 44 26231 156 26267
rect 44 26199 84 26231
rect 116 26199 156 26231
rect 44 26163 156 26199
rect 44 26131 84 26163
rect 116 26131 156 26163
rect 44 26095 156 26131
rect 44 26063 84 26095
rect 116 26063 156 26095
rect 44 26027 156 26063
rect 44 25995 84 26027
rect 116 25995 156 26027
rect 44 25959 156 25995
rect 44 25927 84 25959
rect 116 25927 156 25959
rect 44 25891 156 25927
rect 44 25859 84 25891
rect 116 25859 156 25891
rect 44 25823 156 25859
rect 44 25791 84 25823
rect 116 25791 156 25823
rect 44 25755 156 25791
rect 44 25723 84 25755
rect 116 25723 156 25755
rect 44 25687 156 25723
rect 44 25655 84 25687
rect 116 25655 156 25687
rect 44 25619 156 25655
rect 44 25587 84 25619
rect 116 25587 156 25619
rect 44 25551 156 25587
rect 44 25519 84 25551
rect 116 25519 156 25551
rect 44 25483 156 25519
rect 44 25451 84 25483
rect 116 25451 156 25483
rect 44 25415 156 25451
rect 44 25383 84 25415
rect 116 25383 156 25415
rect 44 25347 156 25383
rect 44 25315 84 25347
rect 116 25315 156 25347
rect 44 25279 156 25315
rect 44 25247 84 25279
rect 116 25247 156 25279
rect 44 25211 156 25247
rect 44 25179 84 25211
rect 116 25179 156 25211
rect 44 25143 156 25179
rect 44 25111 84 25143
rect 116 25111 156 25143
rect 44 25075 156 25111
rect 44 25043 84 25075
rect 116 25043 156 25075
rect 44 25007 156 25043
rect 44 24975 84 25007
rect 116 24975 156 25007
rect 44 24939 156 24975
rect 44 24907 84 24939
rect 116 24907 156 24939
rect 44 24871 156 24907
rect 44 24839 84 24871
rect 116 24839 156 24871
rect 44 24803 156 24839
rect 44 24771 84 24803
rect 116 24771 156 24803
rect 44 24735 156 24771
rect 44 24703 84 24735
rect 116 24703 156 24735
rect 44 24667 156 24703
rect 44 24635 84 24667
rect 116 24635 156 24667
rect 44 24599 156 24635
rect 44 24567 84 24599
rect 116 24567 156 24599
rect 44 24531 156 24567
rect 44 24499 84 24531
rect 116 24499 156 24531
rect 44 24463 156 24499
rect 44 24431 84 24463
rect 116 24431 156 24463
rect 44 24395 156 24431
rect 44 24363 84 24395
rect 116 24363 156 24395
rect 44 24327 156 24363
rect 44 24295 84 24327
rect 116 24295 156 24327
rect 44 24259 156 24295
rect 44 24227 84 24259
rect 116 24227 156 24259
rect 44 24191 156 24227
rect 44 24159 84 24191
rect 116 24159 156 24191
rect 44 24123 156 24159
rect 44 24091 84 24123
rect 116 24091 156 24123
rect 44 24055 156 24091
rect 44 24023 84 24055
rect 116 24023 156 24055
rect 44 23987 156 24023
rect 44 23955 84 23987
rect 116 23955 156 23987
rect 44 23919 156 23955
rect 44 23887 84 23919
rect 116 23887 156 23919
rect 44 23851 156 23887
rect 44 23819 84 23851
rect 116 23819 156 23851
rect 44 23783 156 23819
rect 44 23751 84 23783
rect 116 23751 156 23783
rect 44 23715 156 23751
rect 44 23683 84 23715
rect 116 23683 156 23715
rect 44 23647 156 23683
rect 44 23615 84 23647
rect 116 23615 156 23647
rect 44 23579 156 23615
rect 44 23547 84 23579
rect 116 23547 156 23579
rect 44 23511 156 23547
rect 44 23479 84 23511
rect 116 23479 156 23511
rect 44 23443 156 23479
rect 44 23411 84 23443
rect 116 23411 156 23443
rect 44 23375 156 23411
rect 44 23343 84 23375
rect 116 23343 156 23375
rect 44 23307 156 23343
rect 44 23275 84 23307
rect 116 23275 156 23307
rect 44 23239 156 23275
rect 44 23207 84 23239
rect 116 23207 156 23239
rect 44 23124 156 23207
rect 44 22888 156 22924
rect 44 22856 84 22888
rect 116 22856 156 22888
rect 44 22820 156 22856
rect 44 22788 84 22820
rect 116 22788 156 22820
rect 44 22752 156 22788
rect 44 22720 84 22752
rect 116 22720 156 22752
rect 44 22684 156 22720
rect 44 22652 84 22684
rect 116 22652 156 22684
rect 44 22616 156 22652
rect 44 22584 84 22616
rect 116 22584 156 22616
rect 44 22548 156 22584
rect 44 22516 84 22548
rect 116 22516 156 22548
rect 44 22480 156 22516
rect 44 22448 84 22480
rect 116 22448 156 22480
rect 44 22412 156 22448
rect 44 22380 84 22412
rect 116 22380 156 22412
rect 44 22344 156 22380
rect 44 22312 84 22344
rect 116 22312 156 22344
rect 44 22276 156 22312
rect 44 22244 84 22276
rect 116 22244 156 22276
rect 44 22208 156 22244
rect 44 22176 84 22208
rect 116 22176 156 22208
rect 44 22140 156 22176
rect 44 22108 84 22140
rect 116 22108 156 22140
rect 44 22072 156 22108
rect 44 22040 84 22072
rect 116 22040 156 22072
rect 44 22004 156 22040
rect 44 21972 84 22004
rect 116 21972 156 22004
rect 44 21936 156 21972
rect 44 21904 84 21936
rect 116 21904 156 21936
rect 44 21868 156 21904
rect 44 21836 84 21868
rect 116 21836 156 21868
rect 44 21800 156 21836
rect 44 21768 84 21800
rect 116 21768 156 21800
rect 44 21732 156 21768
rect 44 21700 84 21732
rect 116 21700 156 21732
rect 44 21664 156 21700
rect 44 21632 84 21664
rect 116 21632 156 21664
rect 44 21596 156 21632
rect 44 21564 84 21596
rect 116 21564 156 21596
rect 44 21528 156 21564
rect 44 21496 84 21528
rect 116 21496 156 21528
rect 44 21460 156 21496
rect 44 21428 84 21460
rect 116 21428 156 21460
rect 44 21392 156 21428
rect 44 21360 84 21392
rect 116 21360 156 21392
rect 44 21324 156 21360
rect 44 21292 84 21324
rect 116 21292 156 21324
rect 44 21256 156 21292
rect 44 21224 84 21256
rect 116 21224 156 21256
rect 44 21188 156 21224
rect 44 21156 84 21188
rect 116 21156 156 21188
rect 44 21120 156 21156
rect 44 21088 84 21120
rect 116 21088 156 21120
rect 44 21052 156 21088
rect 44 21020 84 21052
rect 116 21020 156 21052
rect 44 20984 156 21020
rect 44 20952 84 20984
rect 116 20952 156 20984
rect 44 20916 156 20952
rect 44 20884 84 20916
rect 116 20884 156 20916
rect 44 20848 156 20884
rect 44 20816 84 20848
rect 116 20816 156 20848
rect 44 20780 156 20816
rect 44 20748 84 20780
rect 116 20748 156 20780
rect 44 20712 156 20748
rect 44 20680 84 20712
rect 116 20680 156 20712
rect 44 20644 156 20680
rect 44 20612 84 20644
rect 116 20612 156 20644
rect 44 20576 156 20612
rect 44 20544 84 20576
rect 116 20544 156 20576
rect 44 20508 156 20544
rect 44 20476 84 20508
rect 116 20476 156 20508
rect 44 20440 156 20476
rect 44 20408 84 20440
rect 116 20408 156 20440
rect 44 20372 156 20408
rect 44 20340 84 20372
rect 116 20340 156 20372
rect 44 20304 156 20340
rect 44 20272 84 20304
rect 116 20272 156 20304
rect 44 20236 156 20272
rect 44 20204 84 20236
rect 116 20204 156 20236
rect 44 20168 156 20204
rect 44 20136 84 20168
rect 116 20136 156 20168
rect 44 20100 156 20136
rect 44 20068 84 20100
rect 116 20068 156 20100
rect 44 20032 156 20068
rect 44 20000 84 20032
rect 116 20000 156 20032
rect 44 19964 156 20000
rect 44 19932 84 19964
rect 116 19932 156 19964
rect 44 19896 156 19932
rect 44 19864 84 19896
rect 116 19864 156 19896
rect 44 19828 156 19864
rect 44 19796 84 19828
rect 116 19796 156 19828
rect 44 19760 156 19796
rect 44 19728 84 19760
rect 116 19728 156 19760
rect 44 19692 156 19728
rect 44 19660 84 19692
rect 116 19660 156 19692
rect 44 19624 156 19660
rect 44 19592 84 19624
rect 116 19592 156 19624
rect 44 19556 156 19592
rect 44 19524 84 19556
rect 116 19524 156 19556
rect 44 19488 156 19524
rect 44 19456 84 19488
rect 116 19456 156 19488
rect 44 19420 156 19456
rect 44 19388 84 19420
rect 116 19388 156 19420
rect 44 19352 156 19388
rect 44 19320 84 19352
rect 116 19320 156 19352
rect 44 19284 156 19320
rect 44 19252 84 19284
rect 116 19252 156 19284
rect 44 19216 156 19252
rect 44 19184 84 19216
rect 116 19184 156 19216
rect 44 19148 156 19184
rect 44 19116 84 19148
rect 116 19116 156 19148
rect 44 19080 156 19116
rect 44 19048 84 19080
rect 116 19048 156 19080
rect 44 19012 156 19048
rect 44 18980 84 19012
rect 116 18980 156 19012
rect 44 18944 156 18980
rect 44 18912 84 18944
rect 116 18912 156 18944
rect 44 18876 156 18912
rect 44 18844 84 18876
rect 116 18844 156 18876
rect 44 18808 156 18844
rect 44 18776 84 18808
rect 116 18776 156 18808
rect 44 18740 156 18776
rect 44 18708 84 18740
rect 116 18708 156 18740
rect 44 18672 156 18708
rect 44 18640 84 18672
rect 116 18640 156 18672
rect 44 18604 156 18640
rect 44 18572 84 18604
rect 116 18572 156 18604
rect 44 18536 156 18572
rect 44 18504 84 18536
rect 116 18504 156 18536
rect 44 18468 156 18504
rect 44 18436 84 18468
rect 116 18436 156 18468
rect 44 18400 156 18436
rect 44 18368 84 18400
rect 116 18368 156 18400
rect 44 18332 156 18368
rect 44 18300 84 18332
rect 116 18300 156 18332
rect 44 18264 156 18300
rect 44 18232 84 18264
rect 116 18232 156 18264
rect 44 18196 156 18232
rect 44 18164 84 18196
rect 116 18164 156 18196
rect 44 18112 156 18164
rect 44 17870 156 17912
rect 44 17838 84 17870
rect 116 17838 156 17870
rect 44 17802 156 17838
rect 44 17770 84 17802
rect 116 17770 156 17802
rect 44 17734 156 17770
rect 44 17702 84 17734
rect 116 17702 156 17734
rect 44 17666 156 17702
rect 44 17634 84 17666
rect 116 17634 156 17666
rect 44 17598 156 17634
rect 44 17566 84 17598
rect 116 17566 156 17598
rect 44 17530 156 17566
rect 44 17498 84 17530
rect 116 17498 156 17530
rect 44 17462 156 17498
rect 44 17430 84 17462
rect 116 17430 156 17462
rect 44 17394 156 17430
rect 44 17362 84 17394
rect 116 17362 156 17394
rect 44 17326 156 17362
rect 44 17294 84 17326
rect 116 17294 156 17326
rect 44 17258 156 17294
rect 44 17226 84 17258
rect 116 17226 156 17258
rect 44 17190 156 17226
rect 44 17158 84 17190
rect 116 17158 156 17190
rect 44 17122 156 17158
rect 44 17090 84 17122
rect 116 17090 156 17122
rect 44 17054 156 17090
rect 44 17022 84 17054
rect 116 17022 156 17054
rect 44 16986 156 17022
rect 44 16954 84 16986
rect 116 16954 156 16986
rect 44 16918 156 16954
rect 44 16886 84 16918
rect 116 16886 156 16918
rect 44 16850 156 16886
rect 44 16818 84 16850
rect 116 16818 156 16850
rect 44 16782 156 16818
rect 44 16750 84 16782
rect 116 16750 156 16782
rect 44 16714 156 16750
rect 44 16682 84 16714
rect 116 16682 156 16714
rect 44 16646 156 16682
rect 44 16614 84 16646
rect 116 16614 156 16646
rect 44 16578 156 16614
rect 44 16546 84 16578
rect 116 16546 156 16578
rect 44 16510 156 16546
rect 44 16478 84 16510
rect 116 16478 156 16510
rect 44 16442 156 16478
rect 44 16410 84 16442
rect 116 16410 156 16442
rect 44 16374 156 16410
rect 44 16342 84 16374
rect 116 16342 156 16374
rect 44 16306 156 16342
rect 44 16274 84 16306
rect 116 16274 156 16306
rect 44 16238 156 16274
rect 44 16206 84 16238
rect 116 16206 156 16238
rect 44 16170 156 16206
rect 44 16138 84 16170
rect 116 16138 156 16170
rect 44 16102 156 16138
rect 44 16070 84 16102
rect 116 16070 156 16102
rect 44 16034 156 16070
rect 44 16002 84 16034
rect 116 16002 156 16034
rect 44 15966 156 16002
rect 44 15934 84 15966
rect 116 15934 156 15966
rect 44 15898 156 15934
rect 44 15866 84 15898
rect 116 15866 156 15898
rect 44 15830 156 15866
rect 44 15798 84 15830
rect 116 15798 156 15830
rect 44 15762 156 15798
rect 44 15730 84 15762
rect 116 15730 156 15762
rect 44 15694 156 15730
rect 44 15662 84 15694
rect 116 15662 156 15694
rect 44 15626 156 15662
rect 44 15594 84 15626
rect 116 15594 156 15626
rect 44 15558 156 15594
rect 44 15526 84 15558
rect 116 15526 156 15558
rect 44 15490 156 15526
rect 44 15458 84 15490
rect 116 15458 156 15490
rect 44 15422 156 15458
rect 44 15390 84 15422
rect 116 15390 156 15422
rect 44 15354 156 15390
rect 44 15322 84 15354
rect 116 15322 156 15354
rect 44 15286 156 15322
rect 44 15254 84 15286
rect 116 15254 156 15286
rect 44 15218 156 15254
rect 44 15186 84 15218
rect 116 15186 156 15218
rect 44 15150 156 15186
rect 44 15118 84 15150
rect 116 15118 156 15150
rect 44 15082 156 15118
rect 44 15050 84 15082
rect 116 15050 156 15082
rect 44 15014 156 15050
rect 44 14982 84 15014
rect 116 14982 156 15014
rect 44 14946 156 14982
rect 44 14914 84 14946
rect 116 14914 156 14946
rect 44 14878 156 14914
rect 44 14846 84 14878
rect 116 14846 156 14878
rect 44 14810 156 14846
rect 44 14778 84 14810
rect 116 14778 156 14810
rect 44 14742 156 14778
rect 44 14710 84 14742
rect 116 14710 156 14742
rect 44 14674 156 14710
rect 44 14642 84 14674
rect 116 14642 156 14674
rect 44 14606 156 14642
rect 44 14574 84 14606
rect 116 14574 156 14606
rect 44 14538 156 14574
rect 44 14506 84 14538
rect 116 14506 156 14538
rect 44 14470 156 14506
rect 44 14438 84 14470
rect 116 14438 156 14470
rect 44 14402 156 14438
rect 44 14370 84 14402
rect 116 14370 156 14402
rect 44 14334 156 14370
rect 44 14302 84 14334
rect 116 14302 156 14334
rect 44 14266 156 14302
rect 44 14234 84 14266
rect 116 14234 156 14266
rect 44 14198 156 14234
rect 44 14166 84 14198
rect 116 14166 156 14198
rect 44 14130 156 14166
rect 44 14098 84 14130
rect 116 14098 156 14130
rect 44 14062 156 14098
rect 44 14030 84 14062
rect 116 14030 156 14062
rect 44 13994 156 14030
rect 44 13962 84 13994
rect 116 13962 156 13994
rect 44 13926 156 13962
rect 44 13894 84 13926
rect 116 13894 156 13926
rect 44 13858 156 13894
rect 44 13826 84 13858
rect 116 13826 156 13858
rect 44 13790 156 13826
rect 44 13758 84 13790
rect 116 13758 156 13790
rect 44 13722 156 13758
rect 44 13690 84 13722
rect 116 13690 156 13722
rect 44 13654 156 13690
rect 44 13622 84 13654
rect 116 13622 156 13654
rect 44 13586 156 13622
rect 44 13554 84 13586
rect 116 13554 156 13586
rect 44 13518 156 13554
rect 44 13486 84 13518
rect 116 13486 156 13518
rect 44 13450 156 13486
rect 44 13418 84 13450
rect 116 13418 156 13450
rect 44 13382 156 13418
rect 44 13350 84 13382
rect 116 13350 156 13382
rect 44 13314 156 13350
rect 44 13282 84 13314
rect 116 13282 156 13314
rect 44 13246 156 13282
rect 44 13214 84 13246
rect 116 13214 156 13246
rect 44 13178 156 13214
rect 44 13146 84 13178
rect 116 13146 156 13178
rect 44 13110 156 13146
rect 44 13078 84 13110
rect 116 13078 156 13110
rect 44 13000 156 13078
<< nsubdiff >>
rect 44 33416 156 33430
rect 44 33384 84 33416
rect 116 33384 156 33416
rect 44 33370 156 33384
rect 44 29716 156 29730
rect 44 29684 84 29716
rect 116 29684 156 29716
rect 44 29670 156 29684
rect 44 6800 156 12200
rect 44 1200 156 6600
<< psubdiffcont >>
rect 84 31452 116 31484
rect 84 27967 116 27999
rect 84 22856 116 22888
rect 84 17838 116 17870
<< nsubdiffcont >>
rect 84 33384 116 33416
rect 84 29684 116 29716
<< metal1 >>
rect 84 31384 116 31416
rect 84 31316 116 31348
rect 84 31248 116 31280
rect 84 31180 116 31212
rect 84 31112 116 31144
rect 84 27899 116 27931
rect 84 27831 116 27863
rect 84 27763 116 27795
rect 84 27695 116 27727
rect 84 27627 116 27659
rect 84 27559 116 27591
rect 84 27491 116 27523
rect 84 27423 116 27455
rect 84 27355 116 27387
rect 84 27287 116 27319
rect 84 27219 116 27251
rect 84 27151 116 27183
rect 84 27083 116 27115
rect 84 27015 116 27047
rect 84 26947 116 26979
rect 84 26879 116 26911
rect 84 26811 116 26843
rect 84 26743 116 26775
rect 84 26675 116 26707
rect 84 26607 116 26639
rect 84 26539 116 26571
rect 84 26471 116 26503
rect 84 26403 116 26435
rect 84 26335 116 26367
rect 84 26267 116 26299
rect 84 26199 116 26231
rect 84 26131 116 26163
rect 84 26063 116 26095
rect 84 25995 116 26027
rect 84 25927 116 25959
rect 84 25859 116 25891
rect 84 25791 116 25823
rect 84 25723 116 25755
rect 84 25655 116 25687
rect 84 25587 116 25619
rect 84 25519 116 25551
rect 84 25451 116 25483
rect 84 25383 116 25415
rect 84 25315 116 25347
rect 84 25247 116 25279
rect 84 25179 116 25211
rect 84 25111 116 25143
rect 84 25043 116 25075
rect 84 24975 116 25007
rect 84 24907 116 24939
rect 84 24839 116 24871
rect 84 24771 116 24803
rect 84 24703 116 24735
rect 84 24635 116 24667
rect 84 24567 116 24599
rect 84 24499 116 24531
rect 84 24431 116 24463
rect 84 24363 116 24395
rect 84 24295 116 24327
rect 84 24227 116 24259
rect 84 24159 116 24191
rect 84 24091 116 24123
rect 84 24023 116 24055
rect 84 23955 116 23987
rect 84 23887 116 23919
rect 84 23819 116 23851
rect 84 23751 116 23783
rect 84 23683 116 23715
rect 84 23615 116 23647
rect 84 23547 116 23579
rect 84 23479 116 23511
rect 84 23411 116 23443
rect 84 23343 116 23375
rect 84 23275 116 23307
rect 84 23207 116 23239
rect 84 22788 116 22820
rect 84 22720 116 22752
rect 84 22652 116 22684
rect 84 22584 116 22616
rect 84 22516 116 22548
rect 84 22448 116 22480
rect 84 22380 116 22412
rect 84 22312 116 22344
rect 84 22244 116 22276
rect 84 22176 116 22208
rect 84 22108 116 22140
rect 84 22040 116 22072
rect 84 21972 116 22004
rect 84 21904 116 21936
rect 84 21836 116 21868
rect 84 21768 116 21800
rect 84 21700 116 21732
rect 84 21632 116 21664
rect 84 21564 116 21596
rect 84 21496 116 21528
rect 84 21428 116 21460
rect 84 21360 116 21392
rect 84 21292 116 21324
rect 84 21224 116 21256
rect 84 21156 116 21188
rect 84 21088 116 21120
rect 84 21020 116 21052
rect 84 20952 116 20984
rect 84 20884 116 20916
rect 84 20816 116 20848
rect 84 20748 116 20780
rect 84 20680 116 20712
rect 84 20612 116 20644
rect 84 20544 116 20576
rect 84 20476 116 20508
rect 84 20408 116 20440
rect 84 20340 116 20372
rect 84 20272 116 20304
rect 84 20204 116 20236
rect 84 20136 116 20168
rect 84 20068 116 20100
rect 84 20000 116 20032
rect 84 19932 116 19964
rect 84 19864 116 19896
rect 84 19796 116 19828
rect 84 19728 116 19760
rect 84 19660 116 19692
rect 84 19592 116 19624
rect 84 19524 116 19556
rect 84 19456 116 19488
rect 84 19388 116 19420
rect 84 19320 116 19352
rect 84 19252 116 19284
rect 84 19184 116 19216
rect 84 19116 116 19148
rect 84 19048 116 19080
rect 84 18980 116 19012
rect 84 18912 116 18944
rect 84 18844 116 18876
rect 84 18776 116 18808
rect 84 18708 116 18740
rect 84 18640 116 18672
rect 84 18572 116 18604
rect 84 18504 116 18536
rect 84 18436 116 18468
rect 84 18368 116 18400
rect 84 18300 116 18332
rect 84 18232 116 18264
rect 84 18164 116 18196
rect 84 17770 116 17802
rect 84 17702 116 17734
rect 84 17634 116 17666
rect 84 17566 116 17598
rect 84 17498 116 17530
rect 84 17430 116 17462
rect 84 17362 116 17394
rect 84 17294 116 17326
rect 84 17226 116 17258
rect 84 17158 116 17190
rect 84 17090 116 17122
rect 84 17022 116 17054
rect 84 16954 116 16986
rect 84 16886 116 16918
rect 84 16818 116 16850
rect 84 16750 116 16782
rect 84 16682 116 16714
rect 84 16614 116 16646
rect 84 16546 116 16578
rect 84 16478 116 16510
rect 84 16410 116 16442
rect 84 16342 116 16374
rect 84 16274 116 16306
rect 84 16206 116 16238
rect 84 16138 116 16170
rect 84 16070 116 16102
rect 84 16002 116 16034
rect 84 15934 116 15966
rect 84 15866 116 15898
rect 84 15798 116 15830
rect 84 15730 116 15762
rect 84 15662 116 15694
rect 84 15594 116 15626
rect 84 15526 116 15558
rect 84 15458 116 15490
rect 84 15390 116 15422
rect 84 15322 116 15354
rect 84 15254 116 15286
rect 84 15186 116 15218
rect 84 15118 116 15150
rect 84 15050 116 15082
rect 84 14982 116 15014
rect 84 14914 116 14946
rect 84 14846 116 14878
rect 84 14778 116 14810
rect 84 14710 116 14742
rect 84 14642 116 14674
rect 84 14574 116 14606
rect 84 14506 116 14538
rect 84 14438 116 14470
rect 84 14370 116 14402
rect 84 14302 116 14334
rect 84 14234 116 14266
rect 84 14166 116 14198
rect 84 14098 116 14130
rect 84 14030 116 14062
rect 84 13962 116 13994
rect 84 13894 116 13926
rect 84 13826 116 13858
rect 84 13758 116 13790
rect 84 13690 116 13722
rect 84 13622 116 13654
rect 84 13554 116 13586
rect 84 13486 116 13518
rect 84 13418 116 13450
rect 84 13350 116 13382
rect 84 13282 116 13314
rect 84 13214 116 13246
rect 84 13146 116 13178
rect 84 13078 116 13110
rect 0 33384 84 33416
rect 116 33384 200 33416
rect 84 31484 116 31500
rect 84 31416 116 31452
rect 0 31384 84 31416
rect 116 31384 200 31416
rect 84 31348 116 31384
rect 84 31280 116 31316
rect 84 31212 116 31248
rect 84 31144 116 31180
rect 84 31090 116 31112
rect 0 29684 84 29716
rect 116 29684 200 29716
rect 0 27999 200 28034
rect 0 27967 84 27999
rect 116 27967 200 27999
rect 0 27931 200 27967
rect 0 27899 84 27931
rect 116 27899 200 27931
rect 0 27863 200 27899
rect 0 27831 84 27863
rect 116 27831 200 27863
rect 0 27795 200 27831
rect 0 27763 84 27795
rect 116 27763 200 27795
rect 0 27727 200 27763
rect 0 27695 84 27727
rect 116 27695 200 27727
rect 0 27659 200 27695
rect 0 27627 84 27659
rect 116 27627 200 27659
rect 0 27591 200 27627
rect 0 27559 84 27591
rect 116 27559 200 27591
rect 0 27523 200 27559
rect 0 27491 84 27523
rect 116 27491 200 27523
rect 0 27455 200 27491
rect 0 27423 84 27455
rect 116 27423 200 27455
rect 0 27387 200 27423
rect 0 27355 84 27387
rect 116 27355 200 27387
rect 0 27319 200 27355
rect 0 27287 84 27319
rect 116 27287 200 27319
rect 0 27251 200 27287
rect 0 27219 84 27251
rect 116 27219 200 27251
rect 0 27183 200 27219
rect 0 27151 84 27183
rect 116 27151 200 27183
rect 0 27115 200 27151
rect 0 27083 84 27115
rect 116 27083 200 27115
rect 0 27047 200 27083
rect 0 27015 84 27047
rect 116 27015 200 27047
rect 0 26979 200 27015
rect 0 26947 84 26979
rect 116 26947 200 26979
rect 0 26911 200 26947
rect 0 26879 84 26911
rect 116 26879 200 26911
rect 0 26843 200 26879
rect 0 26811 84 26843
rect 116 26811 200 26843
rect 0 26775 200 26811
rect 0 26743 84 26775
rect 116 26743 200 26775
rect 0 26707 200 26743
rect 0 26675 84 26707
rect 116 26675 200 26707
rect 0 26639 200 26675
rect 0 26607 84 26639
rect 116 26607 200 26639
rect 0 26571 200 26607
rect 0 26539 84 26571
rect 116 26539 200 26571
rect 0 26503 200 26539
rect 0 26471 84 26503
rect 116 26471 200 26503
rect 0 26435 200 26471
rect 0 26403 84 26435
rect 116 26403 200 26435
rect 0 26367 200 26403
rect 0 26335 84 26367
rect 116 26335 200 26367
rect 0 26299 200 26335
rect 0 26267 84 26299
rect 116 26267 200 26299
rect 0 26231 200 26267
rect 0 26199 84 26231
rect 116 26199 200 26231
rect 0 26163 200 26199
rect 0 26131 84 26163
rect 116 26131 200 26163
rect 0 26095 200 26131
rect 0 26063 84 26095
rect 116 26063 200 26095
rect 0 26027 200 26063
rect 0 25995 84 26027
rect 116 25995 200 26027
rect 0 25959 200 25995
rect 0 25927 84 25959
rect 116 25927 200 25959
rect 0 25891 200 25927
rect 0 25859 84 25891
rect 116 25859 200 25891
rect 0 25823 200 25859
rect 0 25791 84 25823
rect 116 25791 200 25823
rect 0 25755 200 25791
rect 0 25723 84 25755
rect 116 25723 200 25755
rect 0 25687 200 25723
rect 0 25655 84 25687
rect 116 25655 200 25687
rect 0 25619 200 25655
rect 0 25587 84 25619
rect 116 25587 200 25619
rect 0 25551 200 25587
rect 0 25519 84 25551
rect 116 25519 200 25551
rect 0 25483 200 25519
rect 0 25451 84 25483
rect 116 25451 200 25483
rect 0 25415 200 25451
rect 0 25383 84 25415
rect 116 25383 200 25415
rect 0 25347 200 25383
rect 0 25315 84 25347
rect 116 25315 200 25347
rect 0 25279 200 25315
rect 0 25247 84 25279
rect 116 25247 200 25279
rect 0 25211 200 25247
rect 0 25179 84 25211
rect 116 25179 200 25211
rect 0 25143 200 25179
rect 0 25111 84 25143
rect 116 25111 200 25143
rect 0 25075 200 25111
rect 0 25043 84 25075
rect 116 25043 200 25075
rect 0 25007 200 25043
rect 0 24975 84 25007
rect 116 24975 200 25007
rect 0 24939 200 24975
rect 0 24907 84 24939
rect 116 24907 200 24939
rect 0 24871 200 24907
rect 0 24839 84 24871
rect 116 24839 200 24871
rect 0 24803 200 24839
rect 0 24771 84 24803
rect 116 24771 200 24803
rect 0 24735 200 24771
rect 0 24703 84 24735
rect 116 24703 200 24735
rect 0 24667 200 24703
rect 0 24635 84 24667
rect 116 24635 200 24667
rect 0 24599 200 24635
rect 0 24567 84 24599
rect 116 24567 200 24599
rect 0 24531 200 24567
rect 0 24499 84 24531
rect 116 24499 200 24531
rect 0 24463 200 24499
rect 0 24431 84 24463
rect 116 24431 200 24463
rect 0 24395 200 24431
rect 0 24363 84 24395
rect 116 24363 200 24395
rect 0 24327 200 24363
rect 0 24295 84 24327
rect 116 24295 200 24327
rect 0 24259 200 24295
rect 0 24227 84 24259
rect 116 24227 200 24259
rect 0 24191 200 24227
rect 0 24159 84 24191
rect 116 24159 200 24191
rect 0 24123 200 24159
rect 0 24091 84 24123
rect 116 24091 200 24123
rect 0 24055 200 24091
rect 0 24023 84 24055
rect 116 24023 200 24055
rect 0 23987 200 24023
rect 0 23955 84 23987
rect 116 23955 200 23987
rect 0 23919 200 23955
rect 0 23887 84 23919
rect 116 23887 200 23919
rect 0 23851 200 23887
rect 0 23819 84 23851
rect 116 23819 200 23851
rect 0 23783 200 23819
rect 0 23751 84 23783
rect 116 23751 200 23783
rect 0 23715 200 23751
rect 0 23683 84 23715
rect 116 23683 200 23715
rect 0 23647 200 23683
rect 0 23615 84 23647
rect 116 23615 200 23647
rect 0 23579 200 23615
rect 0 23547 84 23579
rect 116 23547 200 23579
rect 0 23511 200 23547
rect 0 23479 84 23511
rect 116 23479 200 23511
rect 0 23443 200 23479
rect 0 23411 84 23443
rect 116 23411 200 23443
rect 0 23375 200 23411
rect 0 23343 84 23375
rect 116 23343 200 23375
rect 0 23307 200 23343
rect 0 23275 84 23307
rect 116 23275 200 23307
rect 0 23239 200 23275
rect 0 23207 84 23239
rect 116 23207 200 23239
rect 0 23124 200 23207
rect 0 22888 200 22924
rect 0 22856 84 22888
rect 116 22856 200 22888
rect 0 22820 200 22856
rect 0 22788 84 22820
rect 116 22788 200 22820
rect 0 22752 200 22788
rect 0 22720 84 22752
rect 116 22720 200 22752
rect 0 22684 200 22720
rect 0 22652 84 22684
rect 116 22652 200 22684
rect 0 22616 200 22652
rect 0 22584 84 22616
rect 116 22584 200 22616
rect 0 22548 200 22584
rect 0 22516 84 22548
rect 116 22516 200 22548
rect 0 22480 200 22516
rect 0 22448 84 22480
rect 116 22448 200 22480
rect 0 22412 200 22448
rect 0 22380 84 22412
rect 116 22380 200 22412
rect 0 22344 200 22380
rect 0 22312 84 22344
rect 116 22312 200 22344
rect 0 22276 200 22312
rect 0 22244 84 22276
rect 116 22244 200 22276
rect 0 22208 200 22244
rect 0 22176 84 22208
rect 116 22176 200 22208
rect 0 22140 200 22176
rect 0 22108 84 22140
rect 116 22108 200 22140
rect 0 22072 200 22108
rect 0 22040 84 22072
rect 116 22040 200 22072
rect 0 22004 200 22040
rect 0 21972 84 22004
rect 116 21972 200 22004
rect 0 21936 200 21972
rect 0 21904 84 21936
rect 116 21904 200 21936
rect 0 21868 200 21904
rect 0 21836 84 21868
rect 116 21836 200 21868
rect 0 21800 200 21836
rect 0 21768 84 21800
rect 116 21768 200 21800
rect 0 21732 200 21768
rect 0 21700 84 21732
rect 116 21700 200 21732
rect 0 21664 200 21700
rect 0 21632 84 21664
rect 116 21632 200 21664
rect 0 21596 200 21632
rect 0 21564 84 21596
rect 116 21564 200 21596
rect 0 21528 200 21564
rect 0 21496 84 21528
rect 116 21496 200 21528
rect 0 21460 200 21496
rect 0 21428 84 21460
rect 116 21428 200 21460
rect 0 21392 200 21428
rect 0 21360 84 21392
rect 116 21360 200 21392
rect 0 21324 200 21360
rect 0 21292 84 21324
rect 116 21292 200 21324
rect 0 21256 200 21292
rect 0 21224 84 21256
rect 116 21224 200 21256
rect 0 21188 200 21224
rect 0 21156 84 21188
rect 116 21156 200 21188
rect 0 21120 200 21156
rect 0 21088 84 21120
rect 116 21088 200 21120
rect 0 21052 200 21088
rect 0 21020 84 21052
rect 116 21020 200 21052
rect 0 20984 200 21020
rect 0 20952 84 20984
rect 116 20952 200 20984
rect 0 20916 200 20952
rect 0 20884 84 20916
rect 116 20884 200 20916
rect 0 20848 200 20884
rect 0 20816 84 20848
rect 116 20816 200 20848
rect 0 20780 200 20816
rect 0 20748 84 20780
rect 116 20748 200 20780
rect 0 20712 200 20748
rect 0 20680 84 20712
rect 116 20680 200 20712
rect 0 20644 200 20680
rect 0 20612 84 20644
rect 116 20612 200 20644
rect 0 20576 200 20612
rect 0 20544 84 20576
rect 116 20544 200 20576
rect 0 20508 200 20544
rect 0 20476 84 20508
rect 116 20476 200 20508
rect 0 20440 200 20476
rect 0 20408 84 20440
rect 116 20408 200 20440
rect 0 20372 200 20408
rect 0 20340 84 20372
rect 116 20340 200 20372
rect 0 20304 200 20340
rect 0 20272 84 20304
rect 116 20272 200 20304
rect 0 20236 200 20272
rect 0 20204 84 20236
rect 116 20204 200 20236
rect 0 20168 200 20204
rect 0 20136 84 20168
rect 116 20136 200 20168
rect 0 20100 200 20136
rect 0 20068 84 20100
rect 116 20068 200 20100
rect 0 20032 200 20068
rect 0 20000 84 20032
rect 116 20000 200 20032
rect 0 19964 200 20000
rect 0 19932 84 19964
rect 116 19932 200 19964
rect 0 19896 200 19932
rect 0 19864 84 19896
rect 116 19864 200 19896
rect 0 19828 200 19864
rect 0 19796 84 19828
rect 116 19796 200 19828
rect 0 19760 200 19796
rect 0 19728 84 19760
rect 116 19728 200 19760
rect 0 19692 200 19728
rect 0 19660 84 19692
rect 116 19660 200 19692
rect 0 19624 200 19660
rect 0 19592 84 19624
rect 116 19592 200 19624
rect 0 19556 200 19592
rect 0 19524 84 19556
rect 116 19524 200 19556
rect 0 19488 200 19524
rect 0 19456 84 19488
rect 116 19456 200 19488
rect 0 19420 200 19456
rect 0 19388 84 19420
rect 116 19388 200 19420
rect 0 19352 200 19388
rect 0 19320 84 19352
rect 116 19320 200 19352
rect 0 19284 200 19320
rect 0 19252 84 19284
rect 116 19252 200 19284
rect 0 19216 200 19252
rect 0 19184 84 19216
rect 116 19184 200 19216
rect 0 19148 200 19184
rect 0 19116 84 19148
rect 116 19116 200 19148
rect 0 19080 200 19116
rect 0 19048 84 19080
rect 116 19048 200 19080
rect 0 19012 200 19048
rect 0 18980 84 19012
rect 116 18980 200 19012
rect 0 18944 200 18980
rect 0 18912 84 18944
rect 116 18912 200 18944
rect 0 18876 200 18912
rect 0 18844 84 18876
rect 116 18844 200 18876
rect 0 18808 200 18844
rect 0 18776 84 18808
rect 116 18776 200 18808
rect 0 18740 200 18776
rect 0 18708 84 18740
rect 116 18708 200 18740
rect 0 18672 200 18708
rect 0 18640 84 18672
rect 116 18640 200 18672
rect 0 18604 200 18640
rect 0 18572 84 18604
rect 116 18572 200 18604
rect 0 18536 200 18572
rect 0 18504 84 18536
rect 116 18504 200 18536
rect 0 18468 200 18504
rect 0 18436 84 18468
rect 116 18436 200 18468
rect 0 18400 200 18436
rect 0 18368 84 18400
rect 116 18368 200 18400
rect 0 18332 200 18368
rect 0 18300 84 18332
rect 116 18300 200 18332
rect 0 18264 200 18300
rect 0 18232 84 18264
rect 116 18232 200 18264
rect 0 18196 200 18232
rect 0 18164 84 18196
rect 116 18164 200 18196
rect 0 18112 200 18164
rect 0 17870 200 17912
rect 0 17838 84 17870
rect 116 17838 200 17870
rect 0 17802 200 17838
rect 0 17770 84 17802
rect 116 17770 200 17802
rect 0 17734 200 17770
rect 0 17702 84 17734
rect 116 17702 200 17734
rect 0 17666 200 17702
rect 0 17634 84 17666
rect 116 17634 200 17666
rect 0 17598 200 17634
rect 0 17566 84 17598
rect 116 17566 200 17598
rect 0 17530 200 17566
rect 0 17498 84 17530
rect 116 17498 200 17530
rect 0 17462 200 17498
rect 0 17430 84 17462
rect 116 17430 200 17462
rect 0 17394 200 17430
rect 0 17362 84 17394
rect 116 17362 200 17394
rect 0 17326 200 17362
rect 0 17294 84 17326
rect 116 17294 200 17326
rect 0 17258 200 17294
rect 0 17226 84 17258
rect 116 17226 200 17258
rect 0 17190 200 17226
rect 0 17158 84 17190
rect 116 17158 200 17190
rect 0 17122 200 17158
rect 0 17090 84 17122
rect 116 17090 200 17122
rect 0 17054 200 17090
rect 0 17022 84 17054
rect 116 17022 200 17054
rect 0 16986 200 17022
rect 0 16954 84 16986
rect 116 16954 200 16986
rect 0 16918 200 16954
rect 0 16886 84 16918
rect 116 16886 200 16918
rect 0 16850 200 16886
rect 0 16818 84 16850
rect 116 16818 200 16850
rect 0 16782 200 16818
rect 0 16750 84 16782
rect 116 16750 200 16782
rect 0 16714 200 16750
rect 0 16682 84 16714
rect 116 16682 200 16714
rect 0 16646 200 16682
rect 0 16614 84 16646
rect 116 16614 200 16646
rect 0 16578 200 16614
rect 0 16546 84 16578
rect 116 16546 200 16578
rect 0 16510 200 16546
rect 0 16478 84 16510
rect 116 16478 200 16510
rect 0 16442 200 16478
rect 0 16410 84 16442
rect 116 16410 200 16442
rect 0 16374 200 16410
rect 0 16342 84 16374
rect 116 16342 200 16374
rect 0 16306 200 16342
rect 0 16274 84 16306
rect 116 16274 200 16306
rect 0 16238 200 16274
rect 0 16206 84 16238
rect 116 16206 200 16238
rect 0 16170 200 16206
rect 0 16138 84 16170
rect 116 16138 200 16170
rect 0 16102 200 16138
rect 0 16070 84 16102
rect 116 16070 200 16102
rect 0 16034 200 16070
rect 0 16002 84 16034
rect 116 16002 200 16034
rect 0 15966 200 16002
rect 0 15934 84 15966
rect 116 15934 200 15966
rect 0 15898 200 15934
rect 0 15866 84 15898
rect 116 15866 200 15898
rect 0 15830 200 15866
rect 0 15798 84 15830
rect 116 15798 200 15830
rect 0 15762 200 15798
rect 0 15730 84 15762
rect 116 15730 200 15762
rect 0 15694 200 15730
rect 0 15662 84 15694
rect 116 15662 200 15694
rect 0 15626 200 15662
rect 0 15594 84 15626
rect 116 15594 200 15626
rect 0 15558 200 15594
rect 0 15526 84 15558
rect 116 15526 200 15558
rect 0 15490 200 15526
rect 0 15458 84 15490
rect 116 15458 200 15490
rect 0 15422 200 15458
rect 0 15390 84 15422
rect 116 15390 200 15422
rect 0 15354 200 15390
rect 0 15322 84 15354
rect 116 15322 200 15354
rect 0 15286 200 15322
rect 0 15254 84 15286
rect 116 15254 200 15286
rect 0 15218 200 15254
rect 0 15186 84 15218
rect 116 15186 200 15218
rect 0 15150 200 15186
rect 0 15118 84 15150
rect 116 15118 200 15150
rect 0 15082 200 15118
rect 0 15050 84 15082
rect 116 15050 200 15082
rect 0 15014 200 15050
rect 0 14982 84 15014
rect 116 14982 200 15014
rect 0 14946 200 14982
rect 0 14914 84 14946
rect 116 14914 200 14946
rect 0 14878 200 14914
rect 0 14846 84 14878
rect 116 14846 200 14878
rect 0 14810 200 14846
rect 0 14778 84 14810
rect 116 14778 200 14810
rect 0 14742 200 14778
rect 0 14710 84 14742
rect 116 14710 200 14742
rect 0 14674 200 14710
rect 0 14642 84 14674
rect 116 14642 200 14674
rect 0 14606 200 14642
rect 0 14574 84 14606
rect 116 14574 200 14606
rect 0 14538 200 14574
rect 0 14506 84 14538
rect 116 14506 200 14538
rect 0 14470 200 14506
rect 0 14438 84 14470
rect 116 14438 200 14470
rect 0 14402 200 14438
rect 0 14370 84 14402
rect 116 14370 200 14402
rect 0 14334 200 14370
rect 0 14302 84 14334
rect 116 14302 200 14334
rect 0 14266 200 14302
rect 0 14234 84 14266
rect 116 14234 200 14266
rect 0 14198 200 14234
rect 0 14166 84 14198
rect 116 14166 200 14198
rect 0 14130 200 14166
rect 0 14098 84 14130
rect 116 14098 200 14130
rect 0 14062 200 14098
rect 0 14030 84 14062
rect 116 14030 200 14062
rect 0 13994 200 14030
rect 0 13962 84 13994
rect 116 13962 200 13994
rect 0 13926 200 13962
rect 0 13894 84 13926
rect 116 13894 200 13926
rect 0 13858 200 13894
rect 0 13826 84 13858
rect 116 13826 200 13858
rect 0 13790 200 13826
rect 0 13758 84 13790
rect 116 13758 200 13790
rect 0 13722 200 13758
rect 0 13690 84 13722
rect 116 13690 200 13722
rect 0 13654 200 13690
rect 0 13622 84 13654
rect 116 13622 200 13654
rect 0 13586 200 13622
rect 0 13554 84 13586
rect 116 13554 200 13586
rect 0 13518 200 13554
rect 0 13486 84 13518
rect 116 13486 200 13518
rect 0 13450 200 13486
rect 0 13418 84 13450
rect 116 13418 200 13450
rect 0 13382 200 13418
rect 0 13350 84 13382
rect 116 13350 200 13382
rect 0 13314 200 13350
rect 0 13282 84 13314
rect 116 13282 200 13314
rect 0 13246 200 13282
rect 0 13214 84 13246
rect 116 13214 200 13246
rect 0 13178 200 13214
rect 0 13146 84 13178
rect 116 13146 200 13178
rect 0 13110 200 13146
rect 0 13078 84 13110
rect 116 13078 200 13110
rect 0 13000 200 13078
rect 0 6800 200 12200
rect 0 1200 200 6600
<< metal3 >>
rect 0 32000 200 35600
rect 0 28000 200 31600
rect 0 25200 200 26800
rect 0 18700 200 23800
rect 0 13200 200 18300
rect 0 6900 200 12000
rect 0 1400 200 6500
<< metal4 >>
rect 0 32440 200 35600
rect 0 28000 200 31160
rect 0 25200 200 26800
rect 0 18700 200 23800
rect 0 13200 200 18300
rect 0 6900 200 12000
rect 0 1400 200 6500
<< metal5 >>
rect 0 32000 200 35600
rect 0 28000 200 31600
rect 0 25200 200 26800
rect 0 18700 200 23800
rect 0 13200 200 18300
rect 0 6900 200 12000
rect 0 1400 200 6500
<< metal6 >>
rect -68 32000 268 35600
rect -68 28000 268 31600
rect -68 25200 268 26800
rect -68 18700 268 23800
rect -68 13200 268 18300
rect -68 6900 268 12000
rect -68 1400 268 6500
<< metal7 >>
rect -100 25500 300 26500
rect -100 19000 300 23500
rect -100 13500 300 18000
rect -100 7200 300 11700
rect -100 1700 300 6200
<< labels >>
rlabel metal3 s 0 32000 200 35600 4 vdd
port 2 nsew
rlabel metal3 s 0 28000 200 31600 4 vss
port 1 nsew
rlabel metal3 s 0 18700 200 23800 4 iovdd
port 4 nsew
rlabel metal3 s 0 13200 200 18300 4 iovdd
port 4 nsew
rlabel metal3 s 0 6900 200 12000 4 iovss
port 3 nsew
rlabel metal3 s 0 25200 200 26800 4 iovss
port 3 nsew
rlabel metal3 s 0 1400 200 6500 4 iovss
port 3 nsew
rlabel metal4 s 0 28000 200 31160 4 vdd
port 2 nsew
rlabel metal4 s 0 32440 200 35600 4 vss
port 1 nsew
rlabel metal4 s 0 18700 200 23800 4 iovdd
port 4 nsew
rlabel metal4 s 0 13200 200 18300 4 iovdd
port 4 nsew
rlabel metal4 s 0 6900 200 12000 4 iovss
port 3 nsew
rlabel metal4 s 0 25200 200 26800 4 iovss
port 3 nsew
rlabel metal4 s 0 1400 200 6500 4 iovss
port 3 nsew
rlabel metal5 s 0 28000 200 31600 4 vdd
port 2 nsew
rlabel metal5 s 0 32000 200 35600 4 vss
port 1 nsew
rlabel metal5 s 0 18700 200 23800 4 iovdd
port 4 nsew
rlabel metal5 s 0 13200 200 18300 4 iovdd
port 4 nsew
rlabel metal5 s 0 6900 200 12000 4 iovss
port 3 nsew
rlabel metal5 s 0 25200 200 26800 4 iovss
port 3 nsew
rlabel metal5 s 0 1400 200 6500 4 iovss
port 3 nsew
rlabel metal6 s 0 28000 200 31600 4 vdd
port 2 nsew
rlabel metal6 s 0 32000 200 35600 4 vss
port 1 nsew
rlabel metal6 s 0 18700 200 23800 4 iovdd
port 4 nsew
rlabel metal6 s 0 13200 200 18300 4 iovdd
port 4 nsew
rlabel metal6 s 0 6900 200 12000 4 iovss
port 3 nsew
rlabel metal6 s 0 25200 200 26800 4 iovss
port 3 nsew
rlabel metal6 s 0 1400 200 6500 4 iovss
port 3 nsew
rlabel metal7 s 0 13500 200 18000 4 iovdd
port 4 nsew
rlabel metal7 s 0 19000 200 23500 4 iovdd
port 4 nsew
rlabel metal7 s 0 7200 200 11700 4 iovss
port 3 nsew
rlabel metal7 s 0 25500 200 26500 4 iovss
port 3 nsew
rlabel metal7 s 0 1700 200 6200 4 iovss
port 3 nsew
flabel comment s 97 13068 97 13068 0 FreeSans 400 0 0 0 sub!
flabel comment s 97 18219 97 18219 0 FreeSans 400 0 0 0 sub!
flabel comment s 97 23261 97 23261 0 FreeSans 400 0 0 0 sub!
flabel comment s 105 31405 105 31405 0 FreeSans 400 0 0 0 sub!
flabel metal1 s 74 13128 136 13164 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 74 18270 136 18306 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 74 23148 136 23184 0 FreeSans 400 0 0 0 iovss
port 3 nsew
flabel metal1 s 78 31392 139 31409 0 FreeSans 400 0 0 0 vss
port 1 nsew
<< properties >>
string device primitive
string FIXED_BBOX 0 0 200 36000
string GDS_END 63482776
string GDS_FILE sg13g2_io.gds
string GDS_START 63459466
<< end >>
