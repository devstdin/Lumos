magic
tech ihp-sg13g2
timestamp 1757240632
<< error_p >>
rect -33 80 -28 85
rect 28 80 33 85
rect 136 80 141 85
rect 197 80 202 85
rect 305 80 310 85
rect 366 80 371 85
rect 474 80 479 85
rect 535 80 540 85
rect 643 80 648 85
rect 704 80 709 85
rect 812 80 817 85
rect 873 80 878 85
rect 981 80 986 85
rect 1042 80 1047 85
rect 1150 80 1155 85
rect 1211 80 1216 85
rect 1319 80 1324 85
rect 1380 80 1385 85
rect 1488 80 1493 85
rect 1549 80 1554 85
rect 1657 80 1662 85
rect 1718 80 1723 85
rect 1826 80 1831 85
rect 1887 80 1892 85
rect 1995 80 2000 85
rect 2056 80 2061 85
rect 2164 80 2169 85
rect 2225 80 2230 85
rect 2333 80 2338 85
rect 2394 80 2399 85
rect 2502 80 2507 85
rect 2563 80 2568 85
rect 2671 80 2676 85
rect 2732 80 2737 85
rect 2840 80 2845 85
rect 2901 80 2906 85
rect 3009 80 3014 85
rect 3070 80 3075 85
rect 3178 80 3183 85
rect 3239 80 3244 85
rect 3347 80 3352 85
rect 3408 80 3413 85
rect 3516 80 3521 85
rect 3577 80 3582 85
rect -38 75 -33 80
rect 33 75 38 80
rect 131 75 136 80
rect 202 75 207 80
rect 300 75 305 80
rect 371 75 376 80
rect 469 75 474 80
rect 540 75 545 80
rect 638 75 643 80
rect 709 75 714 80
rect 807 75 812 80
rect 878 75 883 80
rect 976 75 981 80
rect 1047 75 1052 80
rect 1145 75 1150 80
rect 1216 75 1221 80
rect 1314 75 1319 80
rect 1385 75 1390 80
rect 1483 75 1488 80
rect 1554 75 1559 80
rect 1652 75 1657 80
rect 1723 75 1728 80
rect 1821 75 1826 80
rect 1892 75 1897 80
rect 1990 75 1995 80
rect 2061 75 2066 80
rect 2159 75 2164 80
rect 2230 75 2235 80
rect 2328 75 2333 80
rect 2399 75 2404 80
rect 2497 75 2502 80
rect 2568 75 2573 80
rect 2666 75 2671 80
rect 2737 75 2742 80
rect 2835 75 2840 80
rect 2906 75 2911 80
rect 3004 75 3009 80
rect 3075 75 3080 80
rect 3173 75 3178 80
rect 3244 75 3249 80
rect 3342 75 3347 80
rect 3413 75 3418 80
rect 3511 75 3516 80
rect 3582 75 3587 80
rect -38 64 -33 69
rect 33 64 38 69
rect 131 64 136 69
rect 202 64 207 69
rect 300 64 305 69
rect 371 64 376 69
rect 469 64 474 69
rect 540 64 545 69
rect 638 64 643 69
rect 709 64 714 69
rect 807 64 812 69
rect 878 64 883 69
rect 976 64 981 69
rect 1047 64 1052 69
rect 1145 64 1150 69
rect 1216 64 1221 69
rect 1314 64 1319 69
rect 1385 64 1390 69
rect 1483 64 1488 69
rect 1554 64 1559 69
rect 1652 64 1657 69
rect 1723 64 1728 69
rect 1821 64 1826 69
rect 1892 64 1897 69
rect 1990 64 1995 69
rect 2061 64 2066 69
rect 2159 64 2164 69
rect 2230 64 2235 69
rect 2328 64 2333 69
rect 2399 64 2404 69
rect 2497 64 2502 69
rect 2568 64 2573 69
rect 2666 64 2671 69
rect 2737 64 2742 69
rect 2835 64 2840 69
rect 2906 64 2911 69
rect 3004 64 3009 69
rect 3075 64 3080 69
rect 3173 64 3178 69
rect 3244 64 3249 69
rect 3342 64 3347 69
rect 3413 64 3418 69
rect 3511 64 3516 69
rect 3582 64 3587 69
rect -33 59 -28 64
rect 28 59 33 64
rect 136 59 141 64
rect 197 59 202 64
rect 305 59 310 64
rect 366 59 371 64
rect 474 59 479 64
rect 535 59 540 64
rect 643 59 648 64
rect 704 59 709 64
rect 812 59 817 64
rect 873 59 878 64
rect 981 59 986 64
rect 1042 59 1047 64
rect 1150 59 1155 64
rect 1211 59 1216 64
rect 1319 59 1324 64
rect 1380 59 1385 64
rect 1488 59 1493 64
rect 1549 59 1554 64
rect 1657 59 1662 64
rect 1718 59 1723 64
rect 1826 59 1831 64
rect 1887 59 1892 64
rect 1995 59 2000 64
rect 2056 59 2061 64
rect 2164 59 2169 64
rect 2225 59 2230 64
rect 2333 59 2338 64
rect 2394 59 2399 64
rect 2502 59 2507 64
rect 2563 59 2568 64
rect 2671 59 2676 64
rect 2732 59 2737 64
rect 2840 59 2845 64
rect 2901 59 2906 64
rect 3009 59 3014 64
rect 3070 59 3075 64
rect 3178 59 3183 64
rect 3239 59 3244 64
rect 3347 59 3352 64
rect 3408 59 3413 64
rect 3516 59 3521 64
rect 3577 59 3582 64
rect -67 43 -62 48
rect -56 43 -51 48
rect 51 43 56 48
rect 62 43 67 48
rect 102 43 107 48
rect 113 43 118 48
rect 220 43 225 48
rect 231 43 236 48
rect 271 43 276 48
rect 282 43 287 48
rect 389 43 394 48
rect 400 43 405 48
rect 440 43 445 48
rect 451 43 456 48
rect 558 43 563 48
rect 569 43 574 48
rect 609 43 614 48
rect 620 43 625 48
rect 727 43 732 48
rect 738 43 743 48
rect 778 43 783 48
rect 789 43 794 48
rect 896 43 901 48
rect 907 43 912 48
rect 947 43 952 48
rect 958 43 963 48
rect 1065 43 1070 48
rect 1076 43 1081 48
rect 1116 43 1121 48
rect 1127 43 1132 48
rect 1234 43 1239 48
rect 1245 43 1250 48
rect 1285 43 1290 48
rect 1296 43 1301 48
rect 1403 43 1408 48
rect 1414 43 1419 48
rect 1454 43 1459 48
rect 1465 43 1470 48
rect 1572 43 1577 48
rect 1583 43 1588 48
rect 1623 43 1628 48
rect 1634 43 1639 48
rect 1741 43 1746 48
rect 1752 43 1757 48
rect 1792 43 1797 48
rect 1803 43 1808 48
rect 1910 43 1915 48
rect 1921 43 1926 48
rect 1961 43 1966 48
rect 1972 43 1977 48
rect 2079 43 2084 48
rect 2090 43 2095 48
rect 2130 43 2135 48
rect 2141 43 2146 48
rect 2248 43 2253 48
rect 2259 43 2264 48
rect 2299 43 2304 48
rect 2310 43 2315 48
rect 2417 43 2422 48
rect 2428 43 2433 48
rect 2468 43 2473 48
rect 2479 43 2484 48
rect 2586 43 2591 48
rect 2597 43 2602 48
rect 2637 43 2642 48
rect 2648 43 2653 48
rect 2755 43 2760 48
rect 2766 43 2771 48
rect 2806 43 2811 48
rect 2817 43 2822 48
rect 2924 43 2929 48
rect 2935 43 2940 48
rect 2975 43 2980 48
rect 2986 43 2991 48
rect 3093 43 3098 48
rect 3104 43 3109 48
rect 3144 43 3149 48
rect 3155 43 3160 48
rect 3262 43 3267 48
rect 3273 43 3278 48
rect 3313 43 3318 48
rect 3324 43 3329 48
rect 3431 43 3436 48
rect 3442 43 3447 48
rect 3482 43 3487 48
rect 3493 43 3498 48
rect 3600 43 3605 48
rect 3611 43 3616 48
rect -72 38 -67 43
rect -51 38 -46 43
rect 46 38 51 43
rect 67 38 72 43
rect 97 38 102 43
rect 118 38 123 43
rect 215 38 220 43
rect 236 38 241 43
rect 266 38 271 43
rect 287 38 292 43
rect 384 38 389 43
rect 405 38 410 43
rect 435 38 440 43
rect 456 38 461 43
rect 553 38 558 43
rect 574 38 579 43
rect 604 38 609 43
rect 625 38 630 43
rect 722 38 727 43
rect 743 38 748 43
rect 773 38 778 43
rect 794 38 799 43
rect 891 38 896 43
rect 912 38 917 43
rect 942 38 947 43
rect 963 38 968 43
rect 1060 38 1065 43
rect 1081 38 1086 43
rect 1111 38 1116 43
rect 1132 38 1137 43
rect 1229 38 1234 43
rect 1250 38 1255 43
rect 1280 38 1285 43
rect 1301 38 1306 43
rect 1398 38 1403 43
rect 1419 38 1424 43
rect 1449 38 1454 43
rect 1470 38 1475 43
rect 1567 38 1572 43
rect 1588 38 1593 43
rect 1618 38 1623 43
rect 1639 38 1644 43
rect 1736 38 1741 43
rect 1757 38 1762 43
rect 1787 38 1792 43
rect 1808 38 1813 43
rect 1905 38 1910 43
rect 1926 38 1931 43
rect 1956 38 1961 43
rect 1977 38 1982 43
rect 2074 38 2079 43
rect 2095 38 2100 43
rect 2125 38 2130 43
rect 2146 38 2151 43
rect 2243 38 2248 43
rect 2264 38 2269 43
rect 2294 38 2299 43
rect 2315 38 2320 43
rect 2412 38 2417 43
rect 2433 38 2438 43
rect 2463 38 2468 43
rect 2484 38 2489 43
rect 2581 38 2586 43
rect 2602 38 2607 43
rect 2632 38 2637 43
rect 2653 38 2658 43
rect 2750 38 2755 43
rect 2771 38 2776 43
rect 2801 38 2806 43
rect 2822 38 2827 43
rect 2919 38 2924 43
rect 2940 38 2945 43
rect 2970 38 2975 43
rect 2991 38 2996 43
rect 3088 38 3093 43
rect 3109 38 3114 43
rect 3139 38 3144 43
rect 3160 38 3165 43
rect 3257 38 3262 43
rect 3278 38 3283 43
rect 3308 38 3313 43
rect 3329 38 3334 43
rect 3426 38 3431 43
rect 3447 38 3452 43
rect 3477 38 3482 43
rect 3498 38 3503 43
rect 3595 38 3600 43
rect 3616 38 3621 43
rect -72 -43 -67 -38
rect -51 -43 -46 -38
rect 46 -43 51 -38
rect 67 -43 72 -38
rect 97 -43 102 -38
rect 118 -43 123 -38
rect 215 -43 220 -38
rect 236 -43 241 -38
rect 266 -43 271 -38
rect 287 -43 292 -38
rect 384 -43 389 -38
rect 405 -43 410 -38
rect 435 -43 440 -38
rect 456 -43 461 -38
rect 553 -43 558 -38
rect 574 -43 579 -38
rect 604 -43 609 -38
rect 625 -43 630 -38
rect 722 -43 727 -38
rect 743 -43 748 -38
rect 773 -43 778 -38
rect 794 -43 799 -38
rect 891 -43 896 -38
rect 912 -43 917 -38
rect 942 -43 947 -38
rect 963 -43 968 -38
rect 1060 -43 1065 -38
rect 1081 -43 1086 -38
rect 1111 -43 1116 -38
rect 1132 -43 1137 -38
rect 1229 -43 1234 -38
rect 1250 -43 1255 -38
rect 1280 -43 1285 -38
rect 1301 -43 1306 -38
rect 1398 -43 1403 -38
rect 1419 -43 1424 -38
rect 1449 -43 1454 -38
rect 1470 -43 1475 -38
rect 1567 -43 1572 -38
rect 1588 -43 1593 -38
rect 1618 -43 1623 -38
rect 1639 -43 1644 -38
rect 1736 -43 1741 -38
rect 1757 -43 1762 -38
rect 1787 -43 1792 -38
rect 1808 -43 1813 -38
rect 1905 -43 1910 -38
rect 1926 -43 1931 -38
rect 1956 -43 1961 -38
rect 1977 -43 1982 -38
rect 2074 -43 2079 -38
rect 2095 -43 2100 -38
rect 2125 -43 2130 -38
rect 2146 -43 2151 -38
rect 2243 -43 2248 -38
rect 2264 -43 2269 -38
rect 2294 -43 2299 -38
rect 2315 -43 2320 -38
rect 2412 -43 2417 -38
rect 2433 -43 2438 -38
rect 2463 -43 2468 -38
rect 2484 -43 2489 -38
rect 2581 -43 2586 -38
rect 2602 -43 2607 -38
rect 2632 -43 2637 -38
rect 2653 -43 2658 -38
rect 2750 -43 2755 -38
rect 2771 -43 2776 -38
rect 2801 -43 2806 -38
rect 2822 -43 2827 -38
rect 2919 -43 2924 -38
rect 2940 -43 2945 -38
rect 2970 -43 2975 -38
rect 2991 -43 2996 -38
rect 3088 -43 3093 -38
rect 3109 -43 3114 -38
rect 3139 -43 3144 -38
rect 3160 -43 3165 -38
rect 3257 -43 3262 -38
rect 3278 -43 3283 -38
rect 3308 -43 3313 -38
rect 3329 -43 3334 -38
rect 3426 -43 3431 -38
rect 3447 -43 3452 -38
rect 3477 -43 3482 -38
rect 3498 -43 3503 -38
rect 3595 -43 3600 -38
rect 3616 -43 3621 -38
rect -67 -48 -62 -43
rect -56 -48 -51 -43
rect 51 -48 56 -43
rect 62 -48 67 -43
rect 102 -48 107 -43
rect 113 -48 118 -43
rect 220 -48 225 -43
rect 231 -48 236 -43
rect 271 -48 276 -43
rect 282 -48 287 -43
rect 389 -48 394 -43
rect 400 -48 405 -43
rect 440 -48 445 -43
rect 451 -48 456 -43
rect 558 -48 563 -43
rect 569 -48 574 -43
rect 609 -48 614 -43
rect 620 -48 625 -43
rect 727 -48 732 -43
rect 738 -48 743 -43
rect 778 -48 783 -43
rect 789 -48 794 -43
rect 896 -48 901 -43
rect 907 -48 912 -43
rect 947 -48 952 -43
rect 958 -48 963 -43
rect 1065 -48 1070 -43
rect 1076 -48 1081 -43
rect 1116 -48 1121 -43
rect 1127 -48 1132 -43
rect 1234 -48 1239 -43
rect 1245 -48 1250 -43
rect 1285 -48 1290 -43
rect 1296 -48 1301 -43
rect 1403 -48 1408 -43
rect 1414 -48 1419 -43
rect 1454 -48 1459 -43
rect 1465 -48 1470 -43
rect 1572 -48 1577 -43
rect 1583 -48 1588 -43
rect 1623 -48 1628 -43
rect 1634 -48 1639 -43
rect 1741 -48 1746 -43
rect 1752 -48 1757 -43
rect 1792 -48 1797 -43
rect 1803 -48 1808 -43
rect 1910 -48 1915 -43
rect 1921 -48 1926 -43
rect 1961 -48 1966 -43
rect 1972 -48 1977 -43
rect 2079 -48 2084 -43
rect 2090 -48 2095 -43
rect 2130 -48 2135 -43
rect 2141 -48 2146 -43
rect 2248 -48 2253 -43
rect 2259 -48 2264 -43
rect 2299 -48 2304 -43
rect 2310 -48 2315 -43
rect 2417 -48 2422 -43
rect 2428 -48 2433 -43
rect 2468 -48 2473 -43
rect 2479 -48 2484 -43
rect 2586 -48 2591 -43
rect 2597 -48 2602 -43
rect 2637 -48 2642 -43
rect 2648 -48 2653 -43
rect 2755 -48 2760 -43
rect 2766 -48 2771 -43
rect 2806 -48 2811 -43
rect 2817 -48 2822 -43
rect 2924 -48 2929 -43
rect 2935 -48 2940 -43
rect 2975 -48 2980 -43
rect 2986 -48 2991 -43
rect 3093 -48 3098 -43
rect 3104 -48 3109 -43
rect 3144 -48 3149 -43
rect 3155 -48 3160 -43
rect 3262 -48 3267 -43
rect 3273 -48 3278 -43
rect 3313 -48 3318 -43
rect 3324 -48 3329 -43
rect 3431 -48 3436 -43
rect 3442 -48 3447 -43
rect 3482 -48 3487 -43
rect 3493 -48 3498 -43
rect 3600 -48 3605 -43
rect 3611 -48 3616 -43
rect -33 -64 -28 -59
rect 28 -64 33 -59
rect 136 -64 141 -59
rect 197 -64 202 -59
rect 305 -64 310 -59
rect 366 -64 371 -59
rect 474 -64 479 -59
rect 535 -64 540 -59
rect 643 -64 648 -59
rect 704 -64 709 -59
rect 812 -64 817 -59
rect 873 -64 878 -59
rect 981 -64 986 -59
rect 1042 -64 1047 -59
rect 1150 -64 1155 -59
rect 1211 -64 1216 -59
rect 1319 -64 1324 -59
rect 1380 -64 1385 -59
rect 1488 -64 1493 -59
rect 1549 -64 1554 -59
rect 1657 -64 1662 -59
rect 1718 -64 1723 -59
rect 1826 -64 1831 -59
rect 1887 -64 1892 -59
rect 1995 -64 2000 -59
rect 2056 -64 2061 -59
rect 2164 -64 2169 -59
rect 2225 -64 2230 -59
rect 2333 -64 2338 -59
rect 2394 -64 2399 -59
rect 2502 -64 2507 -59
rect 2563 -64 2568 -59
rect 2671 -64 2676 -59
rect 2732 -64 2737 -59
rect 2840 -64 2845 -59
rect 2901 -64 2906 -59
rect 3009 -64 3014 -59
rect 3070 -64 3075 -59
rect 3178 -64 3183 -59
rect 3239 -64 3244 -59
rect 3347 -64 3352 -59
rect 3408 -64 3413 -59
rect 3516 -64 3521 -59
rect 3577 -64 3582 -59
rect -38 -69 -33 -64
rect 33 -69 38 -64
rect 131 -69 136 -64
rect 202 -69 207 -64
rect 300 -69 305 -64
rect 371 -69 376 -64
rect 469 -69 474 -64
rect 540 -69 545 -64
rect 638 -69 643 -64
rect 709 -69 714 -64
rect 807 -69 812 -64
rect 878 -69 883 -64
rect 976 -69 981 -64
rect 1047 -69 1052 -64
rect 1145 -69 1150 -64
rect 1216 -69 1221 -64
rect 1314 -69 1319 -64
rect 1385 -69 1390 -64
rect 1483 -69 1488 -64
rect 1554 -69 1559 -64
rect 1652 -69 1657 -64
rect 1723 -69 1728 -64
rect 1821 -69 1826 -64
rect 1892 -69 1897 -64
rect 1990 -69 1995 -64
rect 2061 -69 2066 -64
rect 2159 -69 2164 -64
rect 2230 -69 2235 -64
rect 2328 -69 2333 -64
rect 2399 -69 2404 -64
rect 2497 -69 2502 -64
rect 2568 -69 2573 -64
rect 2666 -69 2671 -64
rect 2737 -69 2742 -64
rect 2835 -69 2840 -64
rect 2906 -69 2911 -64
rect 3004 -69 3009 -64
rect 3075 -69 3080 -64
rect 3173 -69 3178 -64
rect 3244 -69 3249 -64
rect 3342 -69 3347 -64
rect 3413 -69 3418 -64
rect 3511 -69 3516 -64
rect 3582 -69 3587 -64
rect -38 -80 -33 -75
rect 33 -80 38 -75
rect 131 -80 136 -75
rect 202 -80 207 -75
rect 300 -80 305 -75
rect 371 -80 376 -75
rect 469 -80 474 -75
rect 540 -80 545 -75
rect 638 -80 643 -75
rect 709 -80 714 -75
rect 807 -80 812 -75
rect 878 -80 883 -75
rect 976 -80 981 -75
rect 1047 -80 1052 -75
rect 1145 -80 1150 -75
rect 1216 -80 1221 -75
rect 1314 -80 1319 -75
rect 1385 -80 1390 -75
rect 1483 -80 1488 -75
rect 1554 -80 1559 -75
rect 1652 -80 1657 -75
rect 1723 -80 1728 -75
rect 1821 -80 1826 -75
rect 1892 -80 1897 -75
rect 1990 -80 1995 -75
rect 2061 -80 2066 -75
rect 2159 -80 2164 -75
rect 2230 -80 2235 -75
rect 2328 -80 2333 -75
rect 2399 -80 2404 -75
rect 2497 -80 2502 -75
rect 2568 -80 2573 -75
rect 2666 -80 2671 -75
rect 2737 -80 2742 -75
rect 2835 -80 2840 -75
rect 2906 -80 2911 -75
rect 3004 -80 3009 -75
rect 3075 -80 3080 -75
rect 3173 -80 3178 -75
rect 3244 -80 3249 -75
rect 3342 -80 3347 -75
rect 3413 -80 3418 -75
rect 3511 -80 3516 -75
rect 3582 -80 3587 -75
rect -33 -85 -28 -80
rect 28 -85 33 -80
rect 136 -85 141 -80
rect 197 -85 202 -80
rect 305 -85 310 -80
rect 366 -85 371 -80
rect 474 -85 479 -80
rect 535 -85 540 -80
rect 643 -85 648 -80
rect 704 -85 709 -80
rect 812 -85 817 -80
rect 873 -85 878 -80
rect 981 -85 986 -80
rect 1042 -85 1047 -80
rect 1150 -85 1155 -80
rect 1211 -85 1216 -80
rect 1319 -85 1324 -80
rect 1380 -85 1385 -80
rect 1488 -85 1493 -80
rect 1549 -85 1554 -80
rect 1657 -85 1662 -80
rect 1718 -85 1723 -80
rect 1826 -85 1831 -80
rect 1887 -85 1892 -80
rect 1995 -85 2000 -80
rect 2056 -85 2061 -80
rect 2164 -85 2169 -80
rect 2225 -85 2230 -80
rect 2333 -85 2338 -80
rect 2394 -85 2399 -80
rect 2502 -85 2507 -80
rect 2563 -85 2568 -80
rect 2671 -85 2676 -80
rect 2732 -85 2737 -80
rect 2840 -85 2845 -80
rect 2901 -85 2906 -80
rect 3009 -85 3014 -80
rect 3070 -85 3075 -80
rect 3178 -85 3183 -80
rect 3239 -85 3244 -80
rect 3347 -85 3352 -80
rect 3408 -85 3413 -80
rect 3516 -85 3521 -80
rect 3577 -85 3582 -80
<< nwell >>
rect -247 -87 3796 212
rect -136 -112 3685 -87
<< hvpmos >>
rect -40 -50 40 50
rect 129 -50 209 50
rect 298 -50 378 50
rect 467 -50 547 50
rect 636 -50 716 50
rect 805 -50 885 50
rect 974 -50 1054 50
rect 1143 -50 1223 50
rect 1312 -50 1392 50
rect 1481 -50 1561 50
rect 1650 -50 1730 50
rect 1819 -50 1899 50
rect 1988 -50 2068 50
rect 2157 -50 2237 50
rect 2326 -50 2406 50
rect 2495 -50 2575 50
rect 2664 -50 2744 50
rect 2833 -50 2913 50
rect 3002 -50 3082 50
rect 3171 -50 3251 50
rect 3340 -50 3420 50
rect 3509 -50 3589 50
<< hvpdiff >>
rect -74 43 -40 50
rect -74 -43 -67 43
rect -51 -43 -40 43
rect -74 -50 -40 -43
rect 40 43 74 50
rect 40 -43 51 43
rect 67 -43 74 43
rect 40 -50 74 -43
rect 95 43 129 50
rect 95 -43 102 43
rect 118 -43 129 43
rect 95 -50 129 -43
rect 209 43 243 50
rect 209 -43 220 43
rect 236 -43 243 43
rect 209 -50 243 -43
rect 264 43 298 50
rect 264 -43 271 43
rect 287 -43 298 43
rect 264 -50 298 -43
rect 378 43 412 50
rect 378 -43 389 43
rect 405 -43 412 43
rect 378 -50 412 -43
rect 433 43 467 50
rect 433 -43 440 43
rect 456 -43 467 43
rect 433 -50 467 -43
rect 547 43 581 50
rect 547 -43 558 43
rect 574 -43 581 43
rect 547 -50 581 -43
rect 602 43 636 50
rect 602 -43 609 43
rect 625 -43 636 43
rect 602 -50 636 -43
rect 716 43 750 50
rect 716 -43 727 43
rect 743 -43 750 43
rect 716 -50 750 -43
rect 771 43 805 50
rect 771 -43 778 43
rect 794 -43 805 43
rect 771 -50 805 -43
rect 885 43 919 50
rect 885 -43 896 43
rect 912 -43 919 43
rect 885 -50 919 -43
rect 940 43 974 50
rect 940 -43 947 43
rect 963 -43 974 43
rect 940 -50 974 -43
rect 1054 43 1088 50
rect 1054 -43 1065 43
rect 1081 -43 1088 43
rect 1054 -50 1088 -43
rect 1109 43 1143 50
rect 1109 -43 1116 43
rect 1132 -43 1143 43
rect 1109 -50 1143 -43
rect 1223 43 1257 50
rect 1223 -43 1234 43
rect 1250 -43 1257 43
rect 1223 -50 1257 -43
rect 1278 43 1312 50
rect 1278 -43 1285 43
rect 1301 -43 1312 43
rect 1278 -50 1312 -43
rect 1392 43 1426 50
rect 1392 -43 1403 43
rect 1419 -43 1426 43
rect 1392 -50 1426 -43
rect 1447 43 1481 50
rect 1447 -43 1454 43
rect 1470 -43 1481 43
rect 1447 -50 1481 -43
rect 1561 43 1595 50
rect 1561 -43 1572 43
rect 1588 -43 1595 43
rect 1561 -50 1595 -43
rect 1616 43 1650 50
rect 1616 -43 1623 43
rect 1639 -43 1650 43
rect 1616 -50 1650 -43
rect 1730 43 1764 50
rect 1730 -43 1741 43
rect 1757 -43 1764 43
rect 1730 -50 1764 -43
rect 1785 43 1819 50
rect 1785 -43 1792 43
rect 1808 -43 1819 43
rect 1785 -50 1819 -43
rect 1899 43 1933 50
rect 1899 -43 1910 43
rect 1926 -43 1933 43
rect 1899 -50 1933 -43
rect 1954 43 1988 50
rect 1954 -43 1961 43
rect 1977 -43 1988 43
rect 1954 -50 1988 -43
rect 2068 43 2102 50
rect 2068 -43 2079 43
rect 2095 -43 2102 43
rect 2068 -50 2102 -43
rect 2123 43 2157 50
rect 2123 -43 2130 43
rect 2146 -43 2157 43
rect 2123 -50 2157 -43
rect 2237 43 2271 50
rect 2237 -43 2248 43
rect 2264 -43 2271 43
rect 2237 -50 2271 -43
rect 2292 43 2326 50
rect 2292 -43 2299 43
rect 2315 -43 2326 43
rect 2292 -50 2326 -43
rect 2406 43 2440 50
rect 2406 -43 2417 43
rect 2433 -43 2440 43
rect 2406 -50 2440 -43
rect 2461 43 2495 50
rect 2461 -43 2468 43
rect 2484 -43 2495 43
rect 2461 -50 2495 -43
rect 2575 43 2609 50
rect 2575 -43 2586 43
rect 2602 -43 2609 43
rect 2575 -50 2609 -43
rect 2630 43 2664 50
rect 2630 -43 2637 43
rect 2653 -43 2664 43
rect 2630 -50 2664 -43
rect 2744 43 2778 50
rect 2744 -43 2755 43
rect 2771 -43 2778 43
rect 2744 -50 2778 -43
rect 2799 43 2833 50
rect 2799 -43 2806 43
rect 2822 -43 2833 43
rect 2799 -50 2833 -43
rect 2913 43 2947 50
rect 2913 -43 2924 43
rect 2940 -43 2947 43
rect 2913 -50 2947 -43
rect 2968 43 3002 50
rect 2968 -43 2975 43
rect 2991 -43 3002 43
rect 2968 -50 3002 -43
rect 3082 43 3116 50
rect 3082 -43 3093 43
rect 3109 -43 3116 43
rect 3082 -50 3116 -43
rect 3137 43 3171 50
rect 3137 -43 3144 43
rect 3160 -43 3171 43
rect 3137 -50 3171 -43
rect 3251 43 3285 50
rect 3251 -43 3262 43
rect 3278 -43 3285 43
rect 3251 -50 3285 -43
rect 3306 43 3340 50
rect 3306 -43 3313 43
rect 3329 -43 3340 43
rect 3306 -50 3340 -43
rect 3420 43 3454 50
rect 3420 -43 3431 43
rect 3447 -43 3454 43
rect 3420 -50 3454 -43
rect 3475 43 3509 50
rect 3475 -43 3482 43
rect 3498 -43 3509 43
rect 3475 -50 3509 -43
rect 3589 43 3623 50
rect 3589 -43 3600 43
rect 3616 -43 3623 43
rect 3589 -50 3623 -43
<< hvpdiffc >>
rect -67 -43 -51 43
rect 51 -43 67 43
rect 102 -43 118 43
rect 220 -43 236 43
rect 271 -43 287 43
rect 389 -43 405 43
rect 440 -43 456 43
rect 558 -43 574 43
rect 609 -43 625 43
rect 727 -43 743 43
rect 778 -43 794 43
rect 896 -43 912 43
rect 947 -43 963 43
rect 1065 -43 1081 43
rect 1116 -43 1132 43
rect 1234 -43 1250 43
rect 1285 -43 1301 43
rect 1403 -43 1419 43
rect 1454 -43 1470 43
rect 1572 -43 1588 43
rect 1623 -43 1639 43
rect 1741 -43 1757 43
rect 1792 -43 1808 43
rect 1910 -43 1926 43
rect 1961 -43 1977 43
rect 2079 -43 2095 43
rect 2130 -43 2146 43
rect 2248 -43 2264 43
rect 2299 -43 2315 43
rect 2417 -43 2433 43
rect 2468 -43 2484 43
rect 2586 -43 2602 43
rect 2637 -43 2653 43
rect 2755 -43 2771 43
rect 2806 -43 2822 43
rect 2924 -43 2940 43
rect 2975 -43 2991 43
rect 3093 -43 3109 43
rect 3144 -43 3160 43
rect 3262 -43 3278 43
rect 3313 -43 3329 43
rect 3431 -43 3447 43
rect 3482 -43 3498 43
rect 3600 -43 3616 43
<< nsubdiff >>
rect -185 143 3734 150
rect -185 127 -148 143
rect 3697 127 3734 143
rect -185 120 3734 127
rect -185 113 -155 120
rect -185 -18 -178 113
rect -162 -18 -155 113
rect 3704 113 3734 120
rect -185 -25 -155 -18
rect 3704 -18 3711 113
rect 3727 -18 3734 113
rect 3704 -25 3734 -18
<< nsubdiffcont >>
rect -148 127 3697 143
rect -178 -18 -162 113
rect 3711 -18 3727 113
<< poly >>
rect -40 80 40 87
rect -40 64 -33 80
rect 33 64 40 80
rect -40 50 40 64
rect 129 80 209 87
rect 129 64 136 80
rect 202 64 209 80
rect 129 50 209 64
rect 298 80 378 87
rect 298 64 305 80
rect 371 64 378 80
rect 298 50 378 64
rect 467 80 547 87
rect 467 64 474 80
rect 540 64 547 80
rect 467 50 547 64
rect 636 80 716 87
rect 636 64 643 80
rect 709 64 716 80
rect 636 50 716 64
rect 805 80 885 87
rect 805 64 812 80
rect 878 64 885 80
rect 805 50 885 64
rect 974 80 1054 87
rect 974 64 981 80
rect 1047 64 1054 80
rect 974 50 1054 64
rect 1143 80 1223 87
rect 1143 64 1150 80
rect 1216 64 1223 80
rect 1143 50 1223 64
rect 1312 80 1392 87
rect 1312 64 1319 80
rect 1385 64 1392 80
rect 1312 50 1392 64
rect 1481 80 1561 87
rect 1481 64 1488 80
rect 1554 64 1561 80
rect 1481 50 1561 64
rect 1650 80 1730 87
rect 1650 64 1657 80
rect 1723 64 1730 80
rect 1650 50 1730 64
rect 1819 80 1899 87
rect 1819 64 1826 80
rect 1892 64 1899 80
rect 1819 50 1899 64
rect 1988 80 2068 87
rect 1988 64 1995 80
rect 2061 64 2068 80
rect 1988 50 2068 64
rect 2157 80 2237 87
rect 2157 64 2164 80
rect 2230 64 2237 80
rect 2157 50 2237 64
rect 2326 80 2406 87
rect 2326 64 2333 80
rect 2399 64 2406 80
rect 2326 50 2406 64
rect 2495 80 2575 87
rect 2495 64 2502 80
rect 2568 64 2575 80
rect 2495 50 2575 64
rect 2664 80 2744 87
rect 2664 64 2671 80
rect 2737 64 2744 80
rect 2664 50 2744 64
rect 2833 80 2913 87
rect 2833 64 2840 80
rect 2906 64 2913 80
rect 2833 50 2913 64
rect 3002 80 3082 87
rect 3002 64 3009 80
rect 3075 64 3082 80
rect 3002 50 3082 64
rect 3171 80 3251 87
rect 3171 64 3178 80
rect 3244 64 3251 80
rect 3171 50 3251 64
rect 3340 80 3420 87
rect 3340 64 3347 80
rect 3413 64 3420 80
rect 3340 50 3420 64
rect 3509 80 3589 87
rect 3509 64 3516 80
rect 3582 64 3589 80
rect 3509 50 3589 64
rect -40 -64 40 -50
rect -40 -80 -33 -64
rect 33 -80 40 -64
rect -40 -87 40 -80
rect 129 -64 209 -50
rect 129 -80 136 -64
rect 202 -80 209 -64
rect 129 -87 209 -80
rect 298 -64 378 -50
rect 298 -80 305 -64
rect 371 -80 378 -64
rect 298 -87 378 -80
rect 467 -64 547 -50
rect 467 -80 474 -64
rect 540 -80 547 -64
rect 467 -87 547 -80
rect 636 -64 716 -50
rect 636 -80 643 -64
rect 709 -80 716 -64
rect 636 -87 716 -80
rect 805 -64 885 -50
rect 805 -80 812 -64
rect 878 -80 885 -64
rect 805 -87 885 -80
rect 974 -64 1054 -50
rect 974 -80 981 -64
rect 1047 -80 1054 -64
rect 974 -87 1054 -80
rect 1143 -64 1223 -50
rect 1143 -80 1150 -64
rect 1216 -80 1223 -64
rect 1143 -87 1223 -80
rect 1312 -64 1392 -50
rect 1312 -80 1319 -64
rect 1385 -80 1392 -64
rect 1312 -87 1392 -80
rect 1481 -64 1561 -50
rect 1481 -80 1488 -64
rect 1554 -80 1561 -64
rect 1481 -87 1561 -80
rect 1650 -64 1730 -50
rect 1650 -80 1657 -64
rect 1723 -80 1730 -64
rect 1650 -87 1730 -80
rect 1819 -64 1899 -50
rect 1819 -80 1826 -64
rect 1892 -80 1899 -64
rect 1819 -87 1899 -80
rect 1988 -64 2068 -50
rect 1988 -80 1995 -64
rect 2061 -80 2068 -64
rect 1988 -87 2068 -80
rect 2157 -64 2237 -50
rect 2157 -80 2164 -64
rect 2230 -80 2237 -64
rect 2157 -87 2237 -80
rect 2326 -64 2406 -50
rect 2326 -80 2333 -64
rect 2399 -80 2406 -64
rect 2326 -87 2406 -80
rect 2495 -64 2575 -50
rect 2495 -80 2502 -64
rect 2568 -80 2575 -64
rect 2495 -87 2575 -80
rect 2664 -64 2744 -50
rect 2664 -80 2671 -64
rect 2737 -80 2744 -64
rect 2664 -87 2744 -80
rect 2833 -64 2913 -50
rect 2833 -80 2840 -64
rect 2906 -80 2913 -64
rect 2833 -87 2913 -80
rect 3002 -64 3082 -50
rect 3002 -80 3009 -64
rect 3075 -80 3082 -64
rect 3002 -87 3082 -80
rect 3171 -64 3251 -50
rect 3171 -80 3178 -64
rect 3244 -80 3251 -64
rect 3171 -87 3251 -80
rect 3340 -64 3420 -50
rect 3340 -80 3347 -64
rect 3413 -80 3420 -64
rect 3340 -87 3420 -80
rect 3509 -64 3589 -50
rect 3509 -80 3516 -64
rect 3582 -80 3589 -64
rect 3509 -87 3589 -80
<< polycont >>
rect -33 64 33 80
rect 136 64 202 80
rect 305 64 371 80
rect 474 64 540 80
rect 643 64 709 80
rect 812 64 878 80
rect 981 64 1047 80
rect 1150 64 1216 80
rect 1319 64 1385 80
rect 1488 64 1554 80
rect 1657 64 1723 80
rect 1826 64 1892 80
rect 1995 64 2061 80
rect 2164 64 2230 80
rect 2333 64 2399 80
rect 2502 64 2568 80
rect 2671 64 2737 80
rect 2840 64 2906 80
rect 3009 64 3075 80
rect 3178 64 3244 80
rect 3347 64 3413 80
rect 3516 64 3582 80
rect -33 -80 33 -64
rect 136 -80 202 -64
rect 305 -80 371 -64
rect 474 -80 540 -64
rect 643 -80 709 -64
rect 812 -80 878 -64
rect 981 -80 1047 -64
rect 1150 -80 1216 -64
rect 1319 -80 1385 -64
rect 1488 -80 1554 -64
rect 1657 -80 1723 -64
rect 1826 -80 1892 -64
rect 1995 -80 2061 -64
rect 2164 -80 2230 -64
rect 2333 -80 2399 -64
rect 2502 -80 2568 -64
rect 2671 -80 2737 -64
rect 2840 -80 2906 -64
rect 3009 -80 3075 -64
rect 3178 -80 3244 -64
rect 3347 -80 3413 -64
rect 3516 -80 3582 -64
<< metal1 >>
rect -183 143 3732 148
rect -183 127 -148 143
rect 3697 127 3732 143
rect -183 122 3732 127
rect -183 113 -157 122
rect -183 -18 -178 113
rect -162 -18 -157 113
rect 3706 113 3732 122
rect -183 -23 -157 -18
rect 3706 -18 3711 113
rect 3727 -18 3732 113
rect 3706 -23 3732 -18
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 1 l 0.8 nf 1 nx 22 dx 0.21 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 0
<< end >>
