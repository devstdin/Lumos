magic
tech ihp-sg13g2
timestamp 1748514137
<< error_p >>
rect -93 280 -88 285
rect 88 280 93 285
rect 235 280 240 285
rect 416 280 421 285
rect 563 280 568 285
rect 744 280 749 285
rect 891 280 896 285
rect 1072 280 1077 285
rect 1219 280 1224 285
rect 1400 280 1405 285
rect 1547 280 1552 285
rect 1728 280 1733 285
rect -98 275 -93 280
rect 93 275 98 280
rect 230 275 235 280
rect 421 275 426 280
rect 558 275 563 280
rect 749 275 754 280
rect 886 275 891 280
rect 1077 275 1082 280
rect 1214 275 1219 280
rect 1405 275 1410 280
rect 1542 275 1547 280
rect 1733 275 1738 280
rect -98 264 -93 269
rect 93 264 98 269
rect 230 264 235 269
rect 421 264 426 269
rect 558 264 563 269
rect 749 264 754 269
rect 886 264 891 269
rect 1077 264 1082 269
rect 1214 264 1219 269
rect 1405 264 1410 269
rect 1542 264 1547 269
rect 1733 264 1738 269
rect -93 259 -88 264
rect 88 259 93 264
rect 235 259 240 264
rect 416 259 421 264
rect 563 259 568 264
rect 744 259 749 264
rect 891 259 896 264
rect 1072 259 1077 264
rect 1219 259 1224 264
rect 1400 259 1405 264
rect 1547 259 1552 264
rect 1728 259 1733 264
rect -127 243 -122 248
rect -116 243 -111 248
rect 111 243 116 248
rect 122 243 127 248
rect 201 243 206 248
rect 212 243 217 248
rect 439 243 444 248
rect 450 243 455 248
rect 529 243 534 248
rect 540 243 545 248
rect 767 243 772 248
rect 778 243 783 248
rect 857 243 862 248
rect 868 243 873 248
rect 1095 243 1100 248
rect 1106 243 1111 248
rect 1185 243 1190 248
rect 1196 243 1201 248
rect 1423 243 1428 248
rect 1434 243 1439 248
rect 1513 243 1518 248
rect 1524 243 1529 248
rect 1751 243 1756 248
rect 1762 243 1767 248
rect -132 238 -127 243
rect -111 238 -106 243
rect 106 238 111 243
rect 127 238 132 243
rect 196 238 201 243
rect 217 238 222 243
rect 434 238 439 243
rect 455 238 460 243
rect 524 238 529 243
rect 545 238 550 243
rect 762 238 767 243
rect 783 238 788 243
rect 852 238 857 243
rect 873 238 878 243
rect 1090 238 1095 243
rect 1111 238 1116 243
rect 1180 238 1185 243
rect 1201 238 1206 243
rect 1418 238 1423 243
rect 1439 238 1444 243
rect 1508 238 1513 243
rect 1529 238 1534 243
rect 1746 238 1751 243
rect 1767 238 1772 243
rect -132 -243 -127 -238
rect -111 -243 -106 -238
rect 106 -243 111 -238
rect 127 -243 132 -238
rect 196 -243 201 -238
rect 217 -243 222 -238
rect 434 -243 439 -238
rect 455 -243 460 -238
rect 524 -243 529 -238
rect 545 -243 550 -238
rect 762 -243 767 -238
rect 783 -243 788 -238
rect 852 -243 857 -238
rect 873 -243 878 -238
rect 1090 -243 1095 -238
rect 1111 -243 1116 -238
rect 1180 -243 1185 -238
rect 1201 -243 1206 -238
rect 1418 -243 1423 -238
rect 1439 -243 1444 -238
rect 1508 -243 1513 -238
rect 1529 -243 1534 -238
rect 1746 -243 1751 -238
rect 1767 -243 1772 -238
rect -127 -248 -122 -243
rect -116 -248 -111 -243
rect 111 -248 116 -243
rect 122 -248 127 -243
rect 201 -248 206 -243
rect 212 -248 217 -243
rect 439 -248 444 -243
rect 450 -248 455 -243
rect 529 -248 534 -243
rect 540 -248 545 -243
rect 767 -248 772 -243
rect 778 -248 783 -243
rect 857 -248 862 -243
rect 868 -248 873 -243
rect 1095 -248 1100 -243
rect 1106 -248 1111 -243
rect 1185 -248 1190 -243
rect 1196 -248 1201 -243
rect 1423 -248 1428 -243
rect 1434 -248 1439 -243
rect 1513 -248 1518 -243
rect 1524 -248 1529 -243
rect 1751 -248 1756 -243
rect 1762 -248 1767 -243
rect -93 -264 -88 -259
rect 88 -264 93 -259
rect 235 -264 240 -259
rect 416 -264 421 -259
rect 563 -264 568 -259
rect 744 -264 749 -259
rect 891 -264 896 -259
rect 1072 -264 1077 -259
rect 1219 -264 1224 -259
rect 1400 -264 1405 -259
rect 1547 -264 1552 -259
rect 1728 -264 1733 -259
rect -98 -269 -93 -264
rect 93 -269 98 -264
rect 230 -269 235 -264
rect 421 -269 426 -264
rect 558 -269 563 -264
rect 749 -269 754 -264
rect 886 -269 891 -264
rect 1077 -269 1082 -264
rect 1214 -269 1219 -264
rect 1405 -269 1410 -264
rect 1542 -269 1547 -264
rect 1733 -269 1738 -264
rect -98 -280 -93 -275
rect 93 -280 98 -275
rect 230 -280 235 -275
rect 421 -280 426 -275
rect 558 -280 563 -275
rect 749 -280 754 -275
rect 886 -280 891 -275
rect 1077 -280 1082 -275
rect 1214 -280 1219 -275
rect 1405 -280 1410 -275
rect 1542 -280 1547 -275
rect 1733 -280 1738 -275
rect -93 -285 -88 -280
rect 88 -285 93 -280
rect 235 -285 240 -280
rect 416 -285 421 -280
rect 563 -285 568 -280
rect 744 -285 749 -280
rect 891 -285 896 -280
rect 1072 -285 1077 -280
rect 1219 -285 1224 -280
rect 1400 -285 1405 -280
rect 1547 -285 1552 -280
rect 1728 -285 1733 -280
<< nwell >>
rect -280 -401 1920 401
<< hvpmos >>
rect -100 -250 100 250
rect 228 -250 428 250
rect 556 -250 756 250
rect 884 -250 1084 250
rect 1212 -250 1412 250
rect 1540 -250 1740 250
<< hvpdiff >>
rect -134 243 -100 250
rect -134 -243 -127 243
rect -111 -243 -100 243
rect -134 -250 -100 -243
rect 100 243 134 250
rect 100 -243 111 243
rect 127 -243 134 243
rect 100 -250 134 -243
rect 194 243 228 250
rect 194 -243 201 243
rect 217 -243 228 243
rect 194 -250 228 -243
rect 428 243 462 250
rect 428 -243 439 243
rect 455 -243 462 243
rect 428 -250 462 -243
rect 522 243 556 250
rect 522 -243 529 243
rect 545 -243 556 243
rect 522 -250 556 -243
rect 756 243 790 250
rect 756 -243 767 243
rect 783 -243 790 243
rect 756 -250 790 -243
rect 850 243 884 250
rect 850 -243 857 243
rect 873 -243 884 243
rect 850 -250 884 -243
rect 1084 243 1118 250
rect 1084 -243 1095 243
rect 1111 -243 1118 243
rect 1084 -250 1118 -243
rect 1178 243 1212 250
rect 1178 -243 1185 243
rect 1201 -243 1212 243
rect 1178 -250 1212 -243
rect 1412 243 1446 250
rect 1412 -243 1423 243
rect 1439 -243 1446 243
rect 1412 -250 1446 -243
rect 1506 243 1540 250
rect 1506 -243 1513 243
rect 1529 -243 1540 243
rect 1506 -250 1540 -243
rect 1740 243 1774 250
rect 1740 -243 1751 243
rect 1767 -243 1774 243
rect 1740 -250 1774 -243
<< hvpdiffc >>
rect -127 -243 -111 243
rect 111 -243 127 243
rect 201 -243 217 243
rect 439 -243 455 243
rect 529 -243 545 243
rect 767 -243 783 243
rect 857 -243 873 243
rect 1095 -243 1111 243
rect 1185 -243 1201 243
rect 1423 -243 1439 243
rect 1513 -243 1529 243
rect 1751 -243 1767 243
<< nsubdiff >>
rect -218 332 1858 339
rect -218 316 -181 332
rect 1821 316 1858 332
rect -218 309 1858 316
rect -218 302 -188 309
rect -218 -302 -211 302
rect -195 -302 -188 302
rect 1828 302 1858 309
rect -218 -309 -188 -302
rect 1828 -302 1835 302
rect 1851 -302 1858 302
rect 1828 -309 1858 -302
rect -218 -316 1858 -309
rect -218 -332 -181 -316
rect 1821 -332 1858 -316
rect -218 -339 1858 -332
<< nsubdiffcont >>
rect -181 316 1821 332
rect -211 -302 -195 302
rect 1835 -302 1851 302
rect -181 -332 1821 -316
<< poly >>
rect -100 280 100 287
rect -100 264 -93 280
rect 93 264 100 280
rect -100 250 100 264
rect 228 280 428 287
rect 228 264 235 280
rect 421 264 428 280
rect 228 250 428 264
rect 556 280 756 287
rect 556 264 563 280
rect 749 264 756 280
rect 556 250 756 264
rect 884 280 1084 287
rect 884 264 891 280
rect 1077 264 1084 280
rect 884 250 1084 264
rect 1212 280 1412 287
rect 1212 264 1219 280
rect 1405 264 1412 280
rect 1212 250 1412 264
rect 1540 280 1740 287
rect 1540 264 1547 280
rect 1733 264 1740 280
rect 1540 250 1740 264
rect -100 -264 100 -250
rect -100 -280 -93 -264
rect 93 -280 100 -264
rect -100 -287 100 -280
rect 228 -264 428 -250
rect 228 -280 235 -264
rect 421 -280 428 -264
rect 228 -287 428 -280
rect 556 -264 756 -250
rect 556 -280 563 -264
rect 749 -280 756 -264
rect 556 -287 756 -280
rect 884 -264 1084 -250
rect 884 -280 891 -264
rect 1077 -280 1084 -264
rect 884 -287 1084 -280
rect 1212 -264 1412 -250
rect 1212 -280 1219 -264
rect 1405 -280 1412 -264
rect 1212 -287 1412 -280
rect 1540 -264 1740 -250
rect 1540 -280 1547 -264
rect 1733 -280 1740 -264
rect 1540 -287 1740 -280
<< polycont >>
rect -93 264 93 280
rect 235 264 421 280
rect 563 264 749 280
rect 891 264 1077 280
rect 1219 264 1405 280
rect 1547 264 1733 280
rect -93 -280 93 -264
rect 235 -280 421 -264
rect 563 -280 749 -264
rect 891 -280 1077 -264
rect 1219 -280 1405 -264
rect 1547 -280 1733 -264
<< metal1 >>
rect -216 332 1856 337
rect -216 316 -181 332
rect 1821 316 1856 332
rect -216 311 1856 316
rect -216 302 -190 311
rect -216 -302 -211 302
rect -195 -302 -190 302
rect 1830 302 1856 311
rect -216 -311 -190 -302
rect 1830 -302 1835 302
rect 1851 -302 1856 302
rect 1830 -311 1856 -302
rect -216 -316 1856 -311
rect -216 -332 -181 -316
rect 1821 -332 1856 -316
rect -216 -337 1856 -332
<< properties >>
string gencell hvpmos
string library sg13g2_devstdin
string parameters w 5 l 2 nf 1 nx 6 dx 0.6 ny 1 dy 0.21 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1 glc 1 grc 1 gtc 1 gbc 1
<< end >>
