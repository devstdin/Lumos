magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752513657
<< metal1 >>
rect 13749 -469 16789 -201
rect 13749 -2812 13941 -469
rect 14251 -621 14623 -569
rect 14947 -621 15319 -569
rect 15643 -621 16015 -569
rect 16339 -621 16711 -569
rect 14121 -1006 14225 -653
rect 14121 -1186 14131 -1006
rect 14215 -1186 14225 -1006
rect 14121 -2625 14225 -1186
rect 14387 -1549 14487 -621
rect 14387 -1729 14397 -1549
rect 14478 -1729 14487 -1549
rect 14387 -2657 14487 -1729
rect 14649 -2092 14753 -653
rect 14649 -2272 14659 -2092
rect 14743 -2272 14753 -2092
rect 14649 -2625 14753 -2272
rect 14817 -1006 14921 -653
rect 14817 -1186 14827 -1006
rect 14911 -1186 14921 -1006
rect 14817 -2625 14921 -1186
rect 15083 -1549 15183 -621
rect 15083 -1729 15093 -1549
rect 15174 -1729 15183 -1549
rect 15083 -2657 15183 -1729
rect 15345 -2092 15449 -653
rect 15345 -2272 15355 -2092
rect 15439 -2272 15449 -2092
rect 15345 -2625 15449 -2272
rect 15513 -1006 15617 -653
rect 15513 -1186 15523 -1006
rect 15607 -1186 15617 -1006
rect 15513 -2625 15617 -1186
rect 15779 -1549 15879 -621
rect 15779 -1729 15789 -1549
rect 15870 -1729 15879 -1549
rect 15779 -2657 15879 -1729
rect 16041 -2092 16145 -653
rect 16041 -2272 16051 -2092
rect 16135 -2272 16145 -2092
rect 16041 -2625 16145 -2272
rect 16209 -1006 16313 -653
rect 16209 -1186 16219 -1006
rect 16303 -1186 16313 -1006
rect 16209 -2625 16313 -1186
rect 16475 -1549 16575 -621
rect 16475 -1729 16485 -1549
rect 16566 -1729 16575 -1549
rect 16475 -2657 16575 -1729
rect 16737 -2092 16841 -653
rect 16737 -2272 16747 -2092
rect 16831 -2272 16841 -2092
rect 16737 -2625 16841 -2272
rect 14251 -2709 14623 -2657
rect 14947 -2709 15319 -2657
rect 15643 -2709 16015 -2657
rect 16339 -2709 16711 -2657
rect 13749 -2830 16789 -2812
rect 13405 -3152 16789 -2830
rect 16965 -2998 17294 -2988
rect 16965 -3142 16975 -2998
rect 17155 -3142 17294 -2998
rect 16965 -3152 17294 -3142
rect 13405 -3308 14083 -3152
rect 14161 -3276 17133 -3224
rect 13405 -5280 14135 -3308
rect 15547 -4204 15747 -3276
rect 17211 -3308 17294 -3152
rect 15547 -4384 15557 -4204
rect 15737 -4384 15747 -4204
rect 13405 -5492 14083 -5280
rect 15547 -5312 15747 -4384
rect 17159 -5280 17294 -3308
rect 14161 -5460 17133 -5312
rect 13405 -7464 14135 -5492
rect 13405 -7676 14083 -7464
rect 15547 -7496 15747 -5460
rect 17211 -5492 17294 -5280
rect 17159 -7464 17294 -5492
rect 14161 -7644 17133 -7496
rect 13405 -9648 14135 -7676
rect 13405 -9860 14083 -9648
rect 15547 -9680 15747 -7644
rect 17211 -7676 17294 -7464
rect 17159 -9648 17294 -7676
rect 14161 -9828 17133 -9680
rect 13405 -11832 14135 -9860
rect 13405 -12044 14083 -11832
rect 15547 -11864 15747 -9828
rect 17211 -9860 17294 -9648
rect 17159 -11832 17294 -9860
rect 14161 -12012 17133 -11864
rect 13405 -14016 14135 -12044
rect 13405 -14228 14083 -14016
rect 15547 -14048 15747 -12012
rect 17211 -12044 17294 -11832
rect 17159 -14016 17294 -12044
rect 14161 -14196 17133 -14048
rect 13405 -16200 14135 -14228
rect 13405 -16388 14079 -16200
rect 15547 -16232 15747 -14196
rect 17211 -14228 17294 -14016
rect 17159 -16200 17294 -14228
rect 14161 -16284 17133 -16232
rect 17380 -16388 17938 -2852
rect 13405 -17053 17938 -16388
<< via1 >>
rect 14131 -1186 14215 -1006
rect 14397 -1729 14478 -1549
rect 14659 -2272 14743 -2092
rect 14827 -1186 14911 -1006
rect 15093 -1729 15174 -1549
rect 15355 -2272 15439 -2092
rect 15523 -1186 15607 -1006
rect 15789 -1729 15870 -1549
rect 16051 -2272 16135 -2092
rect 16219 -1186 16303 -1006
rect 16485 -1729 16566 -1549
rect 16747 -2272 16831 -2092
rect 16975 -3142 17155 -2998
rect 15557 -4384 15737 -4204
<< metal2 >>
rect 17053 -995 17940 -810
rect 16965 -996 17940 -995
rect 14121 -1006 17940 -996
rect 14121 -1186 14131 -1006
rect 14215 -1186 14827 -1006
rect 14911 -1186 15523 -1006
rect 15607 -1186 16219 -1006
rect 16303 -1186 17940 -1006
rect 14121 -1196 17940 -1186
rect 17053 -1384 17940 -1196
rect 13299 -1549 17938 -1539
rect 13299 -1729 14397 -1549
rect 14478 -1729 15093 -1549
rect 15174 -1729 15789 -1549
rect 15870 -1729 16485 -1549
rect 16566 -1729 17938 -1549
rect 13299 -1739 17938 -1729
rect 14121 -2092 17165 -2082
rect 14121 -2272 14659 -2092
rect 14743 -2272 15355 -2092
rect 15439 -2272 16051 -2092
rect 16135 -2272 16747 -2092
rect 16831 -2272 17165 -2092
rect 14121 -2282 17165 -2272
rect 16965 -2998 17165 -2282
rect 16965 -3142 16975 -2998
rect 17155 -3142 17165 -2998
rect 16965 -3152 17165 -3142
rect 13299 -4204 17938 -4194
rect 13299 -4384 15557 -4204
rect 15737 -4384 17938 -4204
rect 13299 -4394 17938 -4384
use hvnmos_QQE73P  hvnmos_QQE73P_2
timestamp 1748519341
transform 1 0 14437 0 1 -1639
box -544 -1222 2356 1222
use lvnmos_533TXK  lvnmos_533TXK_2
timestamp 1747683008
transform 1 0 15647 0 1 -15214
box -1754 -1218 1754 11994
<< labels >>
flabel metal2 17366 -1384 17940 -810 0 FreeSans 800 0 0 0 ISINK
port 6 nsew
flabel metal2 17549 -1739 17938 -1539 0 FreeSans 800 0 0 0 VSINKT
port 7 nsew
flabel metal2 17567 -4394 17938 -4194 0 FreeSans 800 0 0 0 VSINKB
port 9 nsew
flabel metal1 17646 -17053 17938 -16442 0 FreeSans 800 0 0 0 VSS
port 10 nsew
<< end >>
