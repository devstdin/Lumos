magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752866318
<< error_p >>
rect -36 544 -26 554
rect 26 544 36 554
rect 242 544 252 554
rect 304 544 314 554
rect 520 544 530 554
rect 582 544 592 554
rect 798 544 808 554
rect 860 544 870 554
rect -46 534 46 544
rect 232 534 324 544
rect 510 534 602 544
rect 788 534 880 544
rect -36 522 36 534
rect 242 522 314 534
rect 520 522 592 534
rect 798 522 870 534
rect -46 512 46 522
rect 232 512 324 522
rect 510 512 602 522
rect 788 512 880 522
rect -36 502 -26 512
rect 26 502 36 512
rect 242 502 252 512
rect 304 502 314 512
rect 520 502 530 512
rect 582 502 592 512
rect 798 502 808 512
rect 860 502 870 512
rect -104 470 -94 480
rect -82 470 -72 480
rect 72 470 82 480
rect 94 470 104 480
rect 174 470 184 480
rect 196 470 206 480
rect 350 470 360 480
rect 372 470 382 480
rect 452 470 462 480
rect 474 470 484 480
rect 628 470 638 480
rect 650 470 660 480
rect 730 470 740 480
rect 752 470 762 480
rect 906 470 916 480
rect 928 470 938 480
rect -114 460 -104 470
rect -72 460 -62 470
rect 62 460 72 470
rect 104 460 114 470
rect 164 460 174 470
rect 206 460 216 470
rect 340 460 350 470
rect 382 460 392 470
rect 442 460 452 470
rect 484 460 494 470
rect 618 460 628 470
rect 660 460 670 470
rect 720 460 730 470
rect 762 460 772 470
rect 896 460 906 470
rect 938 460 948 470
rect -114 298 -104 308
rect -72 298 -62 308
rect 62 298 72 308
rect 104 298 114 308
rect 164 298 174 308
rect 206 298 216 308
rect 340 298 350 308
rect 382 298 392 308
rect 442 298 452 308
rect 484 298 494 308
rect 618 298 628 308
rect 660 298 670 308
rect 720 298 730 308
rect 762 298 772 308
rect 896 298 906 308
rect 938 298 948 308
rect -104 288 -94 298
rect -82 288 -72 298
rect 72 288 82 298
rect 94 288 104 298
rect 174 288 184 298
rect 196 288 206 298
rect 350 288 360 298
rect 372 288 382 298
rect 452 288 462 298
rect 474 288 484 298
rect 628 288 638 298
rect 650 288 660 298
rect 730 288 740 298
rect 752 288 762 298
rect 906 288 916 298
rect 928 288 938 298
rect -36 256 -26 266
rect 26 256 36 266
rect 242 256 252 266
rect 304 256 314 266
rect 520 256 530 266
rect 582 256 592 266
rect 798 256 808 266
rect 860 256 870 266
rect -46 246 46 256
rect 232 246 324 256
rect 510 246 602 256
rect 788 246 880 256
rect -36 234 36 246
rect 242 234 314 246
rect 520 234 592 246
rect 798 234 870 246
rect -46 224 46 234
rect 232 224 324 234
rect 510 224 602 234
rect 788 224 880 234
rect -36 214 -26 224
rect 26 214 36 224
rect 242 214 252 224
rect 304 214 314 224
rect 520 214 530 224
rect 582 214 592 224
rect 798 214 808 224
rect 860 214 870 224
rect -36 160 -26 170
rect 26 160 36 170
rect 242 160 252 170
rect 304 160 314 170
rect 520 160 530 170
rect 582 160 592 170
rect 798 160 808 170
rect 860 160 870 170
rect -46 150 46 160
rect 232 150 324 160
rect 510 150 602 160
rect 788 150 880 160
rect -36 138 36 150
rect 242 138 314 150
rect 520 138 592 150
rect 798 138 870 150
rect -46 128 46 138
rect 232 128 324 138
rect 510 128 602 138
rect 788 128 880 138
rect -36 118 -26 128
rect 26 118 36 128
rect 242 118 252 128
rect 304 118 314 128
rect 520 118 530 128
rect 582 118 592 128
rect 798 118 808 128
rect 860 118 870 128
rect -104 86 -94 96
rect -82 86 -72 96
rect 72 86 82 96
rect 94 86 104 96
rect 174 86 184 96
rect 196 86 206 96
rect 350 86 360 96
rect 372 86 382 96
rect 452 86 462 96
rect 474 86 484 96
rect 628 86 638 96
rect 650 86 660 96
rect 730 86 740 96
rect 752 86 762 96
rect 906 86 916 96
rect 928 86 938 96
rect -114 76 -104 86
rect -72 76 -62 86
rect 62 76 72 86
rect 104 76 114 86
rect 164 76 174 86
rect 206 76 216 86
rect 340 76 350 86
rect 382 76 392 86
rect 442 76 452 86
rect 484 76 494 86
rect 618 76 628 86
rect 660 76 670 86
rect 720 76 730 86
rect 762 76 772 86
rect 896 76 906 86
rect 938 76 948 86
rect -114 -86 -104 -76
rect -72 -86 -62 -76
rect 62 -86 72 -76
rect 104 -86 114 -76
rect 164 -86 174 -76
rect 206 -86 216 -76
rect 340 -86 350 -76
rect 382 -86 392 -76
rect 442 -86 452 -76
rect 484 -86 494 -76
rect 618 -86 628 -76
rect 660 -86 670 -76
rect 720 -86 730 -76
rect 762 -86 772 -76
rect 896 -86 906 -76
rect 938 -86 948 -76
rect -104 -96 -94 -86
rect -82 -96 -72 -86
rect 72 -96 82 -86
rect 94 -96 104 -86
rect 174 -96 184 -86
rect 196 -96 206 -86
rect 350 -96 360 -86
rect 372 -96 382 -86
rect 452 -96 462 -86
rect 474 -96 484 -86
rect 628 -96 638 -86
rect 650 -96 660 -86
rect 730 -96 740 -86
rect 752 -96 762 -86
rect 906 -96 916 -86
rect 928 -96 938 -86
rect -36 -128 -26 -118
rect 26 -128 36 -118
rect 242 -128 252 -118
rect 304 -128 314 -118
rect 520 -128 530 -118
rect 582 -128 592 -118
rect 798 -128 808 -118
rect 860 -128 870 -118
rect -46 -138 46 -128
rect 232 -138 324 -128
rect 510 -138 602 -128
rect 788 -138 880 -128
rect -36 -150 36 -138
rect 242 -150 314 -138
rect 520 -150 592 -138
rect 798 -150 870 -138
rect -46 -160 46 -150
rect 232 -160 324 -150
rect 510 -160 602 -150
rect 788 -160 880 -150
rect -36 -170 -26 -160
rect 26 -170 36 -160
rect 242 -170 252 -160
rect 304 -170 314 -160
rect 520 -170 530 -160
rect 582 -170 592 -160
rect 798 -170 808 -160
rect 860 -170 870 -160
<< nmos >>
rect -50 284 50 484
rect 228 284 328 484
rect 506 284 606 484
rect 784 284 884 484
rect -50 -100 50 100
rect 228 -100 328 100
rect 506 -100 606 100
rect 784 -100 884 100
<< ndiff >>
rect -118 470 -50 484
rect -118 298 -104 470
rect -72 298 -50 470
rect -118 284 -50 298
rect 50 470 118 484
rect 50 298 72 470
rect 104 298 118 470
rect 50 284 118 298
rect 160 470 228 484
rect 160 298 174 470
rect 206 298 228 470
rect 160 284 228 298
rect 328 470 396 484
rect 328 298 350 470
rect 382 298 396 470
rect 328 284 396 298
rect 438 470 506 484
rect 438 298 452 470
rect 484 298 506 470
rect 438 284 506 298
rect 606 470 674 484
rect 606 298 628 470
rect 660 298 674 470
rect 606 284 674 298
rect 716 470 784 484
rect 716 298 730 470
rect 762 298 784 470
rect 716 284 784 298
rect 884 470 952 484
rect 884 298 906 470
rect 938 298 952 470
rect 884 284 952 298
rect -118 86 -50 100
rect -118 -86 -104 86
rect -72 -86 -50 86
rect -118 -100 -50 -86
rect 50 86 118 100
rect 50 -86 72 86
rect 104 -86 118 86
rect 50 -100 118 -86
rect 160 86 228 100
rect 160 -86 174 86
rect 206 -86 228 86
rect 160 -100 228 -86
rect 328 86 396 100
rect 328 -86 350 86
rect 382 -86 396 86
rect 328 -100 396 -86
rect 438 86 506 100
rect 438 -86 452 86
rect 484 -86 506 86
rect 438 -100 506 -86
rect 606 86 674 100
rect 606 -86 628 86
rect 660 -86 674 86
rect 606 -100 674 -86
rect 716 86 784 100
rect 716 -86 730 86
rect 762 -86 784 86
rect 716 -100 784 -86
rect 884 86 952 100
rect 884 -86 906 86
rect 938 -86 952 86
rect 884 -100 952 -86
<< ndiffc >>
rect -104 298 -72 470
rect 72 298 104 470
rect 174 298 206 470
rect 350 298 382 470
rect 452 298 484 470
rect 628 298 660 470
rect 730 298 762 470
rect 906 298 938 470
rect -104 -86 -72 86
rect 72 -86 104 86
rect 174 -86 206 86
rect 350 -86 382 86
rect 452 -86 484 86
rect 628 -86 660 86
rect 730 -86 762 86
rect 906 -86 938 86
<< psubdiff >>
rect -241 646 1075 660
rect -241 614 -167 646
rect 1001 614 1075 646
rect -241 600 1075 614
rect -241 586 -181 600
rect -241 -202 -227 586
rect -195 -202 -181 586
rect 1015 586 1075 600
rect -241 -216 -181 -202
rect 1015 -202 1029 586
rect 1061 -202 1075 586
rect 1015 -216 1075 -202
rect -241 -230 1075 -216
rect -241 -262 -167 -230
rect 1001 -262 1075 -230
rect -241 -276 1075 -262
<< psubdiffcont >>
rect -167 614 1001 646
rect -227 -202 -195 586
rect 1029 -202 1061 586
rect -167 -262 1001 -230
<< poly >>
rect -50 544 50 558
rect -50 512 -36 544
rect 36 512 50 544
rect -50 484 50 512
rect 228 544 328 558
rect 228 512 242 544
rect 314 512 328 544
rect 228 484 328 512
rect 506 544 606 558
rect 506 512 520 544
rect 592 512 606 544
rect 506 484 606 512
rect 784 544 884 558
rect 784 512 798 544
rect 870 512 884 544
rect 784 484 884 512
rect -50 256 50 284
rect -50 224 -36 256
rect 36 224 50 256
rect -50 210 50 224
rect 228 256 328 284
rect 228 224 242 256
rect 314 224 328 256
rect 228 210 328 224
rect 506 256 606 284
rect 506 224 520 256
rect 592 224 606 256
rect 506 210 606 224
rect 784 256 884 284
rect 784 224 798 256
rect 870 224 884 256
rect 784 210 884 224
rect -50 160 50 174
rect -50 128 -36 160
rect 36 128 50 160
rect -50 100 50 128
rect 228 160 328 174
rect 228 128 242 160
rect 314 128 328 160
rect 228 100 328 128
rect 506 160 606 174
rect 506 128 520 160
rect 592 128 606 160
rect 506 100 606 128
rect 784 160 884 174
rect 784 128 798 160
rect 870 128 884 160
rect 784 100 884 128
rect -50 -128 50 -100
rect -50 -160 -36 -128
rect 36 -160 50 -128
rect -50 -174 50 -160
rect 228 -128 328 -100
rect 228 -160 242 -128
rect 314 -160 328 -128
rect 228 -174 328 -160
rect 506 -128 606 -100
rect 506 -160 520 -128
rect 592 -160 606 -128
rect 506 -174 606 -160
rect 784 -128 884 -100
rect 784 -160 798 -128
rect 870 -160 884 -128
rect 784 -174 884 -160
<< polycont >>
rect -36 512 36 544
rect 242 512 314 544
rect 520 512 592 544
rect 798 512 870 544
rect -36 224 36 256
rect 242 224 314 256
rect 520 224 592 256
rect 798 224 870 256
rect -36 128 36 160
rect 242 128 314 160
rect 520 128 592 160
rect 798 128 870 160
rect -36 -160 36 -128
rect 242 -160 314 -128
rect 520 -160 592 -128
rect 798 -160 870 -128
<< metal1 >>
rect -237 646 1071 656
rect -237 614 -167 646
rect 1001 614 1071 646
rect -237 604 1071 614
rect -237 586 -185 604
rect -237 -202 -227 586
rect -195 -202 -185 586
rect 1019 586 1071 604
rect -237 -220 -185 -202
rect 1019 -202 1029 586
rect 1061 -202 1071 586
rect 1019 -220 1071 -202
rect -237 -230 1071 -220
rect -237 -262 -167 -230
rect 1001 -262 1071 -230
rect -237 -272 1071 -262
<< properties >>
string gencell lvnmos
string library sg13g2_devstdin
string parameters w 1 l 0.5 nf 1 nx 4 dx 0.21 ny 2 dy 0.18 wmin 0.50 lmin 0.50 class mosfet gcontcov_t 100 gcontcov_b 100 dcontcov_l 100 dcontcov_r 100 guard_distf 1.5 glc 1 grc 1 gtc 1 gbc 1
<< end >>
