magic
tech ihp-sg13g2
timestamp 1747597098
<< nwell >>
rect -325 -325 325 325
<< psubdiff >>
rect -379 372 379 379
rect -379 356 -342 372
rect 342 356 379 372
rect -379 349 379 356
rect -379 342 -349 349
rect -379 -342 -372 342
rect -356 -342 -349 342
rect 349 342 379 349
rect -379 -349 -349 -342
rect 349 -342 356 342
rect 372 -342 379 342
rect 349 -349 379 -342
rect -379 -356 379 -349
rect -379 -372 -342 -356
rect 342 -372 379 -356
rect -379 -379 379 -372
<< nsubdiff >>
rect -301 294 301 301
rect -301 278 -264 294
rect 264 278 301 294
rect -301 271 301 278
rect -301 264 -271 271
rect -301 -264 -294 264
rect -278 -264 -271 264
rect 271 264 301 271
rect -301 -271 -271 -264
rect 271 -264 278 264
rect 294 -264 301 264
rect 271 -271 301 -264
rect -301 -278 301 -271
rect -301 -294 -264 -278
rect 264 -294 301 -278
rect -301 -301 301 -294
<< psubdiffcont >>
rect -342 356 342 372
rect -372 -342 -356 342
rect 356 -342 372 342
rect -342 -372 342 -356
<< nsubdiffcont >>
rect -264 278 264 294
rect -294 -264 -278 264
rect 278 -264 294 264
rect -264 -294 264 -278
<< pdiode >>
rect -250 243 250 250
rect -250 -243 -243 243
rect 243 -243 250 243
rect -250 -250 250 -243
<< pdiodecont >>
rect -243 -243 243 243
<< metal1 >>
rect -377 372 377 377
rect -377 356 -342 372
rect 342 356 377 372
rect -377 351 377 356
rect -377 342 -351 351
rect -377 -342 -372 342
rect -356 -342 -351 342
rect 351 342 377 351
rect -299 294 299 299
rect -299 278 -264 294
rect 264 278 299 294
rect -299 273 299 278
rect -299 264 -273 273
rect -299 -264 -294 264
rect -278 -264 -273 264
rect 273 264 299 273
rect -299 -273 -273 -264
rect 273 -264 278 264
rect 294 -264 299 264
rect 273 -273 299 -264
rect -299 -278 299 -273
rect -299 -294 -264 -278
rect 264 -294 299 -278
rect -299 -299 299 -294
rect -377 -351 -351 -342
rect 351 -342 356 342
rect 372 -342 377 342
rect 351 -351 377 -342
rect -377 -356 377 -351
rect -377 -372 -342 -356
rect 342 -372 377 -356
rect -377 -377 377 -372
<< properties >>
string gencell dpantenna
string library sg13g2_devstdin
string parameters w 5 l 5 nx 1 dx 0.18 ny 1 dy 0.18 wmin 0.50 lmin 0.50 class diode contcov 0 glc 1 grc 1 gtc 1 gbc 1
<< end >>
