magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755542813
<< checkpaint >>
rect -2124 -3692 3470 5854
<< nwell >>
rect -124 2500 1470 3854
<< pwell >>
rect -5 1756 543 2402
rect -26 1644 1372 1756
<< nmos >>
rect 89 1826 115 2376
<< pmos >>
rect 89 2624 115 3574
<< hvnmos >>
rect 359 1846 449 2376
<< hvpmos >>
rect 359 2624 449 3554
<< ndiff >>
rect 21 2355 89 2376
rect 21 2323 35 2355
rect 67 2323 89 2355
rect 21 2287 89 2323
rect 21 2255 35 2287
rect 67 2255 89 2287
rect 21 2219 89 2255
rect 21 2187 35 2219
rect 67 2187 89 2219
rect 21 2151 89 2187
rect 21 2119 35 2151
rect 67 2119 89 2151
rect 21 2083 89 2119
rect 21 2051 35 2083
rect 67 2051 89 2083
rect 21 2015 89 2051
rect 21 1983 35 2015
rect 67 1983 89 2015
rect 21 1947 89 1983
rect 21 1915 35 1947
rect 67 1915 89 1947
rect 21 1879 89 1915
rect 21 1847 35 1879
rect 67 1847 89 1879
rect 21 1826 89 1847
rect 115 2355 183 2376
rect 115 2323 137 2355
rect 169 2323 183 2355
rect 115 2287 183 2323
rect 115 2255 137 2287
rect 169 2255 183 2287
rect 115 2219 183 2255
rect 115 2187 137 2219
rect 169 2187 183 2219
rect 115 2151 183 2187
rect 115 2119 137 2151
rect 169 2119 183 2151
rect 115 2083 183 2119
rect 115 2051 137 2083
rect 169 2051 183 2083
rect 115 2015 183 2051
rect 115 1983 137 2015
rect 169 1983 183 2015
rect 115 1947 183 1983
rect 115 1915 137 1947
rect 169 1915 183 1947
rect 115 1879 183 1915
rect 115 1847 137 1879
rect 169 1847 183 1879
rect 115 1826 183 1847
<< pdiff >>
rect 21 3557 89 3574
rect 21 3525 35 3557
rect 67 3525 89 3557
rect 21 3489 89 3525
rect 21 3457 35 3489
rect 67 3457 89 3489
rect 21 3421 89 3457
rect 21 3389 35 3421
rect 67 3389 89 3421
rect 21 3353 89 3389
rect 21 3321 35 3353
rect 67 3321 89 3353
rect 21 3285 89 3321
rect 21 3253 35 3285
rect 67 3253 89 3285
rect 21 3217 89 3253
rect 21 3185 35 3217
rect 67 3185 89 3217
rect 21 3149 89 3185
rect 21 3117 35 3149
rect 67 3117 89 3149
rect 21 3081 89 3117
rect 21 3049 35 3081
rect 67 3049 89 3081
rect 21 3013 89 3049
rect 21 2981 35 3013
rect 67 2981 89 3013
rect 21 2945 89 2981
rect 21 2913 35 2945
rect 67 2913 89 2945
rect 21 2877 89 2913
rect 21 2845 35 2877
rect 67 2845 89 2877
rect 21 2809 89 2845
rect 21 2777 35 2809
rect 67 2777 89 2809
rect 21 2741 89 2777
rect 21 2709 35 2741
rect 67 2709 89 2741
rect 21 2673 89 2709
rect 21 2641 35 2673
rect 67 2641 89 2673
rect 21 2624 89 2641
rect 115 3557 183 3574
rect 115 3525 137 3557
rect 169 3525 183 3557
rect 115 3489 183 3525
rect 115 3457 137 3489
rect 169 3457 183 3489
rect 115 3421 183 3457
rect 115 3389 137 3421
rect 169 3389 183 3421
rect 115 3353 183 3389
rect 115 3321 137 3353
rect 169 3321 183 3353
rect 115 3285 183 3321
rect 115 3253 137 3285
rect 169 3253 183 3285
rect 115 3217 183 3253
rect 115 3185 137 3217
rect 169 3185 183 3217
rect 115 3149 183 3185
rect 115 3117 137 3149
rect 169 3117 183 3149
rect 115 3081 183 3117
rect 115 3049 137 3081
rect 169 3049 183 3081
rect 115 3013 183 3049
rect 115 2981 137 3013
rect 169 2981 183 3013
rect 115 2945 183 2981
rect 115 2913 137 2945
rect 169 2913 183 2945
rect 115 2877 183 2913
rect 115 2845 137 2877
rect 169 2845 183 2877
rect 115 2809 183 2845
rect 115 2777 137 2809
rect 169 2777 183 2809
rect 115 2741 183 2777
rect 115 2709 137 2741
rect 169 2709 183 2741
rect 115 2673 183 2709
rect 115 2641 137 2673
rect 169 2641 183 2673
rect 115 2624 183 2641
<< hvndiff >>
rect 291 2331 359 2376
rect 291 2299 305 2331
rect 337 2299 359 2331
rect 291 2263 359 2299
rect 291 2231 305 2263
rect 337 2231 359 2263
rect 291 2195 359 2231
rect 291 2163 305 2195
rect 337 2163 359 2195
rect 291 2127 359 2163
rect 291 2095 305 2127
rect 337 2095 359 2127
rect 291 2059 359 2095
rect 291 2027 305 2059
rect 337 2027 359 2059
rect 291 1991 359 2027
rect 291 1959 305 1991
rect 337 1959 359 1991
rect 291 1923 359 1959
rect 291 1891 305 1923
rect 337 1891 359 1923
rect 291 1846 359 1891
rect 449 2331 517 2376
rect 449 2299 471 2331
rect 503 2299 517 2331
rect 449 2263 517 2299
rect 449 2231 471 2263
rect 503 2231 517 2263
rect 449 2195 517 2231
rect 449 2163 471 2195
rect 503 2163 517 2195
rect 449 2127 517 2163
rect 449 2095 471 2127
rect 503 2095 517 2127
rect 449 2059 517 2095
rect 449 2027 471 2059
rect 503 2027 517 2059
rect 449 1991 517 2027
rect 449 1959 471 1991
rect 503 1959 517 1991
rect 449 1923 517 1959
rect 449 1891 471 1923
rect 503 1891 517 1923
rect 449 1846 517 1891
<< hvpdiff >>
rect 291 3513 359 3554
rect 291 3481 305 3513
rect 337 3481 359 3513
rect 291 3445 359 3481
rect 291 3413 305 3445
rect 337 3413 359 3445
rect 291 3377 359 3413
rect 291 3345 305 3377
rect 337 3345 359 3377
rect 291 3309 359 3345
rect 291 3277 305 3309
rect 337 3277 359 3309
rect 291 3241 359 3277
rect 291 3209 305 3241
rect 337 3209 359 3241
rect 291 3173 359 3209
rect 291 3141 305 3173
rect 337 3141 359 3173
rect 291 3105 359 3141
rect 291 3073 305 3105
rect 337 3073 359 3105
rect 291 3037 359 3073
rect 291 3005 305 3037
rect 337 3005 359 3037
rect 291 2969 359 3005
rect 291 2937 305 2969
rect 337 2937 359 2969
rect 291 2901 359 2937
rect 291 2869 305 2901
rect 337 2869 359 2901
rect 291 2833 359 2869
rect 291 2801 305 2833
rect 337 2801 359 2833
rect 291 2765 359 2801
rect 291 2733 305 2765
rect 337 2733 359 2765
rect 291 2697 359 2733
rect 291 2665 305 2697
rect 337 2665 359 2697
rect 291 2624 359 2665
rect 449 3513 517 3554
rect 449 3481 471 3513
rect 503 3481 517 3513
rect 449 3445 517 3481
rect 449 3413 471 3445
rect 503 3413 517 3445
rect 449 3377 517 3413
rect 449 3345 471 3377
rect 503 3345 517 3377
rect 449 3309 517 3345
rect 449 3277 471 3309
rect 503 3277 517 3309
rect 449 3241 517 3277
rect 449 3209 471 3241
rect 503 3209 517 3241
rect 449 3173 517 3209
rect 449 3141 471 3173
rect 503 3141 517 3173
rect 449 3105 517 3141
rect 449 3073 471 3105
rect 503 3073 517 3105
rect 449 3037 517 3073
rect 449 3005 471 3037
rect 503 3005 517 3037
rect 449 2969 517 3005
rect 449 2937 471 2969
rect 503 2937 517 2969
rect 449 2901 517 2937
rect 449 2869 471 2901
rect 503 2869 517 2901
rect 449 2833 517 2869
rect 449 2801 471 2833
rect 503 2801 517 2833
rect 449 2765 517 2801
rect 449 2733 471 2765
rect 503 2733 517 2765
rect 449 2697 517 2733
rect 449 2665 471 2697
rect 503 2665 517 2697
rect 449 2624 517 2665
<< ndiffc >>
rect 35 2323 67 2355
rect 35 2255 67 2287
rect 35 2187 67 2219
rect 35 2119 67 2151
rect 35 2051 67 2083
rect 35 1983 67 2015
rect 35 1915 67 1947
rect 35 1847 67 1879
rect 137 2323 169 2355
rect 137 2255 169 2287
rect 137 2187 169 2219
rect 137 2119 169 2151
rect 137 2051 169 2083
rect 137 1983 169 2015
rect 137 1915 169 1947
rect 137 1847 169 1879
<< pdiffc >>
rect 35 3525 67 3557
rect 35 3457 67 3489
rect 35 3389 67 3421
rect 35 3321 67 3353
rect 35 3253 67 3285
rect 35 3185 67 3217
rect 35 3117 67 3149
rect 35 3049 67 3081
rect 35 2981 67 3013
rect 35 2913 67 2945
rect 35 2845 67 2877
rect 35 2777 67 2809
rect 35 2709 67 2741
rect 35 2641 67 2673
rect 137 3525 169 3557
rect 137 3457 169 3489
rect 137 3389 169 3421
rect 137 3321 169 3353
rect 137 3253 169 3285
rect 137 3185 169 3217
rect 137 3117 169 3149
rect 137 3049 169 3081
rect 137 2981 169 3013
rect 137 2913 169 2945
rect 137 2845 169 2877
rect 137 2777 169 2809
rect 137 2709 169 2741
rect 137 2641 169 2673
<< hvndiffc >>
rect 305 2299 337 2331
rect 305 2231 337 2263
rect 305 2163 337 2195
rect 305 2095 337 2127
rect 305 2027 337 2059
rect 305 1959 337 1991
rect 305 1891 337 1923
rect 471 2299 503 2331
rect 471 2231 503 2263
rect 471 2163 503 2195
rect 471 2095 503 2127
rect 471 2027 503 2059
rect 471 1959 503 1991
rect 471 1891 503 1923
<< hvpdiffc >>
rect 305 3481 337 3513
rect 305 3413 337 3445
rect 305 3345 337 3377
rect 305 3277 337 3309
rect 305 3209 337 3241
rect 305 3141 337 3173
rect 305 3073 337 3105
rect 305 3005 337 3037
rect 305 2937 337 2969
rect 305 2869 337 2901
rect 305 2801 337 2833
rect 305 2733 337 2765
rect 305 2665 337 2697
rect 471 3481 503 3513
rect 471 3413 503 3445
rect 471 3345 503 3377
rect 471 3277 503 3309
rect 471 3209 503 3241
rect 471 3141 503 3173
rect 471 3073 503 3105
rect 471 3005 503 3037
rect 471 2937 503 2969
rect 471 2869 503 2901
rect 471 2801 503 2833
rect 471 2733 503 2765
rect 471 2665 503 2697
<< psubdiff >>
rect 0 1716 1346 1730
rect 0 1684 45 1716
rect 77 1684 113 1716
rect 145 1684 181 1716
rect 213 1684 249 1716
rect 281 1684 317 1716
rect 349 1684 385 1716
rect 417 1684 453 1716
rect 485 1684 521 1716
rect 553 1684 589 1716
rect 621 1684 657 1716
rect 689 1684 725 1716
rect 757 1684 793 1716
rect 825 1684 861 1716
rect 893 1684 929 1716
rect 961 1684 997 1716
rect 1029 1684 1065 1716
rect 1097 1684 1133 1716
rect 1165 1684 1201 1716
rect 1233 1684 1269 1716
rect 1301 1684 1346 1716
rect 0 1670 1346 1684
<< nsubdiff >>
rect 0 3716 1346 3730
rect 0 3684 45 3716
rect 77 3684 113 3716
rect 145 3684 181 3716
rect 213 3684 249 3716
rect 281 3684 317 3716
rect 349 3684 385 3716
rect 417 3684 453 3716
rect 485 3684 521 3716
rect 553 3684 589 3716
rect 621 3684 657 3716
rect 689 3684 725 3716
rect 757 3684 793 3716
rect 825 3684 861 3716
rect 893 3684 929 3716
rect 961 3684 997 3716
rect 1029 3684 1065 3716
rect 1097 3684 1133 3716
rect 1165 3684 1201 3716
rect 1233 3684 1269 3716
rect 1301 3684 1346 3716
rect 0 3670 1346 3684
<< psubdiffcont >>
rect 45 1684 77 1716
rect 113 1684 145 1716
rect 181 1684 213 1716
rect 249 1684 281 1716
rect 317 1684 349 1716
rect 385 1684 417 1716
rect 453 1684 485 1716
rect 521 1684 553 1716
rect 589 1684 621 1716
rect 657 1684 689 1716
rect 725 1684 757 1716
rect 793 1684 825 1716
rect 861 1684 893 1716
rect 929 1684 961 1716
rect 997 1684 1029 1716
rect 1065 1684 1097 1716
rect 1133 1684 1165 1716
rect 1201 1684 1233 1716
rect 1269 1684 1301 1716
<< nsubdiffcont >>
rect 45 3684 77 3716
rect 113 3684 145 3716
rect 181 3684 213 3716
rect 249 3684 281 3716
rect 317 3684 349 3716
rect 385 3684 417 3716
rect 453 3684 485 3716
rect 521 3684 553 3716
rect 589 3684 621 3716
rect 657 3684 689 3716
rect 725 3684 757 3716
rect 793 3684 825 3716
rect 861 3684 893 3716
rect 929 3684 961 3716
rect 997 3684 1029 3716
rect 1065 3684 1097 3716
rect 1133 3684 1165 3716
rect 1201 3684 1233 3716
rect 1269 3684 1301 3716
<< poly >>
rect 89 3574 115 3610
rect 359 3554 449 3590
rect 89 2530 115 2624
rect 89 2516 175 2530
rect 89 2484 129 2516
rect 161 2484 175 2516
rect 89 2470 175 2484
rect 359 2516 449 2624
rect 359 2484 403 2516
rect 435 2484 449 2516
rect 89 2376 115 2470
rect 359 2376 449 2484
rect 89 1790 115 1826
rect 359 1810 449 1846
<< polycont >>
rect 129 2484 161 2516
rect 403 2484 435 2516
<< metal1 >>
rect 0 3716 1346 3721
rect 0 3684 45 3716
rect 77 3684 113 3716
rect 145 3684 181 3716
rect 213 3684 249 3716
rect 281 3684 317 3716
rect 349 3684 385 3716
rect 417 3684 453 3716
rect 485 3684 521 3716
rect 553 3684 589 3716
rect 621 3684 657 3716
rect 689 3684 725 3716
rect 757 3684 793 3716
rect 825 3684 861 3716
rect 893 3684 929 3716
rect 961 3684 997 3716
rect 1029 3684 1065 3716
rect 1097 3684 1133 3716
rect 1165 3684 1201 3716
rect 1233 3684 1269 3716
rect 1301 3684 1346 3716
rect 0 3679 1346 3684
rect 35 3557 67 3573
rect 35 3489 67 3525
rect 35 3421 67 3457
rect 35 3353 67 3389
rect 35 3285 67 3321
rect 35 3217 67 3253
rect 35 3149 67 3185
rect 35 3081 67 3117
rect 35 3013 67 3049
rect 35 2945 67 2981
rect 35 2877 67 2913
rect 35 2809 67 2845
rect 35 2741 67 2777
rect 35 2673 67 2709
rect 35 2355 67 2641
rect 137 3557 337 3679
rect 169 3525 337 3557
rect 137 3513 337 3525
rect 137 3489 305 3513
rect 169 3481 305 3489
rect 169 3457 337 3481
rect 137 3445 337 3457
rect 137 3421 305 3445
rect 169 3413 305 3421
rect 169 3389 337 3413
rect 137 3377 337 3389
rect 137 3353 305 3377
rect 169 3345 305 3353
rect 169 3321 337 3345
rect 137 3309 337 3321
rect 137 3285 305 3309
rect 169 3277 305 3285
rect 169 3253 337 3277
rect 137 3241 337 3253
rect 137 3217 305 3241
rect 169 3209 305 3217
rect 169 3185 337 3209
rect 137 3173 337 3185
rect 137 3149 305 3173
rect 169 3141 305 3149
rect 169 3117 337 3141
rect 137 3105 337 3117
rect 137 3081 305 3105
rect 169 3073 305 3081
rect 169 3049 337 3073
rect 137 3037 337 3049
rect 137 3013 305 3037
rect 169 3005 305 3013
rect 169 2981 337 3005
rect 137 2969 337 2981
rect 137 2945 305 2969
rect 169 2937 305 2945
rect 169 2913 337 2937
rect 137 2901 337 2913
rect 137 2877 305 2901
rect 169 2869 305 2877
rect 169 2845 337 2869
rect 137 2833 337 2845
rect 137 2809 305 2833
rect 169 2801 305 2809
rect 169 2777 337 2801
rect 137 2765 337 2777
rect 137 2741 305 2765
rect 169 2733 305 2741
rect 169 2709 337 2733
rect 137 2697 337 2709
rect 137 2673 305 2697
rect 169 2665 305 2673
rect 169 2649 337 2665
rect 471 3513 539 3529
rect 503 3481 539 3513
rect 471 3445 539 3481
rect 503 3413 539 3445
rect 471 3377 539 3413
rect 503 3345 539 3377
rect 471 3309 539 3345
rect 503 3277 539 3309
rect 471 3241 539 3277
rect 503 3209 539 3241
rect 471 3173 539 3209
rect 503 3141 539 3173
rect 471 3105 539 3141
rect 503 3073 539 3105
rect 471 3037 539 3073
rect 503 3005 539 3037
rect 471 2969 539 3005
rect 503 2937 539 2969
rect 471 2901 539 2937
rect 503 2869 539 2901
rect 471 2833 539 2869
rect 503 2801 539 2833
rect 471 2765 539 2801
rect 503 2733 539 2765
rect 471 2697 539 2733
rect 503 2665 539 2697
rect 471 2649 539 2665
rect 137 2625 169 2641
rect 503 2629 539 2649
rect 503 2620 545 2629
rect 503 2580 504 2620
rect 544 2580 545 2620
rect 503 2571 545 2580
rect 119 2520 267 2521
rect 119 2516 128 2520
rect 113 2484 128 2516
rect 119 2480 128 2484
rect 168 2480 267 2520
rect 119 2479 267 2480
rect 303 2520 451 2521
rect 303 2480 402 2520
rect 442 2480 451 2520
rect 303 2479 451 2480
rect 35 2287 67 2323
rect 35 2219 67 2255
rect 35 2151 67 2187
rect 35 2083 67 2119
rect 35 2015 67 2051
rect 35 1947 67 1983
rect 35 1879 67 1915
rect 35 1831 67 1847
rect 137 2355 169 2371
rect 503 2347 539 2571
rect 169 2331 337 2347
rect 169 2323 305 2331
rect 137 2299 305 2323
rect 137 2287 337 2299
rect 169 2263 337 2287
rect 169 2255 305 2263
rect 137 2231 305 2255
rect 137 2219 337 2231
rect 169 2195 337 2219
rect 169 2187 305 2195
rect 137 2163 305 2187
rect 137 2151 337 2163
rect 169 2127 337 2151
rect 169 2119 305 2127
rect 137 2095 305 2119
rect 137 2083 337 2095
rect 169 2059 337 2083
rect 169 2051 305 2059
rect 137 2027 305 2051
rect 137 2015 337 2027
rect 169 1991 337 2015
rect 169 1983 305 1991
rect 137 1959 305 1983
rect 137 1947 337 1959
rect 169 1923 337 1947
rect 169 1915 305 1923
rect 137 1891 305 1915
rect 137 1879 337 1891
rect 169 1847 337 1879
rect 471 2331 539 2347
rect 503 2299 539 2331
rect 471 2263 539 2299
rect 503 2231 539 2263
rect 471 2195 539 2231
rect 503 2163 539 2195
rect 471 2127 539 2163
rect 503 2095 539 2127
rect 471 2059 539 2095
rect 503 2027 539 2059
rect 471 1991 539 2027
rect 503 1959 539 1991
rect 471 1923 539 1959
rect 503 1891 539 1923
rect 471 1875 539 1891
rect 137 1721 337 1847
rect 0 1716 1346 1721
rect 0 1684 45 1716
rect 77 1684 113 1716
rect 145 1684 181 1716
rect 213 1684 249 1716
rect 281 1684 317 1716
rect 349 1684 385 1716
rect 417 1684 453 1716
rect 485 1684 521 1716
rect 553 1684 589 1716
rect 621 1684 657 1716
rect 689 1684 725 1716
rect 757 1684 793 1716
rect 825 1684 861 1716
rect 893 1684 929 1716
rect 961 1684 997 1716
rect 1029 1684 1065 1716
rect 1097 1684 1133 1716
rect 1165 1684 1201 1716
rect 1233 1684 1269 1716
rect 1301 1684 1346 1716
rect 0 1679 1346 1684
rect 0 -21 1346 21
<< via1 >>
rect 504 2580 544 2620
rect 128 2516 168 2520
rect 128 2484 129 2516
rect 129 2484 161 2516
rect 161 2484 168 2516
rect 128 2480 168 2484
rect 402 2516 442 2520
rect 402 2484 403 2516
rect 403 2484 435 2516
rect 435 2484 442 2516
rect 402 2480 442 2484
<< metal2 >>
rect 128 2620 544 2629
rect 128 2580 504 2620
rect 128 2571 544 2580
rect 128 2520 168 2571
rect 128 2471 168 2480
rect 402 2520 442 2529
rect 402 30 442 2480
rect 204 -1666 372 -1416
rect 535 -1582 909 -1360
use sg13g2_SecondaryProtection  sg13g2_SecondaryProtection_0
timestamp 1755542813
transform 1 0 0 0 1 -1666
box -124 -26 1448 1820
<< labels >>
flabel metal2 s 535 -1582 909 -1360 0 FreeSans 800 0 0 0 iovss
port 4 nsew
rlabel metal2 s 204 -1666 372 -1416 4 pad
port 5 nsew
rlabel metal1 s 0 -21 1346 21 4 iovdd
port 3 nsew
rlabel metal1 s 0 3679 1346 3721 4 vdd
port 1 nsew
rlabel metal1 s 0 1679 1346 1721 4 vss
port 2 nsew
rlabel metal1 s 35 1831 67 3573 4 core
port 6 nsew
flabel comment s 1224 1697 1224 1697 0 FreeSans 1600 0 0 0 sub!
<< properties >>
string device primitive
string GDS_END 17361714
string GDS_FILE sg13g2_io.gds
string GDS_START 17351042
<< end >>
