magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 1 56 447 292
rect -26 -56 506 56
<< nmos >>
rect 95 156 121 266
rect 203 118 229 266
rect 305 118 331 266
<< pmos >>
rect 95 412 121 580
rect 203 412 229 636
rect 305 412 331 636
<< ndiff >>
rect 27 226 95 266
rect 27 194 41 226
rect 73 194 95 226
rect 27 156 95 194
rect 121 174 203 266
rect 121 156 149 174
rect 135 142 149 156
rect 181 142 203 174
rect 135 118 203 142
rect 229 118 305 266
rect 331 252 421 266
rect 331 220 375 252
rect 407 220 421 252
rect 331 164 421 220
rect 331 132 375 164
rect 407 132 421 164
rect 331 118 421 132
<< pdiff >>
rect 135 622 203 636
rect 135 590 149 622
rect 181 590 203 622
rect 135 580 203 590
rect 27 566 95 580
rect 27 534 41 566
rect 73 534 95 566
rect 27 498 95 534
rect 27 466 41 498
rect 73 466 95 498
rect 27 412 95 466
rect 121 550 203 580
rect 121 518 149 550
rect 181 518 203 550
rect 121 412 203 518
rect 229 622 305 636
rect 229 590 251 622
rect 283 590 305 622
rect 229 550 305 590
rect 229 518 251 550
rect 283 518 305 550
rect 229 412 305 518
rect 331 622 399 636
rect 331 590 353 622
rect 385 590 399 622
rect 331 412 399 590
<< ndiffc >>
rect 41 194 73 226
rect 149 142 181 174
rect 375 220 407 252
rect 375 132 407 164
<< pdiffc >>
rect 149 590 181 622
rect 41 534 73 566
rect 41 466 73 498
rect 149 518 181 550
rect 251 590 283 622
rect 251 518 283 550
rect 353 590 385 622
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 203 636 229 672
rect 305 636 331 672
rect 95 580 121 616
rect 95 370 121 412
rect 61 352 121 370
rect 203 366 229 412
rect 305 366 331 412
rect 61 320 75 352
rect 107 320 121 352
rect 61 304 121 320
rect 181 352 241 366
rect 181 320 195 352
rect 227 320 241 352
rect 181 304 241 320
rect 305 352 387 366
rect 305 320 319 352
rect 351 320 387 352
rect 305 304 387 320
rect 95 266 121 304
rect 203 266 229 304
rect 305 266 331 304
rect 95 120 121 156
rect 203 82 229 118
rect 305 82 331 118
<< polycont >>
rect 75 320 107 352
rect 195 320 227 352
rect 319 320 351 352
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 139 622 191 712
rect 139 590 149 622
rect 181 590 191 622
rect 31 566 83 576
rect 31 534 41 566
rect 73 534 83 566
rect 31 498 83 534
rect 139 550 191 590
rect 139 518 149 550
rect 181 518 191 550
rect 139 508 191 518
rect 241 622 293 632
rect 241 590 251 622
rect 283 590 293 622
rect 241 550 293 590
rect 343 622 395 712
rect 343 590 353 622
rect 385 590 395 622
rect 343 580 395 590
rect 241 518 251 550
rect 283 540 293 550
rect 283 518 432 540
rect 241 508 432 518
rect 31 466 41 498
rect 73 471 83 498
rect 73 466 309 471
rect 31 434 309 466
rect 39 352 120 367
rect 39 320 75 352
rect 107 320 120 352
rect 39 306 120 320
rect 168 352 241 367
rect 168 320 195 352
rect 227 320 241 352
rect 168 306 241 320
rect 277 366 309 434
rect 277 352 361 366
rect 277 320 319 352
rect 351 320 361 352
rect 277 304 361 320
rect 277 270 309 304
rect 31 238 309 270
rect 400 263 432 508
rect 349 252 432 263
rect 31 226 83 238
rect 31 194 41 226
rect 73 194 83 226
rect 31 184 83 194
rect 349 220 375 252
rect 407 220 432 252
rect 138 174 192 188
rect 138 142 149 174
rect 181 142 192 174
rect 138 44 192 142
rect 349 164 432 220
rect 349 132 375 164
rect 407 132 432 164
rect 349 122 432 132
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 59 306 120 367 0 FreeSans 400 0 0 0 A_N
port 3 nsew
flabel metal1 s 349 122 432 263 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 168 306 241 367 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 186618
string GDS_FILE 6_final.gds
string GDS_START 182290
<< end >>
