magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754861848
<< nwell >>
rect -48 350 1296 834
<< pwell >>
rect 1 56 1236 292
rect -26 -56 1274 56
<< nmos >>
rect 96 118 122 266
rect 198 118 224 266
rect 300 118 326 266
rect 402 118 428 266
rect 504 118 530 266
rect 606 118 632 266
rect 708 118 734 266
rect 810 118 836 266
rect 912 118 938 266
rect 1014 118 1040 266
rect 1116 118 1142 266
<< pmos >>
rect 96 412 122 636
rect 198 412 224 636
rect 300 412 326 636
rect 402 412 428 636
rect 504 412 530 636
rect 606 412 632 636
rect 708 412 734 636
rect 810 412 836 636
rect 912 412 938 636
rect 1014 412 1040 636
rect 1116 412 1142 636
<< ndiff >>
rect 27 232 96 266
rect 27 200 42 232
rect 74 200 96 232
rect 27 164 96 200
rect 27 132 42 164
rect 74 132 96 164
rect 27 118 96 132
rect 122 164 198 266
rect 122 132 144 164
rect 176 132 198 164
rect 122 118 198 132
rect 224 232 300 266
rect 224 200 246 232
rect 278 200 300 232
rect 224 164 300 200
rect 224 132 246 164
rect 278 132 300 164
rect 224 118 300 132
rect 326 164 402 266
rect 326 132 348 164
rect 380 132 402 164
rect 326 118 402 132
rect 428 232 504 266
rect 428 200 450 232
rect 482 200 504 232
rect 428 164 504 200
rect 428 132 450 164
rect 482 132 504 164
rect 428 118 504 132
rect 530 164 606 266
rect 530 132 552 164
rect 584 132 606 164
rect 530 118 606 132
rect 632 232 708 266
rect 632 200 654 232
rect 686 200 708 232
rect 632 164 708 200
rect 632 132 654 164
rect 686 132 708 164
rect 632 118 708 132
rect 734 164 810 266
rect 734 132 756 164
rect 788 132 810 164
rect 734 118 810 132
rect 836 232 912 266
rect 836 200 858 232
rect 890 200 912 232
rect 836 164 912 200
rect 836 132 858 164
rect 890 132 912 164
rect 836 118 912 132
rect 938 164 1014 266
rect 938 132 960 164
rect 992 132 1014 164
rect 938 118 1014 132
rect 1040 232 1116 266
rect 1040 200 1062 232
rect 1094 200 1116 232
rect 1040 164 1116 200
rect 1040 132 1062 164
rect 1094 132 1116 164
rect 1040 118 1116 132
rect 1142 232 1210 266
rect 1142 200 1164 232
rect 1196 200 1210 232
rect 1142 164 1210 200
rect 1142 132 1164 164
rect 1196 132 1210 164
rect 1142 118 1210 132
<< pdiff >>
rect 28 622 96 636
rect 28 590 42 622
rect 74 590 96 622
rect 28 554 96 590
rect 28 522 42 554
rect 74 522 96 554
rect 28 486 96 522
rect 28 454 42 486
rect 74 454 96 486
rect 28 412 96 454
rect 122 622 198 636
rect 122 590 144 622
rect 176 590 198 622
rect 122 554 198 590
rect 122 522 144 554
rect 176 522 198 554
rect 122 412 198 522
rect 224 622 300 636
rect 224 590 246 622
rect 278 590 300 622
rect 224 554 300 590
rect 224 522 246 554
rect 278 522 300 554
rect 224 486 300 522
rect 224 454 246 486
rect 278 454 300 486
rect 224 412 300 454
rect 326 622 402 636
rect 326 590 348 622
rect 380 590 402 622
rect 326 554 402 590
rect 326 522 348 554
rect 380 522 402 554
rect 326 412 402 522
rect 428 622 504 636
rect 428 590 450 622
rect 482 590 504 622
rect 428 554 504 590
rect 428 522 450 554
rect 482 522 504 554
rect 428 486 504 522
rect 428 454 450 486
rect 482 454 504 486
rect 428 412 504 454
rect 530 622 606 636
rect 530 590 552 622
rect 584 590 606 622
rect 530 554 606 590
rect 530 522 552 554
rect 584 522 606 554
rect 530 412 606 522
rect 632 622 708 636
rect 632 590 654 622
rect 686 590 708 622
rect 632 554 708 590
rect 632 522 654 554
rect 686 522 708 554
rect 632 486 708 522
rect 632 454 654 486
rect 686 454 708 486
rect 632 412 708 454
rect 734 622 810 636
rect 734 590 756 622
rect 788 590 810 622
rect 734 554 810 590
rect 734 522 756 554
rect 788 522 810 554
rect 734 412 810 522
rect 836 622 912 636
rect 836 590 858 622
rect 890 590 912 622
rect 836 554 912 590
rect 836 522 858 554
rect 890 522 912 554
rect 836 486 912 522
rect 836 454 858 486
rect 890 454 912 486
rect 836 412 912 454
rect 938 622 1014 636
rect 938 590 960 622
rect 992 590 1014 622
rect 938 554 1014 590
rect 938 522 960 554
rect 992 522 1014 554
rect 938 412 1014 522
rect 1040 622 1116 636
rect 1040 590 1062 622
rect 1094 590 1116 622
rect 1040 554 1116 590
rect 1040 522 1062 554
rect 1094 522 1116 554
rect 1040 486 1116 522
rect 1040 454 1062 486
rect 1094 454 1116 486
rect 1040 412 1116 454
rect 1142 622 1211 636
rect 1142 590 1164 622
rect 1196 590 1211 622
rect 1142 554 1211 590
rect 1142 522 1164 554
rect 1196 522 1211 554
rect 1142 486 1211 522
rect 1142 454 1164 486
rect 1196 454 1211 486
rect 1142 412 1211 454
<< ndiffc >>
rect 42 200 74 232
rect 42 132 74 164
rect 144 132 176 164
rect 246 200 278 232
rect 246 132 278 164
rect 348 132 380 164
rect 450 200 482 232
rect 450 132 482 164
rect 552 132 584 164
rect 654 200 686 232
rect 654 132 686 164
rect 756 132 788 164
rect 858 200 890 232
rect 858 132 890 164
rect 960 132 992 164
rect 1062 200 1094 232
rect 1062 132 1094 164
rect 1164 200 1196 232
rect 1164 132 1196 164
<< pdiffc >>
rect 42 590 74 622
rect 42 522 74 554
rect 42 454 74 486
rect 144 590 176 622
rect 144 522 176 554
rect 246 590 278 622
rect 246 522 278 554
rect 246 454 278 486
rect 348 590 380 622
rect 348 522 380 554
rect 450 590 482 622
rect 450 522 482 554
rect 450 454 482 486
rect 552 590 584 622
rect 552 522 584 554
rect 654 590 686 622
rect 654 522 686 554
rect 654 454 686 486
rect 756 590 788 622
rect 756 522 788 554
rect 858 590 890 622
rect 858 522 890 554
rect 858 454 890 486
rect 960 590 992 622
rect 960 522 992 554
rect 1062 590 1094 622
rect 1062 522 1094 554
rect 1062 454 1094 486
rect 1164 590 1196 622
rect 1164 522 1196 554
rect 1164 454 1196 486
<< psubdiff >>
rect 0 16 1248 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1248 16
rect 0 -30 1248 -16
<< nsubdiff >>
rect 0 772 1248 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1248 772
rect 0 726 1248 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
<< poly >>
rect 96 636 122 672
rect 198 636 224 672
rect 300 636 326 672
rect 402 636 428 672
rect 504 636 530 672
rect 606 636 632 672
rect 708 636 734 672
rect 810 636 836 672
rect 912 636 938 672
rect 1014 636 1040 672
rect 1116 636 1142 672
rect 96 380 122 412
rect 198 380 224 412
rect 300 380 326 412
rect 96 363 326 380
rect 402 370 428 412
rect 504 370 530 412
rect 606 370 632 412
rect 708 370 734 412
rect 810 370 836 412
rect 912 370 938 412
rect 1014 370 1040 412
rect 1116 370 1142 412
rect 96 331 124 363
rect 156 331 192 363
rect 224 331 260 363
rect 292 331 326 363
rect 96 314 326 331
rect 96 266 122 314
rect 198 266 224 314
rect 300 266 326 314
rect 385 353 1142 370
rect 385 321 402 353
rect 434 321 470 353
rect 502 321 538 353
rect 570 321 606 353
rect 638 321 674 353
rect 706 321 742 353
rect 774 321 810 353
rect 842 321 878 353
rect 910 321 946 353
rect 978 321 1142 353
rect 385 304 1142 321
rect 385 298 428 304
rect 402 266 428 298
rect 504 266 530 304
rect 606 266 632 304
rect 708 266 734 304
rect 810 266 836 304
rect 912 266 938 304
rect 1014 266 1040 304
rect 1116 266 1142 304
rect 96 82 122 118
rect 198 82 224 118
rect 300 82 326 118
rect 402 82 428 118
rect 504 82 530 118
rect 606 82 632 118
rect 708 82 734 118
rect 810 82 836 118
rect 912 82 938 118
rect 1014 82 1040 118
rect 1116 82 1142 118
<< polycont >>
rect 124 331 156 363
rect 192 331 224 363
rect 260 331 292 363
rect 402 321 434 353
rect 470 321 502 353
rect 538 321 570 353
rect 606 321 638 353
rect 674 321 706 353
rect 742 321 774 353
rect 810 321 842 353
rect 878 321 910 353
rect 946 321 978 353
<< metal1 >>
rect 0 772 1248 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1248 772
rect 0 712 1248 740
rect 32 622 84 632
rect 32 590 42 622
rect 74 590 84 622
rect 32 554 84 590
rect 32 522 42 554
rect 74 522 84 554
rect 32 486 84 522
rect 134 622 186 712
rect 134 590 144 622
rect 176 590 186 622
rect 134 554 186 590
rect 134 522 144 554
rect 176 522 186 554
rect 134 512 186 522
rect 236 622 288 632
rect 236 590 246 622
rect 278 590 288 622
rect 236 554 288 590
rect 236 522 246 554
rect 278 522 288 554
rect 32 454 42 486
rect 74 476 84 486
rect 236 486 288 522
rect 338 622 390 712
rect 338 590 348 622
rect 380 590 390 622
rect 338 554 390 590
rect 338 522 348 554
rect 380 522 390 554
rect 338 512 390 522
rect 440 622 492 632
rect 440 590 450 622
rect 482 590 492 622
rect 440 554 492 590
rect 440 522 450 554
rect 482 522 492 554
rect 236 476 246 486
rect 74 454 246 476
rect 278 476 288 486
rect 440 486 492 522
rect 542 622 594 712
rect 542 590 552 622
rect 584 590 594 622
rect 542 554 594 590
rect 542 522 552 554
rect 584 522 594 554
rect 542 512 594 522
rect 644 622 696 632
rect 644 590 654 622
rect 686 590 696 622
rect 644 554 696 590
rect 644 522 654 554
rect 686 522 696 554
rect 278 454 388 476
rect 32 444 388 454
rect 440 454 450 486
rect 482 476 492 486
rect 644 486 696 522
rect 746 622 798 712
rect 746 590 756 622
rect 788 590 798 622
rect 746 554 798 590
rect 746 522 756 554
rect 788 522 798 554
rect 746 512 798 522
rect 848 622 900 632
rect 848 590 858 622
rect 890 590 900 622
rect 848 554 900 590
rect 848 522 858 554
rect 890 522 900 554
rect 644 476 654 486
rect 482 454 654 476
rect 686 476 696 486
rect 848 486 900 522
rect 950 622 1002 712
rect 950 590 960 622
rect 992 590 1002 622
rect 950 554 1002 590
rect 950 522 960 554
rect 992 522 1002 554
rect 950 512 1002 522
rect 1052 622 1104 632
rect 1052 590 1062 622
rect 1094 590 1104 622
rect 1052 554 1104 590
rect 1052 522 1062 554
rect 1094 522 1104 554
rect 848 476 858 486
rect 686 454 858 476
rect 890 476 900 486
rect 1052 486 1104 522
rect 1052 476 1062 486
rect 890 454 1062 476
rect 1094 454 1104 486
rect 440 444 1104 454
rect 1154 622 1206 712
rect 1154 590 1164 622
rect 1196 590 1206 622
rect 1154 554 1206 590
rect 1154 522 1164 554
rect 1196 522 1206 554
rect 1154 486 1206 522
rect 1154 454 1164 486
rect 1196 454 1206 486
rect 1154 444 1206 454
rect 114 363 302 373
rect 114 331 124 363
rect 156 331 192 363
rect 224 331 260 363
rect 292 331 302 363
rect 114 300 302 331
rect 354 363 388 444
rect 1052 363 1104 444
rect 354 353 995 363
rect 354 321 402 353
rect 434 321 470 353
rect 502 321 538 353
rect 570 321 606 353
rect 638 321 674 353
rect 706 321 742 353
rect 774 321 810 353
rect 842 321 878 353
rect 910 321 946 353
rect 978 321 995 353
rect 354 311 995 321
rect 354 242 388 311
rect 1052 310 1190 363
rect 1052 242 1104 310
rect 32 232 388 242
rect 32 200 42 232
rect 74 210 246 232
rect 74 200 84 210
rect 32 164 84 200
rect 236 200 246 210
rect 278 210 388 232
rect 440 232 1104 242
rect 278 200 288 210
rect 32 132 42 164
rect 74 132 84 164
rect 32 122 84 132
rect 134 164 186 174
rect 134 132 144 164
rect 176 132 186 164
rect 134 44 186 132
rect 236 164 288 200
rect 440 200 450 232
rect 482 210 654 232
rect 482 200 492 210
rect 236 132 246 164
rect 278 132 288 164
rect 236 122 288 132
rect 338 164 390 174
rect 338 132 348 164
rect 380 132 390 164
rect 338 44 390 132
rect 440 164 492 200
rect 644 200 654 210
rect 686 210 858 232
rect 686 200 696 210
rect 440 132 450 164
rect 482 132 492 164
rect 440 122 492 132
rect 542 164 594 174
rect 542 132 552 164
rect 584 132 594 164
rect 542 44 594 132
rect 644 164 696 200
rect 848 200 858 210
rect 890 210 1062 232
rect 890 200 900 210
rect 644 132 654 164
rect 686 132 696 164
rect 644 122 696 132
rect 746 164 798 174
rect 746 132 756 164
rect 788 132 798 164
rect 746 44 798 132
rect 848 164 900 200
rect 1052 200 1062 210
rect 1094 200 1104 232
rect 848 132 858 164
rect 890 132 900 164
rect 848 122 900 132
rect 950 164 1002 174
rect 950 132 960 164
rect 992 132 1002 164
rect 950 44 1002 132
rect 1052 164 1104 200
rect 1052 132 1062 164
rect 1094 132 1104 164
rect 1052 122 1104 132
rect 1154 232 1206 242
rect 1154 200 1164 232
rect 1196 200 1206 232
rect 1154 164 1206 200
rect 1154 132 1164 164
rect 1196 132 1206 164
rect 1154 44 1206 132
rect 0 16 1248 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1248 16
rect 0 -44 1248 -16
<< labels >>
flabel metal1 s 1104 310 1190 363 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 712 1248 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 114 300 302 373 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 -44 1248 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 756
string GDS_END 121754
string GDS_FILE 6_final.gds
string GDS_START 111554
<< end >>
